/* Verilog module written by vlog2Verilog (qflow) */

module ALU_wrapper(
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    output Done_o,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input clk,
    input reset
);

wire VDD = 1'b1;
wire GND = 1'b0;

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire BI_0_bF$buf0 ;
wire BI_0_bF$buf1 ;
wire BI_0_bF$buf2 ;
wire BI_0_bF$buf3 ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire [2:0] _926_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _923_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire ABCmd_i_2_bF$buf0 ;
wire ABCmd_i_2_bF$buf1 ;
wire ABCmd_i_2_bF$buf2 ;
wire ABCmd_i_2_bF$buf3 ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _878_ ;
wire _458_ ;
wire _32__bF$buf0 ;
wire _32__bF$buf1 ;
wire _32__bF$buf2 ;
wire _32__bF$buf3 ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire Done_o ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire BI_4_bF$buf0 ;
wire BI_4_bF$buf1 ;
wire BI_4_bF$buf2 ;
wire BI_4_bF$buf3 ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire _919_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _898_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _895_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _913_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _723__bF$buf0 ;
wire _723__bF$buf1 ;
wire _723__bF$buf2 ;
wire _723__bF$buf3 ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _904_ ;
wire _713_ ;
wire [7:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire BI_1_bF$buf0 ;
wire BI_1_bF$buf1 ;
wire BI_1_bF$buf2 ;
wire BI_1_bF$buf3 ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [2:0] state ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire [7:0] _924_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire BI_3_bF$buf0 ;
wire BI_3_bF$buf1 ;
wire BI_3_bF$buf2 ;
wire BI_3_bF$buf3 ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _897_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _912_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert32 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf0)
);

BUFX2 BUFX2_insert31 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf1)
);

BUFX2 BUFX2_insert30 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf2)
);

BUFX2 BUFX2_insert29 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf3)
);

BUFX2 BUFX2_insert28 (
    .A(BI[1]),
    .Y(BI_1_bF$buf0)
);

BUFX2 BUFX2_insert27 (
    .A(BI[1]),
    .Y(BI_1_bF$buf1)
);

BUFX2 BUFX2_insert26 (
    .A(BI[1]),
    .Y(BI_1_bF$buf2)
);

BUFX2 BUFX2_insert25 (
    .A(BI[1]),
    .Y(BI_1_bF$buf3)
);

BUFX2 BUFX2_insert24 (
    .A(BI[4]),
    .Y(BI_4_bF$buf0)
);

BUFX2 BUFX2_insert23 (
    .A(BI[4]),
    .Y(BI_4_bF$buf1)
);

BUFX2 BUFX2_insert22 (
    .A(BI[4]),
    .Y(BI_4_bF$buf2)
);

BUFX2 BUFX2_insert21 (
    .A(BI[4]),
    .Y(BI_4_bF$buf3)
);

BUFX2 BUFX2_insert20 (
    .A(_32_),
    .Y(_32__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .A(_32_),
    .Y(_32__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .A(_32_),
    .Y(_32__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .A(_32_),
    .Y(_32__bF$buf3)
);

CLKBUF1 CLKBUF1_insert16 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert15 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf4)
);

BUFX2 BUFX2_insert11 (
    .A(_723_),
    .Y(_723__bF$buf0)
);

BUFX2 BUFX2_insert10 (
    .A(_723_),
    .Y(_723__bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .A(_723_),
    .Y(_723__bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .A(_723_),
    .Y(_723__bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .A(BI[0]),
    .Y(BI_0_bF$buf0)
);

BUFX2 BUFX2_insert6 (
    .A(BI[0]),
    .Y(BI_0_bF$buf1)
);

BUFX2 BUFX2_insert5 (
    .A(BI[0]),
    .Y(BI_0_bF$buf2)
);

BUFX2 BUFX2_insert4 (
    .A(BI[0]),
    .Y(BI_0_bF$buf3)
);

BUFX2 BUFX2_insert3 (
    .A(BI[3]),
    .Y(BI_3_bF$buf0)
);

BUFX2 BUFX2_insert2 (
    .A(BI[3]),
    .Y(BI_3_bF$buf1)
);

BUFX2 BUFX2_insert1 (
    .A(BI[3]),
    .Y(BI_3_bF$buf2)
);

BUFX2 BUFX2_insert0 (
    .A(BI[3]),
    .Y(BI_3_bF$buf3)
);

NAND2X1 _1000_ (
    .A(BI[2]),
    .B(AI[2]),
    .Y(_68_)
);

INVX1 _1001_ (
    .A(_68_),
    .Y(_69_)
);

NAND2X1 _1002_ (
    .A(BI_1_bF$buf3),
    .B(AI[4]),
    .Y(_70_)
);

OR2X2 _1003_ (
    .A(_63_),
    .B(_70_),
    .Y(_71_)
);

AOI22X1 _1004_ (
    .A(BI_0_bF$buf3),
    .B(AI[4]),
    .C(BI_1_bF$buf2),
    .D(AI[3]),
    .Y(_72_)
);

INVX1 _1005_ (
    .A(_72_),
    .Y(_73_)
);

NAND3X1 _1006_ (
    .A(_73_),
    .B(_69_),
    .C(_71_),
    .Y(_74_)
);

NOR2X1 _1007_ (
    .A(_63_),
    .B(_70_),
    .Y(_75_)
);

OAI21X1 _1008_ (
    .A(_72_),
    .B(_75_),
    .C(_68_),
    .Y(_76_)
);

NAND3X1 _1009_ (
    .A(_76_),
    .B(_67_),
    .C(_74_),
    .Y(_77_)
);

INVX1 _1010_ (
    .A(_59_),
    .Y(_78_)
);

NAND2X1 _1011_ (
    .A(BI_4_bF$buf3),
    .B(AI[1]),
    .Y(_79_)
);

INVX2 _1012_ (
    .A(BI_4_bF$buf2),
    .Y(_80_)
);

NAND2X1 _1013_ (
    .A(BI_3_bF$buf3),
    .B(AI[1]),
    .Y(_81_)
);

OAI21X1 _1014_ (
    .A(_57_),
    .B(_80_),
    .C(_81_),
    .Y(_82_)
);

OAI21X1 _1015_ (
    .A(_79_),
    .B(_78_),
    .C(_82_),
    .Y(_83_)
);

AOI21X1 _1016_ (
    .A(_74_),
    .B(_76_),
    .C(_67_),
    .Y(_84_)
);

OAI21X1 _1017_ (
    .A(_83_),
    .B(_84_),
    .C(_77_),
    .Y(_85_)
);

OAI21X1 _1018_ (
    .A(_68_),
    .B(_72_),
    .C(_71_),
    .Y(_86_)
);

AND2X2 _1019_ (
    .A(BI_0_bF$buf2),
    .B(AI[5]),
    .Y(_87_)
);

NAND3X1 _1020_ (
    .A(BI_1_bF$buf1),
    .B(AI[4]),
    .C(_87_),
    .Y(_88_)
);

AOI22X1 _1021_ (
    .A(BI_0_bF$buf1),
    .B(AI[5]),
    .C(BI_1_bF$buf0),
    .D(AI[4]),
    .Y(_89_)
);

INVX1 _1022_ (
    .A(_89_),
    .Y(_90_)
);

NAND2X1 _1023_ (
    .A(BI[2]),
    .B(AI[3]),
    .Y(_91_)
);

INVX1 _1024_ (
    .A(_91_),
    .Y(_92_)
);

NAND3X1 _1025_ (
    .A(_90_),
    .B(_92_),
    .C(_88_),
    .Y(_93_)
);

NAND2X1 _1026_ (
    .A(BI_0_bF$buf0),
    .B(AI[5]),
    .Y(_94_)
);

NOR2X1 _1027_ (
    .A(_70_),
    .B(_94_),
    .Y(_95_)
);

OAI21X1 _1028_ (
    .A(_89_),
    .B(_95_),
    .C(_91_),
    .Y(_96_)
);

NAND3X1 _1029_ (
    .A(_93_),
    .B(_96_),
    .C(_86_),
    .Y(_97_)
);

AOI21X1 _1030_ (
    .A(_69_),
    .B(_73_),
    .C(_75_),
    .Y(_98_)
);

OAI21X1 _1031_ (
    .A(_89_),
    .B(_95_),
    .C(_92_),
    .Y(_99_)
);

NAND3X1 _1032_ (
    .A(_90_),
    .B(_91_),
    .C(_88_),
    .Y(_100_)
);

NAND3X1 _1033_ (
    .A(_100_),
    .B(_99_),
    .C(_98_),
    .Y(_101_)
);

NAND2X1 _1034_ (
    .A(AI[0]),
    .B(BI[5]),
    .Y(_102_)
);

INVX1 _1035_ (
    .A(_102_),
    .Y(_103_)
);

AND2X2 _1036_ (
    .A(BI_3_bF$buf2),
    .B(AI[2]),
    .Y(_104_)
);

NAND2X1 _1037_ (
    .A(_60_),
    .B(_104_),
    .Y(_105_)
);

INVX1 _1038_ (
    .A(AI[2]),
    .Y(_106_)
);

OAI21X1 _1039_ (
    .A(_58_),
    .B(_106_),
    .C(_79_),
    .Y(_107_)
);

NAND3X1 _1040_ (
    .A(_107_),
    .B(_103_),
    .C(_105_),
    .Y(_108_)
);

OAI21X1 _1041_ (
    .A(_58_),
    .B(_106_),
    .C(_60_),
    .Y(_109_)
);

INVX1 _1042_ (
    .A(AI[1]),
    .Y(_110_)
);

OAI21X1 _1043_ (
    .A(_80_),
    .B(_110_),
    .C(_104_),
    .Y(_111_)
);

NAND3X1 _1044_ (
    .A(_102_),
    .B(_109_),
    .C(_111_),
    .Y(_112_)
);

AND2X2 _1045_ (
    .A(_112_),
    .B(_108_),
    .Y(_113_)
);

NAND3X1 _1046_ (
    .A(_97_),
    .B(_101_),
    .C(_113_),
    .Y(_114_)
);

AOI21X1 _1047_ (
    .A(_99_),
    .B(_100_),
    .C(_98_),
    .Y(_115_)
);

AOI21X1 _1048_ (
    .A(_96_),
    .B(_93_),
    .C(_86_),
    .Y(_116_)
);

NAND2X1 _1049_ (
    .A(_108_),
    .B(_112_),
    .Y(_117_)
);

OAI21X1 _1050_ (
    .A(_115_),
    .B(_116_),
    .C(_117_),
    .Y(_118_)
);

NAND3X1 _1051_ (
    .A(_114_),
    .B(_118_),
    .C(_85_),
    .Y(_119_)
);

AOI21X1 _1052_ (
    .A(_118_),
    .B(_114_),
    .C(_85_),
    .Y(_120_)
);

OAI21X1 _1053_ (
    .A(_61_),
    .B(_120_),
    .C(_119_),
    .Y(_121_)
);

AOI21X1 _1054_ (
    .A(_101_),
    .B(_113_),
    .C(_115_),
    .Y(_122_)
);

OAI21X1 _1055_ (
    .A(_89_),
    .B(_91_),
    .C(_88_),
    .Y(_123_)
);

AND2X2 _1056_ (
    .A(BI_1_bF$buf3),
    .B(AI[6]),
    .Y(_124_)
);

NAND2X1 _1057_ (
    .A(_87_),
    .B(_124_),
    .Y(_125_)
);

INVX1 _1058_ (
    .A(BI_1_bF$buf2),
    .Y(_126_)
);

INVX2 _1059_ (
    .A(AI[5]),
    .Y(_127_)
);

NAND2X1 _1060_ (
    .A(BI_0_bF$buf3),
    .B(AI[6]),
    .Y(_128_)
);

OAI21X1 _1061_ (
    .A(_126_),
    .B(_127_),
    .C(_128_),
    .Y(_129_)
);

NAND2X1 _1062_ (
    .A(BI[2]),
    .B(AI[4]),
    .Y(_130_)
);

INVX1 _1063_ (
    .A(_130_),
    .Y(_131_)
);

NAND3X1 _1064_ (
    .A(_129_),
    .B(_131_),
    .C(_125_),
    .Y(_132_)
);

NAND2X1 _1065_ (
    .A(BI_1_bF$buf1),
    .B(AI[6]),
    .Y(_133_)
);

NOR2X1 _1066_ (
    .A(_94_),
    .B(_133_),
    .Y(_134_)
);

AOI22X1 _1067_ (
    .A(BI_0_bF$buf2),
    .B(AI[6]),
    .C(BI_1_bF$buf0),
    .D(AI[5]),
    .Y(_135_)
);

OAI21X1 _1068_ (
    .A(_135_),
    .B(_134_),
    .C(_130_),
    .Y(_136_)
);

AOI21X1 _1069_ (
    .A(_136_),
    .B(_132_),
    .C(_123_),
    .Y(_137_)
);

AOI21X1 _1070_ (
    .A(_90_),
    .B(_92_),
    .C(_95_),
    .Y(_138_)
);

OAI21X1 _1071_ (
    .A(_135_),
    .B(_134_),
    .C(_131_),
    .Y(_139_)
);

NAND3X1 _1072_ (
    .A(_129_),
    .B(_130_),
    .C(_125_),
    .Y(_140_)
);

AOI21X1 _1073_ (
    .A(_139_),
    .B(_140_),
    .C(_138_),
    .Y(_141_)
);

NAND2X1 _1074_ (
    .A(BI[5]),
    .B(AI[1]),
    .Y(_142_)
);

INVX1 _1075_ (
    .A(_142_),
    .Y(_143_)
);

AND2X2 _1076_ (
    .A(BI_4_bF$buf1),
    .B(AI[2]),
    .Y(_144_)
);

AND2X2 _1077_ (
    .A(BI_3_bF$buf1),
    .B(AI[3]),
    .Y(_145_)
);

NAND2X1 _1078_ (
    .A(_144_),
    .B(_145_),
    .Y(_146_)
);

INVX2 _1079_ (
    .A(AI[3]),
    .Y(_147_)
);

NAND2X1 _1080_ (
    .A(BI_4_bF$buf0),
    .B(AI[2]),
    .Y(_148_)
);

OAI21X1 _1081_ (
    .A(_58_),
    .B(_147_),
    .C(_148_),
    .Y(_149_)
);

NAND3X1 _1082_ (
    .A(_149_),
    .B(_143_),
    .C(_146_),
    .Y(_150_)
);

OAI21X1 _1083_ (
    .A(_58_),
    .B(_147_),
    .C(_144_),
    .Y(_151_)
);

OAI21X1 _1084_ (
    .A(_80_),
    .B(_106_),
    .C(_145_),
    .Y(_152_)
);

NAND3X1 _1085_ (
    .A(_142_),
    .B(_151_),
    .C(_152_),
    .Y(_153_)
);

AND2X2 _1086_ (
    .A(_153_),
    .B(_150_),
    .Y(_154_)
);

OAI21X1 _1087_ (
    .A(_137_),
    .B(_141_),
    .C(_154_),
    .Y(_155_)
);

NAND3X1 _1088_ (
    .A(_140_),
    .B(_139_),
    .C(_138_),
    .Y(_156_)
);

NAND3X1 _1089_ (
    .A(_123_),
    .B(_132_),
    .C(_136_),
    .Y(_157_)
);

NAND2X1 _1090_ (
    .A(_150_),
    .B(_153_),
    .Y(_158_)
);

NAND3X1 _1091_ (
    .A(_158_),
    .B(_157_),
    .C(_156_),
    .Y(_159_)
);

NAND3X1 _1092_ (
    .A(_159_),
    .B(_122_),
    .C(_155_),
    .Y(_160_)
);

OAI21X1 _1093_ (
    .A(_117_),
    .B(_116_),
    .C(_97_),
    .Y(_161_)
);

NAND3X1 _1094_ (
    .A(_157_),
    .B(_156_),
    .C(_154_),
    .Y(_162_)
);

OAI21X1 _1095_ (
    .A(_137_),
    .B(_141_),
    .C(_158_),
    .Y(_163_)
);

NAND3X1 _1096_ (
    .A(_162_),
    .B(_163_),
    .C(_161_),
    .Y(_164_)
);

INVX4 _1097_ (
    .A(BI[6]),
    .Y(_165_)
);

NOR2X1 _1098_ (
    .A(_57_),
    .B(_165_),
    .Y(_166_)
);

OAI21X1 _1099_ (
    .A(_81_),
    .B(_148_),
    .C(_108_),
    .Y(_167_)
);

NAND2X1 _1100_ (
    .A(_166_),
    .B(_167_),
    .Y(_168_)
);

OR2X2 _1101_ (
    .A(_167_),
    .B(_166_),
    .Y(_169_)
);

AND2X2 _1102_ (
    .A(_169_),
    .B(_168_),
    .Y(_170_)
);

NAND3X1 _1103_ (
    .A(_160_),
    .B(_164_),
    .C(_170_),
    .Y(_171_)
);

AOI21X1 _1104_ (
    .A(_163_),
    .B(_162_),
    .C(_161_),
    .Y(_172_)
);

AOI21X1 _1105_ (
    .A(_155_),
    .B(_159_),
    .C(_122_),
    .Y(_173_)
);

NAND2X1 _1106_ (
    .A(_168_),
    .B(_169_),
    .Y(_174_)
);

OAI21X1 _1107_ (
    .A(_173_),
    .B(_172_),
    .C(_174_),
    .Y(_175_)
);

NAND3X1 _1108_ (
    .A(_171_),
    .B(_175_),
    .C(_121_),
    .Y(_176_)
);

INVX1 _1109_ (
    .A(_168_),
    .Y(_177_)
);

OAI21X1 _1110_ (
    .A(_174_),
    .B(_172_),
    .C(_164_),
    .Y(_178_)
);

AOI21X1 _1111_ (
    .A(_156_),
    .B(_154_),
    .C(_141_),
    .Y(_179_)
);

OAI21X1 _1112_ (
    .A(_135_),
    .B(_130_),
    .C(_125_),
    .Y(_180_)
);

NAND3X1 _1113_ (
    .A(BI_0_bF$buf1),
    .B(\u_ALU8.AI7 ),
    .C(_124_),
    .Y(_181_)
);

AOI22X1 _1114_ (
    .A(BI_0_bF$buf0),
    .B(\u_ALU8.AI7 ),
    .C(BI_1_bF$buf3),
    .D(AI[6]),
    .Y(_182_)
);

INVX1 _1115_ (
    .A(_182_),
    .Y(_183_)
);

NAND2X1 _1116_ (
    .A(BI[2]),
    .B(AI[5]),
    .Y(_184_)
);

INVX1 _1117_ (
    .A(_184_),
    .Y(_185_)
);

NAND3X1 _1118_ (
    .A(_183_),
    .B(_185_),
    .C(_181_),
    .Y(_186_)
);

NAND2X1 _1119_ (
    .A(BI_1_bF$buf2),
    .B(\u_ALU8.AI7 ),
    .Y(_187_)
);

NOR2X1 _1120_ (
    .A(_128_),
    .B(_187_),
    .Y(_188_)
);

OAI21X1 _1121_ (
    .A(_182_),
    .B(_188_),
    .C(_184_),
    .Y(_189_)
);

AOI21X1 _1122_ (
    .A(_189_),
    .B(_186_),
    .C(_180_),
    .Y(_190_)
);

OAI21X1 _1123_ (
    .A(_182_),
    .B(_188_),
    .C(_185_),
    .Y(_191_)
);

NAND3X1 _1124_ (
    .A(_183_),
    .B(_184_),
    .C(_181_),
    .Y(_192_)
);

AOI22X1 _1125_ (
    .A(_125_),
    .B(_132_),
    .C(_191_),
    .D(_192_),
    .Y(_193_)
);

NAND2X1 _1126_ (
    .A(BI[5]),
    .B(AI[2]),
    .Y(_194_)
);

INVX1 _1127_ (
    .A(_194_),
    .Y(_195_)
);

AND2X2 _1128_ (
    .A(BI_4_bF$buf3),
    .B(AI[3]),
    .Y(_196_)
);

AND2X2 _1129_ (
    .A(BI_3_bF$buf0),
    .B(AI[4]),
    .Y(_197_)
);

NAND2X1 _1130_ (
    .A(_196_),
    .B(_197_),
    .Y(_198_)
);

AOI22X1 _1131_ (
    .A(BI_3_bF$buf3),
    .B(AI[4]),
    .C(BI_4_bF$buf2),
    .D(AI[3]),
    .Y(_199_)
);

INVX1 _1132_ (
    .A(_199_),
    .Y(_200_)
);

NAND3X1 _1133_ (
    .A(_195_),
    .B(_200_),
    .C(_198_),
    .Y(_201_)
);

INVX1 _1134_ (
    .A(AI[4]),
    .Y(_202_)
);

OAI21X1 _1135_ (
    .A(_58_),
    .B(_202_),
    .C(_196_),
    .Y(_203_)
);

OAI21X1 _1136_ (
    .A(_80_),
    .B(_147_),
    .C(_197_),
    .Y(_204_)
);

NAND3X1 _1137_ (
    .A(_194_),
    .B(_203_),
    .C(_204_),
    .Y(_205_)
);

AND2X2 _1138_ (
    .A(_205_),
    .B(_201_),
    .Y(_206_)
);

OAI21X1 _1139_ (
    .A(_193_),
    .B(_190_),
    .C(_206_),
    .Y(_207_)
);

AOI21X1 _1140_ (
    .A(_129_),
    .B(_131_),
    .C(_134_),
    .Y(_208_)
);

NAND3X1 _1141_ (
    .A(_192_),
    .B(_191_),
    .C(_208_),
    .Y(_209_)
);

NAND3X1 _1142_ (
    .A(_180_),
    .B(_186_),
    .C(_189_),
    .Y(_210_)
);

NAND2X1 _1143_ (
    .A(_201_),
    .B(_205_),
    .Y(_211_)
);

NAND3X1 _1144_ (
    .A(_211_),
    .B(_210_),
    .C(_209_),
    .Y(_212_)
);

NAND3X1 _1145_ (
    .A(_212_),
    .B(_207_),
    .C(_179_),
    .Y(_213_)
);

OAI21X1 _1146_ (
    .A(_158_),
    .B(_137_),
    .C(_157_),
    .Y(_214_)
);

NAND3X1 _1147_ (
    .A(_210_),
    .B(_209_),
    .C(_206_),
    .Y(_215_)
);

OAI21X1 _1148_ (
    .A(_193_),
    .B(_190_),
    .C(_211_),
    .Y(_216_)
);

NAND3X1 _1149_ (
    .A(_215_),
    .B(_214_),
    .C(_216_),
    .Y(_217_)
);

NAND2X1 _1150_ (
    .A(AI[0]),
    .B(BI[7]),
    .Y(_218_)
);

INVX1 _1151_ (
    .A(_218_),
    .Y(_219_)
);

AOI22X1 _1152_ (
    .A(_104_),
    .B(_196_),
    .C(_149_),
    .D(_143_),
    .Y(_220_)
);

INVX1 _1153_ (
    .A(_220_),
    .Y(_221_)
);

OAI21X1 _1154_ (
    .A(_165_),
    .B(_110_),
    .C(_221_),
    .Y(_222_)
);

NOR2X1 _1155_ (
    .A(_165_),
    .B(_110_),
    .Y(_223_)
);

NAND2X1 _1156_ (
    .A(_223_),
    .B(_220_),
    .Y(_224_)
);

NAND3X1 _1157_ (
    .A(_219_),
    .B(_224_),
    .C(_222_),
    .Y(_225_)
);

NAND2X1 _1158_ (
    .A(_223_),
    .B(_221_),
    .Y(_226_)
);

OAI21X1 _1159_ (
    .A(_165_),
    .B(_110_),
    .C(_220_),
    .Y(_227_)
);

NAND3X1 _1160_ (
    .A(_218_),
    .B(_227_),
    .C(_226_),
    .Y(_228_)
);

NAND2X1 _1161_ (
    .A(_228_),
    .B(_225_),
    .Y(_229_)
);

NAND3X1 _1162_ (
    .A(_229_),
    .B(_213_),
    .C(_217_),
    .Y(_230_)
);

AOI21X1 _1163_ (
    .A(_216_),
    .B(_215_),
    .C(_214_),
    .Y(_231_)
);

AOI21X1 _1164_ (
    .A(_207_),
    .B(_212_),
    .C(_179_),
    .Y(_232_)
);

NAND3X1 _1165_ (
    .A(_219_),
    .B(_227_),
    .C(_226_),
    .Y(_233_)
);

NAND3X1 _1166_ (
    .A(_218_),
    .B(_224_),
    .C(_222_),
    .Y(_234_)
);

NAND2X1 _1167_ (
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

OAI21X1 _1168_ (
    .A(_231_),
    .B(_232_),
    .C(_235_),
    .Y(_236_)
);

AOI21X1 _1169_ (
    .A(_236_),
    .B(_230_),
    .C(_178_),
    .Y(_237_)
);

AOI21X1 _1170_ (
    .A(_160_),
    .B(_170_),
    .C(_173_),
    .Y(_238_)
);

OAI21X1 _1171_ (
    .A(_231_),
    .B(_232_),
    .C(_229_),
    .Y(_239_)
);

NAND3X1 _1172_ (
    .A(_235_),
    .B(_213_),
    .C(_217_),
    .Y(_240_)
);

AOI21X1 _1173_ (
    .A(_239_),
    .B(_240_),
    .C(_238_),
    .Y(_241_)
);

OAI21X1 _1174_ (
    .A(_241_),
    .B(_237_),
    .C(_177_),
    .Y(_242_)
);

NAND3X1 _1175_ (
    .A(_240_),
    .B(_239_),
    .C(_238_),
    .Y(_243_)
);

NAND3X1 _1176_ (
    .A(_230_),
    .B(_236_),
    .C(_178_),
    .Y(_244_)
);

NAND3X1 _1177_ (
    .A(_168_),
    .B(_243_),
    .C(_244_),
    .Y(_245_)
);

AOI21X1 _1178_ (
    .A(_242_),
    .B(_245_),
    .C(_176_),
    .Y(_246_)
);

INVX1 _1179_ (
    .A(_246_),
    .Y(_247_)
);

INVX1 _1180_ (
    .A(_61_),
    .Y(_248_)
);

NOR2X1 _1181_ (
    .A(_62_),
    .B(_63_),
    .Y(_249_)
);

INVX1 _1182_ (
    .A(_65_),
    .Y(_250_)
);

INVX1 _1183_ (
    .A(BI_0_bF$buf3),
    .Y(_251_)
);

OAI21X1 _1184_ (
    .A(_251_),
    .B(_147_),
    .C(_62_),
    .Y(_252_)
);

AOI21X1 _1185_ (
    .A(_250_),
    .B(_252_),
    .C(_249_),
    .Y(_253_)
);

OAI21X1 _1186_ (
    .A(_72_),
    .B(_75_),
    .C(_69_),
    .Y(_254_)
);

NAND3X1 _1187_ (
    .A(_68_),
    .B(_73_),
    .C(_71_),
    .Y(_255_)
);

AOI21X1 _1188_ (
    .A(_255_),
    .B(_254_),
    .C(_253_),
    .Y(_256_)
);

AND2X2 _1189_ (
    .A(_61_),
    .B(_82_),
    .Y(_257_)
);

NAND3X1 _1190_ (
    .A(_254_),
    .B(_253_),
    .C(_255_),
    .Y(_258_)
);

AOI21X1 _1191_ (
    .A(_257_),
    .B(_258_),
    .C(_256_),
    .Y(_259_)
);

OAI21X1 _1192_ (
    .A(_115_),
    .B(_116_),
    .C(_113_),
    .Y(_260_)
);

NAND3X1 _1193_ (
    .A(_117_),
    .B(_97_),
    .C(_101_),
    .Y(_261_)
);

NAND3X1 _1194_ (
    .A(_261_),
    .B(_260_),
    .C(_259_),
    .Y(_262_)
);

NAND3X1 _1195_ (
    .A(_248_),
    .B(_262_),
    .C(_119_),
    .Y(_263_)
);

OAI21X1 _1196_ (
    .A(_173_),
    .B(_172_),
    .C(_170_),
    .Y(_264_)
);

NAND3X1 _1197_ (
    .A(_174_),
    .B(_160_),
    .C(_164_),
    .Y(_265_)
);

AOI22X1 _1198_ (
    .A(_119_),
    .B(_263_),
    .C(_264_),
    .D(_265_),
    .Y(_266_)
);

NAND3X1 _1199_ (
    .A(_177_),
    .B(_243_),
    .C(_244_),
    .Y(_267_)
);

OAI21X1 _1200_ (
    .A(_241_),
    .B(_237_),
    .C(_168_),
    .Y(_268_)
);

AOI21X1 _1201_ (
    .A(_268_),
    .B(_267_),
    .C(_266_),
    .Y(_269_)
);

NAND3X1 _1202_ (
    .A(_257_),
    .B(_258_),
    .C(_77_),
    .Y(_270_)
);

NAND3X1 _1203_ (
    .A(_252_),
    .B(_250_),
    .C(_64_),
    .Y(_271_)
);

NAND2X1 _1204_ (
    .A(BI_0_bF$buf2),
    .B(AI[1]),
    .Y(_272_)
);

NAND2X1 _1205_ (
    .A(AI[0]),
    .B(BI[2]),
    .Y(_273_)
);

AOI22X1 _1206_ (
    .A(BI_0_bF$buf1),
    .B(AI[2]),
    .C(BI_1_bF$buf1),
    .D(AI[1]),
    .Y(_274_)
);

OAI22X1 _1207_ (
    .A(_62_),
    .B(_272_),
    .C(_273_),
    .D(_274_),
    .Y(_275_)
);

OAI21X1 _1208_ (
    .A(_249_),
    .B(_66_),
    .C(_65_),
    .Y(_276_)
);

NAND3X1 _1209_ (
    .A(_275_),
    .B(_276_),
    .C(_271_),
    .Y(_277_)
);

AOI21X1 _1210_ (
    .A(_271_),
    .B(_276_),
    .C(_275_),
    .Y(_278_)
);

OAI21X1 _1211_ (
    .A(_78_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

OAI21X1 _1212_ (
    .A(_256_),
    .B(_84_),
    .C(_83_),
    .Y(_280_)
);

NAND3X1 _1213_ (
    .A(_270_),
    .B(_279_),
    .C(_280_),
    .Y(_281_)
);

INVX1 _1214_ (
    .A(_281_),
    .Y(_282_)
);

AOI22X1 _1215_ (
    .A(_77_),
    .B(_270_),
    .C(_260_),
    .D(_261_),
    .Y(_283_)
);

OAI21X1 _1216_ (
    .A(_283_),
    .B(_120_),
    .C(_61_),
    .Y(_284_)
);

NAND3X1 _1217_ (
    .A(_263_),
    .B(_282_),
    .C(_284_),
    .Y(_285_)
);

AOI21X1 _1218_ (
    .A(_175_),
    .B(_171_),
    .C(_121_),
    .Y(_286_)
);

NOR3X1 _1219_ (
    .A(_285_),
    .B(_266_),
    .C(_286_),
    .Y(_287_)
);

INVX1 _1220_ (
    .A(_278_),
    .Y(_288_)
);

NAND3X1 _1221_ (
    .A(_59_),
    .B(_277_),
    .C(_288_),
    .Y(_289_)
);

INVX1 _1222_ (
    .A(_273_),
    .Y(_290_)
);

NOR2X1 _1223_ (
    .A(_62_),
    .B(_272_),
    .Y(_291_)
);

NOR2X1 _1224_ (
    .A(_274_),
    .B(_291_),
    .Y(_292_)
);

NAND2X1 _1225_ (
    .A(_290_),
    .B(_292_),
    .Y(_293_)
);

NAND2X1 _1226_ (
    .A(AI[0]),
    .B(BI_1_bF$buf0),
    .Y(_294_)
);

NOR2X1 _1227_ (
    .A(_272_),
    .B(_294_),
    .Y(_295_)
);

OAI21X1 _1228_ (
    .A(_274_),
    .B(_291_),
    .C(_273_),
    .Y(_296_)
);

NAND3X1 _1229_ (
    .A(_295_),
    .B(_296_),
    .C(_293_),
    .Y(_297_)
);

INVX1 _1230_ (
    .A(_297_),
    .Y(_298_)
);

INVX1 _1231_ (
    .A(_277_),
    .Y(_299_)
);

OAI21X1 _1232_ (
    .A(_278_),
    .B(_299_),
    .C(_78_),
    .Y(_300_)
);

NAND3X1 _1233_ (
    .A(_298_),
    .B(_300_),
    .C(_289_),
    .Y(_301_)
);

AOI21X1 _1234_ (
    .A(_280_),
    .B(_270_),
    .C(_279_),
    .Y(_302_)
);

NOR3X1 _1235_ (
    .A(_302_),
    .B(_301_),
    .C(_282_),
    .Y(_303_)
);

OAI21X1 _1236_ (
    .A(_283_),
    .B(_120_),
    .C(_248_),
    .Y(_304_)
);

NAND3X1 _1237_ (
    .A(_61_),
    .B(_262_),
    .C(_119_),
    .Y(_305_)
);

NAND3X1 _1238_ (
    .A(_281_),
    .B(_305_),
    .C(_304_),
    .Y(_306_)
);

NAND3X1 _1239_ (
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_307_)
);

INVX1 _1240_ (
    .A(_307_),
    .Y(_308_)
);

OAI21X1 _1241_ (
    .A(_266_),
    .B(_286_),
    .C(_285_),
    .Y(_309_)
);

AOI21X1 _1242_ (
    .A(_308_),
    .B(_309_),
    .C(_287_),
    .Y(_310_)
);

OAI21X1 _1243_ (
    .A(_269_),
    .B(_310_),
    .C(_247_),
    .Y(_311_)
);

AOI21X1 _1244_ (
    .A(_177_),
    .B(_243_),
    .C(_241_),
    .Y(_312_)
);

NAND2X1 _1245_ (
    .A(_226_),
    .B(_233_),
    .Y(_313_)
);

OAI21X1 _1246_ (
    .A(_235_),
    .B(_231_),
    .C(_217_),
    .Y(_314_)
);

NAND2X1 _1247_ (
    .A(BI[7]),
    .B(AI[1]),
    .Y(_315_)
);

INVX1 _1248_ (
    .A(_315_),
    .Y(_316_)
);

NOR2X1 _1249_ (
    .A(_106_),
    .B(_165_),
    .Y(_317_)
);

OAI21X1 _1250_ (
    .A(_194_),
    .B(_199_),
    .C(_198_),
    .Y(_318_)
);

NAND2X1 _1251_ (
    .A(_317_),
    .B(_318_),
    .Y(_319_)
);

OR2X2 _1252_ (
    .A(_318_),
    .B(_317_),
    .Y(_320_)
);

NAND3X1 _1253_ (
    .A(_316_),
    .B(_319_),
    .C(_320_),
    .Y(_321_)
);

AND2X2 _1254_ (
    .A(_318_),
    .B(_317_),
    .Y(_322_)
);

NOR2X1 _1255_ (
    .A(_317_),
    .B(_318_),
    .Y(_323_)
);

OAI21X1 _1256_ (
    .A(_323_),
    .B(_322_),
    .C(_315_),
    .Y(_324_)
);

NAND2X1 _1257_ (
    .A(_324_),
    .B(_321_),
    .Y(_325_)
);

AOI21X1 _1258_ (
    .A(_206_),
    .B(_209_),
    .C(_193_),
    .Y(_326_)
);

NAND2X1 _1259_ (
    .A(BI[5]),
    .B(AI[3]),
    .Y(_327_)
);

AND2X2 _1260_ (
    .A(BI_4_bF$buf1),
    .B(AI[4]),
    .Y(_328_)
);

OAI21X1 _1261_ (
    .A(_127_),
    .B(_58_),
    .C(_328_),
    .Y(_329_)
);

AND2X2 _1262_ (
    .A(AI[5]),
    .B(BI_3_bF$buf2),
    .Y(_330_)
);

OAI21X1 _1263_ (
    .A(_80_),
    .B(_202_),
    .C(_330_),
    .Y(_331_)
);

NAND3X1 _1264_ (
    .A(_327_),
    .B(_329_),
    .C(_331_),
    .Y(_332_)
);

INVX1 _1265_ (
    .A(_327_),
    .Y(_333_)
);

NAND2X1 _1266_ (
    .A(_328_),
    .B(_330_),
    .Y(_334_)
);

AOI22X1 _1267_ (
    .A(AI[5]),
    .B(BI_3_bF$buf1),
    .C(BI_4_bF$buf0),
    .D(AI[4]),
    .Y(_335_)
);

INVX1 _1268_ (
    .A(_335_),
    .Y(_336_)
);

NAND3X1 _1269_ (
    .A(_333_),
    .B(_336_),
    .C(_334_),
    .Y(_337_)
);

NAND2X1 _1270_ (
    .A(_337_),
    .B(_332_),
    .Y(_338_)
);

AOI21X1 _1271_ (
    .A(_183_),
    .B(_185_),
    .C(_188_),
    .Y(_339_)
);

NAND2X1 _1272_ (
    .A(\u_ALU8.AI7 ),
    .B(BI[2]),
    .Y(_340_)
);

INVX1 _1273_ (
    .A(_340_),
    .Y(_341_)
);

AOI22X1 _1274_ (
    .A(BI_1_bF$buf3),
    .B(\u_ALU8.AI7 ),
    .C(BI[2]),
    .D(AI[6]),
    .Y(_342_)
);

AOI21X1 _1275_ (
    .A(_341_),
    .B(_124_),
    .C(_342_),
    .Y(_343_)
);

NAND2X1 _1276_ (
    .A(_343_),
    .B(_339_),
    .Y(_344_)
);

OAI21X1 _1277_ (
    .A(_182_),
    .B(_184_),
    .C(_181_),
    .Y(_345_)
);

INVX1 _1278_ (
    .A(_342_),
    .Y(_346_)
);

OAI21X1 _1279_ (
    .A(_133_),
    .B(_340_),
    .C(_346_),
    .Y(_347_)
);

NAND2X1 _1280_ (
    .A(_347_),
    .B(_345_),
    .Y(_348_)
);

NAND3X1 _1281_ (
    .A(_348_),
    .B(_338_),
    .C(_344_),
    .Y(_349_)
);

AND2X2 _1282_ (
    .A(_332_),
    .B(_337_),
    .Y(_350_)
);

NAND2X1 _1283_ (
    .A(_343_),
    .B(_345_),
    .Y(_351_)
);

NAND2X1 _1284_ (
    .A(_347_),
    .B(_339_),
    .Y(_352_)
);

NAND3X1 _1285_ (
    .A(_351_),
    .B(_352_),
    .C(_350_),
    .Y(_353_)
);

NAND3X1 _1286_ (
    .A(_349_),
    .B(_353_),
    .C(_326_),
    .Y(_354_)
);

OAI21X1 _1287_ (
    .A(_211_),
    .B(_190_),
    .C(_210_),
    .Y(_355_)
);

AOI22X1 _1288_ (
    .A(_332_),
    .B(_337_),
    .C(_352_),
    .D(_351_),
    .Y(_356_)
);

AOI21X1 _1289_ (
    .A(_344_),
    .B(_348_),
    .C(_338_),
    .Y(_357_)
);

OAI21X1 _1290_ (
    .A(_356_),
    .B(_357_),
    .C(_355_),
    .Y(_358_)
);

NAND3X1 _1291_ (
    .A(_325_),
    .B(_358_),
    .C(_354_),
    .Y(_359_)
);

AND2X2 _1292_ (
    .A(_321_),
    .B(_324_),
    .Y(_360_)
);

NAND3X1 _1293_ (
    .A(_349_),
    .B(_353_),
    .C(_355_),
    .Y(_361_)
);

OAI21X1 _1294_ (
    .A(_356_),
    .B(_357_),
    .C(_326_),
    .Y(_362_)
);

NAND3X1 _1295_ (
    .A(_362_),
    .B(_361_),
    .C(_360_),
    .Y(_363_)
);

NAND3X1 _1296_ (
    .A(_359_),
    .B(_363_),
    .C(_314_),
    .Y(_364_)
);

AOI21X1 _1297_ (
    .A(_213_),
    .B(_229_),
    .C(_232_),
    .Y(_365_)
);

AOI22X1 _1298_ (
    .A(_321_),
    .B(_324_),
    .C(_361_),
    .D(_362_),
    .Y(_366_)
);

AOI21X1 _1299_ (
    .A(_354_),
    .B(_358_),
    .C(_325_),
    .Y(_367_)
);

OAI21X1 _1300_ (
    .A(_366_),
    .B(_367_),
    .C(_365_),
    .Y(_368_)
);

AOI21X1 _1301_ (
    .A(_364_),
    .B(_368_),
    .C(_313_),
    .Y(_369_)
);

INVX1 _1302_ (
    .A(_313_),
    .Y(_370_)
);

NAND3X1 _1303_ (
    .A(_359_),
    .B(_363_),
    .C(_365_),
    .Y(_371_)
);

OAI21X1 _1304_ (
    .A(_366_),
    .B(_367_),
    .C(_314_),
    .Y(_372_)
);

AOI21X1 _1305_ (
    .A(_371_),
    .B(_372_),
    .C(_370_),
    .Y(_373_)
);

OAI21X1 _1306_ (
    .A(_369_),
    .B(_373_),
    .C(_312_),
    .Y(_374_)
);

OAI21X1 _1307_ (
    .A(_168_),
    .B(_237_),
    .C(_244_),
    .Y(_375_)
);

NAND3X1 _1308_ (
    .A(_370_),
    .B(_372_),
    .C(_371_),
    .Y(_376_)
);

NAND3X1 _1309_ (
    .A(_313_),
    .B(_368_),
    .C(_364_),
    .Y(_377_)
);

NAND3X1 _1310_ (
    .A(_376_),
    .B(_377_),
    .C(_375_),
    .Y(_378_)
);

AND2X2 _1311_ (
    .A(_374_),
    .B(_378_),
    .Y(_379_)
);

NAND2X1 _1312_ (
    .A(_379_),
    .B(_311_),
    .Y(_380_)
);

NAND3X1 _1313_ (
    .A(_176_),
    .B(_245_),
    .C(_242_),
    .Y(_381_)
);

INVX1 _1314_ (
    .A(_285_),
    .Y(_382_)
);

NAND2X1 _1315_ (
    .A(_171_),
    .B(_175_),
    .Y(_383_)
);

NAND3X1 _1316_ (
    .A(_119_),
    .B(_263_),
    .C(_383_),
    .Y(_384_)
);

NAND3X1 _1317_ (
    .A(_176_),
    .B(_382_),
    .C(_384_),
    .Y(_385_)
);

AOI21X1 _1318_ (
    .A(_384_),
    .B(_176_),
    .C(_382_),
    .Y(_386_)
);

OAI21X1 _1319_ (
    .A(_307_),
    .B(_386_),
    .C(_385_),
    .Y(_387_)
);

AOI21X1 _1320_ (
    .A(_387_),
    .B(_381_),
    .C(_246_),
    .Y(_388_)
);

NAND2X1 _1321_ (
    .A(_378_),
    .B(_374_),
    .Y(_389_)
);

NAND2X1 _1322_ (
    .A(_389_),
    .B(_388_),
    .Y(_390_)
);

AND2X2 _1323_ (
    .A(_390_),
    .B(_380_),
    .Y(_391_)
);

NOR2X1 _1324_ (
    .A(ABCmd_i[7]),
    .B(HC),
    .Y(_392_)
);

NOR2X1 _1325_ (
    .A(_392_),
    .B(_733_),
    .Y(_393_)
);

OAI21X1 _1326_ (
    .A(_54_),
    .B(_391_),
    .C(_393_),
    .Y(_394_)
);

AOI21X1 _1327_ (
    .A(BI_0_bF$buf0),
    .B(AI[0]),
    .C(_54_),
    .Y(_395_)
);

OAI21X1 _1328_ (
    .A(ACC[0]),
    .B(ABCmd_i[7]),
    .C(_733_),
    .Y(_396_)
);

OAI21X1 _1329_ (
    .A(_395_),
    .B(_396_),
    .C(_394_),
    .Y(_397_)
);

NAND2X1 _1330_ (
    .A(_718_),
    .B(_397_),
    .Y(_398_)
);

OAI21X1 _1331_ (
    .A(_56_),
    .B(_718_),
    .C(_398_),
    .Y(_9_)
);

INVX1 _1332_ (
    .A(_924_[1]),
    .Y(_399_)
);

INVX1 _1333_ (
    .A(AN),
    .Y(_400_)
);

OAI21X1 _1334_ (
    .A(state[1]),
    .B(_730_),
    .C(ABCmd_i[7]),
    .Y(_401_)
);

OAI21X1 _1335_ (
    .A(_400_),
    .B(_733_),
    .C(_401_),
    .Y(_402_)
);

AOI21X1 _1336_ (
    .A(_359_),
    .B(_363_),
    .C(_314_),
    .Y(_403_)
);

OAI21X1 _1337_ (
    .A(_370_),
    .B(_403_),
    .C(_364_),
    .Y(_404_)
);

OAI21X1 _1338_ (
    .A(_315_),
    .B(_323_),
    .C(_319_),
    .Y(_405_)
);

AOI21X1 _1339_ (
    .A(_349_),
    .B(_353_),
    .C(_355_),
    .Y(_406_)
);

OAI21X1 _1340_ (
    .A(_325_),
    .B(_406_),
    .C(_361_),
    .Y(_407_)
);

NAND2X1 _1341_ (
    .A(AI[2]),
    .B(BI[7]),
    .Y(_408_)
);

INVX1 _1342_ (
    .A(_408_),
    .Y(_409_)
);

NOR2X1 _1343_ (
    .A(_147_),
    .B(_165_),
    .Y(_410_)
);

OAI21X1 _1344_ (
    .A(_327_),
    .B(_335_),
    .C(_334_),
    .Y(_411_)
);

NAND2X1 _1345_ (
    .A(_410_),
    .B(_411_),
    .Y(_412_)
);

OR2X2 _1346_ (
    .A(_411_),
    .B(_410_),
    .Y(_413_)
);

NAND3X1 _1347_ (
    .A(_409_),
    .B(_412_),
    .C(_413_),
    .Y(_414_)
);

AND2X2 _1348_ (
    .A(_411_),
    .B(_410_),
    .Y(_415_)
);

NOR2X1 _1349_ (
    .A(_410_),
    .B(_411_),
    .Y(_416_)
);

OAI21X1 _1350_ (
    .A(_416_),
    .B(_415_),
    .C(_408_),
    .Y(_417_)
);

NAND2X1 _1351_ (
    .A(_417_),
    .B(_414_),
    .Y(_418_)
);

NOR2X1 _1352_ (
    .A(_347_),
    .B(_339_),
    .Y(_419_)
);

AOI21X1 _1353_ (
    .A(_350_),
    .B(_352_),
    .C(_419_),
    .Y(_420_)
);

NAND2X1 _1354_ (
    .A(AI[4]),
    .B(BI[5]),
    .Y(_421_)
);

INVX1 _1355_ (
    .A(_421_),
    .Y(_422_)
);

AND2X2 _1356_ (
    .A(AI[5]),
    .B(BI_4_bF$buf3),
    .Y(_423_)
);

AND2X2 _1357_ (
    .A(AI[6]),
    .B(BI_3_bF$buf0),
    .Y(_424_)
);

NAND2X1 _1358_ (
    .A(_423_),
    .B(_424_),
    .Y(_425_)
);

AOI22X1 _1359_ (
    .A(AI[6]),
    .B(BI_3_bF$buf3),
    .C(AI[5]),
    .D(BI_4_bF$buf2),
    .Y(_426_)
);

INVX1 _1360_ (
    .A(_426_),
    .Y(_427_)
);

AOI21X1 _1361_ (
    .A(_425_),
    .B(_427_),
    .C(_422_),
    .Y(_428_)
);

INVX2 _1362_ (
    .A(AI[6]),
    .Y(_429_)
);

OAI21X1 _1363_ (
    .A(_429_),
    .B(_58_),
    .C(_423_),
    .Y(_430_)
);

OAI21X1 _1364_ (
    .A(_127_),
    .B(_80_),
    .C(_424_),
    .Y(_431_)
);

AOI21X1 _1365_ (
    .A(_430_),
    .B(_431_),
    .C(_421_),
    .Y(_432_)
);

OAI22X1 _1366_ (
    .A(_124_),
    .B(_340_),
    .C(_428_),
    .D(_432_),
    .Y(_433_)
);

NAND3X1 _1367_ (
    .A(_421_),
    .B(_430_),
    .C(_431_),
    .Y(_434_)
);

NAND3X1 _1368_ (
    .A(_422_),
    .B(_427_),
    .C(_425_),
    .Y(_435_)
);

NOR2X1 _1369_ (
    .A(_340_),
    .B(_124_),
    .Y(_436_)
);

NAND3X1 _1370_ (
    .A(_436_),
    .B(_435_),
    .C(_434_),
    .Y(_437_)
);

NAND2X1 _1371_ (
    .A(_437_),
    .B(_433_),
    .Y(_438_)
);

NOR2X1 _1372_ (
    .A(_438_),
    .B(_420_),
    .Y(_439_)
);

NOR2X1 _1373_ (
    .A(_343_),
    .B(_345_),
    .Y(_440_)
);

OAI21X1 _1374_ (
    .A(_338_),
    .B(_440_),
    .C(_351_),
    .Y(_441_)
);

AOI21X1 _1375_ (
    .A(_433_),
    .B(_437_),
    .C(_441_),
    .Y(_442_)
);

OAI21X1 _1376_ (
    .A(_442_),
    .B(_439_),
    .C(_418_),
    .Y(_443_)
);

AND2X2 _1377_ (
    .A(_414_),
    .B(_417_),
    .Y(_444_)
);

NAND3X1 _1378_ (
    .A(_433_),
    .B(_437_),
    .C(_441_),
    .Y(_445_)
);

NAND2X1 _1379_ (
    .A(_438_),
    .B(_420_),
    .Y(_446_)
);

NAND3X1 _1380_ (
    .A(_445_),
    .B(_446_),
    .C(_444_),
    .Y(_447_)
);

NAND3X1 _1381_ (
    .A(_447_),
    .B(_443_),
    .C(_407_),
    .Y(_448_)
);

NOR3X1 _1382_ (
    .A(_356_),
    .B(_357_),
    .C(_326_),
    .Y(_449_)
);

AOI21X1 _1383_ (
    .A(_360_),
    .B(_362_),
    .C(_449_),
    .Y(_450_)
);

AOI21X1 _1384_ (
    .A(_446_),
    .B(_445_),
    .C(_444_),
    .Y(_451_)
);

NAND3X1 _1385_ (
    .A(_433_),
    .B(_437_),
    .C(_420_),
    .Y(_452_)
);

OAI21X1 _1386_ (
    .A(_419_),
    .B(_357_),
    .C(_438_),
    .Y(_453_)
);

AOI21X1 _1387_ (
    .A(_452_),
    .B(_453_),
    .C(_418_),
    .Y(_454_)
);

OAI21X1 _1388_ (
    .A(_451_),
    .B(_454_),
    .C(_450_),
    .Y(_455_)
);

NAND3X1 _1389_ (
    .A(_405_),
    .B(_448_),
    .C(_455_),
    .Y(_456_)
);

INVX1 _1390_ (
    .A(_405_),
    .Y(_457_)
);

NAND3X1 _1391_ (
    .A(_443_),
    .B(_447_),
    .C(_450_),
    .Y(_458_)
);

OAI21X1 _1392_ (
    .A(_454_),
    .B(_451_),
    .C(_407_),
    .Y(_459_)
);

NAND3X1 _1393_ (
    .A(_457_),
    .B(_459_),
    .C(_458_),
    .Y(_460_)
);

AOI21X1 _1394_ (
    .A(_456_),
    .B(_460_),
    .C(_404_),
    .Y(_461_)
);

NAND3X1 _1395_ (
    .A(_457_),
    .B(_448_),
    .C(_455_),
    .Y(_462_)
);

NAND3X1 _1396_ (
    .A(_405_),
    .B(_459_),
    .C(_458_),
    .Y(_463_)
);

AOI22X1 _1397_ (
    .A(_364_),
    .B(_377_),
    .C(_463_),
    .D(_462_),
    .Y(_464_)
);

NOR2X1 _1398_ (
    .A(_464_),
    .B(_461_),
    .Y(_465_)
);

AOI21X1 _1399_ (
    .A(_380_),
    .B(_378_),
    .C(_465_),
    .Y(_466_)
);

OAI21X1 _1400_ (
    .A(_389_),
    .B(_388_),
    .C(_378_),
    .Y(_467_)
);

INVX1 _1401_ (
    .A(_364_),
    .Y(_468_)
);

AOI21X1 _1402_ (
    .A(_313_),
    .B(_368_),
    .C(_468_),
    .Y(_469_)
);

NAND3X1 _1403_ (
    .A(_462_),
    .B(_463_),
    .C(_469_),
    .Y(_470_)
);

NAND3X1 _1404_ (
    .A(_456_),
    .B(_460_),
    .C(_404_),
    .Y(_471_)
);

NAND2X1 _1405_ (
    .A(_471_),
    .B(_470_),
    .Y(_472_)
);

OAI21X1 _1406_ (
    .A(_472_),
    .B(_467_),
    .C(ABCmd_i[7]),
    .Y(_473_)
);

OAI21X1 _1407_ (
    .A(_466_),
    .B(_473_),
    .C(_402_),
    .Y(_474_)
);

AND2X2 _1408_ (
    .A(_272_),
    .B(_294_),
    .Y(_475_)
);

NAND2X1 _1409_ (
    .A(ACC[1]),
    .B(_54_),
    .Y(_476_)
);

OAI21X1 _1410_ (
    .A(_272_),
    .B(_294_),
    .C(ABCmd_i[7]),
    .Y(_477_)
);

OAI21X1 _1411_ (
    .A(_477_),
    .B(_475_),
    .C(_476_),
    .Y(_478_)
);

AOI21X1 _1412_ (
    .A(_478_),
    .B(_721_),
    .C(_730_),
    .Y(_479_)
);

AOI22X1 _1413_ (
    .A(_399_),
    .B(_730_),
    .C(_474_),
    .D(_479_),
    .Y(_10_)
);

OAI21X1 _1414_ (
    .A(state[0]),
    .B(_717_),
    .C(_924_[2]),
    .Y(_480_)
);

NAND3X1 _1415_ (
    .A(_379_),
    .B(_465_),
    .C(_311_),
    .Y(_481_)
);

AOI21X1 _1416_ (
    .A(_378_),
    .B(_471_),
    .C(_461_),
    .Y(_482_)
);

INVX1 _1417_ (
    .A(_482_),
    .Y(_483_)
);

OAI21X1 _1418_ (
    .A(_408_),
    .B(_416_),
    .C(_412_),
    .Y(_484_)
);

INVX1 _1419_ (
    .A(_484_),
    .Y(_485_)
);

AOI21X1 _1420_ (
    .A(_444_),
    .B(_446_),
    .C(_439_),
    .Y(_486_)
);

NAND2X1 _1421_ (
    .A(AI[3]),
    .B(BI[7]),
    .Y(_487_)
);

INVX1 _1422_ (
    .A(_487_),
    .Y(_488_)
);

NOR2X1 _1423_ (
    .A(_202_),
    .B(_165_),
    .Y(_489_)
);

OAI21X1 _1424_ (
    .A(_421_),
    .B(_426_),
    .C(_425_),
    .Y(_490_)
);

NAND2X1 _1425_ (
    .A(_489_),
    .B(_490_),
    .Y(_491_)
);

OR2X2 _1426_ (
    .A(_490_),
    .B(_489_),
    .Y(_492_)
);

NAND3X1 _1427_ (
    .A(_488_),
    .B(_491_),
    .C(_492_),
    .Y(_493_)
);

AND2X2 _1428_ (
    .A(_490_),
    .B(_489_),
    .Y(_494_)
);

NOR2X1 _1429_ (
    .A(_489_),
    .B(_490_),
    .Y(_495_)
);

OAI21X1 _1430_ (
    .A(_495_),
    .B(_494_),
    .C(_487_),
    .Y(_496_)
);

NAND2X1 _1431_ (
    .A(_496_),
    .B(_493_),
    .Y(_497_)
);

NAND2X1 _1432_ (
    .A(_124_),
    .B(_341_),
    .Y(_498_)
);

NAND2X1 _1433_ (
    .A(AI[5]),
    .B(BI[5]),
    .Y(_499_)
);

INVX1 _1434_ (
    .A(_499_),
    .Y(_500_)
);

NAND2X1 _1435_ (
    .A(AI[6]),
    .B(BI_3_bF$buf2),
    .Y(_501_)
);

NAND2X1 _1436_ (
    .A(\u_ALU8.AI7 ),
    .B(BI_4_bF$buf1),
    .Y(_502_)
);

NOR2X1 _1437_ (
    .A(_501_),
    .B(_502_),
    .Y(_503_)
);

INVX1 _1438_ (
    .A(_503_),
    .Y(_504_)
);

AOI22X1 _1439_ (
    .A(\u_ALU8.AI7 ),
    .B(BI_3_bF$buf1),
    .C(AI[6]),
    .D(BI_4_bF$buf0),
    .Y(_505_)
);

INVX1 _1440_ (
    .A(_505_),
    .Y(_506_)
);

NAND3X1 _1441_ (
    .A(_500_),
    .B(_506_),
    .C(_504_),
    .Y(_507_)
);

OAI21X1 _1442_ (
    .A(_505_),
    .B(_503_),
    .C(_499_),
    .Y(_508_)
);

NAND2X1 _1443_ (
    .A(_508_),
    .B(_507_),
    .Y(_509_)
);

AOI21X1 _1444_ (
    .A(_498_),
    .B(_437_),
    .C(_509_),
    .Y(_510_)
);

NAND3X1 _1445_ (
    .A(_498_),
    .B(_437_),
    .C(_509_),
    .Y(_511_)
);

INVX1 _1446_ (
    .A(_511_),
    .Y(_512_)
);

OAI21X1 _1447_ (
    .A(_510_),
    .B(_512_),
    .C(_497_),
    .Y(_513_)
);

AND2X2 _1448_ (
    .A(_493_),
    .B(_496_),
    .Y(_514_)
);

NAND2X1 _1449_ (
    .A(_498_),
    .B(_437_),
    .Y(_515_)
);

NAND3X1 _1450_ (
    .A(_507_),
    .B(_508_),
    .C(_515_),
    .Y(_516_)
);

NAND3X1 _1451_ (
    .A(_516_),
    .B(_511_),
    .C(_514_),
    .Y(_517_)
);

NAND3X1 _1452_ (
    .A(_513_),
    .B(_517_),
    .C(_486_),
    .Y(_518_)
);

OAI21X1 _1453_ (
    .A(_418_),
    .B(_442_),
    .C(_445_),
    .Y(_519_)
);

AOI22X1 _1454_ (
    .A(_493_),
    .B(_496_),
    .C(_516_),
    .D(_511_),
    .Y(_520_)
);

OR2X2 _1455_ (
    .A(_515_),
    .B(_509_),
    .Y(_521_)
);

NAND2X1 _1456_ (
    .A(_509_),
    .B(_515_),
    .Y(_522_)
);

AOI21X1 _1457_ (
    .A(_521_),
    .B(_522_),
    .C(_497_),
    .Y(_523_)
);

OAI21X1 _1458_ (
    .A(_520_),
    .B(_523_),
    .C(_519_),
    .Y(_524_)
);

NAND3X1 _1459_ (
    .A(_485_),
    .B(_524_),
    .C(_518_),
    .Y(_525_)
);

NAND3X1 _1460_ (
    .A(_513_),
    .B(_517_),
    .C(_519_),
    .Y(_526_)
);

OAI21X1 _1461_ (
    .A(_520_),
    .B(_523_),
    .C(_486_),
    .Y(_527_)
);

NAND3X1 _1462_ (
    .A(_484_),
    .B(_526_),
    .C(_527_),
    .Y(_528_)
);

NAND2X1 _1463_ (
    .A(_528_),
    .B(_525_),
    .Y(_529_)
);

NAND3X1 _1464_ (
    .A(_448_),
    .B(_456_),
    .C(_529_),
    .Y(_530_)
);

AOI21X1 _1465_ (
    .A(_443_),
    .B(_447_),
    .C(_407_),
    .Y(_531_)
);

OAI21X1 _1466_ (
    .A(_457_),
    .B(_531_),
    .C(_448_),
    .Y(_532_)
);

NAND3X1 _1467_ (
    .A(_525_),
    .B(_528_),
    .C(_532_),
    .Y(_533_)
);

NAND2X1 _1468_ (
    .A(_533_),
    .B(_530_),
    .Y(_534_)
);

AOI21X1 _1469_ (
    .A(_481_),
    .B(_483_),
    .C(_534_),
    .Y(_535_)
);

NAND2X1 _1470_ (
    .A(_379_),
    .B(_465_),
    .Y(_536_)
);

OAI21X1 _1471_ (
    .A(_388_),
    .B(_536_),
    .C(_483_),
    .Y(_537_)
);

INVX1 _1472_ (
    .A(_534_),
    .Y(_538_)
);

NOR2X1 _1473_ (
    .A(_538_),
    .B(_537_),
    .Y(_539_)
);

OAI21X1 _1474_ (
    .A(_535_),
    .B(_539_),
    .C(ABCmd_i[7]),
    .Y(_540_)
);

NOR2X1 _1475_ (
    .A(ABCmd_i[7]),
    .B(AZ),
    .Y(_541_)
);

NOR2X1 _1476_ (
    .A(_541_),
    .B(_733_),
    .Y(_542_)
);

AOI21X1 _1477_ (
    .A(_293_),
    .B(_296_),
    .C(_295_),
    .Y(_543_)
);

OAI21X1 _1478_ (
    .A(_543_),
    .B(_298_),
    .C(ABCmd_i[7]),
    .Y(_544_)
);

NOR2X1 _1479_ (
    .A(ABCmd_i[7]),
    .B(ACC[2]),
    .Y(_545_)
);

NOR2X1 _1480_ (
    .A(_545_),
    .B(_25_),
    .Y(_546_)
);

AOI22X1 _1481_ (
    .A(_544_),
    .B(_546_),
    .C(_540_),
    .D(_542_),
    .Y(_547_)
);

OAI21X1 _1482_ (
    .A(_730_),
    .B(_547_),
    .C(_480_),
    .Y(_11_)
);

INVX1 _1483_ (
    .A(_924_[3]),
    .Y(_548_)
);

INVX1 _1484_ (
    .A(AV),
    .Y(_549_)
);

OAI21X1 _1485_ (
    .A(_549_),
    .B(_733_),
    .C(_401_),
    .Y(_550_)
);

INVX1 _1486_ (
    .A(_533_),
    .Y(_551_)
);

OAI21X1 _1487_ (
    .A(_487_),
    .B(_495_),
    .C(_491_),
    .Y(_552_)
);

INVX1 _1488_ (
    .A(_552_),
    .Y(_553_)
);

AOI21X1 _1489_ (
    .A(_514_),
    .B(_511_),
    .C(_510_),
    .Y(_554_)
);

NAND2X1 _1490_ (
    .A(AI[4]),
    .B(BI[7]),
    .Y(_555_)
);

INVX1 _1491_ (
    .A(_555_),
    .Y(_556_)
);

NOR2X1 _1492_ (
    .A(_127_),
    .B(_165_),
    .Y(_557_)
);

OAI22X1 _1493_ (
    .A(_501_),
    .B(_502_),
    .C(_499_),
    .D(_505_),
    .Y(_558_)
);

NAND2X1 _1494_ (
    .A(_557_),
    .B(_558_),
    .Y(_559_)
);

OR2X2 _1495_ (
    .A(_558_),
    .B(_557_),
    .Y(_560_)
);

NAND3X1 _1496_ (
    .A(_556_),
    .B(_559_),
    .C(_560_),
    .Y(_561_)
);

INVX2 _1497_ (
    .A(BI[7]),
    .Y(_562_)
);

NAND2X1 _1498_ (
    .A(_559_),
    .B(_560_),
    .Y(_563_)
);

OAI21X1 _1499_ (
    .A(_202_),
    .B(_562_),
    .C(_563_),
    .Y(_564_)
);

NAND2X1 _1500_ (
    .A(AI[6]),
    .B(BI_4_bF$buf3),
    .Y(_565_)
);

NAND2X1 _1501_ (
    .A(\u_ALU8.AI7 ),
    .B(BI[5]),
    .Y(_566_)
);

NOR2X1 _1502_ (
    .A(_565_),
    .B(_566_),
    .Y(_567_)
);

INVX1 _1503_ (
    .A(_567_),
    .Y(_568_)
);

INVX1 _1504_ (
    .A(BI[5]),
    .Y(_569_)
);

OAI21X1 _1505_ (
    .A(_429_),
    .B(_569_),
    .C(_502_),
    .Y(_570_)
);

AND2X2 _1506_ (
    .A(_568_),
    .B(_570_),
    .Y(_571_)
);

AOI21X1 _1507_ (
    .A(_564_),
    .B(_561_),
    .C(_571_),
    .Y(_572_)
);

INVX1 _1508_ (
    .A(_572_),
    .Y(_573_)
);

NAND3X1 _1509_ (
    .A(_571_),
    .B(_561_),
    .C(_564_),
    .Y(_574_)
);

NAND3X1 _1510_ (
    .A(_573_),
    .B(_574_),
    .C(_554_),
    .Y(_575_)
);

OAI21X1 _1511_ (
    .A(_497_),
    .B(_512_),
    .C(_516_),
    .Y(_576_)
);

INVX1 _1512_ (
    .A(_574_),
    .Y(_577_)
);

OAI21X1 _1513_ (
    .A(_572_),
    .B(_577_),
    .C(_576_),
    .Y(_578_)
);

NAND3X1 _1514_ (
    .A(_553_),
    .B(_578_),
    .C(_575_),
    .Y(_579_)
);

NAND3X1 _1515_ (
    .A(_574_),
    .B(_576_),
    .C(_573_),
    .Y(_580_)
);

OAI21X1 _1516_ (
    .A(_572_),
    .B(_577_),
    .C(_554_),
    .Y(_581_)
);

NAND3X1 _1517_ (
    .A(_552_),
    .B(_580_),
    .C(_581_),
    .Y(_582_)
);

NAND2X1 _1518_ (
    .A(_582_),
    .B(_579_),
    .Y(_583_)
);

NAND3X1 _1519_ (
    .A(_526_),
    .B(_528_),
    .C(_583_),
    .Y(_584_)
);

AOI21X1 _1520_ (
    .A(_517_),
    .B(_513_),
    .C(_519_),
    .Y(_585_)
);

OAI21X1 _1521_ (
    .A(_485_),
    .B(_585_),
    .C(_526_),
    .Y(_586_)
);

NAND3X1 _1522_ (
    .A(_579_),
    .B(_582_),
    .C(_586_),
    .Y(_587_)
);

NAND2X1 _1523_ (
    .A(_587_),
    .B(_584_),
    .Y(_588_)
);

NOR3X1 _1524_ (
    .A(_551_),
    .B(_588_),
    .C(_535_),
    .Y(_589_)
);

AOI21X1 _1525_ (
    .A(_537_),
    .B(_538_),
    .C(_551_),
    .Y(_590_)
);

INVX1 _1526_ (
    .A(_588_),
    .Y(_591_)
);

OAI21X1 _1527_ (
    .A(_591_),
    .B(_590_),
    .C(ABCmd_i[7]),
    .Y(_592_)
);

OAI21X1 _1528_ (
    .A(_589_),
    .B(_592_),
    .C(_550_),
    .Y(_593_)
);

NAND2X1 _1529_ (
    .A(_300_),
    .B(_289_),
    .Y(_594_)
);

NAND2X1 _1530_ (
    .A(_297_),
    .B(_594_),
    .Y(_595_)
);

NAND2X1 _1531_ (
    .A(_301_),
    .B(_595_),
    .Y(_596_)
);

NAND2X1 _1532_ (
    .A(ACC[3]),
    .B(_54_),
    .Y(_597_)
);

OAI21X1 _1533_ (
    .A(_54_),
    .B(_596_),
    .C(_597_),
    .Y(_598_)
);

AOI21X1 _1534_ (
    .A(_598_),
    .B(_721_),
    .C(_730_),
    .Y(_599_)
);

AOI22X1 _1535_ (
    .A(_548_),
    .B(_730_),
    .C(_593_),
    .D(_599_),
    .Y(_12_)
);

INVX1 _1536_ (
    .A(_924_[4]),
    .Y(_600_)
);

NAND2X1 _1537_ (
    .A(_580_),
    .B(_582_),
    .Y(_601_)
);

INVX1 _1538_ (
    .A(_601_),
    .Y(_602_)
);

OAI21X1 _1539_ (
    .A(_555_),
    .B(_563_),
    .C(_559_),
    .Y(_603_)
);

INVX1 _1540_ (
    .A(_603_),
    .Y(_604_)
);

INVX1 _1541_ (
    .A(\u_ALU8.AI7 ),
    .Y(_605_)
);

NOR2X1 _1542_ (
    .A(_127_),
    .B(_562_),
    .Y(_606_)
);

NOR2X1 _1543_ (
    .A(_429_),
    .B(_165_),
    .Y(_607_)
);

NOR2X1 _1544_ (
    .A(_607_),
    .B(_567_),
    .Y(_608_)
);

AOI21X1 _1545_ (
    .A(BI[6]),
    .B(_567_),
    .C(_608_),
    .Y(_609_)
);

NAND2X1 _1546_ (
    .A(_606_),
    .B(_609_),
    .Y(_610_)
);

NOR2X1 _1547_ (
    .A(_165_),
    .B(_568_),
    .Y(_611_)
);

OAI22X1 _1548_ (
    .A(_127_),
    .B(_562_),
    .C(_608_),
    .D(_611_),
    .Y(_612_)
);

NAND2X1 _1549_ (
    .A(_612_),
    .B(_610_),
    .Y(_613_)
);

OAI21X1 _1550_ (
    .A(_605_),
    .B(_569_),
    .C(_613_),
    .Y(_614_)
);

INVX1 _1551_ (
    .A(_566_),
    .Y(_615_)
);

NAND3X1 _1552_ (
    .A(_615_),
    .B(_612_),
    .C(_610_),
    .Y(_616_)
);

NAND2X1 _1553_ (
    .A(_616_),
    .B(_614_),
    .Y(_617_)
);

NOR2X1 _1554_ (
    .A(_574_),
    .B(_617_),
    .Y(_618_)
);

AOI21X1 _1555_ (
    .A(_614_),
    .B(_616_),
    .C(_577_),
    .Y(_619_)
);

OAI21X1 _1556_ (
    .A(_619_),
    .B(_618_),
    .C(_604_),
    .Y(_620_)
);

OR2X2 _1557_ (
    .A(_617_),
    .B(_574_),
    .Y(_621_)
);

INVX1 _1558_ (
    .A(_619_),
    .Y(_622_)
);

NAND3X1 _1559_ (
    .A(_603_),
    .B(_621_),
    .C(_622_),
    .Y(_623_)
);

NAND2X1 _1560_ (
    .A(_620_),
    .B(_623_),
    .Y(_624_)
);

NAND2X1 _1561_ (
    .A(_624_),
    .B(_602_),
    .Y(_625_)
);

NAND3X1 _1562_ (
    .A(_620_),
    .B(_623_),
    .C(_601_),
    .Y(_626_)
);

NAND2X1 _1563_ (
    .A(_626_),
    .B(_625_),
    .Y(_627_)
);

NOR2X1 _1564_ (
    .A(_389_),
    .B(_472_),
    .Y(_628_)
);

NOR2X1 _1565_ (
    .A(_588_),
    .B(_534_),
    .Y(_629_)
);

NAND3X1 _1566_ (
    .A(_311_),
    .B(_629_),
    .C(_628_),
    .Y(_630_)
);

NAND2X1 _1567_ (
    .A(_587_),
    .B(_533_),
    .Y(_631_)
);

AOI22X1 _1568_ (
    .A(_584_),
    .B(_631_),
    .C(_629_),
    .D(_482_),
    .Y(_632_)
);

AOI21X1 _1569_ (
    .A(_632_),
    .B(_630_),
    .C(_627_),
    .Y(_633_)
);

INVX1 _1570_ (
    .A(_627_),
    .Y(_634_)
);

NAND2X1 _1571_ (
    .A(_584_),
    .B(_631_),
    .Y(_635_)
);

OAI21X1 _1572_ (
    .A(_534_),
    .B(_588_),
    .C(_635_),
    .Y(_636_)
);

AOI21X1 _1573_ (
    .A(_584_),
    .B(_631_),
    .C(_482_),
    .Y(_637_)
);

OAI21X1 _1574_ (
    .A(_388_),
    .B(_536_),
    .C(_637_),
    .Y(_638_)
);

AOI21X1 _1575_ (
    .A(_638_),
    .B(_636_),
    .C(_634_),
    .Y(_639_)
);

OAI21X1 _1576_ (
    .A(_639_),
    .B(_633_),
    .C(ABCmd_i[7]),
    .Y(_640_)
);

OR2X2 _1577_ (
    .A(ABCmd_i[7]),
    .B(CO),
    .Y(_641_)
);

NAND3X1 _1578_ (
    .A(_25_),
    .B(_641_),
    .C(_640_),
    .Y(_642_)
);

INVX1 _1579_ (
    .A(_303_),
    .Y(_643_)
);

OAI21X1 _1580_ (
    .A(_302_),
    .B(_282_),
    .C(_301_),
    .Y(_644_)
);

NAND2X1 _1581_ (
    .A(_644_),
    .B(_643_),
    .Y(_645_)
);

NAND2X1 _1582_ (
    .A(ACC[4]),
    .B(_54_),
    .Y(_646_)
);

OAI21X1 _1583_ (
    .A(_54_),
    .B(_645_),
    .C(_646_),
    .Y(_647_)
);

AOI21X1 _1584_ (
    .A(_647_),
    .B(_721_),
    .C(_730_),
    .Y(_648_)
);

AOI22X1 _1585_ (
    .A(_600_),
    .B(_730_),
    .C(_642_),
    .D(_648_),
    .Y(_13_)
);

INVX1 _1586_ (
    .A(_924_[5]),
    .Y(_649_)
);

AOI21X1 _1587_ (
    .A(_609_),
    .B(_606_),
    .C(_611_),
    .Y(_650_)
);

NOR2X1 _1588_ (
    .A(_605_),
    .B(_562_),
    .Y(_651_)
);

NAND2X1 _1589_ (
    .A(_607_),
    .B(_651_),
    .Y(_652_)
);

OAI22X1 _1590_ (
    .A(_605_),
    .B(_165_),
    .C(_429_),
    .D(_562_),
    .Y(_653_)
);

NAND2X1 _1591_ (
    .A(_653_),
    .B(_652_),
    .Y(_654_)
);

OR2X2 _1592_ (
    .A(_616_),
    .B(_654_),
    .Y(_655_)
);

OAI21X1 _1593_ (
    .A(_566_),
    .B(_613_),
    .C(_654_),
    .Y(_656_)
);

NAND2X1 _1594_ (
    .A(_656_),
    .B(_655_),
    .Y(_657_)
);

NAND2X1 _1595_ (
    .A(_650_),
    .B(_657_),
    .Y(_658_)
);

OR2X2 _1596_ (
    .A(_657_),
    .B(_650_),
    .Y(_659_)
);

NAND2X1 _1597_ (
    .A(_658_),
    .B(_659_),
    .Y(_660_)
);

NAND3X1 _1598_ (
    .A(_621_),
    .B(_623_),
    .C(_660_),
    .Y(_661_)
);

OAI21X1 _1599_ (
    .A(_604_),
    .B(_619_),
    .C(_621_),
    .Y(_662_)
);

NAND3X1 _1600_ (
    .A(_658_),
    .B(_659_),
    .C(_662_),
    .Y(_663_)
);

NAND2X1 _1601_ (
    .A(_663_),
    .B(_661_),
    .Y(_664_)
);

NOR2X1 _1602_ (
    .A(_664_),
    .B(_627_),
    .Y(_665_)
);

NAND3X1 _1603_ (
    .A(_636_),
    .B(_665_),
    .C(_638_),
    .Y(_666_)
);

NAND3X1 _1604_ (
    .A(_634_),
    .B(_636_),
    .C(_638_),
    .Y(_667_)
);

NAND3X1 _1605_ (
    .A(_626_),
    .B(_664_),
    .C(_667_),
    .Y(_668_)
);

INVX1 _1606_ (
    .A(_401_),
    .Y(_669_)
);

OR2X2 _1607_ (
    .A(_664_),
    .B(_626_),
    .Y(_670_)
);

AND2X2 _1608_ (
    .A(_670_),
    .B(_669_),
    .Y(_671_)
);

NAND3X1 _1609_ (
    .A(_666_),
    .B(_671_),
    .C(_668_),
    .Y(_672_)
);

AOI21X1 _1610_ (
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_673_)
);

OAI21X1 _1611_ (
    .A(_673_),
    .B(_308_),
    .C(ABCmd_i[7]),
    .Y(_674_)
);

INVX1 _1612_ (
    .A(ACC[5]),
    .Y(_675_)
);

AOI21X1 _1613_ (
    .A(_54_),
    .B(_675_),
    .C(state[1]),
    .Y(_676_)
);

AOI21X1 _1614_ (
    .A(_674_),
    .B(_676_),
    .C(_730_),
    .Y(_677_)
);

AOI22X1 _1615_ (
    .A(_649_),
    .B(_730_),
    .C(_672_),
    .D(_677_),
    .Y(_14_)
);

INVX1 _1616_ (
    .A(_924_[6]),
    .Y(_678_)
);

OAI21X1 _1617_ (
    .A(_626_),
    .B(_664_),
    .C(_663_),
    .Y(_679_)
);

INVX1 _1618_ (
    .A(_679_),
    .Y(_680_)
);

OAI21X1 _1619_ (
    .A(_650_),
    .B(_657_),
    .C(_655_),
    .Y(_681_)
);

INVX1 _1620_ (
    .A(_681_),
    .Y(_682_)
);

OAI21X1 _1621_ (
    .A(_429_),
    .B(_165_),
    .C(_651_),
    .Y(_683_)
);

OR2X2 _1622_ (
    .A(_682_),
    .B(_683_),
    .Y(_684_)
);

NAND2X1 _1623_ (
    .A(_683_),
    .B(_682_),
    .Y(_685_)
);

NAND2X1 _1624_ (
    .A(_685_),
    .B(_684_),
    .Y(_686_)
);

NAND3X1 _1625_ (
    .A(_686_),
    .B(_680_),
    .C(_666_),
    .Y(_687_)
);

OR2X2 _1626_ (
    .A(_627_),
    .B(_664_),
    .Y(_688_)
);

AOI21X1 _1627_ (
    .A(_632_),
    .B(_630_),
    .C(_688_),
    .Y(_689_)
);

INVX1 _1628_ (
    .A(_686_),
    .Y(_690_)
);

OAI21X1 _1629_ (
    .A(_679_),
    .B(_689_),
    .C(_690_),
    .Y(_691_)
);

NAND3X1 _1630_ (
    .A(_669_),
    .B(_687_),
    .C(_691_),
    .Y(_692_)
);

NAND3X1 _1631_ (
    .A(_309_),
    .B(_385_),
    .C(_308_),
    .Y(_693_)
);

OAI21X1 _1632_ (
    .A(_287_),
    .B(_386_),
    .C(_307_),
    .Y(_694_)
);

NAND2X1 _1633_ (
    .A(_693_),
    .B(_694_),
    .Y(_695_)
);

NAND2X1 _1634_ (
    .A(ACC[6]),
    .B(_54_),
    .Y(_696_)
);

OAI21X1 _1635_ (
    .A(_54_),
    .B(_695_),
    .C(_696_),
    .Y(_697_)
);

AOI21X1 _1636_ (
    .A(_697_),
    .B(_721_),
    .C(_730_),
    .Y(_698_)
);

AOI22X1 _1637_ (
    .A(_678_),
    .B(_730_),
    .C(_692_),
    .D(_698_),
    .Y(_15_)
);

INVX1 _1638_ (
    .A(_924_[7]),
    .Y(_699_)
);

AOI21X1 _1639_ (
    .A(_666_),
    .B(_680_),
    .C(_686_),
    .Y(_700_)
);

OAI21X1 _1640_ (
    .A(_683_),
    .B(_682_),
    .C(_652_),
    .Y(_701_)
);

OAI21X1 _1641_ (
    .A(_701_),
    .B(_700_),
    .C(_669_),
    .Y(_702_)
);

NAND3X1 _1642_ (
    .A(_381_),
    .B(_247_),
    .C(_387_),
    .Y(_703_)
);

OAI21X1 _1643_ (
    .A(_246_),
    .B(_269_),
    .C(_310_),
    .Y(_704_)
);

NAND2X1 _1644_ (
    .A(_704_),
    .B(_703_),
    .Y(_705_)
);

NAND2X1 _1645_ (
    .A(AN),
    .B(_54_),
    .Y(_706_)
);

OAI21X1 _1646_ (
    .A(_54_),
    .B(_705_),
    .C(_706_),
    .Y(_707_)
);

AOI21X1 _1647_ (
    .A(_707_),
    .B(_721_),
    .C(_730_),
    .Y(_708_)
);

AOI22X1 _1648_ (
    .A(_699_),
    .B(_730_),
    .C(_702_),
    .D(_708_),
    .Y(_16_)
);

NAND2X1 _1649_ (
    .A(AI[0]),
    .B(_723__bF$buf3),
    .Y(_709_)
);

OAI21X1 _1650_ (
    .A(_40_),
    .B(_723__bF$buf2),
    .C(_709_),
    .Y(_17_)
);

NAND2X1 _1651_ (
    .A(AI[1]),
    .B(_723__bF$buf1),
    .Y(_710_)
);

OAI21X1 _1652_ (
    .A(_42_),
    .B(_723__bF$buf0),
    .C(_710_),
    .Y(_18_)
);

NAND2X1 _1653_ (
    .A(AI[2]),
    .B(_723__bF$buf3),
    .Y(_711_)
);

OAI21X1 _1654_ (
    .A(_44_),
    .B(_723__bF$buf2),
    .C(_711_),
    .Y(_19_)
);

NAND2X1 _1655_ (
    .A(AI[3]),
    .B(_723__bF$buf1),
    .Y(_712_)
);

OAI21X1 _1656_ (
    .A(_46_),
    .B(_723__bF$buf0),
    .C(_712_),
    .Y(_20_)
);

NAND2X1 _1657_ (
    .A(AI[4]),
    .B(_723__bF$buf3),
    .Y(_713_)
);

OAI21X1 _1658_ (
    .A(_48_),
    .B(_723__bF$buf2),
    .C(_713_),
    .Y(_21_)
);

NAND2X1 _1659_ (
    .A(AI[5]),
    .B(_723__bF$buf1),
    .Y(_714_)
);

OAI21X1 _1660_ (
    .A(_50_),
    .B(_723__bF$buf0),
    .C(_714_),
    .Y(_22_)
);

NAND2X1 _1661_ (
    .A(AI[6]),
    .B(_723__bF$buf3),
    .Y(_715_)
);

OAI21X1 _1662_ (
    .A(_52_),
    .B(_723__bF$buf2),
    .C(_715_),
    .Y(_23_)
);

NAND2X1 _1663_ (
    .A(\u_ALU8.AI7 ),
    .B(_723__bF$buf1),
    .Y(_716_)
);

OAI21X1 _1664_ (
    .A(_54_),
    .B(_723__bF$buf0),
    .C(_716_),
    .Y(_24_)
);

DFFPOSX1 _1665_ (
    .CLK(clk_bF$buf4),
    .D(_1_),
    .Q(BI[0])
);

DFFPOSX1 _1666_ (
    .CLK(clk_bF$buf3),
    .D(_2_),
    .Q(BI[1])
);

DFFPOSX1 _1667_ (
    .CLK(clk_bF$buf2),
    .D(_3_),
    .Q(BI[2])
);

DFFPOSX1 _1668_ (
    .CLK(clk_bF$buf1),
    .D(_4_),
    .Q(BI[3])
);

DFFPOSX1 _1669_ (
    .CLK(clk_bF$buf0),
    .D(_5_),
    .Q(BI[4])
);

DFFPOSX1 _1670_ (
    .CLK(clk_bF$buf4),
    .D(_6_),
    .Q(BI[5])
);

DFFPOSX1 _1671_ (
    .CLK(clk_bF$buf3),
    .D(_7_),
    .Q(BI[6])
);

DFFPOSX1 _1672_ (
    .CLK(clk_bF$buf2),
    .D(_8_),
    .Q(BI[7])
);

DFFPOSX1 _1673_ (
    .CLK(clk_bF$buf1),
    .D(_9_),
    .Q(_924_[0])
);

DFFPOSX1 _1674_ (
    .CLK(clk_bF$buf0),
    .D(_10_),
    .Q(_924_[1])
);

DFFPOSX1 _1675_ (
    .CLK(clk_bF$buf4),
    .D(_11_),
    .Q(_924_[2])
);

DFFPOSX1 _1676_ (
    .CLK(clk_bF$buf3),
    .D(_12_),
    .Q(_924_[3])
);

DFFPOSX1 _1677_ (
    .CLK(clk_bF$buf2),
    .D(_13_),
    .Q(_924_[4])
);

DFFPOSX1 _1678_ (
    .CLK(clk_bF$buf1),
    .D(_14_),
    .Q(_924_[5])
);

DFFPOSX1 _1679_ (
    .CLK(clk_bF$buf0),
    .D(_15_),
    .Q(_924_[6])
);

DFFPOSX1 _1680_ (
    .CLK(clk_bF$buf4),
    .D(_16_),
    .Q(_924_[7])
);

DFFPOSX1 _1681_ (
    .CLK(clk_bF$buf3),
    .D(_17_),
    .Q(AI[0])
);

DFFPOSX1 _1682_ (
    .CLK(clk_bF$buf2),
    .D(_18_),
    .Q(AI[1])
);

DFFPOSX1 _1683_ (
    .CLK(clk_bF$buf1),
    .D(_19_),
    .Q(AI[2])
);

DFFPOSX1 _1684_ (
    .CLK(clk_bF$buf0),
    .D(_20_),
    .Q(AI[3])
);

DFFPOSX1 _1685_ (
    .CLK(clk_bF$buf4),
    .D(_21_),
    .Q(AI[4])
);

DFFPOSX1 _1686_ (
    .CLK(clk_bF$buf3),
    .D(_22_),
    .Q(AI[5])
);

DFFPOSX1 _1687_ (
    .CLK(clk_bF$buf2),
    .D(_23_),
    .Q(AI[6])
);

DFFPOSX1 _1688_ (
    .CLK(clk_bF$buf1),
    .D(_24_),
    .Q(\u_ALU8.AI7 )
);

DFFSR _1689_ (
    .CLK(clk_bF$buf0),
    .D(_926_[0]),
    .Q(state[0]),
    .R(VDD),
    .S(_0_)
);

DFFSR _1690_ (
    .CLK(clk_bF$buf4),
    .D(_926_[1]),
    .Q(state[1]),
    .R(_0_),
    .S(VDD)
);

DFFSR _1691_ (
    .CLK(clk_bF$buf3),
    .D(_926_[2]),
    .Q(state[2]),
    .R(_0_),
    .S(VDD)
);

INVX1 _1692_ (
    .A(ABCmd_i_2_bF$buf3),
    .Y(_862_)
);

INVX4 _1693_ (
    .A(ABCmd_i[3]),
    .Y(_863_)
);

OAI21X1 _1694_ (
    .A(_862_),
    .B(_863_),
    .C(ABCmd_i[4]),
    .Y(_864_)
);

NOR2X1 _1695_ (
    .A(ABCmd_i[5]),
    .B(_864_),
    .Y(_865_)
);

INVX1 _1696_ (
    .A(_865_),
    .Y(_866_)
);

INVX2 _1697_ (
    .A(ABCmd_i[1]),
    .Y(_867_)
);

NAND2X1 _1698_ (
    .A(ABCmd_i[0]),
    .B(_867_),
    .Y(_868_)
);

INVX2 _1699_ (
    .A(ABCmd_i[0]),
    .Y(_869_)
);

NAND2X1 _1700_ (
    .A(BI_0_bF$buf3),
    .B(_869_),
    .Y(_870_)
);

NAND2X1 _1701_ (
    .A(AI[0]),
    .B(ABCmd_i[1]),
    .Y(_871_)
);

AOI22X1 _1702_ (
    .A(BI_0_bF$buf2),
    .B(_871_),
    .C(_868_),
    .D(_870_),
    .Y(_872_)
);

INVX2 _1703_ (
    .A(ABCmd_i[5]),
    .Y(_873_)
);

INVX1 _1704_ (
    .A(BI_0_bF$buf1),
    .Y(_874_)
);

INVX1 _1705_ (
    .A(AI[0]),
    .Y(_875_)
);

OAI21X1 _1706_ (
    .A(ABCmd_i[0]),
    .B(_874_),
    .C(_875_),
    .Y(_876_)
);

NAND2X1 _1707_ (
    .A(_873_),
    .B(_876_),
    .Y(_877_)
);

NAND2X1 _1708_ (
    .A(AI[1]),
    .B(ABCmd_i[5]),
    .Y(_878_)
);

OAI21X1 _1709_ (
    .A(_872_),
    .B(_877_),
    .C(_878_),
    .Y(_879_)
);

OAI21X1 _1710_ (
    .A(BI_0_bF$buf0),
    .B(ABCmd_i_2_bF$buf2),
    .C(_863_),
    .Y(_880_)
);

AOI21X1 _1711_ (
    .A(BI_0_bF$buf3),
    .B(ABCmd_i_2_bF$buf1),
    .C(_880_),
    .Y(_881_)
);

NOR2X1 _1712_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(_863_),
    .Y(_882_)
);

OAI21X1 _1713_ (
    .A(_882_),
    .B(_881_),
    .C(_879_),
    .Y(_883_)
);

OAI21X1 _1714_ (
    .A(_879_),
    .B(_881_),
    .C(_883_),
    .Y(_884_)
);

OR2X2 _1715_ (
    .A(_884_),
    .B(_866_),
    .Y(_885_)
);

OAI21X1 _1716_ (
    .A(ABCmd_i[5]),
    .B(_864_),
    .C(_884_),
    .Y(_886_)
);

NAND2X1 _1717_ (
    .A(_886_),
    .B(_885_),
    .Y(_887_)
);

INVX1 _1718_ (
    .A(_887_),
    .Y(ACC[0])
);

NOR2X1 _1719_ (
    .A(_881_),
    .B(_879_),
    .Y(_888_)
);

OAI21X1 _1720_ (
    .A(_866_),
    .B(_888_),
    .C(_883_),
    .Y(_889_)
);

NAND2X1 _1721_ (
    .A(ABCmd_i[5]),
    .B(AI[2]),
    .Y(_890_)
);

NAND3X1 _1722_ (
    .A(AI[1]),
    .B(BI_1_bF$buf2),
    .C(_869_),
    .Y(_891_)
);

AOI22X1 _1723_ (
    .A(_867_),
    .B(BI_1_bF$buf1),
    .C(_891_),
    .D(_868_),
    .Y(_892_)
);

INVX1 _1724_ (
    .A(BI_1_bF$buf0),
    .Y(_893_)
);

NOR2X1 _1725_ (
    .A(ABCmd_i[0]),
    .B(_893_),
    .Y(_894_)
);

OAI21X1 _1726_ (
    .A(AI[1]),
    .B(_894_),
    .C(_873_),
    .Y(_895_)
);

OAI21X1 _1727_ (
    .A(_892_),
    .B(_895_),
    .C(_890_),
    .Y(_896_)
);

OAI21X1 _1728_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI_1_bF$buf3),
    .C(_863_),
    .Y(_897_)
);

AOI21X1 _1729_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_1_bF$buf2),
    .C(_897_),
    .Y(_898_)
);

INVX1 _1730_ (
    .A(_898_),
    .Y(_899_)
);

OAI21X1 _1731_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_863_),
    .C(_899_),
    .Y(_900_)
);

MUX2X1 _1732_ (
    .A(_900_),
    .B(_899_),
    .S(_896_),
    .Y(_901_)
);

NAND2X1 _1733_ (
    .A(_901_),
    .B(_889_),
    .Y(_902_)
);

INVX1 _1734_ (
    .A(_881_),
    .Y(_903_)
);

OAI21X1 _1735_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(_863_),
    .C(_903_),
    .Y(_904_)
);

MUX2X1 _1736_ (
    .A(ABCmd_i[1]),
    .B(_874_),
    .S(ABCmd_i[0]),
    .Y(_905_)
);

OAI21X1 _1737_ (
    .A(_875_),
    .B(_867_),
    .C(BI_0_bF$buf2),
    .Y(_906_)
);

NAND2X1 _1738_ (
    .A(_906_),
    .B(_905_),
    .Y(_907_)
);

NAND3X1 _1739_ (
    .A(_873_),
    .B(_876_),
    .C(_907_),
    .Y(_908_)
);

NAND3X1 _1740_ (
    .A(_878_),
    .B(_903_),
    .C(_908_),
    .Y(_909_)
);

AOI22X1 _1741_ (
    .A(_879_),
    .B(_904_),
    .C(_909_),
    .D(_865_),
    .Y(_910_)
);

OAI21X1 _1742_ (
    .A(_882_),
    .B(_898_),
    .C(_896_),
    .Y(_911_)
);

OAI21X1 _1743_ (
    .A(_896_),
    .B(_898_),
    .C(_911_),
    .Y(_912_)
);

NAND2X1 _1744_ (
    .A(_910_),
    .B(_912_),
    .Y(_913_)
);

NAND2X1 _1745_ (
    .A(_913_),
    .B(_902_),
    .Y(_914_)
);

INVX1 _1746_ (
    .A(_914_),
    .Y(ACC[1])
);

NOR2X1 _1747_ (
    .A(_898_),
    .B(_896_),
    .Y(_915_)
);

OAI21X1 _1748_ (
    .A(_915_),
    .B(_910_),
    .C(_911_),
    .Y(_916_)
);

NAND2X1 _1749_ (
    .A(ABCmd_i[5]),
    .B(AI[3]),
    .Y(_917_)
);

INVX1 _1750_ (
    .A(BI[2]),
    .Y(_918_)
);

NOR2X1 _1751_ (
    .A(ABCmd_i[0]),
    .B(_918_),
    .Y(_919_)
);

NAND2X1 _1752_ (
    .A(AI[2]),
    .B(_919_),
    .Y(_920_)
);

AOI22X1 _1753_ (
    .A(_867_),
    .B(BI[2]),
    .C(_920_),
    .D(_868_),
    .Y(_921_)
);

OAI21X1 _1754_ (
    .A(AI[2]),
    .B(_919_),
    .C(_873_),
    .Y(_922_)
);

OAI21X1 _1755_ (
    .A(_922_),
    .B(_921_),
    .C(_917_),
    .Y(_923_)
);

OAI21X1 _1756_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[2]),
    .C(_863_),
    .Y(_734_)
);

AOI21X1 _1757_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI[2]),
    .C(_734_),
    .Y(_735_)
);

INVX1 _1758_ (
    .A(_735_),
    .Y(_736_)
);

OAI21X1 _1759_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_863_),
    .C(_736_),
    .Y(_737_)
);

MUX2X1 _1760_ (
    .A(_737_),
    .B(_736_),
    .S(_923_),
    .Y(_738_)
);

NAND2X1 _1761_ (
    .A(_738_),
    .B(_916_),
    .Y(_739_)
);

OAI21X1 _1762_ (
    .A(_882_),
    .B(_735_),
    .C(_923_),
    .Y(_740_)
);

OAI21X1 _1763_ (
    .A(_923_),
    .B(_735_),
    .C(_740_),
    .Y(_741_)
);

NAND3X1 _1764_ (
    .A(_911_),
    .B(_741_),
    .C(_902_),
    .Y(_742_)
);

NAND2X1 _1765_ (
    .A(_739_),
    .B(_742_),
    .Y(_743_)
);

INVX1 _1766_ (
    .A(_743_),
    .Y(ACC[2])
);

INVX1 _1767_ (
    .A(_740_),
    .Y(_744_)
);

AND2X2 _1768_ (
    .A(_916_),
    .B(_738_),
    .Y(_745_)
);

NAND2X1 _1769_ (
    .A(ABCmd_i[5]),
    .B(AI[4]),
    .Y(_746_)
);

AND2X2 _1770_ (
    .A(_869_),
    .B(BI_3_bF$buf0),
    .Y(_747_)
);

NAND2X1 _1771_ (
    .A(AI[3]),
    .B(_747_),
    .Y(_748_)
);

AOI22X1 _1772_ (
    .A(_867_),
    .B(BI_3_bF$buf3),
    .C(_748_),
    .D(_868_),
    .Y(_749_)
);

OAI21X1 _1773_ (
    .A(AI[3]),
    .B(_747_),
    .C(_873_),
    .Y(_750_)
);

OAI21X1 _1774_ (
    .A(_750_),
    .B(_749_),
    .C(_746_),
    .Y(_751_)
);

OAI21X1 _1775_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI_3_bF$buf2),
    .C(_863_),
    .Y(_752_)
);

AOI21X1 _1776_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI_3_bF$buf1),
    .C(_752_),
    .Y(_753_)
);

OAI21X1 _1777_ (
    .A(_882_),
    .B(_753_),
    .C(_751_),
    .Y(_754_)
);

OAI21X1 _1778_ (
    .A(_751_),
    .B(_753_),
    .C(_754_),
    .Y(_755_)
);

INVX1 _1779_ (
    .A(_755_),
    .Y(_756_)
);

OAI21X1 _1780_ (
    .A(_744_),
    .B(_745_),
    .C(_756_),
    .Y(_757_)
);

NAND3X1 _1781_ (
    .A(_740_),
    .B(_755_),
    .C(_739_),
    .Y(_758_)
);

NAND2X1 _1782_ (
    .A(_758_),
    .B(_757_),
    .Y(_759_)
);

INVX1 _1783_ (
    .A(_759_),
    .Y(ACC[3])
);

INVX1 _1784_ (
    .A(ABCmd_i[6]),
    .Y(_760_)
);

AOI21X1 _1785_ (
    .A(_743_),
    .B(_914_),
    .C(_760_),
    .Y(_761_)
);

NAND3X1 _1786_ (
    .A(_757_),
    .B(_758_),
    .C(_761_),
    .Y(_762_)
);

NAND2X1 _1787_ (
    .A(_740_),
    .B(_739_),
    .Y(_763_)
);

INVX1 _1788_ (
    .A(_754_),
    .Y(_764_)
);

AOI21X1 _1789_ (
    .A(_763_),
    .B(_756_),
    .C(_764_),
    .Y(_765_)
);

NAND2X1 _1790_ (
    .A(ABCmd_i[5]),
    .B(AI[5]),
    .Y(_766_)
);

AND2X2 _1791_ (
    .A(_869_),
    .B(BI_4_bF$buf2),
    .Y(_767_)
);

NAND2X1 _1792_ (
    .A(AI[4]),
    .B(_767_),
    .Y(_768_)
);

AOI22X1 _1793_ (
    .A(_867_),
    .B(BI_4_bF$buf1),
    .C(_768_),
    .D(_868_),
    .Y(_769_)
);

OAI21X1 _1794_ (
    .A(AI[4]),
    .B(_767_),
    .C(_873_),
    .Y(_770_)
);

OAI21X1 _1795_ (
    .A(_770_),
    .B(_769_),
    .C(_766_),
    .Y(_771_)
);

OAI21X1 _1796_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_4_bF$buf0),
    .C(_863_),
    .Y(_772_)
);

AOI21X1 _1797_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(BI_4_bF$buf3),
    .C(_772_),
    .Y(_773_)
);

OAI21X1 _1798_ (
    .A(_882_),
    .B(_773_),
    .C(_771_),
    .Y(_774_)
);

OAI21X1 _1799_ (
    .A(_771_),
    .B(_773_),
    .C(_774_),
    .Y(_775_)
);

AOI21X1 _1800_ (
    .A(_762_),
    .B(_765_),
    .C(_775_),
    .Y(_776_)
);

NOR2X1 _1801_ (
    .A(_738_),
    .B(_916_),
    .Y(_777_)
);

OAI21X1 _1802_ (
    .A(_777_),
    .B(_745_),
    .C(_914_),
    .Y(_778_)
);

NAND2X1 _1803_ (
    .A(ABCmd_i[6]),
    .B(_778_),
    .Y(_779_)
);

OAI21X1 _1804_ (
    .A(_759_),
    .B(_779_),
    .C(_765_),
    .Y(HC)
);

INVX1 _1805_ (
    .A(_775_),
    .Y(_780_)
);

NOR2X1 _1806_ (
    .A(_780_),
    .B(HC),
    .Y(_781_)
);

NOR2X1 _1807_ (
    .A(_776_),
    .B(_781_),
    .Y(ACC[4])
);

INVX1 _1808_ (
    .A(_774_),
    .Y(_782_)
);

NAND2X1 _1809_ (
    .A(ABCmd_i[5]),
    .B(AI[6]),
    .Y(_783_)
);

AND2X2 _1810_ (
    .A(_869_),
    .B(BI[5]),
    .Y(_784_)
);

NAND2X1 _1811_ (
    .A(AI[5]),
    .B(_784_),
    .Y(_785_)
);

AOI22X1 _1812_ (
    .A(_867_),
    .B(BI[5]),
    .C(_785_),
    .D(_868_),
    .Y(_786_)
);

OAI21X1 _1813_ (
    .A(AI[5]),
    .B(_784_),
    .C(_873_),
    .Y(_787_)
);

OAI21X1 _1814_ (
    .A(_787_),
    .B(_786_),
    .C(_783_),
    .Y(_788_)
);

OAI21X1 _1815_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[5]),
    .C(_863_),
    .Y(_789_)
);

AOI21X1 _1816_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[5]),
    .C(_789_),
    .Y(_790_)
);

OAI21X1 _1817_ (
    .A(_882_),
    .B(_790_),
    .C(_788_),
    .Y(_791_)
);

OAI21X1 _1818_ (
    .A(_788_),
    .B(_790_),
    .C(_791_),
    .Y(_792_)
);

OAI21X1 _1819_ (
    .A(_782_),
    .B(_776_),
    .C(_792_),
    .Y(_793_)
);

AOI21X1 _1820_ (
    .A(HC),
    .B(_780_),
    .C(_782_),
    .Y(_794_)
);

INVX1 _1821_ (
    .A(_792_),
    .Y(_795_)
);

NAND2X1 _1822_ (
    .A(_795_),
    .B(_794_),
    .Y(_796_)
);

NAND2X1 _1823_ (
    .A(_793_),
    .B(_796_),
    .Y(ACC[5])
);

OAI21X1 _1824_ (
    .A(_792_),
    .B(_794_),
    .C(_791_),
    .Y(_797_)
);

INVX1 _1825_ (
    .A(\u_ALU8.AI7 ),
    .Y(_798_)
);

AND2X2 _1826_ (
    .A(_869_),
    .B(BI[6]),
    .Y(_799_)
);

NAND2X1 _1827_ (
    .A(AI[6]),
    .B(_799_),
    .Y(_800_)
);

AOI22X1 _1828_ (
    .A(_867_),
    .B(BI[6]),
    .C(_800_),
    .D(_868_),
    .Y(_801_)
);

OAI21X1 _1829_ (
    .A(AI[6]),
    .B(_799_),
    .C(_873_),
    .Y(_802_)
);

OAI22X1 _1830_ (
    .A(_873_),
    .B(_798_),
    .C(_802_),
    .D(_801_),
    .Y(_803_)
);

OAI21X1 _1831_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI[6]),
    .C(_863_),
    .Y(_804_)
);

AOI21X1 _1832_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(BI[6]),
    .C(_804_),
    .Y(_805_)
);

OAI21X1 _1833_ (
    .A(_882_),
    .B(_805_),
    .C(_803_),
    .Y(_806_)
);

OAI21X1 _1834_ (
    .A(_803_),
    .B(_805_),
    .C(_806_),
    .Y(_807_)
);

NAND2X1 _1835_ (
    .A(_807_),
    .B(_797_),
    .Y(_808_)
);

OAI21X1 _1836_ (
    .A(_782_),
    .B(_776_),
    .C(_795_),
    .Y(_809_)
);

INVX1 _1837_ (
    .A(_807_),
    .Y(_810_)
);

NAND3X1 _1838_ (
    .A(_791_),
    .B(_810_),
    .C(_809_),
    .Y(_811_)
);

NAND2X1 _1839_ (
    .A(_811_),
    .B(_808_),
    .Y(ACC[6])
);

INVX1 _1840_ (
    .A(_806_),
    .Y(_812_)
);

AOI21X1 _1841_ (
    .A(_809_),
    .B(_791_),
    .C(_807_),
    .Y(_813_)
);

NAND2X1 _1842_ (
    .A(ABCmd_i[5]),
    .B(ABCmd_i[4]),
    .Y(_814_)
);

AND2X2 _1843_ (
    .A(_869_),
    .B(BI[7]),
    .Y(_815_)
);

NAND2X1 _1844_ (
    .A(\u_ALU8.AI7 ),
    .B(_815_),
    .Y(_816_)
);

AOI22X1 _1845_ (
    .A(_867_),
    .B(BI[7]),
    .C(_816_),
    .D(_868_),
    .Y(_817_)
);

OAI21X1 _1846_ (
    .A(\u_ALU8.AI7 ),
    .B(_815_),
    .C(_873_),
    .Y(_818_)
);

OAI21X1 _1847_ (
    .A(_818_),
    .B(_817_),
    .C(_814_),
    .Y(_819_)
);

OAI21X1 _1848_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[7]),
    .C(_863_),
    .Y(_820_)
);

AOI21X1 _1849_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[7]),
    .C(_820_),
    .Y(_821_)
);

OAI21X1 _1850_ (
    .A(_882_),
    .B(_821_),
    .C(_819_),
    .Y(_822_)
);

OAI21X1 _1851_ (
    .A(_819_),
    .B(_821_),
    .C(_822_),
    .Y(_823_)
);

OAI21X1 _1852_ (
    .A(_812_),
    .B(_813_),
    .C(_823_),
    .Y(_824_)
);

NAND2X1 _1853_ (
    .A(_810_),
    .B(_797_),
    .Y(_825_)
);

INVX1 _1854_ (
    .A(_823_),
    .Y(_826_)
);

NAND3X1 _1855_ (
    .A(_806_),
    .B(_826_),
    .C(_825_),
    .Y(_827_)
);

NAND2X1 _1856_ (
    .A(_827_),
    .B(_824_),
    .Y(AN)
);

NOR2X1 _1857_ (
    .A(ACC[0]),
    .B(_778_),
    .Y(_828_)
);

NAND2X1 _1858_ (
    .A(_759_),
    .B(_828_),
    .Y(_829_)
);

NOR2X1 _1859_ (
    .A(_829_),
    .B(ACC[4]),
    .Y(_830_)
);

INVX1 _1860_ (
    .A(ACC[5]),
    .Y(_831_)
);

NAND3X1 _1861_ (
    .A(_811_),
    .B(_808_),
    .C(_831_),
    .Y(_832_)
);

NOR2X1 _1862_ (
    .A(_832_),
    .B(AN),
    .Y(_833_)
);

AND2X2 _1863_ (
    .A(_833_),
    .B(_830_),
    .Y(AZ)
);

NAND3X1 _1864_ (
    .A(_806_),
    .B(_823_),
    .C(_825_),
    .Y(_834_)
);

OAI21X1 _1865_ (
    .A(_812_),
    .B(_813_),
    .C(_826_),
    .Y(_835_)
);

NAND2X1 _1866_ (
    .A(_834_),
    .B(_835_),
    .Y(_836_)
);

OAI21X1 _1867_ (
    .A(ACC[5]),
    .B(ACC[6]),
    .C(ABCmd_i[6]),
    .Y(_837_)
);

NOR2X1 _1868_ (
    .A(_875_),
    .B(_873_),
    .Y(_838_)
);

OAI21X1 _1869_ (
    .A(_806_),
    .B(_823_),
    .C(_822_),
    .Y(_839_)
);

INVX1 _1870_ (
    .A(_839_),
    .Y(_840_)
);

NAND3X1 _1871_ (
    .A(_810_),
    .B(_826_),
    .C(_797_),
    .Y(_841_)
);

NAND3X1 _1872_ (
    .A(_838_),
    .B(_840_),
    .C(_841_),
    .Y(_842_)
);

INVX1 _1873_ (
    .A(_838_),
    .Y(_843_)
);

NAND2X1 _1874_ (
    .A(_826_),
    .B(_810_),
    .Y(_844_)
);

AOI21X1 _1875_ (
    .A(_809_),
    .B(_791_),
    .C(_844_),
    .Y(_845_)
);

OAI21X1 _1876_ (
    .A(_839_),
    .B(_845_),
    .C(_843_),
    .Y(_846_)
);

AND2X2 _1877_ (
    .A(_846_),
    .B(_842_),
    .Y(_847_)
);

OAI21X1 _1878_ (
    .A(_836_),
    .B(_837_),
    .C(_847_),
    .Y(CO)
);

NAND3X1 _1879_ (
    .A(ABCmd_i[6]),
    .B(_832_),
    .C(AN),
    .Y(_848_)
);

INVX1 _1880_ (
    .A(_821_),
    .Y(_849_)
);

NAND2X1 _1881_ (
    .A(_882_),
    .B(_819_),
    .Y(_850_)
);

AOI21X1 _1882_ (
    .A(_850_),
    .B(_849_),
    .C(_798_),
    .Y(_851_)
);

NAND2X1 _1883_ (
    .A(_849_),
    .B(_850_),
    .Y(_852_)
);

NOR2X1 _1884_ (
    .A(\u_ALU8.AI7 ),
    .B(_852_),
    .Y(_853_)
);

NOR2X1 _1885_ (
    .A(_851_),
    .B(_853_),
    .Y(_854_)
);

NAND3X1 _1886_ (
    .A(_827_),
    .B(_854_),
    .C(_824_),
    .Y(_855_)
);

INVX1 _1887_ (
    .A(_854_),
    .Y(_856_)
);

NAND3X1 _1888_ (
    .A(_834_),
    .B(_856_),
    .C(_835_),
    .Y(_857_)
);

NAND2X1 _1889_ (
    .A(_855_),
    .B(_857_),
    .Y(_858_)
);

NAND3X1 _1890_ (
    .A(_847_),
    .B(_848_),
    .C(_858_),
    .Y(_859_)
);

AND2X2 _1891_ (
    .A(_855_),
    .B(_857_),
    .Y(_860_)
);

NAND2X1 _1892_ (
    .A(CO),
    .B(_860_),
    .Y(_861_)
);

NAND2X1 _1893_ (
    .A(_859_),
    .B(_861_),
    .Y(AV)
);

BUFX2 _1894_ (
    .A(_924_[0]),
    .Y(ACC_o[0])
);

BUFX2 _1895_ (
    .A(_924_[1]),
    .Y(ACC_o[1])
);

BUFX2 _1896_ (
    .A(_924_[2]),
    .Y(ACC_o[2])
);

BUFX2 _1897_ (
    .A(_924_[3]),
    .Y(ACC_o[3])
);

BUFX2 _1898_ (
    .A(_924_[4]),
    .Y(ACC_o[4])
);

BUFX2 _1899_ (
    .A(_924_[5]),
    .Y(ACC_o[5])
);

BUFX2 _1900_ (
    .A(_924_[6]),
    .Y(ACC_o[6])
);

BUFX2 _1901_ (
    .A(_924_[7]),
    .Y(ACC_o[7])
);

BUFX2 _1902_ (
    .A(_925_),
    .Y(Done_o)
);

INVX1 _927_ (
    .A(state[2]),
    .Y(_717_)
);

NOR2X1 _928_ (
    .A(state[0]),
    .B(_717_),
    .Y(_718_)
);

NAND2X1 _929_ (
    .A(state[1]),
    .B(_718_),
    .Y(_719_)
);

INVX1 _930_ (
    .A(_719_),
    .Y(_925_)
);

INVX1 _931_ (
    .A(state[0]),
    .Y(_720_)
);

INVX2 _932_ (
    .A(state[1]),
    .Y(_721_)
);

NOR2X1 _933_ (
    .A(state[2]),
    .B(_721_),
    .Y(_722_)
);

NAND2X1 _934_ (
    .A(_720_),
    .B(_722_),
    .Y(_723_)
);

INVX1 _935_ (
    .A(_723__bF$buf3),
    .Y(_724_)
);

NOR2X1 _936_ (
    .A(state[2]),
    .B(_720_),
    .Y(_725_)
);

AOI21X1 _937_ (
    .A(_721_),
    .B(_725_),
    .C(_925_),
    .Y(_726_)
);

NOR2X1 _938_ (
    .A(LoadCmd_i),
    .B(_726_),
    .Y(_727_)
);

OAI21X1 _939_ (
    .A(_724_),
    .B(_727_),
    .C(LoadB_i),
    .Y(_728_)
);

INVX1 _940_ (
    .A(LoadA_i),
    .Y(_729_)
);

INVX4 _941_ (
    .A(_718_),
    .Y(_730_)
);

OAI21X1 _942_ (
    .A(state[1]),
    .B(state[0]),
    .C(_717_),
    .Y(_731_)
);

INVX1 _943_ (
    .A(LoadB_i),
    .Y(_732_)
);

NOR2X1 _944_ (
    .A(state[1]),
    .B(_730_),
    .Y(_733_)
);

INVX1 _945_ (
    .A(_733_),
    .Y(_25_)
);

INVX1 _946_ (
    .A(LoadCmd_i),
    .Y(_26_)
);

OAI21X1 _947_ (
    .A(_725_),
    .B(_925_),
    .C(_26_),
    .Y(_27_)
);

OAI21X1 _948_ (
    .A(_732_),
    .B(_25_),
    .C(_27_),
    .Y(_28_)
);

AOI22X1 _949_ (
    .A(_730_),
    .B(_731_),
    .C(_28_),
    .D(_729_),
    .Y(_29_)
);

NAND2X1 _950_ (
    .A(_29_),
    .B(_728_),
    .Y(_926_[0])
);

OAI21X1 _951_ (
    .A(LoadA_i),
    .B(LoadB_i),
    .C(_26_),
    .Y(_30_)
);

OAI21X1 _952_ (
    .A(_30_),
    .B(_726_),
    .C(_25_),
    .Y(_31_)
);

NAND2X1 _953_ (
    .A(state[1]),
    .B(_725_),
    .Y(_32_)
);

NOR2X1 _954_ (
    .A(LoadA_i),
    .B(_26_),
    .Y(_33_)
);

NOR2X1 _955_ (
    .A(LoadB_i),
    .B(_26_),
    .Y(_34_)
);

OAI22X1 _956_ (
    .A(_33_),
    .B(_32__bF$buf3),
    .C(_723__bF$buf2),
    .D(_34_),
    .Y(_35_)
);

OR2X2 _957_ (
    .A(_31_),
    .B(_35_),
    .Y(_926_[1])
);

INVX1 _958_ (
    .A(_32__bF$buf2),
    .Y(_36_)
);

AOI22X1 _959_ (
    .A(_36_),
    .B(_33_),
    .C(_724_),
    .D(_34_),
    .Y(_37_)
);

NAND3X1 _960_ (
    .A(_729_),
    .B(_732_),
    .C(_733_),
    .Y(_38_)
);

AND2X2 _961_ (
    .A(_37_),
    .B(_38_),
    .Y(_39_)
);

OAI21X1 _962_ (
    .A(_26_),
    .B(_726_),
    .C(_39_),
    .Y(_926_[2])
);

INVX1 _963_ (
    .A(reset),
    .Y(_0_)
);

INVX1 _964_ (
    .A(ABCmd_i[0]),
    .Y(_40_)
);

NAND2X1 _965_ (
    .A(BI_0_bF$buf1),
    .B(_32__bF$buf1),
    .Y(_41_)
);

OAI21X1 _966_ (
    .A(_40_),
    .B(_32__bF$buf0),
    .C(_41_),
    .Y(_1_)
);

INVX1 _967_ (
    .A(ABCmd_i[1]),
    .Y(_42_)
);

NAND2X1 _968_ (
    .A(BI_1_bF$buf1),
    .B(_32__bF$buf3),
    .Y(_43_)
);

OAI21X1 _969_ (
    .A(_42_),
    .B(_32__bF$buf2),
    .C(_43_),
    .Y(_2_)
);

INVX1 _970_ (
    .A(ABCmd_i_2_bF$buf2),
    .Y(_44_)
);

NAND2X1 _971_ (
    .A(BI[2]),
    .B(_32__bF$buf1),
    .Y(_45_)
);

OAI21X1 _972_ (
    .A(_44_),
    .B(_32__bF$buf0),
    .C(_45_),
    .Y(_3_)
);

INVX1 _973_ (
    .A(ABCmd_i[3]),
    .Y(_46_)
);

NAND2X1 _974_ (
    .A(BI_3_bF$buf0),
    .B(_32__bF$buf3),
    .Y(_47_)
);

OAI21X1 _975_ (
    .A(_46_),
    .B(_32__bF$buf2),
    .C(_47_),
    .Y(_4_)
);

INVX1 _976_ (
    .A(ABCmd_i[4]),
    .Y(_48_)
);

NAND2X1 _977_ (
    .A(BI_4_bF$buf2),
    .B(_32__bF$buf1),
    .Y(_49_)
);

OAI21X1 _978_ (
    .A(_48_),
    .B(_32__bF$buf0),
    .C(_49_),
    .Y(_5_)
);

INVX1 _979_ (
    .A(ABCmd_i[5]),
    .Y(_50_)
);

NAND2X1 _980_ (
    .A(BI[5]),
    .B(_32__bF$buf3),
    .Y(_51_)
);

OAI21X1 _981_ (
    .A(_50_),
    .B(_32__bF$buf2),
    .C(_51_),
    .Y(_6_)
);

INVX1 _982_ (
    .A(ABCmd_i[6]),
    .Y(_52_)
);

NAND2X1 _983_ (
    .A(BI[6]),
    .B(_32__bF$buf1),
    .Y(_53_)
);

OAI21X1 _984_ (
    .A(_52_),
    .B(_32__bF$buf0),
    .C(_53_),
    .Y(_7_)
);

INVX4 _985_ (
    .A(ABCmd_i[7]),
    .Y(_54_)
);

NAND2X1 _986_ (
    .A(BI[7]),
    .B(_32__bF$buf3),
    .Y(_55_)
);

OAI21X1 _987_ (
    .A(_54_),
    .B(_32__bF$buf2),
    .C(_55_),
    .Y(_8_)
);

INVX1 _988_ (
    .A(_924_[0]),
    .Y(_56_)
);

INVX1 _989_ (
    .A(AI[0]),
    .Y(_57_)
);

INVX2 _990_ (
    .A(BI_3_bF$buf3),
    .Y(_58_)
);

NOR2X1 _991_ (
    .A(_57_),
    .B(_58_),
    .Y(_59_)
);

AND2X2 _992_ (
    .A(BI_4_bF$buf1),
    .B(AI[1]),
    .Y(_60_)
);

NAND2X1 _993_ (
    .A(_60_),
    .B(_59_),
    .Y(_61_)
);

NAND2X1 _994_ (
    .A(BI_1_bF$buf0),
    .B(AI[2]),
    .Y(_62_)
);

NAND2X1 _995_ (
    .A(BI_0_bF$buf0),
    .B(AI[3]),
    .Y(_63_)
);

OR2X2 _996_ (
    .A(_62_),
    .B(_63_),
    .Y(_64_)
);

NAND2X1 _997_ (
    .A(BI[2]),
    .B(AI[1]),
    .Y(_65_)
);

AND2X2 _998_ (
    .A(_62_),
    .B(_63_),
    .Y(_66_)
);

OAI21X1 _999_ (
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

endmodule
