* NGSPICE file created from fir_pe.ext - technology: scmos

.subckt NAND2X1 A B Y vdd gnd
M1000 a_26_14# A gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.600001p ps=16.2u
M1001 vdd B Y vdd pfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1002 Y B a_26_14# gnd nfet w=6u l=0.6u
+  ad=16.2p pd=17.400002u as=2.7p ps=6.9u
M1003 Y A vdd vdd pfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
.ends

.subckt OAI22X1 A B C D Y vdd gnd
M1000 Y D a_6_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1001 vdd C a_64_166# vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=5.4p ps=12.900001u
M1002 Y B a_24_166# vdd pfet w=12u l=0.6u
+  ad=23.400002p pd=15.900001u as=5.4p ps=12.900001u
M1003 gnd A a_6_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
M1004 a_64_166# D Y vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.900001u as=23.400002p ps=15.900001u
M1005 a_24_166# A vdd vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.900001u as=25.200003p ps=28.200003u
M1006 a_6_14# C Y gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1007 a_6_14# B gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
.ends

.subckt DFFPOSX1 D CLK Q vdd gnd
M1000 a_189_226# CLK a_165_14# vdd pfet w=3u l=0.6u
+  ad=0.9p pd=3.6u as=6.075p ps=8.400001u
M1001 a_87_10# a_59_14# vdd vdd pfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1002 a_59_14# CLK a_49_206# vdd pfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=5.4p ps=7.8u
M1003 a_87_10# a_59_14# gnd gnd nfet w=3u l=0.6u
+  ad=6.300001p pd=10.200001u as=4.05p ps=5.7u
M1004 a_165_14# a_11_14# a_161_206# vdd pfet w=6u l=0.6u
+  ad=6.075p pd=8.400001u as=1.8p ps=6.6u
M1005 gnd CLK a_11_14# gnd nfet w=6u l=0.6u
+  ad=5.85p pd=8.400001u as=12.600001p ps=16.2u
M1006 gnd a_87_10# a_81_14# gnd nfet w=3u l=0.6u
+  ad=4.05p pd=5.7u as=1.35p ps=3.9u
M1007 Q a_165_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=6.975p ps=8.700001u
M1008 a_157_14# a_87_10# gnd gnd nfet w=3u l=0.6u
+  ad=0.9p pd=3.6u as=6.300001p ps=10.200001u
M1009 vdd CLK a_11_14# vdd pfet w=12u l=0.6u
+  ad=11.250001p pd=14.400001u as=25.200003p ps=28.200003u
M1010 a_49_206# D vdd vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=11.250001p ps=14.400001u
M1011 vdd Q a_189_226# vdd pfet w=3u l=0.6u
+  ad=10.125001p pd=14.700001u as=0.9p ps=3.6u
M1012 a_165_14# CLK a_157_14# gnd nfet w=3u l=0.6u
+  ad=4.05p pd=5.7u as=0.9p ps=3.6u
M1013 a_49_14# D gnd gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=5.85p ps=8.400001u
M1014 a_85_206# a_11_14# a_59_14# vdd pfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=7.200001p ps=8.400001u
M1015 Q a_165_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=10.125001p ps=14.700001u
M1016 vdd a_87_10# a_85_206# vdd pfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=3.6p ps=7.2u
M1017 a_59_14# a_11_14# a_49_14# gnd nfet w=3u l=0.6u
+  ad=4.05p pd=5.7u as=1.35p ps=3.9u
M1018 a_161_206# a_87_10# vdd vdd pfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=12.600001p ps=16.2u
M1019 a_187_14# a_11_14# a_165_14# gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=4.05p ps=5.7u
M1020 gnd Q a_187_14# gnd nfet w=3u l=0.6u
+  ad=6.975p pd=8.700001u as=1.35p ps=3.9u
M1021 a_81_14# CLK a_59_14# gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=4.05p ps=5.7u
.ends

.subckt OAI21X1 A B C Y vdd gnd
M1000 Y C a_6_14# gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1001 Y B a_26_166# vdd pfet w=12u l=0.6u
+  ad=12.150001p pd=14.400001u as=9p ps=13.500001u
M1002 vdd C Y vdd pfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=12.150001p ps=14.400001u
M1003 gnd A a_6_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
M1004 a_6_14# B gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1005 a_26_166# A vdd vdd pfet w=12u l=0.6u
+  ad=9p pd=13.500001u as=25.200003p ps=28.200003u
.ends

.subckt INVX1 A Y vdd gnd
M1000 Y A gnd gnd nfet w=3u l=0.6u
+  ad=6.300001p pd=10.200001u as=6.300001p ps=10.200001u
M1001 Y A vdd vdd pfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=12.600001p ps=16.2u
.ends

.subckt XNOR2X1 A B Y vdd gnd
M1000 a_74_166# A Y vdd pfet w=12u l=0.6u
+  ad=3.6p pd=12.6u as=14.400002p ps=14.400001u
M1001 a_29_58# B vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=16.2p ps=14.700001u
M1002 gnd A a_6_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
M1003 vdd A a_6_14# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=25.200003p ps=28.200003u
M1004 Y A a_44_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=1.8p ps=6.6u
M1005 a_29_58# B gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=8.1p ps=8.700001u
M1006 vdd B a_74_166# vdd pfet w=12u l=0.6u
+  ad=16.2p pd=14.700001u as=3.6p ps=12.6u
M1007 Y a_6_14# a_44_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=5.4p ps=12.900001u
M1008 a_44_14# a_29_58# gnd gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=7.200001p ps=8.400001u
M1009 a_72_14# a_6_14# Y gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=7.200001p ps=8.400001u
M1010 a_44_166# a_29_58# vdd vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.900001u as=14.400002p ps=14.400001u
M1011 gnd B a_72_14# gnd nfet w=6u l=0.6u
+  ad=8.1p pd=8.700001u as=2.7p ps=6.9u
.ends

.subckt NOR2X1 A B Y vdd gnd
M1000 Y A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.300001p ps=10.200001u
M1001 a_24_166# A vdd vdd pfet w=12u l=0.6u
+  ad=9p pd=13.500001u as=25.200003p ps=28.200003u
M1002 gnd B Y gnd nfet w=3u l=0.6u
+  ad=6.300001p pd=10.200001u as=3.6p ps=5.4u
M1003 Y B a_24_166# vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=9p ps=13.500001u
.ends

.subckt NAND3X1 A B C Y vdd gnd
M1000 a_24_14# A gnd gnd nfet w=9u l=0.6u
+  ad=4.05p pd=9.900001u as=18.900002p ps=22.2u
M1001 vdd B Y vdd pfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1002 a_34_14# B a_24_14# gnd nfet w=9u l=0.6u
+  ad=6.750001p pd=10.500001u as=4.05p ps=9.900001u
M1003 Y C a_34_14# gnd nfet w=9u l=0.6u
+  ad=18.900002p pd=22.2u as=6.750001p ps=10.500001u
M1004 Y C vdd vdd pfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1005 Y A vdd vdd pfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
.ends

.subckt BUFX2 A Y vdd gnd
M1000 gnd A a_6_14# gnd nfet w=3u l=0.6u
+  ad=6.075p pd=8.400001u as=6.300001p ps=10.200001u
M1001 Y a_6_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=6.075p ps=8.400001u
M1002 Y a_6_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=12.150001p ps=14.400001u
M1003 vdd A a_6_14# vdd pfet w=6u l=0.6u
+  ad=12.150001p pd=14.400001u as=12.600001p ps=16.2u
.ends

.subckt AOI21X1 A B C Y vdd gnd
M1000 a_28_14# A gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.600001p ps=16.2u
M1001 Y C a_6_166# vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=14.400002p ps=14.400001u
M1002 Y B a_28_14# gnd nfet w=6u l=0.6u
+  ad=6.075p pd=8.400001u as=2.7p ps=6.9u
M1003 vdd A a_6_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=25.200003p ps=28.200003u
M1004 gnd C Y gnd nfet w=3u l=0.6u
+  ad=6.300001p pd=10.200001u as=6.075p ps=8.400001u
M1005 a_6_166# B vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
.ends

.subckt AOI22X1 A B C D Y vdd gnd
M1000 a_26_14# A gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.600001p ps=16.2u
M1001 Y D a_6_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1002 vdd A a_6_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=25.200003p ps=28.200003u
M1003 Y B a_26_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=2.7p ps=6.9u
M1004 a_56_14# D Y gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=7.200001p ps=8.400001u
M1005 a_6_166# C Y vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=14.400002p ps=14.400001u
M1006 a_6_166# B vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1007 gnd C a_56_14# gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=2.7p ps=6.9u
.ends

.subckt AND2X2 A B Y vdd gnd
M1000 a_24_14# A a_6_14# gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.600001p ps=16.2u
M1001 Y a_6_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=11.700001p ps=14.400001u
M1002 vdd B a_6_14# vdd pfet w=6u l=0.6u
+  ad=11.700001p pd=14.400001u as=7.200001p ps=8.400001u
M1003 gnd B a_24_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=2.7p ps=6.9u
M1004 Y a_6_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1005 a_6_14# A vdd vdd pfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
.ends

.subckt XOR2X1 A B Y vdd gnd
M1000 a_74_166# a_6_14# Y vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.900001u as=14.400002p ps=14.400001u
M1001 a_28_58# B vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=14.400002p ps=14.400001u
M1002 a_74_14# A Y gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=7.200001p ps=8.400001u
M1003 gnd A a_6_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
M1004 vdd A a_6_14# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=25.200003p ps=28.200003u
M1005 gnd B a_74_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=2.7p ps=6.9u
M1006 a_28_58# B gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1007 Y A a_44_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=5.4p ps=12.900001u
M1008 a_44_14# a_28_58# gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=7.200001p ps=8.400001u
M1009 vdd B a_74_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=5.4p ps=12.900001u
M1010 Y a_6_14# a_44_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=2.7p ps=6.9u
M1011 a_44_166# a_28_58# vdd vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.900001u as=14.400002p ps=14.400001u
.ends

.subckt OR2X2 A B Y vdd gnd
M1000 Y a_6_166# gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=6.300001p ps=8.400001u
M1001 vdd B a_24_166# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=5.4p ps=12.900001u
M1002 a_6_166# A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.300001p ps=10.200001u
M1003 a_24_166# A a_6_166# vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.900001u as=25.200003p ps=28.200003u
M1004 Y a_6_166# vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=14.400002p ps=14.400001u
M1005 gnd B a_6_166# gnd nfet w=3u l=0.6u
+  ad=6.300001p pd=8.400001u as=3.6p ps=5.4u
.ends

.subckt CLKBUF1 A Y vdd gnd
M1000 a_64_14# a_24_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1001 Y a_104_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1002 a_104_14# a_64_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1003 Y a_104_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1004 a_24_14# A gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
M1005 a_64_14# a_24_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1006 a_24_14# A vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=25.200003p ps=28.200003u
M1007 gnd a_24_14# a_64_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1008 a_104_14# a_64_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1009 gnd a_104_14# Y gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1010 vdd a_104_14# Y vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=14.400002p ps=14.400001u
M1011 gnd A a_24_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1012 vdd a_64_14# a_104_14# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1013 gnd a_64_14# a_104_14# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1014 vdd a_24_14# a_64_14# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1015 vdd A a_24_14# vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
.ends

.subckt INVX2 A Y vdd gnd
M1000 Y A gnd gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=12.600001p ps=16.2u
M1001 Y A vdd vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=25.200003p ps=28.200003u
.ends

.subckt INVX8 A Y vdd gnd
M1000 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1001 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=12.600001p ps=16.2u
M1002 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
M1003 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=25.200003p ps=28.200003u
M1004 gnd A Y gnd nfet w=6u l=0.6u
+  ad=12.600001p pd=16.2u as=7.200001p ps=8.400001u
M1005 gnd A Y gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=7.200001p ps=8.400001u
M1006 vdd A Y vdd pfet w=12u l=0.6u
+  ad=25.200003p pd=28.200003u as=14.400002p ps=14.400001u
M1007 vdd A Y vdd pfet w=12u l=0.6u
+  ad=14.400002p pd=14.400001u as=14.400002p ps=14.400001u
.ends

.subckt fir_pe gnd vdd Cin[5] Cin[4] Cin[3] Cin[2] Cin[1] Cin[0] Rdy Vld Xin[3] Xin[2]
+ Xin[1] Xin[0] Xout[3] Xout[2] Xout[1] Xout[0] Yin[3] Yin[2] Yin[1] Yin[0] Yout[3]
+ Yout[2] Yout[1] Yout[0] clk
X_1270_ _1270_/A _1270_/B _1275_/C vdd gnd NAND2X1
X_1399_ _738_/B _817_/A _1399_/C _1399_/D _1500_/D vdd gnd OAI22X1
X_1468_ _804_/Y _1508_/CLK _802_/A vdd gnd DFFPOSX1
X_981_ _985_/A _985_/B _984_/A _982_/C vdd gnd OAI21X1
X_1253_ _1257_/B _1254_/A vdd gnd INVX1
X_1322_ _1322_/A _1329_/A _1324_/B vdd gnd XNOR2X1
X_1184_ _1390_/C _1184_/B _1184_/C _1481_/D vdd gnd OAI21X1
X_964_ _969_/D _969_/C _965_/A vdd gnd NAND2X1
X_895_ _933_/D _895_/B _895_/C _904_/B vdd gnd OAI21X1
X_1305_ _1307_/A _1306_/A _1309_/A vdd gnd NOR2X1
X_1236_ _1236_/A _1236_/B _1483_/D vdd gnd NAND2X1
X_1167_ _1202_/B _1173_/B _1174_/C _1192_/A vdd gnd NAND3X1
X_1098_ _1212_/B _1098_/B _1099_/B vdd gnd NAND2X1
XBUFX2_insert0 _1526_/Q _841_/C vdd gnd BUFX2
X_947_ _947_/A _947_/B _947_/C _952_/A vdd gnd AOI21X1
X_878_ _878_/A _915_/C vdd gnd INVX1
X_1021_ _974_/A _1089_/C _1036_/B _1025_/A vdd gnd NAND3X1
X_1219_ _1356_/B _817_/A _1219_/C _1482_/D vdd gnd OAI21X1
X_732_ _732_/A _733_/B vdd gnd INVX1
X_801_ _813_/A _801_/B _801_/C _801_/Y vdd gnd OAI21X1
X_1004_ _990_/A Cin[2] _998_/Y _999_/Y _1010_/B vdd gnd AOI22X1
X_1484_ _1484_/D _1508_/CLK _1484_/Q vdd gnd DFFPOSX1
X_1398_ _810_/B _1402_/B _813_/A _1399_/C vdd gnd OAI21X1
X_1467_ _801_/Y _1509_/CLK _799_/A vdd gnd DFFPOSX1
X_980_ _980_/A Cin[4] _984_/A vdd gnd AND2X2
X_1321_ _1328_/B _1321_/B _1329_/A vdd gnd NOR2X1
X_1252_ _1252_/A _1252_/B _1252_/C _1254_/B vdd gnd AOI21X1
X_1183_ _1481_/Q _1390_/C _1184_/C vdd gnd NAND2X1
X_1519_ _1519_/D _1521_/CLK _977_/A vdd gnd DFFPOSX1
X_894_ _933_/C _894_/B _894_/C _904_/A vdd gnd NAND3X1
X_963_ _969_/A _969_/B _965_/B vdd gnd NAND2X1
X_1235_ _807_/A _1235_/B _1235_/C _1236_/B vdd gnd NAND3X1
X_1166_ _1193_/C _1169_/C _1169_/A _1202_/B vdd gnd NAND3X1
X_1304_ _1304_/A _1326_/C _1307_/A vdd gnd AND2X2
XBUFX2_insert1 _1526_/Q _816_/B vdd gnd BUFX2
X_1097_ _1480_/Q _1390_/C _1147_/C vdd gnd NAND2X1
X_946_ _946_/A _989_/B _989_/A _952_/B vdd gnd AOI21X1
X_877_ _877_/A _917_/A vdd gnd INVX1
X_1020_ _1020_/A _1020_/B _976_/Y _1036_/B vdd gnd OAI21X1
X_1149_ _1191_/A _1214_/B _1149_/C _1182_/A vdd gnd AOI21X1
X_1218_ _807_/A _1218_/B _1232_/C _1219_/C vdd gnd NAND3X1
X_731_ _743_/C _741_/A vdd gnd INVX1
X_800_ _813_/A _800_/B _801_/C vdd gnd NAND2X1
X_929_ _929_/A _929_/B _931_/C vdd gnd NAND2X1
X_1003_ _947_/C _1003_/B _946_/A _1078_/C vdd gnd OAI21X1
X_1483_ _1483_/D _1509_/CLK _1483_/Q vdd gnd DFFPOSX1
X_1535_ _745_/Y Yout[3] vdd gnd BUFX2
X_1397_ _808_/A _1401_/C _1399_/D vdd gnd NOR2X1
X_1466_ _798_/Y _1509_/CLK _796_/A vdd gnd DFFPOSX1
X_1320_ _1328_/C _1321_/B vdd gnd INVX1
X_1182_ _1182_/A _1214_/C _1184_/B vdd gnd XOR2X1
X_1251_ _1251_/A _1251_/B _1251_/C _1252_/C vdd gnd OAI21X1
X_1449_ _757_/A _979_/A _1449_/C _1520_/D vdd gnd OAI21X1
X_1518_ _1518_/D _1521_/CLK _922_/A vdd gnd DFFPOSX1
X_893_ _893_/A _893_/B _893_/C _904_/C vdd gnd AOI21X1
X_962_ _971_/A _971_/C _962_/C _969_/B vdd gnd NAND3X1
X_1303_ _781_/A _966_/A _1326_/C vdd gnd NAND2X1
X_1165_ _1165_/A _998_/B _1169_/C vdd gnd NOR2X1
X_1234_ _1241_/B _1234_/B _1235_/B vdd gnd NAND2X1
X_1096_ _967_/A _1096_/B _1096_/C _1479_/D vdd gnd OAI21X1
XBUFX2_insert2 _1526_/Q _813_/A vdd gnd BUFX2
X_945_ _951_/B _951_/C _952_/C _957_/B vdd gnd NAND3X1
X_876_ _876_/A _917_/B _876_/C _876_/D _876_/Y vdd gnd OAI22X1
X_1148_ _1214_/A _1149_/C vdd gnd INVX1
X_1079_ _987_/Y _1079_/B _1079_/C _1101_/C vdd gnd OAI21X1
X_1217_ _1217_/A _1252_/A _1217_/C _1232_/C vdd gnd OAI21X1
X_730_ _730_/A _730_/B _730_/C _730_/Y vdd gnd OAI21X1
X_928_ _928_/A _931_/B vdd gnd INVX1
X_1002_ _990_/A _994_/B _994_/A _992_/B _1003_/B vdd gnd AOI22X1
X_859_ _859_/A _859_/B _859_/C _879_/C vdd gnd OAI21X1
X_1482_ _1482_/D _1509_/CLK _1482_/Q vdd gnd DFFPOSX1
X_1465_ _795_/Y _1515_/CLK _793_/A vdd gnd DFFPOSX1
X_1534_ _741_/Y Yout[2] vdd gnd BUFX2
X_1396_ _1402_/B _1401_/C vdd gnd INVX1
X_1250_ _1251_/B _1252_/B vdd gnd INVX1
X_1181_ _1189_/A _1188_/A _1214_/C vdd gnd AND2X2
X_1448_ _748_/A Xin[2] _1449_/C vdd gnd NAND2X1
X_1517_ _1517_/D _1517_/CLK _776_/B vdd gnd DFFPOSX1
X_1379_ _1381_/A _1395_/A _1383_/A vdd gnd NOR2X1
X_961_ _961_/A _961_/B _961_/C _962_/C vdd gnd OAI21X1
X_892_ _905_/C _905_/B _905_/A _955_/B vdd gnd AOI21X1
X_1302_ _781_/A _966_/A _1304_/A vdd gnd OR2X2
X_1233_ _1233_/A _1242_/B _1241_/A _1234_/B vdd gnd OAI21X1
X_1095_ _1479_/Q _967_/A _1096_/C vdd gnd NAND2X1
X_1164_ _998_/B _1165_/A _1164_/C _1173_/B vdd gnd OAI21X1
XBUFX2_insert3 _1526_/Q _917_/B vdd gnd BUFX2
X_944_ _989_/A _989_/B _946_/A _951_/C vdd gnd NAND3X1
X_875_ _917_/B _878_/A _876_/D vdd gnd NAND2X1
X_1216_ _1233_/A _1217_/C vdd gnd INVX1
X_1078_ _1078_/A _995_/Y _1078_/C _1079_/B vdd gnd AOI21X1
X_1147_ _1390_/C _1147_/B _1147_/C _1480_/D vdd gnd OAI21X1
X_927_ _928_/A _927_/B _927_/C _950_/A vdd gnd NAND3X1
X_858_ _879_/B _879_/A _871_/C _868_/B vdd gnd NAND3X1
X_1001_ _995_/Y _1078_/A _989_/Y _1016_/B vdd gnd NAND3X1
X_789_ _789_/A _789_/B _789_/C _789_/Y vdd gnd OAI21X1
XCLKBUF1_insert10 clk _1522_/CLK vdd gnd CLKBUF1
X_1481_ _1481_/D _1515_/CLK _1481_/Q vdd gnd DFFPOSX1
X_1395_ _1395_/A _1395_/B _1395_/C _1402_/B vdd gnd AOI21X1
X_1464_ _792_/Y _1515_/CLK _790_/A vdd gnd DFFPOSX1
X_1533_ _736_/Y Yout[1] vdd gnd BUFX2
X_1180_ _1192_/B _1180_/B _1180_/C _1188_/A vdd gnd NAND3X1
X_1516_ _1516_/D _1521_/CLK _773_/B vdd gnd DFFPOSX1
X_1378_ _1384_/C _1378_/B _1381_/A vdd gnd AND2X2
X_1447_ _748_/A _924_/A _1447_/C _1519_/D vdd gnd OAI21X1
X_960_ _970_/A _970_/B _970_/C _971_/C vdd gnd NAND3X1
X_891_ _933_/D _895_/B _933_/C _905_/C vdd gnd OAI21X1
X_1232_ _1241_/A _1232_/B _1232_/C _1235_/C vdd gnd NAND3X1
X_1301_ _780_/B _917_/A _1301_/C _1306_/A vdd gnd OAI21X1
X_1094_ _1094_/A _1100_/A _1096_/B vdd gnd XOR2X1
X_1163_ _1193_/C _1169_/A _1164_/C vdd gnd NAND2X1
XBUFX2_insert4 _1526_/Q _789_/A vdd gnd BUFX2
X_874_ _874_/A _874_/B _874_/C _878_/A vdd gnd NAND3X1
X_943_ _943_/A _999_/B _988_/A _989_/B vdd gnd OAI21X1
X_1146_ _1191_/A _1187_/B _1147_/B vdd gnd XOR2X1
X_1215_ _1215_/A _1215_/B _1215_/C _1252_/A vdd gnd AOI21X1
X_1077_ _1101_/B _1101_/A _1085_/C _1091_/C vdd gnd NAND3X1
X_1000_ _999_/Y _996_/Y _998_/Y _1078_/A vdd gnd NAND3X1
X_857_ _893_/A _893_/B _881_/C _879_/B vdd gnd NAND3X1
X_788_ _789_/A _788_/B _789_/C vdd gnd NAND2X1
X_926_ _979_/A _985_/B _929_/A _927_/C vdd gnd OAI21X1
XCLKBUF1_insert11 clk _1509_/CLK vdd gnd CLKBUF1
X_1129_ _1129_/A _1129_/B _1129_/C _1130_/B vdd gnd AOI21X1
X_1480_ _1480_/D _1515_/CLK _1480_/Q vdd gnd DFFPOSX1
X_909_ _909_/A _910_/C vdd gnd INVX1
X_1532_ _730_/Y Yout[0] vdd gnd BUFX2
X_1394_ _1394_/A _1394_/B _1395_/B vdd gnd NOR2X1
X_1463_ _789_/Y _1517_/CLK _787_/A vdd gnd DFFPOSX1
X_1515_ _1515_/D _1515_/CLK _770_/B vdd gnd DFFPOSX1
X_1377_ _1392_/B _1384_/C vdd gnd INVX1
X_1446_ _748_/A Xin[1] _1447_/C vdd gnd NAND2X1
X_890_ _933_/A _988_/A _895_/B vdd gnd NOR2X1
X_1231_ _1241_/B _1232_/B vdd gnd INVX1
X_1300_ _735_/D _1310_/B _1309_/C vdd gnd NAND2X1
X_1162_ _759_/A _1225_/B _1162_/C _1169_/A vdd gnd OAI21X1
X_1093_ _1212_/B _1212_/A _1100_/A vdd gnd NAND2X1
XBUFX2_insert5 _1526_/Q _817_/A vdd gnd BUFX2
X_1429_ _1437_/B _1435_/B _1429_/C _1510_/D vdd gnd OAI21X1
X_873_ _874_/B _874_/C _874_/A _876_/C vdd gnd AOI21X1
X_942_ _942_/A _998_/A _946_/A vdd gnd NAND2X1
X_1214_ _1214_/A _1214_/B _1214_/C _1215_/C vdd gnd NAND3X1
X_1145_ _1214_/A _1214_/B _1187_/B vdd gnd NAND2X1
X_1076_ _1130_/C _1106_/A _1106_/B _1101_/A vdd gnd NAND3X1
X_925_ Cin[3] _985_/B vdd gnd INVX2
X_856_ _881_/B _893_/B vdd gnd INVX1
X_787_ _787_/A _789_/B vdd gnd INVX1
XCLKBUF1_insert12 clk _1521_/CLK vdd gnd CLKBUF1
X_1059_ _1120_/A _1113_/A vdd gnd INVX1
X_1128_ _1178_/A _1178_/B _1138_/C _1143_/A vdd gnd NAND3X1
X_908_ _912_/A _908_/B _908_/C _969_/D vdd gnd NAND3X1
X_839_ _839_/A _874_/A vdd gnd INVX1
X_1462_ _786_/Y _1479_/CLK _784_/A vdd gnd DFFPOSX1
X_1531_ _757_/Y Xout[3] vdd gnd BUFX2
X_1393_ _1393_/A _1395_/C vdd gnd INVX1
X_1445_ _748_/A _901_/A _1445_/C _1518_/D vdd gnd OAI21X1
X_1514_ _1514_/D _1515_/CLK _767_/A vdd gnd DFFPOSX1
X_1376_ _804_/B _1376_/B _1392_/B vdd gnd NOR2X1
X_1092_ _1092_/A _1092_/B _1092_/C _1212_/B vdd gnd NAND3X1
X_1230_ _1239_/B _1239_/A _1241_/B vdd gnd XOR2X1
X_1161_ _1193_/A _1227_/B _1161_/C _1162_/C vdd gnd OAI21X1
XBUFX2_insert6 _1526_/Q _807_/A vdd gnd BUFX2
X_1428_ _728_/A _728_/B _779_/B _1429_/C vdd gnd OAI21X1
X_1359_ _1374_/B _1362_/A _1361_/B vdd gnd AND2X2
X_941_ _994_/A _993_/B _998_/A vdd gnd AND2X2
X_872_ _919_/B _909_/A _910_/B _874_/C vdd gnd NAND3X1
X_1213_ _969_/Y _1213_/B _1213_/C _1215_/A vdd gnd NAND3X1
X_1075_ _1075_/A _1133_/B _1075_/C _1106_/B vdd gnd OAI21X1
X_1144_ _1144_/A _1144_/B _1144_/C _1214_/B vdd gnd OAI21X1
X_924_ _924_/A _979_/B _929_/B _927_/B vdd gnd OAI21X1
X_855_ _865_/C _883_/A _881_/C vdd gnd NAND2X1
X_786_ _841_/C _786_/B _786_/C _786_/Y vdd gnd OAI21X1
XCLKBUF1_insert13 clk _1517_/CLK vdd gnd CLKBUF1
X_1127_ _1168_/B _1168_/A _1152_/C _1178_/B vdd gnd NAND3X1
X_1058_ _1120_/B _1133_/A _1120_/A _1129_/A vdd gnd OAI21X1
X_907_ _921_/B _955_/C _921_/A _912_/A vdd gnd NAND3X1
X_838_ _840_/C _840_/B _840_/A _839_/A vdd gnd NAND3X1
X_769_ _769_/A _771_/B vdd gnd INVX1
X_1392_ _1392_/A _1392_/B _1392_/C _1393_/A vdd gnd AOI21X1
X_1461_ _783_/Y _1479_/CLK _781_/A vdd gnd DFFPOSX1
X_1530_ _754_/Y Xout[2] vdd gnd BUFX2
X_1375_ _804_/B _1376_/B _1378_/B vdd gnd NAND2X1
X_1444_ _728_/A Xin[0] _1445_/C vdd gnd NAND2X1
X_1513_ _1513_/D _1517_/CLK _788_/B vdd gnd DFFPOSX1
X_1091_ _1102_/A _1091_/B _1091_/C _1092_/C vdd gnd NAND3X1
X_1160_ _997_/A Cin[4] _1227_/B vdd gnd NAND2X1
X_1427_ _765_/B _1435_/B vdd gnd INVX1
X_1358_ _1373_/B _1362_/A vdd gnd INVX1
X_1289_ _780_/B _917_/A _1291_/A vdd gnd NAND2X1
X_940_ _947_/C _989_/A vdd gnd INVX1
X_871_ _871_/A _871_/B _871_/C _910_/B vdd gnd OAI21X1
X_1212_ _1212_/A _1212_/B _1213_/B vdd gnd AND2X2
X_1143_ _1143_/A _1143_/B _1179_/A _1144_/B vdd gnd AOI21X1
X_1074_ _1129_/C _1129_/B _1129_/A _1130_/C vdd gnd NAND3X1
X_854_ _978_/A _884_/B _883_/A vdd gnd AND2X2
X_923_ _980_/A Cin[3] _929_/B vdd gnd AND2X2
X_785_ _841_/C _785_/B _786_/C vdd gnd NAND2X1
XCLKBUF1_insert14 clk _1508_/CLK vdd gnd CLKBUF1
X_1126_ _1133_/C _1132_/B _1168_/B vdd gnd NAND2X1
X_1057_ _997_/A _997_/B _755_/A _993_/B _1120_/B vdd gnd AOI22X1
X_906_ _955_/A _921_/B vdd gnd INVX1
X_837_ _847_/B _847_/A _859_/C _840_/B vdd gnd NAND3X1
X_768_ _817_/A _768_/B _768_/C _768_/Y vdd gnd OAI21X1
X_1109_ _994_/A Cin[4] _1150_/B vdd gnd AND2X2
X_1391_ _733_/B _1404_/A _1391_/C _1391_/D _1499_/D vdd gnd AOI22X1
X_1460_ _780_/Y _1479_/CLK _778_/A vdd gnd DFFPOSX1
X_1512_ _1512_/D _1517_/CLK _785_/B vdd gnd DFFPOSX1
X_1443_ _744_/A _1443_/B _1443_/C _1517_/D vdd gnd AOI21X1
X_1374_ _1374_/A _1374_/B _1374_/C _1395_/A vdd gnd OAI21X1
X_1090_ _1090_/A _1102_/C _1090_/C _1092_/B vdd gnd NAND3X1
X_1357_ _1357_/A _1372_/B _1373_/B vdd gnd NOR2X1
X_1426_ _1443_/B _1426_/B _1426_/C _1509_/D vdd gnd AOI21X1
X_1288_ _729_/D _1310_/B _1299_/C vdd gnd NAND2X1
X_870_ _879_/C _879_/B _879_/A _909_/A vdd gnd NAND3X1
X_1142_ _1142_/A _1179_/C _1142_/C _1144_/A vdd gnd AOI21X1
X_1211_ _1233_/A _1242_/B _1218_/B vdd gnd NAND2X1
X_999_ _999_/A _999_/B _999_/C _999_/Y vdd gnd OAI21X1
X_1073_ _1073_/A _1103_/B _1106_/A vdd gnd AND2X2
X_1409_ Yin[1] _1439_/B vdd gnd INVX1
X_853_ _881_/A _893_/A vdd gnd INVX1
X_784_ _784_/A _786_/B vdd gnd INVX1
X_922_ _922_/A Cin[5] _928_/A vdd gnd NAND2X1
X_1125_ _1133_/A _1133_/B _1132_/A _1152_/C vdd gnd OAI21X1
X_1056_ _994_/C _1195_/A _1133_/A vdd gnd NOR2X1
X_905_ _905_/A _905_/B _905_/C _955_/C vdd gnd NAND3X1
X_767_ _767_/A _817_/A _768_/C vdd gnd NAND2X1
X_836_ _924_/A _862_/B _836_/C _847_/B vdd gnd OAI21X1
X_1108_ _985_/A _1225_/B _1150_/D vdd gnd NOR2X1
X_1039_ _1079_/C _1040_/C vdd gnd INVX1
X_1390_ _1390_/A _1394_/A _1390_/C _1391_/D vdd gnd AOI21X1
X_819_ _977_/A _864_/A _826_/A vdd gnd NAND2X1
X_1442_ _744_/A _776_/B _1443_/C vdd gnd NOR2X1
X_1511_ _1511_/D _1517_/CLK _782_/B vdd gnd DFFPOSX1
X_1373_ _1373_/A _1373_/B _1374_/A vdd gnd NAND2X1
X_1425_ _800_/B _1426_/B _1426_/C vdd gnd NOR2X1
X_1356_ _798_/B _1356_/B _1372_/B vdd gnd NOR2X1
X_1287_ _1310_/B _1287_/B _1287_/C _1489_/D vdd gnd OAI21X1
X_1141_ _1141_/A _1144_/C vdd gnd INVX1
X_1072_ _1130_/A _1081_/B _1081_/A _1101_/B vdd gnd NAND3X1
X_998_ _998_/A _998_/B _998_/Y vdd gnd NAND2X1
X_1210_ _1241_/A _1241_/C _1233_/A vdd gnd NAND2X1
X_1408_ _1437_/B _1417_/B _1408_/C _1502_/D vdd gnd OAI21X1
X_1339_ _1339_/A _1352_/B vdd gnd INVX1
X_921_ _921_/A _921_/B _921_/C _961_/C vdd gnd AOI21X1
X_783_ _841_/C _783_/B _783_/C _783_/Y vdd gnd OAI21X1
X_852_ _881_/B _893_/C _881_/A _879_/A vdd gnd OAI21X1
X_1124_ _1150_/C _1150_/D _1168_/A vdd gnd XOR2X1
X_1055_ _755_/A _997_/B _1195_/A vdd gnd NAND2X1
X_904_ _904_/A _904_/B _904_/C _921_/A vdd gnd NAND3X1
X_766_ _766_/A _768_/B vdd gnd INVX1
X_835_ _980_/A _884_/B _836_/C vdd gnd NAND2X1
X_1038_ _1090_/A _1102_/A vdd gnd INVX1
X_1107_ Cin[5] _1225_/B vdd gnd INVX2
X_818_ _922_/A _831_/B _823_/A vdd gnd NAND2X1
X_749_ _994_/A _943_/A vdd gnd INVX1
X_1441_ _1523_/D _1441_/B _1441_/C _1516_/D vdd gnd AOI21X1
X_1510_ _1510_/D _1517_/CLK _779_/B vdd gnd DFFPOSX1
X_1372_ _1373_/A _1372_/B _1372_/C _1374_/C vdd gnd AOI21X1
X_1355_ _796_/A _1482_/Q _1357_/A vdd gnd NOR2X1
X_1424_ _1441_/B _1426_/B _1424_/C _1508_/D vdd gnd AOI21X1
X_1286_ _744_/B _1310_/B _1287_/C vdd gnd NAND2X1
X_997_ _997_/A _997_/B _998_/B vdd gnd AND2X2
X_1140_ _1141_/A _1177_/B _1140_/C _1214_/A vdd gnd NAND3X1
X_1071_ _1075_/A _1133_/B _1129_/C _1081_/A vdd gnd OAI21X1
X_1338_ _1354_/A _1342_/B vdd gnd INVX1
X_1407_ _803_/B _1417_/B _1408_/C vdd gnd NAND2X1
X_1269_ _1271_/B _1271_/A _1270_/B vdd gnd NOR2X1
X_920_ _971_/A _959_/A vdd gnd INVX1
X_851_ _980_/A _889_/B _978_/A _884_/B _881_/B vdd gnd AOI22X1
X_782_ _789_/A _782_/B _783_/C vdd gnd NAND2X1
X_1054_ _994_/A Cin[2] _1120_/A vdd gnd NAND2X1
X_1123_ _1152_/A _1168_/C _1152_/B _1178_/A vdd gnd OAI21X1
X_834_ _889_/B _862_/B vdd gnd INVX1
X_903_ _955_/B _921_/C _955_/A _908_/C vdd gnd OAI21X1
X_765_ _765_/A _765_/B _765_/C _765_/Y vdd gnd OAI21X1
X_1106_ _1106_/A _1106_/B _1106_/C _1138_/C vdd gnd AOI21X1
X_1037_ _986_/C _987_/A _1090_/A vdd gnd NAND2X1
X_817_ _817_/A _817_/Y vdd gnd INVX8
X_748_ _748_/A _759_/A _748_/C _748_/Y vdd gnd OAI21X1
X_1440_ _728_/A _773_/B _1441_/C vdd gnd NOR2X1
X_1371_ _723_/B _1404_/A _1383_/C vdd gnd NAND2X1
X_1423_ _797_/B _1426_/B _1424_/C vdd gnd NOR2X1
X_1285_ _1294_/B _1285_/B _1287_/B vdd gnd XOR2X1
X_1354_ _1354_/A _1354_/B _1354_/C _1374_/B vdd gnd AOI21X1
X_996_ _996_/A _996_/Y vdd gnd INVX1
X_1070_ _1070_/A _1070_/B _1120_/A _1133_/B vdd gnd AOI21X1
X_1337_ _1339_/A _1354_/A _1341_/A vdd gnd NOR2X1
X_1268_ _769_/A _821_/A _1271_/B vdd gnd NOR2X1
X_1406_ _1526_/D _743_/A _743_/C _1417_/B vdd gnd NAND3X1
X_1199_ _1223_/A _1224_/C _1199_/C _1223_/D vdd gnd OAI21X1
X_850_ _850_/A _933_/A _893_/C vdd gnd NOR2X1
X_781_ _781_/A _783_/B vdd gnd INVX1
X_1122_ _1122_/A _1132_/A _1152_/A vdd gnd NOR2X1
X_979_ _979_/A _979_/B _984_/B _982_/B vdd gnd OAI21X1
X_1053_ _998_/A _998_/B _999_/Y _996_/Y _1075_/C vdd gnd AOI22X1
X_833_ _977_/A _924_/A vdd gnd INVX1
X_764_ Xin[3] _765_/B _765_/C vdd gnd NAND2X1
X_902_ _902_/A _930_/C _902_/C _955_/A vdd gnd OAI21X1
X_1105_ _1130_/C _1106_/C vdd gnd INVX1
X_1036_ _974_/A _1036_/B _1036_/C _1087_/C vdd gnd AOI21X1
X_747_ _748_/A _922_/A _748_/C vdd gnd NAND2X1
X_816_ _816_/A _816_/B _816_/C _816_/Y vdd gnd OAI21X1
X_1019_ _1088_/B _1088_/C _1088_/A _1089_/C vdd gnd NAND3X1
X_1370_ _1370_/A _1370_/B _1370_/C _1497_/D vdd gnd OAI21X1
X_1499_ _1499_/D _1515_/CLK _732_/A vdd gnd DFFPOSX1
X_1422_ _1439_/B _1426_/B _1422_/C _1507_/D vdd gnd AOI21X1
X_1284_ _1294_/A _1293_/A _1285_/B vdd gnd NOR2X1
X_1353_ _1353_/A _1353_/B _1353_/C _1354_/C vdd gnd OAI21X1
XBUFX2_insert30 Cin[1] _994_/B vdd gnd BUFX2
X_995_ _996_/A _995_/B _995_/C _995_/Y vdd gnd NAND3X1
X_1405_ Yin[0] _1437_/B vdd gnd INVX1
X_1267_ _771_/B _1275_/B _1271_/A vdd gnd NOR2X1
X_1336_ _1336_/A _1353_/A _1339_/A vdd gnd AND2X2
X_1198_ _755_/A Cin[4] _1224_/C vdd gnd NAND2X1
X_780_ _917_/B _780_/B _780_/C _780_/Y vdd gnd OAI21X1
X_1121_ _1195_/A _1195_/B _1132_/A vdd gnd XOR2X1
X_978_ _978_/A Cin[3] _984_/B vdd gnd AND2X2
X_1052_ _1103_/B _1073_/A _1130_/A vdd gnd NAND2X1
X_1319_ _787_/A _1479_/Q _1328_/C vdd gnd NAND2X1
X_901_ _901_/A _979_/B _973_/A _902_/C vdd gnd OAI21X1
X_832_ _832_/A _865_/C _859_/C vdd gnd NAND2X1
X_763_ _999_/A _765_/B _763_/C _763_/Y vdd gnd OAI21X1
X_1104_ _1142_/C _1179_/A vdd gnd INVX1
X_1035_ _1089_/C _1036_/C vdd gnd INVX1
X_746_ _990_/A _759_/A vdd gnd INVX2
X_815_ _922_/A _864_/A _841_/C _816_/C vdd gnd NAND3X1
X_1018_ _974_/Y _1029_/B _1029_/A _1025_/B vdd gnd NAND3X1
X_729_ _744_/A _729_/B _765_/B _729_/D _730_/C vdd gnd AOI22X1
X_1498_ _1498_/D _1508_/CLK _723_/B vdd gnd DFFPOSX1
X_1421_ _794_/B _1426_/B _1422_/C vdd gnd NOR2X1
X_1352_ _1352_/A _1352_/B _1354_/B vdd gnd NOR2X1
X_1283_ _777_/B _876_/A _1293_/A vdd gnd NOR2X1
XBUFX2_insert20 _817_/Y _967_/A vdd gnd BUFX2
XBUFX2_insert31 Cin[1] _889_/B vdd gnd BUFX2
X_994_ _994_/A _994_/B _994_/C _995_/C vdd gnd NAND3X1
X_1335_ _790_/A _1480_/Q _1353_/A vdd gnd NAND2X1
X_1404_ _1404_/A _1404_/B _1404_/C _1501_/D vdd gnd OAI21X1
X_1266_ _821_/A _1275_/B vdd gnd INVX1
X_1197_ _765_/A _985_/B _1227_/B _1199_/C vdd gnd OAI21X1
X_977_ _977_/A Cin[5] _983_/A vdd gnd NAND2X1
X_1051_ _1051_/A _1051_/B _1103_/A _1103_/B vdd gnd NAND3X1
X_1120_ _1120_/A _1120_/B _1120_/C _1122_/A vdd gnd OAI21X1
X_1318_ _787_/A _1479_/Q _1328_/B vdd gnd NOR2X1
X_1249_ _1257_/B _1257_/A _1255_/C vdd gnd NOR2X1
X_831_ _980_/A _831_/B _865_/C vdd gnd AND2X2
X_900_ _977_/A Cin[3] _973_/A vdd gnd NAND2X1
X_762_ Xin[2] _765_/B _763_/C vdd gnd NAND2X1
X_1103_ _1103_/A _1103_/B _1142_/C vdd gnd NAND2X1
X_1034_ _1034_/A _1034_/B _1100_/B _1094_/A vdd gnd OAI21X1
X_814_ _814_/A _816_/A vdd gnd INVX1
X_745_ _745_/A _745_/B _745_/C _745_/Y vdd gnd OAI21X1
X_1017_ _1020_/A _1020_/B _1088_/C _1029_/B vdd gnd OAI21X1
X_728_ _728_/A _728_/B _765_/B vdd gnd NOR2X1
X_1497_ _1497_/D _1526_/CLK _743_/B vdd gnd DFFPOSX1
X_1420_ _1437_/B _1426_/B _1420_/C _1506_/D vdd gnd AOI21X1
X_1351_ _739_/B _1370_/A _1361_/C vdd gnd NAND2X1
X_1282_ _775_/A _845_/A _1294_/A vdd gnd NOR2X1
XBUFX2_insert21 _817_/Y _1310_/B vdd gnd BUFX2
XBUFX2_insert32 Cin[1] _997_/B vdd gnd BUFX2
X_993_ _997_/A _993_/B _994_/C vdd gnd NAND2X1
X_1334_ _790_/A _1480_/Q _1336_/A vdd gnd OR2X2
X_1403_ _1403_/A _1403_/B _1404_/B vdd gnd NAND2X1
X_1265_ _1370_/A _1265_/B _1265_/C _1486_/D vdd gnd OAI21X1
X_1196_ _943_/A _1225_/B _1222_/A vdd gnd NOR2X1
X_976_ _976_/A _976_/B _976_/C _976_/Y vdd gnd AOI21X1
X_1050_ _985_/A _979_/B _1050_/C _1051_/A vdd gnd OAI21X1
X_1248_ _1258_/A _1248_/B _1257_/B vdd gnd AND2X2
X_1317_ _786_/B _968_/Y _1317_/C _1322_/A vdd gnd OAI21X1
X_1179_ _1179_/A _1179_/B _1179_/C _1180_/C vdd gnd OAI21X1
X_830_ _977_/A _864_/A _832_/A vdd gnd AND2X2
X_761_ _943_/A _765_/B _761_/C _761_/Y vdd gnd OAI21X1
X_959_ _959_/A _959_/B _959_/C _969_/A vdd gnd NAND3X1
X_1102_ _1102_/A _1102_/B _1102_/C _1141_/A vdd gnd OAI21X1
X_1033_ _968_/Y _917_/B _1033_/C _1033_/D _1478_/D vdd gnd OAI22X1
X_744_ _744_/A _744_/B _765_/B _744_/D _745_/C vdd gnd AOI22X1
X_813_ _813_/A _813_/B _813_/C _813_/Y vdd gnd OAI21X1
X_1016_ _1016_/A _1016_/B _987_/Y _1020_/B vdd gnd AOI21X1
X_727_ _727_/A _728_/B vdd gnd INVX2
X_1496_ _1496_/D _1526_/CLK _739_/B vdd gnd DFFPOSX1
X_1281_ _1281_/A _1281_/B _1281_/C _1294_/B vdd gnd AOI21X1
X_1350_ _1404_/A _1350_/B _1350_/C _1495_/D vdd gnd OAI21X1
X_1479_ _1479_/D _1479_/CLK _1479_/Q vdd gnd DFFPOSX1
XBUFX2_insert22 _817_/Y _1324_/A vdd gnd BUFX2
XBUFX2_insert33 Cin[1] _831_/B vdd gnd BUFX2
X_992_ _997_/A _992_/B _999_/C _995_/B vdd gnd NAND3X1
X_1402_ _810_/B _1402_/B _813_/B _1403_/A vdd gnd OAI21X1
X_1264_ _729_/B _1370_/A _1265_/C vdd gnd NAND2X1
X_1333_ _1333_/A _1333_/B _1354_/A vdd gnd NAND2X1
X_1195_ _1195_/A _1195_/B _1202_/A vdd gnd OR2X2
XCLKBUF1_insert7 clk _1479_/CLK vdd gnd CLKBUF1
X_975_ _975_/A _976_/C vdd gnd INVX1
X_1178_ _1178_/A _1178_/B _1178_/C _1179_/B vdd gnd AOI21X1
X_1247_ _1247_/A _1257_/C _1247_/C _1248_/B vdd gnd OAI21X1
X_1316_ _1316_/A _1316_/B _1316_/C _1492_/D vdd gnd OAI21X1
X_760_ Xin[1] _765_/B _761_/C vdd gnd NAND2X1
X_1101_ _1101_/A _1101_/B _1101_/C _1102_/B vdd gnd AOI21X1
X_889_ _990_/A _889_/B _988_/A vdd gnd NAND2X1
X_1032_ _917_/B _1100_/B _1033_/C vdd gnd NAND2X1
X_958_ _961_/A _961_/B _970_/C _959_/C vdd gnd OAI21X1
X_812_ _813_/A _812_/B _813_/C vdd gnd NAND2X1
X_743_ _743_/A _743_/B _743_/C _745_/B vdd gnd OAI21X1
X_1015_ _1040_/B _1079_/C _1040_/A _1020_/A vdd gnd AOI21X1
X_726_ _743_/A _726_/B _743_/C _730_/B vdd gnd OAI21X1
X_1495_ _1495_/D _1526_/CLK _734_/B vdd gnd DFFPOSX1
X_1280_ _774_/B _843_/A _1281_/C vdd gnd NOR2X1
X_1478_ _1478_/D _1479_/CLK _968_/A vdd gnd DFFPOSX1
XBUFX2_insert23 _817_/Y _1404_/A vdd gnd BUFX2
X_991_ _994_/A _994_/B _999_/C vdd gnd NAND2X1
X_1401_ _808_/A _811_/A _1401_/C _1403_/B vdd gnd NAND3X1
X_1194_ _1221_/A _1204_/C vdd gnd INVX1
X_1332_ _1332_/A _1332_/B _1332_/C _1333_/B vdd gnd NAND3X1
X_1263_ _1263_/A _1271_/C _1265_/B vdd gnd NAND2X1
XCLKBUF1_insert8 clk _1526_/CLK vdd gnd CLKBUF1
X_974_ _974_/A _974_/Y vdd gnd INVX1
X_1315_ _841_/C _1317_/C _1316_/B vdd gnd NAND2X1
X_1246_ _1246_/A _1257_/C vdd gnd INVX1
X_1177_ _1179_/C _1177_/B _1177_/C _1189_/A vdd gnd NAND3X1
X_957_ _957_/A _957_/B _957_/C _961_/B vdd gnd AOI21X1
X_1031_ _1098_/B _969_/Y _1031_/C _1100_/B vdd gnd NAND3X1
X_888_ _895_/C _894_/B _894_/C _905_/B vdd gnd NAND3X1
X_1100_ _1100_/A _1100_/B _1215_/B _1191_/A vdd gnd OAI21X1
X_1229_ _1243_/B _1243_/A _1239_/B vdd gnd XNOR2X1
X_811_ _811_/A _813_/B vdd gnd INVX1
X_742_ _742_/A _742_/B _745_/A vdd gnd NOR2X1
X_1014_ _957_/C _1014_/B _975_/A _1088_/C vdd gnd OAI21X1
X_725_ _727_/A _744_/A _743_/C vdd gnd NOR2X1
X_1494_ _1494_/D _1526_/CLK _726_/B vdd gnd DFFPOSX1
X_1477_ _967_/Y _1479_/CLK _966_/A vdd gnd DFFPOSX1
XBUFX2_insert24 _817_/Y _1390_/C vdd gnd BUFX2
X_990_ _990_/A Cin[2] _996_/A vdd gnd NAND2X1
X_1331_ _1331_/A _1331_/B _1332_/A vdd gnd NOR2X1
X_1400_ _742_/B _1404_/A _1404_/C vdd gnd NAND2X1
X_1262_ _768_/B _816_/A _1263_/A vdd gnd NAND2X1
X_1193_ _1193_/A _1227_/B _1193_/C _1221_/A vdd gnd OAI21X1
X_1529_ _751_/Y Xout[1] vdd gnd BUFX2
X_973_ _973_/A _985_/C _973_/C _974_/A vdd gnd OAI21X1
XCLKBUF1_insert9 clk _1515_/CLK vdd gnd CLKBUF1
X_1314_ _1329_/B _1314_/B _1317_/C vdd gnd NAND2X1
X_1245_ _1247_/C _1245_/B _1258_/A vdd gnd OR2X2
X_1176_ _1192_/B _1180_/B _1177_/C vdd gnd NAND2X1
X_956_ _976_/B _975_/A _976_/A _961_/A vdd gnd AOI21X1
X_887_ _933_/C _895_/C vdd gnd INVX1
X_1030_ _1030_/A _1030_/B _1034_/A _1031_/C vdd gnd OAI21X1
X_1228_ _1246_/A _1228_/B _1243_/B vdd gnd AND2X2
X_1159_ _994_/A Cin[3] _1193_/A vdd gnd NAND2X1
X_810_ _813_/A _810_/B _810_/C _810_/Y vdd gnd OAI21X1
X_741_ _741_/A _741_/B _741_/C _741_/Y vdd gnd OAI21X1
X_939_ _947_/C _947_/A _947_/B _951_/B vdd gnd NAND3X1
X_1013_ _951_/C _951_/B _951_/A _1014_/B vdd gnd AOI21X1
X_724_ _742_/A _743_/A vdd gnd INVX2
X_1493_ _1493_/D _1522_/CLK _744_/D vdd gnd DFFPOSX1
X_1476_ _917_/Y _1479_/CLK _877_/A vdd gnd DFFPOSX1
XBUFX2_insert25 _1522_/Q _757_/A vdd gnd BUFX2
X_1261_ _1270_/A _1271_/C vdd gnd INVX1
X_1330_ _1330_/A _1332_/B _1330_/C _1333_/A vdd gnd AOI21X1
X_1192_ _1192_/A _1192_/B _1209_/B vdd gnd NAND2X1
X_1459_ _777_/Y _1479_/CLK _775_/A vdd gnd DFFPOSX1
X_1528_ _748_/Y Xout[0] vdd gnd BUFX2
X_972_ _980_/A Cin[4] _985_/C vdd gnd NAND2X1
X_1313_ _1329_/B _1314_/B _1316_/A vdd gnd NOR2X1
X_1244_ _999_/A _979_/B _1244_/C _1245_/B vdd gnd OAI21X1
X_1175_ _1175_/A _1175_/B _1175_/C _1180_/B vdd gnd NAND3X1
X_886_ _980_/A Cin[2] _933_/C vdd gnd NAND2X1
X_955_ _955_/A _955_/B _955_/C _970_/C vdd gnd OAI21X1
X_1158_ _1158_/A _1161_/C _1158_/C _1193_/C vdd gnd NAND3X1
X_1227_ _1247_/A _1227_/B _1246_/A vdd gnd OR2X2
X_1089_ _974_/Y _1089_/B _1089_/C _1092_/A vdd gnd OAI21X1
X_740_ _744_/A _740_/B _765_/B _740_/D _741_/C vdd gnd AOI22X1
X_869_ _902_/A _919_/B vdd gnd INVX1
X_1012_ _1088_/B _1088_/A _976_/Y _1029_/A vdd gnd NAND3X1
X_938_ _990_/A _994_/B _988_/B _947_/B vdd gnd NAND3X1
X_723_ _742_/A _723_/B _730_/A vdd gnd NOR2X1
X_1492_ _1492_/D _1522_/CLK _740_/D vdd gnd DFFPOSX1
X_1475_ _876_/Y _1479_/CLK _845_/A vdd gnd DFFPOSX1
XBUFX2_insert15 Cin[0] _864_/A vdd gnd BUFX2
XBUFX2_insert26 _1522_/Q _728_/A vdd gnd BUFX2
X_1260_ _768_/B _816_/A _1270_/A vdd gnd NOR2X1
X_1191_ _1191_/A _1191_/B _1217_/A _1242_/B vdd gnd AOI21X1
X_1527_ _807_/A Vld vdd gnd BUFX2
X_1389_ _1390_/A _1394_/A _1391_/C vdd gnd OR2X2
X_1458_ _774_/Y _1522_/CLK _772_/A vdd gnd DFFPOSX1
X_971_ _971_/A _971_/B _971_/C _971_/Y vdd gnd OAI21X1
X_1312_ _784_/A _968_/A _1329_/B vdd gnd XOR2X1
X_1243_ _1243_/A _1243_/B _1247_/C vdd gnd NAND2X1
X_1174_ _1174_/A _1174_/B _1174_/C _1175_/C vdd gnd OAI21X1
X_885_ _933_/D _894_/B vdd gnd INVX1
X_954_ _970_/A _970_/B _961_/C _959_/B vdd gnd NAND3X1
X_1226_ _1244_/C _1247_/A vdd gnd INVX1
X_1157_ _999_/A _985_/B _1157_/C _1161_/C vdd gnd OAI21X1
X_1088_ _1088_/A _1088_/B _1088_/C _1089_/B vdd gnd AOI21X1
X_799_ _799_/A _801_/B vdd gnd INVX1
X_1011_ _1079_/C _1040_/B _1040_/A _1088_/A vdd gnd NAND3X1
X_868_ _902_/A _868_/B _868_/C _874_/B vdd gnd NAND3X1
X_937_ _994_/A _992_/B _988_/B vdd gnd NAND2X1
X_1209_ _1209_/A _1209_/B _1241_/C vdd gnd OR2X2
X_1491_ _1491_/D _1522_/CLK _735_/D vdd gnd DFFPOSX1
X_1474_ _844_/Y _1479_/CLK _842_/A vdd gnd DFFPOSX1
XBUFX2_insert16 Cin[0] _884_/B vdd gnd BUFX2
XBUFX2_insert27 _1522_/Q _1523_/D vdd gnd BUFX2
X_1190_ _1251_/A _1217_/A vdd gnd INVX1
X_1457_ _771_/Y _1517_/CLK _769_/A vdd gnd DFFPOSX1
X_1526_ _1526_/D _1526_/CLK _1526_/Q vdd gnd DFFPOSX1
X_1388_ _1392_/A _1394_/A vdd gnd INVX1
X_970_ _970_/A _970_/B _970_/C _971_/B vdd gnd AOI21X1
X_1311_ _1331_/A _1311_/B _1326_/C _1314_/B vdd gnd OAI21X1
X_1173_ _1202_/B _1173_/B _1173_/C _1175_/B vdd gnd NAND3X1
X_1242_ _1251_/B _1242_/B _1251_/C _1257_/A vdd gnd OAI21X1
X_1509_ _1509_/D _1509_/CLK _800_/B vdd gnd DFFPOSX1
X_953_ _975_/A _976_/A _976_/B _970_/B vdd gnd NAND3X1
X_884_ _990_/A _884_/B _978_/A _889_/B _933_/D vdd gnd AOI22X1
X_1225_ _765_/A _1225_/B _1244_/C vdd gnd NOR2X1
X_1156_ _1157_/C _1223_/A _1158_/C vdd gnd OR2X2
X_1087_ _1087_/A _1087_/B _1087_/C _1212_/A vdd gnd OAI21X1
X_936_ _994_/A _992_/B _988_/A _947_/A vdd gnd NAND3X1
X_798_ _817_/A _798_/B _798_/C _798_/Y vdd gnd OAI21X1
X_867_ _871_/A _871_/B _879_/C _868_/C vdd gnd OAI21X1
X_1010_ _1010_/A _1010_/B _989_/Y _1040_/B vdd gnd OAI21X1
X_1208_ _1209_/B _1209_/A _1241_/A vdd gnd NAND2X1
X_1139_ _1142_/C _1179_/C _1142_/A _1177_/B vdd gnd NAND3X1
X_1490_ _1490_/D _1522_/CLK _729_/D vdd gnd DFFPOSX1
X_919_ _929_/A _919_/B _971_/A vdd gnd NAND2X1
X_1473_ _822_/Y _1517_/CLK _821_/A vdd gnd DFFPOSX1
XBUFX2_insert17 Cin[0] _992_/B vdd gnd BUFX2
XBUFX2_insert28 _1522_/Q _748_/A vdd gnd BUFX2
X_1387_ _1387_/A _1392_/C _1392_/A vdd gnd NOR2X1
X_1456_ _768_/Y _1526_/CLK _766_/A vdd gnd DFFPOSX1
X_1525_ _742_/A _1526_/CLK _1526_/D vdd gnd DFFPOSX1
X_1241_ _1241_/A _1241_/B _1241_/C _1251_/B vdd gnd NAND3X1
X_1310_ _740_/D _1310_/B _1316_/C vdd gnd NAND2X1
X_1172_ _1172_/A _1192_/A _1172_/C _1192_/B vdd gnd NAND3X1
X_1439_ _1523_/D _1439_/B _1439_/C _1515_/D vdd gnd AOI21X1
X_1508_ _1508_/D _1508_/CLK _797_/B vdd gnd DFFPOSX1
X_883_ _883_/A _942_/A _894_/C vdd gnd NAND2X1
X_952_ _952_/A _952_/B _952_/C _976_/B vdd gnd OAI21X1
X_1224_ _999_/A _1225_/B _1224_/C _1228_/B vdd gnd OAI21X1
X_1086_ _1090_/C _1102_/C _1090_/A _1087_/A vdd gnd AOI21X1
X_1155_ _997_/A Cin[3] _1223_/A vdd gnd NAND2X1
X_866_ _866_/A _866_/B _881_/A _871_/B vdd gnd AOI21X1
X_935_ _978_/A Cin[2] _947_/C vdd gnd NAND2X1
X_797_ _817_/A _797_/B _798_/C vdd gnd NAND2X1
X_1207_ _1207_/A _1207_/B _1209_/A vdd gnd AND2X2
X_1069_ _765_/A _999_/B _998_/B _1070_/B vdd gnd OAI21X1
X_1138_ _1138_/A _1138_/B _1138_/C _1142_/A vdd gnd OAI21X1
X_918_ _977_/A Cin[4] _929_/A vdd gnd AND2X2
X_849_ _978_/A _884_/B _933_/A vdd gnd NAND2X1
X_1472_ _816_/Y _1517_/CLK _814_/A vdd gnd DFFPOSX1
XBUFX2_insert18 Cin[0] _993_/B vdd gnd BUFX2
XBUFX2_insert29 _1522_/Q _744_/A vdd gnd BUFX2
X_1524_ _727_/A _1526_/CLK _742_/A vdd gnd DFFPOSX1
X_1386_ _807_/B _1386_/B _1392_/C vdd gnd NOR2X1
X_1455_ _765_/Y _1521_/CLK _755_/A vdd gnd DFFPOSX1
X_1240_ _1240_/A _1240_/B _1251_/C vdd gnd NOR2X1
X_1171_ _1174_/A _1174_/B _1173_/C _1172_/C vdd gnd OAI21X1
X_1507_ _1507_/D _1515_/CLK _794_/B vdd gnd DFFPOSX1
X_1438_ _1523_/D _770_/B _1439_/C vdd gnd NOR2X1
X_1369_ _743_/B _1370_/A _1370_/C vdd gnd NAND2X1
X_951_ _951_/A _951_/B _951_/C _975_/A vdd gnd NAND3X1
X_882_ _990_/A _889_/B _942_/A vdd gnd AND2X2
X_1223_ _1223_/A _1224_/C _1223_/C _1223_/D _1243_/A vdd gnd OAI22X1
X_1154_ _994_/A Cin[4] _1157_/C vdd gnd NAND2X1
X_1085_ _1085_/A _1085_/B _1085_/C _1090_/C vdd gnd OAI21X1
X_934_ _951_/A _952_/C vdd gnd INVX1
X_796_ _796_/A _798_/B vdd gnd INVX1
X_865_ _985_/A _999_/B _865_/C _866_/B vdd gnd OAI21X1
X_1206_ _1221_/A _1221_/B _1206_/C _1207_/B vdd gnd NAND3X1
X_1137_ _1178_/B _1178_/A _1178_/C _1179_/C vdd gnd NAND3X1
X_1068_ _999_/A _862_/B _1068_/C _1070_/A vdd gnd OAI21X1
X_917_ _917_/A _917_/B _917_/C _917_/D _917_/Y vdd gnd OAI22X1
X_779_ _841_/C _779_/B _780_/C vdd gnd NAND2X1
X_848_ _977_/A Cin[2] _881_/A vdd gnd NAND2X1
X_1471_ _813_/Y _1509_/CLK _811_/A vdd gnd DFFPOSX1
XBUFX2_insert19 _817_/Y _1370_/A vdd gnd BUFX2
X_1454_ _763_/Y _1521_/CLK _997_/A vdd gnd DFFPOSX1
X_1523_ _1523_/D _1526_/CLK _727_/A vdd gnd DFFPOSX1
X_1385_ _805_/A _1485_/Q _1387_/A vdd gnd NOR2X1
X_1170_ _1202_/B _1174_/B vdd gnd INVX1
X_1437_ _1523_/D _1437_/B _1437_/C _1514_/D vdd gnd AOI21X1
X_1506_ _1506_/D _1515_/CLK _791_/B vdd gnd DFFPOSX1
X_1368_ _1368_/A _1373_/A _1370_/B vdd gnd XOR2X1
X_1299_ _1310_/B _1299_/B _1299_/C _1490_/D vdd gnd OAI21X1
X_950_ _950_/A _973_/C _976_/A vdd gnd AND2X2
X_881_ _881_/A _881_/B _881_/C _905_/A vdd gnd OAI21X1
X_1153_ _759_/A _1225_/B _1158_/A vdd gnd NOR2X1
X_1222_ _1222_/A _1223_/C vdd gnd INVX1
X_1084_ _1101_/C _1101_/B _1101_/A _1102_/C vdd gnd NAND3X1
X_933_ _933_/A _988_/A _933_/C _933_/D _951_/A vdd gnd OAI22X1
X_864_ _864_/A _999_/B vdd gnd INVX1
X_795_ _816_/B _795_/B _795_/C _795_/Y vdd gnd OAI21X1
X_1067_ _1120_/C _1113_/B _1113_/A _1075_/A vdd gnd AOI21X1
X_1205_ _1221_/C _1206_/C vdd gnd INVX1
X_1136_ _1179_/A _1143_/B _1143_/A _1140_/C vdd gnd NAND3X1
X_916_ _917_/B _969_/C _917_/D vdd gnd NAND2X1
X_847_ _847_/A _847_/B _847_/C _871_/C vdd gnd AOI21X1
X_778_ _778_/A _780_/B vdd gnd INVX1
X_1119_ _1133_/C _1132_/B _1168_/C vdd gnd NOR2X1
X_1470_ _810_/Y _1508_/CLK _808_/A vdd gnd DFFPOSX1
X_1453_ _761_/Y _1521_/CLK _994_/A vdd gnd DFFPOSX1
X_1522_ Rdy _1522_/CLK _1522_/Q vdd gnd DFFPOSX1
X_1384_ _1394_/B _1384_/B _1384_/C _1390_/A vdd gnd OAI21X1
X_1436_ _1523_/D _767_/A _1437_/C vdd gnd NOR2X1
X_1367_ _1367_/A _1372_/C _1373_/A vdd gnd NOR2X1
X_1505_ _1505_/D _1509_/CLK _812_/B vdd gnd DFFPOSX1
X_1298_ _1301_/C _1298_/B _1299_/B vdd gnd NAND2X1
X_880_ _902_/A _880_/B _909_/A _908_/B vdd gnd OAI21X1
X_1221_ _1221_/A _1221_/B _1221_/C _1239_/A vdd gnd AOI21X1
X_1083_ _1091_/C _1091_/B _1102_/A _1087_/B vdd gnd AOI21X1
X_1152_ _1152_/A _1152_/B _1152_/C _1174_/C vdd gnd OAI21X1
X_1419_ _791_/B _1426_/B _1420_/C vdd gnd NOR2X1
X_863_ _978_/A _985_/A vdd gnd INVX2
X_932_ _973_/C _950_/A _957_/C vdd gnd NAND2X1
X_794_ _816_/B _794_/B _795_/C vdd gnd NAND2X1
X_1204_ _1221_/C _1204_/B _1204_/C _1207_/A vdd gnd OAI21X1
X_1066_ _996_/A _1066_/B _998_/Y _1129_/C vdd gnd OAI21X1
X_1135_ _1138_/A _1138_/B _1178_/C _1143_/B vdd gnd OAI21X1
X_915_ _969_/D _915_/B _915_/C _969_/C vdd gnd NAND3X1
X_846_ _922_/A Cin[3] _902_/A vdd gnd NAND2X1
X_777_ _917_/B _777_/B _777_/C _777_/Y vdd gnd OAI21X1
X_1049_ _990_/A Cin[3] _1050_/C vdd gnd NAND2X1
X_1118_ _1118_/A _1165_/A _1118_/C _1133_/C vdd gnd OAI21X1
X_829_ _859_/A _847_/A vdd gnd INVX1
X_1383_ _1383_/A _1383_/B _1383_/C _1498_/D vdd gnd OAI21X1
X_1452_ _759_/Y _1521_/CLK _990_/A vdd gnd DFFPOSX1
X_1521_ _1521_/D _1521_/CLK _978_/A vdd gnd DFFPOSX1
X_1504_ _1504_/D _1508_/CLK _809_/B vdd gnd DFFPOSX1
X_1366_ _1366_/A _1372_/C vdd gnd INVX1
X_1435_ _1443_/B _1435_/B _1435_/C _1513_/D vdd gnd OAI21X1
X_1297_ _1297_/A _1332_/C _1301_/C vdd gnd NAND2X1
X_1151_ _1175_/A _1172_/A vdd gnd INVX1
X_1220_ _1483_/Q _1370_/A _1236_/A vdd gnd NAND2X1
X_1082_ _1085_/A _1085_/B _1101_/C _1091_/B vdd gnd OAI21X1
X_1418_ _743_/A _741_/A _1426_/B vdd gnd NOR2X1
X_1349_ _734_/B _1370_/A _1350_/C vdd gnd NAND2X1
X_931_ _931_/A _931_/B _931_/C _973_/C vdd gnd NAND3X1
X_862_ _979_/A _862_/B _883_/A _866_/A vdd gnd OAI21X1
X_793_ _793_/A _795_/B vdd gnd INVX1
X_1134_ _1134_/A _1134_/B _1152_/B _1138_/B vdd gnd AOI21X1
X_1203_ _1221_/B _1204_/B vdd gnd INVX1
X_1065_ _994_/A _994_/B _997_/A _992_/B _1066_/B vdd gnd AOI22X1
X_914_ _969_/D _915_/B _915_/C _917_/C vdd gnd AOI21X1
X_845_ _845_/A _876_/A vdd gnd INVX1
X_776_ _789_/A _776_/B _777_/C vdd gnd NAND2X1
X_1117_ _765_/A _862_/B _1195_/B _1118_/C vdd gnd OAI21X1
X_1048_ _1048_/A _1150_/A _1103_/A vdd gnd NAND2X1
X_759_ _759_/A _765_/B _759_/C _759_/Y vdd gnd OAI21X1
X_828_ _859_/B _847_/C _859_/A _840_/A vdd gnd OAI21X1
X_1520_ _1520_/D _1521_/CLK _980_/A vdd gnd DFFPOSX1
X_1382_ _1394_/B _1384_/B _807_/A _1383_/B vdd gnd OAI21X1
X_1451_ _748_/A _985_/A _1451_/C _1521_/D vdd gnd OAI21X1
X_1503_ _1503_/D _1508_/CLK _806_/B vdd gnd DFFPOSX1
X_1296_ _1331_/B _1296_/B _1298_/B vdd gnd NAND2X1
X_1365_ _799_/A _1483_/Q _1366_/A vdd gnd NAND2X1
X_1434_ _1523_/D _728_/B _788_/B _1435_/C vdd gnd OAI21X1
X_1150_ _1150_/A _1150_/B _1150_/C _1150_/D _1175_/A vdd gnd AOI22X1
X_1081_ _1081_/A _1081_/B _1130_/A _1085_/B vdd gnd AOI21X1
X_1417_ _1443_/B _1417_/B _1417_/C _1505_/D vdd gnd OAI21X1
X_1348_ _1348_/A _1352_/A _1350_/B vdd gnd XOR2X1
X_1279_ _1324_/A _1279_/B _1279_/C _1488_/D vdd gnd OAI21X1
X_930_ _979_/A _985_/B _930_/C _931_/A vdd gnd OAI21X1
X_861_ _980_/A _979_/A vdd gnd INVX2
X_792_ _816_/B _792_/B _792_/C _792_/Y vdd gnd OAI21X1
X_1202_ _1202_/A _1202_/B _1202_/C _1221_/B vdd gnd NAND3X1
X_1064_ _1129_/B _1075_/C _1129_/A _1081_/B vdd gnd NAND3X1
X_1133_ _1133_/A _1133_/B _1133_/C _1134_/A vdd gnd OAI21X1
X_913_ _913_/A _913_/B _913_/C _915_/B vdd gnd OAI21X1
X_775_ _775_/A _777_/B vdd gnd INVX1
X_844_ _844_/A _844_/B _844_/Y vdd gnd AND2X2
X_1047_ _1047_/A _1051_/B vdd gnd INVX1
X_1116_ _997_/A Cin[2] _1195_/B vdd gnd NAND2X1
X_827_ _977_/A _831_/B _980_/A _864_/A _859_/B vdd gnd AOI22X1
X_758_ Xin[0] _765_/B _759_/C vdd gnd NAND2X1
X_1450_ _728_/A Xin[3] _1451_/C vdd gnd NAND2X1
X_1381_ _1381_/A _1394_/B vdd gnd INVX1
X_1433_ _1441_/B _1435_/B _1433_/C _1512_/D vdd gnd OAI21X1
X_1502_ _1502_/D _1515_/CLK _803_/B vdd gnd DFFPOSX1
X_1364_ _799_/A _1483_/Q _1367_/A vdd gnd NOR2X1
X_1295_ _1332_/C _1296_/B vdd gnd INVX1
X_1080_ _1106_/B _1130_/C _1106_/A _1085_/A vdd gnd AOI21X1
X_1347_ _1347_/A _1352_/A vdd gnd INVX1
X_1416_ _812_/B _1417_/B _1417_/C vdd gnd NAND2X1
X_1278_ _740_/B _1324_/A _1279_/C vdd gnd NAND2X1
X_860_ _881_/C _893_/B _893_/A _871_/A vdd gnd AOI21X1
X_791_ _816_/B _791_/B _792_/C vdd gnd NAND2X1
X_1201_ _1202_/A _1202_/B _1202_/C _1221_/C vdd gnd AOI21X1
X_989_ _989_/A _989_/B _989_/C _989_/Y vdd gnd AOI21X1
X_1063_ _1113_/A _1113_/B _1120_/C _1129_/B vdd gnd NAND3X1
X_1132_ _1132_/A _1132_/B _1134_/B vdd gnd NAND2X1
X_912_ _912_/A _913_/B vdd gnd INVX1
X_843_ _843_/A _967_/A _844_/B vdd gnd NAND2X1
X_774_ _789_/A _774_/B _774_/C _774_/Y vdd gnd OAI21X1
X_1046_ _1047_/A _1046_/B _1046_/C _1073_/A vdd gnd NAND3X1
X_1115_ _755_/A Cin[2] _1165_/A vdd gnd NAND2X1
X_826_ _826_/A _850_/A _847_/C vdd gnd NOR2X1
X_757_ _757_/A _765_/A _757_/C _757_/Y vdd gnd OAI21X1
X_1029_ _1029_/A _1029_/B _974_/Y _1030_/B vdd gnd AOI21X1
X_1380_ _1395_/A _1384_/B vdd gnd INVX1
X_809_ _813_/A _809_/B _810_/C vdd gnd NAND2X1
X_1363_ _1372_/B _1363_/B _1368_/A vdd gnd NOR2X1
X_1432_ _728_/A _728_/B _785_/B _1433_/C vdd gnd OAI21X1
X_1501_ _1501_/D _1509_/CLK _742_/B vdd gnd DFFPOSX1
X_1294_ _1294_/A _1294_/B _1294_/C _1332_/C vdd gnd OAI21X1
X_1346_ _1353_/B _1346_/B _1347_/A vdd gnd NOR2X1
X_1415_ Yin[3] _1443_/B vdd gnd INVX1
X_1277_ _1281_/A _1281_/B _1279_/B vdd gnd XNOR2X1
X_790_ _790_/A _792_/B vdd gnd INVX1
X_988_ _988_/A _988_/B _989_/C vdd gnd NOR2X1
X_1200_ _1223_/D _1222_/A _1202_/C vdd gnd XOR2X1
X_1131_ _1152_/C _1168_/B _1168_/A _1138_/A vdd gnd AOI21X1
X_1062_ _1120_/B _1113_/B vdd gnd INVX1
X_1329_ _1329_/A _1329_/B _1332_/B vdd gnd AND2X2
X_911_ _921_/A _955_/C _921_/B _913_/A vdd gnd AOI21X1
X_842_ _842_/A _843_/A vdd gnd INVX1
X_773_ _789_/A _773_/B _774_/C vdd gnd NAND2X1
X_1114_ _997_/A _997_/B _1118_/A vdd gnd NAND2X1
X_1045_ _759_/A _985_/B _1048_/A _1046_/C vdd gnd OAI21X1
X_756_ _757_/A _978_/A _757_/C vdd gnd NAND2X1
X_825_ _980_/A _831_/B _850_/A vdd gnd NAND2X1
X_1028_ _1036_/B _1089_/C _974_/A _1030_/A vdd gnd AOI21X1
X_808_ _808_/A _810_/B vdd gnd INVX1
X_739_ _743_/A _739_/B _739_/C _741_/B vdd gnd OAI21X1
X_1500_ _1500_/D _1509_/CLK _737_/A vdd gnd DFFPOSX1
X_1362_ _1362_/A _1374_/B _1363_/B vdd gnd NOR2X1
X_1293_ _1293_/A _1294_/C vdd gnd INVX1
X_1431_ _1439_/B _1435_/B _1431_/C _1511_/D vdd gnd OAI21X1
X_1345_ _1353_/C _1346_/B vdd gnd INVX1
X_1276_ _772_/A _842_/A _1281_/B vdd gnd XOR2X1
X_1414_ _1441_/B _1417_/B _1414_/C _1504_/D vdd gnd OAI21X1
X_987_ _987_/A _987_/B _987_/Y vdd gnd NAND2X1
X_1130_ _1130_/A _1130_/B _1130_/C _1178_/C vdd gnd OAI21X1
X_1061_ _998_/B _1068_/C _1120_/C vdd gnd NAND2X1
X_1259_ _1386_/B _1390_/C _1259_/C _1259_/D _1485_/D vdd gnd AOI22X1
X_1328_ _1328_/A _1328_/B _1328_/C _1330_/C vdd gnd OAI21X1
X_910_ _919_/B _910_/B _910_/C _913_/C vdd gnd AOI21X1
X_772_ _772_/A _774_/B vdd gnd INVX1
X_841_ _841_/A _874_/A _841_/C _844_/A vdd gnd OAI21X1
X_1113_ _1113_/A _1113_/B _1133_/A _1132_/B vdd gnd AOI21X1
X_1044_ _978_/A Cin[4] _1048_/A vdd gnd AND2X2
X_755_ _755_/A _765_/A vdd gnd INVX2
X_824_ _922_/A Cin[2] _859_/A vdd gnd NAND2X1
X_1027_ _959_/A _962_/C _1027_/C _1034_/A vdd gnd AOI21X1
X_738_ _743_/A _738_/B _739_/C vdd gnd NAND2X1
X_807_ _807_/A _807_/B _807_/C _807_/Y vdd gnd OAI21X1
X_1430_ _728_/A _728_/B _782_/B _1431_/C vdd gnd OAI21X1
X_1292_ _1297_/A _1331_/B vdd gnd INVX1
X_1361_ _1361_/A _1361_/B _1361_/C _1496_/D vdd gnd OAI21X1
X_1413_ _809_/B _1417_/B _1414_/C vdd gnd NAND2X1
X_1344_ _793_/A _1481_/Q _1353_/C vdd gnd NAND2X1
X_1275_ _771_/B _1275_/B _1275_/C _1281_/A vdd gnd OAI21X1
X_986_ _986_/A _986_/B _986_/C _987_/A vdd gnd NAND3X1
X_1060_ _755_/A _993_/B _1068_/C vdd gnd AND2X2
X_1258_ _1258_/A _816_/B _1259_/D vdd gnd AND2X2
X_1189_ _1189_/A _1189_/B _1251_/A vdd gnd NAND2X1
X_1327_ _784_/A _968_/A _1328_/A vdd gnd NAND2X1
X_840_ _840_/A _840_/B _840_/C _841_/A vdd gnd AOI21X1
X_771_ _789_/A _771_/B _771_/C _771_/Y vdd gnd OAI21X1
X_1112_ _1150_/C _1150_/D _1152_/B vdd gnd XNOR2X1
X_969_ _969_/A _969_/B _969_/C _969_/D _969_/Y vdd gnd AOI22X1
X_1043_ _985_/A _979_/B _1150_/A _1046_/B vdd gnd OAI21X1
X_823_ _823_/A _826_/A _840_/C vdd gnd NOR2X1
X_754_ _757_/A _999_/A _754_/C _754_/Y vdd gnd OAI21X1
X_1026_ _971_/C _1027_/C vdd gnd INVX1
X_806_ _807_/A _806_/B _807_/C vdd gnd NAND2X1
X_737_ _737_/A _738_/B vdd gnd INVX1
X_1009_ _995_/Y _1078_/C _1078_/A _1079_/C vdd gnd NAND3X1
X_1360_ _1362_/A _1374_/B _813_/A _1361_/A vdd gnd OAI21X1
X_1291_ _1291_/A _1326_/A _1297_/A vdd gnd AND2X2
X_1489_ _1489_/D _1522_/CLK _744_/B vdd gnd DFFPOSX1
X_1343_ _793_/A _1481_/Q _1353_/B vdd gnd NOR2X1
X_1412_ Yin[2] _1441_/B vdd gnd INVX1
X_1274_ _1324_/A _1274_/B _1274_/C _1487_/D vdd gnd OAI21X1
X_985_ _985_/A _985_/B _985_/C _986_/A vdd gnd OAI21X1
X_1326_ _1326_/A _1331_/A _1326_/C _1330_/A vdd gnd OAI21X1
X_1257_ _1257_/A _1257_/B _1257_/C _1259_/C vdd gnd AOI21X1
X_1188_ _1188_/A _1214_/A _1189_/B vdd gnd NAND2X1
X_770_ _789_/A _770_/B _771_/C vdd gnd NAND2X1
X_968_ _968_/A _968_/Y vdd gnd INVX1
X_1111_ _1150_/A _1150_/B _1111_/C _1150_/C vdd gnd AOI21X1
X_899_ Cin[4] _979_/B vdd gnd INVX2
X_1042_ _990_/A Cin[3] _1150_/A vdd gnd AND2X2
X_1309_ _1309_/A _1309_/B _1309_/C _1491_/D vdd gnd OAI21X1
X_822_ _967_/A _822_/B _822_/C _822_/Y vdd gnd OAI21X1
X_753_ _757_/A _980_/A _754_/C vdd gnd NAND2X1
X_1025_ _1025_/A _1025_/B _971_/Y _1098_/B vdd gnd NAND3X1
X_805_ _805_/A _807_/B vdd gnd INVX1
X_736_ _741_/A _736_/B _736_/C _736_/Y vdd gnd OAI21X1
X_1008_ _987_/B _987_/A _1040_/A vdd gnd AND2X2
X_1290_ _778_/A _877_/A _1326_/A vdd gnd NAND2X1
X_1488_ _1488_/D _1522_/CLK _740_/B vdd gnd DFFPOSX1
X_1273_ _735_/B _1324_/A _1274_/C vdd gnd NAND2X1
X_1342_ _1352_/B _1342_/B _1353_/A _1348_/A vdd gnd OAI21X1
X_1411_ _1439_/B _1417_/B _1411_/C _1503_/D vdd gnd OAI21X1
X_984_ _984_/A _984_/B _986_/C vdd gnd NAND2X1
X_1256_ _1485_/Q _1386_/B vdd gnd INVX1
X_1325_ _726_/B _1404_/A _1341_/C vdd gnd NAND2X1
X_1187_ _1187_/A _1187_/B _1191_/B vdd gnd NOR2X1
X_898_ _922_/A _901_/A vdd gnd INVX1
X_1110_ _990_/A Cin[4] _994_/A Cin[3] _1111_/C vdd gnd AOI22X1
X_967_ _967_/A _967_/B _967_/C _967_/Y vdd gnd OAI21X1
X_1041_ _980_/A Cin[5] _1047_/A vdd gnd NAND2X1
X_1239_ _1239_/A _1239_/B _1241_/A _1240_/B vdd gnd AOI21X1
X_1308_ _1331_/A _1311_/B _841_/C _1309_/B vdd gnd OAI21X1
X_752_ _997_/A _999_/A vdd gnd INVX2
X_821_ _821_/A _967_/A _822_/C vdd gnd NAND2X1
X_1024_ _969_/Y _1213_/C _1033_/D vdd gnd NOR2X1
X_735_ _744_/A _735_/B _765_/B _735_/D _736_/C vdd gnd AOI22X1
X_804_ _816_/B _804_/B _804_/C _804_/Y vdd gnd OAI21X1
X_1007_ _987_/Y _1016_/B _1016_/A _1088_/B vdd gnd NAND3X1
X_1487_ _1487_/D _1522_/CLK _735_/B vdd gnd DFFPOSX1
X_1410_ _806_/B _1417_/B _1411_/C vdd gnd NAND2X1
X_1272_ _1272_/A _1275_/C _1274_/B vdd gnd NAND2X1
X_1341_ _1341_/A _1341_/B _1341_/C _1494_/D vdd gnd OAI21X1
X_983_ _983_/A _986_/B vdd gnd INVX1
X_1255_ _1376_/B _807_/A _1255_/C _1255_/D _1484_/D vdd gnd OAI22X1
X_1186_ _1188_/A _1189_/A _1187_/A vdd gnd NAND2X1
X_1324_ _1324_/A _1324_/B _1324_/C _1493_/D vdd gnd OAI21X1
X_1040_ _1040_/A _1040_/B _1040_/C _1085_/C vdd gnd AOI21X1
X_897_ _977_/A Cin[4] _930_/C vdd gnd NAND2X1
X_966_ _966_/A _967_/A _967_/C vdd gnd NAND2X1
X_1238_ _1239_/A _1239_/B _1240_/A vdd gnd NOR2X1
X_1307_ _1307_/A _1331_/A vdd gnd INVX1
X_1169_ _1169_/A _1193_/C _1169_/C _1174_/A vdd gnd AOI21X1
X_820_ _823_/A _826_/A _822_/B vdd gnd XNOR2X1
X_751_ _757_/A _943_/A _751_/C _751_/Y vdd gnd OAI21X1
X_949_ _957_/C _957_/B _957_/A _970_/A vdd gnd NAND3X1
X_1023_ _1034_/B _971_/Y _1213_/C vdd gnd XNOR2X1
X_803_ _816_/B _803_/B _804_/C vdd gnd NAND2X1
X_734_ _743_/A _734_/B _734_/C _736_/B vdd gnd OAI21X1
X_1006_ _1010_/A _1010_/B _1078_/C _1016_/A vdd gnd OAI21X1
X_1486_ _1486_/D _1526_/CLK _729_/B vdd gnd DFFPOSX1
X_1340_ _1352_/B _1342_/B _817_/A _1341_/B vdd gnd OAI21X1
X_1271_ _1271_/A _1271_/B _1271_/C _1272_/A vdd gnd OAI21X1
X_1469_ _807_/Y _1508_/CLK _805_/A vdd gnd DFFPOSX1
X_982_ _983_/A _982_/B _982_/C _987_/B vdd gnd NAND3X1
X_1323_ _744_/D _1324_/A _1324_/C vdd gnd NAND2X1
X_1185_ _1482_/Q _1356_/B vdd gnd INVX1
X_1254_ _1254_/A _1254_/B _807_/A _1255_/D vdd gnd OAI21X1
X_965_ _965_/A _965_/B _967_/B vdd gnd XNOR2X1
X_896_ _904_/B _904_/A _904_/C _921_/C vdd gnd AOI21X1
X_1306_ _1306_/A _1311_/B vdd gnd INVX1
X_1237_ _1484_/Q _1376_/B vdd gnd INVX1
X_1168_ _1168_/A _1168_/B _1168_/C _1173_/C vdd gnd AOI21X1
X_1099_ _1212_/A _1099_/B _1215_/B vdd gnd NAND2X1
X_750_ _757_/A _977_/A _751_/C vdd gnd NAND2X1
X_948_ _952_/A _952_/B _951_/A _957_/A vdd gnd OAI21X1
X_879_ _879_/A _879_/B _879_/C _880_/B vdd gnd AOI21X1
X_1022_ _1025_/A _1025_/B _1034_/B vdd gnd NAND2X1
X_802_ _802_/A _804_/B vdd gnd INVX1
X_733_ _743_/A _733_/B _734_/C vdd gnd NAND2X1
X_1005_ _995_/B _995_/C _996_/A _1010_/A vdd gnd AOI21X1
X_1485_ _1485_/D _1508_/CLK _1485_/Q vdd gnd DFFPOSX1
.ends

