magic
tech scmos
magscale 1 2
timestamp 1727401709
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 22 14 26 74
rect 30 14 34 74
rect 38 14 42 74
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 60 206 64 246
<< ndiffusion >>
rect 20 14 22 74
rect 26 14 30 74
rect 34 14 38 74
rect 42 72 56 74
rect 42 14 44 72
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 210 46 246
rect 58 210 60 246
rect 44 206 60 210
rect 64 206 66 246
<< ndcontact >>
rect 8 14 20 74
rect 44 14 56 72
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 46 210 58 246
rect 66 206 78 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 194 24 206
rect 40 194 44 206
rect 10 190 24 194
rect 30 190 44 194
rect 10 163 16 190
rect 10 103 16 151
rect 30 149 36 190
rect 10 90 26 103
rect 22 74 26 90
rect 30 74 34 137
rect 60 103 64 206
rect 38 91 44 103
rect 56 91 64 103
rect 38 74 42 91
rect 22 10 26 14
rect 30 10 34 14
rect 38 10 42 14
<< polycontact >>
rect 4 151 16 163
rect 24 137 36 149
rect 44 91 56 103
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 6 246 18 252
rect 46 246 58 252
rect 28 204 38 206
rect 66 204 72 206
rect 28 198 72 204
rect 3 163 17 177
rect 66 157 72 198
rect 63 143 77 157
rect 23 123 37 137
rect 43 103 57 117
rect 66 81 72 143
rect 44 72 72 81
rect 56 70 72 72
rect 8 8 20 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 3 163 17 177
rect 63 143 77 157
rect 23 123 37 137
rect 43 103 57 117
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 23 123 37 137 0 B
port 1 nsew signal input
rlabel metal1 43 103 57 117 0 C
port 2 nsew signal input
rlabel metal1 63 143 77 157 0 Y
port 3 nsew signal output
rlabel metal1 3 163 17 177 0 A
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
