magic
tech scmos
magscale 1 6
timestamp 1721992760
<< checkpaint >>
rect -156 655 552 936
rect -213 378 552 655
rect 799 465 1500 936
rect 730 405 1500 465
rect -156 -144 552 378
rect 631 147 1500 405
rect 769 142 1500 147
rect 799 -144 1500 142
<< error_s >>
rect -387 762 1518 798
rect -387 -18 1518 18
<< polysilicon >>
rect -207 497 -141 534
rect -93 498 -25 535
rect 866 502 932 538
rect 750 462 816 498
<< polycontact >>
rect -243 497 -207 534
rect -25 498 11 535
rect 932 502 968 538
rect 714 462 750 498
<< metal1 >>
rect -387 756 1518 804
rect -363 366 -321 408
rect -233 366 -171 408
rect 1182 366 1201 438
rect -233 348 -211 366
rect 1290 348 1326 366
rect -291 306 -211 348
rect -99 324 48 342
rect 234 293 258 313
rect 78 261 226 285
rect 444 235 480 348
rect 537 318 606 340
rect 850 327 967 345
rect 1446 306 1488 348
rect 438 193 480 235
rect -385 -24 1518 24
<< m2contact >>
rect -249 534 -207 576
rect 649 558 691 600
rect 11 498 53 540
rect 510 498 552 540
rect 708 498 750 540
rect 932 538 974 580
rect 1170 438 1212 480
rect 126 366 168 408
rect 342 366 384 408
rect 1081 366 1123 408
rect 1290 366 1332 408
rect 1386 366 1428 408
rect 282 306 324 348
rect 226 251 268 293
rect 1021 306 1063 348
rect 1230 306 1272 348
<< metal2 >>
rect -207 558 649 576
rect 691 558 932 576
rect 53 498 510 516
rect 552 498 708 516
rect 150 462 1170 480
rect 150 408 168 462
rect 366 426 1099 444
rect 366 408 384 426
rect 1081 408 1099 426
rect 1152 389 1290 408
rect 1152 348 1170 389
rect 1332 389 1386 408
rect 176 319 282 337
rect 176 234 194 319
rect 1063 330 1170 348
rect 1230 288 1248 306
rect 268 267 788 285
rect 896 270 1248 288
rect -61 216 194 234
use INVX1  INVX1_0 ~/ETRI050_DesignKit/devel/digital_ETRI050_m1d
timestamp 1702308830
transform 1 0 588 0 1 0
box -39 -24 159 816
use INVX1  INVX1_1
timestamp 1702308830
transform 1 0 1380 0 1 0
box -39 -24 159 816
use INVX1  INVX1_2
timestamp 1702308830
transform 1 0 -369 0 1 0
box -39 -24 159 816
use INVX1  INVX1_3
timestamp 1702308830
transform 1 0 432 0 1 0
box -39 -24 159 816
use NAND2X1  NAND2X1_0 ~/ETRI050_DesignKit/devel/digital_ETRI050_m1d
timestamp 1721984330
transform 1 0 216 0 1 0
box -36 -24 216 816
use NAND2X1  NAND2X1_1
timestamp 1721984330
transform 1 0 1164 0 1 0
box -36 -24 216 816
use NAND2X1  NAND2X1_2
timestamp 1721984330
transform 1 0 0 0 1 0
box -36 -24 216 816
use NAND2X1  NAND2X1_3
timestamp 1721984330
transform 1 0 955 0 1 0
box -36 -24 216 816
use SWITCH2X1  SWITCH2X1_0
timestamp 1721969656
transform 1 0 -201 0 1 6
box -50 -30 216 810
use SWITCH2X1  SWITCH2X1_1
timestamp 1721969656
transform -1 0 926 0 1 6
box -50 -30 216 810
<< labels >>
rlabel metal1 438 193 480 235 0 CLK
port 3 nsew
rlabel metal1 1446 306 1488 348 0 Q
port 4 nsew
rlabel metal1 -363 366 -321 408 0 D
port 0 nsew
rlabel metal1 -387 756 1518 804 0 vdd
port 5 nsew
rlabel metal1 -385 -24 1518 24 0 gnd
port 6 nsew
rlabel metal1 566 330 566 330 0 C_Bar
rlabel space 676 367 676 367 0 C
rlabel metal1 -231 329 -231 329 0 D_Bar
rlabel m2contact 126 366 168 408 0 S
port 2 nsew
rlabel m2contact 342 366 384 408 0 R
port 1 nsew
<< end >>
