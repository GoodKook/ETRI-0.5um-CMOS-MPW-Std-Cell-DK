magic
tech scmos
magscale 1 2
timestamp 1728306572
<< nwell >>
rect -13 134 112 252
<< ntransistor >>
rect 21 14 25 54
rect 29 14 33 54
rect 51 14 55 34
<< ptransistor >>
rect 21 186 25 226
rect 41 186 45 226
rect 61 186 65 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 14 29 54
rect 33 14 35 54
rect 47 14 51 34
rect 55 14 57 34
<< pdiffusion >>
rect 19 186 21 226
rect 25 186 27 226
rect 39 186 41 226
rect 45 186 47 226
rect 59 186 61 226
rect 65 186 67 226
<< ndcontact >>
rect 7 14 19 54
rect 35 14 47 54
rect 57 14 69 34
<< pdcontact >>
rect 7 186 19 226
rect 27 186 39 226
rect 47 186 59 226
rect 67 186 79 226
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 234 106 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 61 226 65 230
rect 21 89 25 186
rect 16 77 25 89
rect 41 109 45 186
rect 61 182 65 186
rect 61 178 69 182
rect 41 97 44 109
rect 41 87 45 97
rect 21 54 25 77
rect 29 80 45 87
rect 29 54 33 80
rect 65 72 69 178
rect 57 60 69 72
rect 51 34 55 60
rect 21 10 25 14
rect 29 10 33 14
rect 51 10 55 14
<< polycontact >>
rect 4 77 16 89
rect 44 97 56 109
rect 45 60 57 72
<< metal1 >>
rect -6 246 106 248
rect -6 232 106 234
rect 7 226 19 232
rect 47 226 59 232
rect 28 69 35 186
rect 68 111 75 186
rect 7 60 45 69
rect 7 54 19 60
rect 68 42 75 97
rect 57 34 75 42
rect 35 8 47 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 3 89 17 103
rect 43 109 57 123
rect 63 97 77 111
<< metal2 >>
rect 43 123 57 137
rect 3 103 17 117
rect 63 83 77 97
<< m1p >>
rect -6 232 106 248
rect -6 -8 106 8
<< m2p >>
rect 43 123 57 137
rect 3 103 17 117
rect 63 83 77 97
<< labels >>
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 106 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal2 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal2 43 123 57 137 0 B
port 1 nsew signal input
rlabel metal2 63 83 77 97 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
