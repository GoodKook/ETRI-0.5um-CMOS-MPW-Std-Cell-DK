magic
tech scmos
magscale 1 30
timestamp 1771034720
<< checkpaint >>
rect 18300 370350 361700 370850
rect 9650 369850 370350 370350
rect 9150 360700 370350 369850
rect 9150 181835 370850 360700
rect 6771 175958 370850 181835
rect 205 160774 370850 175958
rect 6771 143081 370850 160774
rect 0 102896 370850 143081
rect -13866 102380 370850 102896
rect -25613 89180 370850 102380
rect -24170 89077 370850 89180
rect -17472 83925 370850 89077
rect 0 47900 370850 83925
rect 6771 31724 370850 47900
rect -4457 18300 370850 31724
rect -4457 9150 370350 18300
rect -4457 8670 185015 9150
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
use apple_1_WozMon_PIA_Core  apple_1_WozMon_PIA_Core_0
timestamp 1771034318
transform 1 0 63960 0 1 65430
box -930 -360 184230 180945
use IOFILLER18  IOFILLER18_0
timestamp 1725930584
transform 0 -1 360600 -1 0 76146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 360598 -1 0 62646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 360600 -1 0 103146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 360600 -1 0 89646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 360602 -1 0 130146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 360600 -1 0 116646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 74345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 101345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 128345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 19399 -1 0 76155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 19399 -1 0 62655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 19400 -1 0 103155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 19400 -1 0 89655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 74345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 19397 -1 0 116655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 19400 -1 0 130155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60845 0 -1 360601
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 101345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87844 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 128345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_24
timestamp 1725930584
transform 0 1 19400 -1 0 143655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_25
timestamp 1725930584
transform 0 1 19400 -1 0 157155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_26
timestamp 1725930584
transform 0 1 19400 -1 0 170655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_27
timestamp 1725930584
transform 0 1 19400 -1 0 184155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_28
timestamp 1725930584
transform 0 1 19400 -1 0 197655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_29
timestamp 1725930584
transform 0 1 19400 -1 0 211155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_30
timestamp 1725930584
transform 0 1 19400 -1 0 224655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_31
timestamp 1725930584
transform 0 1 19400 -1 0 238155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_32
timestamp 1725930584
transform 0 1 19400 -1 0 251655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_33
timestamp 1725930584
transform 0 1 19400 -1 0 265155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_34
timestamp 1725930584
transform 0 1 19400 -1 0 278655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_35
timestamp 1725930584
transform 0 1 19400 -1 0 292155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_36
timestamp 1725930584
transform 0 1 19400 -1 0 305655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_37
timestamp 1725930584
transform 0 1 19400 -1 0 319155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_38
timestamp 1725930584
transform 0 -1 360602 -1 0 143646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_39
timestamp 1725930584
transform 0 -1 360602 -1 0 157146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_40
timestamp 1725930584
transform 0 -1 360602 -1 0 170646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_41
timestamp 1725930584
transform 0 -1 360602 -1 0 184146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_42
timestamp 1725930584
transform 0 -1 360602 -1 0 197646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_43
timestamp 1725930584
transform 0 -1 360602 -1 0 211146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_44
timestamp 1725930584
transform 0 -1 360602 -1 0 224646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_45
timestamp 1725930584
transform 0 -1 360602 -1 0 238146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_46
timestamp 1725930584
transform 0 -1 360602 -1 0 251646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_47
timestamp 1725930584
transform 0 -1 360602 -1 0 265146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_48
timestamp 1725930584
transform 0 -1 360602 -1 0 278646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_49
timestamp 1725930584
transform 0 -1 360602 -1 0 292146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_50
timestamp 1725930584
transform 0 -1 360602 -1 0 305646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_51
timestamp 1725930584
transform 0 -1 360602 -1 0 319146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_52
timestamp 1725930584
transform 1 0 141845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_53
timestamp 1725930584
transform 1 0 155345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_54
timestamp 1725930584
transform 1 0 168845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_55
timestamp 1725930584
transform 1 0 182345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_56
timestamp 1725930584
transform 1 0 195845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_57
timestamp 1725930584
transform 1 0 209345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_58
timestamp 1725930584
transform 1 0 222845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_59
timestamp 1725930584
transform 1 0 236345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_60
timestamp 1725930584
transform 1 0 249845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_61
timestamp 1725930584
transform 1 0 263345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_62
timestamp 1725930584
transform 1 0 276845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_63
timestamp 1725930584
transform 1 0 290345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_64
timestamp 1725930584
transform 1 0 303845 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_65
timestamp 1725930584
transform 1 0 317345 0 1 19400
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_66
timestamp 1725930584
transform 1 0 141845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_67
timestamp 1725930584
transform 1 0 155345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_68
timestamp 1725930584
transform 1 0 168845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_69
timestamp 1725930584
transform 1 0 182345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_70
timestamp 1725930584
transform 1 0 195845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_71
timestamp 1725930584
transform 1 0 209345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_72
timestamp 1725930584
transform 1 0 222845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_73
timestamp 1725930584
transform 1 0 236345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_74
timestamp 1725930584
transform 1 0 249845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_75
timestamp 1725930584
transform 1 0 263345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_76
timestamp 1725930584
transform 1 0 276845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_77
timestamp 1725930584
transform 1 0 290345 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_78
timestamp 1725930584
transform 1 0 303845 0 -1 360600
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_79
timestamp 1725930584
transform 1 0 317345 0 -1 360600
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 44121 0 1 19400
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 330860 0 1 19400
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1569139307
transform 1 0 330845 0 -1 360600
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 44138 0 -1 360600
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 19400 -1 0 49155
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 19400 -1 0 335879
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1569139307
transform 0 -1 360600 -1 0 49155
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1569139307
transform 0 -1 360600 -1 0 335846
box -35 0 5035 25060
use PIC  PAD_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 49000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_1
timestamp 1569139307
transform 1 0 62500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_2
timestamp 1569139307
transform 1 0 76000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_3
timestamp 1569139307
transform 1 0 89500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_4
timestamp 1569139307
transform 1 0 103000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_5
timestamp 1569139307
transform 1 0 116500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_6
timestamp 1569139307
transform 1 0 130000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_7
timestamp 1569139307
transform 1 0 143500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_8
timestamp 1569139307
transform 1 0 157000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_9
timestamp 1569139307
transform 1 0 170500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_10
timestamp 1569139307
transform 1 0 184000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_11
timestamp 1569139307
transform 1 0 197500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_12
timestamp 1569139307
transform 1 0 211000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_13
timestamp 1569139307
transform 1 0 224500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_14
timestamp 1569139307
transform 1 0 238000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_15
timestamp 1569139307
transform 1 0 251500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_16
timestamp 1569139307
transform 1 0 265000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_17
timestamp 1569139307
transform 1 0 278500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_18
timestamp 1569139307
transform 1 0 292000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_19
timestamp 1569139307
transform 1 0 305500 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_20
timestamp 1569139307
transform 1 0 319000 0 1 19400
box -100 -9150 12100 25300
use PIC  PAD_21
timestamp 1569139307
transform 0 -1 360600 1 0 49000
box -100 -9150 12100 25300
use PIC  PAD_22
timestamp 1569139307
transform 0 -1 360600 1 0 62500
box -100 -9150 12100 25300
use PIC  PAD_23
timestamp 1569139307
transform 0 -1 360600 1 0 76000
box -100 -9150 12100 25300
use PIC  PAD_24
timestamp 1569139307
transform 0 -1 360600 1 0 89500
box -100 -9150 12100 25300
use PIC  PAD_25
timestamp 1569139307
transform 0 -1 360600 1 0 103000
box -100 -9150 12100 25300
use PIC  PAD_26
timestamp 1569139307
transform 0 -1 360600 1 0 116500
box -100 -9150 12100 25300
use PIC  PAD_27
timestamp 1569139307
transform 0 -1 360600 1 0 130000
box -100 -9150 12100 25300
use PIC  PAD_28
timestamp 1569139307
transform 0 -1 360600 1 0 143500
box -100 -9150 12100 25300
use PIC  PAD_29
timestamp 1569139307
transform 0 -1 360600 1 0 157000
box -100 -9150 12100 25300
use PIC  PAD_30
timestamp 1569139307
transform 0 -1 360600 1 0 170500
box -100 -9150 12100 25300
use PIC  PAD_31
timestamp 1569139307
transform 0 -1 360600 1 0 184000
box -100 -9150 12100 25300
use PIC  PAD_32
timestamp 1569139307
transform 0 -1 360600 1 0 197500
box -100 -9150 12100 25300
use PIC  PAD_33
timestamp 1569139307
transform 0 -1 360600 1 0 211000
box -100 -9150 12100 25300
use PIC  PAD_34
timestamp 1569139307
transform 0 -1 360600 1 0 224500
box -100 -9150 12100 25300
use PIC  PAD_35
timestamp 1569139307
transform 0 -1 360600 1 0 238000
box -100 -9150 12100 25300
use PIC  PAD_36
timestamp 1569139307
transform 0 -1 360600 1 0 251500
box -100 -9150 12100 25300
use PIC  PAD_37
timestamp 1569139307
transform 0 -1 360600 1 0 265000
box -100 -9150 12100 25300
use PIC  PAD_38
timestamp 1569139307
transform 0 -1 360600 1 0 278500
box -100 -9150 12100 25300
use PIC  PAD_39
timestamp 1569139307
transform 0 -1 360600 1 0 292000
box -100 -9150 12100 25300
use PIC  PAD_40
timestamp 1569139307
transform 0 -1 360600 1 0 305500
box -100 -9150 12100 25300
use PIC  PAD_41
timestamp 1569139307
transform 0 -1 360600 1 0 319000
box -100 -9150 12100 25300
use PIC  PAD_42
timestamp 1569139307
transform 1 0 319000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_43
timestamp 1569139307
transform 1 0 305500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_44
timestamp 1569139307
transform 1 0 292000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_45
timestamp 1569139307
transform 1 0 278500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_46
timestamp 1569139307
transform 1 0 265000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_47
timestamp 1569139307
transform 1 0 251500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_48
timestamp 1569139307
transform 1 0 238000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_49
timestamp 1569139307
transform 1 0 224500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_50
timestamp 1569139307
transform 1 0 211000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_51
timestamp 1569139307
transform 1 0 197500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_52
timestamp 1569139307
transform 1 0 184000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_53
timestamp 1569139307
transform 1 0 170500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_54
timestamp 1569139307
transform 1 0 157000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_55
timestamp 1569139307
transform 1 0 143500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_56
timestamp 1569139307
transform 1 0 130000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_57
timestamp 1569139307
transform 1 0 116500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_58
timestamp 1569139307
transform 1 0 103000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_59
timestamp 1569139307
transform 1 0 89500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_60
timestamp 1569139307
transform 1 0 76000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_61
timestamp 1569139307
transform 1 0 62500 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_62
timestamp 1569139307
transform 1 0 49000 0 -1 360600
box -100 -9150 12100 25300
use PIC  PAD_63
timestamp 1569139307
transform 0 1 19400 -1 0 331000
box -100 -9150 12100 25300
use PIC  PAD_64
timestamp 1569139307
transform 0 1 19400 -1 0 317500
box -100 -9150 12100 25300
use PIC  PAD_65
timestamp 1569139307
transform 0 1 19400 -1 0 304000
box -100 -9150 12100 25300
use PIC  PAD_66
timestamp 1569139307
transform 0 1 19400 -1 0 290500
box -100 -9150 12100 25300
use PIC  PAD_67
timestamp 1569139307
transform 0 1 19400 -1 0 277000
box -100 -9150 12100 25300
use PIC  PAD_68
timestamp 1569139307
transform 0 1 19400 -1 0 263500
box -100 -9150 12100 25300
use PIC  PAD_69
timestamp 1569139307
transform 0 1 19400 -1 0 250000
box -100 -9150 12100 25300
use PIC  PAD_70
timestamp 1569139307
transform 0 1 19400 -1 0 236500
box -100 -9150 12100 25300
use PIC  PAD_71
timestamp 1569139307
transform 0 1 19400 -1 0 223000
box -100 -9150 12100 25300
use PIC  PAD_72
timestamp 1569139307
transform 0 1 19400 -1 0 209500
box -100 -9150 12100 25300
use PIC  PAD_73
timestamp 1569139307
transform 0 1 19400 -1 0 196000
box -100 -9150 12100 25300
use PIC  PAD_74
timestamp 1569139307
transform 0 1 19400 -1 0 182500
box -100 -9150 12100 25300
use PIC  PAD_75
timestamp 1569139307
transform 0 1 19400 -1 0 169000
box -100 -9150 12100 25300
use PIC  PAD_76
timestamp 1569139307
transform 0 1 19400 -1 0 155500
box -100 -9150 12100 25300
use PIC  PAD_77
timestamp 1569139307
transform 0 1 19400 -1 0 142000
box -100 -9150 12100 25300
use PIC  PAD_78
timestamp 1569139307
transform 0 1 19400 -1 0 128500
box -100 -9150 12100 25300
use PIC  PAD_79
timestamp 1569139307
transform 0 1 19400 -1 0 115000
box -100 -9150 12100 25300
use PIC  PAD_80
timestamp 1569139307
transform 0 1 19400 -1 0 101500
box -100 -9150 12100 25300
use PIC  PAD_81
timestamp 1569139307
transform 0 1 19400 -1 0 88000
box -100 -9150 12100 25300
use PIC  PAD_82
timestamp 1569139307
transform 0 1 19400 -1 0 74500
box -100 -9150 12100 25300
use PIC  PAD_83
timestamp 1569139307
transform 0 1 19400 -1 0 61000
box -100 -9150 12100 25300
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 19400 0 1 19400
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 0 -1 360600 1 0 19400
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1569139307
transform -1 0 360600 0 -1 360600
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1569139307
transform 1 0 19400 0 -1 360600
box 0 0 25300 25300
<< end >>
