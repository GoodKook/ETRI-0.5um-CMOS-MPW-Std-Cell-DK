magic
tech scmos
magscale 1 2
timestamp 1727732734
<< nwell >>
rect -13 134 253 252
<< ntransistor >>
rect 25 14 29 54
rect 45 14 49 34
rect 55 14 59 34
rect 77 14 81 34
rect 87 14 91 34
rect 109 14 113 34
rect 153 14 157 34
rect 161 14 165 34
rect 183 14 187 34
rect 193 14 197 34
rect 215 14 219 54
<< ptransistor >>
rect 25 146 29 226
rect 45 186 49 226
rect 61 186 65 226
rect 81 186 85 226
rect 93 186 97 226
rect 113 186 117 226
rect 157 186 161 226
rect 165 186 169 226
rect 185 206 189 226
rect 193 206 197 226
rect 215 146 219 226
<< ndiffusion >>
rect 23 14 25 54
rect 29 34 39 54
rect 202 34 215 54
rect 29 14 31 34
rect 43 14 45 34
rect 49 14 55 34
rect 59 14 63 34
rect 75 14 77 34
rect 81 14 87 34
rect 91 14 93 34
rect 105 14 109 34
rect 113 14 115 34
rect 151 14 153 34
rect 157 14 161 34
rect 165 14 167 34
rect 179 14 183 34
rect 187 14 193 34
rect 197 14 199 34
rect 211 14 215 34
rect 219 14 221 54
<< pdiffusion >>
rect 23 146 25 226
rect 29 186 31 226
rect 43 186 45 226
rect 49 186 61 226
rect 65 186 67 226
rect 79 186 81 226
rect 85 186 93 226
rect 97 186 99 226
rect 111 186 113 226
rect 117 186 119 226
rect 155 186 157 226
rect 161 186 165 226
rect 169 206 171 226
rect 183 206 185 226
rect 189 206 193 226
rect 197 206 201 226
rect 213 206 215 226
rect 169 186 180 206
rect 29 146 38 186
rect 206 146 215 206
rect 219 146 221 226
<< ndcontact >>
rect 11 14 23 54
rect 31 14 43 34
rect 63 14 75 34
rect 93 14 105 34
rect 115 14 127 34
rect 139 14 151 34
rect 167 14 179 34
rect 199 14 211 34
rect 221 14 233 54
<< pdcontact >>
rect 11 146 23 226
rect 31 186 43 226
rect 67 186 79 226
rect 99 186 111 226
rect 119 186 131 226
rect 143 186 155 226
rect 171 206 183 226
rect 201 206 213 226
rect 221 146 233 226
<< psubstratepcontact >>
rect -6 -6 246 6
<< nsubstratencontact >>
rect -6 234 246 246
<< polysilicon >>
rect 25 226 29 230
rect 45 226 49 230
rect 61 226 65 230
rect 81 226 85 230
rect 93 226 97 230
rect 113 226 117 230
rect 157 226 161 230
rect 165 226 169 230
rect 185 226 189 230
rect 193 226 197 230
rect 215 226 219 230
rect 25 103 29 146
rect 45 104 49 186
rect 61 127 65 186
rect 81 146 85 186
rect 93 180 97 186
rect 85 134 88 146
rect 61 119 68 127
rect 25 54 29 91
rect 45 34 49 92
rect 64 90 68 119
rect 84 70 88 134
rect 55 66 88 70
rect 55 34 59 66
rect 93 58 97 168
rect 113 160 117 186
rect 157 182 161 186
rect 125 180 161 182
rect 137 178 161 180
rect 79 46 81 58
rect 77 34 81 46
rect 87 46 89 58
rect 87 34 91 46
rect 109 34 113 148
rect 125 42 129 168
rect 165 154 169 186
rect 185 166 189 206
rect 193 180 197 206
rect 193 176 201 180
rect 163 59 169 154
rect 197 147 201 176
rect 193 141 201 147
rect 193 95 197 141
rect 215 134 219 146
rect 217 122 219 134
rect 163 55 187 59
rect 149 50 165 51
rect 137 46 165 50
rect 125 38 157 42
rect 153 34 157 38
rect 161 34 165 46
rect 183 34 187 55
rect 193 34 197 83
rect 215 54 219 122
rect 25 10 29 14
rect 45 10 49 14
rect 55 10 59 14
rect 77 10 81 14
rect 87 10 91 14
rect 109 10 113 14
rect 153 10 157 14
rect 161 10 165 14
rect 183 10 187 14
rect 193 10 197 14
rect 215 10 219 14
<< polycontact >>
rect 93 168 105 180
rect 73 134 85 146
rect 24 91 36 103
rect 44 92 56 104
rect 64 78 76 90
rect 105 148 117 160
rect 125 168 137 180
rect 67 46 79 58
rect 89 46 101 58
rect 153 154 165 166
rect 177 154 189 166
rect 137 50 149 62
rect 205 122 217 134
rect 191 83 203 95
<< metal1 >>
rect -6 246 246 248
rect -6 232 246 234
rect 31 226 43 232
rect 99 226 111 232
rect 143 226 155 232
rect 201 226 213 232
rect 67 180 75 186
rect 119 180 131 186
rect 57 166 75 180
rect 105 173 125 180
rect 171 172 183 206
rect 67 160 75 166
rect 67 152 105 160
rect 123 156 153 162
rect 11 138 73 146
rect 11 54 17 138
rect 123 142 129 156
rect 171 148 177 166
rect 85 136 129 142
rect 137 142 177 148
rect 56 96 97 102
rect 137 97 143 142
rect 197 134 211 142
rect 225 97 233 146
rect 30 86 36 91
rect 30 78 64 86
rect 83 83 97 96
rect 123 83 143 97
rect 203 83 233 97
rect 69 70 76 78
rect 137 70 143 83
rect 69 64 143 70
rect 69 58 76 64
rect 137 62 143 64
rect 101 46 122 53
rect 225 54 233 83
rect 50 34 57 40
rect 115 34 122 46
rect 172 40 183 48
rect 172 34 179 40
rect 50 28 63 34
rect 31 8 43 14
rect 93 8 105 14
rect 139 8 151 14
rect 199 8 211 14
rect -6 6 246 8
rect -6 -8 246 -6
<< m2contact >>
rect 43 166 57 180
rect 183 172 197 186
rect 183 134 197 148
rect 43 40 57 54
rect 183 40 197 54
<< metal2 >>
rect 48 54 56 166
rect 183 148 191 172
rect 183 54 191 134
<< m1p >>
rect 83 83 97 97
rect 123 83 137 97
rect 203 83 217 97
<< labels >>
rlabel metal1 -6 -8 246 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 203 83 217 97 0 Q
port 2 nsew signal output
rlabel metal1 -6 232 246 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 83 83 97 97 0 D
port 0 nsew signal input
rlabel metal1 123 83 137 97 0 CLK
port 1 nsew clock input
<< properties >>
string FIXED_BBOX 0 0 240 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
