magic
tech scmos
timestamp 1728341909
<< nwell >>
rect -6 67 16 126
<< psubstratepcontact >>
rect -3 -3 13 3
<< nsubstratencontact >>
rect -3 117 13 123
<< metal1 >>
rect -3 123 13 124
rect -3 116 13 117
rect -3 3 13 4
rect -3 -4 13 -3
<< m1p >>
rect -3 116 13 124
<< labels >>
rlabel nsubstratencontact 3 119 3 119 0 vdd
port 0 nsew power bidirectional abutment
rlabel metal1 -3 -4 13 4 0 gnd
port 1 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 10 120
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
