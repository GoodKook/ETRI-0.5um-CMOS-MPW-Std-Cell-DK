magic
tech scmos
magscale 1 2
timestamp 1728304878
<< nwell >>
rect -12 134 92 252
<< ntransistor >>
rect 21 14 25 54
rect 41 14 45 54
<< ptransistor >>
rect 21 146 25 226
rect 41 146 45 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 14 27 54
rect 39 14 41 54
rect 45 14 47 54
<< pdiffusion >>
rect 7 224 21 226
rect 19 146 21 224
rect 25 146 27 226
rect 39 146 41 226
rect 45 146 47 226
<< ndcontact >>
rect 7 14 19 54
rect 27 14 39 54
rect 47 14 59 54
<< pdcontact >>
rect 7 146 19 224
rect 27 146 39 226
rect 47 146 59 226
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 234 86 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 21 142 25 146
rect 41 142 45 146
rect 21 138 45 142
rect 21 89 25 138
rect 16 77 25 89
rect 21 62 25 77
rect 21 58 45 62
rect 21 54 25 58
rect 41 54 45 58
rect 21 10 25 14
rect 41 10 45 14
<< polycontact >>
rect 4 77 16 89
<< metal1 >>
rect -6 246 86 248
rect -6 232 86 234
rect 7 224 19 232
rect 47 226 59 232
rect 29 103 38 146
rect 29 89 43 103
rect 29 54 38 89
rect 7 8 19 14
rect 47 8 59 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 3 89 17 103
rect 43 89 57 103
<< metal2 >>
rect 3 103 17 117
rect 43 103 57 117
<< m1p >>
rect -6 232 86 248
rect -6 -8 86 8
<< m2p >>
rect 3 103 17 117
rect 43 103 57 117
<< labels >>
rlabel metal1 -6 -8 86 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 86 248 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal2 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal2 43 103 57 117 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
