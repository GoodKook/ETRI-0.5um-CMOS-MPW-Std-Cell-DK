magic
tech scmos
magscale 1 2
timestamp 1727495070
<< nwell >>
rect -6 152 86 272
<< ntransistor >>
rect 20 14 24 34
rect 40 14 44 34
<< ptransistor >>
rect 20 166 24 246
rect 34 166 38 246
<< ndiffusion >>
rect 18 14 20 34
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 46 34
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 34 246
rect 38 166 40 246
<< ndcontact >>
rect 6 14 18 34
rect 26 14 38 34
rect 46 14 58 34
<< pdcontact >>
rect 6 166 18 246
rect 40 166 52 246
<< psubstratepcontact >>
rect 0 -6 80 6
<< nsubstratencontact >>
rect 0 254 80 266
<< polysilicon >>
rect 20 246 24 250
rect 34 246 38 250
rect 20 109 24 166
rect 34 161 38 166
rect 34 156 44 161
rect 16 97 24 109
rect 20 34 24 97
rect 40 34 44 156
rect 20 10 24 14
rect 40 10 44 14
<< polycontact >>
rect 4 97 16 109
rect 44 97 56 109
<< metal1 >>
rect 0 266 80 268
rect 0 252 80 254
rect 6 246 18 252
rect 28 166 40 174
rect 28 117 34 166
rect 28 34 34 103
rect 6 8 18 14
rect 46 8 58 14
rect 0 6 80 8
rect 0 -8 80 -6
<< m2contact >>
rect 23 103 37 117
rect 3 83 17 97
rect 43 83 57 97
<< metal2 >>
rect 23 117 37 137
rect 3 63 17 83
rect 43 63 57 83
<< m2p >>
rect 23 123 37 137
rect 3 63 17 77
rect 43 63 57 77
<< labels >>
rlabel metal2 3 63 17 77 0 A
port 0 nsew signal input
rlabel metal2 43 63 57 77 0 B
port 1 nsew signal input
rlabel metal2 23 123 37 137 0 Y
port 2 nsew signal output
rlabel metal1 0 266 80 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 254 80 266 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 252 80 254 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 6 80 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -6 80 6 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -8 80 -6 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
