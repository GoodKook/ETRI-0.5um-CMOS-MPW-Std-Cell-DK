magic
tech scmos
magscale 1 2
timestamp 1756332915
<< nwell >>
rect -3 6144 6742 6356
rect 989 6140 1025 6144
rect -2 5664 6742 5876
rect 1089 5660 1125 5664
rect 3489 5396 3525 5400
rect -3 5278 6742 5396
rect -2 5184 6742 5278
rect 2255 5180 2291 5184
rect 2989 5180 3025 5184
rect 2415 4916 2451 4920
rect -2 4704 6742 4916
rect 2295 4700 2331 4704
rect 509 4436 545 4440
rect 4855 4436 4891 4440
rect 5235 4436 5271 4440
rect -2 4224 6742 4436
rect -2 3838 6743 3956
rect -2 3744 6742 3838
rect -2 3382 6742 3476
rect -2 3264 6743 3382
rect 5362 3256 5437 3264
rect 4723 2996 4798 3004
rect 5962 2996 6037 3004
rect -2 2784 6742 2996
rect 1889 2780 1925 2784
rect 5822 2776 5897 2784
rect 5942 2776 6017 2784
rect 6062 2776 6137 2784
rect 2162 2516 2237 2524
rect 2282 2516 2357 2524
rect 2642 2516 2717 2524
rect 2863 2516 2938 2524
rect 4722 2516 4797 2524
rect -3 2304 6742 2516
rect 3982 2296 4057 2304
rect 4102 2296 4177 2304
rect 4222 2296 4297 2304
rect 4502 2296 4577 2304
rect 4643 2296 4718 2304
rect 4742 2296 4817 2304
rect 4942 2296 5017 2304
rect 5363 2296 5438 2304
rect 5462 2296 5537 2304
rect 5582 2296 5657 2304
rect 6103 2296 6178 2304
rect 6223 2296 6298 2304
rect 1002 2036 1077 2044
rect 1943 2036 2018 2044
rect 2063 2036 2138 2044
rect 2682 2036 2757 2044
rect 2823 2036 2898 2044
rect 5189 2036 5225 2040
rect 6342 2036 6417 2044
rect -2 1824 6742 2036
rect 6182 1816 6257 1824
rect 6302 1816 6377 1824
rect 1423 1556 1498 1564
rect 1543 1556 1618 1564
rect 1663 1556 1738 1564
rect 2002 1556 2077 1564
rect 2823 1556 2898 1564
rect 4303 1556 4378 1564
rect 4423 1556 4498 1564
rect 4522 1556 4597 1564
rect 4642 1556 4717 1564
rect 4762 1556 4837 1564
rect 4882 1556 4957 1564
rect 5602 1556 5677 1564
rect 6303 1556 6378 1564
rect -2 1344 6742 1556
rect 1643 1336 1718 1344
rect 2282 1336 2357 1344
rect 2423 1336 2498 1344
rect 3163 1336 3238 1344
rect 4522 1336 4597 1344
rect 5662 1336 5737 1344
rect 3323 1076 3398 1084
rect 3422 1076 3497 1084
rect 3862 1076 3937 1084
rect 4003 1076 4078 1084
rect 5689 1076 5725 1080
rect -3 958 6742 1076
rect -2 864 6742 958
rect 29 860 65 864
rect 1802 856 1877 864
rect 3123 856 3198 864
rect 3243 856 3318 864
rect 3522 856 3597 864
rect 3723 856 3798 864
rect 4062 856 4137 864
rect 4962 856 5037 864
rect 5103 856 5178 864
rect 5023 596 5098 604
rect 5522 596 5597 604
rect -2 502 6742 596
rect -3 384 6742 502
rect -3 -2 6742 116
<< ntransistor >>
rect 35 6436 39 6476
rect 55 6456 59 6476
rect 65 6456 69 6476
rect 87 6456 91 6476
rect 97 6456 101 6476
rect 119 6456 123 6476
rect 165 6456 169 6476
rect 173 6456 177 6476
rect 193 6456 197 6476
rect 203 6456 207 6476
rect 225 6436 229 6476
rect 285 6436 289 6476
rect 305 6436 309 6476
rect 325 6436 329 6476
rect 373 6436 377 6476
rect 383 6436 387 6476
rect 473 6436 477 6476
rect 483 6436 487 6476
rect 533 6436 537 6476
rect 543 6436 547 6476
rect 611 6436 615 6476
rect 633 6456 637 6476
rect 643 6456 647 6476
rect 663 6456 667 6476
rect 671 6456 675 6476
rect 717 6456 721 6476
rect 739 6456 743 6476
rect 749 6456 753 6476
rect 771 6456 775 6476
rect 781 6456 785 6476
rect 801 6436 805 6476
rect 851 6456 855 6476
rect 914 6436 918 6476
rect 922 6436 926 6476
rect 942 6436 946 6476
rect 950 6436 954 6476
rect 1045 6456 1049 6476
rect 1091 6436 1095 6476
rect 1113 6456 1117 6476
rect 1123 6456 1127 6476
rect 1143 6456 1147 6476
rect 1151 6456 1155 6476
rect 1197 6456 1201 6476
rect 1219 6456 1223 6476
rect 1229 6456 1233 6476
rect 1251 6456 1255 6476
rect 1261 6456 1265 6476
rect 1281 6436 1285 6476
rect 1331 6436 1335 6476
rect 1351 6436 1355 6476
rect 1371 6436 1375 6476
rect 1391 6436 1395 6476
rect 1465 6436 1469 6476
rect 1485 6436 1489 6476
rect 1505 6436 1509 6476
rect 1575 6436 1579 6476
rect 1595 6436 1599 6476
rect 1605 6436 1609 6476
rect 1665 6456 1669 6476
rect 1711 6436 1715 6476
rect 1733 6456 1737 6476
rect 1743 6456 1747 6476
rect 1763 6456 1767 6476
rect 1771 6456 1775 6476
rect 1817 6456 1821 6476
rect 1839 6456 1843 6476
rect 1849 6456 1853 6476
rect 1871 6456 1875 6476
rect 1881 6456 1885 6476
rect 1901 6436 1905 6476
rect 1951 6436 1955 6476
rect 1971 6436 1975 6476
rect 1991 6436 1995 6476
rect 2053 6436 2057 6476
rect 2063 6436 2067 6476
rect 2145 6436 2149 6476
rect 2165 6436 2169 6476
rect 2185 6436 2189 6476
rect 2252 6456 2256 6476
rect 2274 6436 2278 6476
rect 2282 6436 2286 6476
rect 2353 6436 2357 6476
rect 2363 6436 2367 6476
rect 2425 6456 2429 6476
rect 2445 6456 2449 6476
rect 2491 6456 2495 6476
rect 2511 6456 2515 6476
rect 2573 6436 2577 6476
rect 2583 6436 2587 6476
rect 2688 6416 2692 6476
rect 2696 6416 2700 6476
rect 2704 6416 2708 6476
rect 2753 6436 2757 6476
rect 2763 6436 2767 6476
rect 2868 6416 2872 6476
rect 2876 6416 2880 6476
rect 2884 6416 2888 6476
rect 2945 6436 2949 6476
rect 2965 6436 2969 6476
rect 2985 6436 2989 6476
rect 3045 6436 3049 6476
rect 3065 6436 3069 6476
rect 3085 6436 3089 6476
rect 3145 6456 3149 6476
rect 3205 6456 3209 6476
rect 3254 6436 3258 6476
rect 3262 6436 3266 6476
rect 3284 6456 3288 6476
rect 3351 6436 3355 6476
rect 3371 6436 3375 6476
rect 3391 6436 3395 6476
rect 3472 6456 3476 6476
rect 3494 6436 3498 6476
rect 3502 6436 3506 6476
rect 3572 6456 3576 6476
rect 3594 6436 3598 6476
rect 3602 6436 3606 6476
rect 3652 6416 3656 6476
rect 3660 6416 3664 6476
rect 3668 6416 3672 6476
rect 3765 6436 3769 6476
rect 3785 6436 3789 6476
rect 3805 6436 3809 6476
rect 3851 6436 3855 6476
rect 3871 6436 3875 6476
rect 3891 6436 3895 6476
rect 3951 6456 3955 6476
rect 4013 6436 4017 6476
rect 4023 6436 4027 6476
rect 4115 6436 4119 6476
rect 4135 6436 4139 6476
rect 4145 6436 4149 6476
rect 4193 6436 4197 6476
rect 4203 6436 4207 6476
rect 4308 6416 4312 6476
rect 4316 6416 4320 6476
rect 4324 6416 4328 6476
rect 4408 6416 4412 6476
rect 4416 6416 4420 6476
rect 4424 6416 4428 6476
rect 4508 6416 4512 6476
rect 4516 6416 4520 6476
rect 4524 6416 4528 6476
rect 4571 6456 4575 6476
rect 4634 6436 4638 6476
rect 4642 6436 4646 6476
rect 4664 6456 4668 6476
rect 4734 6436 4738 6476
rect 4742 6436 4746 6476
rect 4764 6456 4768 6476
rect 4831 6436 4835 6476
rect 4851 6436 4855 6476
rect 4871 6436 4875 6476
rect 4945 6436 4949 6476
rect 4965 6436 4969 6476
rect 4985 6436 4989 6476
rect 5031 6436 5035 6476
rect 5051 6436 5055 6476
rect 5071 6436 5075 6476
rect 5168 6416 5172 6476
rect 5176 6416 5180 6476
rect 5184 6416 5188 6476
rect 5268 6416 5272 6476
rect 5276 6416 5280 6476
rect 5284 6416 5288 6476
rect 5368 6416 5372 6476
rect 5376 6416 5380 6476
rect 5384 6416 5388 6476
rect 5434 6436 5438 6476
rect 5442 6436 5446 6476
rect 5464 6456 5468 6476
rect 5552 6456 5556 6476
rect 5574 6436 5578 6476
rect 5582 6436 5586 6476
rect 5645 6456 5649 6476
rect 5694 6436 5698 6476
rect 5702 6436 5706 6476
rect 5724 6456 5728 6476
rect 5792 6416 5796 6476
rect 5800 6416 5804 6476
rect 5808 6416 5812 6476
rect 5912 6456 5916 6476
rect 5934 6436 5938 6476
rect 5942 6436 5946 6476
rect 6005 6456 6009 6476
rect 6072 6456 6076 6476
rect 6094 6436 6098 6476
rect 6102 6436 6106 6476
rect 6165 6436 6169 6476
rect 6185 6436 6189 6476
rect 6205 6436 6209 6476
rect 6272 6456 6276 6476
rect 6294 6436 6298 6476
rect 6302 6436 6306 6476
rect 6352 6416 6356 6476
rect 6360 6416 6364 6476
rect 6368 6416 6372 6476
rect 6488 6416 6492 6476
rect 6496 6416 6500 6476
rect 6504 6416 6508 6476
rect 6551 6456 6555 6476
rect 6614 6436 6618 6476
rect 6622 6436 6626 6476
rect 6642 6436 6646 6476
rect 6650 6436 6654 6476
rect 31 6024 35 6064
rect 53 6024 57 6044
rect 63 6024 67 6044
rect 83 6024 87 6044
rect 91 6024 95 6044
rect 137 6024 141 6044
rect 159 6024 163 6044
rect 169 6024 173 6044
rect 191 6024 195 6044
rect 201 6024 205 6044
rect 221 6024 225 6064
rect 292 6024 296 6044
rect 314 6024 318 6064
rect 322 6024 326 6064
rect 393 6024 397 6064
rect 403 6024 407 6064
rect 451 6024 455 6044
rect 471 6024 475 6044
rect 553 6024 557 6064
rect 563 6024 567 6064
rect 611 6024 615 6064
rect 631 6024 635 6064
rect 651 6024 655 6064
rect 725 6024 729 6064
rect 745 6024 749 6064
rect 765 6024 769 6064
rect 811 6024 815 6044
rect 831 6024 835 6044
rect 912 6024 916 6044
rect 934 6024 938 6064
rect 942 6024 946 6064
rect 991 6024 995 6044
rect 1011 6024 1015 6044
rect 1031 6024 1035 6064
rect 1105 6024 1109 6044
rect 1151 6024 1155 6044
rect 1171 6024 1175 6044
rect 1245 6024 1249 6064
rect 1265 6024 1269 6064
rect 1285 6024 1289 6064
rect 1345 6024 1349 6044
rect 1405 6024 1409 6044
rect 1451 6024 1455 6044
rect 1471 6024 1475 6044
rect 1531 6024 1535 6044
rect 1551 6024 1555 6044
rect 1611 6024 1615 6044
rect 1671 6024 1675 6044
rect 1691 6024 1695 6044
rect 1751 6024 1755 6044
rect 1771 6024 1775 6044
rect 1831 6024 1835 6064
rect 1851 6024 1855 6064
rect 1871 6024 1875 6064
rect 1931 6024 1935 6044
rect 2012 6024 2016 6044
rect 2034 6024 2038 6064
rect 2042 6024 2046 6064
rect 2091 6024 2095 6044
rect 2165 6024 2169 6064
rect 2185 6024 2189 6064
rect 2205 6024 2209 6064
rect 2251 6024 2255 6044
rect 2325 6024 2329 6064
rect 2345 6024 2349 6064
rect 2365 6024 2369 6064
rect 2448 6024 2452 6084
rect 2456 6024 2460 6084
rect 2464 6024 2468 6084
rect 2532 6024 2536 6044
rect 2554 6024 2558 6064
rect 2562 6024 2566 6064
rect 2625 6024 2629 6044
rect 2645 6024 2649 6044
rect 2728 6024 2732 6084
rect 2736 6024 2740 6084
rect 2744 6024 2748 6084
rect 2826 6024 2830 6064
rect 2834 6024 2838 6064
rect 2854 6024 2858 6064
rect 2862 6024 2866 6064
rect 2925 6024 2929 6044
rect 2972 6024 2976 6084
rect 2980 6024 2984 6084
rect 2988 6024 2992 6084
rect 3092 6024 3096 6044
rect 3114 6024 3118 6064
rect 3122 6024 3126 6064
rect 3208 6024 3212 6084
rect 3216 6024 3220 6084
rect 3224 6024 3228 6084
rect 3292 6024 3296 6044
rect 3314 6024 3318 6064
rect 3322 6024 3326 6064
rect 3385 6024 3389 6044
rect 3468 6024 3472 6084
rect 3476 6024 3480 6084
rect 3484 6024 3488 6084
rect 3532 6024 3536 6084
rect 3540 6024 3544 6084
rect 3548 6024 3552 6084
rect 3631 6024 3635 6044
rect 3694 6024 3698 6064
rect 3702 6024 3706 6064
rect 3724 6024 3728 6044
rect 3813 6024 3817 6064
rect 3823 6024 3827 6064
rect 3873 6024 3877 6064
rect 3883 6024 3887 6064
rect 3965 6024 3969 6064
rect 3985 6024 3989 6064
rect 4005 6024 4009 6064
rect 4051 6024 4055 6064
rect 4071 6024 4075 6064
rect 4091 6024 4095 6064
rect 4165 6024 4169 6044
rect 4185 6024 4189 6044
rect 4231 6024 4235 6044
rect 4313 6024 4317 6064
rect 4323 6024 4327 6064
rect 4371 6024 4375 6064
rect 4381 6024 4385 6064
rect 4401 6024 4405 6064
rect 4485 6024 4489 6064
rect 4505 6024 4509 6064
rect 4525 6024 4529 6064
rect 4592 6024 4596 6044
rect 4614 6024 4618 6064
rect 4622 6024 4626 6064
rect 4672 6024 4676 6084
rect 4680 6024 4684 6084
rect 4688 6024 4692 6084
rect 4792 6024 4796 6044
rect 4814 6024 4818 6064
rect 4822 6024 4826 6064
rect 4908 6024 4912 6084
rect 4916 6024 4920 6084
rect 4924 6024 4928 6084
rect 4972 6024 4976 6084
rect 4980 6024 4984 6084
rect 4988 6024 4992 6084
rect 5085 6024 5089 6064
rect 5105 6024 5109 6064
rect 5125 6024 5129 6064
rect 5193 6024 5197 6064
rect 5203 6024 5207 6064
rect 5251 6024 5255 6064
rect 5261 6024 5265 6064
rect 5281 6024 5285 6064
rect 5351 6024 5355 6064
rect 5371 6024 5375 6064
rect 5391 6024 5395 6064
rect 5472 6024 5476 6044
rect 5494 6024 5498 6064
rect 5502 6024 5506 6064
rect 5588 6024 5592 6084
rect 5596 6024 5600 6084
rect 5604 6024 5608 6084
rect 5652 6024 5656 6084
rect 5660 6024 5664 6084
rect 5668 6024 5672 6084
rect 5772 6024 5776 6044
rect 5794 6024 5798 6064
rect 5802 6024 5806 6064
rect 5852 6024 5856 6084
rect 5860 6024 5864 6084
rect 5868 6024 5872 6084
rect 5951 6024 5955 6064
rect 5971 6024 5975 6064
rect 5991 6024 5995 6064
rect 6051 6024 6055 6064
rect 6071 6024 6075 6064
rect 6091 6024 6095 6064
rect 6152 6024 6156 6084
rect 6160 6024 6164 6084
rect 6168 6024 6172 6084
rect 6252 6024 6256 6084
rect 6260 6024 6264 6084
rect 6268 6024 6272 6084
rect 6388 6024 6392 6084
rect 6396 6024 6400 6084
rect 6404 6024 6408 6084
rect 6472 6024 6476 6044
rect 6494 6024 6498 6064
rect 6502 6024 6506 6064
rect 6551 6024 6555 6044
rect 6611 6024 6615 6044
rect 43 5956 47 5996
rect 65 5976 69 5996
rect 113 5956 117 5996
rect 123 5956 127 5996
rect 193 5956 197 5996
rect 203 5956 207 5996
rect 292 5976 296 5996
rect 314 5956 318 5996
rect 322 5956 326 5996
rect 393 5956 397 5996
rect 403 5956 407 5996
rect 451 5976 455 5996
rect 525 5976 529 5996
rect 545 5976 549 5996
rect 591 5976 595 5996
rect 611 5976 615 5996
rect 671 5956 675 5996
rect 691 5956 695 5996
rect 711 5956 715 5996
rect 785 5976 789 5996
rect 831 5976 835 5996
rect 851 5976 855 5996
rect 933 5956 937 5996
rect 943 5956 947 5996
rect 1005 5956 1009 5996
rect 1025 5956 1029 5996
rect 1045 5956 1049 5996
rect 1091 5976 1095 5996
rect 1111 5976 1115 5996
rect 1185 5976 1189 5996
rect 1231 5956 1235 5996
rect 1253 5976 1257 5996
rect 1263 5976 1267 5996
rect 1283 5976 1287 5996
rect 1291 5976 1295 5996
rect 1337 5976 1341 5996
rect 1359 5976 1363 5996
rect 1369 5976 1373 5996
rect 1391 5976 1395 5996
rect 1401 5976 1405 5996
rect 1421 5956 1425 5996
rect 1473 5956 1477 5996
rect 1483 5956 1487 5996
rect 1588 5936 1592 5996
rect 1596 5936 1600 5996
rect 1604 5936 1608 5996
rect 1665 5956 1669 5996
rect 1685 5956 1689 5996
rect 1705 5956 1709 5996
rect 1765 5976 1769 5996
rect 1785 5976 1789 5996
rect 1868 5936 1872 5996
rect 1876 5936 1880 5996
rect 1884 5936 1888 5996
rect 1931 5976 1935 5996
rect 2005 5956 2009 5996
rect 2025 5956 2029 5996
rect 2045 5956 2049 5996
rect 2092 5936 2096 5996
rect 2100 5936 2104 5996
rect 2108 5936 2112 5996
rect 2212 5976 2216 5996
rect 2234 5956 2238 5996
rect 2242 5956 2246 5996
rect 2291 5956 2295 5996
rect 2311 5956 2315 5996
rect 2331 5956 2335 5996
rect 2413 5956 2417 5996
rect 2423 5956 2427 5996
rect 2508 5936 2512 5996
rect 2516 5936 2520 5996
rect 2524 5936 2528 5996
rect 2592 5976 2596 5996
rect 2614 5956 2618 5996
rect 2622 5956 2626 5996
rect 2673 5956 2677 5996
rect 2683 5956 2687 5996
rect 2788 5936 2792 5996
rect 2796 5936 2800 5996
rect 2804 5936 2808 5996
rect 2888 5936 2892 5996
rect 2896 5936 2900 5996
rect 2904 5936 2908 5996
rect 2988 5936 2992 5996
rect 2996 5936 3000 5996
rect 3004 5936 3008 5996
rect 3088 5936 3092 5996
rect 3096 5936 3100 5996
rect 3104 5936 3108 5996
rect 3152 5936 3156 5996
rect 3160 5936 3164 5996
rect 3168 5936 3172 5996
rect 3265 5956 3269 5996
rect 3285 5956 3289 5996
rect 3305 5956 3309 5996
rect 3351 5956 3355 5996
rect 3371 5956 3375 5996
rect 3391 5956 3395 5996
rect 3472 5976 3476 5996
rect 3494 5956 3498 5996
rect 3502 5956 3506 5996
rect 3565 5956 3569 5996
rect 3585 5956 3589 5996
rect 3605 5956 3609 5996
rect 3688 5936 3692 5996
rect 3696 5936 3700 5996
rect 3704 5936 3708 5996
rect 3754 5956 3758 5996
rect 3762 5956 3766 5996
rect 3784 5976 3788 5996
rect 3888 5936 3892 5996
rect 3896 5936 3900 5996
rect 3904 5936 3908 5996
rect 3972 5976 3976 5996
rect 3994 5956 3998 5996
rect 4002 5956 4006 5996
rect 4088 5936 4092 5996
rect 4096 5936 4100 5996
rect 4104 5936 4108 5996
rect 4172 5976 4176 5996
rect 4194 5956 4198 5996
rect 4202 5956 4206 5996
rect 4252 5936 4256 5996
rect 4260 5936 4264 5996
rect 4268 5936 4272 5996
rect 4353 5956 4357 5996
rect 4363 5956 4367 5996
rect 4445 5956 4449 5996
rect 4465 5956 4469 5996
rect 4485 5956 4489 5996
rect 4545 5976 4549 5996
rect 4565 5976 4569 5996
rect 4611 5956 4615 5996
rect 4621 5956 4625 5996
rect 4641 5956 4645 5996
rect 4732 5976 4736 5996
rect 4754 5956 4758 5996
rect 4762 5956 4766 5996
rect 4813 5956 4817 5996
rect 4823 5956 4827 5996
rect 4905 5976 4909 5996
rect 4988 5936 4992 5996
rect 4996 5936 5000 5996
rect 5004 5936 5008 5996
rect 5054 5956 5058 5996
rect 5062 5956 5066 5996
rect 5084 5976 5088 5996
rect 5151 5956 5155 5996
rect 5171 5956 5175 5996
rect 5191 5956 5195 5996
rect 5251 5956 5255 5996
rect 5271 5956 5275 5996
rect 5291 5956 5295 5996
rect 5354 5956 5358 5996
rect 5362 5956 5366 5996
rect 5382 5956 5386 5996
rect 5390 5956 5394 5996
rect 5493 5956 5497 5996
rect 5503 5956 5507 5996
rect 5551 5976 5555 5996
rect 5648 5936 5652 5996
rect 5656 5936 5660 5996
rect 5664 5936 5668 5996
rect 5714 5956 5718 5996
rect 5722 5956 5726 5996
rect 5744 5976 5748 5996
rect 5825 5956 5829 5996
rect 5845 5956 5849 5996
rect 5865 5956 5869 5996
rect 5911 5956 5915 5996
rect 5931 5956 5935 5996
rect 5951 5956 5955 5996
rect 6025 5956 6029 5996
rect 6045 5956 6049 5996
rect 6065 5956 6069 5996
rect 6114 5956 6118 5996
rect 6122 5956 6126 5996
rect 6142 5956 6146 5996
rect 6150 5956 6154 5996
rect 6253 5956 6257 5996
rect 6263 5956 6267 5996
rect 6311 5956 6315 5996
rect 6321 5956 6325 5996
rect 6341 5956 6345 5996
rect 6411 5956 6415 5996
rect 6431 5956 6435 5996
rect 6451 5956 6455 5996
rect 6512 5936 6516 5996
rect 6520 5936 6524 5996
rect 6528 5936 6532 5996
rect 6613 5956 6617 5996
rect 6623 5956 6627 5996
rect 43 5544 47 5584
rect 65 5544 69 5564
rect 123 5544 127 5584
rect 145 5544 149 5564
rect 191 5544 195 5584
rect 213 5544 217 5564
rect 223 5544 227 5564
rect 243 5544 247 5564
rect 251 5544 255 5564
rect 297 5544 301 5564
rect 319 5544 323 5564
rect 329 5544 333 5564
rect 351 5544 355 5564
rect 361 5544 365 5564
rect 381 5544 385 5584
rect 445 5544 449 5564
rect 465 5544 469 5564
rect 514 5544 518 5584
rect 522 5544 526 5584
rect 544 5544 548 5564
rect 613 5544 617 5584
rect 623 5544 627 5584
rect 691 5544 695 5584
rect 701 5544 705 5584
rect 721 5544 725 5584
rect 793 5544 797 5584
rect 803 5544 807 5584
rect 873 5544 877 5584
rect 883 5544 887 5584
rect 951 5544 955 5564
rect 971 5544 975 5564
rect 1031 5544 1035 5564
rect 1091 5544 1095 5564
rect 1111 5544 1115 5564
rect 1131 5544 1135 5584
rect 1191 5544 1195 5564
rect 1211 5544 1215 5564
rect 1271 5544 1275 5564
rect 1331 5544 1335 5564
rect 1351 5544 1355 5564
rect 1411 5544 1415 5564
rect 1471 5544 1475 5584
rect 1493 5544 1497 5564
rect 1503 5544 1507 5564
rect 1523 5544 1527 5564
rect 1531 5544 1535 5564
rect 1577 5544 1581 5564
rect 1599 5544 1603 5564
rect 1609 5544 1613 5564
rect 1631 5544 1635 5564
rect 1641 5544 1645 5564
rect 1661 5544 1665 5584
rect 1711 5544 1715 5584
rect 1731 5544 1735 5584
rect 1751 5544 1755 5584
rect 1771 5544 1775 5584
rect 1845 5544 1849 5584
rect 1865 5544 1869 5584
rect 1885 5544 1889 5584
rect 1953 5544 1957 5584
rect 1963 5544 1967 5584
rect 2011 5544 2015 5564
rect 2092 5544 2096 5564
rect 2114 5544 2118 5584
rect 2122 5544 2126 5584
rect 2171 5544 2175 5564
rect 2191 5544 2195 5564
rect 2253 5544 2257 5584
rect 2263 5544 2267 5584
rect 2405 5544 2409 5564
rect 2425 5544 2429 5564
rect 2445 5544 2449 5564
rect 2533 5544 2537 5584
rect 2543 5544 2547 5584
rect 2628 5544 2632 5604
rect 2636 5544 2640 5604
rect 2644 5544 2648 5604
rect 2728 5544 2732 5604
rect 2736 5544 2740 5604
rect 2744 5544 2748 5604
rect 2793 5544 2797 5584
rect 2803 5544 2807 5584
rect 2871 5544 2875 5584
rect 2891 5544 2895 5584
rect 2911 5544 2915 5584
rect 3008 5544 3012 5604
rect 3016 5544 3020 5604
rect 3024 5544 3028 5604
rect 3074 5544 3078 5584
rect 3082 5544 3086 5584
rect 3104 5544 3108 5564
rect 3185 5544 3189 5584
rect 3205 5544 3209 5584
rect 3225 5544 3229 5584
rect 3285 5544 3289 5564
rect 3332 5544 3336 5604
rect 3340 5544 3344 5604
rect 3348 5544 3352 5604
rect 3468 5544 3472 5604
rect 3476 5544 3480 5604
rect 3484 5544 3488 5604
rect 3568 5544 3572 5604
rect 3576 5544 3580 5604
rect 3584 5544 3588 5604
rect 3645 5544 3649 5564
rect 3705 5544 3709 5584
rect 3725 5544 3729 5584
rect 3745 5544 3749 5584
rect 3805 5544 3809 5564
rect 3825 5544 3829 5564
rect 3871 5544 3875 5584
rect 3891 5544 3895 5584
rect 3911 5544 3915 5584
rect 3985 5544 3989 5564
rect 4066 5544 4070 5584
rect 4074 5544 4078 5584
rect 4094 5544 4098 5584
rect 4102 5544 4106 5584
rect 4165 5544 4169 5584
rect 4185 5544 4189 5584
rect 4205 5544 4209 5584
rect 4288 5544 4292 5604
rect 4296 5544 4300 5604
rect 4304 5544 4308 5604
rect 4351 5544 4355 5564
rect 4425 5544 4429 5584
rect 4445 5544 4449 5584
rect 4465 5544 4469 5584
rect 4535 5544 4539 5584
rect 4555 5544 4559 5584
rect 4565 5544 4569 5584
rect 4613 5544 4617 5584
rect 4623 5544 4627 5584
rect 4705 5544 4709 5584
rect 4725 5544 4729 5584
rect 4745 5544 4749 5584
rect 4791 5544 4795 5584
rect 4811 5544 4815 5584
rect 4831 5544 4835 5584
rect 4928 5544 4932 5604
rect 4936 5544 4940 5604
rect 4944 5544 4948 5604
rect 4994 5544 4998 5584
rect 5002 5544 5006 5584
rect 5024 5544 5028 5564
rect 5091 5544 5095 5584
rect 5111 5544 5115 5584
rect 5131 5544 5135 5584
rect 5192 5544 5196 5604
rect 5200 5544 5204 5604
rect 5208 5544 5212 5604
rect 5293 5544 5297 5584
rect 5303 5544 5307 5584
rect 5372 5544 5376 5604
rect 5380 5544 5384 5604
rect 5388 5544 5392 5604
rect 5474 5544 5478 5584
rect 5482 5544 5486 5584
rect 5504 5544 5508 5564
rect 5573 5544 5577 5584
rect 5583 5544 5587 5584
rect 5673 5544 5677 5584
rect 5683 5544 5687 5584
rect 5734 5544 5738 5584
rect 5742 5544 5746 5584
rect 5762 5544 5766 5584
rect 5770 5544 5774 5584
rect 5865 5544 5869 5584
rect 5885 5544 5889 5584
rect 5905 5544 5909 5584
rect 5951 5544 5955 5564
rect 6014 5544 6018 5584
rect 6022 5544 6026 5584
rect 6042 5544 6046 5584
rect 6050 5544 6054 5584
rect 6132 5544 6136 5604
rect 6140 5544 6144 5604
rect 6148 5544 6152 5604
rect 6245 5544 6249 5564
rect 6294 5544 6298 5584
rect 6302 5544 6306 5584
rect 6324 5544 6328 5564
rect 6392 5544 6396 5604
rect 6400 5544 6404 5604
rect 6408 5544 6412 5604
rect 6492 5544 6496 5604
rect 6500 5544 6504 5604
rect 6508 5544 6512 5604
rect 6592 5544 6596 5604
rect 6600 5544 6604 5604
rect 6608 5544 6612 5604
rect 31 5476 35 5516
rect 53 5496 57 5516
rect 63 5496 67 5516
rect 83 5496 87 5516
rect 91 5496 95 5516
rect 137 5496 141 5516
rect 159 5496 163 5516
rect 169 5496 173 5516
rect 191 5496 195 5516
rect 201 5496 205 5516
rect 221 5476 225 5516
rect 273 5476 277 5516
rect 283 5476 287 5516
rect 372 5496 376 5516
rect 394 5476 398 5516
rect 402 5476 406 5516
rect 473 5476 477 5516
rect 483 5476 487 5516
rect 555 5476 559 5516
rect 575 5476 579 5516
rect 585 5476 589 5516
rect 631 5496 635 5516
rect 651 5496 655 5516
rect 711 5496 715 5516
rect 731 5496 735 5516
rect 793 5476 797 5516
rect 803 5476 807 5516
rect 873 5476 877 5516
rect 883 5476 887 5516
rect 951 5496 955 5516
rect 1014 5476 1018 5516
rect 1022 5476 1026 5516
rect 1044 5496 1048 5516
rect 1146 5476 1150 5516
rect 1154 5476 1158 5516
rect 1174 5476 1178 5516
rect 1182 5476 1186 5516
rect 1231 5476 1235 5516
rect 1253 5496 1257 5516
rect 1263 5496 1267 5516
rect 1283 5496 1287 5516
rect 1291 5496 1295 5516
rect 1337 5496 1341 5516
rect 1359 5496 1363 5516
rect 1369 5496 1373 5516
rect 1391 5496 1395 5516
rect 1401 5496 1405 5516
rect 1421 5476 1425 5516
rect 1508 5456 1512 5516
rect 1516 5456 1520 5516
rect 1524 5456 1528 5516
rect 1608 5456 1612 5516
rect 1616 5456 1620 5516
rect 1624 5456 1628 5516
rect 1685 5496 1689 5516
rect 1745 5476 1749 5516
rect 1765 5476 1769 5516
rect 1785 5476 1789 5516
rect 1855 5476 1859 5516
rect 1875 5476 1879 5516
rect 1885 5476 1889 5516
rect 1953 5476 1957 5516
rect 1963 5476 1967 5516
rect 2025 5476 2029 5516
rect 2045 5476 2049 5516
rect 2065 5476 2069 5516
rect 2113 5476 2117 5516
rect 2123 5476 2127 5516
rect 2205 5496 2209 5516
rect 2265 5476 2269 5516
rect 2285 5476 2289 5516
rect 2305 5476 2309 5516
rect 2351 5496 2355 5516
rect 2371 5496 2375 5516
rect 2445 5496 2449 5516
rect 2512 5496 2516 5516
rect 2534 5476 2538 5516
rect 2542 5476 2546 5516
rect 2591 5476 2595 5516
rect 2611 5476 2615 5516
rect 2631 5476 2635 5516
rect 2693 5476 2697 5516
rect 2703 5476 2707 5516
rect 2808 5456 2812 5516
rect 2816 5456 2820 5516
rect 2824 5456 2828 5516
rect 2893 5476 2897 5516
rect 2903 5476 2907 5516
rect 2965 5496 2969 5516
rect 2985 5496 2989 5516
rect 3031 5476 3035 5516
rect 3051 5476 3055 5516
rect 3071 5476 3075 5516
rect 3153 5476 3157 5516
rect 3163 5476 3167 5516
rect 3211 5476 3215 5516
rect 3231 5476 3235 5516
rect 3251 5476 3255 5516
rect 3335 5476 3339 5516
rect 3355 5476 3359 5516
rect 3365 5476 3369 5516
rect 3411 5496 3415 5516
rect 3431 5496 3435 5516
rect 3491 5496 3495 5516
rect 3511 5496 3515 5516
rect 3531 5476 3535 5516
rect 3591 5476 3595 5516
rect 3611 5476 3615 5516
rect 3631 5476 3635 5516
rect 3705 5496 3709 5516
rect 3725 5496 3729 5516
rect 3771 5476 3775 5516
rect 3791 5476 3795 5516
rect 3811 5476 3815 5516
rect 3831 5476 3835 5516
rect 3905 5496 3909 5516
rect 3925 5496 3929 5516
rect 3971 5476 3975 5516
rect 3991 5476 3995 5516
rect 4011 5476 4015 5516
rect 4108 5456 4112 5516
rect 4116 5456 4120 5516
rect 4124 5456 4128 5516
rect 4193 5476 4197 5516
rect 4203 5476 4207 5516
rect 4251 5496 4255 5516
rect 4325 5476 4329 5516
rect 4345 5476 4349 5516
rect 4365 5476 4369 5516
rect 4433 5476 4437 5516
rect 4443 5476 4447 5516
rect 4493 5476 4497 5516
rect 4503 5476 4507 5516
rect 4585 5476 4589 5516
rect 4605 5476 4609 5516
rect 4625 5476 4629 5516
rect 4685 5476 4689 5516
rect 4705 5476 4709 5516
rect 4725 5476 4729 5516
rect 4795 5476 4799 5516
rect 4815 5476 4819 5516
rect 4825 5476 4829 5516
rect 4885 5476 4889 5516
rect 4905 5476 4909 5516
rect 4925 5476 4929 5516
rect 4993 5476 4997 5516
rect 5003 5476 5007 5516
rect 5075 5476 5079 5516
rect 5095 5476 5099 5516
rect 5105 5476 5109 5516
rect 5153 5476 5157 5516
rect 5163 5476 5167 5516
rect 5231 5476 5235 5516
rect 5251 5476 5255 5516
rect 5271 5476 5275 5516
rect 5355 5476 5359 5516
rect 5375 5476 5379 5516
rect 5385 5476 5389 5516
rect 5431 5476 5435 5516
rect 5451 5476 5455 5516
rect 5471 5476 5475 5516
rect 5533 5476 5537 5516
rect 5543 5476 5547 5516
rect 5612 5456 5616 5516
rect 5620 5456 5624 5516
rect 5628 5456 5632 5516
rect 5735 5476 5739 5516
rect 5755 5476 5759 5516
rect 5765 5476 5769 5516
rect 5846 5476 5850 5516
rect 5854 5476 5858 5516
rect 5874 5476 5878 5516
rect 5882 5476 5886 5516
rect 5933 5476 5937 5516
rect 5943 5476 5947 5516
rect 6012 5456 6016 5516
rect 6020 5456 6024 5516
rect 6028 5456 6032 5516
rect 6114 5476 6118 5516
rect 6122 5476 6126 5516
rect 6144 5496 6148 5516
rect 6225 5476 6229 5516
rect 6245 5476 6249 5516
rect 6265 5476 6269 5516
rect 6311 5476 6315 5516
rect 6331 5476 6335 5516
rect 6351 5476 6355 5516
rect 6425 5476 6429 5516
rect 6445 5476 6449 5516
rect 6465 5476 6469 5516
rect 6548 5456 6552 5516
rect 6556 5456 6560 5516
rect 6564 5456 6568 5516
rect 6632 5496 6636 5516
rect 6654 5476 6658 5516
rect 6662 5476 6666 5516
rect 43 5064 47 5104
rect 65 5064 69 5084
rect 111 5064 115 5104
rect 133 5064 137 5084
rect 143 5064 147 5084
rect 163 5064 167 5084
rect 171 5064 175 5084
rect 217 5064 221 5084
rect 239 5064 243 5084
rect 249 5064 253 5084
rect 271 5064 275 5084
rect 281 5064 285 5084
rect 301 5064 305 5104
rect 353 5064 357 5104
rect 363 5064 367 5104
rect 452 5064 456 5084
rect 474 5064 478 5104
rect 482 5064 486 5104
rect 553 5064 557 5104
rect 563 5064 567 5104
rect 615 5064 619 5104
rect 635 5064 639 5084
rect 645 5064 649 5084
rect 667 5064 671 5084
rect 677 5064 681 5084
rect 699 5064 703 5084
rect 745 5064 749 5084
rect 753 5064 757 5084
rect 773 5064 777 5084
rect 783 5064 787 5084
rect 805 5064 809 5104
rect 853 5064 857 5104
rect 863 5064 867 5104
rect 945 5064 949 5104
rect 965 5064 969 5104
rect 985 5064 989 5104
rect 1045 5064 1049 5104
rect 1065 5064 1069 5104
rect 1085 5064 1089 5104
rect 1155 5064 1159 5104
rect 1175 5064 1179 5104
rect 1185 5064 1189 5104
rect 1231 5064 1235 5104
rect 1253 5064 1257 5084
rect 1263 5064 1267 5084
rect 1283 5064 1287 5084
rect 1291 5064 1295 5084
rect 1337 5064 1341 5084
rect 1359 5064 1363 5084
rect 1369 5064 1373 5084
rect 1391 5064 1395 5084
rect 1401 5064 1405 5084
rect 1421 5064 1425 5104
rect 1493 5064 1497 5104
rect 1503 5064 1507 5104
rect 1553 5064 1557 5104
rect 1563 5064 1567 5104
rect 1631 5064 1635 5104
rect 1653 5064 1657 5084
rect 1663 5064 1667 5084
rect 1683 5064 1687 5084
rect 1691 5064 1695 5084
rect 1737 5064 1741 5084
rect 1759 5064 1763 5084
rect 1769 5064 1773 5084
rect 1791 5064 1795 5084
rect 1801 5064 1805 5084
rect 1821 5064 1825 5104
rect 1906 5064 1910 5104
rect 1914 5064 1918 5104
rect 1934 5064 1938 5104
rect 1942 5064 1946 5104
rect 1991 5064 1995 5084
rect 2075 5064 2079 5104
rect 2095 5064 2099 5104
rect 2105 5064 2109 5104
rect 2153 5064 2157 5104
rect 2163 5064 2167 5104
rect 2245 5064 2249 5104
rect 2265 5064 2269 5084
rect 2285 5064 2289 5084
rect 2353 5064 2357 5104
rect 2363 5064 2367 5104
rect 2448 5064 2452 5124
rect 2456 5064 2460 5124
rect 2464 5064 2468 5124
rect 2525 5064 2529 5084
rect 2545 5064 2549 5084
rect 2591 5064 2595 5084
rect 2675 5064 2679 5104
rect 2695 5064 2699 5104
rect 2705 5064 2709 5104
rect 2751 5064 2755 5084
rect 2771 5064 2775 5084
rect 2853 5064 2857 5104
rect 2863 5064 2867 5104
rect 2933 5064 2937 5104
rect 2943 5064 2947 5104
rect 2991 5064 2995 5084
rect 3011 5064 3015 5084
rect 3031 5064 3035 5104
rect 3115 5064 3119 5104
rect 3135 5064 3139 5104
rect 3145 5064 3149 5104
rect 3193 5064 3197 5104
rect 3203 5064 3207 5104
rect 3308 5064 3312 5124
rect 3316 5064 3320 5124
rect 3324 5064 3328 5124
rect 3385 5064 3389 5084
rect 3452 5064 3456 5084
rect 3474 5064 3478 5104
rect 3482 5064 3486 5104
rect 3545 5064 3549 5084
rect 3565 5064 3569 5084
rect 3611 5064 3615 5104
rect 3631 5064 3635 5104
rect 3651 5064 3655 5104
rect 3725 5064 3729 5104
rect 3745 5064 3749 5104
rect 3765 5064 3769 5104
rect 3811 5064 3815 5084
rect 3831 5064 3835 5084
rect 3893 5064 3897 5104
rect 3903 5064 3907 5104
rect 3993 5064 3997 5104
rect 4003 5064 4007 5104
rect 4051 5064 4055 5104
rect 4071 5064 4075 5104
rect 4091 5064 4095 5104
rect 4173 5064 4177 5104
rect 4183 5064 4187 5104
rect 4255 5064 4259 5104
rect 4275 5064 4279 5104
rect 4285 5064 4289 5104
rect 4353 5064 4357 5104
rect 4363 5064 4367 5104
rect 4425 5064 4429 5104
rect 4445 5064 4449 5104
rect 4465 5064 4469 5104
rect 4525 5064 4529 5104
rect 4545 5064 4549 5104
rect 4565 5064 4569 5104
rect 4613 5064 4617 5104
rect 4623 5064 4627 5104
rect 4693 5064 4697 5104
rect 4703 5064 4707 5104
rect 4771 5064 4775 5084
rect 4868 5064 4872 5124
rect 4876 5064 4880 5124
rect 4884 5064 4888 5124
rect 4931 5064 4935 5104
rect 4951 5064 4955 5104
rect 4971 5064 4975 5104
rect 5031 5064 5035 5104
rect 5093 5064 5097 5104
rect 5103 5064 5107 5104
rect 5171 5064 5175 5104
rect 5191 5064 5195 5104
rect 5253 5064 5257 5104
rect 5263 5064 5267 5104
rect 5331 5064 5335 5104
rect 5351 5064 5355 5104
rect 5371 5064 5375 5104
rect 5432 5064 5436 5124
rect 5440 5064 5444 5124
rect 5448 5064 5452 5124
rect 5532 5064 5536 5124
rect 5540 5064 5544 5124
rect 5548 5064 5552 5124
rect 5631 5064 5635 5084
rect 5692 5064 5696 5124
rect 5700 5064 5704 5124
rect 5708 5064 5712 5124
rect 5791 5064 5795 5104
rect 5811 5064 5815 5104
rect 5831 5064 5835 5104
rect 5913 5064 5917 5104
rect 5923 5064 5927 5104
rect 5972 5064 5976 5124
rect 5980 5064 5984 5124
rect 5988 5064 5992 5124
rect 6073 5064 6077 5104
rect 6083 5064 6087 5104
rect 6172 5064 6176 5084
rect 6194 5064 6198 5104
rect 6202 5064 6206 5104
rect 6265 5064 6269 5084
rect 6348 5064 6352 5124
rect 6356 5064 6360 5124
rect 6364 5064 6368 5124
rect 6448 5064 6452 5124
rect 6456 5064 6460 5124
rect 6464 5064 6468 5124
rect 6511 5064 6515 5084
rect 6608 5064 6612 5124
rect 6616 5064 6620 5124
rect 6624 5064 6628 5124
rect 6673 5064 6677 5104
rect 6683 5064 6687 5104
rect 43 4996 47 5036
rect 65 5016 69 5036
rect 123 4996 127 5036
rect 145 5016 149 5036
rect 213 4996 217 5036
rect 223 4996 227 5036
rect 271 4996 275 5036
rect 293 5016 297 5036
rect 303 5016 307 5036
rect 323 5016 327 5036
rect 331 5016 335 5036
rect 377 5016 381 5036
rect 399 5016 403 5036
rect 409 5016 413 5036
rect 431 5016 435 5036
rect 441 5016 445 5036
rect 461 4996 465 5036
rect 532 5016 536 5036
rect 554 4996 558 5036
rect 562 4996 566 5036
rect 633 4996 637 5036
rect 643 4996 647 5036
rect 693 4996 697 5036
rect 703 4996 707 5036
rect 793 4996 797 5036
rect 803 4996 807 5036
rect 851 4996 855 5036
rect 873 5016 877 5036
rect 883 5016 887 5036
rect 903 5016 907 5036
rect 911 5016 915 5036
rect 957 5016 961 5036
rect 979 5016 983 5036
rect 989 5016 993 5036
rect 1011 5016 1015 5036
rect 1021 5016 1025 5036
rect 1041 4996 1045 5036
rect 1103 4996 1107 5036
rect 1125 5016 1129 5036
rect 1192 5016 1196 5036
rect 1214 4996 1218 5036
rect 1222 4996 1226 5036
rect 1293 4996 1297 5036
rect 1303 4996 1307 5036
rect 1363 4996 1367 5036
rect 1385 5016 1389 5036
rect 1433 4996 1437 5036
rect 1443 4996 1447 5036
rect 1533 4996 1537 5036
rect 1543 4996 1547 5036
rect 1605 4996 1609 5036
rect 1625 4996 1629 5036
rect 1645 4996 1649 5036
rect 1713 4996 1717 5036
rect 1723 4996 1727 5036
rect 1785 4996 1789 5036
rect 1805 4996 1809 5036
rect 1825 4996 1829 5036
rect 1873 4996 1877 5036
rect 1883 4996 1887 5036
rect 1965 4996 1969 5036
rect 1985 4996 1989 5036
rect 2005 4996 2009 5036
rect 2065 4996 2069 5036
rect 2085 4996 2089 5036
rect 2105 4996 2109 5036
rect 2175 4996 2179 5036
rect 2195 4996 2199 5036
rect 2205 4996 2209 5036
rect 2251 5016 2255 5036
rect 2325 5016 2329 5036
rect 2345 5016 2349 5036
rect 2405 4996 2409 5036
rect 2425 5016 2429 5036
rect 2445 5016 2449 5036
rect 2513 4996 2517 5036
rect 2523 4996 2527 5036
rect 2585 4996 2589 5036
rect 2605 4996 2609 5036
rect 2625 4996 2629 5036
rect 2685 4996 2689 5036
rect 2705 4996 2709 5036
rect 2725 4996 2729 5036
rect 2785 5016 2789 5036
rect 2831 4996 2835 5036
rect 2851 4996 2855 5036
rect 2871 4996 2875 5036
rect 2945 4996 2949 5036
rect 2965 4996 2969 5036
rect 2985 4996 2989 5036
rect 3045 4996 3049 5036
rect 3065 4996 3069 5036
rect 3085 4996 3089 5036
rect 3145 5016 3149 5036
rect 3165 5016 3169 5036
rect 3225 4996 3229 5036
rect 3293 4996 3297 5036
rect 3303 4996 3307 5036
rect 3365 4996 3369 5036
rect 3385 4996 3389 5036
rect 3405 4996 3409 5036
rect 3455 4996 3459 5036
rect 3475 5016 3479 5036
rect 3485 5016 3489 5036
rect 3507 5016 3511 5036
rect 3517 5016 3521 5036
rect 3539 5016 3543 5036
rect 3585 5016 3589 5036
rect 3593 5016 3597 5036
rect 3613 5016 3617 5036
rect 3623 5016 3627 5036
rect 3645 4996 3649 5036
rect 3691 4996 3695 5036
rect 3711 4996 3715 5036
rect 3731 4996 3735 5036
rect 3812 5016 3816 5036
rect 3834 4996 3838 5036
rect 3842 4996 3846 5036
rect 3928 4976 3932 5036
rect 3936 4976 3940 5036
rect 3944 4976 3948 5036
rect 4012 5016 4016 5036
rect 4034 4996 4038 5036
rect 4042 4996 4046 5036
rect 4105 4996 4109 5036
rect 4175 4996 4179 5036
rect 4195 4996 4199 5036
rect 4205 4996 4209 5036
rect 4273 4996 4277 5036
rect 4283 4996 4287 5036
rect 4331 4996 4335 5036
rect 4341 4996 4345 5036
rect 4361 4996 4365 5036
rect 4445 4996 4449 5036
rect 4465 4996 4469 5036
rect 4485 4996 4489 5036
rect 4532 4976 4536 5036
rect 4540 4976 4544 5036
rect 4548 4976 4552 5036
rect 4631 4996 4635 5036
rect 4651 4996 4655 5036
rect 4671 4996 4675 5036
rect 4753 4996 4757 5036
rect 4763 4996 4767 5036
rect 4835 4996 4839 5036
rect 4855 4996 4859 5036
rect 4865 4996 4869 5036
rect 4933 4996 4937 5036
rect 4943 4996 4947 5036
rect 4993 4996 4997 5036
rect 5003 4996 5007 5036
rect 5071 4996 5075 5036
rect 5081 4996 5085 5036
rect 5101 4996 5105 5036
rect 5193 4996 5197 5036
rect 5203 4996 5207 5036
rect 5275 4996 5279 5036
rect 5295 4996 5299 5036
rect 5305 4996 5309 5036
rect 5351 4996 5355 5036
rect 5361 4996 5365 5036
rect 5381 4996 5385 5036
rect 5486 4996 5490 5036
rect 5494 4996 5498 5036
rect 5514 4996 5518 5036
rect 5522 4996 5526 5036
rect 5593 4996 5597 5036
rect 5603 4996 5607 5036
rect 5652 4976 5656 5036
rect 5660 4976 5664 5036
rect 5668 4976 5672 5036
rect 5772 5016 5776 5036
rect 5794 4996 5798 5036
rect 5802 4996 5806 5036
rect 5888 4976 5892 5036
rect 5896 4976 5900 5036
rect 5904 4976 5908 5036
rect 5973 4996 5977 5036
rect 5983 4996 5987 5036
rect 6034 4996 6038 5036
rect 6042 4996 6046 5036
rect 6062 4996 6066 5036
rect 6070 4996 6074 5036
rect 6188 4976 6192 5036
rect 6196 4976 6200 5036
rect 6204 4976 6208 5036
rect 6251 4996 6255 5036
rect 6271 4996 6275 5036
rect 6291 4996 6295 5036
rect 6388 4976 6392 5036
rect 6396 4976 6400 5036
rect 6404 4976 6408 5036
rect 6488 4976 6492 5036
rect 6496 4976 6500 5036
rect 6504 4976 6508 5036
rect 6553 4996 6557 5036
rect 6563 4996 6567 5036
rect 6645 5016 6649 5036
rect 31 4584 35 4624
rect 51 4584 55 4624
rect 71 4584 75 4624
rect 91 4584 95 4624
rect 111 4584 115 4624
rect 131 4584 135 4624
rect 151 4584 155 4624
rect 171 4584 175 4624
rect 245 4584 249 4604
rect 265 4584 269 4604
rect 325 4584 329 4604
rect 392 4584 396 4604
rect 414 4584 418 4624
rect 422 4584 426 4624
rect 485 4584 489 4604
rect 545 4584 549 4604
rect 565 4584 569 4604
rect 635 4584 639 4624
rect 655 4584 659 4624
rect 665 4584 669 4624
rect 711 4584 715 4604
rect 731 4584 735 4604
rect 803 4584 807 4624
rect 825 4584 829 4604
rect 893 4584 897 4624
rect 903 4584 907 4624
rect 951 4584 955 4624
rect 973 4584 977 4604
rect 983 4584 987 4604
rect 1003 4584 1007 4604
rect 1011 4584 1015 4604
rect 1057 4584 1061 4604
rect 1079 4584 1083 4604
rect 1089 4584 1093 4604
rect 1111 4584 1115 4604
rect 1121 4584 1125 4604
rect 1141 4584 1145 4624
rect 1205 4584 1209 4624
rect 1225 4584 1229 4624
rect 1245 4584 1249 4624
rect 1313 4584 1317 4624
rect 1323 4584 1327 4624
rect 1373 4584 1377 4624
rect 1383 4584 1387 4624
rect 1465 4584 1469 4624
rect 1485 4584 1489 4624
rect 1505 4584 1509 4624
rect 1551 4584 1555 4604
rect 1571 4584 1575 4604
rect 1631 4584 1635 4604
rect 1651 4584 1655 4604
rect 1711 4584 1715 4604
rect 1771 4584 1775 4604
rect 1791 4584 1795 4604
rect 1851 4584 1855 4624
rect 1871 4584 1875 4624
rect 1891 4584 1895 4624
rect 1951 4584 1955 4624
rect 1973 4584 1977 4604
rect 1983 4584 1987 4604
rect 2003 4584 2007 4604
rect 2011 4584 2015 4604
rect 2057 4584 2061 4604
rect 2079 4584 2083 4604
rect 2089 4584 2093 4604
rect 2111 4584 2115 4604
rect 2121 4584 2125 4604
rect 2141 4584 2145 4624
rect 2213 4584 2217 4624
rect 2223 4584 2227 4624
rect 2285 4584 2289 4624
rect 2305 4584 2309 4604
rect 2325 4584 2329 4604
rect 2373 4584 2377 4624
rect 2383 4584 2387 4624
rect 2451 4584 2455 4604
rect 2471 4584 2475 4604
rect 2534 4584 2538 4624
rect 2542 4584 2546 4624
rect 2564 4584 2568 4604
rect 2645 4584 2649 4604
rect 2691 4584 2695 4624
rect 2713 4584 2717 4604
rect 2723 4584 2727 4604
rect 2743 4584 2747 4604
rect 2751 4584 2755 4604
rect 2797 4584 2801 4604
rect 2819 4584 2823 4604
rect 2829 4584 2833 4604
rect 2851 4584 2855 4604
rect 2861 4584 2865 4604
rect 2881 4584 2885 4624
rect 2931 4584 2935 4624
rect 2951 4584 2955 4624
rect 2971 4584 2975 4624
rect 3031 4584 3035 4624
rect 3053 4584 3057 4604
rect 3063 4584 3067 4604
rect 3083 4584 3087 4604
rect 3091 4584 3095 4604
rect 3137 4584 3141 4604
rect 3159 4584 3163 4604
rect 3169 4584 3173 4604
rect 3191 4584 3195 4604
rect 3201 4584 3205 4604
rect 3221 4584 3225 4624
rect 3271 4584 3275 4624
rect 3293 4584 3297 4604
rect 3303 4584 3307 4604
rect 3323 4584 3327 4604
rect 3331 4584 3335 4604
rect 3377 4584 3381 4604
rect 3399 4584 3403 4604
rect 3409 4584 3413 4604
rect 3431 4584 3435 4604
rect 3441 4584 3445 4604
rect 3461 4584 3465 4624
rect 3525 4584 3529 4624
rect 3545 4584 3549 4624
rect 3565 4584 3569 4624
rect 3625 4584 3629 4624
rect 3693 4584 3697 4624
rect 3703 4584 3707 4624
rect 3765 4584 3769 4624
rect 3785 4584 3789 4624
rect 3805 4584 3809 4624
rect 3855 4584 3859 4624
rect 3875 4584 3879 4604
rect 3885 4584 3889 4604
rect 3907 4584 3911 4604
rect 3917 4584 3921 4604
rect 3939 4584 3943 4604
rect 3985 4584 3989 4604
rect 3993 4584 3997 4604
rect 4013 4584 4017 4604
rect 4023 4584 4027 4604
rect 4045 4584 4049 4624
rect 4105 4584 4109 4624
rect 4173 4584 4177 4624
rect 4183 4584 4187 4624
rect 4231 4584 4235 4624
rect 4253 4584 4257 4604
rect 4263 4584 4267 4604
rect 4283 4584 4287 4604
rect 4291 4584 4295 4604
rect 4337 4584 4341 4604
rect 4359 4584 4363 4604
rect 4369 4584 4373 4604
rect 4391 4584 4395 4604
rect 4401 4584 4405 4604
rect 4421 4584 4425 4624
rect 4508 4584 4512 4644
rect 4516 4584 4520 4644
rect 4524 4584 4528 4644
rect 4571 4584 4575 4604
rect 4631 4584 4635 4624
rect 4705 4584 4709 4604
rect 4751 4584 4755 4624
rect 4771 4584 4775 4624
rect 4791 4584 4795 4624
rect 4851 4584 4855 4604
rect 4871 4584 4875 4604
rect 4933 4584 4937 4624
rect 4943 4584 4947 4624
rect 5013 4584 5017 4624
rect 5023 4584 5027 4624
rect 5113 4584 5117 4624
rect 5123 4584 5127 4624
rect 5171 4584 5175 4624
rect 5191 4584 5195 4624
rect 5211 4584 5215 4624
rect 5285 4584 5289 4624
rect 5305 4584 5309 4624
rect 5325 4584 5329 4624
rect 5345 4584 5349 4624
rect 5393 4584 5397 4624
rect 5403 4584 5407 4624
rect 5493 4584 5497 4624
rect 5503 4584 5507 4624
rect 5552 4584 5556 4644
rect 5560 4584 5564 4644
rect 5568 4584 5572 4644
rect 5673 4584 5677 4624
rect 5683 4584 5687 4624
rect 5732 4584 5736 4644
rect 5740 4584 5744 4644
rect 5748 4584 5752 4644
rect 5845 4584 5849 4604
rect 5892 4584 5896 4644
rect 5900 4584 5904 4644
rect 5908 4584 5912 4644
rect 6015 4584 6019 4624
rect 6035 4584 6039 4624
rect 6045 4584 6049 4624
rect 6091 4584 6095 4624
rect 6111 4584 6115 4624
rect 6131 4584 6135 4624
rect 6213 4584 6217 4624
rect 6223 4584 6227 4624
rect 6274 4584 6278 4624
rect 6282 4584 6286 4624
rect 6304 4584 6308 4604
rect 6372 4584 6376 4644
rect 6380 4584 6384 4644
rect 6388 4584 6392 4644
rect 6495 4584 6499 4624
rect 6515 4584 6519 4624
rect 6525 4584 6529 4624
rect 6608 4584 6612 4644
rect 6616 4584 6620 4644
rect 6624 4584 6628 4644
rect 45 4536 49 4556
rect 105 4536 109 4556
rect 125 4536 129 4556
rect 185 4536 189 4556
rect 231 4516 235 4556
rect 251 4516 255 4556
rect 271 4516 275 4556
rect 345 4536 349 4556
rect 365 4536 369 4556
rect 411 4516 415 4556
rect 431 4516 435 4556
rect 451 4516 455 4556
rect 511 4536 515 4556
rect 531 4536 535 4556
rect 551 4516 555 4556
rect 614 4516 618 4556
rect 622 4516 626 4556
rect 644 4536 648 4556
rect 725 4536 729 4556
rect 771 4536 775 4556
rect 791 4536 795 4556
rect 851 4536 855 4556
rect 911 4536 915 4556
rect 931 4536 935 4556
rect 991 4536 995 4556
rect 1051 4516 1055 4556
rect 1071 4516 1075 4556
rect 1091 4516 1095 4556
rect 1111 4516 1115 4556
rect 1131 4516 1135 4556
rect 1151 4516 1155 4556
rect 1171 4516 1175 4556
rect 1191 4516 1195 4556
rect 1251 4536 1255 4556
rect 1273 4516 1277 4556
rect 1345 4536 1349 4556
rect 1405 4536 1409 4556
rect 1425 4536 1429 4556
rect 1493 4516 1497 4556
rect 1503 4516 1507 4556
rect 1553 4516 1557 4556
rect 1563 4516 1567 4556
rect 1645 4516 1649 4556
rect 1665 4516 1669 4556
rect 1685 4516 1689 4556
rect 1705 4516 1709 4556
rect 1755 4516 1759 4556
rect 1775 4536 1779 4556
rect 1785 4536 1789 4556
rect 1807 4536 1811 4556
rect 1817 4536 1821 4556
rect 1839 4536 1843 4556
rect 1885 4536 1889 4556
rect 1893 4536 1897 4556
rect 1913 4536 1917 4556
rect 1923 4536 1927 4556
rect 1945 4516 1949 4556
rect 1993 4516 1997 4556
rect 2003 4516 2007 4556
rect 2071 4516 2075 4556
rect 2093 4536 2097 4556
rect 2103 4536 2107 4556
rect 2123 4536 2127 4556
rect 2131 4536 2135 4556
rect 2177 4536 2181 4556
rect 2199 4536 2203 4556
rect 2209 4536 2213 4556
rect 2231 4536 2235 4556
rect 2241 4536 2245 4556
rect 2261 4516 2265 4556
rect 2311 4536 2315 4556
rect 2371 4536 2375 4556
rect 2391 4536 2395 4556
rect 2451 4536 2455 4556
rect 2471 4536 2475 4556
rect 2531 4536 2535 4556
rect 2591 4516 2595 4556
rect 2613 4536 2617 4556
rect 2623 4536 2627 4556
rect 2643 4536 2647 4556
rect 2651 4536 2655 4556
rect 2697 4536 2701 4556
rect 2719 4536 2723 4556
rect 2729 4536 2733 4556
rect 2751 4536 2755 4556
rect 2761 4536 2765 4556
rect 2781 4516 2785 4556
rect 2831 4516 2835 4556
rect 2851 4516 2855 4556
rect 2871 4516 2875 4556
rect 2933 4516 2937 4556
rect 2943 4516 2947 4556
rect 3025 4536 3029 4556
rect 3071 4516 3075 4556
rect 3091 4516 3095 4556
rect 3111 4516 3115 4556
rect 3171 4516 3175 4556
rect 3193 4536 3197 4556
rect 3203 4536 3207 4556
rect 3223 4536 3227 4556
rect 3231 4536 3235 4556
rect 3277 4536 3281 4556
rect 3299 4536 3303 4556
rect 3309 4536 3313 4556
rect 3331 4536 3335 4556
rect 3341 4536 3345 4556
rect 3361 4516 3365 4556
rect 3411 4516 3415 4556
rect 3431 4516 3435 4556
rect 3451 4516 3455 4556
rect 3525 4516 3529 4556
rect 3545 4516 3549 4556
rect 3565 4516 3569 4556
rect 3615 4516 3619 4556
rect 3635 4536 3639 4556
rect 3645 4536 3649 4556
rect 3667 4536 3671 4556
rect 3677 4536 3681 4556
rect 3699 4536 3703 4556
rect 3745 4536 3749 4556
rect 3753 4536 3757 4556
rect 3773 4536 3777 4556
rect 3783 4536 3787 4556
rect 3805 4516 3809 4556
rect 3851 4516 3855 4556
rect 3871 4516 3875 4556
rect 3891 4516 3895 4556
rect 3955 4516 3959 4556
rect 3975 4536 3979 4556
rect 3985 4536 3989 4556
rect 4007 4536 4011 4556
rect 4017 4536 4021 4556
rect 4039 4536 4043 4556
rect 4085 4536 4089 4556
rect 4093 4536 4097 4556
rect 4113 4536 4117 4556
rect 4123 4536 4127 4556
rect 4145 4516 4149 4556
rect 4228 4496 4232 4556
rect 4236 4496 4240 4556
rect 4244 4496 4248 4556
rect 4291 4516 4295 4556
rect 4311 4516 4315 4556
rect 4331 4516 4335 4556
rect 4405 4536 4409 4556
rect 4425 4536 4429 4556
rect 4492 4536 4496 4556
rect 4514 4516 4518 4556
rect 4522 4516 4526 4556
rect 4572 4496 4576 4556
rect 4580 4496 4584 4556
rect 4588 4496 4592 4556
rect 4685 4536 4689 4556
rect 4731 4516 4735 4556
rect 4751 4516 4755 4556
rect 4771 4516 4775 4556
rect 4845 4516 4849 4556
rect 4865 4536 4869 4556
rect 4885 4536 4889 4556
rect 4953 4516 4957 4556
rect 4963 4516 4967 4556
rect 5048 4496 5052 4556
rect 5056 4496 5060 4556
rect 5064 4496 5068 4556
rect 5111 4516 5115 4556
rect 5131 4516 5135 4556
rect 5151 4516 5155 4556
rect 5225 4516 5229 4556
rect 5245 4536 5249 4556
rect 5265 4536 5269 4556
rect 5311 4516 5315 4556
rect 5331 4516 5335 4556
rect 5351 4516 5355 4556
rect 5411 4536 5415 4556
rect 5508 4496 5512 4556
rect 5516 4496 5520 4556
rect 5524 4496 5528 4556
rect 5573 4516 5577 4556
rect 5583 4516 5587 4556
rect 5651 4516 5655 4556
rect 5671 4516 5675 4556
rect 5691 4516 5695 4556
rect 5773 4516 5777 4556
rect 5783 4516 5787 4556
rect 5868 4496 5872 4556
rect 5876 4496 5880 4556
rect 5884 4496 5888 4556
rect 5945 4516 5949 4556
rect 5965 4516 5969 4556
rect 5985 4516 5989 4556
rect 6031 4536 6035 4556
rect 6105 4536 6109 4556
rect 6152 4496 6156 4556
rect 6160 4496 6164 4556
rect 6168 4496 6172 4556
rect 6265 4516 6269 4556
rect 6285 4516 6289 4556
rect 6305 4516 6309 4556
rect 6352 4496 6356 4556
rect 6360 4496 6364 4556
rect 6368 4496 6372 4556
rect 6452 4496 6456 4556
rect 6460 4496 6464 4556
rect 6468 4496 6472 4556
rect 6551 4516 6555 4556
rect 6571 4516 6575 4556
rect 6591 4516 6595 4556
rect 6651 4536 6655 4556
rect 43 4104 47 4144
rect 65 4104 69 4124
rect 125 4104 129 4144
rect 145 4104 149 4144
rect 165 4104 169 4144
rect 211 4104 215 4144
rect 231 4104 235 4144
rect 251 4104 255 4144
rect 315 4104 319 4144
rect 335 4104 339 4124
rect 345 4104 349 4124
rect 367 4104 371 4124
rect 377 4104 381 4124
rect 399 4104 403 4124
rect 445 4104 449 4124
rect 453 4104 457 4124
rect 473 4104 477 4124
rect 483 4104 487 4124
rect 505 4104 509 4144
rect 553 4104 557 4144
rect 563 4104 567 4144
rect 666 4104 670 4144
rect 674 4104 678 4144
rect 694 4104 698 4144
rect 702 4104 706 4144
rect 765 4104 769 4124
rect 811 4104 815 4144
rect 833 4104 837 4124
rect 843 4104 847 4124
rect 863 4104 867 4124
rect 871 4104 875 4124
rect 917 4104 921 4124
rect 939 4104 943 4124
rect 949 4104 953 4124
rect 971 4104 975 4124
rect 981 4104 985 4124
rect 1001 4104 1005 4144
rect 1053 4104 1057 4144
rect 1063 4104 1067 4144
rect 1131 4104 1135 4144
rect 1153 4104 1157 4124
rect 1163 4104 1167 4124
rect 1183 4104 1187 4124
rect 1191 4104 1195 4124
rect 1237 4104 1241 4124
rect 1259 4104 1263 4124
rect 1269 4104 1273 4124
rect 1291 4104 1295 4124
rect 1301 4104 1305 4124
rect 1321 4104 1325 4144
rect 1373 4104 1377 4144
rect 1383 4104 1387 4144
rect 1451 4104 1455 4124
rect 1525 4104 1529 4144
rect 1545 4104 1549 4144
rect 1565 4104 1569 4144
rect 1632 4104 1636 4124
rect 1654 4104 1658 4144
rect 1662 4104 1666 4144
rect 1733 4104 1737 4144
rect 1743 4104 1747 4144
rect 1793 4104 1797 4144
rect 1803 4104 1807 4144
rect 1871 4104 1875 4144
rect 1893 4104 1897 4124
rect 1903 4104 1907 4124
rect 1923 4104 1927 4124
rect 1931 4104 1935 4124
rect 1977 4104 1981 4124
rect 1999 4104 2003 4124
rect 2009 4104 2013 4124
rect 2031 4104 2035 4124
rect 2041 4104 2045 4124
rect 2061 4104 2065 4144
rect 2113 4104 2117 4144
rect 2123 4104 2127 4144
rect 2205 4104 2209 4144
rect 2225 4104 2229 4144
rect 2245 4104 2249 4144
rect 2295 4104 2299 4144
rect 2315 4104 2319 4124
rect 2325 4104 2329 4124
rect 2347 4104 2351 4124
rect 2357 4104 2361 4124
rect 2379 4104 2383 4124
rect 2425 4104 2429 4124
rect 2433 4104 2437 4124
rect 2453 4104 2457 4124
rect 2463 4104 2467 4124
rect 2485 4104 2489 4144
rect 2545 4104 2549 4124
rect 2565 4104 2569 4124
rect 2611 4104 2615 4124
rect 2671 4104 2675 4144
rect 2691 4104 2695 4144
rect 2711 4104 2715 4144
rect 2773 4104 2777 4144
rect 2783 4104 2787 4144
rect 2865 4104 2869 4144
rect 2885 4104 2889 4144
rect 2905 4104 2909 4144
rect 2951 4104 2955 4124
rect 3011 4104 3015 4124
rect 3031 4104 3035 4124
rect 3105 4104 3109 4124
rect 3151 4104 3155 4144
rect 3173 4104 3177 4124
rect 3183 4104 3187 4124
rect 3203 4104 3207 4124
rect 3211 4104 3215 4124
rect 3257 4104 3261 4124
rect 3279 4104 3283 4124
rect 3289 4104 3293 4124
rect 3311 4104 3315 4124
rect 3321 4104 3325 4124
rect 3341 4104 3345 4144
rect 3391 4104 3395 4144
rect 3411 4104 3415 4144
rect 3431 4104 3435 4144
rect 3451 4104 3455 4144
rect 3513 4104 3517 4144
rect 3523 4104 3527 4144
rect 3591 4104 3595 4144
rect 3611 4104 3615 4144
rect 3631 4104 3635 4144
rect 3651 4104 3655 4144
rect 3671 4104 3675 4144
rect 3691 4104 3695 4144
rect 3711 4104 3715 4144
rect 3731 4104 3735 4144
rect 3793 4104 3797 4144
rect 3803 4104 3807 4144
rect 3873 4104 3877 4144
rect 3883 4104 3887 4144
rect 3973 4104 3977 4144
rect 3983 4104 3987 4144
rect 4031 4104 4035 4124
rect 4105 4104 4109 4144
rect 4125 4104 4129 4144
rect 4145 4104 4149 4144
rect 4191 4104 4195 4144
rect 4211 4104 4215 4144
rect 4231 4104 4235 4144
rect 4295 4104 4299 4144
rect 4315 4104 4319 4124
rect 4325 4104 4329 4124
rect 4347 4104 4351 4124
rect 4357 4104 4361 4124
rect 4379 4104 4383 4124
rect 4425 4104 4429 4124
rect 4433 4104 4437 4124
rect 4453 4104 4457 4124
rect 4463 4104 4467 4124
rect 4485 4104 4489 4144
rect 4545 4104 4549 4144
rect 4565 4104 4569 4144
rect 4585 4104 4589 4144
rect 4635 4104 4639 4144
rect 4655 4104 4659 4124
rect 4665 4104 4669 4124
rect 4687 4104 4691 4124
rect 4697 4104 4701 4124
rect 4719 4104 4723 4124
rect 4765 4104 4769 4124
rect 4773 4104 4777 4124
rect 4793 4104 4797 4124
rect 4803 4104 4807 4124
rect 4825 4104 4829 4144
rect 4885 4104 4889 4144
rect 4952 4104 4956 4124
rect 4974 4104 4978 4144
rect 4982 4104 4986 4144
rect 5032 4104 5036 4164
rect 5040 4104 5044 4164
rect 5048 4104 5052 4164
rect 5145 4104 5149 4124
rect 5191 4104 5195 4144
rect 5211 4104 5215 4144
rect 5231 4104 5235 4144
rect 5295 4104 5299 4144
rect 5315 4104 5319 4124
rect 5325 4104 5329 4124
rect 5347 4104 5351 4124
rect 5357 4104 5361 4124
rect 5379 4104 5383 4124
rect 5425 4104 5429 4124
rect 5433 4104 5437 4124
rect 5453 4104 5457 4124
rect 5463 4104 5467 4124
rect 5485 4104 5489 4144
rect 5533 4104 5537 4144
rect 5543 4104 5547 4144
rect 5611 4104 5615 4124
rect 5671 4104 5675 4144
rect 5691 4104 5695 4144
rect 5711 4104 5715 4144
rect 5795 4104 5799 4144
rect 5815 4104 5819 4144
rect 5825 4104 5829 4144
rect 5872 4104 5876 4164
rect 5880 4104 5884 4164
rect 5888 4104 5892 4164
rect 5985 4104 5989 4144
rect 6031 4104 6035 4144
rect 6051 4104 6055 4144
rect 6071 4104 6075 4144
rect 6131 4104 6135 4124
rect 6153 4104 6157 4144
rect 6213 4104 6217 4144
rect 6223 4104 6227 4144
rect 6315 4104 6319 4144
rect 6335 4104 6339 4144
rect 6345 4104 6349 4144
rect 6393 4104 6397 4144
rect 6403 4104 6407 4144
rect 6471 4104 6475 4124
rect 6552 4104 6556 4124
rect 6574 4104 6578 4144
rect 6582 4104 6586 4144
rect 6632 4104 6636 4164
rect 6640 4104 6644 4164
rect 6648 4104 6652 4164
rect 43 4036 47 4076
rect 65 4056 69 4076
rect 111 4036 115 4076
rect 133 4056 137 4076
rect 143 4056 147 4076
rect 163 4056 167 4076
rect 171 4056 175 4076
rect 217 4056 221 4076
rect 239 4056 243 4076
rect 249 4056 253 4076
rect 271 4056 275 4076
rect 281 4056 285 4076
rect 301 4036 305 4076
rect 353 4036 357 4076
rect 363 4036 367 4076
rect 452 4056 456 4076
rect 474 4036 478 4076
rect 482 4036 486 4076
rect 553 4036 557 4076
rect 563 4036 567 4076
rect 633 4036 637 4076
rect 643 4036 647 4076
rect 703 4036 707 4076
rect 725 4056 729 4076
rect 771 4036 775 4076
rect 793 4056 797 4076
rect 803 4056 807 4076
rect 823 4056 827 4076
rect 831 4056 835 4076
rect 877 4056 881 4076
rect 899 4056 903 4076
rect 909 4056 913 4076
rect 931 4056 935 4076
rect 941 4056 945 4076
rect 961 4036 965 4076
rect 1033 4036 1037 4076
rect 1043 4036 1047 4076
rect 1093 4036 1097 4076
rect 1103 4036 1107 4076
rect 1173 4036 1177 4076
rect 1183 4036 1187 4076
rect 1272 4056 1276 4076
rect 1294 4036 1298 4076
rect 1302 4036 1306 4076
rect 1351 4036 1355 4076
rect 1373 4056 1377 4076
rect 1383 4056 1387 4076
rect 1403 4056 1407 4076
rect 1411 4056 1415 4076
rect 1457 4056 1461 4076
rect 1479 4056 1483 4076
rect 1489 4056 1493 4076
rect 1511 4056 1515 4076
rect 1521 4056 1525 4076
rect 1541 4036 1545 4076
rect 1613 4036 1617 4076
rect 1623 4036 1627 4076
rect 1671 4056 1675 4076
rect 1693 4036 1697 4076
rect 1753 4036 1757 4076
rect 1763 4036 1767 4076
rect 1831 4036 1835 4076
rect 1853 4056 1857 4076
rect 1863 4056 1867 4076
rect 1883 4056 1887 4076
rect 1891 4056 1895 4076
rect 1937 4056 1941 4076
rect 1959 4056 1963 4076
rect 1969 4056 1973 4076
rect 1991 4056 1995 4076
rect 2001 4056 2005 4076
rect 2021 4036 2025 4076
rect 2073 4036 2077 4076
rect 2083 4036 2087 4076
rect 2165 4036 2169 4076
rect 2185 4036 2189 4076
rect 2205 4036 2209 4076
rect 2273 4036 2277 4076
rect 2283 4036 2287 4076
rect 2333 4036 2337 4076
rect 2343 4036 2347 4076
rect 2425 4056 2429 4076
rect 2485 4036 2489 4076
rect 2505 4036 2509 4076
rect 2525 4036 2529 4076
rect 2571 4056 2575 4076
rect 2591 4056 2595 4076
rect 2665 4056 2669 4076
rect 2685 4056 2689 4076
rect 2731 4056 2735 4076
rect 2805 4056 2809 4076
rect 2873 4036 2877 4076
rect 2883 4036 2887 4076
rect 2931 4056 2935 4076
rect 2951 4056 2955 4076
rect 3011 4036 3015 4076
rect 3031 4036 3035 4076
rect 3051 4036 3055 4076
rect 3111 4056 3115 4076
rect 3171 4056 3175 4076
rect 3191 4056 3195 4076
rect 3273 4036 3277 4076
rect 3283 4036 3287 4076
rect 3353 4036 3357 4076
rect 3363 4036 3367 4076
rect 3415 4036 3419 4076
rect 3435 4056 3439 4076
rect 3445 4056 3449 4076
rect 3467 4056 3471 4076
rect 3477 4056 3481 4076
rect 3499 4056 3503 4076
rect 3545 4056 3549 4076
rect 3553 4056 3557 4076
rect 3573 4056 3577 4076
rect 3583 4056 3587 4076
rect 3605 4036 3609 4076
rect 3665 4056 3669 4076
rect 3715 4036 3719 4076
rect 3735 4056 3739 4076
rect 3745 4056 3749 4076
rect 3767 4056 3771 4076
rect 3777 4056 3781 4076
rect 3799 4056 3803 4076
rect 3845 4056 3849 4076
rect 3853 4056 3857 4076
rect 3873 4056 3877 4076
rect 3883 4056 3887 4076
rect 3905 4036 3909 4076
rect 3988 4016 3992 4076
rect 3996 4016 4000 4076
rect 4004 4016 4008 4076
rect 4053 4036 4057 4076
rect 4063 4036 4067 4076
rect 4145 4036 4149 4076
rect 4165 4036 4169 4076
rect 4185 4036 4189 4076
rect 4231 4056 4235 4076
rect 4251 4056 4255 4076
rect 4325 4056 4329 4076
rect 4393 4036 4397 4076
rect 4403 4036 4407 4076
rect 4465 4036 4469 4076
rect 4485 4036 4489 4076
rect 4505 4036 4509 4076
rect 4555 4036 4559 4076
rect 4575 4056 4579 4076
rect 4585 4056 4589 4076
rect 4607 4056 4611 4076
rect 4617 4056 4621 4076
rect 4639 4056 4643 4076
rect 4685 4056 4689 4076
rect 4693 4056 4697 4076
rect 4713 4056 4717 4076
rect 4723 4056 4727 4076
rect 4745 4036 4749 4076
rect 4813 4036 4817 4076
rect 4823 4036 4827 4076
rect 4885 4036 4889 4076
rect 4905 4036 4909 4076
rect 4925 4036 4929 4076
rect 4975 4036 4979 4076
rect 4995 4056 4999 4076
rect 5005 4056 5009 4076
rect 5027 4056 5031 4076
rect 5037 4056 5041 4076
rect 5059 4056 5063 4076
rect 5105 4056 5109 4076
rect 5113 4056 5117 4076
rect 5133 4056 5137 4076
rect 5143 4056 5147 4076
rect 5165 4036 5169 4076
rect 5233 4036 5237 4076
rect 5243 4036 5247 4076
rect 5305 4036 5309 4076
rect 5325 4036 5329 4076
rect 5345 4036 5349 4076
rect 5413 4036 5417 4076
rect 5423 4036 5427 4076
rect 5471 4036 5475 4076
rect 5491 4036 5495 4076
rect 5511 4036 5515 4076
rect 5585 4056 5589 4076
rect 5635 4036 5639 4076
rect 5655 4056 5659 4076
rect 5665 4056 5669 4076
rect 5687 4056 5691 4076
rect 5697 4056 5701 4076
rect 5719 4056 5723 4076
rect 5765 4056 5769 4076
rect 5773 4056 5777 4076
rect 5793 4056 5797 4076
rect 5803 4056 5807 4076
rect 5825 4036 5829 4076
rect 5871 4056 5875 4076
rect 5968 4016 5972 4076
rect 5976 4016 5980 4076
rect 5984 4016 5988 4076
rect 6031 4036 6035 4076
rect 6053 4056 6057 4076
rect 6063 4056 6067 4076
rect 6083 4056 6087 4076
rect 6091 4056 6095 4076
rect 6137 4056 6141 4076
rect 6159 4056 6163 4076
rect 6169 4056 6173 4076
rect 6191 4056 6195 4076
rect 6201 4056 6205 4076
rect 6221 4036 6225 4076
rect 6271 4036 6275 4076
rect 6293 4056 6297 4076
rect 6303 4056 6307 4076
rect 6323 4056 6327 4076
rect 6331 4056 6335 4076
rect 6377 4056 6381 4076
rect 6399 4056 6403 4076
rect 6409 4056 6413 4076
rect 6431 4056 6435 4076
rect 6441 4056 6445 4076
rect 6461 4036 6465 4076
rect 6511 4036 6515 4076
rect 6533 4056 6537 4076
rect 6543 4056 6547 4076
rect 6563 4056 6567 4076
rect 6571 4056 6575 4076
rect 6617 4056 6621 4076
rect 6639 4056 6643 4076
rect 6649 4056 6653 4076
rect 6671 4056 6675 4076
rect 6681 4056 6685 4076
rect 6701 4036 6705 4076
rect 43 3624 47 3664
rect 65 3624 69 3644
rect 123 3624 127 3664
rect 145 3624 149 3644
rect 213 3624 217 3664
rect 223 3624 227 3664
rect 271 3624 275 3664
rect 293 3624 297 3644
rect 303 3624 307 3644
rect 323 3624 327 3644
rect 331 3624 335 3644
rect 377 3624 381 3644
rect 399 3624 403 3644
rect 409 3624 413 3644
rect 431 3624 435 3644
rect 441 3624 445 3644
rect 461 3624 465 3664
rect 532 3624 536 3644
rect 554 3624 558 3664
rect 562 3624 566 3664
rect 633 3624 637 3664
rect 643 3624 647 3664
rect 693 3624 697 3664
rect 703 3624 707 3664
rect 793 3624 797 3664
rect 803 3624 807 3664
rect 851 3624 855 3664
rect 873 3624 877 3644
rect 883 3624 887 3644
rect 903 3624 907 3644
rect 911 3624 915 3644
rect 957 3624 961 3644
rect 979 3624 983 3644
rect 989 3624 993 3644
rect 1011 3624 1015 3644
rect 1021 3624 1025 3644
rect 1041 3624 1045 3664
rect 1094 3624 1098 3664
rect 1102 3624 1106 3664
rect 1124 3624 1128 3644
rect 1213 3624 1217 3664
rect 1223 3624 1227 3664
rect 1271 3624 1275 3644
rect 1293 3624 1297 3664
rect 1372 3624 1376 3644
rect 1394 3624 1398 3664
rect 1402 3624 1406 3664
rect 1473 3624 1477 3664
rect 1483 3624 1487 3664
rect 1533 3624 1537 3664
rect 1543 3624 1547 3664
rect 1611 3624 1615 3644
rect 1631 3624 1635 3644
rect 1691 3624 1695 3664
rect 1713 3624 1717 3644
rect 1723 3624 1727 3644
rect 1743 3624 1747 3644
rect 1751 3624 1755 3644
rect 1797 3624 1801 3644
rect 1819 3624 1823 3644
rect 1829 3624 1833 3644
rect 1851 3624 1855 3644
rect 1861 3624 1865 3644
rect 1881 3624 1885 3664
rect 1953 3624 1957 3664
rect 1963 3624 1967 3664
rect 2011 3624 2015 3644
rect 2031 3624 2035 3644
rect 2091 3624 2095 3644
rect 2151 3624 2155 3664
rect 2171 3624 2175 3664
rect 2191 3624 2195 3664
rect 2265 3624 2269 3664
rect 2285 3624 2289 3664
rect 2305 3624 2309 3664
rect 2372 3624 2376 3644
rect 2394 3624 2398 3664
rect 2402 3624 2406 3664
rect 2451 3624 2455 3644
rect 2525 3624 2529 3644
rect 2571 3624 2575 3664
rect 2591 3624 2595 3664
rect 2611 3624 2615 3664
rect 2672 3624 2676 3684
rect 2680 3624 2684 3684
rect 2688 3624 2692 3684
rect 2785 3624 2789 3644
rect 2853 3624 2857 3664
rect 2863 3624 2867 3664
rect 2911 3624 2915 3664
rect 2931 3624 2935 3664
rect 2951 3624 2955 3664
rect 3011 3624 3015 3664
rect 3031 3624 3035 3664
rect 3051 3624 3055 3664
rect 3114 3624 3118 3664
rect 3122 3624 3126 3664
rect 3144 3624 3148 3644
rect 3246 3624 3250 3664
rect 3254 3624 3258 3664
rect 3274 3624 3278 3664
rect 3282 3624 3286 3664
rect 3353 3624 3357 3664
rect 3363 3624 3367 3664
rect 3433 3624 3437 3664
rect 3443 3624 3447 3664
rect 3495 3624 3499 3664
rect 3515 3624 3519 3644
rect 3525 3624 3529 3644
rect 3547 3624 3551 3644
rect 3557 3624 3561 3644
rect 3579 3624 3583 3644
rect 3625 3624 3629 3644
rect 3633 3624 3637 3644
rect 3653 3624 3657 3644
rect 3663 3624 3667 3644
rect 3685 3624 3689 3664
rect 3753 3624 3757 3664
rect 3763 3624 3767 3664
rect 3846 3624 3850 3664
rect 3854 3624 3858 3664
rect 3874 3624 3878 3664
rect 3882 3624 3886 3664
rect 3931 3624 3935 3644
rect 3993 3624 3997 3664
rect 4003 3624 4007 3664
rect 4071 3624 4075 3664
rect 4091 3624 4095 3664
rect 4111 3624 4115 3664
rect 4175 3624 4179 3664
rect 4195 3624 4199 3644
rect 4205 3624 4209 3644
rect 4227 3624 4231 3644
rect 4237 3624 4241 3644
rect 4259 3624 4263 3644
rect 4305 3624 4309 3644
rect 4313 3624 4317 3644
rect 4333 3624 4337 3644
rect 4343 3624 4347 3644
rect 4365 3624 4369 3664
rect 4413 3624 4417 3664
rect 4423 3624 4427 3664
rect 4513 3624 4517 3664
rect 4523 3624 4527 3664
rect 4585 3624 4589 3664
rect 4605 3624 4609 3664
rect 4625 3624 4629 3664
rect 4645 3624 4649 3664
rect 4665 3624 4669 3664
rect 4685 3624 4689 3664
rect 4705 3624 4709 3664
rect 4725 3624 4729 3664
rect 4775 3624 4779 3664
rect 4795 3624 4799 3644
rect 4805 3624 4809 3644
rect 4827 3624 4831 3644
rect 4837 3624 4841 3644
rect 4859 3624 4863 3644
rect 4905 3624 4909 3644
rect 4913 3624 4917 3644
rect 4933 3624 4937 3644
rect 4943 3624 4947 3644
rect 4965 3624 4969 3664
rect 5011 3624 5015 3664
rect 5031 3624 5035 3664
rect 5051 3624 5055 3664
rect 5133 3624 5137 3664
rect 5143 3624 5147 3664
rect 5213 3624 5217 3664
rect 5223 3624 5227 3664
rect 5285 3624 5289 3644
rect 5331 3624 5335 3664
rect 5351 3624 5355 3664
rect 5371 3624 5375 3664
rect 5391 3624 5395 3664
rect 5411 3624 5415 3664
rect 5431 3624 5435 3664
rect 5451 3624 5455 3664
rect 5471 3624 5475 3664
rect 5531 3624 5535 3664
rect 5553 3624 5557 3644
rect 5563 3624 5567 3644
rect 5583 3624 5587 3644
rect 5591 3624 5595 3644
rect 5637 3624 5641 3644
rect 5659 3624 5663 3644
rect 5669 3624 5673 3644
rect 5691 3624 5695 3644
rect 5701 3624 5705 3644
rect 5721 3624 5725 3664
rect 5785 3624 5789 3644
rect 5833 3624 5837 3664
rect 5843 3624 5847 3664
rect 5913 3624 5917 3664
rect 5923 3624 5927 3664
rect 6005 3624 6009 3644
rect 6051 3624 6055 3644
rect 6071 3624 6075 3644
rect 6145 3624 6149 3644
rect 6165 3624 6169 3644
rect 6214 3624 6218 3664
rect 6222 3624 6226 3664
rect 6244 3624 6248 3644
rect 6311 3624 6315 3664
rect 6333 3624 6337 3644
rect 6343 3624 6347 3644
rect 6363 3624 6367 3644
rect 6371 3624 6375 3644
rect 6417 3624 6421 3644
rect 6439 3624 6443 3644
rect 6449 3624 6453 3644
rect 6471 3624 6475 3644
rect 6481 3624 6485 3644
rect 6501 3624 6505 3664
rect 6551 3624 6555 3664
rect 6571 3624 6575 3664
rect 6591 3624 6595 3664
rect 6653 3624 6657 3664
rect 6663 3624 6667 3664
rect 43 3556 47 3596
rect 65 3576 69 3596
rect 111 3556 115 3596
rect 133 3576 137 3596
rect 143 3576 147 3596
rect 163 3576 167 3596
rect 171 3576 175 3596
rect 217 3576 221 3596
rect 239 3576 243 3596
rect 249 3576 253 3596
rect 271 3576 275 3596
rect 281 3576 285 3596
rect 301 3556 305 3596
rect 353 3556 357 3596
rect 363 3556 367 3596
rect 431 3576 435 3596
rect 453 3556 457 3596
rect 532 3576 536 3596
rect 554 3556 558 3596
rect 562 3556 566 3596
rect 633 3556 637 3596
rect 643 3556 647 3596
rect 703 3556 707 3596
rect 725 3576 729 3596
rect 771 3576 775 3596
rect 793 3556 797 3596
rect 853 3556 857 3596
rect 863 3556 867 3596
rect 943 3556 947 3596
rect 965 3576 969 3596
rect 1025 3576 1029 3596
rect 1083 3556 1087 3596
rect 1105 3576 1109 3596
rect 1163 3556 1167 3596
rect 1185 3576 1189 3596
rect 1231 3556 1235 3596
rect 1253 3576 1257 3596
rect 1263 3576 1267 3596
rect 1283 3576 1287 3596
rect 1291 3576 1295 3596
rect 1337 3576 1341 3596
rect 1359 3576 1363 3596
rect 1369 3576 1373 3596
rect 1391 3576 1395 3596
rect 1401 3576 1405 3596
rect 1421 3556 1425 3596
rect 1485 3576 1489 3596
rect 1505 3576 1509 3596
rect 1551 3556 1555 3596
rect 1573 3576 1577 3596
rect 1583 3576 1587 3596
rect 1603 3576 1607 3596
rect 1611 3576 1615 3596
rect 1657 3576 1661 3596
rect 1679 3576 1683 3596
rect 1689 3576 1693 3596
rect 1711 3576 1715 3596
rect 1721 3576 1725 3596
rect 1741 3556 1745 3596
rect 1815 3556 1819 3596
rect 1835 3556 1839 3596
rect 1845 3556 1849 3596
rect 1905 3576 1909 3596
rect 1965 3556 1969 3596
rect 1985 3556 1989 3596
rect 2005 3556 2009 3596
rect 2051 3576 2055 3596
rect 2071 3576 2075 3596
rect 2145 3576 2149 3596
rect 2215 3556 2219 3596
rect 2235 3556 2239 3596
rect 2245 3556 2249 3596
rect 2305 3576 2309 3596
rect 2325 3576 2329 3596
rect 2371 3556 2375 3596
rect 2393 3576 2397 3596
rect 2403 3576 2407 3596
rect 2423 3576 2427 3596
rect 2431 3576 2435 3596
rect 2477 3576 2481 3596
rect 2499 3576 2503 3596
rect 2509 3576 2513 3596
rect 2531 3576 2535 3596
rect 2541 3576 2545 3596
rect 2561 3556 2565 3596
rect 2611 3576 2615 3596
rect 2631 3576 2635 3596
rect 2691 3556 2695 3596
rect 2711 3556 2715 3596
rect 2731 3556 2735 3596
rect 2805 3576 2809 3596
rect 2873 3556 2877 3596
rect 2883 3556 2887 3596
rect 2931 3556 2935 3596
rect 2951 3556 2955 3596
rect 2971 3556 2975 3596
rect 3034 3556 3038 3596
rect 3042 3556 3046 3596
rect 3064 3576 3068 3596
rect 3131 3556 3135 3596
rect 3226 3556 3230 3596
rect 3234 3556 3238 3596
rect 3254 3556 3258 3596
rect 3262 3556 3266 3596
rect 3325 3576 3329 3596
rect 3371 3556 3375 3596
rect 3393 3576 3397 3596
rect 3403 3576 3407 3596
rect 3423 3576 3427 3596
rect 3431 3576 3435 3596
rect 3477 3576 3481 3596
rect 3499 3576 3503 3596
rect 3509 3576 3513 3596
rect 3531 3576 3535 3596
rect 3541 3576 3545 3596
rect 3561 3556 3565 3596
rect 3646 3556 3650 3596
rect 3654 3556 3658 3596
rect 3674 3556 3678 3596
rect 3682 3556 3686 3596
rect 3731 3556 3735 3596
rect 3753 3576 3757 3596
rect 3763 3576 3767 3596
rect 3783 3576 3787 3596
rect 3791 3576 3795 3596
rect 3837 3576 3841 3596
rect 3859 3576 3863 3596
rect 3869 3576 3873 3596
rect 3891 3576 3895 3596
rect 3901 3576 3905 3596
rect 3921 3556 3925 3596
rect 3985 3576 3989 3596
rect 4031 3556 4035 3596
rect 4053 3576 4057 3596
rect 4063 3576 4067 3596
rect 4083 3576 4087 3596
rect 4091 3576 4095 3596
rect 4137 3576 4141 3596
rect 4159 3576 4163 3596
rect 4169 3576 4173 3596
rect 4191 3576 4195 3596
rect 4201 3576 4205 3596
rect 4221 3556 4225 3596
rect 4285 3576 4289 3596
rect 4345 3576 4349 3596
rect 4393 3556 4397 3596
rect 4403 3556 4407 3596
rect 4475 3556 4479 3596
rect 4495 3576 4499 3596
rect 4505 3576 4509 3596
rect 4527 3576 4531 3596
rect 4537 3576 4541 3596
rect 4559 3576 4563 3596
rect 4605 3576 4609 3596
rect 4613 3576 4617 3596
rect 4633 3576 4637 3596
rect 4643 3576 4647 3596
rect 4665 3556 4669 3596
rect 4725 3576 4729 3596
rect 4771 3556 4775 3596
rect 4793 3576 4797 3596
rect 4803 3576 4807 3596
rect 4823 3576 4827 3596
rect 4831 3576 4835 3596
rect 4877 3576 4881 3596
rect 4899 3576 4903 3596
rect 4909 3576 4913 3596
rect 4931 3576 4935 3596
rect 4941 3576 4945 3596
rect 4961 3556 4965 3596
rect 5046 3556 5050 3596
rect 5054 3556 5058 3596
rect 5074 3556 5078 3596
rect 5082 3556 5086 3596
rect 5145 3576 5149 3596
rect 5191 3556 5195 3596
rect 5213 3576 5217 3596
rect 5223 3576 5227 3596
rect 5243 3576 5247 3596
rect 5251 3576 5255 3596
rect 5297 3576 5301 3596
rect 5319 3576 5323 3596
rect 5329 3576 5333 3596
rect 5351 3576 5355 3596
rect 5361 3576 5365 3596
rect 5381 3556 5385 3596
rect 5431 3556 5435 3596
rect 5453 3576 5457 3596
rect 5463 3576 5467 3596
rect 5483 3576 5487 3596
rect 5491 3576 5495 3596
rect 5537 3576 5541 3596
rect 5559 3576 5563 3596
rect 5569 3576 5573 3596
rect 5591 3576 5595 3596
rect 5601 3576 5605 3596
rect 5621 3556 5625 3596
rect 5671 3556 5675 3596
rect 5691 3556 5695 3596
rect 5711 3556 5715 3596
rect 5771 3556 5775 3596
rect 5791 3556 5795 3596
rect 5811 3556 5815 3596
rect 5885 3576 5889 3596
rect 5966 3556 5970 3596
rect 5974 3556 5978 3596
rect 5994 3556 5998 3596
rect 6002 3556 6006 3596
rect 6053 3556 6057 3596
rect 6063 3556 6067 3596
rect 6145 3576 6149 3596
rect 6211 3576 6215 3596
rect 6231 3576 6235 3596
rect 6251 3576 6255 3596
rect 6385 3576 6389 3596
rect 6431 3556 6435 3596
rect 6453 3576 6457 3596
rect 6463 3576 6467 3596
rect 6483 3576 6487 3596
rect 6491 3576 6495 3596
rect 6537 3576 6541 3596
rect 6559 3576 6563 3596
rect 6569 3576 6573 3596
rect 6591 3576 6595 3596
rect 6601 3576 6605 3596
rect 6621 3556 6625 3596
rect 43 3144 47 3184
rect 65 3144 69 3164
rect 111 3144 115 3184
rect 133 3144 137 3164
rect 143 3144 147 3164
rect 163 3144 167 3164
rect 171 3144 175 3164
rect 217 3144 221 3164
rect 239 3144 243 3164
rect 249 3144 253 3164
rect 271 3144 275 3164
rect 281 3144 285 3164
rect 301 3144 305 3184
rect 353 3144 357 3184
rect 363 3144 367 3184
rect 452 3144 456 3164
rect 474 3144 478 3184
rect 482 3144 486 3184
rect 553 3144 557 3184
rect 563 3144 567 3184
rect 611 3144 615 3164
rect 672 3144 676 3204
rect 680 3144 684 3204
rect 688 3144 692 3204
rect 773 3144 777 3184
rect 783 3144 787 3184
rect 865 3144 869 3184
rect 885 3144 889 3184
rect 905 3144 909 3184
rect 951 3144 955 3164
rect 1011 3144 1015 3164
rect 1031 3144 1035 3164
rect 1091 3144 1095 3184
rect 1111 3144 1115 3184
rect 1131 3144 1135 3184
rect 1191 3144 1195 3184
rect 1211 3144 1215 3184
rect 1231 3144 1235 3184
rect 1293 3144 1297 3184
rect 1303 3144 1307 3184
rect 1371 3144 1375 3184
rect 1393 3144 1397 3164
rect 1403 3144 1407 3164
rect 1423 3144 1427 3164
rect 1431 3144 1435 3164
rect 1477 3144 1481 3164
rect 1499 3144 1503 3164
rect 1509 3144 1513 3164
rect 1531 3144 1535 3164
rect 1541 3144 1545 3164
rect 1561 3144 1565 3184
rect 1635 3144 1639 3184
rect 1655 3144 1659 3184
rect 1665 3144 1669 3184
rect 1732 3144 1736 3164
rect 1754 3144 1758 3184
rect 1762 3144 1766 3184
rect 1848 3144 1852 3204
rect 1856 3144 1860 3204
rect 1864 3144 1868 3204
rect 1914 3144 1918 3184
rect 1922 3144 1926 3184
rect 1944 3144 1948 3164
rect 2015 3144 2019 3184
rect 2035 3144 2039 3164
rect 2045 3144 2049 3164
rect 2067 3144 2071 3164
rect 2077 3144 2081 3164
rect 2099 3144 2103 3164
rect 2145 3144 2149 3164
rect 2153 3144 2157 3164
rect 2173 3144 2177 3164
rect 2183 3144 2187 3164
rect 2205 3144 2209 3184
rect 2253 3144 2257 3184
rect 2263 3144 2267 3184
rect 2331 3144 2335 3164
rect 2351 3144 2355 3164
rect 2425 3144 2429 3164
rect 2445 3144 2449 3164
rect 2505 3144 2509 3184
rect 2525 3144 2529 3184
rect 2545 3144 2549 3184
rect 2591 3144 2595 3164
rect 2655 3144 2659 3184
rect 2675 3144 2679 3164
rect 2685 3144 2689 3164
rect 2707 3144 2711 3164
rect 2717 3144 2721 3164
rect 2739 3144 2743 3164
rect 2785 3144 2789 3164
rect 2793 3144 2797 3164
rect 2813 3144 2817 3164
rect 2823 3144 2827 3164
rect 2845 3144 2849 3184
rect 2893 3144 2897 3184
rect 2903 3144 2907 3184
rect 2993 3144 2997 3184
rect 3003 3144 3007 3184
rect 3065 3144 3069 3184
rect 3085 3144 3089 3184
rect 3105 3144 3109 3184
rect 3173 3144 3177 3184
rect 3183 3144 3187 3184
rect 3245 3144 3249 3164
rect 3305 3144 3309 3184
rect 3325 3144 3329 3184
rect 3345 3144 3349 3184
rect 3391 3144 3395 3164
rect 3465 3144 3469 3164
rect 3485 3144 3489 3164
rect 3552 3144 3556 3164
rect 3574 3144 3578 3184
rect 3582 3144 3586 3184
rect 3645 3144 3649 3164
rect 3665 3144 3669 3164
rect 3711 3144 3715 3184
rect 3733 3144 3737 3164
rect 3743 3144 3747 3164
rect 3763 3144 3767 3164
rect 3771 3144 3775 3164
rect 3817 3144 3821 3164
rect 3839 3144 3843 3164
rect 3849 3144 3853 3164
rect 3871 3144 3875 3164
rect 3881 3144 3885 3164
rect 3901 3144 3905 3184
rect 3954 3144 3958 3184
rect 3962 3144 3966 3184
rect 3982 3144 3986 3184
rect 3990 3144 3994 3184
rect 4106 3144 4110 3184
rect 4114 3144 4118 3184
rect 4134 3144 4138 3184
rect 4142 3144 4146 3184
rect 4195 3144 4199 3184
rect 4215 3144 4219 3164
rect 4225 3144 4229 3164
rect 4247 3144 4251 3164
rect 4257 3144 4261 3164
rect 4279 3144 4283 3164
rect 4325 3144 4329 3164
rect 4333 3144 4337 3164
rect 4353 3144 4357 3164
rect 4363 3144 4367 3164
rect 4385 3144 4389 3184
rect 4431 3144 4435 3164
rect 4451 3144 4455 3164
rect 4514 3144 4518 3184
rect 4522 3144 4526 3184
rect 4542 3144 4546 3184
rect 4550 3144 4554 3184
rect 4631 3144 4635 3164
rect 4651 3144 4655 3164
rect 4711 3144 4715 3164
rect 4731 3144 4735 3164
rect 4791 3144 4795 3164
rect 4854 3144 4858 3184
rect 4862 3144 4866 3184
rect 4882 3144 4886 3184
rect 4890 3144 4894 3184
rect 4974 3144 4978 3184
rect 4982 3144 4986 3184
rect 5004 3144 5008 3164
rect 5071 3144 5075 3184
rect 5093 3144 5097 3164
rect 5103 3144 5107 3164
rect 5123 3144 5127 3164
rect 5131 3144 5135 3164
rect 5177 3144 5181 3164
rect 5199 3144 5203 3164
rect 5209 3144 5213 3164
rect 5231 3144 5235 3164
rect 5241 3144 5245 3164
rect 5261 3144 5265 3184
rect 5325 3144 5329 3164
rect 5371 3152 5375 3172
rect 5391 3152 5395 3192
rect 5401 3152 5405 3192
rect 5421 3152 5425 3192
rect 5431 3152 5435 3192
rect 5505 3144 5509 3164
rect 5555 3144 5559 3184
rect 5575 3144 5579 3164
rect 5585 3144 5589 3164
rect 5607 3144 5611 3164
rect 5617 3144 5621 3164
rect 5639 3144 5643 3164
rect 5685 3144 5689 3164
rect 5693 3144 5697 3164
rect 5713 3144 5717 3164
rect 5723 3144 5727 3164
rect 5745 3144 5749 3184
rect 5805 3144 5809 3184
rect 5825 3144 5829 3184
rect 5845 3144 5849 3184
rect 5905 3144 5909 3164
rect 5972 3144 5976 3164
rect 5994 3144 5998 3184
rect 6002 3144 6006 3184
rect 6051 3144 6055 3184
rect 6071 3144 6075 3184
rect 6091 3144 6095 3184
rect 6173 3144 6177 3184
rect 6183 3144 6187 3184
rect 6252 3144 6256 3164
rect 6274 3144 6278 3184
rect 6282 3144 6286 3184
rect 6353 3144 6357 3184
rect 6363 3144 6367 3184
rect 6411 3144 6415 3184
rect 6431 3144 6435 3184
rect 6451 3144 6455 3184
rect 6511 3144 6515 3184
rect 6533 3144 6537 3164
rect 6543 3144 6547 3164
rect 6563 3144 6567 3164
rect 6571 3144 6575 3164
rect 6617 3144 6621 3164
rect 6639 3144 6643 3164
rect 6649 3144 6653 3164
rect 6671 3144 6675 3164
rect 6681 3144 6685 3164
rect 6701 3144 6705 3184
rect 31 3076 35 3116
rect 51 3076 55 3116
rect 71 3076 75 3116
rect 91 3076 95 3116
rect 111 3076 115 3116
rect 131 3076 135 3116
rect 151 3076 155 3116
rect 171 3076 175 3116
rect 243 3076 247 3116
rect 265 3096 269 3116
rect 315 3076 319 3116
rect 335 3096 339 3116
rect 345 3096 349 3116
rect 367 3096 371 3116
rect 377 3096 381 3116
rect 399 3096 403 3116
rect 445 3096 449 3116
rect 453 3096 457 3116
rect 473 3096 477 3116
rect 483 3096 487 3116
rect 505 3076 509 3116
rect 573 3076 577 3116
rect 583 3076 587 3116
rect 633 3076 637 3116
rect 643 3076 647 3116
rect 725 3076 729 3116
rect 745 3076 749 3116
rect 765 3076 769 3116
rect 833 3076 837 3116
rect 843 3076 847 3116
rect 913 3076 917 3116
rect 923 3076 927 3116
rect 974 3076 978 3116
rect 982 3076 986 3116
rect 1004 3096 1008 3116
rect 1071 3076 1075 3116
rect 1093 3096 1097 3116
rect 1103 3096 1107 3116
rect 1123 3096 1127 3116
rect 1131 3096 1135 3116
rect 1177 3096 1181 3116
rect 1199 3096 1203 3116
rect 1209 3096 1213 3116
rect 1231 3096 1235 3116
rect 1241 3096 1245 3116
rect 1261 3076 1265 3116
rect 1333 3076 1337 3116
rect 1343 3076 1347 3116
rect 1391 3076 1395 3116
rect 1413 3096 1417 3116
rect 1423 3096 1427 3116
rect 1443 3096 1447 3116
rect 1451 3096 1455 3116
rect 1497 3096 1501 3116
rect 1519 3096 1523 3116
rect 1529 3096 1533 3116
rect 1551 3096 1555 3116
rect 1561 3096 1565 3116
rect 1581 3076 1585 3116
rect 1645 3096 1649 3116
rect 1705 3076 1709 3116
rect 1725 3076 1729 3116
rect 1745 3076 1749 3116
rect 1805 3096 1809 3116
rect 1825 3096 1829 3116
rect 1895 3076 1899 3116
rect 1915 3076 1919 3116
rect 1925 3076 1929 3116
rect 1971 3076 1975 3116
rect 1991 3076 1995 3116
rect 2011 3076 2015 3116
rect 2092 3096 2096 3116
rect 2114 3076 2118 3116
rect 2122 3076 2126 3116
rect 2173 3076 2177 3116
rect 2183 3076 2187 3116
rect 2265 3096 2269 3116
rect 2311 3076 2315 3116
rect 2321 3076 2325 3116
rect 2341 3076 2345 3116
rect 2415 3076 2419 3116
rect 2435 3096 2439 3116
rect 2445 3096 2449 3116
rect 2467 3096 2471 3116
rect 2477 3096 2481 3116
rect 2499 3096 2503 3116
rect 2545 3096 2549 3116
rect 2553 3096 2557 3116
rect 2573 3096 2577 3116
rect 2583 3096 2587 3116
rect 2605 3076 2609 3116
rect 2651 3096 2655 3116
rect 2711 3096 2715 3116
rect 2731 3096 2735 3116
rect 2805 3096 2809 3116
rect 2865 3076 2869 3116
rect 2885 3076 2889 3116
rect 2905 3076 2909 3116
rect 2951 3076 2955 3116
rect 3048 3056 3052 3116
rect 3056 3056 3060 3116
rect 3064 3056 3068 3116
rect 3133 3076 3137 3116
rect 3143 3076 3147 3116
rect 3205 3076 3209 3116
rect 3225 3076 3229 3116
rect 3245 3076 3249 3116
rect 3293 3076 3297 3116
rect 3303 3076 3307 3116
rect 3373 3076 3377 3116
rect 3383 3076 3387 3116
rect 3451 3076 3455 3116
rect 3471 3076 3475 3116
rect 3491 3076 3495 3116
rect 3551 3076 3555 3116
rect 3561 3076 3565 3116
rect 3581 3076 3585 3116
rect 3686 3076 3690 3116
rect 3694 3076 3698 3116
rect 3714 3076 3718 3116
rect 3722 3076 3726 3116
rect 3785 3076 3789 3116
rect 3805 3076 3809 3116
rect 3855 3076 3859 3116
rect 3875 3096 3879 3116
rect 3885 3096 3889 3116
rect 3907 3096 3911 3116
rect 3917 3096 3921 3116
rect 3939 3096 3943 3116
rect 3985 3096 3989 3116
rect 3993 3096 3997 3116
rect 4013 3096 4017 3116
rect 4023 3096 4027 3116
rect 4045 3076 4049 3116
rect 4091 3076 4095 3116
rect 4111 3076 4115 3116
rect 4131 3076 4135 3116
rect 4228 3056 4232 3116
rect 4236 3056 4240 3116
rect 4244 3056 4248 3116
rect 4295 3076 4299 3116
rect 4315 3096 4319 3116
rect 4325 3096 4329 3116
rect 4347 3096 4351 3116
rect 4357 3096 4361 3116
rect 4379 3096 4383 3116
rect 4425 3096 4429 3116
rect 4433 3096 4437 3116
rect 4453 3096 4457 3116
rect 4463 3096 4467 3116
rect 4485 3076 4489 3116
rect 4545 3076 4549 3116
rect 4565 3076 4569 3116
rect 4585 3076 4589 3116
rect 4605 3076 4609 3116
rect 4665 3096 4669 3116
rect 4725 3068 4729 3108
rect 4735 3068 4739 3108
rect 4755 3068 4759 3108
rect 4765 3068 4769 3108
rect 4785 3088 4789 3108
rect 4834 3076 4838 3116
rect 4842 3076 4846 3116
rect 4862 3076 4866 3116
rect 4870 3076 4874 3116
rect 4965 3096 4969 3116
rect 5014 3076 5018 3116
rect 5022 3076 5026 3116
rect 5042 3076 5046 3116
rect 5050 3076 5054 3116
rect 5131 3096 5135 3116
rect 5191 3096 5195 3116
rect 5211 3096 5215 3116
rect 5275 3076 5279 3116
rect 5295 3096 5299 3116
rect 5305 3096 5309 3116
rect 5327 3096 5331 3116
rect 5337 3096 5341 3116
rect 5359 3096 5363 3116
rect 5405 3096 5409 3116
rect 5413 3096 5417 3116
rect 5433 3096 5437 3116
rect 5443 3096 5447 3116
rect 5465 3076 5469 3116
rect 5525 3096 5529 3116
rect 5545 3096 5549 3116
rect 5591 3076 5595 3116
rect 5611 3076 5615 3116
rect 5631 3076 5635 3116
rect 5728 3056 5732 3116
rect 5736 3056 5740 3116
rect 5744 3056 5748 3116
rect 5805 3076 5809 3116
rect 5825 3076 5829 3116
rect 5845 3076 5849 3116
rect 5865 3076 5869 3116
rect 5911 3096 5915 3116
rect 5971 3088 5975 3108
rect 5991 3068 5995 3108
rect 6001 3068 6005 3108
rect 6021 3068 6025 3108
rect 6031 3068 6035 3108
rect 6112 3096 6116 3116
rect 6134 3076 6138 3116
rect 6142 3076 6146 3116
rect 6205 3096 6209 3116
rect 6225 3096 6229 3116
rect 6271 3096 6275 3116
rect 6366 3076 6370 3116
rect 6374 3076 6378 3116
rect 6394 3076 6398 3116
rect 6402 3076 6406 3116
rect 6465 3096 6469 3116
rect 6511 3096 6515 3116
rect 6571 3076 6575 3116
rect 6591 3076 6595 3116
rect 6611 3076 6615 3116
rect 31 2664 35 2684
rect 105 2664 109 2684
rect 125 2664 129 2684
rect 175 2664 179 2704
rect 195 2664 199 2684
rect 205 2664 209 2684
rect 227 2664 231 2684
rect 237 2664 241 2684
rect 259 2664 263 2684
rect 305 2664 309 2684
rect 313 2664 317 2684
rect 333 2664 337 2684
rect 343 2664 347 2684
rect 365 2664 369 2704
rect 411 2664 415 2684
rect 485 2664 489 2684
rect 505 2664 509 2684
rect 555 2664 559 2704
rect 575 2664 579 2684
rect 585 2664 589 2684
rect 607 2664 611 2684
rect 617 2664 621 2684
rect 639 2664 643 2684
rect 685 2664 689 2684
rect 693 2664 697 2684
rect 713 2664 717 2684
rect 723 2664 727 2684
rect 745 2664 749 2704
rect 803 2664 807 2704
rect 825 2664 829 2684
rect 871 2664 875 2704
rect 891 2664 895 2704
rect 953 2664 957 2704
rect 963 2664 967 2704
rect 1033 2664 1037 2704
rect 1043 2664 1047 2704
rect 1111 2664 1115 2684
rect 1174 2664 1178 2704
rect 1182 2664 1186 2704
rect 1202 2664 1206 2704
rect 1210 2664 1214 2704
rect 1312 2664 1316 2684
rect 1334 2664 1338 2704
rect 1342 2664 1346 2704
rect 1405 2664 1409 2684
rect 1465 2664 1469 2704
rect 1485 2664 1489 2704
rect 1505 2664 1509 2704
rect 1551 2664 1555 2684
rect 1571 2664 1575 2684
rect 1633 2664 1637 2704
rect 1643 2664 1647 2704
rect 1711 2664 1715 2684
rect 1731 2664 1735 2684
rect 1805 2664 1809 2704
rect 1825 2664 1829 2704
rect 1845 2664 1849 2704
rect 1891 2664 1895 2684
rect 1911 2664 1915 2684
rect 1931 2664 1935 2704
rect 1991 2664 1995 2704
rect 2011 2664 2015 2704
rect 2031 2664 2035 2704
rect 2112 2664 2116 2684
rect 2134 2664 2138 2704
rect 2142 2664 2146 2704
rect 2195 2664 2199 2704
rect 2215 2664 2219 2684
rect 2225 2664 2229 2684
rect 2247 2664 2251 2684
rect 2257 2664 2261 2684
rect 2279 2664 2283 2684
rect 2325 2664 2329 2684
rect 2333 2664 2337 2684
rect 2353 2664 2357 2684
rect 2363 2664 2367 2684
rect 2385 2664 2389 2704
rect 2433 2664 2437 2704
rect 2443 2664 2447 2704
rect 2511 2664 2515 2684
rect 2585 2664 2589 2684
rect 2635 2664 2639 2704
rect 2655 2664 2659 2684
rect 2665 2664 2669 2684
rect 2687 2664 2691 2684
rect 2697 2664 2701 2684
rect 2719 2664 2723 2684
rect 2765 2664 2769 2684
rect 2773 2664 2777 2684
rect 2793 2664 2797 2684
rect 2803 2664 2807 2684
rect 2825 2664 2829 2704
rect 2871 2664 2875 2704
rect 2891 2664 2895 2704
rect 2911 2664 2915 2704
rect 2992 2664 2996 2684
rect 3014 2664 3018 2704
rect 3022 2664 3026 2704
rect 3071 2664 3075 2704
rect 3093 2664 3097 2684
rect 3103 2664 3107 2684
rect 3123 2664 3127 2684
rect 3131 2664 3135 2684
rect 3177 2664 3181 2684
rect 3199 2664 3203 2684
rect 3209 2664 3213 2684
rect 3231 2664 3235 2684
rect 3241 2664 3245 2684
rect 3261 2664 3265 2704
rect 3311 2664 3315 2684
rect 3371 2664 3375 2704
rect 3391 2664 3395 2704
rect 3411 2664 3415 2704
rect 3431 2664 3435 2704
rect 3491 2664 3495 2704
rect 3511 2664 3515 2704
rect 3531 2664 3535 2704
rect 3605 2664 3609 2704
rect 3625 2664 3629 2704
rect 3645 2664 3649 2704
rect 3665 2664 3669 2704
rect 3711 2664 3715 2704
rect 3731 2664 3735 2704
rect 3751 2664 3755 2704
rect 3825 2664 3829 2704
rect 3845 2664 3849 2704
rect 3865 2664 3869 2704
rect 3885 2664 3889 2704
rect 3945 2664 3949 2684
rect 3991 2664 3995 2684
rect 4011 2664 4015 2684
rect 4071 2664 4075 2684
rect 4091 2664 4095 2684
rect 4172 2664 4176 2684
rect 4194 2664 4198 2704
rect 4202 2664 4206 2704
rect 4251 2664 4255 2704
rect 4271 2664 4275 2704
rect 4291 2664 4295 2704
rect 4388 2664 4392 2724
rect 4396 2664 4400 2724
rect 4404 2664 4408 2724
rect 4455 2664 4459 2704
rect 4475 2664 4479 2684
rect 4485 2664 4489 2684
rect 4507 2664 4511 2684
rect 4517 2664 4521 2684
rect 4539 2664 4543 2684
rect 4585 2664 4589 2684
rect 4593 2664 4597 2684
rect 4613 2664 4617 2684
rect 4623 2664 4627 2684
rect 4645 2664 4649 2704
rect 4691 2664 4695 2684
rect 4751 2664 4755 2684
rect 4771 2664 4775 2684
rect 4831 2664 4835 2704
rect 4851 2664 4855 2704
rect 4871 2664 4875 2704
rect 4945 2664 4949 2684
rect 4965 2664 4969 2684
rect 5025 2664 5029 2704
rect 5045 2664 5049 2704
rect 5065 2664 5069 2704
rect 5085 2664 5089 2704
rect 5134 2664 5138 2704
rect 5142 2664 5146 2704
rect 5164 2664 5168 2684
rect 5231 2664 5235 2684
rect 5253 2664 5257 2704
rect 5311 2664 5315 2704
rect 5331 2664 5335 2704
rect 5351 2664 5355 2704
rect 5425 2664 5429 2704
rect 5445 2664 5449 2704
rect 5465 2664 5469 2704
rect 5485 2664 5489 2704
rect 5545 2664 5549 2684
rect 5595 2664 5599 2704
rect 5615 2664 5619 2684
rect 5625 2664 5629 2684
rect 5647 2664 5651 2684
rect 5657 2664 5661 2684
rect 5679 2664 5683 2684
rect 5725 2664 5729 2684
rect 5733 2664 5737 2684
rect 5753 2664 5757 2684
rect 5763 2664 5767 2684
rect 5785 2664 5789 2704
rect 5831 2672 5835 2692
rect 5851 2672 5855 2712
rect 5861 2672 5865 2712
rect 5881 2672 5885 2712
rect 5891 2672 5895 2712
rect 5951 2672 5955 2692
rect 5971 2672 5975 2712
rect 5981 2672 5985 2712
rect 6001 2672 6005 2712
rect 6011 2672 6015 2712
rect 6071 2672 6075 2692
rect 6091 2672 6095 2712
rect 6101 2672 6105 2712
rect 6121 2672 6125 2712
rect 6131 2672 6135 2712
rect 6215 2664 6219 2704
rect 6235 2664 6239 2704
rect 6245 2664 6249 2704
rect 6305 2664 6309 2704
rect 6325 2664 6329 2704
rect 6371 2664 6375 2704
rect 6381 2664 6385 2704
rect 6401 2664 6405 2704
rect 6471 2664 6475 2704
rect 6493 2664 6497 2684
rect 6503 2664 6507 2684
rect 6523 2664 6527 2684
rect 6531 2664 6535 2684
rect 6577 2664 6581 2684
rect 6599 2664 6603 2684
rect 6609 2664 6613 2684
rect 6631 2664 6635 2684
rect 6641 2664 6645 2684
rect 6661 2664 6665 2704
rect 31 2596 35 2636
rect 53 2616 57 2636
rect 63 2616 67 2636
rect 83 2616 87 2636
rect 91 2616 95 2636
rect 137 2616 141 2636
rect 159 2616 163 2636
rect 169 2616 173 2636
rect 191 2616 195 2636
rect 201 2616 205 2636
rect 221 2596 225 2636
rect 283 2596 287 2636
rect 305 2616 309 2636
rect 351 2596 355 2636
rect 373 2616 377 2636
rect 383 2616 387 2636
rect 403 2616 407 2636
rect 411 2616 415 2636
rect 457 2616 461 2636
rect 479 2616 483 2636
rect 489 2616 493 2636
rect 511 2616 515 2636
rect 521 2616 525 2636
rect 541 2596 545 2636
rect 612 2616 616 2636
rect 634 2596 638 2636
rect 642 2596 646 2636
rect 693 2596 697 2636
rect 703 2596 707 2636
rect 793 2596 797 2636
rect 803 2596 807 2636
rect 865 2596 869 2636
rect 885 2596 889 2636
rect 905 2596 909 2636
rect 925 2596 929 2636
rect 945 2596 949 2636
rect 965 2596 969 2636
rect 985 2596 989 2636
rect 1005 2596 1009 2636
rect 1051 2596 1055 2636
rect 1073 2616 1077 2636
rect 1083 2616 1087 2636
rect 1103 2616 1107 2636
rect 1111 2616 1115 2636
rect 1157 2616 1161 2636
rect 1179 2616 1183 2636
rect 1189 2616 1193 2636
rect 1211 2616 1215 2636
rect 1221 2616 1225 2636
rect 1241 2596 1245 2636
rect 1313 2596 1317 2636
rect 1323 2596 1327 2636
rect 1371 2616 1375 2636
rect 1391 2616 1395 2636
rect 1451 2616 1455 2636
rect 1525 2596 1529 2636
rect 1545 2596 1549 2636
rect 1565 2596 1569 2636
rect 1615 2596 1619 2636
rect 1635 2616 1639 2636
rect 1645 2616 1649 2636
rect 1667 2616 1671 2636
rect 1677 2616 1681 2636
rect 1699 2616 1703 2636
rect 1745 2616 1749 2636
rect 1753 2616 1757 2636
rect 1773 2616 1777 2636
rect 1783 2616 1787 2636
rect 1805 2596 1809 2636
rect 1851 2616 1855 2636
rect 1911 2616 1915 2636
rect 1971 2596 1975 2636
rect 1991 2596 1995 2636
rect 2011 2596 2015 2636
rect 2031 2596 2035 2636
rect 2091 2616 2095 2636
rect 2111 2616 2115 2636
rect 2171 2608 2175 2628
rect 2191 2588 2195 2628
rect 2201 2588 2205 2628
rect 2221 2588 2225 2628
rect 2231 2588 2235 2628
rect 2291 2608 2295 2628
rect 2311 2588 2315 2628
rect 2321 2588 2325 2628
rect 2341 2588 2345 2628
rect 2351 2588 2355 2628
rect 2415 2596 2419 2636
rect 2435 2616 2439 2636
rect 2445 2616 2449 2636
rect 2467 2616 2471 2636
rect 2477 2616 2481 2636
rect 2499 2616 2503 2636
rect 2545 2616 2549 2636
rect 2553 2616 2557 2636
rect 2573 2616 2577 2636
rect 2583 2616 2587 2636
rect 2605 2596 2609 2636
rect 2651 2608 2655 2628
rect 2671 2588 2675 2628
rect 2681 2588 2685 2628
rect 2701 2588 2705 2628
rect 2711 2588 2715 2628
rect 2785 2616 2789 2636
rect 2805 2616 2809 2636
rect 2865 2588 2869 2628
rect 2875 2588 2879 2628
rect 2895 2588 2899 2628
rect 2905 2588 2909 2628
rect 2925 2608 2929 2628
rect 2985 2596 2989 2636
rect 3005 2596 3009 2636
rect 3025 2596 3029 2636
rect 3045 2596 3049 2636
rect 3105 2616 3109 2636
rect 3155 2596 3159 2636
rect 3175 2616 3179 2636
rect 3185 2616 3189 2636
rect 3207 2616 3211 2636
rect 3217 2616 3221 2636
rect 3239 2616 3243 2636
rect 3285 2616 3289 2636
rect 3293 2616 3297 2636
rect 3313 2616 3317 2636
rect 3323 2616 3327 2636
rect 3345 2596 3349 2636
rect 3391 2616 3395 2636
rect 3411 2616 3415 2636
rect 3493 2596 3497 2636
rect 3503 2596 3507 2636
rect 3551 2616 3555 2636
rect 3612 2576 3616 2636
rect 3620 2576 3624 2636
rect 3628 2576 3632 2636
rect 3712 2576 3716 2636
rect 3720 2576 3724 2636
rect 3728 2576 3732 2636
rect 3848 2576 3852 2636
rect 3856 2576 3860 2636
rect 3864 2576 3868 2636
rect 3911 2596 3915 2636
rect 3931 2596 3935 2636
rect 3951 2596 3955 2636
rect 4014 2596 4018 2636
rect 4022 2596 4026 2636
rect 4044 2616 4048 2636
rect 4125 2616 4129 2636
rect 4145 2616 4149 2636
rect 4205 2596 4209 2636
rect 4225 2596 4229 2636
rect 4245 2596 4249 2636
rect 4265 2596 4269 2636
rect 4315 2596 4319 2636
rect 4335 2616 4339 2636
rect 4345 2616 4349 2636
rect 4367 2616 4371 2636
rect 4377 2616 4381 2636
rect 4399 2616 4403 2636
rect 4445 2616 4449 2636
rect 4453 2616 4457 2636
rect 4473 2616 4477 2636
rect 4483 2616 4487 2636
rect 4505 2596 4509 2636
rect 4565 2616 4569 2636
rect 4625 2596 4629 2636
rect 4645 2596 4649 2636
rect 4665 2596 4669 2636
rect 4685 2596 4689 2636
rect 4731 2608 4735 2628
rect 4751 2588 4755 2628
rect 4761 2588 4765 2628
rect 4781 2588 4785 2628
rect 4791 2588 4795 2628
rect 4851 2596 4855 2636
rect 4873 2616 4877 2636
rect 4883 2616 4887 2636
rect 4903 2616 4907 2636
rect 4911 2616 4915 2636
rect 4957 2616 4961 2636
rect 4979 2616 4983 2636
rect 4989 2616 4993 2636
rect 5011 2616 5015 2636
rect 5021 2616 5025 2636
rect 5041 2596 5045 2636
rect 5091 2616 5095 2636
rect 5151 2596 5155 2636
rect 5171 2596 5175 2636
rect 5191 2596 5195 2636
rect 5211 2596 5215 2636
rect 5271 2596 5275 2636
rect 5291 2596 5295 2636
rect 5311 2596 5315 2636
rect 5371 2616 5375 2636
rect 5391 2616 5395 2636
rect 5465 2616 5469 2636
rect 5485 2616 5489 2636
rect 5531 2596 5535 2636
rect 5551 2596 5555 2636
rect 5571 2596 5575 2636
rect 5591 2596 5595 2636
rect 5611 2596 5615 2636
rect 5631 2596 5635 2636
rect 5651 2596 5655 2636
rect 5671 2596 5675 2636
rect 5745 2616 5749 2636
rect 5765 2616 5769 2636
rect 5811 2596 5815 2636
rect 5831 2596 5835 2636
rect 5851 2596 5855 2636
rect 5925 2596 5929 2636
rect 5945 2596 5949 2636
rect 5965 2596 5969 2636
rect 5985 2596 5989 2636
rect 6045 2616 6049 2636
rect 6091 2596 6095 2636
rect 6113 2616 6117 2636
rect 6123 2616 6127 2636
rect 6143 2616 6147 2636
rect 6151 2616 6155 2636
rect 6197 2616 6201 2636
rect 6219 2616 6223 2636
rect 6229 2616 6233 2636
rect 6251 2616 6255 2636
rect 6261 2616 6265 2636
rect 6281 2596 6285 2636
rect 6366 2596 6370 2636
rect 6374 2596 6378 2636
rect 6394 2596 6398 2636
rect 6402 2596 6406 2636
rect 6451 2596 6455 2636
rect 6471 2596 6475 2636
rect 6531 2616 6535 2636
rect 6594 2596 6598 2636
rect 6602 2596 6606 2636
rect 6622 2596 6626 2636
rect 6630 2596 6634 2636
rect 35 2184 39 2224
rect 55 2184 59 2204
rect 65 2184 69 2204
rect 87 2184 91 2204
rect 97 2184 101 2204
rect 119 2184 123 2204
rect 165 2184 169 2204
rect 173 2184 177 2204
rect 193 2184 197 2204
rect 203 2184 207 2204
rect 225 2184 229 2224
rect 283 2184 287 2224
rect 305 2184 309 2204
rect 365 2184 369 2224
rect 425 2184 429 2204
rect 485 2184 489 2204
rect 505 2184 509 2204
rect 551 2184 555 2224
rect 571 2184 575 2224
rect 591 2184 595 2224
rect 675 2184 679 2224
rect 695 2184 699 2224
rect 705 2184 709 2224
rect 752 2184 756 2244
rect 760 2184 764 2244
rect 768 2184 772 2244
rect 853 2184 857 2224
rect 863 2184 867 2224
rect 931 2184 935 2224
rect 953 2184 957 2204
rect 963 2184 967 2204
rect 983 2184 987 2204
rect 991 2184 995 2204
rect 1037 2184 1041 2204
rect 1059 2184 1063 2204
rect 1069 2184 1073 2204
rect 1091 2184 1095 2204
rect 1101 2184 1105 2204
rect 1121 2184 1125 2224
rect 1171 2184 1175 2204
rect 1235 2184 1239 2224
rect 1255 2184 1259 2204
rect 1265 2184 1269 2204
rect 1287 2184 1291 2204
rect 1297 2184 1301 2204
rect 1319 2184 1323 2204
rect 1365 2184 1369 2204
rect 1373 2184 1377 2204
rect 1393 2184 1397 2204
rect 1403 2184 1407 2204
rect 1425 2184 1429 2224
rect 1485 2184 1489 2204
rect 1531 2184 1535 2224
rect 1551 2184 1555 2224
rect 1571 2184 1575 2224
rect 1591 2184 1595 2224
rect 1651 2184 1655 2224
rect 1671 2184 1675 2224
rect 1691 2184 1695 2224
rect 1765 2184 1769 2204
rect 1785 2184 1789 2204
rect 1845 2184 1849 2204
rect 1865 2184 1869 2204
rect 1925 2184 1929 2224
rect 1945 2184 1949 2224
rect 1965 2184 1969 2224
rect 1985 2184 1989 2224
rect 2045 2184 2049 2204
rect 2095 2184 2099 2224
rect 2115 2184 2119 2204
rect 2125 2184 2129 2204
rect 2147 2184 2151 2204
rect 2157 2184 2161 2204
rect 2179 2184 2183 2204
rect 2225 2184 2229 2204
rect 2233 2184 2237 2204
rect 2253 2184 2257 2204
rect 2263 2184 2267 2204
rect 2285 2184 2289 2224
rect 2345 2184 2349 2204
rect 2365 2184 2369 2204
rect 2411 2184 2415 2224
rect 2431 2184 2435 2224
rect 2451 2184 2455 2224
rect 2548 2184 2552 2244
rect 2556 2184 2560 2244
rect 2564 2184 2568 2244
rect 2632 2184 2636 2204
rect 2654 2184 2658 2224
rect 2662 2184 2666 2224
rect 2711 2184 2715 2224
rect 2731 2184 2735 2224
rect 2751 2184 2755 2224
rect 2825 2184 2829 2204
rect 2845 2184 2849 2204
rect 2891 2184 2895 2224
rect 2913 2184 2917 2204
rect 2923 2184 2927 2204
rect 2943 2184 2947 2204
rect 2951 2184 2955 2204
rect 2997 2184 3001 2204
rect 3019 2184 3023 2204
rect 3029 2184 3033 2204
rect 3051 2184 3055 2204
rect 3061 2184 3065 2204
rect 3081 2184 3085 2224
rect 3131 2184 3135 2224
rect 3151 2184 3155 2224
rect 3171 2184 3175 2224
rect 3245 2184 3249 2224
rect 3265 2184 3269 2224
rect 3285 2184 3289 2224
rect 3305 2184 3309 2224
rect 3365 2184 3369 2204
rect 3385 2184 3389 2204
rect 3445 2184 3449 2204
rect 3505 2184 3509 2204
rect 3525 2184 3529 2204
rect 3575 2184 3579 2224
rect 3595 2184 3599 2204
rect 3605 2184 3609 2204
rect 3627 2184 3631 2204
rect 3637 2184 3641 2204
rect 3659 2184 3663 2204
rect 3705 2184 3709 2204
rect 3713 2184 3717 2204
rect 3733 2184 3737 2204
rect 3743 2184 3747 2204
rect 3765 2184 3769 2224
rect 3813 2184 3817 2224
rect 3823 2184 3827 2224
rect 3892 2184 3896 2244
rect 3900 2184 3904 2244
rect 3908 2184 3912 2244
rect 3991 2192 3995 2212
rect 4011 2192 4015 2232
rect 4021 2192 4025 2232
rect 4041 2192 4045 2232
rect 4051 2192 4055 2232
rect 4111 2192 4115 2212
rect 4131 2192 4135 2232
rect 4141 2192 4145 2232
rect 4161 2192 4165 2232
rect 4171 2192 4175 2232
rect 4231 2192 4235 2212
rect 4251 2192 4255 2232
rect 4261 2192 4265 2232
rect 4281 2192 4285 2232
rect 4291 2192 4295 2232
rect 4351 2184 4355 2204
rect 4373 2184 4377 2224
rect 4445 2184 4449 2204
rect 4465 2184 4469 2204
rect 4511 2192 4515 2212
rect 4531 2192 4535 2232
rect 4541 2192 4545 2232
rect 4561 2192 4565 2232
rect 4571 2192 4575 2232
rect 4645 2192 4649 2232
rect 4655 2192 4659 2232
rect 4675 2192 4679 2232
rect 4685 2192 4689 2232
rect 4705 2192 4709 2212
rect 4751 2192 4755 2212
rect 4771 2192 4775 2232
rect 4781 2192 4785 2232
rect 4801 2192 4805 2232
rect 4811 2192 4815 2232
rect 4871 2184 4875 2204
rect 4891 2184 4895 2204
rect 4951 2192 4955 2212
rect 4971 2192 4975 2232
rect 4981 2192 4985 2232
rect 5001 2192 5005 2232
rect 5011 2192 5015 2232
rect 5092 2184 5096 2204
rect 5114 2184 5118 2224
rect 5122 2184 5126 2224
rect 5171 2184 5175 2204
rect 5231 2184 5235 2224
rect 5251 2184 5255 2224
rect 5271 2184 5275 2224
rect 5291 2184 5295 2224
rect 5365 2192 5369 2232
rect 5375 2192 5379 2232
rect 5395 2192 5399 2232
rect 5405 2192 5409 2232
rect 5425 2192 5429 2212
rect 5471 2192 5475 2212
rect 5491 2192 5495 2232
rect 5501 2192 5505 2232
rect 5521 2192 5525 2232
rect 5531 2192 5535 2232
rect 5591 2192 5595 2212
rect 5611 2192 5615 2232
rect 5621 2192 5625 2232
rect 5641 2192 5645 2232
rect 5651 2192 5655 2232
rect 5748 2184 5752 2244
rect 5756 2184 5760 2244
rect 5764 2184 5768 2244
rect 5848 2184 5852 2244
rect 5856 2184 5860 2244
rect 5864 2184 5868 2244
rect 5925 2184 5929 2204
rect 6006 2184 6010 2224
rect 6014 2184 6018 2224
rect 6034 2184 6038 2224
rect 6042 2184 6046 2224
rect 6105 2192 6109 2232
rect 6115 2192 6119 2232
rect 6135 2192 6139 2232
rect 6145 2192 6149 2232
rect 6165 2192 6169 2212
rect 6225 2192 6229 2232
rect 6235 2192 6239 2232
rect 6255 2192 6259 2232
rect 6265 2192 6269 2232
rect 6285 2192 6289 2212
rect 6331 2184 6335 2204
rect 6391 2184 6395 2224
rect 6411 2184 6415 2224
rect 6431 2184 6435 2224
rect 6493 2184 6497 2224
rect 6503 2184 6507 2224
rect 6574 2184 6578 2224
rect 6582 2184 6586 2224
rect 6604 2184 6608 2204
rect 6671 2184 6675 2204
rect 45 2136 49 2156
rect 65 2136 69 2156
rect 133 2116 137 2156
rect 143 2116 147 2156
rect 228 2096 232 2156
rect 236 2096 240 2156
rect 244 2096 248 2156
rect 328 2096 332 2156
rect 336 2096 340 2156
rect 344 2096 348 2156
rect 413 2116 417 2156
rect 423 2116 427 2156
rect 472 2096 476 2156
rect 480 2096 484 2156
rect 488 2096 492 2156
rect 585 2136 589 2156
rect 605 2136 609 2156
rect 651 2116 655 2156
rect 671 2116 675 2156
rect 691 2116 695 2156
rect 752 2096 756 2156
rect 760 2096 764 2156
rect 768 2096 772 2156
rect 851 2136 855 2156
rect 871 2136 875 2156
rect 953 2116 957 2156
rect 963 2116 967 2156
rect 1011 2128 1015 2148
rect 1031 2108 1035 2148
rect 1041 2108 1045 2148
rect 1061 2108 1065 2148
rect 1071 2108 1075 2148
rect 1135 2116 1139 2156
rect 1155 2136 1159 2156
rect 1165 2136 1169 2156
rect 1187 2136 1191 2156
rect 1197 2136 1201 2156
rect 1219 2136 1223 2156
rect 1265 2136 1269 2156
rect 1273 2136 1277 2156
rect 1293 2136 1297 2156
rect 1303 2136 1307 2156
rect 1325 2116 1329 2156
rect 1371 2136 1375 2156
rect 1431 2116 1435 2156
rect 1451 2116 1455 2156
rect 1471 2116 1475 2156
rect 1491 2116 1495 2156
rect 1565 2116 1569 2156
rect 1585 2116 1589 2156
rect 1605 2116 1609 2156
rect 1665 2116 1669 2156
rect 1685 2116 1689 2156
rect 1705 2116 1709 2156
rect 1765 2136 1769 2156
rect 1785 2136 1789 2156
rect 1845 2116 1849 2156
rect 1865 2116 1869 2156
rect 1885 2116 1889 2156
rect 1945 2108 1949 2148
rect 1955 2108 1959 2148
rect 1975 2108 1979 2148
rect 1985 2108 1989 2148
rect 2005 2128 2009 2148
rect 2065 2108 2069 2148
rect 2075 2108 2079 2148
rect 2095 2108 2099 2148
rect 2105 2108 2109 2148
rect 2125 2128 2129 2148
rect 2175 2116 2179 2156
rect 2195 2136 2199 2156
rect 2205 2136 2209 2156
rect 2227 2136 2231 2156
rect 2237 2136 2241 2156
rect 2259 2136 2263 2156
rect 2305 2136 2309 2156
rect 2313 2136 2317 2156
rect 2333 2136 2337 2156
rect 2343 2136 2347 2156
rect 2365 2116 2369 2156
rect 2425 2116 2429 2156
rect 2445 2116 2449 2156
rect 2465 2116 2469 2156
rect 2511 2136 2515 2156
rect 2531 2136 2535 2156
rect 2628 2096 2632 2156
rect 2636 2096 2640 2156
rect 2644 2096 2648 2156
rect 2691 2128 2695 2148
rect 2711 2108 2715 2148
rect 2721 2108 2725 2148
rect 2741 2108 2745 2148
rect 2751 2108 2755 2148
rect 2825 2108 2829 2148
rect 2835 2108 2839 2148
rect 2855 2108 2859 2148
rect 2865 2108 2869 2148
rect 2885 2128 2889 2148
rect 2931 2136 2935 2156
rect 2991 2116 2995 2156
rect 3011 2116 3015 2156
rect 3031 2116 3035 2156
rect 3051 2116 3055 2156
rect 3132 2136 3136 2156
rect 3154 2116 3158 2156
rect 3162 2116 3166 2156
rect 3211 2136 3215 2156
rect 3271 2116 3275 2156
rect 3291 2116 3295 2156
rect 3311 2116 3315 2156
rect 3331 2116 3335 2156
rect 3391 2136 3395 2156
rect 3411 2136 3415 2156
rect 3475 2116 3479 2156
rect 3495 2136 3499 2156
rect 3505 2136 3509 2156
rect 3527 2136 3531 2156
rect 3537 2136 3541 2156
rect 3559 2136 3563 2156
rect 3605 2136 3609 2156
rect 3613 2136 3617 2156
rect 3633 2136 3637 2156
rect 3643 2136 3647 2156
rect 3665 2116 3669 2156
rect 3725 2136 3729 2156
rect 3745 2136 3749 2156
rect 3805 2116 3809 2156
rect 3825 2116 3829 2156
rect 3845 2116 3849 2156
rect 3865 2116 3869 2156
rect 3925 2136 3929 2156
rect 3971 2116 3975 2156
rect 3991 2116 3995 2156
rect 4011 2116 4015 2156
rect 4073 2116 4077 2156
rect 4083 2116 4087 2156
rect 4165 2136 4169 2156
rect 4185 2136 4189 2156
rect 4235 2116 4239 2156
rect 4255 2136 4259 2156
rect 4265 2136 4269 2156
rect 4287 2136 4291 2156
rect 4297 2136 4301 2156
rect 4319 2136 4323 2156
rect 4365 2136 4369 2156
rect 4373 2136 4377 2156
rect 4393 2136 4397 2156
rect 4403 2136 4407 2156
rect 4425 2116 4429 2156
rect 4471 2136 4475 2156
rect 4531 2116 4535 2156
rect 4551 2116 4555 2156
rect 4571 2116 4575 2156
rect 4591 2116 4595 2156
rect 4651 2136 4655 2156
rect 4671 2136 4675 2156
rect 4745 2116 4749 2156
rect 4765 2116 4769 2156
rect 4785 2116 4789 2156
rect 4845 2136 4849 2156
rect 4865 2136 4869 2156
rect 4911 2116 4915 2156
rect 4931 2116 4935 2156
rect 4951 2116 4955 2156
rect 4971 2116 4975 2156
rect 5053 2116 5057 2156
rect 5063 2116 5067 2156
rect 5125 2136 5129 2156
rect 5145 2136 5149 2156
rect 5191 2136 5195 2156
rect 5211 2136 5215 2156
rect 5231 2116 5235 2156
rect 5305 2116 5309 2156
rect 5325 2116 5329 2156
rect 5345 2116 5349 2156
rect 5365 2116 5369 2156
rect 5411 2116 5415 2156
rect 5431 2116 5435 2156
rect 5451 2116 5455 2156
rect 5471 2116 5475 2156
rect 5545 2136 5549 2156
rect 5565 2136 5569 2156
rect 5625 2116 5629 2156
rect 5645 2116 5649 2156
rect 5665 2116 5669 2156
rect 5685 2116 5689 2156
rect 5745 2136 5749 2156
rect 5793 2116 5797 2156
rect 5803 2116 5807 2156
rect 5871 2116 5875 2156
rect 5893 2136 5897 2156
rect 5903 2136 5907 2156
rect 5923 2136 5927 2156
rect 5931 2136 5935 2156
rect 5977 2136 5981 2156
rect 5999 2136 6003 2156
rect 6009 2136 6013 2156
rect 6031 2136 6035 2156
rect 6041 2136 6045 2156
rect 6061 2116 6065 2156
rect 6115 2116 6119 2156
rect 6135 2136 6139 2156
rect 6145 2136 6149 2156
rect 6167 2136 6171 2156
rect 6177 2136 6181 2156
rect 6199 2136 6203 2156
rect 6245 2136 6249 2156
rect 6253 2136 6257 2156
rect 6273 2136 6277 2156
rect 6283 2136 6287 2156
rect 6305 2116 6309 2156
rect 6351 2128 6355 2148
rect 6371 2108 6375 2148
rect 6381 2108 6385 2148
rect 6401 2108 6405 2148
rect 6411 2108 6415 2148
rect 6474 2116 6478 2156
rect 6482 2116 6486 2156
rect 6504 2136 6508 2156
rect 6571 2116 6575 2156
rect 6591 2116 6595 2156
rect 6611 2116 6615 2156
rect 45 1704 49 1724
rect 91 1704 95 1744
rect 113 1704 117 1724
rect 123 1704 127 1724
rect 143 1704 147 1724
rect 151 1704 155 1724
rect 197 1704 201 1724
rect 219 1704 223 1724
rect 229 1704 233 1724
rect 251 1704 255 1724
rect 261 1704 265 1724
rect 281 1704 285 1744
rect 331 1704 335 1724
rect 351 1704 355 1724
rect 425 1704 429 1724
rect 445 1704 449 1724
rect 505 1704 509 1724
rect 565 1704 569 1744
rect 585 1704 589 1744
rect 605 1704 609 1744
rect 651 1704 655 1744
rect 673 1704 677 1724
rect 683 1704 687 1724
rect 703 1704 707 1724
rect 711 1704 715 1724
rect 757 1704 761 1724
rect 779 1704 783 1724
rect 789 1704 793 1724
rect 811 1704 815 1724
rect 821 1704 825 1724
rect 841 1704 845 1744
rect 928 1704 932 1764
rect 936 1704 940 1764
rect 944 1704 948 1764
rect 991 1704 995 1744
rect 1001 1704 1005 1744
rect 1021 1704 1025 1744
rect 1091 1704 1095 1724
rect 1151 1704 1155 1744
rect 1171 1704 1175 1744
rect 1191 1704 1195 1744
rect 1273 1704 1277 1744
rect 1283 1704 1287 1744
rect 1368 1704 1372 1764
rect 1376 1704 1380 1764
rect 1384 1704 1388 1764
rect 1431 1704 1435 1724
rect 1495 1704 1499 1744
rect 1515 1704 1519 1724
rect 1525 1704 1529 1724
rect 1547 1704 1551 1724
rect 1557 1704 1561 1724
rect 1579 1704 1583 1724
rect 1625 1704 1629 1724
rect 1633 1704 1637 1724
rect 1653 1704 1657 1724
rect 1663 1704 1667 1724
rect 1685 1704 1689 1744
rect 1731 1704 1735 1724
rect 1791 1704 1795 1744
rect 1811 1704 1815 1744
rect 1831 1704 1835 1744
rect 1851 1704 1855 1744
rect 1911 1704 1915 1724
rect 1931 1704 1935 1724
rect 1991 1704 1995 1744
rect 2011 1704 2015 1744
rect 2031 1704 2035 1744
rect 2091 1704 2095 1744
rect 2113 1704 2117 1724
rect 2123 1704 2127 1724
rect 2143 1704 2147 1724
rect 2151 1704 2155 1724
rect 2197 1704 2201 1724
rect 2219 1704 2223 1724
rect 2229 1704 2233 1724
rect 2251 1704 2255 1724
rect 2261 1704 2265 1724
rect 2281 1704 2285 1744
rect 2345 1704 2349 1744
rect 2365 1704 2369 1744
rect 2385 1704 2389 1744
rect 2405 1704 2409 1744
rect 2451 1704 2455 1724
rect 2511 1704 2515 1724
rect 2531 1704 2535 1724
rect 2591 1704 2595 1744
rect 2613 1704 2617 1724
rect 2623 1704 2627 1724
rect 2643 1704 2647 1724
rect 2651 1704 2655 1724
rect 2697 1704 2701 1724
rect 2719 1704 2723 1724
rect 2729 1704 2733 1724
rect 2751 1704 2755 1724
rect 2761 1704 2765 1724
rect 2781 1704 2785 1744
rect 2832 1704 2836 1764
rect 2840 1704 2844 1764
rect 2848 1704 2852 1764
rect 2945 1704 2949 1744
rect 2965 1704 2969 1744
rect 2985 1704 2989 1744
rect 3031 1704 3035 1724
rect 3051 1704 3055 1724
rect 3132 1704 3136 1724
rect 3154 1704 3158 1744
rect 3162 1704 3166 1744
rect 3232 1704 3236 1724
rect 3254 1704 3258 1744
rect 3262 1704 3266 1744
rect 3323 1704 3327 1744
rect 3345 1704 3349 1724
rect 3413 1704 3417 1744
rect 3423 1704 3427 1744
rect 3471 1704 3475 1724
rect 3491 1704 3495 1724
rect 3553 1704 3557 1744
rect 3563 1704 3567 1744
rect 3631 1704 3635 1744
rect 3651 1704 3655 1744
rect 3671 1704 3675 1744
rect 3753 1704 3757 1744
rect 3763 1704 3767 1744
rect 3825 1704 3829 1724
rect 3873 1704 3877 1744
rect 3883 1704 3887 1744
rect 3951 1704 3955 1724
rect 3971 1704 3975 1724
rect 4031 1704 4035 1744
rect 4051 1704 4055 1744
rect 4071 1704 4075 1744
rect 4091 1704 4095 1744
rect 4165 1704 4169 1724
rect 4185 1704 4189 1724
rect 4231 1704 4235 1744
rect 4251 1704 4255 1744
rect 4271 1704 4275 1744
rect 4331 1704 4335 1744
rect 4351 1704 4355 1744
rect 4411 1704 4415 1744
rect 4431 1704 4435 1744
rect 4451 1704 4455 1744
rect 4525 1704 4529 1724
rect 4545 1704 4549 1724
rect 4605 1704 4609 1744
rect 4625 1704 4629 1744
rect 4645 1704 4649 1744
rect 4665 1704 4669 1744
rect 4725 1704 4729 1724
rect 4771 1704 4775 1744
rect 4793 1704 4797 1724
rect 4803 1704 4807 1724
rect 4823 1704 4827 1724
rect 4831 1704 4835 1724
rect 4877 1704 4881 1724
rect 4899 1704 4903 1724
rect 4909 1704 4913 1724
rect 4931 1704 4935 1724
rect 4941 1704 4945 1724
rect 4961 1704 4965 1744
rect 5014 1704 5018 1744
rect 5022 1704 5026 1744
rect 5044 1704 5048 1724
rect 5111 1704 5115 1724
rect 5131 1704 5135 1724
rect 5191 1704 5195 1744
rect 5211 1704 5215 1744
rect 5231 1704 5235 1744
rect 5292 1704 5296 1764
rect 5300 1704 5304 1764
rect 5308 1704 5312 1764
rect 5391 1704 5395 1724
rect 5413 1704 5417 1744
rect 5485 1704 5489 1724
rect 5545 1704 5549 1744
rect 5605 1704 5609 1744
rect 5625 1704 5629 1744
rect 5645 1704 5649 1744
rect 5693 1704 5697 1744
rect 5703 1704 5707 1744
rect 5806 1704 5810 1744
rect 5814 1704 5818 1744
rect 5834 1704 5838 1744
rect 5842 1704 5846 1744
rect 5891 1704 5895 1724
rect 5913 1704 5917 1744
rect 5985 1704 5989 1744
rect 6005 1704 6009 1744
rect 6025 1704 6029 1744
rect 6085 1704 6089 1744
rect 6105 1704 6109 1744
rect 6125 1704 6129 1744
rect 6145 1704 6149 1744
rect 6191 1712 6195 1732
rect 6211 1712 6215 1752
rect 6221 1712 6225 1752
rect 6241 1712 6245 1752
rect 6251 1712 6255 1752
rect 6311 1712 6315 1732
rect 6331 1712 6335 1752
rect 6341 1712 6345 1752
rect 6361 1712 6365 1752
rect 6371 1712 6375 1752
rect 6431 1704 6435 1724
rect 6491 1704 6495 1744
rect 6511 1704 6515 1744
rect 6531 1704 6535 1744
rect 6613 1704 6617 1744
rect 6623 1704 6627 1744
rect 45 1656 49 1676
rect 65 1656 69 1676
rect 125 1636 129 1676
rect 145 1636 149 1676
rect 165 1636 169 1676
rect 185 1636 189 1676
rect 205 1636 209 1676
rect 225 1636 229 1676
rect 245 1636 249 1676
rect 265 1636 269 1676
rect 315 1636 319 1676
rect 335 1656 339 1676
rect 345 1656 349 1676
rect 367 1656 371 1676
rect 377 1656 381 1676
rect 399 1656 403 1676
rect 445 1656 449 1676
rect 453 1656 457 1676
rect 473 1656 477 1676
rect 483 1656 487 1676
rect 505 1636 509 1676
rect 565 1656 569 1676
rect 612 1616 616 1676
rect 620 1616 624 1676
rect 628 1616 632 1676
rect 714 1636 718 1676
rect 722 1636 726 1676
rect 744 1656 748 1676
rect 815 1636 819 1676
rect 835 1656 839 1676
rect 845 1656 849 1676
rect 867 1656 871 1676
rect 877 1656 881 1676
rect 899 1656 903 1676
rect 945 1656 949 1676
rect 953 1656 957 1676
rect 973 1656 977 1676
rect 983 1656 987 1676
rect 1005 1636 1009 1676
rect 1065 1656 1069 1676
rect 1111 1636 1115 1676
rect 1131 1636 1135 1676
rect 1151 1636 1155 1676
rect 1171 1636 1175 1676
rect 1245 1636 1249 1676
rect 1265 1636 1269 1676
rect 1285 1636 1289 1676
rect 1345 1656 1349 1676
rect 1365 1656 1369 1676
rect 1425 1628 1429 1668
rect 1435 1628 1439 1668
rect 1455 1628 1459 1668
rect 1465 1628 1469 1668
rect 1485 1648 1489 1668
rect 1545 1628 1549 1668
rect 1555 1628 1559 1668
rect 1575 1628 1579 1668
rect 1585 1628 1589 1668
rect 1605 1648 1609 1668
rect 1665 1628 1669 1668
rect 1675 1628 1679 1668
rect 1695 1628 1699 1668
rect 1705 1628 1709 1668
rect 1725 1648 1729 1668
rect 1771 1636 1775 1676
rect 1793 1656 1797 1676
rect 1803 1656 1807 1676
rect 1823 1656 1827 1676
rect 1831 1656 1835 1676
rect 1877 1656 1881 1676
rect 1899 1656 1903 1676
rect 1909 1656 1913 1676
rect 1931 1656 1935 1676
rect 1941 1656 1945 1676
rect 1961 1636 1965 1676
rect 2011 1648 2015 1668
rect 2031 1628 2035 1668
rect 2041 1628 2045 1668
rect 2061 1628 2065 1668
rect 2071 1628 2075 1668
rect 2131 1656 2135 1676
rect 2191 1636 2195 1676
rect 2211 1636 2215 1676
rect 2231 1636 2235 1676
rect 2251 1636 2255 1676
rect 2311 1656 2315 1676
rect 2331 1656 2335 1676
rect 2405 1636 2409 1676
rect 2425 1636 2429 1676
rect 2445 1636 2449 1676
rect 2503 1636 2507 1676
rect 2525 1656 2529 1676
rect 2571 1656 2575 1676
rect 2591 1656 2595 1676
rect 2673 1636 2677 1676
rect 2683 1636 2687 1676
rect 2733 1636 2737 1676
rect 2743 1636 2747 1676
rect 2825 1628 2829 1668
rect 2835 1628 2839 1668
rect 2855 1628 2859 1668
rect 2865 1628 2869 1668
rect 2885 1648 2889 1668
rect 2968 1616 2972 1676
rect 2976 1616 2980 1676
rect 2984 1616 2988 1676
rect 3045 1636 3049 1676
rect 3095 1636 3099 1676
rect 3115 1656 3119 1676
rect 3125 1656 3129 1676
rect 3147 1656 3151 1676
rect 3157 1656 3161 1676
rect 3179 1656 3183 1676
rect 3225 1656 3229 1676
rect 3233 1656 3237 1676
rect 3253 1656 3257 1676
rect 3263 1656 3267 1676
rect 3285 1636 3289 1676
rect 3353 1636 3357 1676
rect 3363 1636 3367 1676
rect 3425 1636 3429 1676
rect 3445 1636 3449 1676
rect 3465 1636 3469 1676
rect 3514 1636 3518 1676
rect 3522 1636 3526 1676
rect 3542 1636 3546 1676
rect 3550 1636 3554 1676
rect 3645 1636 3649 1676
rect 3665 1636 3669 1676
rect 3685 1636 3689 1676
rect 3745 1656 3749 1676
rect 3805 1656 3809 1676
rect 3825 1656 3829 1676
rect 3885 1636 3889 1676
rect 3905 1636 3909 1676
rect 3925 1636 3929 1676
rect 3945 1636 3949 1676
rect 4005 1656 4009 1676
rect 4055 1636 4059 1676
rect 4075 1656 4079 1676
rect 4085 1656 4089 1676
rect 4107 1656 4111 1676
rect 4117 1656 4121 1676
rect 4139 1656 4143 1676
rect 4185 1656 4189 1676
rect 4193 1656 4197 1676
rect 4213 1656 4217 1676
rect 4223 1656 4227 1676
rect 4245 1636 4249 1676
rect 4305 1628 4309 1668
rect 4315 1628 4319 1668
rect 4335 1628 4339 1668
rect 4345 1628 4349 1668
rect 4365 1648 4369 1668
rect 4425 1628 4429 1668
rect 4435 1628 4439 1668
rect 4455 1628 4459 1668
rect 4465 1628 4469 1668
rect 4485 1648 4489 1668
rect 4531 1648 4535 1668
rect 4551 1628 4555 1668
rect 4561 1628 4565 1668
rect 4581 1628 4585 1668
rect 4591 1628 4595 1668
rect 4651 1648 4655 1668
rect 4671 1628 4675 1668
rect 4681 1628 4685 1668
rect 4701 1628 4705 1668
rect 4711 1628 4715 1668
rect 4771 1648 4775 1668
rect 4791 1628 4795 1668
rect 4801 1628 4805 1668
rect 4821 1628 4825 1668
rect 4831 1628 4835 1668
rect 4891 1648 4895 1668
rect 4911 1628 4915 1668
rect 4921 1628 4925 1668
rect 4941 1628 4945 1668
rect 4951 1628 4955 1668
rect 5011 1636 5015 1676
rect 5033 1656 5037 1676
rect 5043 1656 5047 1676
rect 5063 1656 5067 1676
rect 5071 1656 5075 1676
rect 5117 1656 5121 1676
rect 5139 1656 5143 1676
rect 5149 1656 5153 1676
rect 5171 1656 5175 1676
rect 5181 1656 5185 1676
rect 5201 1636 5205 1676
rect 5251 1636 5255 1676
rect 5273 1656 5277 1676
rect 5283 1656 5287 1676
rect 5303 1656 5307 1676
rect 5311 1656 5315 1676
rect 5357 1656 5361 1676
rect 5379 1656 5383 1676
rect 5389 1656 5393 1676
rect 5411 1656 5415 1676
rect 5421 1656 5425 1676
rect 5441 1636 5445 1676
rect 5494 1636 5498 1676
rect 5502 1636 5506 1676
rect 5522 1636 5526 1676
rect 5530 1636 5534 1676
rect 5611 1648 5615 1668
rect 5631 1628 5635 1668
rect 5641 1628 5645 1668
rect 5661 1628 5665 1668
rect 5671 1628 5675 1668
rect 5745 1636 5749 1676
rect 5765 1636 5769 1676
rect 5785 1636 5789 1676
rect 5845 1656 5849 1676
rect 5865 1656 5869 1676
rect 5933 1636 5937 1676
rect 5943 1636 5947 1676
rect 6005 1636 6009 1676
rect 6025 1636 6029 1676
rect 6045 1636 6049 1676
rect 6105 1656 6109 1676
rect 6125 1656 6129 1676
rect 6185 1636 6189 1676
rect 6205 1636 6209 1676
rect 6225 1636 6229 1676
rect 6245 1636 6249 1676
rect 6305 1628 6309 1668
rect 6315 1628 6319 1668
rect 6335 1628 6339 1668
rect 6345 1628 6349 1668
rect 6365 1648 6369 1668
rect 6411 1656 6415 1676
rect 6471 1636 6475 1676
rect 6493 1656 6497 1676
rect 6503 1656 6507 1676
rect 6523 1656 6527 1676
rect 6531 1656 6535 1676
rect 6577 1656 6581 1676
rect 6599 1656 6603 1676
rect 6609 1656 6613 1676
rect 6631 1656 6635 1676
rect 6641 1656 6645 1676
rect 6661 1636 6665 1676
rect 31 1224 35 1264
rect 41 1224 45 1264
rect 61 1224 65 1264
rect 131 1224 135 1244
rect 151 1224 155 1244
rect 225 1224 229 1264
rect 245 1224 249 1264
rect 265 1224 269 1264
rect 325 1224 329 1244
rect 345 1224 349 1244
rect 391 1224 395 1244
rect 451 1224 455 1244
rect 533 1224 537 1264
rect 543 1224 547 1264
rect 594 1224 598 1264
rect 602 1224 606 1264
rect 624 1224 628 1244
rect 695 1224 699 1264
rect 715 1224 719 1244
rect 725 1224 729 1244
rect 747 1224 751 1244
rect 757 1224 761 1244
rect 779 1224 783 1244
rect 825 1224 829 1244
rect 833 1224 837 1244
rect 853 1224 857 1244
rect 863 1224 867 1244
rect 885 1224 889 1264
rect 953 1224 957 1264
rect 963 1224 967 1264
rect 1012 1224 1016 1284
rect 1020 1224 1024 1284
rect 1028 1224 1032 1284
rect 1111 1224 1115 1244
rect 1131 1224 1135 1244
rect 1195 1224 1199 1264
rect 1215 1224 1219 1244
rect 1225 1224 1229 1244
rect 1247 1224 1251 1244
rect 1257 1224 1261 1244
rect 1279 1224 1283 1244
rect 1325 1224 1329 1244
rect 1333 1224 1337 1244
rect 1353 1224 1357 1244
rect 1363 1224 1367 1244
rect 1385 1224 1389 1264
rect 1445 1224 1449 1264
rect 1465 1224 1469 1264
rect 1485 1224 1489 1264
rect 1505 1224 1509 1264
rect 1525 1224 1529 1264
rect 1545 1224 1549 1264
rect 1565 1224 1569 1264
rect 1585 1224 1589 1264
rect 1645 1232 1649 1272
rect 1655 1232 1659 1272
rect 1675 1232 1679 1272
rect 1685 1232 1689 1272
rect 1705 1232 1709 1252
rect 1765 1224 1769 1244
rect 1785 1224 1789 1244
rect 1845 1224 1849 1264
rect 1865 1224 1869 1264
rect 1885 1224 1889 1264
rect 1905 1224 1909 1264
rect 1965 1224 1969 1264
rect 1985 1224 1989 1264
rect 2005 1224 2009 1264
rect 2051 1224 2055 1244
rect 2111 1224 2115 1264
rect 2131 1224 2135 1264
rect 2151 1224 2155 1264
rect 2213 1224 2217 1264
rect 2223 1224 2227 1264
rect 2291 1232 2295 1252
rect 2311 1232 2315 1272
rect 2321 1232 2325 1272
rect 2341 1232 2345 1272
rect 2351 1232 2355 1272
rect 2425 1232 2429 1272
rect 2435 1232 2439 1272
rect 2455 1232 2459 1272
rect 2465 1232 2469 1272
rect 2485 1232 2489 1252
rect 2566 1224 2570 1264
rect 2574 1224 2578 1264
rect 2594 1224 2598 1264
rect 2602 1224 2606 1264
rect 2654 1224 2658 1264
rect 2662 1224 2666 1264
rect 2682 1224 2686 1264
rect 2690 1224 2694 1264
rect 2806 1224 2810 1264
rect 2814 1224 2818 1264
rect 2834 1224 2838 1264
rect 2842 1224 2846 1264
rect 2891 1224 2895 1244
rect 2913 1224 2917 1264
rect 3006 1224 3010 1264
rect 3014 1224 3018 1264
rect 3034 1224 3038 1264
rect 3042 1224 3046 1264
rect 3105 1224 3109 1244
rect 3165 1232 3169 1272
rect 3175 1232 3179 1272
rect 3195 1232 3199 1272
rect 3205 1232 3209 1272
rect 3225 1232 3229 1252
rect 3275 1224 3279 1264
rect 3295 1224 3299 1244
rect 3305 1224 3309 1244
rect 3327 1224 3331 1244
rect 3337 1224 3341 1244
rect 3359 1224 3363 1244
rect 3405 1224 3409 1244
rect 3413 1224 3417 1244
rect 3433 1224 3437 1244
rect 3443 1224 3447 1244
rect 3465 1224 3469 1264
rect 3525 1224 3529 1244
rect 3545 1224 3549 1244
rect 3605 1224 3609 1264
rect 3625 1224 3629 1264
rect 3645 1224 3649 1264
rect 3665 1224 3669 1264
rect 3725 1224 3729 1264
rect 3745 1224 3749 1264
rect 3765 1224 3769 1264
rect 3825 1224 3829 1244
rect 3871 1224 3875 1264
rect 3893 1224 3897 1244
rect 3903 1224 3907 1244
rect 3923 1224 3927 1244
rect 3931 1224 3935 1244
rect 3977 1224 3981 1244
rect 3999 1224 4003 1244
rect 4009 1224 4013 1244
rect 4031 1224 4035 1244
rect 4041 1224 4045 1244
rect 4061 1224 4065 1264
rect 4111 1224 4115 1264
rect 4133 1224 4137 1244
rect 4143 1224 4147 1244
rect 4163 1224 4167 1244
rect 4171 1224 4175 1244
rect 4217 1224 4221 1244
rect 4239 1224 4243 1244
rect 4249 1224 4253 1244
rect 4271 1224 4275 1244
rect 4281 1224 4285 1244
rect 4301 1224 4305 1264
rect 4365 1224 4369 1244
rect 4414 1224 4418 1264
rect 4422 1224 4426 1264
rect 4442 1224 4446 1264
rect 4450 1224 4454 1264
rect 4531 1232 4535 1252
rect 4551 1232 4555 1272
rect 4561 1232 4565 1272
rect 4581 1232 4585 1272
rect 4591 1232 4595 1272
rect 4686 1224 4690 1264
rect 4694 1224 4698 1264
rect 4714 1224 4718 1264
rect 4722 1224 4726 1264
rect 4783 1224 4787 1264
rect 4805 1224 4809 1244
rect 4873 1224 4877 1264
rect 4883 1224 4887 1264
rect 4953 1224 4957 1264
rect 4963 1224 4967 1264
rect 5025 1224 5029 1264
rect 5045 1224 5049 1264
rect 5065 1224 5069 1264
rect 5085 1224 5089 1264
rect 5145 1224 5149 1264
rect 5165 1224 5169 1264
rect 5185 1224 5189 1264
rect 5205 1224 5209 1264
rect 5251 1224 5255 1264
rect 5333 1224 5337 1264
rect 5343 1224 5347 1264
rect 5391 1224 5395 1264
rect 5411 1224 5415 1264
rect 5431 1224 5435 1264
rect 5451 1224 5455 1264
rect 5532 1224 5536 1244
rect 5554 1224 5558 1264
rect 5562 1224 5566 1264
rect 5611 1224 5615 1264
rect 5671 1232 5675 1252
rect 5691 1232 5695 1272
rect 5701 1232 5705 1272
rect 5721 1232 5725 1272
rect 5731 1232 5735 1272
rect 5813 1224 5817 1264
rect 5823 1224 5827 1264
rect 5885 1224 5889 1264
rect 5905 1224 5909 1264
rect 5925 1224 5929 1264
rect 5985 1224 5989 1244
rect 6031 1224 6035 1264
rect 6051 1224 6055 1264
rect 6071 1224 6075 1264
rect 6131 1224 6135 1264
rect 6151 1224 6155 1264
rect 6171 1224 6175 1264
rect 6191 1224 6195 1264
rect 6251 1224 6255 1264
rect 6273 1224 6277 1244
rect 6283 1224 6287 1244
rect 6303 1224 6307 1244
rect 6311 1224 6315 1244
rect 6357 1224 6361 1244
rect 6379 1224 6383 1244
rect 6389 1224 6393 1244
rect 6411 1224 6415 1244
rect 6421 1224 6425 1244
rect 6441 1224 6445 1264
rect 6491 1224 6495 1264
rect 6513 1224 6517 1244
rect 6523 1224 6527 1244
rect 6543 1224 6547 1244
rect 6551 1224 6555 1244
rect 6597 1224 6601 1244
rect 6619 1224 6623 1244
rect 6629 1224 6633 1244
rect 6651 1224 6655 1244
rect 6661 1224 6665 1244
rect 6681 1224 6685 1264
rect 31 1156 35 1196
rect 53 1176 57 1196
rect 63 1176 67 1196
rect 83 1176 87 1196
rect 91 1176 95 1196
rect 137 1176 141 1196
rect 159 1176 163 1196
rect 169 1176 173 1196
rect 191 1176 195 1196
rect 201 1176 205 1196
rect 221 1156 225 1196
rect 285 1176 289 1196
rect 331 1156 335 1196
rect 353 1176 357 1196
rect 363 1176 367 1196
rect 383 1176 387 1196
rect 391 1176 395 1196
rect 437 1176 441 1196
rect 459 1176 463 1196
rect 469 1176 473 1196
rect 491 1176 495 1196
rect 501 1176 505 1196
rect 521 1156 525 1196
rect 571 1176 575 1196
rect 632 1136 636 1196
rect 640 1136 644 1196
rect 648 1136 652 1196
rect 731 1176 735 1196
rect 751 1176 755 1196
rect 812 1136 816 1196
rect 820 1136 824 1196
rect 828 1136 832 1196
rect 913 1156 917 1196
rect 923 1156 927 1196
rect 991 1176 995 1196
rect 1055 1156 1059 1196
rect 1075 1176 1079 1196
rect 1085 1176 1089 1196
rect 1107 1176 1111 1196
rect 1117 1176 1121 1196
rect 1139 1176 1143 1196
rect 1185 1176 1189 1196
rect 1193 1176 1197 1196
rect 1213 1176 1217 1196
rect 1223 1176 1227 1196
rect 1245 1156 1249 1196
rect 1291 1156 1295 1196
rect 1311 1156 1315 1196
rect 1331 1156 1335 1196
rect 1351 1156 1355 1196
rect 1371 1156 1375 1196
rect 1391 1156 1395 1196
rect 1411 1156 1415 1196
rect 1431 1156 1435 1196
rect 1495 1156 1499 1196
rect 1515 1176 1519 1196
rect 1525 1176 1529 1196
rect 1547 1176 1551 1196
rect 1557 1176 1561 1196
rect 1579 1176 1583 1196
rect 1625 1176 1629 1196
rect 1633 1176 1637 1196
rect 1653 1176 1657 1196
rect 1663 1176 1667 1196
rect 1685 1156 1689 1196
rect 1745 1176 1749 1196
rect 1765 1176 1769 1196
rect 1825 1156 1829 1196
rect 1845 1156 1849 1196
rect 1865 1156 1869 1196
rect 1885 1156 1889 1196
rect 1945 1156 1949 1196
rect 1965 1156 1969 1196
rect 1985 1156 1989 1196
rect 2045 1156 2049 1196
rect 2065 1156 2069 1196
rect 2085 1156 2089 1196
rect 2145 1176 2149 1196
rect 2165 1176 2169 1196
rect 2225 1156 2229 1196
rect 2245 1156 2249 1196
rect 2265 1156 2269 1196
rect 2285 1156 2289 1196
rect 2335 1156 2339 1196
rect 2355 1176 2359 1196
rect 2365 1176 2369 1196
rect 2387 1176 2391 1196
rect 2397 1176 2401 1196
rect 2419 1176 2423 1196
rect 2465 1176 2469 1196
rect 2473 1176 2477 1196
rect 2493 1176 2497 1196
rect 2503 1176 2507 1196
rect 2525 1156 2529 1196
rect 2585 1176 2589 1196
rect 2631 1156 2635 1196
rect 2651 1156 2655 1196
rect 2671 1156 2675 1196
rect 2743 1156 2747 1196
rect 2765 1176 2769 1196
rect 2811 1176 2815 1196
rect 2906 1156 2910 1196
rect 2914 1156 2918 1196
rect 2934 1156 2938 1196
rect 2942 1156 2946 1196
rect 2995 1156 2999 1196
rect 3015 1176 3019 1196
rect 3025 1176 3029 1196
rect 3047 1176 3051 1196
rect 3057 1176 3061 1196
rect 3079 1176 3083 1196
rect 3125 1176 3129 1196
rect 3133 1176 3137 1196
rect 3153 1176 3157 1196
rect 3163 1176 3167 1196
rect 3185 1156 3189 1196
rect 3233 1156 3237 1196
rect 3243 1156 3247 1196
rect 3325 1148 3329 1188
rect 3335 1148 3339 1188
rect 3355 1148 3359 1188
rect 3365 1148 3369 1188
rect 3385 1168 3389 1188
rect 3431 1168 3435 1188
rect 3451 1148 3455 1188
rect 3461 1148 3465 1188
rect 3481 1148 3485 1188
rect 3491 1148 3495 1188
rect 3563 1156 3567 1196
rect 3585 1176 3589 1196
rect 3635 1156 3639 1196
rect 3655 1176 3659 1196
rect 3665 1176 3669 1196
rect 3687 1176 3691 1196
rect 3697 1176 3701 1196
rect 3719 1176 3723 1196
rect 3765 1176 3769 1196
rect 3773 1176 3777 1196
rect 3793 1176 3797 1196
rect 3803 1176 3807 1196
rect 3825 1156 3829 1196
rect 3871 1168 3875 1188
rect 3891 1148 3895 1188
rect 3901 1148 3905 1188
rect 3921 1148 3925 1188
rect 3931 1148 3935 1188
rect 4005 1148 4009 1188
rect 4015 1148 4019 1188
rect 4035 1148 4039 1188
rect 4045 1148 4049 1188
rect 4065 1168 4069 1188
rect 4111 1176 4115 1196
rect 4171 1156 4175 1196
rect 4191 1156 4195 1196
rect 4211 1156 4215 1196
rect 4231 1156 4235 1196
rect 4291 1176 4295 1196
rect 4311 1176 4315 1196
rect 4385 1156 4389 1196
rect 4405 1156 4409 1196
rect 4425 1156 4429 1196
rect 4492 1176 4496 1196
rect 4514 1156 4518 1196
rect 4522 1156 4526 1196
rect 4575 1156 4579 1196
rect 4595 1176 4599 1196
rect 4605 1176 4609 1196
rect 4627 1176 4631 1196
rect 4637 1176 4641 1196
rect 4659 1176 4663 1196
rect 4705 1176 4709 1196
rect 4713 1176 4717 1196
rect 4733 1176 4737 1196
rect 4743 1176 4747 1196
rect 4765 1156 4769 1196
rect 4811 1156 4815 1196
rect 4831 1156 4835 1196
rect 4851 1156 4855 1196
rect 4871 1156 4875 1196
rect 4945 1176 4949 1196
rect 4965 1176 4969 1196
rect 5025 1156 5029 1196
rect 5045 1156 5049 1196
rect 5065 1156 5069 1196
rect 5125 1176 5129 1196
rect 5145 1176 5149 1196
rect 5191 1176 5195 1196
rect 5211 1176 5215 1196
rect 5271 1176 5275 1196
rect 5291 1176 5295 1196
rect 5363 1156 5367 1196
rect 5385 1176 5389 1196
rect 5431 1176 5435 1196
rect 5451 1176 5455 1196
rect 5511 1176 5515 1196
rect 5531 1176 5535 1196
rect 5594 1156 5598 1196
rect 5602 1156 5606 1196
rect 5624 1176 5628 1196
rect 5691 1176 5695 1196
rect 5711 1176 5715 1196
rect 5731 1156 5735 1196
rect 5805 1176 5809 1196
rect 5825 1176 5829 1196
rect 5871 1156 5875 1196
rect 5891 1156 5895 1196
rect 5911 1156 5915 1196
rect 6008 1136 6012 1196
rect 6016 1136 6020 1196
rect 6024 1136 6028 1196
rect 6071 1156 6075 1196
rect 6091 1156 6095 1196
rect 6111 1156 6115 1196
rect 6185 1176 6189 1196
rect 6205 1176 6209 1196
rect 6251 1176 6255 1196
rect 6271 1176 6275 1196
rect 6331 1156 6335 1196
rect 6353 1176 6357 1196
rect 6363 1176 6367 1196
rect 6383 1176 6387 1196
rect 6391 1176 6395 1196
rect 6437 1176 6441 1196
rect 6459 1176 6463 1196
rect 6469 1176 6473 1196
rect 6491 1176 6495 1196
rect 6501 1176 6505 1196
rect 6521 1156 6525 1196
rect 6571 1156 6575 1196
rect 6591 1156 6595 1196
rect 6611 1156 6615 1196
rect 6631 1156 6635 1196
rect 31 744 35 764
rect 51 744 55 764
rect 71 744 75 784
rect 153 744 157 784
rect 163 744 167 784
rect 211 744 215 784
rect 233 744 237 764
rect 243 744 247 764
rect 263 744 267 764
rect 271 744 275 764
rect 317 744 321 764
rect 339 744 343 764
rect 349 744 353 764
rect 371 744 375 764
rect 381 744 385 764
rect 401 744 405 784
rect 465 744 469 764
rect 525 744 529 764
rect 545 744 549 764
rect 591 744 595 764
rect 611 744 615 764
rect 673 744 677 784
rect 683 744 687 784
rect 752 744 756 804
rect 760 744 764 804
rect 768 744 772 804
rect 851 744 855 784
rect 871 744 875 784
rect 891 744 895 784
rect 911 744 915 784
rect 971 744 975 784
rect 991 744 995 784
rect 1011 744 1015 784
rect 1071 744 1075 784
rect 1091 744 1095 784
rect 1111 744 1115 784
rect 1245 744 1249 764
rect 1265 744 1269 764
rect 1285 744 1289 764
rect 1351 744 1355 784
rect 1371 744 1375 784
rect 1391 744 1395 784
rect 1465 744 1469 764
rect 1515 744 1519 784
rect 1535 744 1539 764
rect 1545 744 1549 764
rect 1567 744 1571 764
rect 1577 744 1581 764
rect 1599 744 1603 764
rect 1645 744 1649 764
rect 1653 744 1657 764
rect 1673 744 1677 764
rect 1683 744 1687 764
rect 1705 744 1709 784
rect 1751 744 1755 764
rect 1811 752 1815 772
rect 1831 752 1835 792
rect 1841 752 1845 792
rect 1861 752 1865 792
rect 1871 752 1875 792
rect 1931 744 1935 784
rect 1951 744 1955 784
rect 1971 744 1975 784
rect 2033 744 2037 784
rect 2043 744 2047 784
rect 2111 744 2115 784
rect 2133 744 2137 764
rect 2143 744 2147 764
rect 2163 744 2167 764
rect 2171 744 2175 764
rect 2217 744 2221 764
rect 2239 744 2243 764
rect 2249 744 2253 764
rect 2271 744 2275 764
rect 2281 744 2285 764
rect 2301 744 2305 784
rect 2351 744 2355 764
rect 2411 744 2415 784
rect 2431 744 2435 784
rect 2451 744 2455 784
rect 2471 744 2475 784
rect 2531 744 2535 764
rect 2551 744 2555 764
rect 2625 744 2629 784
rect 2645 744 2649 784
rect 2665 744 2669 784
rect 2725 744 2729 784
rect 2745 744 2749 784
rect 2765 744 2769 784
rect 2785 744 2789 784
rect 2805 744 2809 784
rect 2825 744 2829 784
rect 2845 744 2849 784
rect 2865 744 2869 784
rect 2914 744 2918 784
rect 2922 744 2926 784
rect 2944 744 2948 764
rect 3032 744 3036 764
rect 3054 744 3058 784
rect 3062 744 3066 784
rect 3125 752 3129 792
rect 3135 752 3139 792
rect 3155 752 3159 792
rect 3165 752 3169 792
rect 3185 752 3189 772
rect 3245 752 3249 792
rect 3255 752 3259 792
rect 3275 752 3279 792
rect 3285 752 3289 792
rect 3305 752 3309 772
rect 3365 744 3369 784
rect 3385 744 3389 784
rect 3405 744 3409 784
rect 3453 744 3457 784
rect 3463 744 3467 784
rect 3531 752 3535 772
rect 3551 752 3555 792
rect 3561 752 3565 792
rect 3581 752 3585 792
rect 3591 752 3595 792
rect 3665 744 3669 764
rect 3725 752 3729 792
rect 3735 752 3739 792
rect 3755 752 3759 792
rect 3765 752 3769 792
rect 3785 752 3789 772
rect 3835 744 3839 784
rect 3855 744 3859 764
rect 3865 744 3869 764
rect 3887 744 3891 764
rect 3897 744 3901 764
rect 3919 744 3923 764
rect 3965 744 3969 764
rect 3973 744 3977 764
rect 3993 744 3997 764
rect 4003 744 4007 764
rect 4025 744 4029 784
rect 4071 752 4075 772
rect 4091 752 4095 792
rect 4101 752 4105 792
rect 4121 752 4125 792
rect 4131 752 4135 792
rect 4194 744 4198 784
rect 4202 744 4206 784
rect 4224 744 4228 764
rect 4291 744 4295 784
rect 4311 744 4315 784
rect 4331 744 4335 784
rect 4428 744 4432 804
rect 4436 744 4440 804
rect 4444 744 4448 804
rect 4491 744 4495 764
rect 4551 744 4555 784
rect 4571 744 4575 784
rect 4591 744 4595 784
rect 4653 744 4657 784
rect 4663 744 4667 784
rect 4745 744 4749 764
rect 4791 744 4795 784
rect 4811 744 4815 784
rect 4831 744 4835 784
rect 4893 744 4897 784
rect 4903 744 4907 784
rect 4971 752 4975 772
rect 4991 752 4995 792
rect 5001 752 5005 792
rect 5021 752 5025 792
rect 5031 752 5035 792
rect 5105 752 5109 792
rect 5115 752 5119 792
rect 5135 752 5139 792
rect 5145 752 5149 792
rect 5165 752 5169 772
rect 5211 744 5215 784
rect 5231 744 5235 784
rect 5251 744 5255 784
rect 5271 744 5275 784
rect 5291 744 5295 784
rect 5311 744 5315 784
rect 5331 744 5335 784
rect 5351 744 5355 784
rect 5414 744 5418 784
rect 5422 744 5426 784
rect 5444 744 5448 764
rect 5525 744 5529 764
rect 5571 744 5575 784
rect 5591 744 5595 784
rect 5611 744 5615 784
rect 5673 744 5677 784
rect 5683 744 5687 784
rect 5751 744 5755 784
rect 5771 744 5775 784
rect 5791 744 5795 784
rect 5888 744 5892 804
rect 5896 744 5900 804
rect 5904 744 5908 804
rect 5955 744 5959 784
rect 5975 744 5979 764
rect 5985 744 5989 764
rect 6007 744 6011 764
rect 6017 744 6021 764
rect 6039 744 6043 764
rect 6085 744 6089 764
rect 6093 744 6097 764
rect 6113 744 6117 764
rect 6123 744 6127 764
rect 6145 744 6149 784
rect 6191 744 6195 784
rect 6211 744 6215 784
rect 6231 744 6235 784
rect 6291 744 6295 784
rect 6311 744 6315 784
rect 6331 744 6335 784
rect 6413 744 6417 784
rect 6423 744 6427 784
rect 6475 744 6479 784
rect 6495 744 6499 764
rect 6505 744 6509 764
rect 6527 744 6531 764
rect 6537 744 6541 764
rect 6559 744 6563 764
rect 6605 744 6609 764
rect 6613 744 6617 764
rect 6633 744 6637 764
rect 6643 744 6647 764
rect 6665 744 6669 784
rect 31 696 35 716
rect 93 676 97 716
rect 103 676 107 716
rect 174 676 178 716
rect 182 676 186 716
rect 204 696 208 716
rect 271 696 275 716
rect 352 696 356 716
rect 374 676 378 716
rect 382 676 386 716
rect 432 656 436 716
rect 440 656 444 716
rect 448 656 452 716
rect 553 676 557 716
rect 563 676 567 716
rect 648 656 652 716
rect 656 656 660 716
rect 664 656 668 716
rect 711 696 715 716
rect 771 696 775 716
rect 845 696 849 716
rect 865 696 869 716
rect 985 696 989 716
rect 1005 696 1009 716
rect 1025 696 1029 716
rect 1095 676 1099 716
rect 1115 696 1119 716
rect 1125 696 1129 716
rect 1147 696 1151 716
rect 1157 696 1161 716
rect 1179 696 1183 716
rect 1225 696 1229 716
rect 1233 696 1237 716
rect 1253 696 1257 716
rect 1263 696 1267 716
rect 1285 676 1289 716
rect 1331 696 1335 716
rect 1353 676 1357 716
rect 1413 676 1417 716
rect 1423 676 1427 716
rect 1495 676 1499 716
rect 1515 696 1519 716
rect 1525 696 1529 716
rect 1547 696 1551 716
rect 1557 696 1561 716
rect 1579 696 1583 716
rect 1625 696 1629 716
rect 1633 696 1637 716
rect 1653 696 1657 716
rect 1663 696 1667 716
rect 1685 676 1689 716
rect 1735 676 1739 716
rect 1755 696 1759 716
rect 1765 696 1769 716
rect 1787 696 1791 716
rect 1797 696 1801 716
rect 1819 696 1823 716
rect 1865 696 1869 716
rect 1873 696 1877 716
rect 1893 696 1897 716
rect 1903 696 1907 716
rect 1925 676 1929 716
rect 1975 676 1979 716
rect 1995 696 1999 716
rect 2005 696 2009 716
rect 2027 696 2031 716
rect 2037 696 2041 716
rect 2059 696 2063 716
rect 2105 696 2109 716
rect 2113 696 2117 716
rect 2133 696 2137 716
rect 2143 696 2147 716
rect 2165 676 2169 716
rect 2215 676 2219 716
rect 2235 696 2239 716
rect 2245 696 2249 716
rect 2267 696 2271 716
rect 2277 696 2281 716
rect 2299 696 2303 716
rect 2345 696 2349 716
rect 2353 696 2357 716
rect 2373 696 2377 716
rect 2383 696 2387 716
rect 2405 676 2409 716
rect 2451 676 2455 716
rect 2473 696 2477 716
rect 2483 696 2487 716
rect 2503 696 2507 716
rect 2511 696 2515 716
rect 2557 696 2561 716
rect 2579 696 2583 716
rect 2589 696 2593 716
rect 2611 696 2615 716
rect 2621 696 2625 716
rect 2641 676 2645 716
rect 2726 676 2730 716
rect 2734 676 2738 716
rect 2754 676 2758 716
rect 2762 676 2766 716
rect 2825 696 2829 716
rect 2892 696 2896 716
rect 2914 676 2918 716
rect 2922 676 2926 716
rect 2971 696 2975 716
rect 3031 676 3035 716
rect 3051 676 3055 716
rect 3071 676 3075 716
rect 3133 676 3137 716
rect 3143 676 3147 716
rect 3212 656 3216 716
rect 3220 656 3224 716
rect 3228 656 3232 716
rect 3311 696 3315 716
rect 3371 676 3375 716
rect 3391 676 3395 716
rect 3411 676 3415 716
rect 3473 676 3477 716
rect 3483 676 3487 716
rect 3554 676 3558 716
rect 3562 676 3566 716
rect 3584 696 3588 716
rect 3651 696 3655 716
rect 3671 696 3675 716
rect 3731 676 3735 716
rect 3751 676 3755 716
rect 3771 676 3775 716
rect 3868 656 3872 716
rect 3876 656 3880 716
rect 3884 656 3888 716
rect 3931 676 3935 716
rect 3953 696 3957 716
rect 3963 696 3967 716
rect 3983 696 3987 716
rect 3991 696 3995 716
rect 4037 696 4041 716
rect 4059 696 4063 716
rect 4069 696 4073 716
rect 4091 696 4095 716
rect 4101 696 4105 716
rect 4121 676 4125 716
rect 4185 696 4189 716
rect 4205 696 4209 716
rect 4251 676 4255 716
rect 4273 696 4277 716
rect 4283 696 4287 716
rect 4303 696 4307 716
rect 4311 696 4315 716
rect 4357 696 4361 716
rect 4379 696 4383 716
rect 4389 696 4393 716
rect 4411 696 4415 716
rect 4421 696 4425 716
rect 4441 676 4445 716
rect 4491 696 4495 716
rect 4554 676 4558 716
rect 4562 676 4566 716
rect 4582 676 4586 716
rect 4590 676 4594 716
rect 4692 696 4696 716
rect 4714 676 4718 716
rect 4722 676 4726 716
rect 4785 676 4789 716
rect 4805 676 4809 716
rect 4825 676 4829 716
rect 4873 676 4877 716
rect 4883 676 4887 716
rect 4965 696 4969 716
rect 5025 668 5029 708
rect 5035 668 5039 708
rect 5055 668 5059 708
rect 5065 668 5069 708
rect 5085 688 5089 708
rect 5132 656 5136 716
rect 5140 656 5144 716
rect 5148 656 5152 716
rect 5231 676 5235 716
rect 5253 696 5257 716
rect 5263 696 5267 716
rect 5283 696 5287 716
rect 5291 696 5295 716
rect 5337 696 5341 716
rect 5359 696 5363 716
rect 5369 696 5373 716
rect 5391 696 5395 716
rect 5401 696 5405 716
rect 5421 676 5425 716
rect 5471 676 5475 716
rect 5531 688 5535 708
rect 5551 668 5555 708
rect 5561 668 5565 708
rect 5581 668 5585 708
rect 5591 668 5595 708
rect 5665 696 5669 716
rect 5685 696 5689 716
rect 5745 696 5749 716
rect 5765 696 5769 716
rect 5825 696 5829 716
rect 5845 696 5849 716
rect 5891 696 5895 716
rect 5911 696 5915 716
rect 5985 696 5989 716
rect 6005 696 6009 716
rect 6051 676 6055 716
rect 6071 676 6075 716
rect 6091 676 6095 716
rect 6151 676 6155 716
rect 6171 676 6175 716
rect 6191 676 6195 716
rect 6273 676 6277 716
rect 6283 676 6287 716
rect 6335 676 6339 716
rect 6355 696 6359 716
rect 6365 696 6369 716
rect 6387 696 6391 716
rect 6397 696 6401 716
rect 6419 696 6423 716
rect 6465 696 6469 716
rect 6473 696 6477 716
rect 6493 696 6497 716
rect 6503 696 6507 716
rect 6525 676 6529 716
rect 6571 696 6575 716
rect 6631 696 6635 716
rect 31 264 35 304
rect 53 264 57 284
rect 63 264 67 284
rect 83 264 87 284
rect 91 264 95 284
rect 137 264 141 284
rect 159 264 163 284
rect 169 264 173 284
rect 191 264 195 284
rect 201 264 205 284
rect 221 264 225 304
rect 275 264 279 304
rect 295 264 299 284
rect 305 264 309 284
rect 327 264 331 284
rect 337 264 341 284
rect 359 264 363 284
rect 405 264 409 284
rect 413 264 417 284
rect 433 264 437 284
rect 443 264 447 284
rect 465 264 469 304
rect 512 264 516 324
rect 520 264 524 324
rect 528 264 532 324
rect 611 264 615 284
rect 631 264 635 284
rect 705 264 709 284
rect 725 264 729 284
rect 773 264 777 304
rect 783 264 787 304
rect 865 264 869 284
rect 915 264 919 304
rect 935 264 939 284
rect 945 264 949 284
rect 967 264 971 284
rect 977 264 981 284
rect 999 264 1003 284
rect 1045 264 1049 284
rect 1053 264 1057 284
rect 1073 264 1077 284
rect 1083 264 1087 284
rect 1105 264 1109 304
rect 1163 264 1167 304
rect 1185 264 1189 284
rect 1231 264 1235 284
rect 1253 264 1257 304
rect 1311 264 1315 284
rect 1333 264 1337 304
rect 1405 264 1409 284
rect 1451 264 1455 304
rect 1471 264 1475 304
rect 1491 264 1495 304
rect 1565 264 1569 284
rect 1611 264 1615 304
rect 1631 264 1635 304
rect 1651 264 1655 304
rect 1715 264 1719 304
rect 1735 264 1739 284
rect 1745 264 1749 284
rect 1767 264 1771 284
rect 1777 264 1781 284
rect 1799 264 1803 284
rect 1845 264 1849 284
rect 1853 264 1857 284
rect 1873 264 1877 284
rect 1883 264 1887 284
rect 1905 264 1909 304
rect 1965 264 1969 284
rect 2025 264 2029 284
rect 2071 264 2075 304
rect 2091 264 2095 304
rect 2111 264 2115 304
rect 2171 264 2175 284
rect 2231 264 2235 304
rect 2251 264 2255 304
rect 2271 264 2275 304
rect 2291 264 2295 304
rect 2365 264 2369 304
rect 2385 264 2389 304
rect 2405 264 2409 304
rect 2451 264 2455 284
rect 2471 264 2475 284
rect 2535 264 2539 304
rect 2555 264 2559 284
rect 2565 264 2569 284
rect 2587 264 2591 284
rect 2597 264 2601 284
rect 2619 264 2623 284
rect 2665 264 2669 284
rect 2673 264 2677 284
rect 2693 264 2697 284
rect 2703 264 2707 284
rect 2725 264 2729 304
rect 2785 264 2789 304
rect 2805 264 2809 304
rect 2825 264 2829 304
rect 2871 264 2875 284
rect 2891 264 2895 284
rect 2955 264 2959 304
rect 2975 264 2979 284
rect 2985 264 2989 284
rect 3007 264 3011 284
rect 3017 264 3021 284
rect 3039 264 3043 284
rect 3085 264 3089 284
rect 3093 264 3097 284
rect 3113 264 3117 284
rect 3123 264 3127 284
rect 3145 264 3149 304
rect 3193 264 3197 304
rect 3203 264 3207 304
rect 3285 264 3289 304
rect 3305 264 3309 304
rect 3325 264 3329 304
rect 3371 264 3375 284
rect 3391 264 3395 284
rect 3472 264 3476 284
rect 3494 264 3498 304
rect 3502 264 3506 304
rect 3551 264 3555 304
rect 3571 264 3575 304
rect 3591 264 3595 304
rect 3651 264 3655 284
rect 3671 264 3675 284
rect 3734 264 3738 304
rect 3742 264 3746 304
rect 3764 264 3768 284
rect 3845 264 3849 284
rect 3865 264 3869 284
rect 3911 264 3915 304
rect 3931 264 3935 304
rect 3951 264 3955 304
rect 4048 264 4052 324
rect 4056 264 4060 324
rect 4064 264 4068 324
rect 4111 264 4115 284
rect 4131 264 4135 284
rect 4191 264 4195 304
rect 4213 264 4217 284
rect 4223 264 4227 284
rect 4243 264 4247 284
rect 4251 264 4255 284
rect 4297 264 4301 284
rect 4319 264 4323 284
rect 4329 264 4333 284
rect 4351 264 4355 284
rect 4361 264 4365 284
rect 4381 264 4385 304
rect 4431 264 4435 284
rect 4451 264 4455 284
rect 4525 264 4529 304
rect 4545 264 4549 304
rect 4565 264 4569 304
rect 4611 264 4615 284
rect 4631 264 4635 284
rect 4705 264 4709 304
rect 4725 264 4729 304
rect 4745 264 4749 304
rect 4765 264 4769 304
rect 4825 264 4829 284
rect 4875 264 4879 304
rect 4895 264 4899 284
rect 4905 264 4909 284
rect 4927 264 4931 284
rect 4937 264 4941 284
rect 4959 264 4963 284
rect 5005 264 5009 284
rect 5013 264 5017 284
rect 5033 264 5037 284
rect 5043 264 5047 284
rect 5065 264 5069 304
rect 5132 264 5136 284
rect 5154 264 5158 304
rect 5162 264 5166 304
rect 5211 264 5215 284
rect 5231 264 5235 284
rect 5305 264 5309 304
rect 5325 264 5329 304
rect 5345 264 5349 304
rect 5391 264 5395 284
rect 5411 264 5415 284
rect 5474 264 5478 304
rect 5482 264 5486 304
rect 5504 264 5508 284
rect 5572 264 5576 324
rect 5580 264 5584 324
rect 5588 264 5592 324
rect 5671 264 5675 304
rect 5691 264 5695 304
rect 5711 264 5715 304
rect 5793 264 5797 304
rect 5803 264 5807 304
rect 5865 264 5869 304
rect 5885 264 5889 304
rect 5905 264 5909 304
rect 5951 264 5955 304
rect 5971 264 5975 304
rect 5991 264 5995 304
rect 6051 264 6055 304
rect 6071 264 6075 304
rect 6091 264 6095 304
rect 6165 264 6169 284
rect 6185 264 6189 284
rect 6245 264 6249 284
rect 6265 264 6269 284
rect 6325 264 6329 304
rect 6345 264 6349 304
rect 6365 264 6369 304
rect 6385 264 6389 304
rect 6435 264 6439 304
rect 6455 264 6459 284
rect 6465 264 6469 284
rect 6487 264 6491 284
rect 6497 264 6501 284
rect 6519 264 6523 284
rect 6565 264 6569 284
rect 6573 264 6577 284
rect 6593 264 6597 284
rect 6603 264 6607 284
rect 6625 264 6629 304
rect 31 196 35 236
rect 53 216 57 236
rect 63 216 67 236
rect 83 216 87 236
rect 91 216 95 236
rect 137 216 141 236
rect 159 216 163 236
rect 169 216 173 236
rect 191 216 195 236
rect 201 216 205 236
rect 221 196 225 236
rect 271 196 275 236
rect 293 216 297 236
rect 303 216 307 236
rect 323 216 327 236
rect 331 216 335 236
rect 377 216 381 236
rect 399 216 403 236
rect 409 216 413 236
rect 431 216 435 236
rect 441 216 445 236
rect 461 196 465 236
rect 523 196 527 236
rect 545 216 549 236
rect 591 216 595 236
rect 613 196 617 236
rect 683 196 687 236
rect 705 216 709 236
rect 751 196 755 236
rect 773 216 777 236
rect 783 216 787 236
rect 803 216 807 236
rect 811 216 815 236
rect 857 216 861 236
rect 879 216 883 236
rect 889 216 893 236
rect 911 216 915 236
rect 921 216 925 236
rect 941 196 945 236
rect 991 216 995 236
rect 1013 196 1017 236
rect 1093 196 1097 236
rect 1103 196 1107 236
rect 1165 196 1169 236
rect 1185 196 1189 236
rect 1205 196 1209 236
rect 1255 196 1259 236
rect 1275 216 1279 236
rect 1285 216 1289 236
rect 1307 216 1311 236
rect 1317 216 1321 236
rect 1339 216 1343 236
rect 1385 216 1389 236
rect 1393 216 1397 236
rect 1413 216 1417 236
rect 1423 216 1427 236
rect 1445 196 1449 236
rect 1505 216 1509 236
rect 1553 196 1557 236
rect 1563 196 1567 236
rect 1645 196 1649 236
rect 1665 196 1669 236
rect 1685 196 1689 236
rect 1731 216 1735 236
rect 1793 196 1797 236
rect 1803 196 1807 236
rect 1873 196 1877 236
rect 1883 196 1887 236
rect 1953 196 1957 236
rect 1963 196 1967 236
rect 2045 196 2049 236
rect 2065 196 2069 236
rect 2085 196 2089 236
rect 2135 196 2139 236
rect 2155 216 2159 236
rect 2165 216 2169 236
rect 2187 216 2191 236
rect 2197 216 2201 236
rect 2219 216 2223 236
rect 2265 216 2269 236
rect 2273 216 2277 236
rect 2293 216 2297 236
rect 2303 216 2307 236
rect 2325 196 2329 236
rect 2373 196 2377 236
rect 2383 196 2387 236
rect 2473 196 2477 236
rect 2483 196 2487 236
rect 2545 196 2549 236
rect 2565 196 2569 236
rect 2585 196 2589 236
rect 2645 216 2649 236
rect 2695 196 2699 236
rect 2715 216 2719 236
rect 2725 216 2729 236
rect 2747 216 2751 236
rect 2757 216 2761 236
rect 2779 216 2783 236
rect 2825 216 2829 236
rect 2833 216 2837 236
rect 2853 216 2857 236
rect 2863 216 2867 236
rect 2885 196 2889 236
rect 2945 196 2949 236
rect 2965 196 2969 236
rect 2985 196 2989 236
rect 3045 216 3049 236
rect 3065 216 3069 236
rect 3125 196 3129 236
rect 3145 196 3149 236
rect 3165 196 3169 236
rect 3185 196 3189 236
rect 3245 216 3249 236
rect 3291 196 3295 236
rect 3313 216 3317 236
rect 3323 216 3327 236
rect 3343 216 3347 236
rect 3351 216 3355 236
rect 3397 216 3401 236
rect 3419 216 3423 236
rect 3429 216 3433 236
rect 3451 216 3455 236
rect 3461 216 3465 236
rect 3481 196 3485 236
rect 3553 196 3557 236
rect 3563 196 3567 236
rect 3625 196 3629 236
rect 3645 196 3649 236
rect 3665 196 3669 236
rect 3711 196 3715 236
rect 3731 196 3735 236
rect 3751 196 3755 236
rect 3811 196 3815 236
rect 3833 216 3837 236
rect 3843 216 3847 236
rect 3863 216 3867 236
rect 3871 216 3875 236
rect 3917 216 3921 236
rect 3939 216 3943 236
rect 3949 216 3953 236
rect 3971 216 3975 236
rect 3981 216 3985 236
rect 4001 196 4005 236
rect 4051 196 4055 236
rect 4071 196 4075 236
rect 4091 196 4095 236
rect 4151 196 4155 236
rect 4171 196 4175 236
rect 4191 196 4195 236
rect 4253 196 4257 236
rect 4263 196 4267 236
rect 4331 196 4335 236
rect 4353 216 4357 236
rect 4363 216 4367 236
rect 4383 216 4387 236
rect 4391 216 4395 236
rect 4437 216 4441 236
rect 4459 216 4463 236
rect 4469 216 4473 236
rect 4491 216 4495 236
rect 4501 216 4505 236
rect 4521 196 4525 236
rect 4571 196 4575 236
rect 4591 196 4595 236
rect 4611 196 4615 236
rect 4671 196 4675 236
rect 4691 196 4695 236
rect 4711 196 4715 236
rect 4773 196 4777 236
rect 4783 196 4787 236
rect 4851 196 4855 236
rect 4873 216 4877 236
rect 4883 216 4887 236
rect 4903 216 4907 236
rect 4911 216 4915 236
rect 4957 216 4961 236
rect 4979 216 4983 236
rect 4989 216 4993 236
rect 5011 216 5015 236
rect 5021 216 5025 236
rect 5041 196 5045 236
rect 5105 196 5109 236
rect 5125 196 5129 236
rect 5145 196 5149 236
rect 5191 196 5195 236
rect 5211 196 5215 236
rect 5231 196 5235 236
rect 5293 196 5297 236
rect 5303 196 5307 236
rect 5371 196 5375 236
rect 5393 216 5397 236
rect 5403 216 5407 236
rect 5423 216 5427 236
rect 5431 216 5435 236
rect 5477 216 5481 236
rect 5499 216 5503 236
rect 5509 216 5513 236
rect 5531 216 5535 236
rect 5541 216 5545 236
rect 5561 196 5565 236
rect 5611 196 5615 236
rect 5633 216 5637 236
rect 5643 216 5647 236
rect 5663 216 5667 236
rect 5671 216 5675 236
rect 5717 216 5721 236
rect 5739 216 5743 236
rect 5749 216 5753 236
rect 5771 216 5775 236
rect 5781 216 5785 236
rect 5801 196 5805 236
rect 5851 196 5855 236
rect 5873 216 5877 236
rect 5883 216 5887 236
rect 5903 216 5907 236
rect 5911 216 5915 236
rect 5957 216 5961 236
rect 5979 216 5983 236
rect 5989 216 5993 236
rect 6011 216 6015 236
rect 6021 216 6025 236
rect 6041 196 6045 236
rect 6105 196 6109 236
rect 6151 196 6155 236
rect 6171 196 6175 236
rect 6191 196 6195 236
rect 6265 196 6269 236
rect 6285 196 6289 236
rect 6305 196 6309 236
rect 6325 196 6329 236
rect 6385 216 6389 236
rect 6431 196 6435 236
rect 6453 216 6457 236
rect 6463 216 6467 236
rect 6483 216 6487 236
rect 6491 216 6495 236
rect 6537 216 6541 236
rect 6559 216 6563 236
rect 6569 216 6573 236
rect 6591 216 6595 236
rect 6601 216 6605 236
rect 6621 196 6625 236
<< ptransistor >>
rect 35 6264 39 6344
rect 55 6264 59 6304
rect 69 6264 73 6304
rect 89 6264 93 6304
rect 101 6264 105 6304
rect 121 6264 125 6304
rect 167 6264 171 6304
rect 175 6264 179 6304
rect 195 6264 199 6284
rect 203 6264 207 6284
rect 225 6264 229 6344
rect 290 6264 294 6304
rect 312 6264 316 6344
rect 320 6264 324 6344
rect 371 6264 375 6304
rect 391 6264 395 6304
rect 465 6264 469 6304
rect 485 6264 489 6304
rect 531 6264 535 6304
rect 551 6264 555 6304
rect 611 6264 615 6344
rect 633 6264 637 6284
rect 641 6264 645 6284
rect 661 6264 665 6304
rect 669 6264 673 6304
rect 715 6264 719 6304
rect 735 6264 739 6304
rect 747 6264 751 6304
rect 767 6264 771 6304
rect 781 6264 785 6304
rect 801 6264 805 6344
rect 851 6264 855 6304
rect 911 6264 915 6344
rect 931 6264 935 6344
rect 951 6264 955 6344
rect 971 6264 975 6344
rect 1045 6264 1049 6304
rect 1091 6264 1095 6344
rect 1113 6264 1117 6284
rect 1121 6264 1125 6284
rect 1141 6264 1145 6304
rect 1149 6264 1153 6304
rect 1195 6264 1199 6304
rect 1215 6264 1219 6304
rect 1227 6264 1231 6304
rect 1247 6264 1251 6304
rect 1261 6264 1265 6304
rect 1281 6264 1285 6344
rect 1331 6264 1335 6344
rect 1341 6264 1345 6344
rect 1371 6264 1375 6344
rect 1381 6264 1385 6344
rect 1470 6264 1474 6304
rect 1492 6264 1496 6344
rect 1500 6264 1504 6344
rect 1561 6264 1565 6344
rect 1583 6264 1587 6304
rect 1605 6264 1609 6304
rect 1665 6264 1669 6304
rect 1711 6264 1715 6344
rect 1733 6264 1737 6284
rect 1741 6264 1745 6284
rect 1761 6264 1765 6304
rect 1769 6264 1773 6304
rect 1815 6264 1819 6304
rect 1835 6264 1839 6304
rect 1847 6264 1851 6304
rect 1867 6264 1871 6304
rect 1881 6264 1885 6304
rect 1901 6264 1905 6344
rect 1956 6264 1960 6344
rect 1964 6264 1968 6344
rect 1986 6264 1990 6304
rect 2051 6264 2055 6304
rect 2071 6264 2075 6304
rect 2150 6264 2154 6304
rect 2172 6264 2176 6344
rect 2180 6264 2184 6344
rect 2245 6264 2249 6344
rect 2265 6264 2269 6344
rect 2285 6264 2289 6344
rect 2345 6264 2349 6304
rect 2365 6264 2369 6304
rect 2437 6264 2441 6344
rect 2445 6264 2449 6344
rect 2491 6264 2495 6344
rect 2499 6264 2503 6344
rect 2571 6264 2575 6304
rect 2591 6264 2595 6304
rect 2665 6264 2669 6304
rect 2685 6264 2689 6304
rect 2705 6264 2709 6304
rect 2751 6264 2755 6304
rect 2771 6264 2775 6304
rect 2845 6264 2849 6304
rect 2865 6264 2869 6304
rect 2885 6264 2889 6304
rect 2950 6264 2954 6304
rect 2972 6264 2976 6344
rect 2980 6264 2984 6344
rect 3050 6264 3054 6304
rect 3072 6264 3076 6344
rect 3080 6264 3084 6344
rect 3145 6264 3149 6304
rect 3205 6264 3209 6304
rect 3251 6264 3255 6344
rect 3271 6264 3275 6344
rect 3291 6264 3295 6344
rect 3356 6264 3360 6344
rect 3364 6264 3368 6344
rect 3386 6264 3390 6304
rect 3465 6264 3469 6344
rect 3485 6264 3489 6344
rect 3505 6264 3509 6344
rect 3565 6264 3569 6344
rect 3585 6264 3589 6344
rect 3605 6264 3609 6344
rect 3651 6264 3655 6304
rect 3671 6264 3675 6304
rect 3691 6264 3695 6304
rect 3770 6264 3774 6304
rect 3792 6264 3796 6344
rect 3800 6264 3804 6344
rect 3856 6264 3860 6344
rect 3864 6264 3868 6344
rect 3886 6264 3890 6304
rect 3951 6264 3955 6304
rect 4011 6264 4015 6304
rect 4031 6264 4035 6304
rect 4101 6264 4105 6344
rect 4123 6264 4127 6304
rect 4145 6264 4149 6304
rect 4191 6264 4195 6304
rect 4211 6264 4215 6304
rect 4285 6264 4289 6304
rect 4305 6264 4309 6304
rect 4325 6264 4329 6304
rect 4385 6264 4389 6304
rect 4405 6264 4409 6304
rect 4425 6264 4429 6304
rect 4485 6264 4489 6304
rect 4505 6264 4509 6304
rect 4525 6264 4529 6304
rect 4571 6264 4575 6304
rect 4631 6264 4635 6344
rect 4651 6264 4655 6344
rect 4671 6264 4675 6344
rect 4731 6264 4735 6344
rect 4751 6264 4755 6344
rect 4771 6264 4775 6344
rect 4836 6264 4840 6344
rect 4844 6264 4848 6344
rect 4866 6264 4870 6304
rect 4950 6264 4954 6304
rect 4972 6264 4976 6344
rect 4980 6264 4984 6344
rect 5036 6264 5040 6344
rect 5044 6264 5048 6344
rect 5066 6264 5070 6304
rect 5145 6264 5149 6304
rect 5165 6264 5169 6304
rect 5185 6264 5189 6304
rect 5245 6264 5249 6304
rect 5265 6264 5269 6304
rect 5285 6264 5289 6304
rect 5345 6264 5349 6304
rect 5365 6264 5369 6304
rect 5385 6264 5389 6304
rect 5431 6264 5435 6344
rect 5451 6264 5455 6344
rect 5471 6264 5475 6344
rect 5545 6264 5549 6344
rect 5565 6264 5569 6344
rect 5585 6264 5589 6344
rect 5645 6264 5649 6304
rect 5691 6264 5695 6344
rect 5711 6264 5715 6344
rect 5731 6264 5735 6344
rect 5791 6264 5795 6304
rect 5811 6264 5815 6304
rect 5831 6264 5835 6304
rect 5905 6264 5909 6344
rect 5925 6264 5929 6344
rect 5945 6264 5949 6344
rect 6005 6264 6009 6304
rect 6065 6264 6069 6344
rect 6085 6264 6089 6344
rect 6105 6264 6109 6344
rect 6170 6264 6174 6304
rect 6192 6264 6196 6344
rect 6200 6264 6204 6344
rect 6265 6264 6269 6344
rect 6285 6264 6289 6344
rect 6305 6264 6309 6344
rect 6351 6264 6355 6304
rect 6371 6264 6375 6304
rect 6391 6264 6395 6304
rect 6465 6264 6469 6304
rect 6485 6264 6489 6304
rect 6505 6264 6509 6304
rect 6551 6264 6555 6304
rect 6611 6264 6615 6344
rect 6631 6264 6635 6344
rect 6651 6264 6655 6344
rect 6671 6264 6675 6344
rect 31 6156 35 6236
rect 53 6216 57 6236
rect 61 6216 65 6236
rect 81 6196 85 6236
rect 89 6196 93 6236
rect 135 6196 139 6236
rect 155 6196 159 6236
rect 167 6196 171 6236
rect 187 6196 191 6236
rect 201 6196 205 6236
rect 221 6156 225 6236
rect 285 6156 289 6236
rect 305 6156 309 6236
rect 325 6156 329 6236
rect 385 6196 389 6236
rect 405 6196 409 6236
rect 451 6156 455 6236
rect 459 6156 463 6236
rect 545 6196 549 6236
rect 565 6196 569 6236
rect 616 6156 620 6236
rect 624 6156 628 6236
rect 646 6196 650 6236
rect 730 6196 734 6236
rect 752 6156 756 6236
rect 760 6156 764 6236
rect 811 6156 815 6236
rect 819 6156 823 6236
rect 905 6156 909 6236
rect 925 6156 929 6236
rect 945 6156 949 6236
rect 991 6156 995 6236
rect 1001 6156 1005 6236
rect 1021 6156 1025 6236
rect 1105 6196 1109 6236
rect 1151 6156 1155 6236
rect 1159 6156 1163 6236
rect 1250 6196 1254 6236
rect 1272 6156 1276 6236
rect 1280 6156 1284 6236
rect 1345 6196 1349 6236
rect 1405 6196 1409 6236
rect 1451 6156 1455 6236
rect 1459 6156 1463 6236
rect 1531 6156 1535 6236
rect 1539 6156 1543 6236
rect 1611 6196 1615 6236
rect 1671 6156 1675 6236
rect 1679 6156 1683 6236
rect 1751 6156 1755 6236
rect 1759 6156 1763 6236
rect 1836 6156 1840 6236
rect 1844 6156 1848 6236
rect 1866 6196 1870 6236
rect 1931 6196 1935 6236
rect 2005 6156 2009 6236
rect 2025 6156 2029 6236
rect 2045 6156 2049 6236
rect 2091 6196 2095 6236
rect 2170 6196 2174 6236
rect 2192 6156 2196 6236
rect 2200 6156 2204 6236
rect 2251 6196 2255 6236
rect 2330 6196 2334 6236
rect 2352 6156 2356 6236
rect 2360 6156 2364 6236
rect 2425 6196 2429 6236
rect 2445 6196 2449 6236
rect 2465 6196 2469 6236
rect 2525 6156 2529 6236
rect 2545 6156 2549 6236
rect 2565 6156 2569 6236
rect 2637 6156 2641 6236
rect 2645 6156 2649 6236
rect 2705 6196 2709 6236
rect 2725 6196 2729 6236
rect 2745 6196 2749 6236
rect 2805 6156 2809 6236
rect 2825 6156 2829 6236
rect 2845 6156 2849 6236
rect 2865 6156 2869 6236
rect 2925 6196 2929 6236
rect 2971 6196 2975 6236
rect 2991 6196 2995 6236
rect 3011 6196 3015 6236
rect 3085 6156 3089 6236
rect 3105 6156 3109 6236
rect 3125 6156 3129 6236
rect 3185 6196 3189 6236
rect 3205 6196 3209 6236
rect 3225 6196 3229 6236
rect 3285 6156 3289 6236
rect 3305 6156 3309 6236
rect 3325 6156 3329 6236
rect 3385 6196 3389 6236
rect 3445 6196 3449 6236
rect 3465 6196 3469 6236
rect 3485 6196 3489 6236
rect 3531 6196 3535 6236
rect 3551 6196 3555 6236
rect 3571 6196 3575 6236
rect 3631 6196 3635 6236
rect 3691 6156 3695 6236
rect 3711 6156 3715 6236
rect 3731 6156 3735 6236
rect 3805 6196 3809 6236
rect 3825 6196 3829 6236
rect 3871 6196 3875 6236
rect 3891 6196 3895 6236
rect 3970 6196 3974 6236
rect 3992 6156 3996 6236
rect 4000 6156 4004 6236
rect 4056 6156 4060 6236
rect 4064 6156 4068 6236
rect 4086 6196 4090 6236
rect 4177 6156 4181 6236
rect 4185 6156 4189 6236
rect 4231 6196 4235 6236
rect 4305 6196 4309 6236
rect 4325 6196 4329 6236
rect 4371 6196 4375 6236
rect 4393 6196 4397 6236
rect 4415 6156 4419 6236
rect 4490 6196 4494 6236
rect 4512 6156 4516 6236
rect 4520 6156 4524 6236
rect 4585 6156 4589 6236
rect 4605 6156 4609 6236
rect 4625 6156 4629 6236
rect 4671 6196 4675 6236
rect 4691 6196 4695 6236
rect 4711 6196 4715 6236
rect 4785 6156 4789 6236
rect 4805 6156 4809 6236
rect 4825 6156 4829 6236
rect 4885 6196 4889 6236
rect 4905 6196 4909 6236
rect 4925 6196 4929 6236
rect 4971 6196 4975 6236
rect 4991 6196 4995 6236
rect 5011 6196 5015 6236
rect 5090 6196 5094 6236
rect 5112 6156 5116 6236
rect 5120 6156 5124 6236
rect 5185 6196 5189 6236
rect 5205 6196 5209 6236
rect 5251 6196 5255 6236
rect 5273 6196 5277 6236
rect 5295 6156 5299 6236
rect 5356 6156 5360 6236
rect 5364 6156 5368 6236
rect 5386 6196 5390 6236
rect 5465 6156 5469 6236
rect 5485 6156 5489 6236
rect 5505 6156 5509 6236
rect 5565 6196 5569 6236
rect 5585 6196 5589 6236
rect 5605 6196 5609 6236
rect 5651 6196 5655 6236
rect 5671 6196 5675 6236
rect 5691 6196 5695 6236
rect 5765 6156 5769 6236
rect 5785 6156 5789 6236
rect 5805 6156 5809 6236
rect 5851 6196 5855 6236
rect 5871 6196 5875 6236
rect 5891 6196 5895 6236
rect 5956 6156 5960 6236
rect 5964 6156 5968 6236
rect 5986 6196 5990 6236
rect 6056 6156 6060 6236
rect 6064 6156 6068 6236
rect 6086 6196 6090 6236
rect 6151 6196 6155 6236
rect 6171 6196 6175 6236
rect 6191 6196 6195 6236
rect 6251 6196 6255 6236
rect 6271 6196 6275 6236
rect 6291 6196 6295 6236
rect 6365 6196 6369 6236
rect 6385 6196 6389 6236
rect 6405 6196 6409 6236
rect 6465 6156 6469 6236
rect 6485 6156 6489 6236
rect 6505 6156 6509 6236
rect 6551 6196 6555 6236
rect 6611 6196 6615 6236
rect 43 5784 47 5864
rect 65 5784 69 5824
rect 111 5784 115 5824
rect 131 5784 135 5824
rect 191 5784 195 5824
rect 211 5784 215 5824
rect 285 5784 289 5864
rect 305 5784 309 5864
rect 325 5784 329 5864
rect 385 5784 389 5824
rect 405 5784 409 5824
rect 451 5784 455 5824
rect 537 5784 541 5864
rect 545 5784 549 5864
rect 591 5784 595 5864
rect 599 5784 603 5864
rect 676 5784 680 5864
rect 684 5784 688 5864
rect 706 5784 710 5824
rect 785 5784 789 5824
rect 831 5784 835 5864
rect 839 5784 843 5864
rect 925 5784 929 5824
rect 945 5784 949 5824
rect 1010 5784 1014 5824
rect 1032 5784 1036 5864
rect 1040 5784 1044 5864
rect 1091 5784 1095 5864
rect 1099 5784 1103 5864
rect 1185 5784 1189 5824
rect 1231 5784 1235 5864
rect 1253 5784 1257 5804
rect 1261 5784 1265 5804
rect 1281 5784 1285 5824
rect 1289 5784 1293 5824
rect 1335 5784 1339 5824
rect 1355 5784 1359 5824
rect 1367 5784 1371 5824
rect 1387 5784 1391 5824
rect 1401 5784 1405 5824
rect 1421 5784 1425 5864
rect 1471 5784 1475 5824
rect 1491 5784 1495 5824
rect 1565 5784 1569 5824
rect 1585 5784 1589 5824
rect 1605 5784 1609 5824
rect 1670 5784 1674 5824
rect 1692 5784 1696 5864
rect 1700 5784 1704 5864
rect 1777 5784 1781 5864
rect 1785 5784 1789 5864
rect 1845 5784 1849 5824
rect 1865 5784 1869 5824
rect 1885 5784 1889 5824
rect 1931 5784 1935 5824
rect 2010 5784 2014 5824
rect 2032 5784 2036 5864
rect 2040 5784 2044 5864
rect 2091 5784 2095 5824
rect 2111 5784 2115 5824
rect 2131 5784 2135 5824
rect 2205 5784 2209 5864
rect 2225 5784 2229 5864
rect 2245 5784 2249 5864
rect 2296 5784 2300 5864
rect 2304 5784 2308 5864
rect 2326 5784 2330 5824
rect 2405 5784 2409 5824
rect 2425 5784 2429 5824
rect 2485 5784 2489 5824
rect 2505 5784 2509 5824
rect 2525 5784 2529 5824
rect 2585 5784 2589 5864
rect 2605 5784 2609 5864
rect 2625 5784 2629 5864
rect 2671 5784 2675 5824
rect 2691 5784 2695 5824
rect 2765 5784 2769 5824
rect 2785 5784 2789 5824
rect 2805 5784 2809 5824
rect 2865 5784 2869 5824
rect 2885 5784 2889 5824
rect 2905 5784 2909 5824
rect 2965 5784 2969 5824
rect 2985 5784 2989 5824
rect 3005 5784 3009 5824
rect 3065 5784 3069 5824
rect 3085 5784 3089 5824
rect 3105 5784 3109 5824
rect 3151 5784 3155 5824
rect 3171 5784 3175 5824
rect 3191 5784 3195 5824
rect 3270 5784 3274 5824
rect 3292 5784 3296 5864
rect 3300 5784 3304 5864
rect 3356 5784 3360 5864
rect 3364 5784 3368 5864
rect 3386 5784 3390 5824
rect 3465 5784 3469 5864
rect 3485 5784 3489 5864
rect 3505 5784 3509 5864
rect 3570 5784 3574 5824
rect 3592 5784 3596 5864
rect 3600 5784 3604 5864
rect 3665 5784 3669 5824
rect 3685 5784 3689 5824
rect 3705 5784 3709 5824
rect 3751 5784 3755 5864
rect 3771 5784 3775 5864
rect 3791 5784 3795 5864
rect 3865 5784 3869 5824
rect 3885 5784 3889 5824
rect 3905 5784 3909 5824
rect 3965 5784 3969 5864
rect 3985 5784 3989 5864
rect 4005 5784 4009 5864
rect 4065 5784 4069 5824
rect 4085 5784 4089 5824
rect 4105 5784 4109 5824
rect 4165 5784 4169 5864
rect 4185 5784 4189 5864
rect 4205 5784 4209 5864
rect 4251 5784 4255 5824
rect 4271 5784 4275 5824
rect 4291 5784 4295 5824
rect 4351 5784 4355 5824
rect 4371 5784 4375 5824
rect 4450 5784 4454 5824
rect 4472 5784 4476 5864
rect 4480 5784 4484 5864
rect 4557 5784 4561 5864
rect 4565 5784 4569 5864
rect 4611 5784 4615 5824
rect 4633 5784 4637 5824
rect 4655 5784 4659 5864
rect 4725 5784 4729 5864
rect 4745 5784 4749 5864
rect 4765 5784 4769 5864
rect 4811 5784 4815 5824
rect 4831 5784 4835 5824
rect 4905 5784 4909 5824
rect 4965 5784 4969 5824
rect 4985 5784 4989 5824
rect 5005 5784 5009 5824
rect 5051 5784 5055 5864
rect 5071 5784 5075 5864
rect 5091 5784 5095 5864
rect 5156 5784 5160 5864
rect 5164 5784 5168 5864
rect 5186 5784 5190 5824
rect 5256 5784 5260 5864
rect 5264 5784 5268 5864
rect 5286 5784 5290 5824
rect 5351 5784 5355 5864
rect 5371 5784 5375 5864
rect 5391 5784 5395 5864
rect 5411 5784 5415 5864
rect 5485 5784 5489 5824
rect 5505 5784 5509 5824
rect 5551 5784 5555 5824
rect 5625 5784 5629 5824
rect 5645 5784 5649 5824
rect 5665 5784 5669 5824
rect 5711 5784 5715 5864
rect 5731 5784 5735 5864
rect 5751 5784 5755 5864
rect 5830 5784 5834 5824
rect 5852 5784 5856 5864
rect 5860 5784 5864 5864
rect 5916 5784 5920 5864
rect 5924 5784 5928 5864
rect 5946 5784 5950 5824
rect 6030 5784 6034 5824
rect 6052 5784 6056 5864
rect 6060 5784 6064 5864
rect 6111 5784 6115 5864
rect 6131 5784 6135 5864
rect 6151 5784 6155 5864
rect 6171 5784 6175 5864
rect 6245 5784 6249 5824
rect 6265 5784 6269 5824
rect 6311 5784 6315 5824
rect 6333 5784 6337 5824
rect 6355 5784 6359 5864
rect 6416 5784 6420 5864
rect 6424 5784 6428 5864
rect 6446 5784 6450 5824
rect 6511 5784 6515 5824
rect 6531 5784 6535 5824
rect 6551 5784 6555 5824
rect 6611 5784 6615 5824
rect 6631 5784 6635 5824
rect 43 5676 47 5756
rect 65 5716 69 5756
rect 123 5676 127 5756
rect 145 5716 149 5756
rect 191 5676 195 5756
rect 213 5736 217 5756
rect 221 5736 225 5756
rect 241 5716 245 5756
rect 249 5716 253 5756
rect 295 5716 299 5756
rect 315 5716 319 5756
rect 327 5716 331 5756
rect 347 5716 351 5756
rect 361 5716 365 5756
rect 381 5676 385 5756
rect 457 5676 461 5756
rect 465 5676 469 5756
rect 511 5676 515 5756
rect 531 5676 535 5756
rect 551 5676 555 5756
rect 611 5716 615 5756
rect 631 5716 635 5756
rect 691 5716 695 5756
rect 713 5716 717 5756
rect 735 5676 739 5756
rect 791 5716 795 5756
rect 811 5716 815 5756
rect 871 5716 875 5756
rect 891 5716 895 5756
rect 951 5676 955 5756
rect 959 5676 963 5756
rect 1031 5716 1035 5756
rect 1091 5676 1095 5756
rect 1101 5676 1105 5756
rect 1121 5676 1125 5756
rect 1191 5676 1195 5756
rect 1199 5676 1203 5756
rect 1271 5716 1275 5756
rect 1331 5676 1335 5756
rect 1339 5676 1343 5756
rect 1411 5716 1415 5756
rect 1471 5676 1475 5756
rect 1493 5736 1497 5756
rect 1501 5736 1505 5756
rect 1521 5716 1525 5756
rect 1529 5716 1533 5756
rect 1575 5716 1579 5756
rect 1595 5716 1599 5756
rect 1607 5716 1611 5756
rect 1627 5716 1631 5756
rect 1641 5716 1645 5756
rect 1661 5676 1665 5756
rect 1711 5676 1715 5756
rect 1721 5676 1725 5756
rect 1751 5676 1755 5756
rect 1761 5676 1765 5756
rect 1850 5716 1854 5756
rect 1872 5676 1876 5756
rect 1880 5676 1884 5756
rect 1945 5716 1949 5756
rect 1965 5716 1969 5756
rect 2011 5716 2015 5756
rect 2085 5676 2089 5756
rect 2105 5676 2109 5756
rect 2125 5676 2129 5756
rect 2171 5676 2175 5756
rect 2179 5676 2183 5756
rect 2251 5716 2255 5756
rect 2271 5716 2275 5756
rect 2341 5688 2345 5748
rect 2361 5688 2365 5748
rect 2405 5696 2409 5756
rect 2425 5696 2429 5756
rect 2445 5696 2449 5756
rect 2465 5696 2469 5756
rect 2525 5716 2529 5756
rect 2545 5716 2549 5756
rect 2605 5716 2609 5756
rect 2625 5716 2629 5756
rect 2645 5716 2649 5756
rect 2705 5716 2709 5756
rect 2725 5716 2729 5756
rect 2745 5716 2749 5756
rect 2791 5716 2795 5756
rect 2811 5716 2815 5756
rect 2876 5676 2880 5756
rect 2884 5676 2888 5756
rect 2906 5716 2910 5756
rect 2985 5716 2989 5756
rect 3005 5716 3009 5756
rect 3025 5716 3029 5756
rect 3071 5676 3075 5756
rect 3091 5676 3095 5756
rect 3111 5676 3115 5756
rect 3190 5716 3194 5756
rect 3212 5676 3216 5756
rect 3220 5676 3224 5756
rect 3285 5716 3289 5756
rect 3331 5716 3335 5756
rect 3351 5716 3355 5756
rect 3371 5716 3375 5756
rect 3445 5716 3449 5756
rect 3465 5716 3469 5756
rect 3485 5716 3489 5756
rect 3545 5716 3549 5756
rect 3565 5716 3569 5756
rect 3585 5716 3589 5756
rect 3645 5716 3649 5756
rect 3710 5716 3714 5756
rect 3732 5676 3736 5756
rect 3740 5676 3744 5756
rect 3817 5676 3821 5756
rect 3825 5676 3829 5756
rect 3876 5676 3880 5756
rect 3884 5676 3888 5756
rect 3906 5716 3910 5756
rect 3985 5716 3989 5756
rect 4045 5676 4049 5756
rect 4065 5676 4069 5756
rect 4085 5676 4089 5756
rect 4105 5676 4109 5756
rect 4170 5716 4174 5756
rect 4192 5676 4196 5756
rect 4200 5676 4204 5756
rect 4265 5716 4269 5756
rect 4285 5716 4289 5756
rect 4305 5716 4309 5756
rect 4351 5716 4355 5756
rect 4430 5716 4434 5756
rect 4452 5676 4456 5756
rect 4460 5676 4464 5756
rect 4521 5676 4525 5756
rect 4543 5716 4547 5756
rect 4565 5716 4569 5756
rect 4611 5716 4615 5756
rect 4631 5716 4635 5756
rect 4710 5716 4714 5756
rect 4732 5676 4736 5756
rect 4740 5676 4744 5756
rect 4796 5676 4800 5756
rect 4804 5676 4808 5756
rect 4826 5716 4830 5756
rect 4905 5716 4909 5756
rect 4925 5716 4929 5756
rect 4945 5716 4949 5756
rect 4991 5676 4995 5756
rect 5011 5676 5015 5756
rect 5031 5676 5035 5756
rect 5096 5676 5100 5756
rect 5104 5676 5108 5756
rect 5126 5716 5130 5756
rect 5191 5716 5195 5756
rect 5211 5716 5215 5756
rect 5231 5716 5235 5756
rect 5291 5716 5295 5756
rect 5311 5716 5315 5756
rect 5371 5716 5375 5756
rect 5391 5716 5395 5756
rect 5411 5716 5415 5756
rect 5471 5676 5475 5756
rect 5491 5676 5495 5756
rect 5511 5676 5515 5756
rect 5571 5716 5575 5756
rect 5591 5716 5595 5756
rect 5665 5716 5669 5756
rect 5685 5716 5689 5756
rect 5731 5676 5735 5756
rect 5751 5676 5755 5756
rect 5771 5676 5775 5756
rect 5791 5676 5795 5756
rect 5870 5716 5874 5756
rect 5892 5676 5896 5756
rect 5900 5676 5904 5756
rect 5951 5716 5955 5756
rect 6011 5676 6015 5756
rect 6031 5676 6035 5756
rect 6051 5676 6055 5756
rect 6071 5676 6075 5756
rect 6131 5716 6135 5756
rect 6151 5716 6155 5756
rect 6171 5716 6175 5756
rect 6245 5716 6249 5756
rect 6291 5676 6295 5756
rect 6311 5676 6315 5756
rect 6331 5676 6335 5756
rect 6391 5716 6395 5756
rect 6411 5716 6415 5756
rect 6431 5716 6435 5756
rect 6491 5716 6495 5756
rect 6511 5716 6515 5756
rect 6531 5716 6535 5756
rect 6591 5716 6595 5756
rect 6611 5716 6615 5756
rect 6631 5716 6635 5756
rect 31 5304 35 5384
rect 53 5304 57 5324
rect 61 5304 65 5324
rect 81 5304 85 5344
rect 89 5304 93 5344
rect 135 5304 139 5344
rect 155 5304 159 5344
rect 167 5304 171 5344
rect 187 5304 191 5344
rect 201 5304 205 5344
rect 221 5304 225 5384
rect 271 5304 275 5344
rect 291 5304 295 5344
rect 365 5304 369 5384
rect 385 5304 389 5384
rect 405 5304 409 5384
rect 465 5304 469 5344
rect 485 5304 489 5344
rect 541 5304 545 5384
rect 563 5304 567 5344
rect 585 5304 589 5344
rect 631 5304 635 5384
rect 639 5304 643 5384
rect 711 5304 715 5384
rect 719 5304 723 5384
rect 791 5304 795 5344
rect 811 5304 815 5344
rect 871 5304 875 5344
rect 891 5304 895 5344
rect 951 5304 955 5344
rect 1011 5304 1015 5384
rect 1031 5304 1035 5384
rect 1051 5304 1055 5384
rect 1125 5304 1129 5384
rect 1145 5304 1149 5384
rect 1165 5304 1169 5384
rect 1185 5304 1189 5384
rect 1231 5304 1235 5384
rect 1253 5304 1257 5324
rect 1261 5304 1265 5324
rect 1281 5304 1285 5344
rect 1289 5304 1293 5344
rect 1335 5304 1339 5344
rect 1355 5304 1359 5344
rect 1367 5304 1371 5344
rect 1387 5304 1391 5344
rect 1401 5304 1405 5344
rect 1421 5304 1425 5384
rect 1485 5304 1489 5344
rect 1505 5304 1509 5344
rect 1525 5304 1529 5344
rect 1585 5304 1589 5344
rect 1605 5304 1609 5344
rect 1625 5304 1629 5344
rect 1685 5304 1689 5344
rect 1750 5304 1754 5344
rect 1772 5304 1776 5384
rect 1780 5304 1784 5384
rect 1841 5304 1845 5384
rect 1863 5304 1867 5344
rect 1885 5304 1889 5344
rect 1945 5304 1949 5344
rect 1965 5304 1969 5344
rect 2030 5304 2034 5344
rect 2052 5304 2056 5384
rect 2060 5304 2064 5384
rect 2111 5304 2115 5344
rect 2131 5304 2135 5344
rect 2205 5304 2209 5344
rect 2270 5304 2274 5344
rect 2292 5304 2296 5384
rect 2300 5304 2304 5384
rect 2351 5304 2355 5384
rect 2359 5304 2363 5384
rect 2445 5304 2449 5344
rect 2505 5304 2509 5384
rect 2525 5304 2529 5384
rect 2545 5304 2549 5384
rect 2596 5304 2600 5384
rect 2604 5304 2608 5384
rect 2626 5304 2630 5344
rect 2691 5304 2695 5344
rect 2711 5304 2715 5344
rect 2785 5304 2789 5344
rect 2805 5304 2809 5344
rect 2825 5304 2829 5344
rect 2885 5304 2889 5344
rect 2905 5304 2909 5344
rect 2977 5304 2981 5384
rect 2985 5304 2989 5384
rect 3036 5304 3040 5384
rect 3044 5304 3048 5384
rect 3066 5304 3070 5344
rect 3145 5304 3149 5344
rect 3165 5304 3169 5344
rect 3216 5304 3220 5384
rect 3224 5304 3228 5384
rect 3246 5304 3250 5344
rect 3321 5304 3325 5384
rect 3343 5304 3347 5344
rect 3365 5304 3369 5344
rect 3411 5304 3415 5384
rect 3419 5304 3423 5384
rect 3491 5304 3495 5384
rect 3501 5304 3505 5384
rect 3521 5304 3525 5384
rect 3596 5304 3600 5384
rect 3604 5304 3608 5384
rect 3626 5304 3630 5344
rect 3717 5304 3721 5384
rect 3725 5304 3729 5384
rect 3771 5304 3775 5384
rect 3781 5304 3785 5384
rect 3811 5304 3815 5384
rect 3821 5304 3825 5384
rect 3917 5304 3921 5384
rect 3925 5304 3929 5384
rect 3976 5304 3980 5384
rect 3984 5304 3988 5384
rect 4006 5304 4010 5344
rect 4085 5304 4089 5344
rect 4105 5304 4109 5344
rect 4125 5304 4129 5344
rect 4185 5304 4189 5344
rect 4205 5304 4209 5344
rect 4251 5304 4255 5344
rect 4330 5304 4334 5344
rect 4352 5304 4356 5384
rect 4360 5304 4364 5384
rect 4425 5304 4429 5344
rect 4445 5304 4449 5344
rect 4491 5304 4495 5344
rect 4511 5304 4515 5344
rect 4590 5304 4594 5344
rect 4612 5304 4616 5384
rect 4620 5304 4624 5384
rect 4690 5304 4694 5344
rect 4712 5304 4716 5384
rect 4720 5304 4724 5384
rect 4781 5304 4785 5384
rect 4803 5304 4807 5344
rect 4825 5304 4829 5344
rect 4890 5304 4894 5344
rect 4912 5304 4916 5384
rect 4920 5304 4924 5384
rect 4985 5304 4989 5344
rect 5005 5304 5009 5344
rect 5061 5304 5065 5384
rect 5083 5304 5087 5344
rect 5105 5304 5109 5344
rect 5151 5304 5155 5344
rect 5171 5304 5175 5344
rect 5236 5304 5240 5384
rect 5244 5304 5248 5384
rect 5266 5304 5270 5344
rect 5341 5304 5345 5384
rect 5363 5304 5367 5344
rect 5385 5304 5389 5344
rect 5436 5304 5440 5384
rect 5444 5304 5448 5384
rect 5466 5304 5470 5344
rect 5531 5304 5535 5344
rect 5551 5304 5555 5344
rect 5611 5304 5615 5344
rect 5631 5304 5635 5344
rect 5651 5304 5655 5344
rect 5721 5304 5725 5384
rect 5743 5304 5747 5344
rect 5765 5304 5769 5344
rect 5825 5304 5829 5384
rect 5845 5304 5849 5384
rect 5865 5304 5869 5384
rect 5885 5304 5889 5384
rect 5931 5304 5935 5344
rect 5951 5304 5955 5344
rect 6011 5304 6015 5344
rect 6031 5304 6035 5344
rect 6051 5304 6055 5344
rect 6111 5304 6115 5384
rect 6131 5304 6135 5384
rect 6151 5304 6155 5384
rect 6230 5304 6234 5344
rect 6252 5304 6256 5384
rect 6260 5304 6264 5384
rect 6316 5304 6320 5384
rect 6324 5304 6328 5384
rect 6346 5304 6350 5344
rect 6430 5304 6434 5344
rect 6452 5304 6456 5384
rect 6460 5304 6464 5384
rect 6525 5304 6529 5344
rect 6545 5304 6549 5344
rect 6565 5304 6569 5344
rect 6625 5304 6629 5384
rect 6645 5304 6649 5384
rect 6665 5304 6669 5384
rect 43 5196 47 5276
rect 65 5236 69 5276
rect 111 5196 115 5276
rect 133 5256 137 5276
rect 141 5256 145 5276
rect 161 5236 165 5276
rect 169 5236 173 5276
rect 215 5236 219 5276
rect 235 5236 239 5276
rect 247 5236 251 5276
rect 267 5236 271 5276
rect 281 5236 285 5276
rect 301 5196 305 5276
rect 351 5236 355 5276
rect 371 5236 375 5276
rect 445 5196 449 5276
rect 465 5196 469 5276
rect 485 5196 489 5276
rect 545 5236 549 5276
rect 565 5236 569 5276
rect 615 5196 619 5276
rect 635 5236 639 5276
rect 649 5236 653 5276
rect 669 5236 673 5276
rect 681 5236 685 5276
rect 701 5236 705 5276
rect 747 5236 751 5276
rect 755 5236 759 5276
rect 775 5256 779 5276
rect 783 5256 787 5276
rect 805 5196 809 5276
rect 851 5236 855 5276
rect 871 5236 875 5276
rect 950 5236 954 5276
rect 972 5196 976 5276
rect 980 5196 984 5276
rect 1050 5236 1054 5276
rect 1072 5196 1076 5276
rect 1080 5196 1084 5276
rect 1141 5196 1145 5276
rect 1163 5236 1167 5276
rect 1185 5236 1189 5276
rect 1231 5196 1235 5276
rect 1253 5256 1257 5276
rect 1261 5256 1265 5276
rect 1281 5236 1285 5276
rect 1289 5236 1293 5276
rect 1335 5236 1339 5276
rect 1355 5236 1359 5276
rect 1367 5236 1371 5276
rect 1387 5236 1391 5276
rect 1401 5236 1405 5276
rect 1421 5196 1425 5276
rect 1485 5236 1489 5276
rect 1505 5236 1509 5276
rect 1551 5236 1555 5276
rect 1571 5236 1575 5276
rect 1631 5196 1635 5276
rect 1653 5256 1657 5276
rect 1661 5256 1665 5276
rect 1681 5236 1685 5276
rect 1689 5236 1693 5276
rect 1735 5236 1739 5276
rect 1755 5236 1759 5276
rect 1767 5236 1771 5276
rect 1787 5236 1791 5276
rect 1801 5236 1805 5276
rect 1821 5196 1825 5276
rect 1885 5196 1889 5276
rect 1905 5196 1909 5276
rect 1925 5196 1929 5276
rect 1945 5196 1949 5276
rect 1991 5236 1995 5276
rect 2061 5196 2065 5276
rect 2083 5236 2087 5276
rect 2105 5236 2109 5276
rect 2151 5236 2155 5276
rect 2171 5236 2175 5276
rect 2255 5196 2259 5276
rect 2275 5196 2279 5276
rect 2285 5196 2289 5276
rect 2345 5236 2349 5276
rect 2365 5236 2369 5276
rect 2425 5236 2429 5276
rect 2445 5236 2449 5276
rect 2465 5236 2469 5276
rect 2537 5196 2541 5276
rect 2545 5196 2549 5276
rect 2591 5236 2595 5276
rect 2661 5196 2665 5276
rect 2683 5236 2687 5276
rect 2705 5236 2709 5276
rect 2751 5196 2755 5276
rect 2759 5196 2763 5276
rect 2845 5236 2849 5276
rect 2865 5236 2869 5276
rect 2925 5236 2929 5276
rect 2945 5236 2949 5276
rect 2991 5196 2995 5276
rect 3001 5196 3005 5276
rect 3021 5196 3025 5276
rect 3101 5196 3105 5276
rect 3123 5236 3127 5276
rect 3145 5236 3149 5276
rect 3191 5236 3195 5276
rect 3211 5236 3215 5276
rect 3285 5236 3289 5276
rect 3305 5236 3309 5276
rect 3325 5236 3329 5276
rect 3385 5236 3389 5276
rect 3445 5196 3449 5276
rect 3465 5196 3469 5276
rect 3485 5196 3489 5276
rect 3557 5196 3561 5276
rect 3565 5196 3569 5276
rect 3616 5196 3620 5276
rect 3624 5196 3628 5276
rect 3646 5236 3650 5276
rect 3730 5236 3734 5276
rect 3752 5196 3756 5276
rect 3760 5196 3764 5276
rect 3811 5196 3815 5276
rect 3819 5196 3823 5276
rect 3891 5236 3895 5276
rect 3911 5236 3915 5276
rect 3985 5236 3989 5276
rect 4005 5236 4009 5276
rect 4056 5196 4060 5276
rect 4064 5196 4068 5276
rect 4086 5236 4090 5276
rect 4165 5236 4169 5276
rect 4185 5236 4189 5276
rect 4241 5196 4245 5276
rect 4263 5236 4267 5276
rect 4285 5236 4289 5276
rect 4345 5236 4349 5276
rect 4365 5236 4369 5276
rect 4430 5236 4434 5276
rect 4452 5196 4456 5276
rect 4460 5196 4464 5276
rect 4530 5236 4534 5276
rect 4552 5196 4556 5276
rect 4560 5196 4564 5276
rect 4611 5236 4615 5276
rect 4631 5236 4635 5276
rect 4691 5236 4695 5276
rect 4711 5236 4715 5276
rect 4771 5236 4775 5276
rect 4845 5236 4849 5276
rect 4865 5236 4869 5276
rect 4885 5236 4889 5276
rect 4936 5196 4940 5276
rect 4944 5196 4948 5276
rect 4966 5236 4970 5276
rect 5031 5196 5035 5276
rect 5091 5236 5095 5276
rect 5111 5236 5115 5276
rect 5171 5196 5175 5276
rect 5191 5196 5195 5276
rect 5251 5236 5255 5276
rect 5271 5236 5275 5276
rect 5336 5196 5340 5276
rect 5344 5196 5348 5276
rect 5366 5236 5370 5276
rect 5431 5236 5435 5276
rect 5451 5236 5455 5276
rect 5471 5236 5475 5276
rect 5531 5236 5535 5276
rect 5551 5236 5555 5276
rect 5571 5236 5575 5276
rect 5631 5236 5635 5276
rect 5691 5236 5695 5276
rect 5711 5236 5715 5276
rect 5731 5236 5735 5276
rect 5796 5196 5800 5276
rect 5804 5196 5808 5276
rect 5826 5236 5830 5276
rect 5905 5236 5909 5276
rect 5925 5236 5929 5276
rect 5971 5236 5975 5276
rect 5991 5236 5995 5276
rect 6011 5236 6015 5276
rect 6071 5236 6075 5276
rect 6091 5236 6095 5276
rect 6165 5196 6169 5276
rect 6185 5196 6189 5276
rect 6205 5196 6209 5276
rect 6265 5236 6269 5276
rect 6325 5236 6329 5276
rect 6345 5236 6349 5276
rect 6365 5236 6369 5276
rect 6425 5236 6429 5276
rect 6445 5236 6449 5276
rect 6465 5236 6469 5276
rect 6511 5236 6515 5276
rect 6585 5236 6589 5276
rect 6605 5236 6609 5276
rect 6625 5236 6629 5276
rect 6671 5236 6675 5276
rect 6691 5236 6695 5276
rect 43 4824 47 4904
rect 65 4824 69 4864
rect 123 4824 127 4904
rect 145 4824 149 4864
rect 205 4824 209 4864
rect 225 4824 229 4864
rect 271 4824 275 4904
rect 293 4824 297 4844
rect 301 4824 305 4844
rect 321 4824 325 4864
rect 329 4824 333 4864
rect 375 4824 379 4864
rect 395 4824 399 4864
rect 407 4824 411 4864
rect 427 4824 431 4864
rect 441 4824 445 4864
rect 461 4824 465 4904
rect 525 4824 529 4904
rect 545 4824 549 4904
rect 565 4824 569 4904
rect 625 4824 629 4864
rect 645 4824 649 4864
rect 691 4824 695 4864
rect 711 4824 715 4864
rect 785 4824 789 4864
rect 805 4824 809 4864
rect 851 4824 855 4904
rect 873 4824 877 4844
rect 881 4824 885 4844
rect 901 4824 905 4864
rect 909 4824 913 4864
rect 955 4824 959 4864
rect 975 4824 979 4864
rect 987 4824 991 4864
rect 1007 4824 1011 4864
rect 1021 4824 1025 4864
rect 1041 4824 1045 4904
rect 1103 4824 1107 4904
rect 1125 4824 1129 4864
rect 1185 4824 1189 4904
rect 1205 4824 1209 4904
rect 1225 4824 1229 4904
rect 1285 4824 1289 4864
rect 1305 4824 1309 4864
rect 1363 4824 1367 4904
rect 1385 4824 1389 4864
rect 1431 4824 1435 4864
rect 1451 4824 1455 4864
rect 1525 4824 1529 4864
rect 1545 4824 1549 4864
rect 1610 4824 1614 4864
rect 1632 4824 1636 4904
rect 1640 4824 1644 4904
rect 1705 4824 1709 4864
rect 1725 4824 1729 4864
rect 1790 4824 1794 4864
rect 1812 4824 1816 4904
rect 1820 4824 1824 4904
rect 1871 4824 1875 4864
rect 1891 4824 1895 4864
rect 1970 4824 1974 4864
rect 1992 4824 1996 4904
rect 2000 4824 2004 4904
rect 2070 4824 2074 4864
rect 2092 4824 2096 4904
rect 2100 4824 2104 4904
rect 2161 4824 2165 4904
rect 2183 4824 2187 4864
rect 2205 4824 2209 4864
rect 2251 4824 2255 4864
rect 2337 4824 2341 4904
rect 2345 4824 2349 4904
rect 2415 4824 2419 4904
rect 2435 4824 2439 4904
rect 2445 4824 2449 4904
rect 2505 4824 2509 4864
rect 2525 4824 2529 4864
rect 2590 4824 2594 4864
rect 2612 4824 2616 4904
rect 2620 4824 2624 4904
rect 2690 4824 2694 4864
rect 2712 4824 2716 4904
rect 2720 4824 2724 4904
rect 2785 4824 2789 4864
rect 2836 4824 2840 4904
rect 2844 4824 2848 4904
rect 2866 4824 2870 4864
rect 2950 4824 2954 4864
rect 2972 4824 2976 4904
rect 2980 4824 2984 4904
rect 3050 4824 3054 4864
rect 3072 4824 3076 4904
rect 3080 4824 3084 4904
rect 3157 4824 3161 4904
rect 3165 4824 3169 4904
rect 3225 4824 3229 4904
rect 3285 4824 3289 4864
rect 3305 4824 3309 4864
rect 3370 4824 3374 4864
rect 3392 4824 3396 4904
rect 3400 4824 3404 4904
rect 3455 4824 3459 4904
rect 3475 4824 3479 4864
rect 3489 4824 3493 4864
rect 3509 4824 3513 4864
rect 3521 4824 3525 4864
rect 3541 4824 3545 4864
rect 3587 4824 3591 4864
rect 3595 4824 3599 4864
rect 3615 4824 3619 4844
rect 3623 4824 3627 4844
rect 3645 4824 3649 4904
rect 3696 4824 3700 4904
rect 3704 4824 3708 4904
rect 3726 4824 3730 4864
rect 3805 4824 3809 4904
rect 3825 4824 3829 4904
rect 3845 4824 3849 4904
rect 3905 4824 3909 4864
rect 3925 4824 3929 4864
rect 3945 4824 3949 4864
rect 4005 4824 4009 4904
rect 4025 4824 4029 4904
rect 4045 4824 4049 4904
rect 4105 4824 4109 4904
rect 4161 4824 4165 4904
rect 4183 4824 4187 4864
rect 4205 4824 4209 4864
rect 4265 4824 4269 4864
rect 4285 4824 4289 4864
rect 4331 4824 4335 4864
rect 4353 4824 4357 4864
rect 4375 4824 4379 4904
rect 4450 4824 4454 4864
rect 4472 4824 4476 4904
rect 4480 4824 4484 4904
rect 4531 4824 4535 4864
rect 4551 4824 4555 4864
rect 4571 4824 4575 4864
rect 4636 4824 4640 4904
rect 4644 4824 4648 4904
rect 4666 4824 4670 4864
rect 4745 4824 4749 4864
rect 4765 4824 4769 4864
rect 4821 4824 4825 4904
rect 4843 4824 4847 4864
rect 4865 4824 4869 4864
rect 4925 4824 4929 4864
rect 4945 4824 4949 4864
rect 4991 4824 4995 4864
rect 5011 4824 5015 4864
rect 5071 4824 5075 4864
rect 5093 4824 5097 4864
rect 5115 4824 5119 4904
rect 5185 4824 5189 4864
rect 5205 4824 5209 4864
rect 5261 4824 5265 4904
rect 5283 4824 5287 4864
rect 5305 4824 5309 4864
rect 5351 4824 5355 4864
rect 5373 4824 5377 4864
rect 5395 4824 5399 4904
rect 5465 4824 5469 4904
rect 5485 4824 5489 4904
rect 5505 4824 5509 4904
rect 5525 4824 5529 4904
rect 5585 4824 5589 4864
rect 5605 4824 5609 4864
rect 5651 4824 5655 4864
rect 5671 4824 5675 4864
rect 5691 4824 5695 4864
rect 5765 4824 5769 4904
rect 5785 4824 5789 4904
rect 5805 4824 5809 4904
rect 5865 4824 5869 4864
rect 5885 4824 5889 4864
rect 5905 4824 5909 4864
rect 5965 4824 5969 4864
rect 5985 4824 5989 4864
rect 6031 4824 6035 4904
rect 6051 4824 6055 4904
rect 6071 4824 6075 4904
rect 6091 4824 6095 4904
rect 6165 4824 6169 4864
rect 6185 4824 6189 4864
rect 6205 4824 6209 4864
rect 6256 4824 6260 4904
rect 6264 4824 6268 4904
rect 6286 4824 6290 4864
rect 6365 4824 6369 4864
rect 6385 4824 6389 4864
rect 6405 4824 6409 4864
rect 6465 4824 6469 4864
rect 6485 4824 6489 4864
rect 6505 4824 6509 4864
rect 6551 4824 6555 4864
rect 6571 4824 6575 4864
rect 6645 4824 6649 4864
rect 31 4716 35 4796
rect 51 4716 55 4796
rect 71 4716 75 4796
rect 91 4716 95 4796
rect 111 4716 115 4796
rect 131 4716 135 4796
rect 151 4716 155 4796
rect 171 4716 175 4796
rect 257 4716 261 4796
rect 265 4716 269 4796
rect 325 4756 329 4796
rect 385 4716 389 4796
rect 405 4716 409 4796
rect 425 4716 429 4796
rect 485 4756 489 4796
rect 557 4716 561 4796
rect 565 4716 569 4796
rect 621 4716 625 4796
rect 643 4756 647 4796
rect 665 4756 669 4796
rect 711 4716 715 4796
rect 719 4716 723 4796
rect 803 4716 807 4796
rect 825 4756 829 4796
rect 885 4756 889 4796
rect 905 4756 909 4796
rect 951 4716 955 4796
rect 973 4776 977 4796
rect 981 4776 985 4796
rect 1001 4756 1005 4796
rect 1009 4756 1013 4796
rect 1055 4756 1059 4796
rect 1075 4756 1079 4796
rect 1087 4756 1091 4796
rect 1107 4756 1111 4796
rect 1121 4756 1125 4796
rect 1141 4716 1145 4796
rect 1210 4756 1214 4796
rect 1232 4716 1236 4796
rect 1240 4716 1244 4796
rect 1305 4756 1309 4796
rect 1325 4756 1329 4796
rect 1371 4756 1375 4796
rect 1391 4756 1395 4796
rect 1470 4756 1474 4796
rect 1492 4716 1496 4796
rect 1500 4716 1504 4796
rect 1551 4716 1555 4796
rect 1559 4716 1563 4796
rect 1631 4716 1635 4796
rect 1639 4716 1643 4796
rect 1711 4756 1715 4796
rect 1771 4716 1775 4796
rect 1779 4716 1783 4796
rect 1856 4716 1860 4796
rect 1864 4716 1868 4796
rect 1886 4756 1890 4796
rect 1951 4716 1955 4796
rect 1973 4776 1977 4796
rect 1981 4776 1985 4796
rect 2001 4756 2005 4796
rect 2009 4756 2013 4796
rect 2055 4756 2059 4796
rect 2075 4756 2079 4796
rect 2087 4756 2091 4796
rect 2107 4756 2111 4796
rect 2121 4756 2125 4796
rect 2141 4716 2145 4796
rect 2205 4756 2209 4796
rect 2225 4756 2229 4796
rect 2295 4716 2299 4796
rect 2315 4716 2319 4796
rect 2325 4716 2329 4796
rect 2371 4756 2375 4796
rect 2391 4756 2395 4796
rect 2451 4716 2455 4796
rect 2459 4716 2463 4796
rect 2531 4716 2535 4796
rect 2551 4716 2555 4796
rect 2571 4716 2575 4796
rect 2645 4756 2649 4796
rect 2691 4716 2695 4796
rect 2713 4776 2717 4796
rect 2721 4776 2725 4796
rect 2741 4756 2745 4796
rect 2749 4756 2753 4796
rect 2795 4756 2799 4796
rect 2815 4756 2819 4796
rect 2827 4756 2831 4796
rect 2847 4756 2851 4796
rect 2861 4756 2865 4796
rect 2881 4716 2885 4796
rect 2936 4716 2940 4796
rect 2944 4716 2948 4796
rect 2966 4756 2970 4796
rect 3031 4716 3035 4796
rect 3053 4776 3057 4796
rect 3061 4776 3065 4796
rect 3081 4756 3085 4796
rect 3089 4756 3093 4796
rect 3135 4756 3139 4796
rect 3155 4756 3159 4796
rect 3167 4756 3171 4796
rect 3187 4756 3191 4796
rect 3201 4756 3205 4796
rect 3221 4716 3225 4796
rect 3271 4716 3275 4796
rect 3293 4776 3297 4796
rect 3301 4776 3305 4796
rect 3321 4756 3325 4796
rect 3329 4756 3333 4796
rect 3375 4756 3379 4796
rect 3395 4756 3399 4796
rect 3407 4756 3411 4796
rect 3427 4756 3431 4796
rect 3441 4756 3445 4796
rect 3461 4716 3465 4796
rect 3530 4756 3534 4796
rect 3552 4716 3556 4796
rect 3560 4716 3564 4796
rect 3625 4716 3629 4796
rect 3685 4756 3689 4796
rect 3705 4756 3709 4796
rect 3770 4756 3774 4796
rect 3792 4716 3796 4796
rect 3800 4716 3804 4796
rect 3855 4716 3859 4796
rect 3875 4756 3879 4796
rect 3889 4756 3893 4796
rect 3909 4756 3913 4796
rect 3921 4756 3925 4796
rect 3941 4756 3945 4796
rect 3987 4756 3991 4796
rect 3995 4756 3999 4796
rect 4015 4776 4019 4796
rect 4023 4776 4027 4796
rect 4045 4716 4049 4796
rect 4105 4716 4109 4796
rect 4165 4756 4169 4796
rect 4185 4756 4189 4796
rect 4231 4716 4235 4796
rect 4253 4776 4257 4796
rect 4261 4776 4265 4796
rect 4281 4756 4285 4796
rect 4289 4756 4293 4796
rect 4335 4756 4339 4796
rect 4355 4756 4359 4796
rect 4367 4756 4371 4796
rect 4387 4756 4391 4796
rect 4401 4756 4405 4796
rect 4421 4716 4425 4796
rect 4485 4756 4489 4796
rect 4505 4756 4509 4796
rect 4525 4756 4529 4796
rect 4571 4756 4575 4796
rect 4631 4716 4635 4796
rect 4705 4756 4709 4796
rect 4756 4716 4760 4796
rect 4764 4716 4768 4796
rect 4786 4756 4790 4796
rect 4851 4716 4855 4796
rect 4859 4716 4863 4796
rect 4931 4756 4935 4796
rect 4951 4756 4955 4796
rect 5011 4756 5015 4796
rect 5031 4756 5035 4796
rect 5105 4756 5109 4796
rect 5125 4756 5129 4796
rect 5176 4716 5180 4796
rect 5184 4716 5188 4796
rect 5206 4756 5210 4796
rect 5295 4716 5299 4796
rect 5305 4716 5309 4796
rect 5335 4716 5339 4796
rect 5345 4716 5349 4796
rect 5391 4756 5395 4796
rect 5411 4756 5415 4796
rect 5485 4756 5489 4796
rect 5505 4756 5509 4796
rect 5551 4756 5555 4796
rect 5571 4756 5575 4796
rect 5591 4756 5595 4796
rect 5665 4756 5669 4796
rect 5685 4756 5689 4796
rect 5731 4756 5735 4796
rect 5751 4756 5755 4796
rect 5771 4756 5775 4796
rect 5845 4756 5849 4796
rect 5891 4756 5895 4796
rect 5911 4756 5915 4796
rect 5931 4756 5935 4796
rect 6001 4716 6005 4796
rect 6023 4756 6027 4796
rect 6045 4756 6049 4796
rect 6096 4716 6100 4796
rect 6104 4716 6108 4796
rect 6126 4756 6130 4796
rect 6205 4756 6209 4796
rect 6225 4756 6229 4796
rect 6271 4716 6275 4796
rect 6291 4716 6295 4796
rect 6311 4716 6315 4796
rect 6371 4756 6375 4796
rect 6391 4756 6395 4796
rect 6411 4756 6415 4796
rect 6481 4716 6485 4796
rect 6503 4756 6507 4796
rect 6525 4756 6529 4796
rect 6585 4756 6589 4796
rect 6605 4756 6609 4796
rect 6625 4756 6629 4796
rect 45 4344 49 4384
rect 117 4344 121 4424
rect 125 4344 129 4424
rect 185 4344 189 4384
rect 236 4344 240 4424
rect 244 4344 248 4424
rect 266 4344 270 4384
rect 357 4344 361 4424
rect 365 4344 369 4424
rect 416 4344 420 4424
rect 424 4344 428 4424
rect 446 4344 450 4384
rect 511 4344 515 4424
rect 521 4344 525 4424
rect 541 4344 545 4424
rect 611 4344 615 4424
rect 631 4344 635 4424
rect 651 4344 655 4424
rect 725 4344 729 4384
rect 771 4344 775 4424
rect 779 4344 783 4424
rect 851 4344 855 4384
rect 911 4344 915 4424
rect 919 4344 923 4424
rect 991 4344 995 4384
rect 1051 4344 1055 4424
rect 1071 4344 1075 4424
rect 1091 4344 1095 4424
rect 1111 4344 1115 4424
rect 1131 4344 1135 4424
rect 1151 4344 1155 4424
rect 1171 4344 1175 4424
rect 1191 4344 1195 4424
rect 1251 4344 1255 4384
rect 1273 4344 1277 4424
rect 1345 4344 1349 4384
rect 1417 4344 1421 4424
rect 1425 4344 1429 4424
rect 1485 4344 1489 4384
rect 1505 4344 1509 4384
rect 1551 4344 1555 4384
rect 1571 4344 1575 4384
rect 1645 4344 1649 4424
rect 1665 4344 1669 4424
rect 1685 4344 1689 4424
rect 1705 4344 1709 4424
rect 1755 4344 1759 4424
rect 1775 4344 1779 4384
rect 1789 4344 1793 4384
rect 1809 4344 1813 4384
rect 1821 4344 1825 4384
rect 1841 4344 1845 4384
rect 1887 4344 1891 4384
rect 1895 4344 1899 4384
rect 1915 4344 1919 4364
rect 1923 4344 1927 4364
rect 1945 4344 1949 4424
rect 1991 4344 1995 4384
rect 2011 4344 2015 4384
rect 2071 4344 2075 4424
rect 2093 4344 2097 4364
rect 2101 4344 2105 4364
rect 2121 4344 2125 4384
rect 2129 4344 2133 4384
rect 2175 4344 2179 4384
rect 2195 4344 2199 4384
rect 2207 4344 2211 4384
rect 2227 4344 2231 4384
rect 2241 4344 2245 4384
rect 2261 4344 2265 4424
rect 2311 4344 2315 4384
rect 2371 4344 2375 4424
rect 2379 4344 2383 4424
rect 2451 4344 2455 4424
rect 2459 4344 2463 4424
rect 2531 4344 2535 4384
rect 2591 4344 2595 4424
rect 2613 4344 2617 4364
rect 2621 4344 2625 4364
rect 2641 4344 2645 4384
rect 2649 4344 2653 4384
rect 2695 4344 2699 4384
rect 2715 4344 2719 4384
rect 2727 4344 2731 4384
rect 2747 4344 2751 4384
rect 2761 4344 2765 4384
rect 2781 4344 2785 4424
rect 2836 4344 2840 4424
rect 2844 4344 2848 4424
rect 2866 4344 2870 4384
rect 2931 4344 2935 4384
rect 2951 4344 2955 4384
rect 3025 4344 3029 4384
rect 3076 4344 3080 4424
rect 3084 4344 3088 4424
rect 3106 4344 3110 4384
rect 3171 4344 3175 4424
rect 3193 4344 3197 4364
rect 3201 4344 3205 4364
rect 3221 4344 3225 4384
rect 3229 4344 3233 4384
rect 3275 4344 3279 4384
rect 3295 4344 3299 4384
rect 3307 4344 3311 4384
rect 3327 4344 3331 4384
rect 3341 4344 3345 4384
rect 3361 4344 3365 4424
rect 3416 4344 3420 4424
rect 3424 4344 3428 4424
rect 3446 4344 3450 4384
rect 3530 4344 3534 4384
rect 3552 4344 3556 4424
rect 3560 4344 3564 4424
rect 3615 4344 3619 4424
rect 3635 4344 3639 4384
rect 3649 4344 3653 4384
rect 3669 4344 3673 4384
rect 3681 4344 3685 4384
rect 3701 4344 3705 4384
rect 3747 4344 3751 4384
rect 3755 4344 3759 4384
rect 3775 4344 3779 4364
rect 3783 4344 3787 4364
rect 3805 4344 3809 4424
rect 3856 4344 3860 4424
rect 3864 4344 3868 4424
rect 3886 4344 3890 4384
rect 3955 4344 3959 4424
rect 3975 4344 3979 4384
rect 3989 4344 3993 4384
rect 4009 4344 4013 4384
rect 4021 4344 4025 4384
rect 4041 4344 4045 4384
rect 4087 4344 4091 4384
rect 4095 4344 4099 4384
rect 4115 4344 4119 4364
rect 4123 4344 4127 4364
rect 4145 4344 4149 4424
rect 4205 4344 4209 4384
rect 4225 4344 4229 4384
rect 4245 4344 4249 4384
rect 4296 4344 4300 4424
rect 4304 4344 4308 4424
rect 4326 4344 4330 4384
rect 4417 4344 4421 4424
rect 4425 4344 4429 4424
rect 4485 4344 4489 4424
rect 4505 4344 4509 4424
rect 4525 4344 4529 4424
rect 4571 4344 4575 4384
rect 4591 4344 4595 4384
rect 4611 4344 4615 4384
rect 4685 4344 4689 4384
rect 4736 4344 4740 4424
rect 4744 4344 4748 4424
rect 4766 4344 4770 4384
rect 4855 4344 4859 4424
rect 4875 4344 4879 4424
rect 4885 4344 4889 4424
rect 4945 4344 4949 4384
rect 4965 4344 4969 4384
rect 5025 4344 5029 4384
rect 5045 4344 5049 4384
rect 5065 4344 5069 4384
rect 5116 4344 5120 4424
rect 5124 4344 5128 4424
rect 5146 4344 5150 4384
rect 5235 4344 5239 4424
rect 5255 4344 5259 4424
rect 5265 4344 5269 4424
rect 5316 4344 5320 4424
rect 5324 4344 5328 4424
rect 5346 4344 5350 4384
rect 5411 4344 5415 4384
rect 5485 4344 5489 4384
rect 5505 4344 5509 4384
rect 5525 4344 5529 4384
rect 5571 4344 5575 4384
rect 5591 4344 5595 4384
rect 5656 4344 5660 4424
rect 5664 4344 5668 4424
rect 5686 4344 5690 4384
rect 5765 4344 5769 4384
rect 5785 4344 5789 4384
rect 5845 4344 5849 4384
rect 5865 4344 5869 4384
rect 5885 4344 5889 4384
rect 5950 4344 5954 4384
rect 5972 4344 5976 4424
rect 5980 4344 5984 4424
rect 6031 4344 6035 4384
rect 6105 4344 6109 4384
rect 6151 4344 6155 4384
rect 6171 4344 6175 4384
rect 6191 4344 6195 4384
rect 6270 4344 6274 4384
rect 6292 4344 6296 4424
rect 6300 4344 6304 4424
rect 6351 4344 6355 4384
rect 6371 4344 6375 4384
rect 6391 4344 6395 4384
rect 6451 4344 6455 4384
rect 6471 4344 6475 4384
rect 6491 4344 6495 4384
rect 6556 4344 6560 4424
rect 6564 4344 6568 4424
rect 6586 4344 6590 4384
rect 6651 4344 6655 4384
rect 43 4236 47 4316
rect 65 4276 69 4316
rect 130 4276 134 4316
rect 152 4236 156 4316
rect 160 4236 164 4316
rect 216 4236 220 4316
rect 224 4236 228 4316
rect 246 4276 250 4316
rect 315 4236 319 4316
rect 335 4276 339 4316
rect 349 4276 353 4316
rect 369 4276 373 4316
rect 381 4276 385 4316
rect 401 4276 405 4316
rect 447 4276 451 4316
rect 455 4276 459 4316
rect 475 4296 479 4316
rect 483 4296 487 4316
rect 505 4236 509 4316
rect 551 4276 555 4316
rect 571 4276 575 4316
rect 645 4236 649 4316
rect 665 4236 669 4316
rect 685 4236 689 4316
rect 705 4236 709 4316
rect 765 4276 769 4316
rect 811 4236 815 4316
rect 833 4296 837 4316
rect 841 4296 845 4316
rect 861 4276 865 4316
rect 869 4276 873 4316
rect 915 4276 919 4316
rect 935 4276 939 4316
rect 947 4276 951 4316
rect 967 4276 971 4316
rect 981 4276 985 4316
rect 1001 4236 1005 4316
rect 1051 4276 1055 4316
rect 1071 4276 1075 4316
rect 1131 4236 1135 4316
rect 1153 4296 1157 4316
rect 1161 4296 1165 4316
rect 1181 4276 1185 4316
rect 1189 4276 1193 4316
rect 1235 4276 1239 4316
rect 1255 4276 1259 4316
rect 1267 4276 1271 4316
rect 1287 4276 1291 4316
rect 1301 4276 1305 4316
rect 1321 4236 1325 4316
rect 1371 4276 1375 4316
rect 1391 4276 1395 4316
rect 1451 4276 1455 4316
rect 1530 4276 1534 4316
rect 1552 4236 1556 4316
rect 1560 4236 1564 4316
rect 1625 4236 1629 4316
rect 1645 4236 1649 4316
rect 1665 4236 1669 4316
rect 1725 4276 1729 4316
rect 1745 4276 1749 4316
rect 1791 4276 1795 4316
rect 1811 4276 1815 4316
rect 1871 4236 1875 4316
rect 1893 4296 1897 4316
rect 1901 4296 1905 4316
rect 1921 4276 1925 4316
rect 1929 4276 1933 4316
rect 1975 4276 1979 4316
rect 1995 4276 1999 4316
rect 2007 4276 2011 4316
rect 2027 4276 2031 4316
rect 2041 4276 2045 4316
rect 2061 4236 2065 4316
rect 2111 4276 2115 4316
rect 2131 4276 2135 4316
rect 2210 4276 2214 4316
rect 2232 4236 2236 4316
rect 2240 4236 2244 4316
rect 2295 4236 2299 4316
rect 2315 4276 2319 4316
rect 2329 4276 2333 4316
rect 2349 4276 2353 4316
rect 2361 4276 2365 4316
rect 2381 4276 2385 4316
rect 2427 4276 2431 4316
rect 2435 4276 2439 4316
rect 2455 4296 2459 4316
rect 2463 4296 2467 4316
rect 2485 4236 2489 4316
rect 2557 4236 2561 4316
rect 2565 4236 2569 4316
rect 2611 4276 2615 4316
rect 2676 4236 2680 4316
rect 2684 4236 2688 4316
rect 2706 4276 2710 4316
rect 2771 4276 2775 4316
rect 2791 4276 2795 4316
rect 2870 4276 2874 4316
rect 2892 4236 2896 4316
rect 2900 4236 2904 4316
rect 2951 4276 2955 4316
rect 3011 4236 3015 4316
rect 3019 4236 3023 4316
rect 3105 4276 3109 4316
rect 3151 4236 3155 4316
rect 3173 4296 3177 4316
rect 3181 4296 3185 4316
rect 3201 4276 3205 4316
rect 3209 4276 3213 4316
rect 3255 4276 3259 4316
rect 3275 4276 3279 4316
rect 3287 4276 3291 4316
rect 3307 4276 3311 4316
rect 3321 4276 3325 4316
rect 3341 4236 3345 4316
rect 3391 4236 3395 4316
rect 3401 4236 3405 4316
rect 3431 4236 3435 4316
rect 3441 4236 3445 4316
rect 3511 4276 3515 4316
rect 3531 4276 3535 4316
rect 3591 4236 3595 4316
rect 3611 4236 3615 4316
rect 3631 4236 3635 4316
rect 3651 4236 3655 4316
rect 3671 4236 3675 4316
rect 3691 4236 3695 4316
rect 3711 4236 3715 4316
rect 3731 4236 3735 4316
rect 3791 4276 3795 4316
rect 3811 4276 3815 4316
rect 3871 4276 3875 4316
rect 3891 4276 3895 4316
rect 3965 4276 3969 4316
rect 3985 4276 3989 4316
rect 4031 4276 4035 4316
rect 4110 4276 4114 4316
rect 4132 4236 4136 4316
rect 4140 4236 4144 4316
rect 4196 4236 4200 4316
rect 4204 4236 4208 4316
rect 4226 4276 4230 4316
rect 4295 4236 4299 4316
rect 4315 4276 4319 4316
rect 4329 4276 4333 4316
rect 4349 4276 4353 4316
rect 4361 4276 4365 4316
rect 4381 4276 4385 4316
rect 4427 4276 4431 4316
rect 4435 4276 4439 4316
rect 4455 4296 4459 4316
rect 4463 4296 4467 4316
rect 4485 4236 4489 4316
rect 4550 4276 4554 4316
rect 4572 4236 4576 4316
rect 4580 4236 4584 4316
rect 4635 4236 4639 4316
rect 4655 4276 4659 4316
rect 4669 4276 4673 4316
rect 4689 4276 4693 4316
rect 4701 4276 4705 4316
rect 4721 4276 4725 4316
rect 4767 4276 4771 4316
rect 4775 4276 4779 4316
rect 4795 4296 4799 4316
rect 4803 4296 4807 4316
rect 4825 4236 4829 4316
rect 4885 4236 4889 4316
rect 4945 4236 4949 4316
rect 4965 4236 4969 4316
rect 4985 4236 4989 4316
rect 5031 4276 5035 4316
rect 5051 4276 5055 4316
rect 5071 4276 5075 4316
rect 5145 4276 5149 4316
rect 5196 4236 5200 4316
rect 5204 4236 5208 4316
rect 5226 4276 5230 4316
rect 5295 4236 5299 4316
rect 5315 4276 5319 4316
rect 5329 4276 5333 4316
rect 5349 4276 5353 4316
rect 5361 4276 5365 4316
rect 5381 4276 5385 4316
rect 5427 4276 5431 4316
rect 5435 4276 5439 4316
rect 5455 4296 5459 4316
rect 5463 4296 5467 4316
rect 5485 4236 5489 4316
rect 5531 4276 5535 4316
rect 5551 4276 5555 4316
rect 5611 4276 5615 4316
rect 5676 4236 5680 4316
rect 5684 4236 5688 4316
rect 5706 4276 5710 4316
rect 5781 4236 5785 4316
rect 5803 4276 5807 4316
rect 5825 4276 5829 4316
rect 5871 4276 5875 4316
rect 5891 4276 5895 4316
rect 5911 4276 5915 4316
rect 5985 4236 5989 4316
rect 6036 4236 6040 4316
rect 6044 4236 6048 4316
rect 6066 4276 6070 4316
rect 6131 4276 6135 4316
rect 6153 4236 6157 4316
rect 6211 4276 6215 4316
rect 6231 4276 6235 4316
rect 6301 4236 6305 4316
rect 6323 4276 6327 4316
rect 6345 4276 6349 4316
rect 6391 4276 6395 4316
rect 6411 4276 6415 4316
rect 6471 4276 6475 4316
rect 6545 4236 6549 4316
rect 6565 4236 6569 4316
rect 6585 4236 6589 4316
rect 6631 4276 6635 4316
rect 6651 4276 6655 4316
rect 6671 4276 6675 4316
rect 43 3864 47 3944
rect 65 3864 69 3904
rect 111 3864 115 3944
rect 133 3864 137 3884
rect 141 3864 145 3884
rect 161 3864 165 3904
rect 169 3864 173 3904
rect 215 3864 219 3904
rect 235 3864 239 3904
rect 247 3864 251 3904
rect 267 3864 271 3904
rect 281 3864 285 3904
rect 301 3864 305 3944
rect 351 3864 355 3904
rect 371 3864 375 3904
rect 445 3864 449 3944
rect 465 3864 469 3944
rect 485 3864 489 3944
rect 545 3864 549 3904
rect 565 3864 569 3904
rect 625 3864 629 3904
rect 645 3864 649 3904
rect 703 3864 707 3944
rect 725 3864 729 3904
rect 771 3864 775 3944
rect 793 3864 797 3884
rect 801 3864 805 3884
rect 821 3864 825 3904
rect 829 3864 833 3904
rect 875 3864 879 3904
rect 895 3864 899 3904
rect 907 3864 911 3904
rect 927 3864 931 3904
rect 941 3864 945 3904
rect 961 3864 965 3944
rect 1025 3864 1029 3904
rect 1045 3864 1049 3904
rect 1091 3864 1095 3904
rect 1111 3864 1115 3904
rect 1171 3864 1175 3904
rect 1191 3864 1195 3904
rect 1265 3864 1269 3944
rect 1285 3864 1289 3944
rect 1305 3864 1309 3944
rect 1351 3864 1355 3944
rect 1373 3864 1377 3884
rect 1381 3864 1385 3884
rect 1401 3864 1405 3904
rect 1409 3864 1413 3904
rect 1455 3864 1459 3904
rect 1475 3864 1479 3904
rect 1487 3864 1491 3904
rect 1507 3864 1511 3904
rect 1521 3864 1525 3904
rect 1541 3864 1545 3944
rect 1605 3864 1609 3904
rect 1625 3864 1629 3904
rect 1671 3864 1675 3904
rect 1693 3864 1697 3944
rect 1751 3864 1755 3904
rect 1771 3864 1775 3904
rect 1831 3864 1835 3944
rect 1853 3864 1857 3884
rect 1861 3864 1865 3884
rect 1881 3864 1885 3904
rect 1889 3864 1893 3904
rect 1935 3864 1939 3904
rect 1955 3864 1959 3904
rect 1967 3864 1971 3904
rect 1987 3864 1991 3904
rect 2001 3864 2005 3904
rect 2021 3864 2025 3944
rect 2071 3864 2075 3904
rect 2091 3864 2095 3904
rect 2170 3864 2174 3904
rect 2192 3864 2196 3944
rect 2200 3864 2204 3944
rect 2265 3864 2269 3904
rect 2285 3864 2289 3904
rect 2331 3864 2335 3904
rect 2351 3864 2355 3904
rect 2425 3864 2429 3904
rect 2490 3864 2494 3904
rect 2512 3864 2516 3944
rect 2520 3864 2524 3944
rect 2571 3864 2575 3944
rect 2579 3864 2583 3944
rect 2677 3864 2681 3944
rect 2685 3864 2689 3944
rect 2731 3864 2735 3904
rect 2805 3864 2809 3904
rect 2865 3864 2869 3904
rect 2885 3864 2889 3904
rect 2931 3864 2935 3944
rect 2939 3864 2943 3944
rect 3016 3864 3020 3944
rect 3024 3864 3028 3944
rect 3046 3864 3050 3904
rect 3111 3864 3115 3904
rect 3171 3864 3175 3944
rect 3179 3864 3183 3944
rect 3265 3864 3269 3904
rect 3285 3864 3289 3904
rect 3345 3864 3349 3904
rect 3365 3864 3369 3904
rect 3415 3864 3419 3944
rect 3435 3864 3439 3904
rect 3449 3864 3453 3904
rect 3469 3864 3473 3904
rect 3481 3864 3485 3904
rect 3501 3864 3505 3904
rect 3547 3864 3551 3904
rect 3555 3864 3559 3904
rect 3575 3864 3579 3884
rect 3583 3864 3587 3884
rect 3605 3864 3609 3944
rect 3665 3864 3669 3904
rect 3715 3864 3719 3944
rect 3735 3864 3739 3904
rect 3749 3864 3753 3904
rect 3769 3864 3773 3904
rect 3781 3864 3785 3904
rect 3801 3864 3805 3904
rect 3847 3864 3851 3904
rect 3855 3864 3859 3904
rect 3875 3864 3879 3884
rect 3883 3864 3887 3884
rect 3905 3864 3909 3944
rect 3965 3864 3969 3904
rect 3985 3864 3989 3904
rect 4005 3864 4009 3904
rect 4051 3864 4055 3904
rect 4071 3864 4075 3904
rect 4150 3864 4154 3904
rect 4172 3864 4176 3944
rect 4180 3864 4184 3944
rect 4231 3864 4235 3944
rect 4239 3864 4243 3944
rect 4325 3864 4329 3904
rect 4385 3864 4389 3904
rect 4405 3864 4409 3904
rect 4470 3864 4474 3904
rect 4492 3864 4496 3944
rect 4500 3864 4504 3944
rect 4555 3864 4559 3944
rect 4575 3864 4579 3904
rect 4589 3864 4593 3904
rect 4609 3864 4613 3904
rect 4621 3864 4625 3904
rect 4641 3864 4645 3904
rect 4687 3864 4691 3904
rect 4695 3864 4699 3904
rect 4715 3864 4719 3884
rect 4723 3864 4727 3884
rect 4745 3864 4749 3944
rect 4805 3864 4809 3904
rect 4825 3864 4829 3904
rect 4890 3864 4894 3904
rect 4912 3864 4916 3944
rect 4920 3864 4924 3944
rect 4975 3864 4979 3944
rect 4995 3864 4999 3904
rect 5009 3864 5013 3904
rect 5029 3864 5033 3904
rect 5041 3864 5045 3904
rect 5061 3864 5065 3904
rect 5107 3864 5111 3904
rect 5115 3864 5119 3904
rect 5135 3864 5139 3884
rect 5143 3864 5147 3884
rect 5165 3864 5169 3944
rect 5225 3864 5229 3904
rect 5245 3864 5249 3904
rect 5310 3864 5314 3904
rect 5332 3864 5336 3944
rect 5340 3864 5344 3944
rect 5405 3864 5409 3904
rect 5425 3864 5429 3904
rect 5476 3864 5480 3944
rect 5484 3864 5488 3944
rect 5506 3864 5510 3904
rect 5585 3864 5589 3904
rect 5635 3864 5639 3944
rect 5655 3864 5659 3904
rect 5669 3864 5673 3904
rect 5689 3864 5693 3904
rect 5701 3864 5705 3904
rect 5721 3864 5725 3904
rect 5767 3864 5771 3904
rect 5775 3864 5779 3904
rect 5795 3864 5799 3884
rect 5803 3864 5807 3884
rect 5825 3864 5829 3944
rect 5871 3864 5875 3904
rect 5945 3864 5949 3904
rect 5965 3864 5969 3904
rect 5985 3864 5989 3904
rect 6031 3864 6035 3944
rect 6053 3864 6057 3884
rect 6061 3864 6065 3884
rect 6081 3864 6085 3904
rect 6089 3864 6093 3904
rect 6135 3864 6139 3904
rect 6155 3864 6159 3904
rect 6167 3864 6171 3904
rect 6187 3864 6191 3904
rect 6201 3864 6205 3904
rect 6221 3864 6225 3944
rect 6271 3864 6275 3944
rect 6293 3864 6297 3884
rect 6301 3864 6305 3884
rect 6321 3864 6325 3904
rect 6329 3864 6333 3904
rect 6375 3864 6379 3904
rect 6395 3864 6399 3904
rect 6407 3864 6411 3904
rect 6427 3864 6431 3904
rect 6441 3864 6445 3904
rect 6461 3864 6465 3944
rect 6511 3864 6515 3944
rect 6533 3864 6537 3884
rect 6541 3864 6545 3884
rect 6561 3864 6565 3904
rect 6569 3864 6573 3904
rect 6615 3864 6619 3904
rect 6635 3864 6639 3904
rect 6647 3864 6651 3904
rect 6667 3864 6671 3904
rect 6681 3864 6685 3904
rect 6701 3864 6705 3944
rect 43 3756 47 3836
rect 65 3796 69 3836
rect 123 3756 127 3836
rect 145 3796 149 3836
rect 205 3796 209 3836
rect 225 3796 229 3836
rect 271 3756 275 3836
rect 293 3816 297 3836
rect 301 3816 305 3836
rect 321 3796 325 3836
rect 329 3796 333 3836
rect 375 3796 379 3836
rect 395 3796 399 3836
rect 407 3796 411 3836
rect 427 3796 431 3836
rect 441 3796 445 3836
rect 461 3756 465 3836
rect 525 3756 529 3836
rect 545 3756 549 3836
rect 565 3756 569 3836
rect 625 3796 629 3836
rect 645 3796 649 3836
rect 691 3796 695 3836
rect 711 3796 715 3836
rect 785 3796 789 3836
rect 805 3796 809 3836
rect 851 3756 855 3836
rect 873 3816 877 3836
rect 881 3816 885 3836
rect 901 3796 905 3836
rect 909 3796 913 3836
rect 955 3796 959 3836
rect 975 3796 979 3836
rect 987 3796 991 3836
rect 1007 3796 1011 3836
rect 1021 3796 1025 3836
rect 1041 3756 1045 3836
rect 1091 3756 1095 3836
rect 1111 3756 1115 3836
rect 1131 3756 1135 3836
rect 1205 3796 1209 3836
rect 1225 3796 1229 3836
rect 1271 3796 1275 3836
rect 1293 3756 1297 3836
rect 1365 3756 1369 3836
rect 1385 3756 1389 3836
rect 1405 3756 1409 3836
rect 1465 3796 1469 3836
rect 1485 3796 1489 3836
rect 1531 3796 1535 3836
rect 1551 3796 1555 3836
rect 1611 3756 1615 3836
rect 1619 3756 1623 3836
rect 1691 3756 1695 3836
rect 1713 3816 1717 3836
rect 1721 3816 1725 3836
rect 1741 3796 1745 3836
rect 1749 3796 1753 3836
rect 1795 3796 1799 3836
rect 1815 3796 1819 3836
rect 1827 3796 1831 3836
rect 1847 3796 1851 3836
rect 1861 3796 1865 3836
rect 1881 3756 1885 3836
rect 1945 3796 1949 3836
rect 1965 3796 1969 3836
rect 2011 3756 2015 3836
rect 2019 3756 2023 3836
rect 2091 3796 2095 3836
rect 2156 3756 2160 3836
rect 2164 3756 2168 3836
rect 2186 3796 2190 3836
rect 2270 3796 2274 3836
rect 2292 3756 2296 3836
rect 2300 3756 2304 3836
rect 2365 3756 2369 3836
rect 2385 3756 2389 3836
rect 2405 3756 2409 3836
rect 2451 3796 2455 3836
rect 2525 3796 2529 3836
rect 2576 3756 2580 3836
rect 2584 3756 2588 3836
rect 2606 3796 2610 3836
rect 2671 3796 2675 3836
rect 2691 3796 2695 3836
rect 2711 3796 2715 3836
rect 2785 3796 2789 3836
rect 2845 3796 2849 3836
rect 2865 3796 2869 3836
rect 2916 3756 2920 3836
rect 2924 3756 2928 3836
rect 2946 3796 2950 3836
rect 3016 3756 3020 3836
rect 3024 3756 3028 3836
rect 3046 3796 3050 3836
rect 3111 3756 3115 3836
rect 3131 3756 3135 3836
rect 3151 3756 3155 3836
rect 3225 3756 3229 3836
rect 3245 3756 3249 3836
rect 3265 3756 3269 3836
rect 3285 3756 3289 3836
rect 3345 3796 3349 3836
rect 3365 3796 3369 3836
rect 3425 3796 3429 3836
rect 3445 3796 3449 3836
rect 3495 3756 3499 3836
rect 3515 3796 3519 3836
rect 3529 3796 3533 3836
rect 3549 3796 3553 3836
rect 3561 3796 3565 3836
rect 3581 3796 3585 3836
rect 3627 3796 3631 3836
rect 3635 3796 3639 3836
rect 3655 3816 3659 3836
rect 3663 3816 3667 3836
rect 3685 3756 3689 3836
rect 3745 3796 3749 3836
rect 3765 3796 3769 3836
rect 3825 3756 3829 3836
rect 3845 3756 3849 3836
rect 3865 3756 3869 3836
rect 3885 3756 3889 3836
rect 3931 3796 3935 3836
rect 3991 3796 3995 3836
rect 4011 3796 4015 3836
rect 4076 3756 4080 3836
rect 4084 3756 4088 3836
rect 4106 3796 4110 3836
rect 4175 3756 4179 3836
rect 4195 3796 4199 3836
rect 4209 3796 4213 3836
rect 4229 3796 4233 3836
rect 4241 3796 4245 3836
rect 4261 3796 4265 3836
rect 4307 3796 4311 3836
rect 4315 3796 4319 3836
rect 4335 3816 4339 3836
rect 4343 3816 4347 3836
rect 4365 3756 4369 3836
rect 4411 3796 4415 3836
rect 4431 3796 4435 3836
rect 4505 3796 4509 3836
rect 4525 3796 4529 3836
rect 4585 3756 4589 3836
rect 4605 3756 4609 3836
rect 4625 3756 4629 3836
rect 4645 3756 4649 3836
rect 4665 3756 4669 3836
rect 4685 3756 4689 3836
rect 4705 3756 4709 3836
rect 4725 3756 4729 3836
rect 4775 3756 4779 3836
rect 4795 3796 4799 3836
rect 4809 3796 4813 3836
rect 4829 3796 4833 3836
rect 4841 3796 4845 3836
rect 4861 3796 4865 3836
rect 4907 3796 4911 3836
rect 4915 3796 4919 3836
rect 4935 3816 4939 3836
rect 4943 3816 4947 3836
rect 4965 3756 4969 3836
rect 5016 3756 5020 3836
rect 5024 3756 5028 3836
rect 5046 3796 5050 3836
rect 5125 3796 5129 3836
rect 5145 3796 5149 3836
rect 5205 3796 5209 3836
rect 5225 3796 5229 3836
rect 5285 3796 5289 3836
rect 5331 3756 5335 3836
rect 5351 3756 5355 3836
rect 5371 3756 5375 3836
rect 5391 3756 5395 3836
rect 5411 3756 5415 3836
rect 5431 3756 5435 3836
rect 5451 3756 5455 3836
rect 5471 3756 5475 3836
rect 5531 3756 5535 3836
rect 5553 3816 5557 3836
rect 5561 3816 5565 3836
rect 5581 3796 5585 3836
rect 5589 3796 5593 3836
rect 5635 3796 5639 3836
rect 5655 3796 5659 3836
rect 5667 3796 5671 3836
rect 5687 3796 5691 3836
rect 5701 3796 5705 3836
rect 5721 3756 5725 3836
rect 5785 3796 5789 3836
rect 5831 3796 5835 3836
rect 5851 3796 5855 3836
rect 5911 3796 5915 3836
rect 5931 3796 5935 3836
rect 6005 3796 6009 3836
rect 6051 3756 6055 3836
rect 6059 3756 6063 3836
rect 6157 3756 6161 3836
rect 6165 3756 6169 3836
rect 6211 3756 6215 3836
rect 6231 3756 6235 3836
rect 6251 3756 6255 3836
rect 6311 3756 6315 3836
rect 6333 3816 6337 3836
rect 6341 3816 6345 3836
rect 6361 3796 6365 3836
rect 6369 3796 6373 3836
rect 6415 3796 6419 3836
rect 6435 3796 6439 3836
rect 6447 3796 6451 3836
rect 6467 3796 6471 3836
rect 6481 3796 6485 3836
rect 6501 3756 6505 3836
rect 6556 3756 6560 3836
rect 6564 3756 6568 3836
rect 6586 3796 6590 3836
rect 6651 3796 6655 3836
rect 6671 3796 6675 3836
rect 43 3384 47 3464
rect 65 3384 69 3424
rect 111 3384 115 3464
rect 133 3384 137 3404
rect 141 3384 145 3404
rect 161 3384 165 3424
rect 169 3384 173 3424
rect 215 3384 219 3424
rect 235 3384 239 3424
rect 247 3384 251 3424
rect 267 3384 271 3424
rect 281 3384 285 3424
rect 301 3384 305 3464
rect 351 3384 355 3424
rect 371 3384 375 3424
rect 431 3384 435 3424
rect 453 3384 457 3464
rect 525 3384 529 3464
rect 545 3384 549 3464
rect 565 3384 569 3464
rect 625 3384 629 3424
rect 645 3384 649 3424
rect 703 3384 707 3464
rect 725 3384 729 3424
rect 771 3384 775 3424
rect 793 3384 797 3464
rect 851 3384 855 3424
rect 871 3384 875 3424
rect 943 3384 947 3464
rect 965 3384 969 3424
rect 1025 3384 1029 3424
rect 1083 3384 1087 3464
rect 1105 3384 1109 3424
rect 1163 3384 1167 3464
rect 1185 3384 1189 3424
rect 1231 3384 1235 3464
rect 1253 3384 1257 3404
rect 1261 3384 1265 3404
rect 1281 3384 1285 3424
rect 1289 3384 1293 3424
rect 1335 3384 1339 3424
rect 1355 3384 1359 3424
rect 1367 3384 1371 3424
rect 1387 3384 1391 3424
rect 1401 3384 1405 3424
rect 1421 3384 1425 3464
rect 1497 3384 1501 3464
rect 1505 3384 1509 3464
rect 1551 3384 1555 3464
rect 1573 3384 1577 3404
rect 1581 3384 1585 3404
rect 1601 3384 1605 3424
rect 1609 3384 1613 3424
rect 1655 3384 1659 3424
rect 1675 3384 1679 3424
rect 1687 3384 1691 3424
rect 1707 3384 1711 3424
rect 1721 3384 1725 3424
rect 1741 3384 1745 3464
rect 1801 3384 1805 3464
rect 1823 3384 1827 3424
rect 1845 3384 1849 3424
rect 1905 3384 1909 3424
rect 1970 3384 1974 3424
rect 1992 3384 1996 3464
rect 2000 3384 2004 3464
rect 2051 3384 2055 3464
rect 2059 3384 2063 3464
rect 2145 3384 2149 3424
rect 2201 3384 2205 3464
rect 2223 3384 2227 3424
rect 2245 3384 2249 3424
rect 2317 3384 2321 3464
rect 2325 3384 2329 3464
rect 2371 3384 2375 3464
rect 2393 3384 2397 3404
rect 2401 3384 2405 3404
rect 2421 3384 2425 3424
rect 2429 3384 2433 3424
rect 2475 3384 2479 3424
rect 2495 3384 2499 3424
rect 2507 3384 2511 3424
rect 2527 3384 2531 3424
rect 2541 3384 2545 3424
rect 2561 3384 2565 3464
rect 2611 3384 2615 3464
rect 2619 3384 2623 3464
rect 2696 3384 2700 3464
rect 2704 3384 2708 3464
rect 2726 3384 2730 3424
rect 2805 3384 2809 3424
rect 2865 3384 2869 3424
rect 2885 3384 2889 3424
rect 2936 3384 2940 3464
rect 2944 3384 2948 3464
rect 2966 3384 2970 3424
rect 3031 3384 3035 3464
rect 3051 3384 3055 3464
rect 3071 3384 3075 3464
rect 3131 3384 3135 3464
rect 3205 3384 3209 3464
rect 3225 3384 3229 3464
rect 3245 3384 3249 3464
rect 3265 3384 3269 3464
rect 3325 3384 3329 3424
rect 3371 3384 3375 3464
rect 3393 3384 3397 3404
rect 3401 3384 3405 3404
rect 3421 3384 3425 3424
rect 3429 3384 3433 3424
rect 3475 3384 3479 3424
rect 3495 3384 3499 3424
rect 3507 3384 3511 3424
rect 3527 3384 3531 3424
rect 3541 3384 3545 3424
rect 3561 3384 3565 3464
rect 3625 3384 3629 3464
rect 3645 3384 3649 3464
rect 3665 3384 3669 3464
rect 3685 3384 3689 3464
rect 3731 3384 3735 3464
rect 3753 3384 3757 3404
rect 3761 3384 3765 3404
rect 3781 3384 3785 3424
rect 3789 3384 3793 3424
rect 3835 3384 3839 3424
rect 3855 3384 3859 3424
rect 3867 3384 3871 3424
rect 3887 3384 3891 3424
rect 3901 3384 3905 3424
rect 3921 3384 3925 3464
rect 3985 3384 3989 3424
rect 4031 3384 4035 3464
rect 4053 3384 4057 3404
rect 4061 3384 4065 3404
rect 4081 3384 4085 3424
rect 4089 3384 4093 3424
rect 4135 3384 4139 3424
rect 4155 3384 4159 3424
rect 4167 3384 4171 3424
rect 4187 3384 4191 3424
rect 4201 3384 4205 3424
rect 4221 3384 4225 3464
rect 4285 3384 4289 3424
rect 4345 3384 4349 3424
rect 4391 3384 4395 3424
rect 4411 3384 4415 3424
rect 4475 3384 4479 3464
rect 4495 3384 4499 3424
rect 4509 3384 4513 3424
rect 4529 3384 4533 3424
rect 4541 3384 4545 3424
rect 4561 3384 4565 3424
rect 4607 3384 4611 3424
rect 4615 3384 4619 3424
rect 4635 3384 4639 3404
rect 4643 3384 4647 3404
rect 4665 3384 4669 3464
rect 4725 3384 4729 3424
rect 4771 3384 4775 3464
rect 4793 3384 4797 3404
rect 4801 3384 4805 3404
rect 4821 3384 4825 3424
rect 4829 3384 4833 3424
rect 4875 3384 4879 3424
rect 4895 3384 4899 3424
rect 4907 3384 4911 3424
rect 4927 3384 4931 3424
rect 4941 3384 4945 3424
rect 4961 3384 4965 3464
rect 5025 3384 5029 3464
rect 5045 3384 5049 3464
rect 5065 3384 5069 3464
rect 5085 3384 5089 3464
rect 5145 3384 5149 3424
rect 5191 3384 5195 3464
rect 5213 3384 5217 3404
rect 5221 3384 5225 3404
rect 5241 3384 5245 3424
rect 5249 3384 5253 3424
rect 5295 3384 5299 3424
rect 5315 3384 5319 3424
rect 5327 3384 5331 3424
rect 5347 3384 5351 3424
rect 5361 3384 5365 3424
rect 5381 3384 5385 3464
rect 5431 3384 5435 3464
rect 5453 3384 5457 3404
rect 5461 3384 5465 3404
rect 5481 3384 5485 3424
rect 5489 3384 5493 3424
rect 5535 3384 5539 3424
rect 5555 3384 5559 3424
rect 5567 3384 5571 3424
rect 5587 3384 5591 3424
rect 5601 3384 5605 3424
rect 5621 3384 5625 3464
rect 5676 3384 5680 3464
rect 5684 3384 5688 3464
rect 5706 3384 5710 3424
rect 5776 3384 5780 3464
rect 5784 3384 5788 3464
rect 5806 3384 5810 3424
rect 5885 3384 5889 3424
rect 5945 3384 5949 3464
rect 5965 3384 5969 3464
rect 5985 3384 5989 3464
rect 6005 3384 6009 3464
rect 6051 3384 6055 3424
rect 6071 3384 6075 3424
rect 6145 3384 6149 3424
rect 6191 3384 6195 3444
rect 6211 3384 6215 3444
rect 6231 3384 6235 3444
rect 6251 3384 6255 3444
rect 6295 3392 6299 3452
rect 6315 3392 6319 3452
rect 6385 3384 6389 3424
rect 6431 3384 6435 3464
rect 6453 3384 6457 3404
rect 6461 3384 6465 3404
rect 6481 3384 6485 3424
rect 6489 3384 6493 3424
rect 6535 3384 6539 3424
rect 6555 3384 6559 3424
rect 6567 3384 6571 3424
rect 6587 3384 6591 3424
rect 6601 3384 6605 3424
rect 6621 3384 6625 3464
rect 43 3276 47 3356
rect 65 3316 69 3356
rect 111 3276 115 3356
rect 133 3336 137 3356
rect 141 3336 145 3356
rect 161 3316 165 3356
rect 169 3316 173 3356
rect 215 3316 219 3356
rect 235 3316 239 3356
rect 247 3316 251 3356
rect 267 3316 271 3356
rect 281 3316 285 3356
rect 301 3276 305 3356
rect 351 3316 355 3356
rect 371 3316 375 3356
rect 445 3276 449 3356
rect 465 3276 469 3356
rect 485 3276 489 3356
rect 545 3316 549 3356
rect 565 3316 569 3356
rect 611 3316 615 3356
rect 671 3316 675 3356
rect 691 3316 695 3356
rect 711 3316 715 3356
rect 771 3316 775 3356
rect 791 3316 795 3356
rect 870 3316 874 3356
rect 892 3276 896 3356
rect 900 3276 904 3356
rect 951 3316 955 3356
rect 1011 3276 1015 3356
rect 1019 3276 1023 3356
rect 1096 3276 1100 3356
rect 1104 3276 1108 3356
rect 1126 3316 1130 3356
rect 1196 3276 1200 3356
rect 1204 3276 1208 3356
rect 1226 3316 1230 3356
rect 1291 3316 1295 3356
rect 1311 3316 1315 3356
rect 1371 3276 1375 3356
rect 1393 3336 1397 3356
rect 1401 3336 1405 3356
rect 1421 3316 1425 3356
rect 1429 3316 1433 3356
rect 1475 3316 1479 3356
rect 1495 3316 1499 3356
rect 1507 3316 1511 3356
rect 1527 3316 1531 3356
rect 1541 3316 1545 3356
rect 1561 3276 1565 3356
rect 1621 3276 1625 3356
rect 1643 3316 1647 3356
rect 1665 3316 1669 3356
rect 1725 3276 1729 3356
rect 1745 3276 1749 3356
rect 1765 3276 1769 3356
rect 1825 3316 1829 3356
rect 1845 3316 1849 3356
rect 1865 3316 1869 3356
rect 1911 3276 1915 3356
rect 1931 3276 1935 3356
rect 1951 3276 1955 3356
rect 2015 3276 2019 3356
rect 2035 3316 2039 3356
rect 2049 3316 2053 3356
rect 2069 3316 2073 3356
rect 2081 3316 2085 3356
rect 2101 3316 2105 3356
rect 2147 3316 2151 3356
rect 2155 3316 2159 3356
rect 2175 3336 2179 3356
rect 2183 3336 2187 3356
rect 2205 3276 2209 3356
rect 2251 3316 2255 3356
rect 2271 3316 2275 3356
rect 2331 3276 2335 3356
rect 2339 3276 2343 3356
rect 2437 3276 2441 3356
rect 2445 3276 2449 3356
rect 2510 3316 2514 3356
rect 2532 3276 2536 3356
rect 2540 3276 2544 3356
rect 2591 3316 2595 3356
rect 2655 3276 2659 3356
rect 2675 3316 2679 3356
rect 2689 3316 2693 3356
rect 2709 3316 2713 3356
rect 2721 3316 2725 3356
rect 2741 3316 2745 3356
rect 2787 3316 2791 3356
rect 2795 3316 2799 3356
rect 2815 3336 2819 3356
rect 2823 3336 2827 3356
rect 2845 3276 2849 3356
rect 2891 3316 2895 3356
rect 2911 3316 2915 3356
rect 2985 3316 2989 3356
rect 3005 3316 3009 3356
rect 3070 3316 3074 3356
rect 3092 3276 3096 3356
rect 3100 3276 3104 3356
rect 3165 3316 3169 3356
rect 3185 3316 3189 3356
rect 3245 3316 3249 3356
rect 3310 3316 3314 3356
rect 3332 3276 3336 3356
rect 3340 3276 3344 3356
rect 3391 3316 3395 3356
rect 3477 3276 3481 3356
rect 3485 3276 3489 3356
rect 3545 3276 3549 3356
rect 3565 3276 3569 3356
rect 3585 3276 3589 3356
rect 3657 3276 3661 3356
rect 3665 3276 3669 3356
rect 3711 3276 3715 3356
rect 3733 3336 3737 3356
rect 3741 3336 3745 3356
rect 3761 3316 3765 3356
rect 3769 3316 3773 3356
rect 3815 3316 3819 3356
rect 3835 3316 3839 3356
rect 3847 3316 3851 3356
rect 3867 3316 3871 3356
rect 3881 3316 3885 3356
rect 3901 3276 3905 3356
rect 3951 3276 3955 3356
rect 3971 3276 3975 3356
rect 3991 3276 3995 3356
rect 4011 3276 4015 3356
rect 4085 3276 4089 3356
rect 4105 3276 4109 3356
rect 4125 3276 4129 3356
rect 4145 3276 4149 3356
rect 4195 3276 4199 3356
rect 4215 3316 4219 3356
rect 4229 3316 4233 3356
rect 4249 3316 4253 3356
rect 4261 3316 4265 3356
rect 4281 3316 4285 3356
rect 4327 3316 4331 3356
rect 4335 3316 4339 3356
rect 4355 3336 4359 3356
rect 4363 3336 4367 3356
rect 4385 3276 4389 3356
rect 4431 3276 4435 3356
rect 4439 3276 4443 3356
rect 4511 3276 4515 3356
rect 4531 3276 4535 3356
rect 4551 3276 4555 3356
rect 4571 3276 4575 3356
rect 4631 3276 4635 3356
rect 4639 3276 4643 3356
rect 4711 3276 4715 3356
rect 4719 3276 4723 3356
rect 4791 3316 4795 3356
rect 4851 3276 4855 3356
rect 4871 3276 4875 3356
rect 4891 3276 4895 3356
rect 4911 3276 4915 3356
rect 4971 3276 4975 3356
rect 4991 3276 4995 3356
rect 5011 3276 5015 3356
rect 5071 3276 5075 3356
rect 5093 3336 5097 3356
rect 5101 3336 5105 3356
rect 5121 3316 5125 3356
rect 5129 3316 5133 3356
rect 5175 3316 5179 3356
rect 5195 3316 5199 3356
rect 5207 3316 5211 3356
rect 5227 3316 5231 3356
rect 5241 3316 5245 3356
rect 5261 3276 5265 3356
rect 5325 3316 5329 3356
rect 5371 3308 5375 3348
rect 5391 3268 5395 3348
rect 5401 3268 5405 3348
rect 5421 3276 5425 3356
rect 5431 3276 5435 3356
rect 5505 3316 5509 3356
rect 5555 3276 5559 3356
rect 5575 3316 5579 3356
rect 5589 3316 5593 3356
rect 5609 3316 5613 3356
rect 5621 3316 5625 3356
rect 5641 3316 5645 3356
rect 5687 3316 5691 3356
rect 5695 3316 5699 3356
rect 5715 3336 5719 3356
rect 5723 3336 5727 3356
rect 5745 3276 5749 3356
rect 5810 3316 5814 3356
rect 5832 3276 5836 3356
rect 5840 3276 5844 3356
rect 5905 3316 5909 3356
rect 5965 3276 5969 3356
rect 5985 3276 5989 3356
rect 6005 3276 6009 3356
rect 6056 3276 6060 3356
rect 6064 3276 6068 3356
rect 6086 3316 6090 3356
rect 6165 3316 6169 3356
rect 6185 3316 6189 3356
rect 6245 3276 6249 3356
rect 6265 3276 6269 3356
rect 6285 3276 6289 3356
rect 6345 3316 6349 3356
rect 6365 3316 6369 3356
rect 6416 3276 6420 3356
rect 6424 3276 6428 3356
rect 6446 3316 6450 3356
rect 6511 3276 6515 3356
rect 6533 3336 6537 3356
rect 6541 3336 6545 3356
rect 6561 3316 6565 3356
rect 6569 3316 6573 3356
rect 6615 3316 6619 3356
rect 6635 3316 6639 3356
rect 6647 3316 6651 3356
rect 6667 3316 6671 3356
rect 6681 3316 6685 3356
rect 6701 3276 6705 3356
rect 31 2904 35 2984
rect 51 2904 55 2984
rect 71 2904 75 2984
rect 91 2904 95 2984
rect 111 2904 115 2984
rect 131 2904 135 2984
rect 151 2904 155 2984
rect 171 2904 175 2984
rect 243 2904 247 2984
rect 265 2904 269 2944
rect 315 2904 319 2984
rect 335 2904 339 2944
rect 349 2904 353 2944
rect 369 2904 373 2944
rect 381 2904 385 2944
rect 401 2904 405 2944
rect 447 2904 451 2944
rect 455 2904 459 2944
rect 475 2904 479 2924
rect 483 2904 487 2924
rect 505 2904 509 2984
rect 565 2904 569 2944
rect 585 2904 589 2944
rect 631 2904 635 2944
rect 651 2904 655 2944
rect 730 2904 734 2944
rect 752 2904 756 2984
rect 760 2904 764 2984
rect 825 2904 829 2944
rect 845 2904 849 2944
rect 905 2904 909 2944
rect 925 2904 929 2944
rect 971 2904 975 2984
rect 991 2904 995 2984
rect 1011 2904 1015 2984
rect 1071 2904 1075 2984
rect 1093 2904 1097 2924
rect 1101 2904 1105 2924
rect 1121 2904 1125 2944
rect 1129 2904 1133 2944
rect 1175 2904 1179 2944
rect 1195 2904 1199 2944
rect 1207 2904 1211 2944
rect 1227 2904 1231 2944
rect 1241 2904 1245 2944
rect 1261 2904 1265 2984
rect 1325 2904 1329 2944
rect 1345 2904 1349 2944
rect 1391 2904 1395 2984
rect 1413 2904 1417 2924
rect 1421 2904 1425 2924
rect 1441 2904 1445 2944
rect 1449 2904 1453 2944
rect 1495 2904 1499 2944
rect 1515 2904 1519 2944
rect 1527 2904 1531 2944
rect 1547 2904 1551 2944
rect 1561 2904 1565 2944
rect 1581 2904 1585 2984
rect 1645 2904 1649 2944
rect 1710 2904 1714 2944
rect 1732 2904 1736 2984
rect 1740 2904 1744 2984
rect 1817 2904 1821 2984
rect 1825 2904 1829 2984
rect 1881 2904 1885 2984
rect 1903 2904 1907 2944
rect 1925 2904 1929 2944
rect 1976 2904 1980 2984
rect 1984 2904 1988 2984
rect 2006 2904 2010 2944
rect 2085 2904 2089 2984
rect 2105 2904 2109 2984
rect 2125 2904 2129 2984
rect 2171 2904 2175 2944
rect 2191 2904 2195 2944
rect 2265 2904 2269 2944
rect 2311 2904 2315 2944
rect 2333 2904 2337 2944
rect 2355 2904 2359 2984
rect 2415 2904 2419 2984
rect 2435 2904 2439 2944
rect 2449 2904 2453 2944
rect 2469 2904 2473 2944
rect 2481 2904 2485 2944
rect 2501 2904 2505 2944
rect 2547 2904 2551 2944
rect 2555 2904 2559 2944
rect 2575 2904 2579 2924
rect 2583 2904 2587 2924
rect 2605 2904 2609 2984
rect 2651 2904 2655 2944
rect 2711 2904 2715 2984
rect 2719 2904 2723 2984
rect 2805 2904 2809 2944
rect 2870 2904 2874 2944
rect 2892 2904 2896 2984
rect 2900 2904 2904 2984
rect 2951 2904 2955 2984
rect 3025 2904 3029 2944
rect 3045 2904 3049 2944
rect 3065 2904 3069 2944
rect 3125 2904 3129 2944
rect 3145 2904 3149 2944
rect 3210 2904 3214 2944
rect 3232 2904 3236 2984
rect 3240 2904 3244 2984
rect 3291 2904 3295 2944
rect 3311 2904 3315 2944
rect 3371 2904 3375 2944
rect 3391 2904 3395 2944
rect 3456 2904 3460 2984
rect 3464 2904 3468 2984
rect 3486 2904 3490 2944
rect 3551 2904 3555 2944
rect 3573 2904 3577 2944
rect 3595 2904 3599 2984
rect 3665 2904 3669 2984
rect 3685 2904 3689 2984
rect 3705 2904 3709 2984
rect 3725 2904 3729 2984
rect 3785 2904 3789 2984
rect 3805 2904 3809 2984
rect 3855 2904 3859 2984
rect 3875 2904 3879 2944
rect 3889 2904 3893 2944
rect 3909 2904 3913 2944
rect 3921 2904 3925 2944
rect 3941 2904 3945 2944
rect 3987 2904 3991 2944
rect 3995 2904 3999 2944
rect 4015 2904 4019 2924
rect 4023 2904 4027 2924
rect 4045 2904 4049 2984
rect 4096 2904 4100 2984
rect 4104 2904 4108 2984
rect 4126 2904 4130 2944
rect 4205 2904 4209 2944
rect 4225 2904 4229 2944
rect 4245 2904 4249 2944
rect 4295 2904 4299 2984
rect 4315 2904 4319 2944
rect 4329 2904 4333 2944
rect 4349 2904 4353 2944
rect 4361 2904 4365 2944
rect 4381 2904 4385 2944
rect 4427 2904 4431 2944
rect 4435 2904 4439 2944
rect 4455 2904 4459 2924
rect 4463 2904 4467 2924
rect 4485 2904 4489 2984
rect 4555 2904 4559 2984
rect 4565 2904 4569 2984
rect 4595 2904 4599 2984
rect 4605 2904 4609 2984
rect 4665 2904 4669 2944
rect 4725 2904 4729 2984
rect 4735 2904 4739 2984
rect 4755 2912 4759 2992
rect 4765 2912 4769 2992
rect 4785 2912 4789 2952
rect 4831 2904 4835 2984
rect 4851 2904 4855 2984
rect 4871 2904 4875 2984
rect 4891 2904 4895 2984
rect 4965 2904 4969 2944
rect 5011 2904 5015 2984
rect 5031 2904 5035 2984
rect 5051 2904 5055 2984
rect 5071 2904 5075 2984
rect 5131 2904 5135 2944
rect 5191 2904 5195 2984
rect 5199 2904 5203 2984
rect 5275 2904 5279 2984
rect 5295 2904 5299 2944
rect 5309 2904 5313 2944
rect 5329 2904 5333 2944
rect 5341 2904 5345 2944
rect 5361 2904 5365 2944
rect 5407 2904 5411 2944
rect 5415 2904 5419 2944
rect 5435 2904 5439 2924
rect 5443 2904 5447 2924
rect 5465 2904 5469 2984
rect 5537 2904 5541 2984
rect 5545 2904 5549 2984
rect 5596 2904 5600 2984
rect 5604 2904 5608 2984
rect 5626 2904 5630 2944
rect 5705 2904 5709 2944
rect 5725 2904 5729 2944
rect 5745 2904 5749 2944
rect 5815 2904 5819 2984
rect 5825 2904 5829 2984
rect 5855 2904 5859 2984
rect 5865 2904 5869 2984
rect 5911 2904 5915 2944
rect 5971 2912 5975 2952
rect 5991 2912 5995 2992
rect 6001 2912 6005 2992
rect 6021 2904 6025 2984
rect 6031 2904 6035 2984
rect 6105 2904 6109 2984
rect 6125 2904 6129 2984
rect 6145 2904 6149 2984
rect 6217 2904 6221 2984
rect 6225 2904 6229 2984
rect 6271 2904 6275 2944
rect 6345 2904 6349 2984
rect 6365 2904 6369 2984
rect 6385 2904 6389 2984
rect 6405 2904 6409 2984
rect 6465 2904 6469 2944
rect 6511 2904 6515 2944
rect 6576 2904 6580 2984
rect 6584 2904 6588 2984
rect 6606 2904 6610 2944
rect 31 2836 35 2876
rect 117 2796 121 2876
rect 125 2796 129 2876
rect 175 2796 179 2876
rect 195 2836 199 2876
rect 209 2836 213 2876
rect 229 2836 233 2876
rect 241 2836 245 2876
rect 261 2836 265 2876
rect 307 2836 311 2876
rect 315 2836 319 2876
rect 335 2856 339 2876
rect 343 2856 347 2876
rect 365 2796 369 2876
rect 411 2836 415 2876
rect 497 2796 501 2876
rect 505 2796 509 2876
rect 555 2796 559 2876
rect 575 2836 579 2876
rect 589 2836 593 2876
rect 609 2836 613 2876
rect 621 2836 625 2876
rect 641 2836 645 2876
rect 687 2836 691 2876
rect 695 2836 699 2876
rect 715 2856 719 2876
rect 723 2856 727 2876
rect 745 2796 749 2876
rect 803 2796 807 2876
rect 825 2836 829 2876
rect 871 2796 875 2876
rect 891 2796 895 2876
rect 951 2836 955 2876
rect 971 2836 975 2876
rect 1031 2836 1035 2876
rect 1051 2836 1055 2876
rect 1111 2836 1115 2876
rect 1171 2796 1175 2876
rect 1191 2796 1195 2876
rect 1211 2796 1215 2876
rect 1231 2796 1235 2876
rect 1305 2796 1309 2876
rect 1325 2796 1329 2876
rect 1345 2796 1349 2876
rect 1405 2836 1409 2876
rect 1470 2836 1474 2876
rect 1492 2796 1496 2876
rect 1500 2796 1504 2876
rect 1551 2796 1555 2876
rect 1559 2796 1563 2876
rect 1631 2836 1635 2876
rect 1651 2836 1655 2876
rect 1711 2796 1715 2876
rect 1719 2796 1723 2876
rect 1810 2836 1814 2876
rect 1832 2796 1836 2876
rect 1840 2796 1844 2876
rect 1891 2796 1895 2876
rect 1901 2796 1905 2876
rect 1921 2796 1925 2876
rect 1996 2796 2000 2876
rect 2004 2796 2008 2876
rect 2026 2836 2030 2876
rect 2105 2796 2109 2876
rect 2125 2796 2129 2876
rect 2145 2796 2149 2876
rect 2195 2796 2199 2876
rect 2215 2836 2219 2876
rect 2229 2836 2233 2876
rect 2249 2836 2253 2876
rect 2261 2836 2265 2876
rect 2281 2836 2285 2876
rect 2327 2836 2331 2876
rect 2335 2836 2339 2876
rect 2355 2856 2359 2876
rect 2363 2856 2367 2876
rect 2385 2796 2389 2876
rect 2431 2836 2435 2876
rect 2451 2836 2455 2876
rect 2511 2836 2515 2876
rect 2585 2836 2589 2876
rect 2635 2796 2639 2876
rect 2655 2836 2659 2876
rect 2669 2836 2673 2876
rect 2689 2836 2693 2876
rect 2701 2836 2705 2876
rect 2721 2836 2725 2876
rect 2767 2836 2771 2876
rect 2775 2836 2779 2876
rect 2795 2856 2799 2876
rect 2803 2856 2807 2876
rect 2825 2796 2829 2876
rect 2876 2796 2880 2876
rect 2884 2796 2888 2876
rect 2906 2836 2910 2876
rect 2985 2796 2989 2876
rect 3005 2796 3009 2876
rect 3025 2796 3029 2876
rect 3071 2796 3075 2876
rect 3093 2856 3097 2876
rect 3101 2856 3105 2876
rect 3121 2836 3125 2876
rect 3129 2836 3133 2876
rect 3175 2836 3179 2876
rect 3195 2836 3199 2876
rect 3207 2836 3211 2876
rect 3227 2836 3231 2876
rect 3241 2836 3245 2876
rect 3261 2796 3265 2876
rect 3311 2836 3315 2876
rect 3371 2796 3375 2876
rect 3381 2796 3385 2876
rect 3411 2796 3415 2876
rect 3421 2796 3425 2876
rect 3496 2796 3500 2876
rect 3504 2796 3508 2876
rect 3526 2836 3530 2876
rect 3615 2796 3619 2876
rect 3625 2796 3629 2876
rect 3655 2796 3659 2876
rect 3665 2796 3669 2876
rect 3716 2796 3720 2876
rect 3724 2796 3728 2876
rect 3746 2836 3750 2876
rect 3835 2796 3839 2876
rect 3845 2796 3849 2876
rect 3875 2796 3879 2876
rect 3885 2796 3889 2876
rect 3945 2836 3949 2876
rect 3991 2796 3995 2876
rect 3999 2796 4003 2876
rect 4071 2796 4075 2876
rect 4079 2796 4083 2876
rect 4165 2796 4169 2876
rect 4185 2796 4189 2876
rect 4205 2796 4209 2876
rect 4256 2796 4260 2876
rect 4264 2796 4268 2876
rect 4286 2836 4290 2876
rect 4365 2836 4369 2876
rect 4385 2836 4389 2876
rect 4405 2836 4409 2876
rect 4455 2796 4459 2876
rect 4475 2836 4479 2876
rect 4489 2836 4493 2876
rect 4509 2836 4513 2876
rect 4521 2836 4525 2876
rect 4541 2836 4545 2876
rect 4587 2836 4591 2876
rect 4595 2836 4599 2876
rect 4615 2856 4619 2876
rect 4623 2856 4627 2876
rect 4645 2796 4649 2876
rect 4691 2836 4695 2876
rect 4751 2796 4755 2876
rect 4759 2796 4763 2876
rect 4836 2796 4840 2876
rect 4844 2796 4848 2876
rect 4866 2836 4870 2876
rect 4957 2796 4961 2876
rect 4965 2796 4969 2876
rect 5035 2796 5039 2876
rect 5045 2796 5049 2876
rect 5075 2796 5079 2876
rect 5085 2796 5089 2876
rect 5131 2796 5135 2876
rect 5151 2796 5155 2876
rect 5171 2796 5175 2876
rect 5231 2836 5235 2876
rect 5253 2796 5257 2876
rect 5316 2796 5320 2876
rect 5324 2796 5328 2876
rect 5346 2836 5350 2876
rect 5435 2796 5439 2876
rect 5445 2796 5449 2876
rect 5475 2796 5479 2876
rect 5485 2796 5489 2876
rect 5545 2836 5549 2876
rect 5595 2796 5599 2876
rect 5615 2836 5619 2876
rect 5629 2836 5633 2876
rect 5649 2836 5653 2876
rect 5661 2836 5665 2876
rect 5681 2836 5685 2876
rect 5727 2836 5731 2876
rect 5735 2836 5739 2876
rect 5755 2856 5759 2876
rect 5763 2856 5767 2876
rect 5785 2796 5789 2876
rect 5831 2828 5835 2868
rect 5851 2788 5855 2868
rect 5861 2788 5865 2868
rect 5881 2796 5885 2876
rect 5891 2796 5895 2876
rect 5951 2828 5955 2868
rect 5971 2788 5975 2868
rect 5981 2788 5985 2868
rect 6001 2796 6005 2876
rect 6011 2796 6015 2876
rect 6071 2828 6075 2868
rect 6091 2788 6095 2868
rect 6101 2788 6105 2868
rect 6121 2796 6125 2876
rect 6131 2796 6135 2876
rect 6201 2796 6205 2876
rect 6223 2836 6227 2876
rect 6245 2836 6249 2876
rect 6305 2796 6309 2876
rect 6325 2796 6329 2876
rect 6371 2836 6375 2876
rect 6393 2836 6397 2876
rect 6415 2796 6419 2876
rect 6471 2796 6475 2876
rect 6493 2856 6497 2876
rect 6501 2856 6505 2876
rect 6521 2836 6525 2876
rect 6529 2836 6533 2876
rect 6575 2836 6579 2876
rect 6595 2836 6599 2876
rect 6607 2836 6611 2876
rect 6627 2836 6631 2876
rect 6641 2836 6645 2876
rect 6661 2796 6665 2876
rect 31 2424 35 2504
rect 53 2424 57 2444
rect 61 2424 65 2444
rect 81 2424 85 2464
rect 89 2424 93 2464
rect 135 2424 139 2464
rect 155 2424 159 2464
rect 167 2424 171 2464
rect 187 2424 191 2464
rect 201 2424 205 2464
rect 221 2424 225 2504
rect 283 2424 287 2504
rect 305 2424 309 2464
rect 351 2424 355 2504
rect 373 2424 377 2444
rect 381 2424 385 2444
rect 401 2424 405 2464
rect 409 2424 413 2464
rect 455 2424 459 2464
rect 475 2424 479 2464
rect 487 2424 491 2464
rect 507 2424 511 2464
rect 521 2424 525 2464
rect 541 2424 545 2504
rect 605 2424 609 2504
rect 625 2424 629 2504
rect 645 2424 649 2504
rect 691 2424 695 2464
rect 711 2424 715 2464
rect 785 2424 789 2464
rect 805 2424 809 2464
rect 865 2424 869 2504
rect 885 2424 889 2504
rect 905 2424 909 2504
rect 925 2424 929 2504
rect 945 2424 949 2504
rect 965 2424 969 2504
rect 985 2424 989 2504
rect 1005 2424 1009 2504
rect 1051 2424 1055 2504
rect 1073 2424 1077 2444
rect 1081 2424 1085 2444
rect 1101 2424 1105 2464
rect 1109 2424 1113 2464
rect 1155 2424 1159 2464
rect 1175 2424 1179 2464
rect 1187 2424 1191 2464
rect 1207 2424 1211 2464
rect 1221 2424 1225 2464
rect 1241 2424 1245 2504
rect 1305 2424 1309 2464
rect 1325 2424 1329 2464
rect 1371 2424 1375 2504
rect 1379 2424 1383 2504
rect 1451 2424 1455 2464
rect 1530 2424 1534 2464
rect 1552 2424 1556 2504
rect 1560 2424 1564 2504
rect 1615 2424 1619 2504
rect 1635 2424 1639 2464
rect 1649 2424 1653 2464
rect 1669 2424 1673 2464
rect 1681 2424 1685 2464
rect 1701 2424 1705 2464
rect 1747 2424 1751 2464
rect 1755 2424 1759 2464
rect 1775 2424 1779 2444
rect 1783 2424 1787 2444
rect 1805 2424 1809 2504
rect 1851 2424 1855 2464
rect 1911 2424 1915 2464
rect 1971 2424 1975 2504
rect 1981 2424 1985 2504
rect 2011 2424 2015 2504
rect 2021 2424 2025 2504
rect 2091 2424 2095 2504
rect 2099 2424 2103 2504
rect 2171 2432 2175 2472
rect 2191 2432 2195 2512
rect 2201 2432 2205 2512
rect 2221 2424 2225 2504
rect 2231 2424 2235 2504
rect 2291 2432 2295 2472
rect 2311 2432 2315 2512
rect 2321 2432 2325 2512
rect 2341 2424 2345 2504
rect 2351 2424 2355 2504
rect 2415 2424 2419 2504
rect 2435 2424 2439 2464
rect 2449 2424 2453 2464
rect 2469 2424 2473 2464
rect 2481 2424 2485 2464
rect 2501 2424 2505 2464
rect 2547 2424 2551 2464
rect 2555 2424 2559 2464
rect 2575 2424 2579 2444
rect 2583 2424 2587 2444
rect 2605 2424 2609 2504
rect 2651 2432 2655 2472
rect 2671 2432 2675 2512
rect 2681 2432 2685 2512
rect 2701 2424 2705 2504
rect 2711 2424 2715 2504
rect 2797 2424 2801 2504
rect 2805 2424 2809 2504
rect 2865 2424 2869 2504
rect 2875 2424 2879 2504
rect 2895 2432 2899 2512
rect 2905 2432 2909 2512
rect 2925 2432 2929 2472
rect 2995 2424 2999 2504
rect 3005 2424 3009 2504
rect 3035 2424 3039 2504
rect 3045 2424 3049 2504
rect 3105 2424 3109 2464
rect 3155 2424 3159 2504
rect 3175 2424 3179 2464
rect 3189 2424 3193 2464
rect 3209 2424 3213 2464
rect 3221 2424 3225 2464
rect 3241 2424 3245 2464
rect 3287 2424 3291 2464
rect 3295 2424 3299 2464
rect 3315 2424 3319 2444
rect 3323 2424 3327 2444
rect 3345 2424 3349 2504
rect 3391 2424 3395 2504
rect 3399 2424 3403 2504
rect 3485 2424 3489 2464
rect 3505 2424 3509 2464
rect 3551 2424 3555 2464
rect 3611 2424 3615 2464
rect 3631 2424 3635 2464
rect 3651 2424 3655 2464
rect 3711 2424 3715 2464
rect 3731 2424 3735 2464
rect 3751 2424 3755 2464
rect 3825 2424 3829 2464
rect 3845 2424 3849 2464
rect 3865 2424 3869 2464
rect 3916 2424 3920 2504
rect 3924 2424 3928 2504
rect 3946 2424 3950 2464
rect 4011 2424 4015 2504
rect 4031 2424 4035 2504
rect 4051 2424 4055 2504
rect 4137 2424 4141 2504
rect 4145 2424 4149 2504
rect 4215 2424 4219 2504
rect 4225 2424 4229 2504
rect 4255 2424 4259 2504
rect 4265 2424 4269 2504
rect 4315 2424 4319 2504
rect 4335 2424 4339 2464
rect 4349 2424 4353 2464
rect 4369 2424 4373 2464
rect 4381 2424 4385 2464
rect 4401 2424 4405 2464
rect 4447 2424 4451 2464
rect 4455 2424 4459 2464
rect 4475 2424 4479 2444
rect 4483 2424 4487 2444
rect 4505 2424 4509 2504
rect 4565 2424 4569 2464
rect 4635 2424 4639 2504
rect 4645 2424 4649 2504
rect 4675 2424 4679 2504
rect 4685 2424 4689 2504
rect 4731 2432 4735 2472
rect 4751 2432 4755 2512
rect 4761 2432 4765 2512
rect 4781 2424 4785 2504
rect 4791 2424 4795 2504
rect 4851 2424 4855 2504
rect 4873 2424 4877 2444
rect 4881 2424 4885 2444
rect 4901 2424 4905 2464
rect 4909 2424 4913 2464
rect 4955 2424 4959 2464
rect 4975 2424 4979 2464
rect 4987 2424 4991 2464
rect 5007 2424 5011 2464
rect 5021 2424 5025 2464
rect 5041 2424 5045 2504
rect 5091 2424 5095 2464
rect 5151 2424 5155 2504
rect 5161 2424 5165 2504
rect 5191 2424 5195 2504
rect 5201 2424 5205 2504
rect 5276 2424 5280 2504
rect 5284 2424 5288 2504
rect 5306 2424 5310 2464
rect 5371 2424 5375 2504
rect 5379 2424 5383 2504
rect 5477 2424 5481 2504
rect 5485 2424 5489 2504
rect 5531 2424 5535 2504
rect 5551 2424 5555 2504
rect 5571 2424 5575 2504
rect 5591 2424 5595 2504
rect 5611 2424 5615 2504
rect 5631 2424 5635 2504
rect 5651 2424 5655 2504
rect 5671 2424 5675 2504
rect 5757 2424 5761 2504
rect 5765 2424 5769 2504
rect 5816 2424 5820 2504
rect 5824 2424 5828 2504
rect 5846 2424 5850 2464
rect 5935 2424 5939 2504
rect 5945 2424 5949 2504
rect 5975 2424 5979 2504
rect 5985 2424 5989 2504
rect 6045 2424 6049 2464
rect 6091 2424 6095 2504
rect 6113 2424 6117 2444
rect 6121 2424 6125 2444
rect 6141 2424 6145 2464
rect 6149 2424 6153 2464
rect 6195 2424 6199 2464
rect 6215 2424 6219 2464
rect 6227 2424 6231 2464
rect 6247 2424 6251 2464
rect 6261 2424 6265 2464
rect 6281 2424 6285 2504
rect 6345 2424 6349 2504
rect 6365 2424 6369 2504
rect 6385 2424 6389 2504
rect 6405 2424 6409 2504
rect 6451 2424 6455 2504
rect 6471 2424 6475 2504
rect 6531 2424 6535 2464
rect 6591 2424 6595 2504
rect 6611 2424 6615 2504
rect 6631 2424 6635 2504
rect 6651 2424 6655 2504
rect 35 2316 39 2396
rect 55 2356 59 2396
rect 69 2356 73 2396
rect 89 2356 93 2396
rect 101 2356 105 2396
rect 121 2356 125 2396
rect 167 2356 171 2396
rect 175 2356 179 2396
rect 195 2376 199 2396
rect 203 2376 207 2396
rect 225 2316 229 2396
rect 283 2316 287 2396
rect 305 2356 309 2396
rect 365 2316 369 2396
rect 425 2356 429 2396
rect 497 2316 501 2396
rect 505 2316 509 2396
rect 556 2316 560 2396
rect 564 2316 568 2396
rect 586 2356 590 2396
rect 661 2316 665 2396
rect 683 2356 687 2396
rect 705 2356 709 2396
rect 751 2356 755 2396
rect 771 2356 775 2396
rect 791 2356 795 2396
rect 851 2356 855 2396
rect 871 2356 875 2396
rect 931 2316 935 2396
rect 953 2376 957 2396
rect 961 2376 965 2396
rect 981 2356 985 2396
rect 989 2356 993 2396
rect 1035 2356 1039 2396
rect 1055 2356 1059 2396
rect 1067 2356 1071 2396
rect 1087 2356 1091 2396
rect 1101 2356 1105 2396
rect 1121 2316 1125 2396
rect 1171 2356 1175 2396
rect 1235 2316 1239 2396
rect 1255 2356 1259 2396
rect 1269 2356 1273 2396
rect 1289 2356 1293 2396
rect 1301 2356 1305 2396
rect 1321 2356 1325 2396
rect 1367 2356 1371 2396
rect 1375 2356 1379 2396
rect 1395 2376 1399 2396
rect 1403 2376 1407 2396
rect 1425 2316 1429 2396
rect 1485 2356 1489 2396
rect 1531 2316 1535 2396
rect 1541 2316 1545 2396
rect 1571 2316 1575 2396
rect 1581 2316 1585 2396
rect 1656 2316 1660 2396
rect 1664 2316 1668 2396
rect 1686 2356 1690 2396
rect 1777 2316 1781 2396
rect 1785 2316 1789 2396
rect 1857 2316 1861 2396
rect 1865 2316 1869 2396
rect 1935 2316 1939 2396
rect 1945 2316 1949 2396
rect 1975 2316 1979 2396
rect 1985 2316 1989 2396
rect 2045 2356 2049 2396
rect 2095 2316 2099 2396
rect 2115 2356 2119 2396
rect 2129 2356 2133 2396
rect 2149 2356 2153 2396
rect 2161 2356 2165 2396
rect 2181 2356 2185 2396
rect 2227 2356 2231 2396
rect 2235 2356 2239 2396
rect 2255 2376 2259 2396
rect 2263 2376 2267 2396
rect 2285 2316 2289 2396
rect 2357 2316 2361 2396
rect 2365 2316 2369 2396
rect 2416 2316 2420 2396
rect 2424 2316 2428 2396
rect 2446 2356 2450 2396
rect 2525 2356 2529 2396
rect 2545 2356 2549 2396
rect 2565 2356 2569 2396
rect 2625 2316 2629 2396
rect 2645 2316 2649 2396
rect 2665 2316 2669 2396
rect 2716 2316 2720 2396
rect 2724 2316 2728 2396
rect 2746 2356 2750 2396
rect 2837 2316 2841 2396
rect 2845 2316 2849 2396
rect 2891 2316 2895 2396
rect 2913 2376 2917 2396
rect 2921 2376 2925 2396
rect 2941 2356 2945 2396
rect 2949 2356 2953 2396
rect 2995 2356 2999 2396
rect 3015 2356 3019 2396
rect 3027 2356 3031 2396
rect 3047 2356 3051 2396
rect 3061 2356 3065 2396
rect 3081 2316 3085 2396
rect 3136 2316 3140 2396
rect 3144 2316 3148 2396
rect 3166 2356 3170 2396
rect 3255 2316 3259 2396
rect 3265 2316 3269 2396
rect 3295 2316 3299 2396
rect 3305 2316 3309 2396
rect 3377 2316 3381 2396
rect 3385 2316 3389 2396
rect 3445 2356 3449 2396
rect 3517 2316 3521 2396
rect 3525 2316 3529 2396
rect 3575 2316 3579 2396
rect 3595 2356 3599 2396
rect 3609 2356 3613 2396
rect 3629 2356 3633 2396
rect 3641 2356 3645 2396
rect 3661 2356 3665 2396
rect 3707 2356 3711 2396
rect 3715 2356 3719 2396
rect 3735 2376 3739 2396
rect 3743 2376 3747 2396
rect 3765 2316 3769 2396
rect 3811 2356 3815 2396
rect 3831 2356 3835 2396
rect 3891 2356 3895 2396
rect 3911 2356 3915 2396
rect 3931 2356 3935 2396
rect 3991 2348 3995 2388
rect 4011 2308 4015 2388
rect 4021 2308 4025 2388
rect 4041 2316 4045 2396
rect 4051 2316 4055 2396
rect 4111 2348 4115 2388
rect 4131 2308 4135 2388
rect 4141 2308 4145 2388
rect 4161 2316 4165 2396
rect 4171 2316 4175 2396
rect 4231 2348 4235 2388
rect 4251 2308 4255 2388
rect 4261 2308 4265 2388
rect 4281 2316 4285 2396
rect 4291 2316 4295 2396
rect 4351 2356 4355 2396
rect 4373 2316 4377 2396
rect 4457 2316 4461 2396
rect 4465 2316 4469 2396
rect 4511 2348 4515 2388
rect 4531 2308 4535 2388
rect 4541 2308 4545 2388
rect 4561 2316 4565 2396
rect 4571 2316 4575 2396
rect 4645 2316 4649 2396
rect 4655 2316 4659 2396
rect 4675 2308 4679 2388
rect 4685 2308 4689 2388
rect 4705 2348 4709 2388
rect 4751 2348 4755 2388
rect 4771 2308 4775 2388
rect 4781 2308 4785 2388
rect 4801 2316 4805 2396
rect 4811 2316 4815 2396
rect 4871 2316 4875 2396
rect 4879 2316 4883 2396
rect 4951 2348 4955 2388
rect 4971 2308 4975 2388
rect 4981 2308 4985 2388
rect 5001 2316 5005 2396
rect 5011 2316 5015 2396
rect 5085 2316 5089 2396
rect 5105 2316 5109 2396
rect 5125 2316 5129 2396
rect 5171 2356 5175 2396
rect 5231 2316 5235 2396
rect 5241 2316 5245 2396
rect 5271 2316 5275 2396
rect 5281 2316 5285 2396
rect 5365 2316 5369 2396
rect 5375 2316 5379 2396
rect 5395 2308 5399 2388
rect 5405 2308 5409 2388
rect 5425 2348 5429 2388
rect 5471 2348 5475 2388
rect 5491 2308 5495 2388
rect 5501 2308 5505 2388
rect 5521 2316 5525 2396
rect 5531 2316 5535 2396
rect 5591 2348 5595 2388
rect 5611 2308 5615 2388
rect 5621 2308 5625 2388
rect 5641 2316 5645 2396
rect 5651 2316 5655 2396
rect 5725 2356 5729 2396
rect 5745 2356 5749 2396
rect 5765 2356 5769 2396
rect 5825 2356 5829 2396
rect 5845 2356 5849 2396
rect 5865 2356 5869 2396
rect 5925 2356 5929 2396
rect 5985 2316 5989 2396
rect 6005 2316 6009 2396
rect 6025 2316 6029 2396
rect 6045 2316 6049 2396
rect 6105 2316 6109 2396
rect 6115 2316 6119 2396
rect 6135 2308 6139 2388
rect 6145 2308 6149 2388
rect 6165 2348 6169 2388
rect 6225 2316 6229 2396
rect 6235 2316 6239 2396
rect 6255 2308 6259 2388
rect 6265 2308 6269 2388
rect 6285 2348 6289 2388
rect 6331 2356 6335 2396
rect 6396 2316 6400 2396
rect 6404 2316 6408 2396
rect 6426 2356 6430 2396
rect 6491 2356 6495 2396
rect 6511 2356 6515 2396
rect 6571 2316 6575 2396
rect 6591 2316 6595 2396
rect 6611 2316 6615 2396
rect 6671 2356 6675 2396
rect 57 1944 61 2024
rect 65 1944 69 2024
rect 125 1944 129 1984
rect 145 1944 149 1984
rect 205 1944 209 1984
rect 225 1944 229 1984
rect 245 1944 249 1984
rect 305 1944 309 1984
rect 325 1944 329 1984
rect 345 1944 349 1984
rect 405 1944 409 1984
rect 425 1944 429 1984
rect 471 1944 475 1984
rect 491 1944 495 1984
rect 511 1944 515 1984
rect 597 1944 601 2024
rect 605 1944 609 2024
rect 656 1944 660 2024
rect 664 1944 668 2024
rect 686 1944 690 1984
rect 751 1944 755 1984
rect 771 1944 775 1984
rect 791 1944 795 1984
rect 851 1944 855 2024
rect 859 1944 863 2024
rect 945 1944 949 1984
rect 965 1944 969 1984
rect 1011 1952 1015 1992
rect 1031 1952 1035 2032
rect 1041 1952 1045 2032
rect 1061 1944 1065 2024
rect 1071 1944 1075 2024
rect 1135 1944 1139 2024
rect 1155 1944 1159 1984
rect 1169 1944 1173 1984
rect 1189 1944 1193 1984
rect 1201 1944 1205 1984
rect 1221 1944 1225 1984
rect 1267 1944 1271 1984
rect 1275 1944 1279 1984
rect 1295 1944 1299 1964
rect 1303 1944 1307 1964
rect 1325 1944 1329 2024
rect 1371 1944 1375 1984
rect 1431 1944 1435 2024
rect 1441 1944 1445 2024
rect 1471 1944 1475 2024
rect 1481 1944 1485 2024
rect 1570 1944 1574 1984
rect 1592 1944 1596 2024
rect 1600 1944 1604 2024
rect 1670 1944 1674 1984
rect 1692 1944 1696 2024
rect 1700 1944 1704 2024
rect 1777 1944 1781 2024
rect 1785 1944 1789 2024
rect 1850 1944 1854 1984
rect 1872 1944 1876 2024
rect 1880 1944 1884 2024
rect 1945 1944 1949 2024
rect 1955 1944 1959 2024
rect 1975 1952 1979 2032
rect 1985 1952 1989 2032
rect 2005 1952 2009 1992
rect 2065 1944 2069 2024
rect 2075 1944 2079 2024
rect 2095 1952 2099 2032
rect 2105 1952 2109 2032
rect 2125 1952 2129 1992
rect 2175 1944 2179 2024
rect 2195 1944 2199 1984
rect 2209 1944 2213 1984
rect 2229 1944 2233 1984
rect 2241 1944 2245 1984
rect 2261 1944 2265 1984
rect 2307 1944 2311 1984
rect 2315 1944 2319 1984
rect 2335 1944 2339 1964
rect 2343 1944 2347 1964
rect 2365 1944 2369 2024
rect 2430 1944 2434 1984
rect 2452 1944 2456 2024
rect 2460 1944 2464 2024
rect 2511 1944 2515 2024
rect 2519 1944 2523 2024
rect 2605 1944 2609 1984
rect 2625 1944 2629 1984
rect 2645 1944 2649 1984
rect 2691 1952 2695 1992
rect 2711 1952 2715 2032
rect 2721 1952 2725 2032
rect 2741 1944 2745 2024
rect 2751 1944 2755 2024
rect 2825 1944 2829 2024
rect 2835 1944 2839 2024
rect 2855 1952 2859 2032
rect 2865 1952 2869 2032
rect 2885 1952 2889 1992
rect 2931 1944 2935 1984
rect 2991 1944 2995 2024
rect 3001 1944 3005 2024
rect 3031 1944 3035 2024
rect 3041 1944 3045 2024
rect 3125 1944 3129 2024
rect 3145 1944 3149 2024
rect 3165 1944 3169 2024
rect 3211 1944 3215 1984
rect 3271 1944 3275 2024
rect 3281 1944 3285 2024
rect 3311 1944 3315 2024
rect 3321 1944 3325 2024
rect 3391 1944 3395 2024
rect 3399 1944 3403 2024
rect 3475 1944 3479 2024
rect 3495 1944 3499 1984
rect 3509 1944 3513 1984
rect 3529 1944 3533 1984
rect 3541 1944 3545 1984
rect 3561 1944 3565 1984
rect 3607 1944 3611 1984
rect 3615 1944 3619 1984
rect 3635 1944 3639 1964
rect 3643 1944 3647 1964
rect 3665 1944 3669 2024
rect 3737 1944 3741 2024
rect 3745 1944 3749 2024
rect 3815 1944 3819 2024
rect 3825 1944 3829 2024
rect 3855 1944 3859 2024
rect 3865 1944 3869 2024
rect 3925 1944 3929 1984
rect 3976 1944 3980 2024
rect 3984 1944 3988 2024
rect 4006 1944 4010 1984
rect 4071 1944 4075 1984
rect 4091 1944 4095 1984
rect 4177 1944 4181 2024
rect 4185 1944 4189 2024
rect 4235 1944 4239 2024
rect 4255 1944 4259 1984
rect 4269 1944 4273 1984
rect 4289 1944 4293 1984
rect 4301 1944 4305 1984
rect 4321 1944 4325 1984
rect 4367 1944 4371 1984
rect 4375 1944 4379 1984
rect 4395 1944 4399 1964
rect 4403 1944 4407 1964
rect 4425 1944 4429 2024
rect 4471 1944 4475 1984
rect 4531 1944 4535 2024
rect 4541 1944 4545 2024
rect 4571 1944 4575 2024
rect 4581 1944 4585 2024
rect 4651 1944 4655 2024
rect 4659 1944 4663 2024
rect 4750 1944 4754 1984
rect 4772 1944 4776 2024
rect 4780 1944 4784 2024
rect 4857 1944 4861 2024
rect 4865 1944 4869 2024
rect 4911 1944 4915 2024
rect 4921 1944 4925 2024
rect 4951 1944 4955 2024
rect 4961 1944 4965 2024
rect 5045 1944 5049 1984
rect 5065 1944 5069 1984
rect 5137 1944 5141 2024
rect 5145 1944 5149 2024
rect 5191 1944 5195 2024
rect 5201 1944 5205 2024
rect 5221 1944 5225 2024
rect 5315 1944 5319 2024
rect 5325 1944 5329 2024
rect 5355 1944 5359 2024
rect 5365 1944 5369 2024
rect 5411 1944 5415 2024
rect 5421 1944 5425 2024
rect 5451 1944 5455 2024
rect 5461 1944 5465 2024
rect 5557 1944 5561 2024
rect 5565 1944 5569 2024
rect 5635 1944 5639 2024
rect 5645 1944 5649 2024
rect 5675 1944 5679 2024
rect 5685 1944 5689 2024
rect 5745 1944 5749 1984
rect 5791 1944 5795 1984
rect 5811 1944 5815 1984
rect 5871 1944 5875 2024
rect 5893 1944 5897 1964
rect 5901 1944 5905 1964
rect 5921 1944 5925 1984
rect 5929 1944 5933 1984
rect 5975 1944 5979 1984
rect 5995 1944 5999 1984
rect 6007 1944 6011 1984
rect 6027 1944 6031 1984
rect 6041 1944 6045 1984
rect 6061 1944 6065 2024
rect 6115 1944 6119 2024
rect 6135 1944 6139 1984
rect 6149 1944 6153 1984
rect 6169 1944 6173 1984
rect 6181 1944 6185 1984
rect 6201 1944 6205 1984
rect 6247 1944 6251 1984
rect 6255 1944 6259 1984
rect 6275 1944 6279 1964
rect 6283 1944 6287 1964
rect 6305 1944 6309 2024
rect 6351 1952 6355 1992
rect 6371 1952 6375 2032
rect 6381 1952 6385 2032
rect 6401 1944 6405 2024
rect 6411 1944 6415 2024
rect 6471 1944 6475 2024
rect 6491 1944 6495 2024
rect 6511 1944 6515 2024
rect 6576 1944 6580 2024
rect 6584 1944 6588 2024
rect 6606 1944 6610 1984
rect 45 1876 49 1916
rect 91 1836 95 1916
rect 113 1896 117 1916
rect 121 1896 125 1916
rect 141 1876 145 1916
rect 149 1876 153 1916
rect 195 1876 199 1916
rect 215 1876 219 1916
rect 227 1876 231 1916
rect 247 1876 251 1916
rect 261 1876 265 1916
rect 281 1836 285 1916
rect 331 1836 335 1916
rect 339 1836 343 1916
rect 437 1836 441 1916
rect 445 1836 449 1916
rect 505 1876 509 1916
rect 570 1876 574 1916
rect 592 1836 596 1916
rect 600 1836 604 1916
rect 651 1836 655 1916
rect 673 1896 677 1916
rect 681 1896 685 1916
rect 701 1876 705 1916
rect 709 1876 713 1916
rect 755 1876 759 1916
rect 775 1876 779 1916
rect 787 1876 791 1916
rect 807 1876 811 1916
rect 821 1876 825 1916
rect 841 1836 845 1916
rect 905 1876 909 1916
rect 925 1876 929 1916
rect 945 1876 949 1916
rect 991 1876 995 1916
rect 1013 1876 1017 1916
rect 1035 1836 1039 1916
rect 1091 1876 1095 1916
rect 1156 1836 1160 1916
rect 1164 1836 1168 1916
rect 1186 1876 1190 1916
rect 1265 1876 1269 1916
rect 1285 1876 1289 1916
rect 1345 1876 1349 1916
rect 1365 1876 1369 1916
rect 1385 1876 1389 1916
rect 1431 1876 1435 1916
rect 1495 1836 1499 1916
rect 1515 1876 1519 1916
rect 1529 1876 1533 1916
rect 1549 1876 1553 1916
rect 1561 1876 1565 1916
rect 1581 1876 1585 1916
rect 1627 1876 1631 1916
rect 1635 1876 1639 1916
rect 1655 1896 1659 1916
rect 1663 1896 1667 1916
rect 1685 1836 1689 1916
rect 1731 1876 1735 1916
rect 1791 1836 1795 1916
rect 1801 1836 1805 1916
rect 1831 1836 1835 1916
rect 1841 1836 1845 1916
rect 1911 1836 1915 1916
rect 1919 1836 1923 1916
rect 1996 1836 2000 1916
rect 2004 1836 2008 1916
rect 2026 1876 2030 1916
rect 2091 1836 2095 1916
rect 2113 1896 2117 1916
rect 2121 1896 2125 1916
rect 2141 1876 2145 1916
rect 2149 1876 2153 1916
rect 2195 1876 2199 1916
rect 2215 1876 2219 1916
rect 2227 1876 2231 1916
rect 2247 1876 2251 1916
rect 2261 1876 2265 1916
rect 2281 1836 2285 1916
rect 2355 1836 2359 1916
rect 2365 1836 2369 1916
rect 2395 1836 2399 1916
rect 2405 1836 2409 1916
rect 2451 1876 2455 1916
rect 2511 1836 2515 1916
rect 2519 1836 2523 1916
rect 2591 1836 2595 1916
rect 2613 1896 2617 1916
rect 2621 1896 2625 1916
rect 2641 1876 2645 1916
rect 2649 1876 2653 1916
rect 2695 1876 2699 1916
rect 2715 1876 2719 1916
rect 2727 1876 2731 1916
rect 2747 1876 2751 1916
rect 2761 1876 2765 1916
rect 2781 1836 2785 1916
rect 2831 1876 2835 1916
rect 2851 1876 2855 1916
rect 2871 1876 2875 1916
rect 2950 1876 2954 1916
rect 2972 1836 2976 1916
rect 2980 1836 2984 1916
rect 3031 1836 3035 1916
rect 3039 1836 3043 1916
rect 3125 1836 3129 1916
rect 3145 1836 3149 1916
rect 3165 1836 3169 1916
rect 3225 1836 3229 1916
rect 3245 1836 3249 1916
rect 3265 1836 3269 1916
rect 3323 1836 3327 1916
rect 3345 1876 3349 1916
rect 3405 1876 3409 1916
rect 3425 1876 3429 1916
rect 3471 1836 3475 1916
rect 3479 1836 3483 1916
rect 3551 1876 3555 1916
rect 3571 1876 3575 1916
rect 3636 1836 3640 1916
rect 3644 1836 3648 1916
rect 3666 1876 3670 1916
rect 3745 1876 3749 1916
rect 3765 1876 3769 1916
rect 3825 1876 3829 1916
rect 3871 1876 3875 1916
rect 3891 1876 3895 1916
rect 3951 1836 3955 1916
rect 3959 1836 3963 1916
rect 4031 1836 4035 1916
rect 4041 1836 4045 1916
rect 4071 1836 4075 1916
rect 4081 1836 4085 1916
rect 4177 1836 4181 1916
rect 4185 1836 4189 1916
rect 4236 1836 4240 1916
rect 4244 1836 4248 1916
rect 4266 1876 4270 1916
rect 4331 1836 4335 1916
rect 4351 1836 4355 1916
rect 4416 1836 4420 1916
rect 4424 1836 4428 1916
rect 4446 1876 4450 1916
rect 4537 1836 4541 1916
rect 4545 1836 4549 1916
rect 4615 1836 4619 1916
rect 4625 1836 4629 1916
rect 4655 1836 4659 1916
rect 4665 1836 4669 1916
rect 4725 1876 4729 1916
rect 4771 1836 4775 1916
rect 4793 1896 4797 1916
rect 4801 1896 4805 1916
rect 4821 1876 4825 1916
rect 4829 1876 4833 1916
rect 4875 1876 4879 1916
rect 4895 1876 4899 1916
rect 4907 1876 4911 1916
rect 4927 1876 4931 1916
rect 4941 1876 4945 1916
rect 4961 1836 4965 1916
rect 5011 1836 5015 1916
rect 5031 1836 5035 1916
rect 5051 1836 5055 1916
rect 5111 1836 5115 1916
rect 5119 1836 5123 1916
rect 5196 1836 5200 1916
rect 5204 1836 5208 1916
rect 5226 1876 5230 1916
rect 5291 1876 5295 1916
rect 5311 1876 5315 1916
rect 5331 1876 5335 1916
rect 5391 1876 5395 1916
rect 5413 1836 5417 1916
rect 5485 1876 5489 1916
rect 5545 1836 5549 1916
rect 5610 1876 5614 1916
rect 5632 1836 5636 1916
rect 5640 1836 5644 1916
rect 5691 1876 5695 1916
rect 5711 1876 5715 1916
rect 5785 1836 5789 1916
rect 5805 1836 5809 1916
rect 5825 1836 5829 1916
rect 5845 1836 5849 1916
rect 5891 1876 5895 1916
rect 5913 1836 5917 1916
rect 5990 1876 5994 1916
rect 6012 1836 6016 1916
rect 6020 1836 6024 1916
rect 6095 1836 6099 1916
rect 6105 1836 6109 1916
rect 6135 1836 6139 1916
rect 6145 1836 6149 1916
rect 6191 1868 6195 1908
rect 6211 1828 6215 1908
rect 6221 1828 6225 1908
rect 6241 1836 6245 1916
rect 6251 1836 6255 1916
rect 6311 1868 6315 1908
rect 6331 1828 6335 1908
rect 6341 1828 6345 1908
rect 6361 1836 6365 1916
rect 6371 1836 6375 1916
rect 6431 1876 6435 1916
rect 6496 1836 6500 1916
rect 6504 1836 6508 1916
rect 6526 1876 6530 1916
rect 6605 1876 6609 1916
rect 6625 1876 6629 1916
rect 57 1464 61 1544
rect 65 1464 69 1544
rect 125 1464 129 1544
rect 145 1464 149 1544
rect 165 1464 169 1544
rect 185 1464 189 1544
rect 205 1464 209 1544
rect 225 1464 229 1544
rect 245 1464 249 1544
rect 265 1464 269 1544
rect 315 1464 319 1544
rect 335 1464 339 1504
rect 349 1464 353 1504
rect 369 1464 373 1504
rect 381 1464 385 1504
rect 401 1464 405 1504
rect 447 1464 451 1504
rect 455 1464 459 1504
rect 475 1464 479 1484
rect 483 1464 487 1484
rect 505 1464 509 1544
rect 565 1464 569 1504
rect 611 1464 615 1504
rect 631 1464 635 1504
rect 651 1464 655 1504
rect 711 1464 715 1544
rect 731 1464 735 1544
rect 751 1464 755 1544
rect 815 1464 819 1544
rect 835 1464 839 1504
rect 849 1464 853 1504
rect 869 1464 873 1504
rect 881 1464 885 1504
rect 901 1464 905 1504
rect 947 1464 951 1504
rect 955 1464 959 1504
rect 975 1464 979 1484
rect 983 1464 987 1484
rect 1005 1464 1009 1544
rect 1065 1464 1069 1504
rect 1111 1464 1115 1544
rect 1121 1464 1125 1544
rect 1151 1464 1155 1544
rect 1161 1464 1165 1544
rect 1250 1464 1254 1504
rect 1272 1464 1276 1544
rect 1280 1464 1284 1544
rect 1357 1464 1361 1544
rect 1365 1464 1369 1544
rect 1425 1464 1429 1544
rect 1435 1464 1439 1544
rect 1455 1472 1459 1552
rect 1465 1472 1469 1552
rect 1485 1472 1489 1512
rect 1545 1464 1549 1544
rect 1555 1464 1559 1544
rect 1575 1472 1579 1552
rect 1585 1472 1589 1552
rect 1605 1472 1609 1512
rect 1665 1464 1669 1544
rect 1675 1464 1679 1544
rect 1695 1472 1699 1552
rect 1705 1472 1709 1552
rect 1725 1472 1729 1512
rect 1771 1464 1775 1544
rect 1793 1464 1797 1484
rect 1801 1464 1805 1484
rect 1821 1464 1825 1504
rect 1829 1464 1833 1504
rect 1875 1464 1879 1504
rect 1895 1464 1899 1504
rect 1907 1464 1911 1504
rect 1927 1464 1931 1504
rect 1941 1464 1945 1504
rect 1961 1464 1965 1544
rect 2011 1472 2015 1512
rect 2031 1472 2035 1552
rect 2041 1472 2045 1552
rect 2061 1464 2065 1544
rect 2071 1464 2075 1544
rect 2131 1464 2135 1504
rect 2191 1464 2195 1544
rect 2201 1464 2205 1544
rect 2231 1464 2235 1544
rect 2241 1464 2245 1544
rect 2311 1464 2315 1544
rect 2319 1464 2323 1544
rect 2410 1464 2414 1504
rect 2432 1464 2436 1544
rect 2440 1464 2444 1544
rect 2503 1464 2507 1544
rect 2525 1464 2529 1504
rect 2571 1464 2575 1544
rect 2579 1464 2583 1544
rect 2665 1464 2669 1504
rect 2685 1464 2689 1504
rect 2731 1464 2735 1504
rect 2751 1464 2755 1504
rect 2825 1464 2829 1544
rect 2835 1464 2839 1544
rect 2855 1472 2859 1552
rect 2865 1472 2869 1552
rect 2885 1472 2889 1512
rect 2945 1464 2949 1504
rect 2965 1464 2969 1504
rect 2985 1464 2989 1504
rect 3045 1464 3049 1544
rect 3095 1464 3099 1544
rect 3115 1464 3119 1504
rect 3129 1464 3133 1504
rect 3149 1464 3153 1504
rect 3161 1464 3165 1504
rect 3181 1464 3185 1504
rect 3227 1464 3231 1504
rect 3235 1464 3239 1504
rect 3255 1464 3259 1484
rect 3263 1464 3267 1484
rect 3285 1464 3289 1544
rect 3345 1464 3349 1504
rect 3365 1464 3369 1504
rect 3430 1464 3434 1504
rect 3452 1464 3456 1544
rect 3460 1464 3464 1544
rect 3511 1464 3515 1544
rect 3531 1464 3535 1544
rect 3551 1464 3555 1544
rect 3571 1464 3575 1544
rect 3650 1464 3654 1504
rect 3672 1464 3676 1544
rect 3680 1464 3684 1544
rect 3745 1464 3749 1504
rect 3817 1464 3821 1544
rect 3825 1464 3829 1544
rect 3895 1464 3899 1544
rect 3905 1464 3909 1544
rect 3935 1464 3939 1544
rect 3945 1464 3949 1544
rect 4005 1464 4009 1504
rect 4055 1464 4059 1544
rect 4075 1464 4079 1504
rect 4089 1464 4093 1504
rect 4109 1464 4113 1504
rect 4121 1464 4125 1504
rect 4141 1464 4145 1504
rect 4187 1464 4191 1504
rect 4195 1464 4199 1504
rect 4215 1464 4219 1484
rect 4223 1464 4227 1484
rect 4245 1464 4249 1544
rect 4305 1464 4309 1544
rect 4315 1464 4319 1544
rect 4335 1472 4339 1552
rect 4345 1472 4349 1552
rect 4365 1472 4369 1512
rect 4425 1464 4429 1544
rect 4435 1464 4439 1544
rect 4455 1472 4459 1552
rect 4465 1472 4469 1552
rect 4485 1472 4489 1512
rect 4531 1472 4535 1512
rect 4551 1472 4555 1552
rect 4561 1472 4565 1552
rect 4581 1464 4585 1544
rect 4591 1464 4595 1544
rect 4651 1472 4655 1512
rect 4671 1472 4675 1552
rect 4681 1472 4685 1552
rect 4701 1464 4705 1544
rect 4711 1464 4715 1544
rect 4771 1472 4775 1512
rect 4791 1472 4795 1552
rect 4801 1472 4805 1552
rect 4821 1464 4825 1544
rect 4831 1464 4835 1544
rect 4891 1472 4895 1512
rect 4911 1472 4915 1552
rect 4921 1472 4925 1552
rect 4941 1464 4945 1544
rect 4951 1464 4955 1544
rect 5011 1464 5015 1544
rect 5033 1464 5037 1484
rect 5041 1464 5045 1484
rect 5061 1464 5065 1504
rect 5069 1464 5073 1504
rect 5115 1464 5119 1504
rect 5135 1464 5139 1504
rect 5147 1464 5151 1504
rect 5167 1464 5171 1504
rect 5181 1464 5185 1504
rect 5201 1464 5205 1544
rect 5251 1464 5255 1544
rect 5273 1464 5277 1484
rect 5281 1464 5285 1484
rect 5301 1464 5305 1504
rect 5309 1464 5313 1504
rect 5355 1464 5359 1504
rect 5375 1464 5379 1504
rect 5387 1464 5391 1504
rect 5407 1464 5411 1504
rect 5421 1464 5425 1504
rect 5441 1464 5445 1544
rect 5491 1464 5495 1544
rect 5511 1464 5515 1544
rect 5531 1464 5535 1544
rect 5551 1464 5555 1544
rect 5611 1472 5615 1512
rect 5631 1472 5635 1552
rect 5641 1472 5645 1552
rect 5661 1464 5665 1544
rect 5671 1464 5675 1544
rect 5750 1464 5754 1504
rect 5772 1464 5776 1544
rect 5780 1464 5784 1544
rect 5857 1464 5861 1544
rect 5865 1464 5869 1544
rect 5925 1464 5929 1504
rect 5945 1464 5949 1504
rect 6010 1464 6014 1504
rect 6032 1464 6036 1544
rect 6040 1464 6044 1544
rect 6117 1464 6121 1544
rect 6125 1464 6129 1544
rect 6195 1464 6199 1544
rect 6205 1464 6209 1544
rect 6235 1464 6239 1544
rect 6245 1464 6249 1544
rect 6305 1464 6309 1544
rect 6315 1464 6319 1544
rect 6335 1472 6339 1552
rect 6345 1472 6349 1552
rect 6365 1472 6369 1512
rect 6411 1464 6415 1504
rect 6471 1464 6475 1544
rect 6493 1464 6497 1484
rect 6501 1464 6505 1484
rect 6521 1464 6525 1504
rect 6529 1464 6533 1504
rect 6575 1464 6579 1504
rect 6595 1464 6599 1504
rect 6607 1464 6611 1504
rect 6627 1464 6631 1504
rect 6641 1464 6645 1504
rect 6661 1464 6665 1544
rect 31 1396 35 1436
rect 53 1396 57 1436
rect 75 1356 79 1436
rect 131 1356 135 1436
rect 139 1356 143 1436
rect 230 1396 234 1436
rect 252 1356 256 1436
rect 260 1356 264 1436
rect 337 1356 341 1436
rect 345 1356 349 1436
rect 391 1396 395 1436
rect 451 1396 455 1436
rect 525 1396 529 1436
rect 545 1396 549 1436
rect 591 1356 595 1436
rect 611 1356 615 1436
rect 631 1356 635 1436
rect 695 1356 699 1436
rect 715 1396 719 1436
rect 729 1396 733 1436
rect 749 1396 753 1436
rect 761 1396 765 1436
rect 781 1396 785 1436
rect 827 1396 831 1436
rect 835 1396 839 1436
rect 855 1416 859 1436
rect 863 1416 867 1436
rect 885 1356 889 1436
rect 945 1396 949 1436
rect 965 1396 969 1436
rect 1011 1396 1015 1436
rect 1031 1396 1035 1436
rect 1051 1396 1055 1436
rect 1111 1356 1115 1436
rect 1119 1356 1123 1436
rect 1195 1356 1199 1436
rect 1215 1396 1219 1436
rect 1229 1396 1233 1436
rect 1249 1396 1253 1436
rect 1261 1396 1265 1436
rect 1281 1396 1285 1436
rect 1327 1396 1331 1436
rect 1335 1396 1339 1436
rect 1355 1416 1359 1436
rect 1363 1416 1367 1436
rect 1385 1356 1389 1436
rect 1445 1356 1449 1436
rect 1465 1356 1469 1436
rect 1485 1356 1489 1436
rect 1505 1356 1509 1436
rect 1525 1356 1529 1436
rect 1545 1356 1549 1436
rect 1565 1356 1569 1436
rect 1585 1356 1589 1436
rect 1645 1356 1649 1436
rect 1655 1356 1659 1436
rect 1675 1348 1679 1428
rect 1685 1348 1689 1428
rect 1705 1388 1709 1428
rect 1777 1356 1781 1436
rect 1785 1356 1789 1436
rect 1855 1356 1859 1436
rect 1865 1356 1869 1436
rect 1895 1356 1899 1436
rect 1905 1356 1909 1436
rect 1970 1396 1974 1436
rect 1992 1356 1996 1436
rect 2000 1356 2004 1436
rect 2051 1396 2055 1436
rect 2116 1356 2120 1436
rect 2124 1356 2128 1436
rect 2146 1396 2150 1436
rect 2211 1396 2215 1436
rect 2231 1396 2235 1436
rect 2291 1388 2295 1428
rect 2311 1348 2315 1428
rect 2321 1348 2325 1428
rect 2341 1356 2345 1436
rect 2351 1356 2355 1436
rect 2425 1356 2429 1436
rect 2435 1356 2439 1436
rect 2455 1348 2459 1428
rect 2465 1348 2469 1428
rect 2485 1388 2489 1428
rect 2545 1356 2549 1436
rect 2565 1356 2569 1436
rect 2585 1356 2589 1436
rect 2605 1356 2609 1436
rect 2651 1356 2655 1436
rect 2671 1356 2675 1436
rect 2691 1356 2695 1436
rect 2711 1356 2715 1436
rect 2785 1356 2789 1436
rect 2805 1356 2809 1436
rect 2825 1356 2829 1436
rect 2845 1356 2849 1436
rect 2891 1396 2895 1436
rect 2913 1356 2917 1436
rect 2985 1356 2989 1436
rect 3005 1356 3009 1436
rect 3025 1356 3029 1436
rect 3045 1356 3049 1436
rect 3105 1396 3109 1436
rect 3165 1356 3169 1436
rect 3175 1356 3179 1436
rect 3195 1348 3199 1428
rect 3205 1348 3209 1428
rect 3225 1388 3229 1428
rect 3275 1356 3279 1436
rect 3295 1396 3299 1436
rect 3309 1396 3313 1436
rect 3329 1396 3333 1436
rect 3341 1396 3345 1436
rect 3361 1396 3365 1436
rect 3407 1396 3411 1436
rect 3415 1396 3419 1436
rect 3435 1416 3439 1436
rect 3443 1416 3447 1436
rect 3465 1356 3469 1436
rect 3537 1356 3541 1436
rect 3545 1356 3549 1436
rect 3615 1356 3619 1436
rect 3625 1356 3629 1436
rect 3655 1356 3659 1436
rect 3665 1356 3669 1436
rect 3730 1396 3734 1436
rect 3752 1356 3756 1436
rect 3760 1356 3764 1436
rect 3825 1396 3829 1436
rect 3871 1356 3875 1436
rect 3893 1416 3897 1436
rect 3901 1416 3905 1436
rect 3921 1396 3925 1436
rect 3929 1396 3933 1436
rect 3975 1396 3979 1436
rect 3995 1396 3999 1436
rect 4007 1396 4011 1436
rect 4027 1396 4031 1436
rect 4041 1396 4045 1436
rect 4061 1356 4065 1436
rect 4111 1356 4115 1436
rect 4133 1416 4137 1436
rect 4141 1416 4145 1436
rect 4161 1396 4165 1436
rect 4169 1396 4173 1436
rect 4215 1396 4219 1436
rect 4235 1396 4239 1436
rect 4247 1396 4251 1436
rect 4267 1396 4271 1436
rect 4281 1396 4285 1436
rect 4301 1356 4305 1436
rect 4365 1396 4369 1436
rect 4411 1356 4415 1436
rect 4431 1356 4435 1436
rect 4451 1356 4455 1436
rect 4471 1356 4475 1436
rect 4531 1388 4535 1428
rect 4551 1348 4555 1428
rect 4561 1348 4565 1428
rect 4581 1356 4585 1436
rect 4591 1356 4595 1436
rect 4665 1356 4669 1436
rect 4685 1356 4689 1436
rect 4705 1356 4709 1436
rect 4725 1356 4729 1436
rect 4783 1356 4787 1436
rect 4805 1396 4809 1436
rect 4865 1396 4869 1436
rect 4885 1396 4889 1436
rect 4945 1396 4949 1436
rect 4965 1396 4969 1436
rect 5035 1356 5039 1436
rect 5045 1356 5049 1436
rect 5075 1356 5079 1436
rect 5085 1356 5089 1436
rect 5155 1356 5159 1436
rect 5165 1356 5169 1436
rect 5195 1356 5199 1436
rect 5205 1356 5209 1436
rect 5251 1356 5255 1436
rect 5325 1396 5329 1436
rect 5345 1396 5349 1436
rect 5391 1356 5395 1436
rect 5401 1356 5405 1436
rect 5431 1356 5435 1436
rect 5441 1356 5445 1436
rect 5525 1356 5529 1436
rect 5545 1356 5549 1436
rect 5565 1356 5569 1436
rect 5611 1356 5615 1436
rect 5671 1388 5675 1428
rect 5691 1348 5695 1428
rect 5701 1348 5705 1428
rect 5721 1356 5725 1436
rect 5731 1356 5735 1436
rect 5805 1396 5809 1436
rect 5825 1396 5829 1436
rect 5890 1396 5894 1436
rect 5912 1356 5916 1436
rect 5920 1356 5924 1436
rect 5985 1396 5989 1436
rect 6036 1356 6040 1436
rect 6044 1356 6048 1436
rect 6066 1396 6070 1436
rect 6131 1356 6135 1436
rect 6141 1356 6145 1436
rect 6171 1356 6175 1436
rect 6181 1356 6185 1436
rect 6251 1356 6255 1436
rect 6273 1416 6277 1436
rect 6281 1416 6285 1436
rect 6301 1396 6305 1436
rect 6309 1396 6313 1436
rect 6355 1396 6359 1436
rect 6375 1396 6379 1436
rect 6387 1396 6391 1436
rect 6407 1396 6411 1436
rect 6421 1396 6425 1436
rect 6441 1356 6445 1436
rect 6491 1356 6495 1436
rect 6513 1416 6517 1436
rect 6521 1416 6525 1436
rect 6541 1396 6545 1436
rect 6549 1396 6553 1436
rect 6595 1396 6599 1436
rect 6615 1396 6619 1436
rect 6627 1396 6631 1436
rect 6647 1396 6651 1436
rect 6661 1396 6665 1436
rect 6681 1356 6685 1436
rect 31 984 35 1064
rect 53 984 57 1004
rect 61 984 65 1004
rect 81 984 85 1024
rect 89 984 93 1024
rect 135 984 139 1024
rect 155 984 159 1024
rect 167 984 171 1024
rect 187 984 191 1024
rect 201 984 205 1024
rect 221 984 225 1064
rect 285 984 289 1024
rect 331 984 335 1064
rect 353 984 357 1004
rect 361 984 365 1004
rect 381 984 385 1024
rect 389 984 393 1024
rect 435 984 439 1024
rect 455 984 459 1024
rect 467 984 471 1024
rect 487 984 491 1024
rect 501 984 505 1024
rect 521 984 525 1064
rect 571 984 575 1024
rect 631 984 635 1024
rect 651 984 655 1024
rect 671 984 675 1024
rect 731 984 735 1064
rect 739 984 743 1064
rect 811 984 815 1024
rect 831 984 835 1024
rect 851 984 855 1024
rect 911 984 915 1024
rect 931 984 935 1024
rect 991 984 995 1024
rect 1055 984 1059 1064
rect 1075 984 1079 1024
rect 1089 984 1093 1024
rect 1109 984 1113 1024
rect 1121 984 1125 1024
rect 1141 984 1145 1024
rect 1187 984 1191 1024
rect 1195 984 1199 1024
rect 1215 984 1219 1004
rect 1223 984 1227 1004
rect 1245 984 1249 1064
rect 1291 984 1295 1064
rect 1311 984 1315 1064
rect 1331 984 1335 1064
rect 1351 984 1355 1064
rect 1371 984 1375 1064
rect 1391 984 1395 1064
rect 1411 984 1415 1064
rect 1431 984 1435 1064
rect 1495 984 1499 1064
rect 1515 984 1519 1024
rect 1529 984 1533 1024
rect 1549 984 1553 1024
rect 1561 984 1565 1024
rect 1581 984 1585 1024
rect 1627 984 1631 1024
rect 1635 984 1639 1024
rect 1655 984 1659 1004
rect 1663 984 1667 1004
rect 1685 984 1689 1064
rect 1757 984 1761 1064
rect 1765 984 1769 1064
rect 1835 984 1839 1064
rect 1845 984 1849 1064
rect 1875 984 1879 1064
rect 1885 984 1889 1064
rect 1950 984 1954 1024
rect 1972 984 1976 1064
rect 1980 984 1984 1064
rect 2050 984 2054 1024
rect 2072 984 2076 1064
rect 2080 984 2084 1064
rect 2157 984 2161 1064
rect 2165 984 2169 1064
rect 2235 984 2239 1064
rect 2245 984 2249 1064
rect 2275 984 2279 1064
rect 2285 984 2289 1064
rect 2335 984 2339 1064
rect 2355 984 2359 1024
rect 2369 984 2373 1024
rect 2389 984 2393 1024
rect 2401 984 2405 1024
rect 2421 984 2425 1024
rect 2467 984 2471 1024
rect 2475 984 2479 1024
rect 2495 984 2499 1004
rect 2503 984 2507 1004
rect 2525 984 2529 1064
rect 2585 984 2589 1024
rect 2636 984 2640 1064
rect 2644 984 2648 1064
rect 2666 984 2670 1024
rect 2743 984 2747 1064
rect 2765 984 2769 1024
rect 2811 984 2815 1024
rect 2885 984 2889 1064
rect 2905 984 2909 1064
rect 2925 984 2929 1064
rect 2945 984 2949 1064
rect 2995 984 2999 1064
rect 3015 984 3019 1024
rect 3029 984 3033 1024
rect 3049 984 3053 1024
rect 3061 984 3065 1024
rect 3081 984 3085 1024
rect 3127 984 3131 1024
rect 3135 984 3139 1024
rect 3155 984 3159 1004
rect 3163 984 3167 1004
rect 3185 984 3189 1064
rect 3231 984 3235 1024
rect 3251 984 3255 1024
rect 3325 984 3329 1064
rect 3335 984 3339 1064
rect 3355 992 3359 1072
rect 3365 992 3369 1072
rect 3385 992 3389 1032
rect 3431 992 3435 1032
rect 3451 992 3455 1072
rect 3461 992 3465 1072
rect 3481 984 3485 1064
rect 3491 984 3495 1064
rect 3563 984 3567 1064
rect 3585 984 3589 1024
rect 3635 984 3639 1064
rect 3655 984 3659 1024
rect 3669 984 3673 1024
rect 3689 984 3693 1024
rect 3701 984 3705 1024
rect 3721 984 3725 1024
rect 3767 984 3771 1024
rect 3775 984 3779 1024
rect 3795 984 3799 1004
rect 3803 984 3807 1004
rect 3825 984 3829 1064
rect 3871 992 3875 1032
rect 3891 992 3895 1072
rect 3901 992 3905 1072
rect 3921 984 3925 1064
rect 3931 984 3935 1064
rect 4005 984 4009 1064
rect 4015 984 4019 1064
rect 4035 992 4039 1072
rect 4045 992 4049 1072
rect 4065 992 4069 1032
rect 4111 984 4115 1024
rect 4171 984 4175 1064
rect 4181 984 4185 1064
rect 4211 984 4215 1064
rect 4221 984 4225 1064
rect 4291 984 4295 1064
rect 4299 984 4303 1064
rect 4390 984 4394 1024
rect 4412 984 4416 1064
rect 4420 984 4424 1064
rect 4485 984 4489 1064
rect 4505 984 4509 1064
rect 4525 984 4529 1064
rect 4575 984 4579 1064
rect 4595 984 4599 1024
rect 4609 984 4613 1024
rect 4629 984 4633 1024
rect 4641 984 4645 1024
rect 4661 984 4665 1024
rect 4707 984 4711 1024
rect 4715 984 4719 1024
rect 4735 984 4739 1004
rect 4743 984 4747 1004
rect 4765 984 4769 1064
rect 4811 984 4815 1064
rect 4821 984 4825 1064
rect 4851 984 4855 1064
rect 4861 984 4865 1064
rect 4957 984 4961 1064
rect 4965 984 4969 1064
rect 5030 984 5034 1024
rect 5052 984 5056 1064
rect 5060 984 5064 1064
rect 5137 984 5141 1064
rect 5145 984 5149 1064
rect 5191 984 5195 1064
rect 5199 984 5203 1064
rect 5271 984 5275 1064
rect 5279 984 5283 1064
rect 5363 984 5367 1064
rect 5385 984 5389 1024
rect 5431 984 5435 1064
rect 5439 984 5443 1064
rect 5511 984 5515 1064
rect 5519 984 5523 1064
rect 5591 984 5595 1064
rect 5611 984 5615 1064
rect 5631 984 5635 1064
rect 5691 984 5695 1064
rect 5701 984 5705 1064
rect 5721 984 5725 1064
rect 5817 984 5821 1064
rect 5825 984 5829 1064
rect 5876 984 5880 1064
rect 5884 984 5888 1064
rect 5906 984 5910 1024
rect 5985 984 5989 1024
rect 6005 984 6009 1024
rect 6025 984 6029 1024
rect 6076 984 6080 1064
rect 6084 984 6088 1064
rect 6106 984 6110 1024
rect 6197 984 6201 1064
rect 6205 984 6209 1064
rect 6251 984 6255 1064
rect 6259 984 6263 1064
rect 6331 984 6335 1064
rect 6353 984 6357 1004
rect 6361 984 6365 1004
rect 6381 984 6385 1024
rect 6389 984 6393 1024
rect 6435 984 6439 1024
rect 6455 984 6459 1024
rect 6467 984 6471 1024
rect 6487 984 6491 1024
rect 6501 984 6505 1024
rect 6521 984 6525 1064
rect 6571 984 6575 1064
rect 6581 984 6585 1064
rect 6611 984 6615 1064
rect 6621 984 6625 1064
rect 31 876 35 956
rect 41 876 45 956
rect 61 876 65 956
rect 145 916 149 956
rect 165 916 169 956
rect 211 876 215 956
rect 233 936 237 956
rect 241 936 245 956
rect 261 916 265 956
rect 269 916 273 956
rect 315 916 319 956
rect 335 916 339 956
rect 347 916 351 956
rect 367 916 371 956
rect 381 916 385 956
rect 401 876 405 956
rect 465 916 469 956
rect 537 876 541 956
rect 545 876 549 956
rect 591 876 595 956
rect 599 876 603 956
rect 671 916 675 956
rect 691 916 695 956
rect 751 916 755 956
rect 771 916 775 956
rect 791 916 795 956
rect 851 876 855 956
rect 861 876 865 956
rect 891 876 895 956
rect 901 876 905 956
rect 976 876 980 956
rect 984 876 988 956
rect 1006 916 1010 956
rect 1076 876 1080 956
rect 1084 876 1088 956
rect 1106 916 1110 956
rect 1181 888 1185 948
rect 1201 888 1205 948
rect 1245 896 1249 956
rect 1265 896 1269 956
rect 1285 896 1289 956
rect 1305 896 1309 956
rect 1356 876 1360 956
rect 1364 876 1368 956
rect 1386 916 1390 956
rect 1465 916 1469 956
rect 1515 876 1519 956
rect 1535 916 1539 956
rect 1549 916 1553 956
rect 1569 916 1573 956
rect 1581 916 1585 956
rect 1601 916 1605 956
rect 1647 916 1651 956
rect 1655 916 1659 956
rect 1675 936 1679 956
rect 1683 936 1687 956
rect 1705 876 1709 956
rect 1751 916 1755 956
rect 1811 908 1815 948
rect 1831 868 1835 948
rect 1841 868 1845 948
rect 1861 876 1865 956
rect 1871 876 1875 956
rect 1936 876 1940 956
rect 1944 876 1948 956
rect 1966 916 1970 956
rect 2031 916 2035 956
rect 2051 916 2055 956
rect 2111 876 2115 956
rect 2133 936 2137 956
rect 2141 936 2145 956
rect 2161 916 2165 956
rect 2169 916 2173 956
rect 2215 916 2219 956
rect 2235 916 2239 956
rect 2247 916 2251 956
rect 2267 916 2271 956
rect 2281 916 2285 956
rect 2301 876 2305 956
rect 2351 916 2355 956
rect 2411 876 2415 956
rect 2421 876 2425 956
rect 2451 876 2455 956
rect 2461 876 2465 956
rect 2531 876 2535 956
rect 2539 876 2543 956
rect 2630 916 2634 956
rect 2652 876 2656 956
rect 2660 876 2664 956
rect 2725 876 2729 956
rect 2745 876 2749 956
rect 2765 876 2769 956
rect 2785 876 2789 956
rect 2805 876 2809 956
rect 2825 876 2829 956
rect 2845 876 2849 956
rect 2865 876 2869 956
rect 2911 876 2915 956
rect 2931 876 2935 956
rect 2951 876 2955 956
rect 3025 876 3029 956
rect 3045 876 3049 956
rect 3065 876 3069 956
rect 3125 876 3129 956
rect 3135 876 3139 956
rect 3155 868 3159 948
rect 3165 868 3169 948
rect 3185 908 3189 948
rect 3245 876 3249 956
rect 3255 876 3259 956
rect 3275 868 3279 948
rect 3285 868 3289 948
rect 3305 908 3309 948
rect 3370 916 3374 956
rect 3392 876 3396 956
rect 3400 876 3404 956
rect 3451 916 3455 956
rect 3471 916 3475 956
rect 3531 908 3535 948
rect 3551 868 3555 948
rect 3561 868 3565 948
rect 3581 876 3585 956
rect 3591 876 3595 956
rect 3665 916 3669 956
rect 3725 876 3729 956
rect 3735 876 3739 956
rect 3755 868 3759 948
rect 3765 868 3769 948
rect 3785 908 3789 948
rect 3835 876 3839 956
rect 3855 916 3859 956
rect 3869 916 3873 956
rect 3889 916 3893 956
rect 3901 916 3905 956
rect 3921 916 3925 956
rect 3967 916 3971 956
rect 3975 916 3979 956
rect 3995 936 3999 956
rect 4003 936 4007 956
rect 4025 876 4029 956
rect 4071 908 4075 948
rect 4091 868 4095 948
rect 4101 868 4105 948
rect 4121 876 4125 956
rect 4131 876 4135 956
rect 4191 876 4195 956
rect 4211 876 4215 956
rect 4231 876 4235 956
rect 4296 876 4300 956
rect 4304 876 4308 956
rect 4326 916 4330 956
rect 4405 916 4409 956
rect 4425 916 4429 956
rect 4445 916 4449 956
rect 4491 916 4495 956
rect 4556 876 4560 956
rect 4564 876 4568 956
rect 4586 916 4590 956
rect 4651 916 4655 956
rect 4671 916 4675 956
rect 4745 916 4749 956
rect 4796 876 4800 956
rect 4804 876 4808 956
rect 4826 916 4830 956
rect 4891 916 4895 956
rect 4911 916 4915 956
rect 4971 908 4975 948
rect 4991 868 4995 948
rect 5001 868 5005 948
rect 5021 876 5025 956
rect 5031 876 5035 956
rect 5105 876 5109 956
rect 5115 876 5119 956
rect 5135 868 5139 948
rect 5145 868 5149 948
rect 5165 908 5169 948
rect 5211 876 5215 956
rect 5231 876 5235 956
rect 5251 876 5255 956
rect 5271 876 5275 956
rect 5291 876 5295 956
rect 5311 876 5315 956
rect 5331 876 5335 956
rect 5351 876 5355 956
rect 5411 876 5415 956
rect 5431 876 5435 956
rect 5451 876 5455 956
rect 5525 916 5529 956
rect 5576 876 5580 956
rect 5584 876 5588 956
rect 5606 916 5610 956
rect 5671 916 5675 956
rect 5691 916 5695 956
rect 5756 876 5760 956
rect 5764 876 5768 956
rect 5786 916 5790 956
rect 5865 916 5869 956
rect 5885 916 5889 956
rect 5905 916 5909 956
rect 5955 876 5959 956
rect 5975 916 5979 956
rect 5989 916 5993 956
rect 6009 916 6013 956
rect 6021 916 6025 956
rect 6041 916 6045 956
rect 6087 916 6091 956
rect 6095 916 6099 956
rect 6115 936 6119 956
rect 6123 936 6127 956
rect 6145 876 6149 956
rect 6196 876 6200 956
rect 6204 876 6208 956
rect 6226 916 6230 956
rect 6296 876 6300 956
rect 6304 876 6308 956
rect 6326 916 6330 956
rect 6405 916 6409 956
rect 6425 916 6429 956
rect 6475 876 6479 956
rect 6495 916 6499 956
rect 6509 916 6513 956
rect 6529 916 6533 956
rect 6541 916 6545 956
rect 6561 916 6565 956
rect 6607 916 6611 956
rect 6615 916 6619 956
rect 6635 936 6639 956
rect 6643 936 6647 956
rect 6665 876 6669 956
rect 31 504 35 544
rect 91 504 95 544
rect 111 504 115 544
rect 171 504 175 584
rect 191 504 195 584
rect 211 504 215 584
rect 271 504 275 544
rect 345 504 349 584
rect 365 504 369 584
rect 385 504 389 584
rect 431 504 435 544
rect 451 504 455 544
rect 471 504 475 544
rect 545 504 549 544
rect 565 504 569 544
rect 625 504 629 544
rect 645 504 649 544
rect 665 504 669 544
rect 711 504 715 544
rect 771 504 775 544
rect 857 504 861 584
rect 865 504 869 584
rect 921 512 925 572
rect 941 512 945 572
rect 985 504 989 564
rect 1005 504 1009 564
rect 1025 504 1029 564
rect 1045 504 1049 564
rect 1095 504 1099 584
rect 1115 504 1119 544
rect 1129 504 1133 544
rect 1149 504 1153 544
rect 1161 504 1165 544
rect 1181 504 1185 544
rect 1227 504 1231 544
rect 1235 504 1239 544
rect 1255 504 1259 524
rect 1263 504 1267 524
rect 1285 504 1289 584
rect 1331 504 1335 544
rect 1353 504 1357 584
rect 1411 504 1415 544
rect 1431 504 1435 544
rect 1495 504 1499 584
rect 1515 504 1519 544
rect 1529 504 1533 544
rect 1549 504 1553 544
rect 1561 504 1565 544
rect 1581 504 1585 544
rect 1627 504 1631 544
rect 1635 504 1639 544
rect 1655 504 1659 524
rect 1663 504 1667 524
rect 1685 504 1689 584
rect 1735 504 1739 584
rect 1755 504 1759 544
rect 1769 504 1773 544
rect 1789 504 1793 544
rect 1801 504 1805 544
rect 1821 504 1825 544
rect 1867 504 1871 544
rect 1875 504 1879 544
rect 1895 504 1899 524
rect 1903 504 1907 524
rect 1925 504 1929 584
rect 1975 504 1979 584
rect 1995 504 1999 544
rect 2009 504 2013 544
rect 2029 504 2033 544
rect 2041 504 2045 544
rect 2061 504 2065 544
rect 2107 504 2111 544
rect 2115 504 2119 544
rect 2135 504 2139 524
rect 2143 504 2147 524
rect 2165 504 2169 584
rect 2215 504 2219 584
rect 2235 504 2239 544
rect 2249 504 2253 544
rect 2269 504 2273 544
rect 2281 504 2285 544
rect 2301 504 2305 544
rect 2347 504 2351 544
rect 2355 504 2359 544
rect 2375 504 2379 524
rect 2383 504 2387 524
rect 2405 504 2409 584
rect 2451 504 2455 584
rect 2473 504 2477 524
rect 2481 504 2485 524
rect 2501 504 2505 544
rect 2509 504 2513 544
rect 2555 504 2559 544
rect 2575 504 2579 544
rect 2587 504 2591 544
rect 2607 504 2611 544
rect 2621 504 2625 544
rect 2641 504 2645 584
rect 2705 504 2709 584
rect 2725 504 2729 584
rect 2745 504 2749 584
rect 2765 504 2769 584
rect 2825 504 2829 544
rect 2885 504 2889 584
rect 2905 504 2909 584
rect 2925 504 2929 584
rect 2971 504 2975 544
rect 3036 504 3040 584
rect 3044 504 3048 584
rect 3066 504 3070 544
rect 3131 504 3135 544
rect 3151 504 3155 544
rect 3211 504 3215 544
rect 3231 504 3235 544
rect 3251 504 3255 544
rect 3311 504 3315 544
rect 3376 504 3380 584
rect 3384 504 3388 584
rect 3406 504 3410 544
rect 3471 504 3475 544
rect 3491 504 3495 544
rect 3551 504 3555 584
rect 3571 504 3575 584
rect 3591 504 3595 584
rect 3651 504 3655 584
rect 3659 504 3663 584
rect 3736 504 3740 584
rect 3744 504 3748 584
rect 3766 504 3770 544
rect 3845 504 3849 544
rect 3865 504 3869 544
rect 3885 504 3889 544
rect 3931 504 3935 584
rect 3953 504 3957 524
rect 3961 504 3965 524
rect 3981 504 3985 544
rect 3989 504 3993 544
rect 4035 504 4039 544
rect 4055 504 4059 544
rect 4067 504 4071 544
rect 4087 504 4091 544
rect 4101 504 4105 544
rect 4121 504 4125 584
rect 4197 504 4201 584
rect 4205 504 4209 584
rect 4251 504 4255 584
rect 4273 504 4277 524
rect 4281 504 4285 524
rect 4301 504 4305 544
rect 4309 504 4313 544
rect 4355 504 4359 544
rect 4375 504 4379 544
rect 4387 504 4391 544
rect 4407 504 4411 544
rect 4421 504 4425 544
rect 4441 504 4445 584
rect 4491 504 4495 544
rect 4551 504 4555 584
rect 4571 504 4575 584
rect 4591 504 4595 584
rect 4611 504 4615 584
rect 4685 504 4689 584
rect 4705 504 4709 584
rect 4725 504 4729 584
rect 4790 504 4794 544
rect 4812 504 4816 584
rect 4820 504 4824 584
rect 4871 504 4875 544
rect 4891 504 4895 544
rect 4965 504 4969 544
rect 5025 504 5029 584
rect 5035 504 5039 584
rect 5055 512 5059 592
rect 5065 512 5069 592
rect 5085 512 5089 552
rect 5131 504 5135 544
rect 5151 504 5155 544
rect 5171 504 5175 544
rect 5231 504 5235 584
rect 5253 504 5257 524
rect 5261 504 5265 524
rect 5281 504 5285 544
rect 5289 504 5293 544
rect 5335 504 5339 544
rect 5355 504 5359 544
rect 5367 504 5371 544
rect 5387 504 5391 544
rect 5401 504 5405 544
rect 5421 504 5425 584
rect 5471 504 5475 584
rect 5531 512 5535 552
rect 5551 512 5555 592
rect 5561 512 5565 592
rect 5581 504 5585 584
rect 5591 504 5595 584
rect 5677 504 5681 584
rect 5685 504 5689 584
rect 5757 504 5761 584
rect 5765 504 5769 584
rect 5837 504 5841 584
rect 5845 504 5849 584
rect 5891 504 5895 584
rect 5899 504 5903 584
rect 5997 504 6001 584
rect 6005 504 6009 584
rect 6056 504 6060 584
rect 6064 504 6068 584
rect 6086 504 6090 544
rect 6156 504 6160 584
rect 6164 504 6168 584
rect 6186 504 6190 544
rect 6265 504 6269 544
rect 6285 504 6289 544
rect 6335 504 6339 584
rect 6355 504 6359 544
rect 6369 504 6373 544
rect 6389 504 6393 544
rect 6401 504 6405 544
rect 6421 504 6425 544
rect 6467 504 6471 544
rect 6475 504 6479 544
rect 6495 504 6499 524
rect 6503 504 6507 524
rect 6525 504 6529 584
rect 6571 504 6575 544
rect 6631 504 6635 544
rect 31 396 35 476
rect 53 456 57 476
rect 61 456 65 476
rect 81 436 85 476
rect 89 436 93 476
rect 135 436 139 476
rect 155 436 159 476
rect 167 436 171 476
rect 187 436 191 476
rect 201 436 205 476
rect 221 396 225 476
rect 275 396 279 476
rect 295 436 299 476
rect 309 436 313 476
rect 329 436 333 476
rect 341 436 345 476
rect 361 436 365 476
rect 407 436 411 476
rect 415 436 419 476
rect 435 456 439 476
rect 443 456 447 476
rect 465 396 469 476
rect 511 436 515 476
rect 531 436 535 476
rect 551 436 555 476
rect 611 396 615 476
rect 619 396 623 476
rect 717 396 721 476
rect 725 396 729 476
rect 771 436 775 476
rect 791 436 795 476
rect 865 436 869 476
rect 915 396 919 476
rect 935 436 939 476
rect 949 436 953 476
rect 969 436 973 476
rect 981 436 985 476
rect 1001 436 1005 476
rect 1047 436 1051 476
rect 1055 436 1059 476
rect 1075 456 1079 476
rect 1083 456 1087 476
rect 1105 396 1109 476
rect 1163 396 1167 476
rect 1185 436 1189 476
rect 1231 436 1235 476
rect 1253 396 1257 476
rect 1311 436 1315 476
rect 1333 396 1337 476
rect 1405 436 1409 476
rect 1456 396 1460 476
rect 1464 396 1468 476
rect 1486 436 1490 476
rect 1565 436 1569 476
rect 1616 396 1620 476
rect 1624 396 1628 476
rect 1646 436 1650 476
rect 1715 396 1719 476
rect 1735 436 1739 476
rect 1749 436 1753 476
rect 1769 436 1773 476
rect 1781 436 1785 476
rect 1801 436 1805 476
rect 1847 436 1851 476
rect 1855 436 1859 476
rect 1875 456 1879 476
rect 1883 456 1887 476
rect 1905 396 1909 476
rect 1965 436 1969 476
rect 2025 436 2029 476
rect 2076 396 2080 476
rect 2084 396 2088 476
rect 2106 436 2110 476
rect 2171 436 2175 476
rect 2231 396 2235 476
rect 2241 396 2245 476
rect 2271 396 2275 476
rect 2281 396 2285 476
rect 2370 436 2374 476
rect 2392 396 2396 476
rect 2400 396 2404 476
rect 2451 396 2455 476
rect 2459 396 2463 476
rect 2535 396 2539 476
rect 2555 436 2559 476
rect 2569 436 2573 476
rect 2589 436 2593 476
rect 2601 436 2605 476
rect 2621 436 2625 476
rect 2667 436 2671 476
rect 2675 436 2679 476
rect 2695 456 2699 476
rect 2703 456 2707 476
rect 2725 396 2729 476
rect 2790 436 2794 476
rect 2812 396 2816 476
rect 2820 396 2824 476
rect 2871 396 2875 476
rect 2879 396 2883 476
rect 2955 396 2959 476
rect 2975 436 2979 476
rect 2989 436 2993 476
rect 3009 436 3013 476
rect 3021 436 3025 476
rect 3041 436 3045 476
rect 3087 436 3091 476
rect 3095 436 3099 476
rect 3115 456 3119 476
rect 3123 456 3127 476
rect 3145 396 3149 476
rect 3191 436 3195 476
rect 3211 436 3215 476
rect 3290 436 3294 476
rect 3312 396 3316 476
rect 3320 396 3324 476
rect 3371 396 3375 476
rect 3379 396 3383 476
rect 3465 396 3469 476
rect 3485 396 3489 476
rect 3505 396 3509 476
rect 3556 396 3560 476
rect 3564 396 3568 476
rect 3586 436 3590 476
rect 3651 396 3655 476
rect 3659 396 3663 476
rect 3731 396 3735 476
rect 3751 396 3755 476
rect 3771 396 3775 476
rect 3857 396 3861 476
rect 3865 396 3869 476
rect 3916 396 3920 476
rect 3924 396 3928 476
rect 3946 436 3950 476
rect 4025 436 4029 476
rect 4045 436 4049 476
rect 4065 436 4069 476
rect 4111 396 4115 476
rect 4119 396 4123 476
rect 4191 396 4195 476
rect 4213 456 4217 476
rect 4221 456 4225 476
rect 4241 436 4245 476
rect 4249 436 4253 476
rect 4295 436 4299 476
rect 4315 436 4319 476
rect 4327 436 4331 476
rect 4347 436 4351 476
rect 4361 436 4365 476
rect 4381 396 4385 476
rect 4431 396 4435 476
rect 4439 396 4443 476
rect 4530 436 4534 476
rect 4552 396 4556 476
rect 4560 396 4564 476
rect 4611 396 4615 476
rect 4619 396 4623 476
rect 4715 396 4719 476
rect 4725 396 4729 476
rect 4755 396 4759 476
rect 4765 396 4769 476
rect 4825 436 4829 476
rect 4875 396 4879 476
rect 4895 436 4899 476
rect 4909 436 4913 476
rect 4929 436 4933 476
rect 4941 436 4945 476
rect 4961 436 4965 476
rect 5007 436 5011 476
rect 5015 436 5019 476
rect 5035 456 5039 476
rect 5043 456 5047 476
rect 5065 396 5069 476
rect 5125 396 5129 476
rect 5145 396 5149 476
rect 5165 396 5169 476
rect 5211 396 5215 476
rect 5219 396 5223 476
rect 5310 436 5314 476
rect 5332 396 5336 476
rect 5340 396 5344 476
rect 5391 396 5395 476
rect 5399 396 5403 476
rect 5471 396 5475 476
rect 5491 396 5495 476
rect 5511 396 5515 476
rect 5571 436 5575 476
rect 5591 436 5595 476
rect 5611 436 5615 476
rect 5676 396 5680 476
rect 5684 396 5688 476
rect 5706 436 5710 476
rect 5785 436 5789 476
rect 5805 436 5809 476
rect 5870 436 5874 476
rect 5892 396 5896 476
rect 5900 396 5904 476
rect 5956 396 5960 476
rect 5964 396 5968 476
rect 5986 436 5990 476
rect 6056 396 6060 476
rect 6064 396 6068 476
rect 6086 436 6090 476
rect 6177 396 6181 476
rect 6185 396 6189 476
rect 6257 396 6261 476
rect 6265 396 6269 476
rect 6335 396 6339 476
rect 6345 396 6349 476
rect 6375 396 6379 476
rect 6385 396 6389 476
rect 6435 396 6439 476
rect 6455 436 6459 476
rect 6469 436 6473 476
rect 6489 436 6493 476
rect 6501 436 6505 476
rect 6521 436 6525 476
rect 6567 436 6571 476
rect 6575 436 6579 476
rect 6595 456 6599 476
rect 6603 456 6607 476
rect 6625 396 6629 476
rect 31 24 35 104
rect 53 24 57 44
rect 61 24 65 44
rect 81 24 85 64
rect 89 24 93 64
rect 135 24 139 64
rect 155 24 159 64
rect 167 24 171 64
rect 187 24 191 64
rect 201 24 205 64
rect 221 24 225 104
rect 271 24 275 104
rect 293 24 297 44
rect 301 24 305 44
rect 321 24 325 64
rect 329 24 333 64
rect 375 24 379 64
rect 395 24 399 64
rect 407 24 411 64
rect 427 24 431 64
rect 441 24 445 64
rect 461 24 465 104
rect 523 24 527 104
rect 545 24 549 64
rect 591 24 595 64
rect 613 24 617 104
rect 683 24 687 104
rect 705 24 709 64
rect 751 24 755 104
rect 773 24 777 44
rect 781 24 785 44
rect 801 24 805 64
rect 809 24 813 64
rect 855 24 859 64
rect 875 24 879 64
rect 887 24 891 64
rect 907 24 911 64
rect 921 24 925 64
rect 941 24 945 104
rect 991 24 995 64
rect 1013 24 1017 104
rect 1085 24 1089 64
rect 1105 24 1109 64
rect 1170 24 1174 64
rect 1192 24 1196 104
rect 1200 24 1204 104
rect 1255 24 1259 104
rect 1275 24 1279 64
rect 1289 24 1293 64
rect 1309 24 1313 64
rect 1321 24 1325 64
rect 1341 24 1345 64
rect 1387 24 1391 64
rect 1395 24 1399 64
rect 1415 24 1419 44
rect 1423 24 1427 44
rect 1445 24 1449 104
rect 1505 24 1509 64
rect 1551 24 1555 64
rect 1571 24 1575 64
rect 1650 24 1654 64
rect 1672 24 1676 104
rect 1680 24 1684 104
rect 1731 24 1735 64
rect 1791 24 1795 64
rect 1811 24 1815 64
rect 1871 24 1875 64
rect 1891 24 1895 64
rect 1951 24 1955 64
rect 1971 24 1975 64
rect 2050 24 2054 64
rect 2072 24 2076 104
rect 2080 24 2084 104
rect 2135 24 2139 104
rect 2155 24 2159 64
rect 2169 24 2173 64
rect 2189 24 2193 64
rect 2201 24 2205 64
rect 2221 24 2225 64
rect 2267 24 2271 64
rect 2275 24 2279 64
rect 2295 24 2299 44
rect 2303 24 2307 44
rect 2325 24 2329 104
rect 2371 24 2375 64
rect 2391 24 2395 64
rect 2465 24 2469 64
rect 2485 24 2489 64
rect 2550 24 2554 64
rect 2572 24 2576 104
rect 2580 24 2584 104
rect 2645 24 2649 64
rect 2695 24 2699 104
rect 2715 24 2719 64
rect 2729 24 2733 64
rect 2749 24 2753 64
rect 2761 24 2765 64
rect 2781 24 2785 64
rect 2827 24 2831 64
rect 2835 24 2839 64
rect 2855 24 2859 44
rect 2863 24 2867 44
rect 2885 24 2889 104
rect 2950 24 2954 64
rect 2972 24 2976 104
rect 2980 24 2984 104
rect 3057 24 3061 104
rect 3065 24 3069 104
rect 3135 24 3139 104
rect 3145 24 3149 104
rect 3175 24 3179 104
rect 3185 24 3189 104
rect 3245 24 3249 64
rect 3291 24 3295 104
rect 3313 24 3317 44
rect 3321 24 3325 44
rect 3341 24 3345 64
rect 3349 24 3353 64
rect 3395 24 3399 64
rect 3415 24 3419 64
rect 3427 24 3431 64
rect 3447 24 3451 64
rect 3461 24 3465 64
rect 3481 24 3485 104
rect 3545 24 3549 64
rect 3565 24 3569 64
rect 3630 24 3634 64
rect 3652 24 3656 104
rect 3660 24 3664 104
rect 3716 24 3720 104
rect 3724 24 3728 104
rect 3746 24 3750 64
rect 3811 24 3815 104
rect 3833 24 3837 44
rect 3841 24 3845 44
rect 3861 24 3865 64
rect 3869 24 3873 64
rect 3915 24 3919 64
rect 3935 24 3939 64
rect 3947 24 3951 64
rect 3967 24 3971 64
rect 3981 24 3985 64
rect 4001 24 4005 104
rect 4056 24 4060 104
rect 4064 24 4068 104
rect 4086 24 4090 64
rect 4156 24 4160 104
rect 4164 24 4168 104
rect 4186 24 4190 64
rect 4251 24 4255 64
rect 4271 24 4275 64
rect 4331 24 4335 104
rect 4353 24 4357 44
rect 4361 24 4365 44
rect 4381 24 4385 64
rect 4389 24 4393 64
rect 4435 24 4439 64
rect 4455 24 4459 64
rect 4467 24 4471 64
rect 4487 24 4491 64
rect 4501 24 4505 64
rect 4521 24 4525 104
rect 4576 24 4580 104
rect 4584 24 4588 104
rect 4606 24 4610 64
rect 4676 24 4680 104
rect 4684 24 4688 104
rect 4706 24 4710 64
rect 4771 24 4775 64
rect 4791 24 4795 64
rect 4851 24 4855 104
rect 4873 24 4877 44
rect 4881 24 4885 44
rect 4901 24 4905 64
rect 4909 24 4913 64
rect 4955 24 4959 64
rect 4975 24 4979 64
rect 4987 24 4991 64
rect 5007 24 5011 64
rect 5021 24 5025 64
rect 5041 24 5045 104
rect 5110 24 5114 64
rect 5132 24 5136 104
rect 5140 24 5144 104
rect 5196 24 5200 104
rect 5204 24 5208 104
rect 5226 24 5230 64
rect 5291 24 5295 64
rect 5311 24 5315 64
rect 5371 24 5375 104
rect 5393 24 5397 44
rect 5401 24 5405 44
rect 5421 24 5425 64
rect 5429 24 5433 64
rect 5475 24 5479 64
rect 5495 24 5499 64
rect 5507 24 5511 64
rect 5527 24 5531 64
rect 5541 24 5545 64
rect 5561 24 5565 104
rect 5611 24 5615 104
rect 5633 24 5637 44
rect 5641 24 5645 44
rect 5661 24 5665 64
rect 5669 24 5673 64
rect 5715 24 5719 64
rect 5735 24 5739 64
rect 5747 24 5751 64
rect 5767 24 5771 64
rect 5781 24 5785 64
rect 5801 24 5805 104
rect 5851 24 5855 104
rect 5873 24 5877 44
rect 5881 24 5885 44
rect 5901 24 5905 64
rect 5909 24 5913 64
rect 5955 24 5959 64
rect 5975 24 5979 64
rect 5987 24 5991 64
rect 6007 24 6011 64
rect 6021 24 6025 64
rect 6041 24 6045 104
rect 6105 24 6109 104
rect 6156 24 6160 104
rect 6164 24 6168 104
rect 6186 24 6190 64
rect 6275 24 6279 104
rect 6285 24 6289 104
rect 6315 24 6319 104
rect 6325 24 6329 104
rect 6385 24 6389 64
rect 6431 24 6435 104
rect 6453 24 6457 44
rect 6461 24 6465 44
rect 6481 24 6485 64
rect 6489 24 6493 64
rect 6535 24 6539 64
rect 6555 24 6559 64
rect 6567 24 6571 64
rect 6587 24 6591 64
rect 6601 24 6605 64
rect 6621 24 6625 104
<< ndiffusion >>
rect 33 6436 35 6476
rect 39 6456 41 6476
rect 53 6456 55 6476
rect 59 6456 65 6476
rect 69 6456 73 6476
rect 85 6456 87 6476
rect 91 6456 97 6476
rect 101 6456 103 6476
rect 115 6456 119 6476
rect 123 6456 125 6476
rect 163 6456 165 6476
rect 169 6456 173 6476
rect 177 6456 179 6476
rect 191 6456 193 6476
rect 197 6456 203 6476
rect 207 6456 209 6476
rect 221 6456 225 6476
rect 39 6436 49 6456
rect 212 6436 225 6456
rect 229 6436 231 6476
rect 283 6436 285 6476
rect 289 6436 291 6476
rect 303 6436 305 6476
rect 309 6448 311 6476
rect 323 6448 325 6476
rect 309 6436 325 6448
rect 329 6436 331 6476
rect 371 6436 373 6476
rect 377 6436 383 6476
rect 387 6436 389 6476
rect 471 6436 473 6476
rect 477 6436 483 6476
rect 487 6436 489 6476
rect 531 6436 533 6476
rect 537 6436 543 6476
rect 547 6436 549 6476
rect 609 6436 611 6476
rect 615 6456 619 6476
rect 631 6456 633 6476
rect 637 6456 643 6476
rect 647 6456 649 6476
rect 661 6456 663 6476
rect 667 6456 671 6476
rect 675 6456 677 6476
rect 715 6456 717 6476
rect 721 6456 725 6476
rect 737 6456 739 6476
rect 743 6456 749 6476
rect 753 6456 755 6476
rect 767 6456 771 6476
rect 775 6456 781 6476
rect 785 6456 787 6476
rect 799 6456 801 6476
rect 615 6436 628 6456
rect 791 6436 801 6456
rect 805 6436 807 6476
rect 849 6456 851 6476
rect 855 6456 857 6476
rect 912 6436 914 6476
rect 918 6436 922 6476
rect 926 6436 928 6476
rect 940 6436 942 6476
rect 946 6436 950 6476
rect 954 6436 956 6476
rect 1043 6456 1045 6476
rect 1049 6456 1051 6476
rect 1089 6436 1091 6476
rect 1095 6456 1099 6476
rect 1111 6456 1113 6476
rect 1117 6456 1123 6476
rect 1127 6456 1129 6476
rect 1141 6456 1143 6476
rect 1147 6456 1151 6476
rect 1155 6456 1157 6476
rect 1195 6456 1197 6476
rect 1201 6456 1205 6476
rect 1217 6456 1219 6476
rect 1223 6456 1229 6476
rect 1233 6456 1235 6476
rect 1247 6456 1251 6476
rect 1255 6456 1261 6476
rect 1265 6456 1267 6476
rect 1279 6456 1281 6476
rect 1095 6436 1108 6456
rect 1271 6436 1281 6456
rect 1285 6436 1287 6476
rect 1329 6436 1331 6476
rect 1335 6446 1337 6476
rect 1349 6446 1351 6476
rect 1335 6436 1351 6446
rect 1355 6436 1357 6476
rect 1369 6436 1371 6476
rect 1375 6464 1391 6476
rect 1375 6436 1377 6464
rect 1389 6436 1391 6464
rect 1395 6436 1397 6476
rect 1463 6436 1465 6476
rect 1469 6436 1471 6476
rect 1483 6436 1485 6476
rect 1489 6448 1491 6476
rect 1503 6448 1505 6476
rect 1489 6436 1505 6448
rect 1509 6436 1511 6476
rect 1573 6436 1575 6476
rect 1579 6436 1581 6476
rect 1593 6436 1595 6476
rect 1599 6436 1605 6476
rect 1609 6436 1611 6476
rect 1663 6456 1665 6476
rect 1669 6456 1671 6476
rect 1709 6436 1711 6476
rect 1715 6456 1719 6476
rect 1731 6456 1733 6476
rect 1737 6456 1743 6476
rect 1747 6456 1749 6476
rect 1761 6456 1763 6476
rect 1767 6456 1771 6476
rect 1775 6456 1777 6476
rect 1815 6456 1817 6476
rect 1821 6456 1825 6476
rect 1837 6456 1839 6476
rect 1843 6456 1849 6476
rect 1853 6456 1855 6476
rect 1867 6456 1871 6476
rect 1875 6456 1881 6476
rect 1885 6456 1887 6476
rect 1899 6456 1901 6476
rect 1715 6436 1728 6456
rect 1891 6436 1901 6456
rect 1905 6436 1907 6476
rect 1949 6436 1951 6476
rect 1955 6448 1957 6476
rect 1969 6448 1971 6476
rect 1955 6436 1971 6448
rect 1975 6436 1977 6476
rect 1989 6436 1991 6476
rect 1995 6436 1997 6476
rect 2051 6436 2053 6476
rect 2057 6436 2063 6476
rect 2067 6436 2069 6476
rect 2143 6436 2145 6476
rect 2149 6436 2151 6476
rect 2163 6436 2165 6476
rect 2169 6448 2171 6476
rect 2183 6448 2185 6476
rect 2169 6436 2185 6448
rect 2189 6436 2191 6476
rect 2250 6456 2252 6476
rect 2256 6456 2260 6476
rect 2272 6436 2274 6476
rect 2278 6436 2282 6476
rect 2286 6436 2288 6476
rect 2351 6436 2353 6476
rect 2357 6436 2363 6476
rect 2367 6436 2369 6476
rect 2423 6456 2425 6476
rect 2429 6456 2431 6476
rect 2443 6456 2445 6476
rect 2449 6456 2451 6476
rect 2489 6456 2491 6476
rect 2495 6456 2497 6476
rect 2509 6456 2511 6476
rect 2515 6456 2517 6476
rect 2571 6436 2573 6476
rect 2577 6436 2583 6476
rect 2587 6436 2589 6476
rect 2686 6418 2688 6476
rect 2674 6416 2688 6418
rect 2692 6416 2696 6476
rect 2700 6416 2704 6476
rect 2708 6416 2710 6476
rect 2751 6436 2753 6476
rect 2757 6436 2763 6476
rect 2767 6436 2769 6476
rect 2866 6418 2868 6476
rect 2854 6416 2868 6418
rect 2872 6416 2876 6476
rect 2880 6416 2884 6476
rect 2888 6416 2890 6476
rect 2943 6436 2945 6476
rect 2949 6436 2951 6476
rect 2963 6436 2965 6476
rect 2969 6448 2971 6476
rect 2983 6448 2985 6476
rect 2969 6436 2985 6448
rect 2989 6436 2991 6476
rect 3043 6436 3045 6476
rect 3049 6436 3051 6476
rect 3063 6436 3065 6476
rect 3069 6448 3071 6476
rect 3083 6448 3085 6476
rect 3069 6436 3085 6448
rect 3089 6436 3091 6476
rect 3143 6456 3145 6476
rect 3149 6456 3151 6476
rect 3203 6456 3205 6476
rect 3209 6456 3211 6476
rect 3252 6436 3254 6476
rect 3258 6436 3262 6476
rect 3266 6436 3268 6476
rect 3280 6456 3284 6476
rect 3288 6456 3290 6476
rect 3349 6436 3351 6476
rect 3355 6448 3357 6476
rect 3369 6448 3371 6476
rect 3355 6436 3371 6448
rect 3375 6436 3377 6476
rect 3389 6436 3391 6476
rect 3395 6436 3397 6476
rect 3470 6456 3472 6476
rect 3476 6456 3480 6476
rect 3492 6436 3494 6476
rect 3498 6436 3502 6476
rect 3506 6436 3508 6476
rect 3570 6456 3572 6476
rect 3576 6456 3580 6476
rect 3592 6436 3594 6476
rect 3598 6436 3602 6476
rect 3606 6436 3608 6476
rect 3650 6416 3652 6476
rect 3656 6416 3660 6476
rect 3664 6416 3668 6476
rect 3672 6418 3674 6476
rect 3763 6436 3765 6476
rect 3769 6436 3771 6476
rect 3783 6436 3785 6476
rect 3789 6448 3791 6476
rect 3803 6448 3805 6476
rect 3789 6436 3805 6448
rect 3809 6436 3811 6476
rect 3849 6436 3851 6476
rect 3855 6448 3857 6476
rect 3869 6448 3871 6476
rect 3855 6436 3871 6448
rect 3875 6436 3877 6476
rect 3889 6436 3891 6476
rect 3895 6436 3897 6476
rect 3949 6456 3951 6476
rect 3955 6456 3957 6476
rect 3672 6416 3686 6418
rect 4011 6436 4013 6476
rect 4017 6436 4023 6476
rect 4027 6436 4029 6476
rect 4113 6436 4115 6476
rect 4119 6436 4121 6476
rect 4133 6436 4135 6476
rect 4139 6436 4145 6476
rect 4149 6436 4151 6476
rect 4191 6436 4193 6476
rect 4197 6436 4203 6476
rect 4207 6436 4209 6476
rect 4306 6418 4308 6476
rect 4294 6416 4308 6418
rect 4312 6416 4316 6476
rect 4320 6416 4324 6476
rect 4328 6416 4330 6476
rect 4406 6418 4408 6476
rect 4394 6416 4408 6418
rect 4412 6416 4416 6476
rect 4420 6416 4424 6476
rect 4428 6416 4430 6476
rect 4506 6418 4508 6476
rect 4494 6416 4508 6418
rect 4512 6416 4516 6476
rect 4520 6416 4524 6476
rect 4528 6416 4530 6476
rect 4569 6456 4571 6476
rect 4575 6456 4577 6476
rect 4632 6436 4634 6476
rect 4638 6436 4642 6476
rect 4646 6436 4648 6476
rect 4660 6456 4664 6476
rect 4668 6456 4670 6476
rect 4732 6436 4734 6476
rect 4738 6436 4742 6476
rect 4746 6436 4748 6476
rect 4760 6456 4764 6476
rect 4768 6456 4770 6476
rect 4829 6436 4831 6476
rect 4835 6448 4837 6476
rect 4849 6448 4851 6476
rect 4835 6436 4851 6448
rect 4855 6436 4857 6476
rect 4869 6436 4871 6476
rect 4875 6436 4877 6476
rect 4943 6436 4945 6476
rect 4949 6436 4951 6476
rect 4963 6436 4965 6476
rect 4969 6448 4971 6476
rect 4983 6448 4985 6476
rect 4969 6436 4985 6448
rect 4989 6436 4991 6476
rect 5029 6436 5031 6476
rect 5035 6448 5037 6476
rect 5049 6448 5051 6476
rect 5035 6436 5051 6448
rect 5055 6436 5057 6476
rect 5069 6436 5071 6476
rect 5075 6436 5077 6476
rect 5166 6418 5168 6476
rect 5154 6416 5168 6418
rect 5172 6416 5176 6476
rect 5180 6416 5184 6476
rect 5188 6416 5190 6476
rect 5266 6418 5268 6476
rect 5254 6416 5268 6418
rect 5272 6416 5276 6476
rect 5280 6416 5284 6476
rect 5288 6416 5290 6476
rect 5366 6418 5368 6476
rect 5354 6416 5368 6418
rect 5372 6416 5376 6476
rect 5380 6416 5384 6476
rect 5388 6416 5390 6476
rect 5432 6436 5434 6476
rect 5438 6436 5442 6476
rect 5446 6436 5448 6476
rect 5460 6456 5464 6476
rect 5468 6456 5470 6476
rect 5550 6456 5552 6476
rect 5556 6456 5560 6476
rect 5572 6436 5574 6476
rect 5578 6436 5582 6476
rect 5586 6436 5588 6476
rect 5643 6456 5645 6476
rect 5649 6456 5651 6476
rect 5692 6436 5694 6476
rect 5698 6436 5702 6476
rect 5706 6436 5708 6476
rect 5720 6456 5724 6476
rect 5728 6456 5730 6476
rect 5790 6416 5792 6476
rect 5796 6416 5800 6476
rect 5804 6416 5808 6476
rect 5812 6418 5814 6476
rect 5910 6456 5912 6476
rect 5916 6456 5920 6476
rect 5812 6416 5826 6418
rect 5932 6436 5934 6476
rect 5938 6436 5942 6476
rect 5946 6436 5948 6476
rect 6003 6456 6005 6476
rect 6009 6456 6011 6476
rect 6070 6456 6072 6476
rect 6076 6456 6080 6476
rect 6092 6436 6094 6476
rect 6098 6436 6102 6476
rect 6106 6436 6108 6476
rect 6163 6436 6165 6476
rect 6169 6436 6171 6476
rect 6183 6436 6185 6476
rect 6189 6448 6191 6476
rect 6203 6448 6205 6476
rect 6189 6436 6205 6448
rect 6209 6436 6211 6476
rect 6270 6456 6272 6476
rect 6276 6456 6280 6476
rect 6292 6436 6294 6476
rect 6298 6436 6302 6476
rect 6306 6436 6308 6476
rect 6350 6416 6352 6476
rect 6356 6416 6360 6476
rect 6364 6416 6368 6476
rect 6372 6418 6374 6476
rect 6372 6416 6386 6418
rect 6486 6418 6488 6476
rect 6474 6416 6488 6418
rect 6492 6416 6496 6476
rect 6500 6416 6504 6476
rect 6508 6416 6510 6476
rect 6549 6456 6551 6476
rect 6555 6456 6557 6476
rect 6612 6436 6614 6476
rect 6618 6436 6622 6476
rect 6626 6436 6628 6476
rect 6640 6436 6642 6476
rect 6646 6436 6650 6476
rect 6654 6436 6656 6476
rect 29 6024 31 6064
rect 35 6044 48 6064
rect 211 6044 221 6064
rect 35 6024 39 6044
rect 51 6024 53 6044
rect 57 6024 63 6044
rect 67 6024 69 6044
rect 81 6024 83 6044
rect 87 6024 91 6044
rect 95 6024 97 6044
rect 135 6024 137 6044
rect 141 6024 145 6044
rect 157 6024 159 6044
rect 163 6024 169 6044
rect 173 6024 175 6044
rect 187 6024 191 6044
rect 195 6024 201 6044
rect 205 6024 207 6044
rect 219 6024 221 6044
rect 225 6024 227 6064
rect 290 6024 292 6044
rect 296 6024 300 6044
rect 312 6024 314 6064
rect 318 6024 322 6064
rect 326 6024 328 6064
rect 391 6024 393 6064
rect 397 6024 403 6064
rect 407 6024 409 6064
rect 449 6024 451 6044
rect 455 6024 457 6044
rect 469 6024 471 6044
rect 475 6024 477 6044
rect 551 6024 553 6064
rect 557 6024 563 6064
rect 567 6024 569 6064
rect 609 6024 611 6064
rect 615 6052 631 6064
rect 615 6024 617 6052
rect 629 6024 631 6052
rect 635 6024 637 6064
rect 649 6024 651 6064
rect 655 6024 657 6064
rect 723 6024 725 6064
rect 729 6024 731 6064
rect 743 6024 745 6064
rect 749 6052 765 6064
rect 749 6024 751 6052
rect 763 6024 765 6052
rect 769 6024 771 6064
rect 809 6024 811 6044
rect 815 6024 817 6044
rect 829 6024 831 6044
rect 835 6024 837 6044
rect 910 6024 912 6044
rect 916 6024 920 6044
rect 932 6024 934 6064
rect 938 6024 942 6064
rect 946 6024 948 6064
rect 1019 6044 1031 6064
rect 989 6024 991 6044
rect 995 6024 997 6044
rect 1009 6024 1011 6044
rect 1015 6024 1017 6044
rect 1029 6024 1031 6044
rect 1035 6024 1037 6064
rect 1103 6024 1105 6044
rect 1109 6024 1111 6044
rect 1149 6024 1151 6044
rect 1155 6024 1157 6044
rect 1169 6024 1171 6044
rect 1175 6024 1177 6044
rect 1243 6024 1245 6064
rect 1249 6024 1251 6064
rect 1263 6024 1265 6064
rect 1269 6052 1285 6064
rect 1269 6024 1271 6052
rect 1283 6024 1285 6052
rect 1289 6024 1291 6064
rect 1343 6024 1345 6044
rect 1349 6024 1351 6044
rect 1403 6024 1405 6044
rect 1409 6024 1411 6044
rect 1449 6024 1451 6044
rect 1455 6024 1457 6044
rect 1469 6024 1471 6044
rect 1475 6024 1477 6044
rect 1529 6024 1531 6044
rect 1535 6024 1537 6044
rect 1549 6024 1551 6044
rect 1555 6024 1557 6044
rect 1609 6024 1611 6044
rect 1615 6024 1617 6044
rect 1669 6024 1671 6044
rect 1675 6024 1677 6044
rect 1689 6024 1691 6044
rect 1695 6024 1697 6044
rect 1749 6024 1751 6044
rect 1755 6024 1757 6044
rect 1769 6024 1771 6044
rect 1775 6024 1777 6044
rect 1829 6024 1831 6064
rect 1835 6052 1851 6064
rect 1835 6024 1837 6052
rect 1849 6024 1851 6052
rect 1855 6024 1857 6064
rect 1869 6024 1871 6064
rect 1875 6024 1877 6064
rect 1929 6024 1931 6044
rect 1935 6024 1937 6044
rect 2010 6024 2012 6044
rect 2016 6024 2020 6044
rect 2032 6024 2034 6064
rect 2038 6024 2042 6064
rect 2046 6024 2048 6064
rect 2089 6024 2091 6044
rect 2095 6024 2097 6044
rect 2163 6024 2165 6064
rect 2169 6024 2171 6064
rect 2183 6024 2185 6064
rect 2189 6052 2205 6064
rect 2189 6024 2191 6052
rect 2203 6024 2205 6052
rect 2209 6024 2211 6064
rect 2434 6082 2448 6084
rect 2249 6024 2251 6044
rect 2255 6024 2257 6044
rect 2323 6024 2325 6064
rect 2329 6024 2331 6064
rect 2343 6024 2345 6064
rect 2349 6052 2365 6064
rect 2349 6024 2351 6052
rect 2363 6024 2365 6052
rect 2369 6024 2371 6064
rect 2446 6024 2448 6082
rect 2452 6024 2456 6084
rect 2460 6024 2464 6084
rect 2468 6024 2470 6084
rect 2530 6024 2532 6044
rect 2536 6024 2540 6044
rect 2552 6024 2554 6064
rect 2558 6024 2562 6064
rect 2566 6024 2568 6064
rect 2714 6082 2728 6084
rect 2623 6024 2625 6044
rect 2629 6024 2631 6044
rect 2643 6024 2645 6044
rect 2649 6024 2651 6044
rect 2726 6024 2728 6082
rect 2732 6024 2736 6084
rect 2740 6024 2744 6084
rect 2748 6024 2750 6084
rect 2824 6024 2826 6064
rect 2830 6024 2834 6064
rect 2838 6024 2840 6064
rect 2852 6024 2854 6064
rect 2858 6024 2862 6064
rect 2866 6024 2868 6064
rect 2923 6024 2925 6044
rect 2929 6024 2931 6044
rect 2970 6024 2972 6084
rect 2976 6024 2980 6084
rect 2984 6024 2988 6084
rect 2992 6082 3006 6084
rect 2992 6024 2994 6082
rect 3194 6082 3208 6084
rect 3090 6024 3092 6044
rect 3096 6024 3100 6044
rect 3112 6024 3114 6064
rect 3118 6024 3122 6064
rect 3126 6024 3128 6064
rect 3206 6024 3208 6082
rect 3212 6024 3216 6084
rect 3220 6024 3224 6084
rect 3228 6024 3230 6084
rect 3290 6024 3292 6044
rect 3296 6024 3300 6044
rect 3312 6024 3314 6064
rect 3318 6024 3322 6064
rect 3326 6024 3328 6064
rect 3454 6082 3468 6084
rect 3383 6024 3385 6044
rect 3389 6024 3391 6044
rect 3466 6024 3468 6082
rect 3472 6024 3476 6084
rect 3480 6024 3484 6084
rect 3488 6024 3490 6084
rect 3530 6024 3532 6084
rect 3536 6024 3540 6084
rect 3544 6024 3548 6084
rect 3552 6082 3566 6084
rect 3552 6024 3554 6082
rect 3629 6024 3631 6044
rect 3635 6024 3637 6044
rect 3692 6024 3694 6064
rect 3698 6024 3702 6064
rect 3706 6024 3708 6064
rect 3720 6024 3724 6044
rect 3728 6024 3730 6044
rect 3811 6024 3813 6064
rect 3817 6024 3823 6064
rect 3827 6024 3829 6064
rect 3871 6024 3873 6064
rect 3877 6024 3883 6064
rect 3887 6024 3889 6064
rect 3963 6024 3965 6064
rect 3969 6024 3971 6064
rect 3983 6024 3985 6064
rect 3989 6052 4005 6064
rect 3989 6024 3991 6052
rect 4003 6024 4005 6052
rect 4009 6024 4011 6064
rect 4049 6024 4051 6064
rect 4055 6052 4071 6064
rect 4055 6024 4057 6052
rect 4069 6024 4071 6052
rect 4075 6024 4077 6064
rect 4089 6024 4091 6064
rect 4095 6024 4097 6064
rect 4163 6024 4165 6044
rect 4169 6024 4171 6044
rect 4183 6024 4185 6044
rect 4189 6024 4191 6044
rect 4229 6024 4231 6044
rect 4235 6024 4237 6044
rect 4311 6024 4313 6064
rect 4317 6024 4323 6064
rect 4327 6024 4329 6064
rect 4369 6024 4371 6064
rect 4375 6024 4381 6064
rect 4385 6024 4387 6064
rect 4399 6024 4401 6064
rect 4405 6024 4407 6064
rect 4483 6024 4485 6064
rect 4489 6024 4491 6064
rect 4503 6024 4505 6064
rect 4509 6052 4525 6064
rect 4509 6024 4511 6052
rect 4523 6024 4525 6052
rect 4529 6024 4531 6064
rect 4590 6024 4592 6044
rect 4596 6024 4600 6044
rect 4612 6024 4614 6064
rect 4618 6024 4622 6064
rect 4626 6024 4628 6064
rect 4670 6024 4672 6084
rect 4676 6024 4680 6084
rect 4684 6024 4688 6084
rect 4692 6082 4706 6084
rect 4692 6024 4694 6082
rect 4894 6082 4908 6084
rect 4790 6024 4792 6044
rect 4796 6024 4800 6044
rect 4812 6024 4814 6064
rect 4818 6024 4822 6064
rect 4826 6024 4828 6064
rect 4906 6024 4908 6082
rect 4912 6024 4916 6084
rect 4920 6024 4924 6084
rect 4928 6024 4930 6084
rect 4970 6024 4972 6084
rect 4976 6024 4980 6084
rect 4984 6024 4988 6084
rect 4992 6082 5006 6084
rect 4992 6024 4994 6082
rect 5083 6024 5085 6064
rect 5089 6024 5091 6064
rect 5103 6024 5105 6064
rect 5109 6052 5125 6064
rect 5109 6024 5111 6052
rect 5123 6024 5125 6052
rect 5129 6024 5131 6064
rect 5191 6024 5193 6064
rect 5197 6024 5203 6064
rect 5207 6024 5209 6064
rect 5249 6024 5251 6064
rect 5255 6024 5261 6064
rect 5265 6024 5267 6064
rect 5279 6024 5281 6064
rect 5285 6024 5287 6064
rect 5349 6024 5351 6064
rect 5355 6052 5371 6064
rect 5355 6024 5357 6052
rect 5369 6024 5371 6052
rect 5375 6024 5377 6064
rect 5389 6024 5391 6064
rect 5395 6024 5397 6064
rect 5574 6082 5588 6084
rect 5470 6024 5472 6044
rect 5476 6024 5480 6044
rect 5492 6024 5494 6064
rect 5498 6024 5502 6064
rect 5506 6024 5508 6064
rect 5586 6024 5588 6082
rect 5592 6024 5596 6084
rect 5600 6024 5604 6084
rect 5608 6024 5610 6084
rect 5650 6024 5652 6084
rect 5656 6024 5660 6084
rect 5664 6024 5668 6084
rect 5672 6082 5686 6084
rect 5672 6024 5674 6082
rect 5770 6024 5772 6044
rect 5776 6024 5780 6044
rect 5792 6024 5794 6064
rect 5798 6024 5802 6064
rect 5806 6024 5808 6064
rect 5850 6024 5852 6084
rect 5856 6024 5860 6084
rect 5864 6024 5868 6084
rect 5872 6082 5886 6084
rect 5872 6024 5874 6082
rect 5949 6024 5951 6064
rect 5955 6052 5971 6064
rect 5955 6024 5957 6052
rect 5969 6024 5971 6052
rect 5975 6024 5977 6064
rect 5989 6024 5991 6064
rect 5995 6024 5997 6064
rect 6049 6024 6051 6064
rect 6055 6052 6071 6064
rect 6055 6024 6057 6052
rect 6069 6024 6071 6052
rect 6075 6024 6077 6064
rect 6089 6024 6091 6064
rect 6095 6024 6097 6064
rect 6150 6024 6152 6084
rect 6156 6024 6160 6084
rect 6164 6024 6168 6084
rect 6172 6082 6186 6084
rect 6172 6024 6174 6082
rect 6250 6024 6252 6084
rect 6256 6024 6260 6084
rect 6264 6024 6268 6084
rect 6272 6082 6286 6084
rect 6272 6024 6274 6082
rect 6374 6082 6388 6084
rect 6386 6024 6388 6082
rect 6392 6024 6396 6084
rect 6400 6024 6404 6084
rect 6408 6024 6410 6084
rect 6470 6024 6472 6044
rect 6476 6024 6480 6044
rect 6492 6024 6494 6064
rect 6498 6024 6502 6064
rect 6506 6024 6508 6064
rect 6549 6024 6551 6044
rect 6555 6024 6557 6044
rect 6609 6024 6611 6044
rect 6615 6024 6617 6044
rect 41 5956 43 5996
rect 47 5956 49 5996
rect 61 5976 65 5996
rect 69 5976 71 5996
rect 111 5956 113 5996
rect 117 5956 123 5996
rect 127 5956 129 5996
rect 191 5956 193 5996
rect 197 5956 203 5996
rect 207 5956 209 5996
rect 290 5976 292 5996
rect 296 5976 300 5996
rect 312 5956 314 5996
rect 318 5956 322 5996
rect 326 5956 328 5996
rect 391 5956 393 5996
rect 397 5956 403 5996
rect 407 5956 409 5996
rect 449 5976 451 5996
rect 455 5976 457 5996
rect 523 5976 525 5996
rect 529 5976 531 5996
rect 543 5976 545 5996
rect 549 5976 551 5996
rect 589 5976 591 5996
rect 595 5976 597 5996
rect 609 5976 611 5996
rect 615 5976 617 5996
rect 669 5956 671 5996
rect 675 5968 677 5996
rect 689 5968 691 5996
rect 675 5956 691 5968
rect 695 5956 697 5996
rect 709 5956 711 5996
rect 715 5956 717 5996
rect 783 5976 785 5996
rect 789 5976 791 5996
rect 829 5976 831 5996
rect 835 5976 837 5996
rect 849 5976 851 5996
rect 855 5976 857 5996
rect 931 5956 933 5996
rect 937 5956 943 5996
rect 947 5956 949 5996
rect 1003 5956 1005 5996
rect 1009 5956 1011 5996
rect 1023 5956 1025 5996
rect 1029 5968 1031 5996
rect 1043 5968 1045 5996
rect 1029 5956 1045 5968
rect 1049 5956 1051 5996
rect 1089 5976 1091 5996
rect 1095 5976 1097 5996
rect 1109 5976 1111 5996
rect 1115 5976 1117 5996
rect 1183 5976 1185 5996
rect 1189 5976 1191 5996
rect 1229 5956 1231 5996
rect 1235 5976 1239 5996
rect 1251 5976 1253 5996
rect 1257 5976 1263 5996
rect 1267 5976 1269 5996
rect 1281 5976 1283 5996
rect 1287 5976 1291 5996
rect 1295 5976 1297 5996
rect 1335 5976 1337 5996
rect 1341 5976 1345 5996
rect 1357 5976 1359 5996
rect 1363 5976 1369 5996
rect 1373 5976 1375 5996
rect 1387 5976 1391 5996
rect 1395 5976 1401 5996
rect 1405 5976 1407 5996
rect 1419 5976 1421 5996
rect 1235 5956 1248 5976
rect 1411 5956 1421 5976
rect 1425 5956 1427 5996
rect 1471 5956 1473 5996
rect 1477 5956 1483 5996
rect 1487 5956 1489 5996
rect 1586 5938 1588 5996
rect 1574 5936 1588 5938
rect 1592 5936 1596 5996
rect 1600 5936 1604 5996
rect 1608 5936 1610 5996
rect 1663 5956 1665 5996
rect 1669 5956 1671 5996
rect 1683 5956 1685 5996
rect 1689 5968 1691 5996
rect 1703 5968 1705 5996
rect 1689 5956 1705 5968
rect 1709 5956 1711 5996
rect 1763 5976 1765 5996
rect 1769 5976 1771 5996
rect 1783 5976 1785 5996
rect 1789 5976 1791 5996
rect 1866 5938 1868 5996
rect 1854 5936 1868 5938
rect 1872 5936 1876 5996
rect 1880 5936 1884 5996
rect 1888 5936 1890 5996
rect 1929 5976 1931 5996
rect 1935 5976 1937 5996
rect 2003 5956 2005 5996
rect 2009 5956 2011 5996
rect 2023 5956 2025 5996
rect 2029 5968 2031 5996
rect 2043 5968 2045 5996
rect 2029 5956 2045 5968
rect 2049 5956 2051 5996
rect 2090 5936 2092 5996
rect 2096 5936 2100 5996
rect 2104 5936 2108 5996
rect 2112 5938 2114 5996
rect 2210 5976 2212 5996
rect 2216 5976 2220 5996
rect 2112 5936 2126 5938
rect 2232 5956 2234 5996
rect 2238 5956 2242 5996
rect 2246 5956 2248 5996
rect 2289 5956 2291 5996
rect 2295 5968 2297 5996
rect 2309 5968 2311 5996
rect 2295 5956 2311 5968
rect 2315 5956 2317 5996
rect 2329 5956 2331 5996
rect 2335 5956 2337 5996
rect 2411 5956 2413 5996
rect 2417 5956 2423 5996
rect 2427 5956 2429 5996
rect 2506 5938 2508 5996
rect 2494 5936 2508 5938
rect 2512 5936 2516 5996
rect 2520 5936 2524 5996
rect 2528 5936 2530 5996
rect 2590 5976 2592 5996
rect 2596 5976 2600 5996
rect 2612 5956 2614 5996
rect 2618 5956 2622 5996
rect 2626 5956 2628 5996
rect 2671 5956 2673 5996
rect 2677 5956 2683 5996
rect 2687 5956 2689 5996
rect 2786 5938 2788 5996
rect 2774 5936 2788 5938
rect 2792 5936 2796 5996
rect 2800 5936 2804 5996
rect 2808 5936 2810 5996
rect 2886 5938 2888 5996
rect 2874 5936 2888 5938
rect 2892 5936 2896 5996
rect 2900 5936 2904 5996
rect 2908 5936 2910 5996
rect 2986 5938 2988 5996
rect 2974 5936 2988 5938
rect 2992 5936 2996 5996
rect 3000 5936 3004 5996
rect 3008 5936 3010 5996
rect 3086 5938 3088 5996
rect 3074 5936 3088 5938
rect 3092 5936 3096 5996
rect 3100 5936 3104 5996
rect 3108 5936 3110 5996
rect 3150 5936 3152 5996
rect 3156 5936 3160 5996
rect 3164 5936 3168 5996
rect 3172 5938 3174 5996
rect 3263 5956 3265 5996
rect 3269 5956 3271 5996
rect 3283 5956 3285 5996
rect 3289 5968 3291 5996
rect 3303 5968 3305 5996
rect 3289 5956 3305 5968
rect 3309 5956 3311 5996
rect 3349 5956 3351 5996
rect 3355 5968 3357 5996
rect 3369 5968 3371 5996
rect 3355 5956 3371 5968
rect 3375 5956 3377 5996
rect 3389 5956 3391 5996
rect 3395 5956 3397 5996
rect 3470 5976 3472 5996
rect 3476 5976 3480 5996
rect 3172 5936 3186 5938
rect 3492 5956 3494 5996
rect 3498 5956 3502 5996
rect 3506 5956 3508 5996
rect 3563 5956 3565 5996
rect 3569 5956 3571 5996
rect 3583 5956 3585 5996
rect 3589 5968 3591 5996
rect 3603 5968 3605 5996
rect 3589 5956 3605 5968
rect 3609 5956 3611 5996
rect 3686 5938 3688 5996
rect 3674 5936 3688 5938
rect 3692 5936 3696 5996
rect 3700 5936 3704 5996
rect 3708 5936 3710 5996
rect 3752 5956 3754 5996
rect 3758 5956 3762 5996
rect 3766 5956 3768 5996
rect 3780 5976 3784 5996
rect 3788 5976 3790 5996
rect 3886 5938 3888 5996
rect 3874 5936 3888 5938
rect 3892 5936 3896 5996
rect 3900 5936 3904 5996
rect 3908 5936 3910 5996
rect 3970 5976 3972 5996
rect 3976 5976 3980 5996
rect 3992 5956 3994 5996
rect 3998 5956 4002 5996
rect 4006 5956 4008 5996
rect 4086 5938 4088 5996
rect 4074 5936 4088 5938
rect 4092 5936 4096 5996
rect 4100 5936 4104 5996
rect 4108 5936 4110 5996
rect 4170 5976 4172 5996
rect 4176 5976 4180 5996
rect 4192 5956 4194 5996
rect 4198 5956 4202 5996
rect 4206 5956 4208 5996
rect 4250 5936 4252 5996
rect 4256 5936 4260 5996
rect 4264 5936 4268 5996
rect 4272 5938 4274 5996
rect 4351 5956 4353 5996
rect 4357 5956 4363 5996
rect 4367 5956 4369 5996
rect 4443 5956 4445 5996
rect 4449 5956 4451 5996
rect 4463 5956 4465 5996
rect 4469 5968 4471 5996
rect 4483 5968 4485 5996
rect 4469 5956 4485 5968
rect 4489 5956 4491 5996
rect 4543 5976 4545 5996
rect 4549 5976 4551 5996
rect 4563 5976 4565 5996
rect 4569 5976 4571 5996
rect 4272 5936 4286 5938
rect 4609 5956 4611 5996
rect 4615 5956 4621 5996
rect 4625 5956 4627 5996
rect 4639 5956 4641 5996
rect 4645 5956 4647 5996
rect 4730 5976 4732 5996
rect 4736 5976 4740 5996
rect 4752 5956 4754 5996
rect 4758 5956 4762 5996
rect 4766 5956 4768 5996
rect 4811 5956 4813 5996
rect 4817 5956 4823 5996
rect 4827 5956 4829 5996
rect 4903 5976 4905 5996
rect 4909 5976 4911 5996
rect 4986 5938 4988 5996
rect 4974 5936 4988 5938
rect 4992 5936 4996 5996
rect 5000 5936 5004 5996
rect 5008 5936 5010 5996
rect 5052 5956 5054 5996
rect 5058 5956 5062 5996
rect 5066 5956 5068 5996
rect 5080 5976 5084 5996
rect 5088 5976 5090 5996
rect 5149 5956 5151 5996
rect 5155 5968 5157 5996
rect 5169 5968 5171 5996
rect 5155 5956 5171 5968
rect 5175 5956 5177 5996
rect 5189 5956 5191 5996
rect 5195 5956 5197 5996
rect 5249 5956 5251 5996
rect 5255 5968 5257 5996
rect 5269 5968 5271 5996
rect 5255 5956 5271 5968
rect 5275 5956 5277 5996
rect 5289 5956 5291 5996
rect 5295 5956 5297 5996
rect 5352 5956 5354 5996
rect 5358 5956 5362 5996
rect 5366 5956 5368 5996
rect 5380 5956 5382 5996
rect 5386 5956 5390 5996
rect 5394 5956 5396 5996
rect 5491 5956 5493 5996
rect 5497 5956 5503 5996
rect 5507 5956 5509 5996
rect 5549 5976 5551 5996
rect 5555 5976 5557 5996
rect 5646 5938 5648 5996
rect 5634 5936 5648 5938
rect 5652 5936 5656 5996
rect 5660 5936 5664 5996
rect 5668 5936 5670 5996
rect 5712 5956 5714 5996
rect 5718 5956 5722 5996
rect 5726 5956 5728 5996
rect 5740 5976 5744 5996
rect 5748 5976 5750 5996
rect 5823 5956 5825 5996
rect 5829 5956 5831 5996
rect 5843 5956 5845 5996
rect 5849 5968 5851 5996
rect 5863 5968 5865 5996
rect 5849 5956 5865 5968
rect 5869 5956 5871 5996
rect 5909 5956 5911 5996
rect 5915 5968 5917 5996
rect 5929 5968 5931 5996
rect 5915 5956 5931 5968
rect 5935 5956 5937 5996
rect 5949 5956 5951 5996
rect 5955 5956 5957 5996
rect 6023 5956 6025 5996
rect 6029 5956 6031 5996
rect 6043 5956 6045 5996
rect 6049 5968 6051 5996
rect 6063 5968 6065 5996
rect 6049 5956 6065 5968
rect 6069 5956 6071 5996
rect 6112 5956 6114 5996
rect 6118 5956 6122 5996
rect 6126 5956 6128 5996
rect 6140 5956 6142 5996
rect 6146 5956 6150 5996
rect 6154 5956 6156 5996
rect 6251 5956 6253 5996
rect 6257 5956 6263 5996
rect 6267 5956 6269 5996
rect 6309 5956 6311 5996
rect 6315 5956 6321 5996
rect 6325 5956 6327 5996
rect 6339 5956 6341 5996
rect 6345 5956 6347 5996
rect 6409 5956 6411 5996
rect 6415 5968 6417 5996
rect 6429 5968 6431 5996
rect 6415 5956 6431 5968
rect 6435 5956 6437 5996
rect 6449 5956 6451 5996
rect 6455 5956 6457 5996
rect 6510 5936 6512 5996
rect 6516 5936 6520 5996
rect 6524 5936 6528 5996
rect 6532 5938 6534 5996
rect 6611 5956 6613 5996
rect 6617 5956 6623 5996
rect 6627 5956 6629 5996
rect 6532 5936 6546 5938
rect 41 5544 43 5584
rect 47 5544 49 5584
rect 61 5544 65 5564
rect 69 5544 71 5564
rect 121 5544 123 5584
rect 127 5544 129 5584
rect 141 5544 145 5564
rect 149 5544 151 5564
rect 189 5544 191 5584
rect 195 5564 208 5584
rect 371 5564 381 5584
rect 195 5544 199 5564
rect 211 5544 213 5564
rect 217 5544 223 5564
rect 227 5544 229 5564
rect 241 5544 243 5564
rect 247 5544 251 5564
rect 255 5544 257 5564
rect 295 5544 297 5564
rect 301 5544 305 5564
rect 317 5544 319 5564
rect 323 5544 329 5564
rect 333 5544 335 5564
rect 347 5544 351 5564
rect 355 5544 361 5564
rect 365 5544 367 5564
rect 379 5544 381 5564
rect 385 5544 387 5584
rect 443 5544 445 5564
rect 449 5544 451 5564
rect 463 5544 465 5564
rect 469 5544 471 5564
rect 512 5544 514 5584
rect 518 5544 522 5584
rect 526 5544 528 5584
rect 540 5544 544 5564
rect 548 5544 550 5564
rect 611 5544 613 5584
rect 617 5544 623 5584
rect 627 5544 629 5584
rect 689 5544 691 5584
rect 695 5544 701 5584
rect 705 5544 707 5584
rect 719 5544 721 5584
rect 725 5544 727 5584
rect 791 5544 793 5584
rect 797 5544 803 5584
rect 807 5544 809 5584
rect 871 5544 873 5584
rect 877 5544 883 5584
rect 887 5544 889 5584
rect 1119 5564 1131 5584
rect 949 5544 951 5564
rect 955 5544 957 5564
rect 969 5544 971 5564
rect 975 5544 977 5564
rect 1029 5544 1031 5564
rect 1035 5544 1037 5564
rect 1089 5544 1091 5564
rect 1095 5544 1097 5564
rect 1109 5544 1111 5564
rect 1115 5544 1117 5564
rect 1129 5544 1131 5564
rect 1135 5544 1137 5584
rect 1189 5544 1191 5564
rect 1195 5544 1197 5564
rect 1209 5544 1211 5564
rect 1215 5544 1217 5564
rect 1269 5544 1271 5564
rect 1275 5544 1277 5564
rect 1329 5544 1331 5564
rect 1335 5544 1337 5564
rect 1349 5544 1351 5564
rect 1355 5544 1357 5564
rect 1409 5544 1411 5564
rect 1415 5544 1417 5564
rect 1469 5544 1471 5584
rect 1475 5564 1488 5584
rect 1651 5564 1661 5584
rect 1475 5544 1479 5564
rect 1491 5544 1493 5564
rect 1497 5544 1503 5564
rect 1507 5544 1509 5564
rect 1521 5544 1523 5564
rect 1527 5544 1531 5564
rect 1535 5544 1537 5564
rect 1575 5544 1577 5564
rect 1581 5544 1585 5564
rect 1597 5544 1599 5564
rect 1603 5544 1609 5564
rect 1613 5544 1615 5564
rect 1627 5544 1631 5564
rect 1635 5544 1641 5564
rect 1645 5544 1647 5564
rect 1659 5544 1661 5564
rect 1665 5544 1667 5584
rect 1709 5544 1711 5584
rect 1715 5574 1731 5584
rect 1715 5544 1717 5574
rect 1729 5544 1731 5574
rect 1735 5544 1737 5584
rect 1749 5544 1751 5584
rect 1755 5556 1757 5584
rect 1769 5556 1771 5584
rect 1755 5544 1771 5556
rect 1775 5544 1777 5584
rect 1843 5544 1845 5584
rect 1849 5544 1851 5584
rect 1863 5544 1865 5584
rect 1869 5572 1885 5584
rect 1869 5544 1871 5572
rect 1883 5544 1885 5572
rect 1889 5544 1891 5584
rect 1951 5544 1953 5584
rect 1957 5544 1963 5584
rect 1967 5544 1969 5584
rect 2009 5544 2011 5564
rect 2015 5544 2017 5564
rect 2090 5544 2092 5564
rect 2096 5544 2100 5564
rect 2112 5544 2114 5584
rect 2118 5544 2122 5584
rect 2126 5544 2128 5584
rect 2169 5544 2171 5564
rect 2175 5544 2177 5564
rect 2189 5544 2191 5564
rect 2195 5544 2197 5564
rect 2251 5544 2253 5584
rect 2257 5544 2263 5584
rect 2267 5544 2269 5584
rect 2614 5602 2628 5604
rect 2403 5544 2405 5564
rect 2409 5544 2411 5564
rect 2423 5544 2425 5564
rect 2429 5544 2431 5564
rect 2443 5544 2445 5564
rect 2449 5544 2451 5564
rect 2531 5544 2533 5584
rect 2537 5544 2543 5584
rect 2547 5544 2549 5584
rect 2626 5544 2628 5602
rect 2632 5544 2636 5604
rect 2640 5544 2644 5604
rect 2648 5544 2650 5604
rect 2714 5602 2728 5604
rect 2726 5544 2728 5602
rect 2732 5544 2736 5604
rect 2740 5544 2744 5604
rect 2748 5544 2750 5604
rect 2994 5602 3008 5604
rect 2791 5544 2793 5584
rect 2797 5544 2803 5584
rect 2807 5544 2809 5584
rect 2869 5544 2871 5584
rect 2875 5572 2891 5584
rect 2875 5544 2877 5572
rect 2889 5544 2891 5572
rect 2895 5544 2897 5584
rect 2909 5544 2911 5584
rect 2915 5544 2917 5584
rect 3006 5544 3008 5602
rect 3012 5544 3016 5604
rect 3020 5544 3024 5604
rect 3028 5544 3030 5604
rect 3072 5544 3074 5584
rect 3078 5544 3082 5584
rect 3086 5544 3088 5584
rect 3100 5544 3104 5564
rect 3108 5544 3110 5564
rect 3183 5544 3185 5584
rect 3189 5544 3191 5584
rect 3203 5544 3205 5584
rect 3209 5572 3225 5584
rect 3209 5544 3211 5572
rect 3223 5544 3225 5572
rect 3229 5544 3231 5584
rect 3283 5544 3285 5564
rect 3289 5544 3291 5564
rect 3330 5544 3332 5604
rect 3336 5544 3340 5604
rect 3344 5544 3348 5604
rect 3352 5602 3366 5604
rect 3352 5544 3354 5602
rect 3454 5602 3468 5604
rect 3466 5544 3468 5602
rect 3472 5544 3476 5604
rect 3480 5544 3484 5604
rect 3488 5544 3490 5604
rect 3554 5602 3568 5604
rect 3566 5544 3568 5602
rect 3572 5544 3576 5604
rect 3580 5544 3584 5604
rect 3588 5544 3590 5604
rect 3643 5544 3645 5564
rect 3649 5544 3651 5564
rect 3703 5544 3705 5584
rect 3709 5544 3711 5584
rect 3723 5544 3725 5584
rect 3729 5572 3745 5584
rect 3729 5544 3731 5572
rect 3743 5544 3745 5572
rect 3749 5544 3751 5584
rect 3803 5544 3805 5564
rect 3809 5544 3811 5564
rect 3823 5544 3825 5564
rect 3829 5544 3831 5564
rect 3869 5544 3871 5584
rect 3875 5572 3891 5584
rect 3875 5544 3877 5572
rect 3889 5544 3891 5572
rect 3895 5544 3897 5584
rect 3909 5544 3911 5584
rect 3915 5544 3917 5584
rect 4274 5602 4288 5604
rect 3983 5544 3985 5564
rect 3989 5544 3991 5564
rect 4064 5544 4066 5584
rect 4070 5544 4074 5584
rect 4078 5544 4080 5584
rect 4092 5544 4094 5584
rect 4098 5544 4102 5584
rect 4106 5544 4108 5584
rect 4163 5544 4165 5584
rect 4169 5544 4171 5584
rect 4183 5544 4185 5584
rect 4189 5572 4205 5584
rect 4189 5544 4191 5572
rect 4203 5544 4205 5572
rect 4209 5544 4211 5584
rect 4286 5544 4288 5602
rect 4292 5544 4296 5604
rect 4300 5544 4304 5604
rect 4308 5544 4310 5604
rect 4914 5602 4928 5604
rect 4349 5544 4351 5564
rect 4355 5544 4357 5564
rect 4423 5544 4425 5584
rect 4429 5544 4431 5584
rect 4443 5544 4445 5584
rect 4449 5572 4465 5584
rect 4449 5544 4451 5572
rect 4463 5544 4465 5572
rect 4469 5544 4471 5584
rect 4533 5544 4535 5584
rect 4539 5544 4541 5584
rect 4553 5544 4555 5584
rect 4559 5544 4565 5584
rect 4569 5544 4571 5584
rect 4611 5544 4613 5584
rect 4617 5544 4623 5584
rect 4627 5544 4629 5584
rect 4703 5544 4705 5584
rect 4709 5544 4711 5584
rect 4723 5544 4725 5584
rect 4729 5572 4745 5584
rect 4729 5544 4731 5572
rect 4743 5544 4745 5572
rect 4749 5544 4751 5584
rect 4789 5544 4791 5584
rect 4795 5572 4811 5584
rect 4795 5544 4797 5572
rect 4809 5544 4811 5572
rect 4815 5544 4817 5584
rect 4829 5544 4831 5584
rect 4835 5544 4837 5584
rect 4926 5544 4928 5602
rect 4932 5544 4936 5604
rect 4940 5544 4944 5604
rect 4948 5544 4950 5604
rect 4992 5544 4994 5584
rect 4998 5544 5002 5584
rect 5006 5544 5008 5584
rect 5020 5544 5024 5564
rect 5028 5544 5030 5564
rect 5089 5544 5091 5584
rect 5095 5572 5111 5584
rect 5095 5544 5097 5572
rect 5109 5544 5111 5572
rect 5115 5544 5117 5584
rect 5129 5544 5131 5584
rect 5135 5544 5137 5584
rect 5190 5544 5192 5604
rect 5196 5544 5200 5604
rect 5204 5544 5208 5604
rect 5212 5602 5226 5604
rect 5212 5544 5214 5602
rect 5291 5544 5293 5584
rect 5297 5544 5303 5584
rect 5307 5544 5309 5584
rect 5370 5544 5372 5604
rect 5376 5544 5380 5604
rect 5384 5544 5388 5604
rect 5392 5602 5406 5604
rect 5392 5544 5394 5602
rect 5472 5544 5474 5584
rect 5478 5544 5482 5584
rect 5486 5544 5488 5584
rect 5500 5544 5504 5564
rect 5508 5544 5510 5564
rect 5571 5544 5573 5584
rect 5577 5544 5583 5584
rect 5587 5544 5589 5584
rect 5671 5544 5673 5584
rect 5677 5544 5683 5584
rect 5687 5544 5689 5584
rect 5732 5544 5734 5584
rect 5738 5544 5742 5584
rect 5746 5544 5748 5584
rect 5760 5544 5762 5584
rect 5766 5544 5770 5584
rect 5774 5544 5776 5584
rect 5863 5544 5865 5584
rect 5869 5544 5871 5584
rect 5883 5544 5885 5584
rect 5889 5572 5905 5584
rect 5889 5544 5891 5572
rect 5903 5544 5905 5572
rect 5909 5544 5911 5584
rect 5949 5544 5951 5564
rect 5955 5544 5957 5564
rect 6012 5544 6014 5584
rect 6018 5544 6022 5584
rect 6026 5544 6028 5584
rect 6040 5544 6042 5584
rect 6046 5544 6050 5584
rect 6054 5544 6056 5584
rect 6130 5544 6132 5604
rect 6136 5544 6140 5604
rect 6144 5544 6148 5604
rect 6152 5602 6166 5604
rect 6152 5544 6154 5602
rect 6243 5544 6245 5564
rect 6249 5544 6251 5564
rect 6292 5544 6294 5584
rect 6298 5544 6302 5584
rect 6306 5544 6308 5584
rect 6320 5544 6324 5564
rect 6328 5544 6330 5564
rect 6390 5544 6392 5604
rect 6396 5544 6400 5604
rect 6404 5544 6408 5604
rect 6412 5602 6426 5604
rect 6412 5544 6414 5602
rect 6490 5544 6492 5604
rect 6496 5544 6500 5604
rect 6504 5544 6508 5604
rect 6512 5602 6526 5604
rect 6512 5544 6514 5602
rect 6590 5544 6592 5604
rect 6596 5544 6600 5604
rect 6604 5544 6608 5604
rect 6612 5602 6626 5604
rect 6612 5544 6614 5602
rect 29 5476 31 5516
rect 35 5496 39 5516
rect 51 5496 53 5516
rect 57 5496 63 5516
rect 67 5496 69 5516
rect 81 5496 83 5516
rect 87 5496 91 5516
rect 95 5496 97 5516
rect 135 5496 137 5516
rect 141 5496 145 5516
rect 157 5496 159 5516
rect 163 5496 169 5516
rect 173 5496 175 5516
rect 187 5496 191 5516
rect 195 5496 201 5516
rect 205 5496 207 5516
rect 219 5496 221 5516
rect 35 5476 48 5496
rect 211 5476 221 5496
rect 225 5476 227 5516
rect 271 5476 273 5516
rect 277 5476 283 5516
rect 287 5476 289 5516
rect 370 5496 372 5516
rect 376 5496 380 5516
rect 392 5476 394 5516
rect 398 5476 402 5516
rect 406 5476 408 5516
rect 471 5476 473 5516
rect 477 5476 483 5516
rect 487 5476 489 5516
rect 553 5476 555 5516
rect 559 5476 561 5516
rect 573 5476 575 5516
rect 579 5476 585 5516
rect 589 5476 591 5516
rect 629 5496 631 5516
rect 635 5496 637 5516
rect 649 5496 651 5516
rect 655 5496 657 5516
rect 709 5496 711 5516
rect 715 5496 717 5516
rect 729 5496 731 5516
rect 735 5496 737 5516
rect 791 5476 793 5516
rect 797 5476 803 5516
rect 807 5476 809 5516
rect 871 5476 873 5516
rect 877 5476 883 5516
rect 887 5476 889 5516
rect 949 5496 951 5516
rect 955 5496 957 5516
rect 1012 5476 1014 5516
rect 1018 5476 1022 5516
rect 1026 5476 1028 5516
rect 1040 5496 1044 5516
rect 1048 5496 1050 5516
rect 1144 5476 1146 5516
rect 1150 5476 1154 5516
rect 1158 5476 1160 5516
rect 1172 5476 1174 5516
rect 1178 5476 1182 5516
rect 1186 5476 1188 5516
rect 1229 5476 1231 5516
rect 1235 5496 1239 5516
rect 1251 5496 1253 5516
rect 1257 5496 1263 5516
rect 1267 5496 1269 5516
rect 1281 5496 1283 5516
rect 1287 5496 1291 5516
rect 1295 5496 1297 5516
rect 1335 5496 1337 5516
rect 1341 5496 1345 5516
rect 1357 5496 1359 5516
rect 1363 5496 1369 5516
rect 1373 5496 1375 5516
rect 1387 5496 1391 5516
rect 1395 5496 1401 5516
rect 1405 5496 1407 5516
rect 1419 5496 1421 5516
rect 1235 5476 1248 5496
rect 1411 5476 1421 5496
rect 1425 5476 1427 5516
rect 1506 5458 1508 5516
rect 1494 5456 1508 5458
rect 1512 5456 1516 5516
rect 1520 5456 1524 5516
rect 1528 5456 1530 5516
rect 1606 5458 1608 5516
rect 1594 5456 1608 5458
rect 1612 5456 1616 5516
rect 1620 5456 1624 5516
rect 1628 5456 1630 5516
rect 1683 5496 1685 5516
rect 1689 5496 1691 5516
rect 1743 5476 1745 5516
rect 1749 5476 1751 5516
rect 1763 5476 1765 5516
rect 1769 5488 1771 5516
rect 1783 5488 1785 5516
rect 1769 5476 1785 5488
rect 1789 5476 1791 5516
rect 1853 5476 1855 5516
rect 1859 5476 1861 5516
rect 1873 5476 1875 5516
rect 1879 5476 1885 5516
rect 1889 5476 1891 5516
rect 1951 5476 1953 5516
rect 1957 5476 1963 5516
rect 1967 5476 1969 5516
rect 2023 5476 2025 5516
rect 2029 5476 2031 5516
rect 2043 5476 2045 5516
rect 2049 5488 2051 5516
rect 2063 5488 2065 5516
rect 2049 5476 2065 5488
rect 2069 5476 2071 5516
rect 2111 5476 2113 5516
rect 2117 5476 2123 5516
rect 2127 5476 2129 5516
rect 2203 5496 2205 5516
rect 2209 5496 2211 5516
rect 2263 5476 2265 5516
rect 2269 5476 2271 5516
rect 2283 5476 2285 5516
rect 2289 5488 2291 5516
rect 2303 5488 2305 5516
rect 2289 5476 2305 5488
rect 2309 5476 2311 5516
rect 2349 5496 2351 5516
rect 2355 5496 2357 5516
rect 2369 5496 2371 5516
rect 2375 5496 2377 5516
rect 2443 5496 2445 5516
rect 2449 5496 2451 5516
rect 2510 5496 2512 5516
rect 2516 5496 2520 5516
rect 2532 5476 2534 5516
rect 2538 5476 2542 5516
rect 2546 5476 2548 5516
rect 2589 5476 2591 5516
rect 2595 5488 2597 5516
rect 2609 5488 2611 5516
rect 2595 5476 2611 5488
rect 2615 5476 2617 5516
rect 2629 5476 2631 5516
rect 2635 5476 2637 5516
rect 2691 5476 2693 5516
rect 2697 5476 2703 5516
rect 2707 5476 2709 5516
rect 2806 5458 2808 5516
rect 2794 5456 2808 5458
rect 2812 5456 2816 5516
rect 2820 5456 2824 5516
rect 2828 5456 2830 5516
rect 2891 5476 2893 5516
rect 2897 5476 2903 5516
rect 2907 5476 2909 5516
rect 2963 5496 2965 5516
rect 2969 5496 2971 5516
rect 2983 5496 2985 5516
rect 2989 5496 2991 5516
rect 3029 5476 3031 5516
rect 3035 5488 3037 5516
rect 3049 5488 3051 5516
rect 3035 5476 3051 5488
rect 3055 5476 3057 5516
rect 3069 5476 3071 5516
rect 3075 5476 3077 5516
rect 3151 5476 3153 5516
rect 3157 5476 3163 5516
rect 3167 5476 3169 5516
rect 3209 5476 3211 5516
rect 3215 5488 3217 5516
rect 3229 5488 3231 5516
rect 3215 5476 3231 5488
rect 3235 5476 3237 5516
rect 3249 5476 3251 5516
rect 3255 5476 3257 5516
rect 3333 5476 3335 5516
rect 3339 5476 3341 5516
rect 3353 5476 3355 5516
rect 3359 5476 3365 5516
rect 3369 5476 3371 5516
rect 3409 5496 3411 5516
rect 3415 5496 3417 5516
rect 3429 5496 3431 5516
rect 3435 5496 3437 5516
rect 3489 5496 3491 5516
rect 3495 5496 3497 5516
rect 3509 5496 3511 5516
rect 3515 5496 3517 5516
rect 3529 5496 3531 5516
rect 3519 5476 3531 5496
rect 3535 5476 3537 5516
rect 3589 5476 3591 5516
rect 3595 5488 3597 5516
rect 3609 5488 3611 5516
rect 3595 5476 3611 5488
rect 3615 5476 3617 5516
rect 3629 5476 3631 5516
rect 3635 5476 3637 5516
rect 3703 5496 3705 5516
rect 3709 5496 3711 5516
rect 3723 5496 3725 5516
rect 3729 5496 3731 5516
rect 3769 5476 3771 5516
rect 3775 5486 3777 5516
rect 3789 5486 3791 5516
rect 3775 5476 3791 5486
rect 3795 5476 3797 5516
rect 3809 5476 3811 5516
rect 3815 5504 3831 5516
rect 3815 5476 3817 5504
rect 3829 5476 3831 5504
rect 3835 5476 3837 5516
rect 3903 5496 3905 5516
rect 3909 5496 3911 5516
rect 3923 5496 3925 5516
rect 3929 5496 3931 5516
rect 3969 5476 3971 5516
rect 3975 5488 3977 5516
rect 3989 5488 3991 5516
rect 3975 5476 3991 5488
rect 3995 5476 3997 5516
rect 4009 5476 4011 5516
rect 4015 5476 4017 5516
rect 4106 5458 4108 5516
rect 4094 5456 4108 5458
rect 4112 5456 4116 5516
rect 4120 5456 4124 5516
rect 4128 5456 4130 5516
rect 4191 5476 4193 5516
rect 4197 5476 4203 5516
rect 4207 5476 4209 5516
rect 4249 5496 4251 5516
rect 4255 5496 4257 5516
rect 4323 5476 4325 5516
rect 4329 5476 4331 5516
rect 4343 5476 4345 5516
rect 4349 5488 4351 5516
rect 4363 5488 4365 5516
rect 4349 5476 4365 5488
rect 4369 5476 4371 5516
rect 4431 5476 4433 5516
rect 4437 5476 4443 5516
rect 4447 5476 4449 5516
rect 4491 5476 4493 5516
rect 4497 5476 4503 5516
rect 4507 5476 4509 5516
rect 4583 5476 4585 5516
rect 4589 5476 4591 5516
rect 4603 5476 4605 5516
rect 4609 5488 4611 5516
rect 4623 5488 4625 5516
rect 4609 5476 4625 5488
rect 4629 5476 4631 5516
rect 4683 5476 4685 5516
rect 4689 5476 4691 5516
rect 4703 5476 4705 5516
rect 4709 5488 4711 5516
rect 4723 5488 4725 5516
rect 4709 5476 4725 5488
rect 4729 5476 4731 5516
rect 4793 5476 4795 5516
rect 4799 5476 4801 5516
rect 4813 5476 4815 5516
rect 4819 5476 4825 5516
rect 4829 5476 4831 5516
rect 4883 5476 4885 5516
rect 4889 5476 4891 5516
rect 4903 5476 4905 5516
rect 4909 5488 4911 5516
rect 4923 5488 4925 5516
rect 4909 5476 4925 5488
rect 4929 5476 4931 5516
rect 4991 5476 4993 5516
rect 4997 5476 5003 5516
rect 5007 5476 5009 5516
rect 5073 5476 5075 5516
rect 5079 5476 5081 5516
rect 5093 5476 5095 5516
rect 5099 5476 5105 5516
rect 5109 5476 5111 5516
rect 5151 5476 5153 5516
rect 5157 5476 5163 5516
rect 5167 5476 5169 5516
rect 5229 5476 5231 5516
rect 5235 5488 5237 5516
rect 5249 5488 5251 5516
rect 5235 5476 5251 5488
rect 5255 5476 5257 5516
rect 5269 5476 5271 5516
rect 5275 5476 5277 5516
rect 5353 5476 5355 5516
rect 5359 5476 5361 5516
rect 5373 5476 5375 5516
rect 5379 5476 5385 5516
rect 5389 5476 5391 5516
rect 5429 5476 5431 5516
rect 5435 5488 5437 5516
rect 5449 5488 5451 5516
rect 5435 5476 5451 5488
rect 5455 5476 5457 5516
rect 5469 5476 5471 5516
rect 5475 5476 5477 5516
rect 5531 5476 5533 5516
rect 5537 5476 5543 5516
rect 5547 5476 5549 5516
rect 5610 5456 5612 5516
rect 5616 5456 5620 5516
rect 5624 5456 5628 5516
rect 5632 5458 5634 5516
rect 5733 5476 5735 5516
rect 5739 5476 5741 5516
rect 5753 5476 5755 5516
rect 5759 5476 5765 5516
rect 5769 5476 5771 5516
rect 5844 5476 5846 5516
rect 5850 5476 5854 5516
rect 5858 5476 5860 5516
rect 5872 5476 5874 5516
rect 5878 5476 5882 5516
rect 5886 5476 5888 5516
rect 5931 5476 5933 5516
rect 5937 5476 5943 5516
rect 5947 5476 5949 5516
rect 5632 5456 5646 5458
rect 6010 5456 6012 5516
rect 6016 5456 6020 5516
rect 6024 5456 6028 5516
rect 6032 5458 6034 5516
rect 6112 5476 6114 5516
rect 6118 5476 6122 5516
rect 6126 5476 6128 5516
rect 6140 5496 6144 5516
rect 6148 5496 6150 5516
rect 6032 5456 6046 5458
rect 6223 5476 6225 5516
rect 6229 5476 6231 5516
rect 6243 5476 6245 5516
rect 6249 5488 6251 5516
rect 6263 5488 6265 5516
rect 6249 5476 6265 5488
rect 6269 5476 6271 5516
rect 6309 5476 6311 5516
rect 6315 5488 6317 5516
rect 6329 5488 6331 5516
rect 6315 5476 6331 5488
rect 6335 5476 6337 5516
rect 6349 5476 6351 5516
rect 6355 5476 6357 5516
rect 6423 5476 6425 5516
rect 6429 5476 6431 5516
rect 6443 5476 6445 5516
rect 6449 5488 6451 5516
rect 6463 5488 6465 5516
rect 6449 5476 6465 5488
rect 6469 5476 6471 5516
rect 6546 5458 6548 5516
rect 6534 5456 6548 5458
rect 6552 5456 6556 5516
rect 6560 5456 6564 5516
rect 6568 5456 6570 5516
rect 6630 5496 6632 5516
rect 6636 5496 6640 5516
rect 6652 5476 6654 5516
rect 6658 5476 6662 5516
rect 6666 5476 6668 5516
rect 41 5064 43 5104
rect 47 5064 49 5104
rect 61 5064 65 5084
rect 69 5064 71 5084
rect 109 5064 111 5104
rect 115 5084 128 5104
rect 291 5084 301 5104
rect 115 5064 119 5084
rect 131 5064 133 5084
rect 137 5064 143 5084
rect 147 5064 149 5084
rect 161 5064 163 5084
rect 167 5064 171 5084
rect 175 5064 177 5084
rect 215 5064 217 5084
rect 221 5064 225 5084
rect 237 5064 239 5084
rect 243 5064 249 5084
rect 253 5064 255 5084
rect 267 5064 271 5084
rect 275 5064 281 5084
rect 285 5064 287 5084
rect 299 5064 301 5084
rect 305 5064 307 5104
rect 351 5064 353 5104
rect 357 5064 363 5104
rect 367 5064 369 5104
rect 450 5064 452 5084
rect 456 5064 460 5084
rect 472 5064 474 5104
rect 478 5064 482 5104
rect 486 5064 488 5104
rect 551 5064 553 5104
rect 557 5064 563 5104
rect 567 5064 569 5104
rect 613 5064 615 5104
rect 619 5084 629 5104
rect 792 5084 805 5104
rect 619 5064 621 5084
rect 633 5064 635 5084
rect 639 5064 645 5084
rect 649 5064 653 5084
rect 665 5064 667 5084
rect 671 5064 677 5084
rect 681 5064 683 5084
rect 695 5064 699 5084
rect 703 5064 705 5084
rect 743 5064 745 5084
rect 749 5064 753 5084
rect 757 5064 759 5084
rect 771 5064 773 5084
rect 777 5064 783 5084
rect 787 5064 789 5084
rect 801 5064 805 5084
rect 809 5064 811 5104
rect 851 5064 853 5104
rect 857 5064 863 5104
rect 867 5064 869 5104
rect 943 5064 945 5104
rect 949 5064 951 5104
rect 963 5064 965 5104
rect 969 5092 985 5104
rect 969 5064 971 5092
rect 983 5064 985 5092
rect 989 5064 991 5104
rect 1043 5064 1045 5104
rect 1049 5064 1051 5104
rect 1063 5064 1065 5104
rect 1069 5092 1085 5104
rect 1069 5064 1071 5092
rect 1083 5064 1085 5092
rect 1089 5064 1091 5104
rect 1153 5064 1155 5104
rect 1159 5064 1161 5104
rect 1173 5064 1175 5104
rect 1179 5064 1185 5104
rect 1189 5064 1191 5104
rect 1229 5064 1231 5104
rect 1235 5084 1248 5104
rect 1411 5084 1421 5104
rect 1235 5064 1239 5084
rect 1251 5064 1253 5084
rect 1257 5064 1263 5084
rect 1267 5064 1269 5084
rect 1281 5064 1283 5084
rect 1287 5064 1291 5084
rect 1295 5064 1297 5084
rect 1335 5064 1337 5084
rect 1341 5064 1345 5084
rect 1357 5064 1359 5084
rect 1363 5064 1369 5084
rect 1373 5064 1375 5084
rect 1387 5064 1391 5084
rect 1395 5064 1401 5084
rect 1405 5064 1407 5084
rect 1419 5064 1421 5084
rect 1425 5064 1427 5104
rect 1491 5064 1493 5104
rect 1497 5064 1503 5104
rect 1507 5064 1509 5104
rect 1551 5064 1553 5104
rect 1557 5064 1563 5104
rect 1567 5064 1569 5104
rect 1629 5064 1631 5104
rect 1635 5084 1648 5104
rect 1811 5084 1821 5104
rect 1635 5064 1639 5084
rect 1651 5064 1653 5084
rect 1657 5064 1663 5084
rect 1667 5064 1669 5084
rect 1681 5064 1683 5084
rect 1687 5064 1691 5084
rect 1695 5064 1697 5084
rect 1735 5064 1737 5084
rect 1741 5064 1745 5084
rect 1757 5064 1759 5084
rect 1763 5064 1769 5084
rect 1773 5064 1775 5084
rect 1787 5064 1791 5084
rect 1795 5064 1801 5084
rect 1805 5064 1807 5084
rect 1819 5064 1821 5084
rect 1825 5064 1827 5104
rect 1904 5064 1906 5104
rect 1910 5064 1914 5104
rect 1918 5064 1920 5104
rect 1932 5064 1934 5104
rect 1938 5064 1942 5104
rect 1946 5064 1948 5104
rect 1989 5064 1991 5084
rect 1995 5064 1997 5084
rect 2073 5064 2075 5104
rect 2079 5064 2081 5104
rect 2093 5064 2095 5104
rect 2099 5064 2105 5104
rect 2109 5064 2111 5104
rect 2151 5064 2153 5104
rect 2157 5064 2163 5104
rect 2167 5064 2169 5104
rect 2243 5064 2245 5104
rect 2249 5084 2261 5104
rect 2434 5122 2448 5124
rect 2249 5064 2251 5084
rect 2263 5064 2265 5084
rect 2269 5064 2271 5084
rect 2283 5064 2285 5084
rect 2289 5064 2291 5084
rect 2351 5064 2353 5104
rect 2357 5064 2363 5104
rect 2367 5064 2369 5104
rect 2446 5064 2448 5122
rect 2452 5064 2456 5124
rect 2460 5064 2464 5124
rect 2468 5064 2470 5124
rect 2523 5064 2525 5084
rect 2529 5064 2531 5084
rect 2543 5064 2545 5084
rect 2549 5064 2551 5084
rect 2589 5064 2591 5084
rect 2595 5064 2597 5084
rect 2673 5064 2675 5104
rect 2679 5064 2681 5104
rect 2693 5064 2695 5104
rect 2699 5064 2705 5104
rect 2709 5064 2711 5104
rect 2749 5064 2751 5084
rect 2755 5064 2757 5084
rect 2769 5064 2771 5084
rect 2775 5064 2777 5084
rect 2851 5064 2853 5104
rect 2857 5064 2863 5104
rect 2867 5064 2869 5104
rect 2931 5064 2933 5104
rect 2937 5064 2943 5104
rect 2947 5064 2949 5104
rect 3294 5122 3308 5124
rect 3019 5084 3031 5104
rect 2989 5064 2991 5084
rect 2995 5064 2997 5084
rect 3009 5064 3011 5084
rect 3015 5064 3017 5084
rect 3029 5064 3031 5084
rect 3035 5064 3037 5104
rect 3113 5064 3115 5104
rect 3119 5064 3121 5104
rect 3133 5064 3135 5104
rect 3139 5064 3145 5104
rect 3149 5064 3151 5104
rect 3191 5064 3193 5104
rect 3197 5064 3203 5104
rect 3207 5064 3209 5104
rect 3306 5064 3308 5122
rect 3312 5064 3316 5124
rect 3320 5064 3324 5124
rect 3328 5064 3330 5124
rect 3383 5064 3385 5084
rect 3389 5064 3391 5084
rect 3450 5064 3452 5084
rect 3456 5064 3460 5084
rect 3472 5064 3474 5104
rect 3478 5064 3482 5104
rect 3486 5064 3488 5104
rect 3543 5064 3545 5084
rect 3549 5064 3551 5084
rect 3563 5064 3565 5084
rect 3569 5064 3571 5084
rect 3609 5064 3611 5104
rect 3615 5092 3631 5104
rect 3615 5064 3617 5092
rect 3629 5064 3631 5092
rect 3635 5064 3637 5104
rect 3649 5064 3651 5104
rect 3655 5064 3657 5104
rect 3723 5064 3725 5104
rect 3729 5064 3731 5104
rect 3743 5064 3745 5104
rect 3749 5092 3765 5104
rect 3749 5064 3751 5092
rect 3763 5064 3765 5092
rect 3769 5064 3771 5104
rect 3809 5064 3811 5084
rect 3815 5064 3817 5084
rect 3829 5064 3831 5084
rect 3835 5064 3837 5084
rect 3891 5064 3893 5104
rect 3897 5064 3903 5104
rect 3907 5064 3909 5104
rect 3991 5064 3993 5104
rect 3997 5064 4003 5104
rect 4007 5064 4009 5104
rect 4049 5064 4051 5104
rect 4055 5092 4071 5104
rect 4055 5064 4057 5092
rect 4069 5064 4071 5092
rect 4075 5064 4077 5104
rect 4089 5064 4091 5104
rect 4095 5064 4097 5104
rect 4171 5064 4173 5104
rect 4177 5064 4183 5104
rect 4187 5064 4189 5104
rect 4253 5064 4255 5104
rect 4259 5064 4261 5104
rect 4273 5064 4275 5104
rect 4279 5064 4285 5104
rect 4289 5064 4291 5104
rect 4351 5064 4353 5104
rect 4357 5064 4363 5104
rect 4367 5064 4369 5104
rect 4423 5064 4425 5104
rect 4429 5064 4431 5104
rect 4443 5064 4445 5104
rect 4449 5092 4465 5104
rect 4449 5064 4451 5092
rect 4463 5064 4465 5092
rect 4469 5064 4471 5104
rect 4523 5064 4525 5104
rect 4529 5064 4531 5104
rect 4543 5064 4545 5104
rect 4549 5092 4565 5104
rect 4549 5064 4551 5092
rect 4563 5064 4565 5092
rect 4569 5064 4571 5104
rect 4611 5064 4613 5104
rect 4617 5064 4623 5104
rect 4627 5064 4629 5104
rect 4691 5064 4693 5104
rect 4697 5064 4703 5104
rect 4707 5064 4709 5104
rect 4854 5122 4868 5124
rect 4769 5064 4771 5084
rect 4775 5064 4777 5084
rect 4866 5064 4868 5122
rect 4872 5064 4876 5124
rect 4880 5064 4884 5124
rect 4888 5064 4890 5124
rect 4929 5064 4931 5104
rect 4935 5092 4951 5104
rect 4935 5064 4937 5092
rect 4949 5064 4951 5092
rect 4955 5064 4957 5104
rect 4969 5064 4971 5104
rect 4975 5064 4977 5104
rect 5029 5064 5031 5104
rect 5035 5064 5037 5104
rect 5091 5064 5093 5104
rect 5097 5064 5103 5104
rect 5107 5064 5109 5104
rect 5169 5064 5171 5104
rect 5175 5064 5177 5104
rect 5189 5064 5191 5104
rect 5195 5064 5197 5104
rect 5251 5064 5253 5104
rect 5257 5064 5263 5104
rect 5267 5064 5269 5104
rect 5329 5064 5331 5104
rect 5335 5092 5351 5104
rect 5335 5064 5337 5092
rect 5349 5064 5351 5092
rect 5355 5064 5357 5104
rect 5369 5064 5371 5104
rect 5375 5064 5377 5104
rect 5430 5064 5432 5124
rect 5436 5064 5440 5124
rect 5444 5064 5448 5124
rect 5452 5122 5466 5124
rect 5452 5064 5454 5122
rect 5530 5064 5532 5124
rect 5536 5064 5540 5124
rect 5544 5064 5548 5124
rect 5552 5122 5566 5124
rect 5552 5064 5554 5122
rect 5629 5064 5631 5084
rect 5635 5064 5637 5084
rect 5690 5064 5692 5124
rect 5696 5064 5700 5124
rect 5704 5064 5708 5124
rect 5712 5122 5726 5124
rect 5712 5064 5714 5122
rect 5789 5064 5791 5104
rect 5795 5092 5811 5104
rect 5795 5064 5797 5092
rect 5809 5064 5811 5092
rect 5815 5064 5817 5104
rect 5829 5064 5831 5104
rect 5835 5064 5837 5104
rect 5911 5064 5913 5104
rect 5917 5064 5923 5104
rect 5927 5064 5929 5104
rect 5970 5064 5972 5124
rect 5976 5064 5980 5124
rect 5984 5064 5988 5124
rect 5992 5122 6006 5124
rect 5992 5064 5994 5122
rect 6071 5064 6073 5104
rect 6077 5064 6083 5104
rect 6087 5064 6089 5104
rect 6170 5064 6172 5084
rect 6176 5064 6180 5084
rect 6192 5064 6194 5104
rect 6198 5064 6202 5104
rect 6206 5064 6208 5104
rect 6334 5122 6348 5124
rect 6263 5064 6265 5084
rect 6269 5064 6271 5084
rect 6346 5064 6348 5122
rect 6352 5064 6356 5124
rect 6360 5064 6364 5124
rect 6368 5064 6370 5124
rect 6434 5122 6448 5124
rect 6446 5064 6448 5122
rect 6452 5064 6456 5124
rect 6460 5064 6464 5124
rect 6468 5064 6470 5124
rect 6594 5122 6608 5124
rect 6509 5064 6511 5084
rect 6515 5064 6517 5084
rect 6606 5064 6608 5122
rect 6612 5064 6616 5124
rect 6620 5064 6624 5124
rect 6628 5064 6630 5124
rect 6671 5064 6673 5104
rect 6677 5064 6683 5104
rect 6687 5064 6689 5104
rect 41 4996 43 5036
rect 47 4996 49 5036
rect 61 5016 65 5036
rect 69 5016 71 5036
rect 121 4996 123 5036
rect 127 4996 129 5036
rect 141 5016 145 5036
rect 149 5016 151 5036
rect 211 4996 213 5036
rect 217 4996 223 5036
rect 227 4996 229 5036
rect 269 4996 271 5036
rect 275 5016 279 5036
rect 291 5016 293 5036
rect 297 5016 303 5036
rect 307 5016 309 5036
rect 321 5016 323 5036
rect 327 5016 331 5036
rect 335 5016 337 5036
rect 375 5016 377 5036
rect 381 5016 385 5036
rect 397 5016 399 5036
rect 403 5016 409 5036
rect 413 5016 415 5036
rect 427 5016 431 5036
rect 435 5016 441 5036
rect 445 5016 447 5036
rect 459 5016 461 5036
rect 275 4996 288 5016
rect 451 4996 461 5016
rect 465 4996 467 5036
rect 530 5016 532 5036
rect 536 5016 540 5036
rect 552 4996 554 5036
rect 558 4996 562 5036
rect 566 4996 568 5036
rect 631 4996 633 5036
rect 637 4996 643 5036
rect 647 4996 649 5036
rect 691 4996 693 5036
rect 697 4996 703 5036
rect 707 4996 709 5036
rect 791 4996 793 5036
rect 797 4996 803 5036
rect 807 4996 809 5036
rect 849 4996 851 5036
rect 855 5016 859 5036
rect 871 5016 873 5036
rect 877 5016 883 5036
rect 887 5016 889 5036
rect 901 5016 903 5036
rect 907 5016 911 5036
rect 915 5016 917 5036
rect 955 5016 957 5036
rect 961 5016 965 5036
rect 977 5016 979 5036
rect 983 5016 989 5036
rect 993 5016 995 5036
rect 1007 5016 1011 5036
rect 1015 5016 1021 5036
rect 1025 5016 1027 5036
rect 1039 5016 1041 5036
rect 855 4996 868 5016
rect 1031 4996 1041 5016
rect 1045 4996 1047 5036
rect 1101 4996 1103 5036
rect 1107 4996 1109 5036
rect 1121 5016 1125 5036
rect 1129 5016 1131 5036
rect 1190 5016 1192 5036
rect 1196 5016 1200 5036
rect 1212 4996 1214 5036
rect 1218 4996 1222 5036
rect 1226 4996 1228 5036
rect 1291 4996 1293 5036
rect 1297 4996 1303 5036
rect 1307 4996 1309 5036
rect 1361 4996 1363 5036
rect 1367 4996 1369 5036
rect 1381 5016 1385 5036
rect 1389 5016 1391 5036
rect 1431 4996 1433 5036
rect 1437 4996 1443 5036
rect 1447 4996 1449 5036
rect 1531 4996 1533 5036
rect 1537 4996 1543 5036
rect 1547 4996 1549 5036
rect 1603 4996 1605 5036
rect 1609 4996 1611 5036
rect 1623 4996 1625 5036
rect 1629 5008 1631 5036
rect 1643 5008 1645 5036
rect 1629 4996 1645 5008
rect 1649 4996 1651 5036
rect 1711 4996 1713 5036
rect 1717 4996 1723 5036
rect 1727 4996 1729 5036
rect 1783 4996 1785 5036
rect 1789 4996 1791 5036
rect 1803 4996 1805 5036
rect 1809 5008 1811 5036
rect 1823 5008 1825 5036
rect 1809 4996 1825 5008
rect 1829 4996 1831 5036
rect 1871 4996 1873 5036
rect 1877 4996 1883 5036
rect 1887 4996 1889 5036
rect 1963 4996 1965 5036
rect 1969 4996 1971 5036
rect 1983 4996 1985 5036
rect 1989 5008 1991 5036
rect 2003 5008 2005 5036
rect 1989 4996 2005 5008
rect 2009 4996 2011 5036
rect 2063 4996 2065 5036
rect 2069 4996 2071 5036
rect 2083 4996 2085 5036
rect 2089 5008 2091 5036
rect 2103 5008 2105 5036
rect 2089 4996 2105 5008
rect 2109 4996 2111 5036
rect 2173 4996 2175 5036
rect 2179 4996 2181 5036
rect 2193 4996 2195 5036
rect 2199 4996 2205 5036
rect 2209 4996 2211 5036
rect 2249 5016 2251 5036
rect 2255 5016 2257 5036
rect 2323 5016 2325 5036
rect 2329 5016 2331 5036
rect 2343 5016 2345 5036
rect 2349 5016 2351 5036
rect 2403 4996 2405 5036
rect 2409 5016 2411 5036
rect 2423 5016 2425 5036
rect 2429 5016 2431 5036
rect 2443 5016 2445 5036
rect 2449 5016 2451 5036
rect 2409 4996 2421 5016
rect 2511 4996 2513 5036
rect 2517 4996 2523 5036
rect 2527 4996 2529 5036
rect 2583 4996 2585 5036
rect 2589 4996 2591 5036
rect 2603 4996 2605 5036
rect 2609 5008 2611 5036
rect 2623 5008 2625 5036
rect 2609 4996 2625 5008
rect 2629 4996 2631 5036
rect 2683 4996 2685 5036
rect 2689 4996 2691 5036
rect 2703 4996 2705 5036
rect 2709 5008 2711 5036
rect 2723 5008 2725 5036
rect 2709 4996 2725 5008
rect 2729 4996 2731 5036
rect 2783 5016 2785 5036
rect 2789 5016 2791 5036
rect 2829 4996 2831 5036
rect 2835 5008 2837 5036
rect 2849 5008 2851 5036
rect 2835 4996 2851 5008
rect 2855 4996 2857 5036
rect 2869 4996 2871 5036
rect 2875 4996 2877 5036
rect 2943 4996 2945 5036
rect 2949 4996 2951 5036
rect 2963 4996 2965 5036
rect 2969 5008 2971 5036
rect 2983 5008 2985 5036
rect 2969 4996 2985 5008
rect 2989 4996 2991 5036
rect 3043 4996 3045 5036
rect 3049 4996 3051 5036
rect 3063 4996 3065 5036
rect 3069 5008 3071 5036
rect 3083 5008 3085 5036
rect 3069 4996 3085 5008
rect 3089 4996 3091 5036
rect 3143 5016 3145 5036
rect 3149 5016 3151 5036
rect 3163 5016 3165 5036
rect 3169 5016 3171 5036
rect 3223 4996 3225 5036
rect 3229 4996 3231 5036
rect 3291 4996 3293 5036
rect 3297 4996 3303 5036
rect 3307 4996 3309 5036
rect 3363 4996 3365 5036
rect 3369 4996 3371 5036
rect 3383 4996 3385 5036
rect 3389 5008 3391 5036
rect 3403 5008 3405 5036
rect 3389 4996 3405 5008
rect 3409 4996 3411 5036
rect 3453 4996 3455 5036
rect 3459 5016 3461 5036
rect 3473 5016 3475 5036
rect 3479 5016 3485 5036
rect 3489 5016 3493 5036
rect 3505 5016 3507 5036
rect 3511 5016 3517 5036
rect 3521 5016 3523 5036
rect 3535 5016 3539 5036
rect 3543 5016 3545 5036
rect 3583 5016 3585 5036
rect 3589 5016 3593 5036
rect 3597 5016 3599 5036
rect 3611 5016 3613 5036
rect 3617 5016 3623 5036
rect 3627 5016 3629 5036
rect 3641 5016 3645 5036
rect 3459 4996 3469 5016
rect 3632 4996 3645 5016
rect 3649 4996 3651 5036
rect 3689 4996 3691 5036
rect 3695 5008 3697 5036
rect 3709 5008 3711 5036
rect 3695 4996 3711 5008
rect 3715 4996 3717 5036
rect 3729 4996 3731 5036
rect 3735 4996 3737 5036
rect 3810 5016 3812 5036
rect 3816 5016 3820 5036
rect 3832 4996 3834 5036
rect 3838 4996 3842 5036
rect 3846 4996 3848 5036
rect 3926 4978 3928 5036
rect 3914 4976 3928 4978
rect 3932 4976 3936 5036
rect 3940 4976 3944 5036
rect 3948 4976 3950 5036
rect 4010 5016 4012 5036
rect 4016 5016 4020 5036
rect 4032 4996 4034 5036
rect 4038 4996 4042 5036
rect 4046 4996 4048 5036
rect 4103 4996 4105 5036
rect 4109 4996 4111 5036
rect 4173 4996 4175 5036
rect 4179 4996 4181 5036
rect 4193 4996 4195 5036
rect 4199 4996 4205 5036
rect 4209 4996 4211 5036
rect 4271 4996 4273 5036
rect 4277 4996 4283 5036
rect 4287 4996 4289 5036
rect 4329 4996 4331 5036
rect 4335 4996 4341 5036
rect 4345 4996 4347 5036
rect 4359 4996 4361 5036
rect 4365 4996 4367 5036
rect 4443 4996 4445 5036
rect 4449 4996 4451 5036
rect 4463 4996 4465 5036
rect 4469 5008 4471 5036
rect 4483 5008 4485 5036
rect 4469 4996 4485 5008
rect 4489 4996 4491 5036
rect 4530 4976 4532 5036
rect 4536 4976 4540 5036
rect 4544 4976 4548 5036
rect 4552 4978 4554 5036
rect 4629 4996 4631 5036
rect 4635 5008 4637 5036
rect 4649 5008 4651 5036
rect 4635 4996 4651 5008
rect 4655 4996 4657 5036
rect 4669 4996 4671 5036
rect 4675 4996 4677 5036
rect 4751 4996 4753 5036
rect 4757 4996 4763 5036
rect 4767 4996 4769 5036
rect 4833 4996 4835 5036
rect 4839 4996 4841 5036
rect 4853 4996 4855 5036
rect 4859 4996 4865 5036
rect 4869 4996 4871 5036
rect 4931 4996 4933 5036
rect 4937 4996 4943 5036
rect 4947 4996 4949 5036
rect 4991 4996 4993 5036
rect 4997 4996 5003 5036
rect 5007 4996 5009 5036
rect 5069 4996 5071 5036
rect 5075 4996 5081 5036
rect 5085 4996 5087 5036
rect 5099 4996 5101 5036
rect 5105 4996 5107 5036
rect 5191 4996 5193 5036
rect 5197 4996 5203 5036
rect 5207 4996 5209 5036
rect 5273 4996 5275 5036
rect 5279 4996 5281 5036
rect 5293 4996 5295 5036
rect 5299 4996 5305 5036
rect 5309 4996 5311 5036
rect 5349 4996 5351 5036
rect 5355 4996 5361 5036
rect 5365 4996 5367 5036
rect 5379 4996 5381 5036
rect 5385 4996 5387 5036
rect 5484 4996 5486 5036
rect 5490 4996 5494 5036
rect 5498 4996 5500 5036
rect 5512 4996 5514 5036
rect 5518 4996 5522 5036
rect 5526 4996 5528 5036
rect 5591 4996 5593 5036
rect 5597 4996 5603 5036
rect 5607 4996 5609 5036
rect 4552 4976 4566 4978
rect 5650 4976 5652 5036
rect 5656 4976 5660 5036
rect 5664 4976 5668 5036
rect 5672 4978 5674 5036
rect 5770 5016 5772 5036
rect 5776 5016 5780 5036
rect 5672 4976 5686 4978
rect 5792 4996 5794 5036
rect 5798 4996 5802 5036
rect 5806 4996 5808 5036
rect 5886 4978 5888 5036
rect 5874 4976 5888 4978
rect 5892 4976 5896 5036
rect 5900 4976 5904 5036
rect 5908 4976 5910 5036
rect 5971 4996 5973 5036
rect 5977 4996 5983 5036
rect 5987 4996 5989 5036
rect 6032 4996 6034 5036
rect 6038 4996 6042 5036
rect 6046 4996 6048 5036
rect 6060 4996 6062 5036
rect 6066 4996 6070 5036
rect 6074 4996 6076 5036
rect 6186 4978 6188 5036
rect 6174 4976 6188 4978
rect 6192 4976 6196 5036
rect 6200 4976 6204 5036
rect 6208 4976 6210 5036
rect 6249 4996 6251 5036
rect 6255 5008 6257 5036
rect 6269 5008 6271 5036
rect 6255 4996 6271 5008
rect 6275 4996 6277 5036
rect 6289 4996 6291 5036
rect 6295 4996 6297 5036
rect 6386 4978 6388 5036
rect 6374 4976 6388 4978
rect 6392 4976 6396 5036
rect 6400 4976 6404 5036
rect 6408 4976 6410 5036
rect 6486 4978 6488 5036
rect 6474 4976 6488 4978
rect 6492 4976 6496 5036
rect 6500 4976 6504 5036
rect 6508 4976 6510 5036
rect 6551 4996 6553 5036
rect 6557 4996 6563 5036
rect 6567 4996 6569 5036
rect 6643 5016 6645 5036
rect 6649 5016 6651 5036
rect 29 4584 31 4624
rect 35 4584 37 4624
rect 49 4584 51 4624
rect 55 4584 57 4624
rect 69 4584 71 4624
rect 75 4584 77 4624
rect 89 4584 91 4624
rect 95 4584 97 4624
rect 109 4584 111 4624
rect 115 4584 117 4624
rect 129 4584 131 4624
rect 135 4584 137 4624
rect 149 4584 151 4624
rect 155 4584 157 4624
rect 169 4584 171 4624
rect 175 4584 177 4624
rect 243 4584 245 4604
rect 249 4584 251 4604
rect 263 4584 265 4604
rect 269 4584 271 4604
rect 323 4584 325 4604
rect 329 4584 331 4604
rect 390 4584 392 4604
rect 396 4584 400 4604
rect 412 4584 414 4624
rect 418 4584 422 4624
rect 426 4584 428 4624
rect 483 4584 485 4604
rect 489 4584 491 4604
rect 543 4584 545 4604
rect 549 4584 551 4604
rect 563 4584 565 4604
rect 569 4584 571 4604
rect 633 4584 635 4624
rect 639 4584 641 4624
rect 653 4584 655 4624
rect 659 4584 665 4624
rect 669 4584 671 4624
rect 709 4584 711 4604
rect 715 4584 717 4604
rect 729 4584 731 4604
rect 735 4584 737 4604
rect 801 4584 803 4624
rect 807 4584 809 4624
rect 821 4584 825 4604
rect 829 4584 831 4604
rect 891 4584 893 4624
rect 897 4584 903 4624
rect 907 4584 909 4624
rect 949 4584 951 4624
rect 955 4604 968 4624
rect 1131 4604 1141 4624
rect 955 4584 959 4604
rect 971 4584 973 4604
rect 977 4584 983 4604
rect 987 4584 989 4604
rect 1001 4584 1003 4604
rect 1007 4584 1011 4604
rect 1015 4584 1017 4604
rect 1055 4584 1057 4604
rect 1061 4584 1065 4604
rect 1077 4584 1079 4604
rect 1083 4584 1089 4604
rect 1093 4584 1095 4604
rect 1107 4584 1111 4604
rect 1115 4584 1121 4604
rect 1125 4584 1127 4604
rect 1139 4584 1141 4604
rect 1145 4584 1147 4624
rect 1203 4584 1205 4624
rect 1209 4584 1211 4624
rect 1223 4584 1225 4624
rect 1229 4612 1245 4624
rect 1229 4584 1231 4612
rect 1243 4584 1245 4612
rect 1249 4584 1251 4624
rect 1311 4584 1313 4624
rect 1317 4584 1323 4624
rect 1327 4584 1329 4624
rect 1371 4584 1373 4624
rect 1377 4584 1383 4624
rect 1387 4584 1389 4624
rect 1463 4584 1465 4624
rect 1469 4584 1471 4624
rect 1483 4584 1485 4624
rect 1489 4612 1505 4624
rect 1489 4584 1491 4612
rect 1503 4584 1505 4612
rect 1509 4584 1511 4624
rect 1549 4584 1551 4604
rect 1555 4584 1557 4604
rect 1569 4584 1571 4604
rect 1575 4584 1577 4604
rect 1629 4584 1631 4604
rect 1635 4584 1637 4604
rect 1649 4584 1651 4604
rect 1655 4584 1657 4604
rect 1709 4584 1711 4604
rect 1715 4584 1717 4604
rect 1769 4584 1771 4604
rect 1775 4584 1777 4604
rect 1789 4584 1791 4604
rect 1795 4584 1797 4604
rect 1849 4584 1851 4624
rect 1855 4612 1871 4624
rect 1855 4584 1857 4612
rect 1869 4584 1871 4612
rect 1875 4584 1877 4624
rect 1889 4584 1891 4624
rect 1895 4584 1897 4624
rect 1949 4584 1951 4624
rect 1955 4604 1968 4624
rect 2131 4604 2141 4624
rect 1955 4584 1959 4604
rect 1971 4584 1973 4604
rect 1977 4584 1983 4604
rect 1987 4584 1989 4604
rect 2001 4584 2003 4604
rect 2007 4584 2011 4604
rect 2015 4584 2017 4604
rect 2055 4584 2057 4604
rect 2061 4584 2065 4604
rect 2077 4584 2079 4604
rect 2083 4584 2089 4604
rect 2093 4584 2095 4604
rect 2107 4584 2111 4604
rect 2115 4584 2121 4604
rect 2125 4584 2127 4604
rect 2139 4584 2141 4604
rect 2145 4584 2147 4624
rect 2211 4584 2213 4624
rect 2217 4584 2223 4624
rect 2227 4584 2229 4624
rect 2283 4584 2285 4624
rect 2289 4604 2301 4624
rect 2289 4584 2291 4604
rect 2303 4584 2305 4604
rect 2309 4584 2311 4604
rect 2323 4584 2325 4604
rect 2329 4584 2331 4604
rect 2371 4584 2373 4624
rect 2377 4584 2383 4624
rect 2387 4584 2389 4624
rect 2449 4584 2451 4604
rect 2455 4584 2457 4604
rect 2469 4584 2471 4604
rect 2475 4584 2477 4604
rect 2532 4584 2534 4624
rect 2538 4584 2542 4624
rect 2546 4584 2548 4624
rect 2560 4584 2564 4604
rect 2568 4584 2570 4604
rect 2643 4584 2645 4604
rect 2649 4584 2651 4604
rect 2689 4584 2691 4624
rect 2695 4604 2708 4624
rect 2871 4604 2881 4624
rect 2695 4584 2699 4604
rect 2711 4584 2713 4604
rect 2717 4584 2723 4604
rect 2727 4584 2729 4604
rect 2741 4584 2743 4604
rect 2747 4584 2751 4604
rect 2755 4584 2757 4604
rect 2795 4584 2797 4604
rect 2801 4584 2805 4604
rect 2817 4584 2819 4604
rect 2823 4584 2829 4604
rect 2833 4584 2835 4604
rect 2847 4584 2851 4604
rect 2855 4584 2861 4604
rect 2865 4584 2867 4604
rect 2879 4584 2881 4604
rect 2885 4584 2887 4624
rect 2929 4584 2931 4624
rect 2935 4612 2951 4624
rect 2935 4584 2937 4612
rect 2949 4584 2951 4612
rect 2955 4584 2957 4624
rect 2969 4584 2971 4624
rect 2975 4584 2977 4624
rect 3029 4584 3031 4624
rect 3035 4604 3048 4624
rect 3211 4604 3221 4624
rect 3035 4584 3039 4604
rect 3051 4584 3053 4604
rect 3057 4584 3063 4604
rect 3067 4584 3069 4604
rect 3081 4584 3083 4604
rect 3087 4584 3091 4604
rect 3095 4584 3097 4604
rect 3135 4584 3137 4604
rect 3141 4584 3145 4604
rect 3157 4584 3159 4604
rect 3163 4584 3169 4604
rect 3173 4584 3175 4604
rect 3187 4584 3191 4604
rect 3195 4584 3201 4604
rect 3205 4584 3207 4604
rect 3219 4584 3221 4604
rect 3225 4584 3227 4624
rect 3269 4584 3271 4624
rect 3275 4604 3288 4624
rect 3451 4604 3461 4624
rect 3275 4584 3279 4604
rect 3291 4584 3293 4604
rect 3297 4584 3303 4604
rect 3307 4584 3309 4604
rect 3321 4584 3323 4604
rect 3327 4584 3331 4604
rect 3335 4584 3337 4604
rect 3375 4584 3377 4604
rect 3381 4584 3385 4604
rect 3397 4584 3399 4604
rect 3403 4584 3409 4604
rect 3413 4584 3415 4604
rect 3427 4584 3431 4604
rect 3435 4584 3441 4604
rect 3445 4584 3447 4604
rect 3459 4584 3461 4604
rect 3465 4584 3467 4624
rect 3523 4584 3525 4624
rect 3529 4584 3531 4624
rect 3543 4584 3545 4624
rect 3549 4612 3565 4624
rect 3549 4584 3551 4612
rect 3563 4584 3565 4612
rect 3569 4584 3571 4624
rect 3623 4584 3625 4624
rect 3629 4584 3631 4624
rect 3691 4584 3693 4624
rect 3697 4584 3703 4624
rect 3707 4584 3709 4624
rect 3763 4584 3765 4624
rect 3769 4584 3771 4624
rect 3783 4584 3785 4624
rect 3789 4612 3805 4624
rect 3789 4584 3791 4612
rect 3803 4584 3805 4612
rect 3809 4584 3811 4624
rect 3853 4584 3855 4624
rect 3859 4604 3869 4624
rect 4032 4604 4045 4624
rect 3859 4584 3861 4604
rect 3873 4584 3875 4604
rect 3879 4584 3885 4604
rect 3889 4584 3893 4604
rect 3905 4584 3907 4604
rect 3911 4584 3917 4604
rect 3921 4584 3923 4604
rect 3935 4584 3939 4604
rect 3943 4584 3945 4604
rect 3983 4584 3985 4604
rect 3989 4584 3993 4604
rect 3997 4584 3999 4604
rect 4011 4584 4013 4604
rect 4017 4584 4023 4604
rect 4027 4584 4029 4604
rect 4041 4584 4045 4604
rect 4049 4584 4051 4624
rect 4103 4584 4105 4624
rect 4109 4584 4111 4624
rect 4171 4584 4173 4624
rect 4177 4584 4183 4624
rect 4187 4584 4189 4624
rect 4229 4584 4231 4624
rect 4235 4604 4248 4624
rect 4494 4642 4508 4644
rect 4411 4604 4421 4624
rect 4235 4584 4239 4604
rect 4251 4584 4253 4604
rect 4257 4584 4263 4604
rect 4267 4584 4269 4604
rect 4281 4584 4283 4604
rect 4287 4584 4291 4604
rect 4295 4584 4297 4604
rect 4335 4584 4337 4604
rect 4341 4584 4345 4604
rect 4357 4584 4359 4604
rect 4363 4584 4369 4604
rect 4373 4584 4375 4604
rect 4387 4584 4391 4604
rect 4395 4584 4401 4604
rect 4405 4584 4407 4604
rect 4419 4584 4421 4604
rect 4425 4584 4427 4624
rect 4506 4584 4508 4642
rect 4512 4584 4516 4644
rect 4520 4584 4524 4644
rect 4528 4584 4530 4644
rect 4569 4584 4571 4604
rect 4575 4584 4577 4604
rect 4629 4584 4631 4624
rect 4635 4584 4637 4624
rect 4703 4584 4705 4604
rect 4709 4584 4711 4604
rect 4749 4584 4751 4624
rect 4755 4612 4771 4624
rect 4755 4584 4757 4612
rect 4769 4584 4771 4612
rect 4775 4584 4777 4624
rect 4789 4584 4791 4624
rect 4795 4584 4797 4624
rect 4849 4584 4851 4604
rect 4855 4584 4857 4604
rect 4869 4584 4871 4604
rect 4875 4584 4877 4604
rect 4931 4584 4933 4624
rect 4937 4584 4943 4624
rect 4947 4584 4949 4624
rect 5011 4584 5013 4624
rect 5017 4584 5023 4624
rect 5027 4584 5029 4624
rect 5111 4584 5113 4624
rect 5117 4584 5123 4624
rect 5127 4584 5129 4624
rect 5169 4584 5171 4624
rect 5175 4612 5191 4624
rect 5175 4584 5177 4612
rect 5189 4584 5191 4612
rect 5195 4584 5197 4624
rect 5209 4584 5211 4624
rect 5215 4584 5217 4624
rect 5283 4584 5285 4624
rect 5289 4596 5291 4624
rect 5303 4596 5305 4624
rect 5289 4584 5305 4596
rect 5309 4584 5311 4624
rect 5323 4584 5325 4624
rect 5329 4614 5345 4624
rect 5329 4584 5331 4614
rect 5343 4584 5345 4614
rect 5349 4584 5351 4624
rect 5391 4584 5393 4624
rect 5397 4584 5403 4624
rect 5407 4584 5409 4624
rect 5491 4584 5493 4624
rect 5497 4584 5503 4624
rect 5507 4584 5509 4624
rect 5550 4584 5552 4644
rect 5556 4584 5560 4644
rect 5564 4584 5568 4644
rect 5572 4642 5586 4644
rect 5572 4584 5574 4642
rect 5671 4584 5673 4624
rect 5677 4584 5683 4624
rect 5687 4584 5689 4624
rect 5730 4584 5732 4644
rect 5736 4584 5740 4644
rect 5744 4584 5748 4644
rect 5752 4642 5766 4644
rect 5752 4584 5754 4642
rect 5843 4584 5845 4604
rect 5849 4584 5851 4604
rect 5890 4584 5892 4644
rect 5896 4584 5900 4644
rect 5904 4584 5908 4644
rect 5912 4642 5926 4644
rect 5912 4584 5914 4642
rect 6013 4584 6015 4624
rect 6019 4584 6021 4624
rect 6033 4584 6035 4624
rect 6039 4584 6045 4624
rect 6049 4584 6051 4624
rect 6089 4584 6091 4624
rect 6095 4612 6111 4624
rect 6095 4584 6097 4612
rect 6109 4584 6111 4612
rect 6115 4584 6117 4624
rect 6129 4584 6131 4624
rect 6135 4584 6137 4624
rect 6211 4584 6213 4624
rect 6217 4584 6223 4624
rect 6227 4584 6229 4624
rect 6272 4584 6274 4624
rect 6278 4584 6282 4624
rect 6286 4584 6288 4624
rect 6300 4584 6304 4604
rect 6308 4584 6310 4604
rect 6370 4584 6372 4644
rect 6376 4584 6380 4644
rect 6384 4584 6388 4644
rect 6392 4642 6406 4644
rect 6392 4584 6394 4642
rect 6594 4642 6608 4644
rect 6493 4584 6495 4624
rect 6499 4584 6501 4624
rect 6513 4584 6515 4624
rect 6519 4584 6525 4624
rect 6529 4584 6531 4624
rect 6606 4584 6608 4642
rect 6612 4584 6616 4644
rect 6620 4584 6624 4644
rect 6628 4584 6630 4644
rect 43 4536 45 4556
rect 49 4536 51 4556
rect 103 4536 105 4556
rect 109 4536 111 4556
rect 123 4536 125 4556
rect 129 4536 131 4556
rect 183 4536 185 4556
rect 189 4536 191 4556
rect 229 4516 231 4556
rect 235 4528 237 4556
rect 249 4528 251 4556
rect 235 4516 251 4528
rect 255 4516 257 4556
rect 269 4516 271 4556
rect 275 4516 277 4556
rect 343 4536 345 4556
rect 349 4536 351 4556
rect 363 4536 365 4556
rect 369 4536 371 4556
rect 409 4516 411 4556
rect 415 4528 417 4556
rect 429 4528 431 4556
rect 415 4516 431 4528
rect 435 4516 437 4556
rect 449 4516 451 4556
rect 455 4516 457 4556
rect 509 4536 511 4556
rect 515 4536 517 4556
rect 529 4536 531 4556
rect 535 4536 537 4556
rect 549 4536 551 4556
rect 539 4516 551 4536
rect 555 4516 557 4556
rect 612 4516 614 4556
rect 618 4516 622 4556
rect 626 4516 628 4556
rect 640 4536 644 4556
rect 648 4536 650 4556
rect 723 4536 725 4556
rect 729 4536 731 4556
rect 769 4536 771 4556
rect 775 4536 777 4556
rect 789 4536 791 4556
rect 795 4536 797 4556
rect 849 4536 851 4556
rect 855 4536 857 4556
rect 909 4536 911 4556
rect 915 4536 917 4556
rect 929 4536 931 4556
rect 935 4536 937 4556
rect 989 4536 991 4556
rect 995 4536 997 4556
rect 1049 4516 1051 4556
rect 1055 4516 1057 4556
rect 1069 4516 1071 4556
rect 1075 4516 1077 4556
rect 1089 4516 1091 4556
rect 1095 4516 1097 4556
rect 1109 4516 1111 4556
rect 1115 4516 1117 4556
rect 1129 4516 1131 4556
rect 1135 4516 1137 4556
rect 1149 4516 1151 4556
rect 1155 4516 1157 4556
rect 1169 4516 1171 4556
rect 1175 4516 1177 4556
rect 1189 4516 1191 4556
rect 1195 4516 1197 4556
rect 1249 4536 1251 4556
rect 1255 4536 1259 4556
rect 1271 4516 1273 4556
rect 1277 4516 1279 4556
rect 1343 4536 1345 4556
rect 1349 4536 1351 4556
rect 1403 4536 1405 4556
rect 1409 4536 1411 4556
rect 1423 4536 1425 4556
rect 1429 4536 1431 4556
rect 1491 4516 1493 4556
rect 1497 4516 1503 4556
rect 1507 4516 1509 4556
rect 1551 4516 1553 4556
rect 1557 4516 1563 4556
rect 1567 4516 1569 4556
rect 1643 4516 1645 4556
rect 1649 4516 1651 4556
rect 1663 4516 1665 4556
rect 1669 4516 1671 4556
rect 1683 4516 1685 4556
rect 1689 4516 1691 4556
rect 1703 4516 1705 4556
rect 1709 4516 1711 4556
rect 1753 4516 1755 4556
rect 1759 4536 1761 4556
rect 1773 4536 1775 4556
rect 1779 4536 1785 4556
rect 1789 4536 1793 4556
rect 1805 4536 1807 4556
rect 1811 4536 1817 4556
rect 1821 4536 1823 4556
rect 1835 4536 1839 4556
rect 1843 4536 1845 4556
rect 1883 4536 1885 4556
rect 1889 4536 1893 4556
rect 1897 4536 1899 4556
rect 1911 4536 1913 4556
rect 1917 4536 1923 4556
rect 1927 4536 1929 4556
rect 1941 4536 1945 4556
rect 1759 4516 1769 4536
rect 1932 4516 1945 4536
rect 1949 4516 1951 4556
rect 1991 4516 1993 4556
rect 1997 4516 2003 4556
rect 2007 4516 2009 4556
rect 2069 4516 2071 4556
rect 2075 4536 2079 4556
rect 2091 4536 2093 4556
rect 2097 4536 2103 4556
rect 2107 4536 2109 4556
rect 2121 4536 2123 4556
rect 2127 4536 2131 4556
rect 2135 4536 2137 4556
rect 2175 4536 2177 4556
rect 2181 4536 2185 4556
rect 2197 4536 2199 4556
rect 2203 4536 2209 4556
rect 2213 4536 2215 4556
rect 2227 4536 2231 4556
rect 2235 4536 2241 4556
rect 2245 4536 2247 4556
rect 2259 4536 2261 4556
rect 2075 4516 2088 4536
rect 2251 4516 2261 4536
rect 2265 4516 2267 4556
rect 2309 4536 2311 4556
rect 2315 4536 2317 4556
rect 2369 4536 2371 4556
rect 2375 4536 2377 4556
rect 2389 4536 2391 4556
rect 2395 4536 2397 4556
rect 2449 4536 2451 4556
rect 2455 4536 2457 4556
rect 2469 4536 2471 4556
rect 2475 4536 2477 4556
rect 2529 4536 2531 4556
rect 2535 4536 2537 4556
rect 2589 4516 2591 4556
rect 2595 4536 2599 4556
rect 2611 4536 2613 4556
rect 2617 4536 2623 4556
rect 2627 4536 2629 4556
rect 2641 4536 2643 4556
rect 2647 4536 2651 4556
rect 2655 4536 2657 4556
rect 2695 4536 2697 4556
rect 2701 4536 2705 4556
rect 2717 4536 2719 4556
rect 2723 4536 2729 4556
rect 2733 4536 2735 4556
rect 2747 4536 2751 4556
rect 2755 4536 2761 4556
rect 2765 4536 2767 4556
rect 2779 4536 2781 4556
rect 2595 4516 2608 4536
rect 2771 4516 2781 4536
rect 2785 4516 2787 4556
rect 2829 4516 2831 4556
rect 2835 4528 2837 4556
rect 2849 4528 2851 4556
rect 2835 4516 2851 4528
rect 2855 4516 2857 4556
rect 2869 4516 2871 4556
rect 2875 4516 2877 4556
rect 2931 4516 2933 4556
rect 2937 4516 2943 4556
rect 2947 4516 2949 4556
rect 3023 4536 3025 4556
rect 3029 4536 3031 4556
rect 3069 4516 3071 4556
rect 3075 4528 3077 4556
rect 3089 4528 3091 4556
rect 3075 4516 3091 4528
rect 3095 4516 3097 4556
rect 3109 4516 3111 4556
rect 3115 4516 3117 4556
rect 3169 4516 3171 4556
rect 3175 4536 3179 4556
rect 3191 4536 3193 4556
rect 3197 4536 3203 4556
rect 3207 4536 3209 4556
rect 3221 4536 3223 4556
rect 3227 4536 3231 4556
rect 3235 4536 3237 4556
rect 3275 4536 3277 4556
rect 3281 4536 3285 4556
rect 3297 4536 3299 4556
rect 3303 4536 3309 4556
rect 3313 4536 3315 4556
rect 3327 4536 3331 4556
rect 3335 4536 3341 4556
rect 3345 4536 3347 4556
rect 3359 4536 3361 4556
rect 3175 4516 3188 4536
rect 3351 4516 3361 4536
rect 3365 4516 3367 4556
rect 3409 4516 3411 4556
rect 3415 4528 3417 4556
rect 3429 4528 3431 4556
rect 3415 4516 3431 4528
rect 3435 4516 3437 4556
rect 3449 4516 3451 4556
rect 3455 4516 3457 4556
rect 3523 4516 3525 4556
rect 3529 4516 3531 4556
rect 3543 4516 3545 4556
rect 3549 4528 3551 4556
rect 3563 4528 3565 4556
rect 3549 4516 3565 4528
rect 3569 4516 3571 4556
rect 3613 4516 3615 4556
rect 3619 4536 3621 4556
rect 3633 4536 3635 4556
rect 3639 4536 3645 4556
rect 3649 4536 3653 4556
rect 3665 4536 3667 4556
rect 3671 4536 3677 4556
rect 3681 4536 3683 4556
rect 3695 4536 3699 4556
rect 3703 4536 3705 4556
rect 3743 4536 3745 4556
rect 3749 4536 3753 4556
rect 3757 4536 3759 4556
rect 3771 4536 3773 4556
rect 3777 4536 3783 4556
rect 3787 4536 3789 4556
rect 3801 4536 3805 4556
rect 3619 4516 3629 4536
rect 3792 4516 3805 4536
rect 3809 4516 3811 4556
rect 3849 4516 3851 4556
rect 3855 4528 3857 4556
rect 3869 4528 3871 4556
rect 3855 4516 3871 4528
rect 3875 4516 3877 4556
rect 3889 4516 3891 4556
rect 3895 4516 3897 4556
rect 3953 4516 3955 4556
rect 3959 4536 3961 4556
rect 3973 4536 3975 4556
rect 3979 4536 3985 4556
rect 3989 4536 3993 4556
rect 4005 4536 4007 4556
rect 4011 4536 4017 4556
rect 4021 4536 4023 4556
rect 4035 4536 4039 4556
rect 4043 4536 4045 4556
rect 4083 4536 4085 4556
rect 4089 4536 4093 4556
rect 4097 4536 4099 4556
rect 4111 4536 4113 4556
rect 4117 4536 4123 4556
rect 4127 4536 4129 4556
rect 4141 4536 4145 4556
rect 3959 4516 3969 4536
rect 4132 4516 4145 4536
rect 4149 4516 4151 4556
rect 4226 4498 4228 4556
rect 4214 4496 4228 4498
rect 4232 4496 4236 4556
rect 4240 4496 4244 4556
rect 4248 4496 4250 4556
rect 4289 4516 4291 4556
rect 4295 4528 4297 4556
rect 4309 4528 4311 4556
rect 4295 4516 4311 4528
rect 4315 4516 4317 4556
rect 4329 4516 4331 4556
rect 4335 4516 4337 4556
rect 4403 4536 4405 4556
rect 4409 4536 4411 4556
rect 4423 4536 4425 4556
rect 4429 4536 4431 4556
rect 4490 4536 4492 4556
rect 4496 4536 4500 4556
rect 4512 4516 4514 4556
rect 4518 4516 4522 4556
rect 4526 4516 4528 4556
rect 4570 4496 4572 4556
rect 4576 4496 4580 4556
rect 4584 4496 4588 4556
rect 4592 4498 4594 4556
rect 4683 4536 4685 4556
rect 4689 4536 4691 4556
rect 4592 4496 4606 4498
rect 4729 4516 4731 4556
rect 4735 4528 4737 4556
rect 4749 4528 4751 4556
rect 4735 4516 4751 4528
rect 4755 4516 4757 4556
rect 4769 4516 4771 4556
rect 4775 4516 4777 4556
rect 4843 4516 4845 4556
rect 4849 4536 4851 4556
rect 4863 4536 4865 4556
rect 4869 4536 4871 4556
rect 4883 4536 4885 4556
rect 4889 4536 4891 4556
rect 4849 4516 4861 4536
rect 4951 4516 4953 4556
rect 4957 4516 4963 4556
rect 4967 4516 4969 4556
rect 5046 4498 5048 4556
rect 5034 4496 5048 4498
rect 5052 4496 5056 4556
rect 5060 4496 5064 4556
rect 5068 4496 5070 4556
rect 5109 4516 5111 4556
rect 5115 4528 5117 4556
rect 5129 4528 5131 4556
rect 5115 4516 5131 4528
rect 5135 4516 5137 4556
rect 5149 4516 5151 4556
rect 5155 4516 5157 4556
rect 5223 4516 5225 4556
rect 5229 4536 5231 4556
rect 5243 4536 5245 4556
rect 5249 4536 5251 4556
rect 5263 4536 5265 4556
rect 5269 4536 5271 4556
rect 5229 4516 5241 4536
rect 5309 4516 5311 4556
rect 5315 4528 5317 4556
rect 5329 4528 5331 4556
rect 5315 4516 5331 4528
rect 5335 4516 5337 4556
rect 5349 4516 5351 4556
rect 5355 4516 5357 4556
rect 5409 4536 5411 4556
rect 5415 4536 5417 4556
rect 5506 4498 5508 4556
rect 5494 4496 5508 4498
rect 5512 4496 5516 4556
rect 5520 4496 5524 4556
rect 5528 4496 5530 4556
rect 5571 4516 5573 4556
rect 5577 4516 5583 4556
rect 5587 4516 5589 4556
rect 5649 4516 5651 4556
rect 5655 4528 5657 4556
rect 5669 4528 5671 4556
rect 5655 4516 5671 4528
rect 5675 4516 5677 4556
rect 5689 4516 5691 4556
rect 5695 4516 5697 4556
rect 5771 4516 5773 4556
rect 5777 4516 5783 4556
rect 5787 4516 5789 4556
rect 5866 4498 5868 4556
rect 5854 4496 5868 4498
rect 5872 4496 5876 4556
rect 5880 4496 5884 4556
rect 5888 4496 5890 4556
rect 5943 4516 5945 4556
rect 5949 4516 5951 4556
rect 5963 4516 5965 4556
rect 5969 4528 5971 4556
rect 5983 4528 5985 4556
rect 5969 4516 5985 4528
rect 5989 4516 5991 4556
rect 6029 4536 6031 4556
rect 6035 4536 6037 4556
rect 6103 4536 6105 4556
rect 6109 4536 6111 4556
rect 6150 4496 6152 4556
rect 6156 4496 6160 4556
rect 6164 4496 6168 4556
rect 6172 4498 6174 4556
rect 6263 4516 6265 4556
rect 6269 4516 6271 4556
rect 6283 4516 6285 4556
rect 6289 4528 6291 4556
rect 6303 4528 6305 4556
rect 6289 4516 6305 4528
rect 6309 4516 6311 4556
rect 6172 4496 6186 4498
rect 6350 4496 6352 4556
rect 6356 4496 6360 4556
rect 6364 4496 6368 4556
rect 6372 4498 6374 4556
rect 6372 4496 6386 4498
rect 6450 4496 6452 4556
rect 6456 4496 6460 4556
rect 6464 4496 6468 4556
rect 6472 4498 6474 4556
rect 6549 4516 6551 4556
rect 6555 4528 6557 4556
rect 6569 4528 6571 4556
rect 6555 4516 6571 4528
rect 6575 4516 6577 4556
rect 6589 4516 6591 4556
rect 6595 4516 6597 4556
rect 6649 4536 6651 4556
rect 6655 4536 6657 4556
rect 6472 4496 6486 4498
rect 41 4104 43 4144
rect 47 4104 49 4144
rect 61 4104 65 4124
rect 69 4104 71 4124
rect 123 4104 125 4144
rect 129 4104 131 4144
rect 143 4104 145 4144
rect 149 4132 165 4144
rect 149 4104 151 4132
rect 163 4104 165 4132
rect 169 4104 171 4144
rect 209 4104 211 4144
rect 215 4132 231 4144
rect 215 4104 217 4132
rect 229 4104 231 4132
rect 235 4104 237 4144
rect 249 4104 251 4144
rect 255 4104 257 4144
rect 313 4104 315 4144
rect 319 4124 329 4144
rect 492 4124 505 4144
rect 319 4104 321 4124
rect 333 4104 335 4124
rect 339 4104 345 4124
rect 349 4104 353 4124
rect 365 4104 367 4124
rect 371 4104 377 4124
rect 381 4104 383 4124
rect 395 4104 399 4124
rect 403 4104 405 4124
rect 443 4104 445 4124
rect 449 4104 453 4124
rect 457 4104 459 4124
rect 471 4104 473 4124
rect 477 4104 483 4124
rect 487 4104 489 4124
rect 501 4104 505 4124
rect 509 4104 511 4144
rect 551 4104 553 4144
rect 557 4104 563 4144
rect 567 4104 569 4144
rect 664 4104 666 4144
rect 670 4104 674 4144
rect 678 4104 680 4144
rect 692 4104 694 4144
rect 698 4104 702 4144
rect 706 4104 708 4144
rect 763 4104 765 4124
rect 769 4104 771 4124
rect 809 4104 811 4144
rect 815 4124 828 4144
rect 991 4124 1001 4144
rect 815 4104 819 4124
rect 831 4104 833 4124
rect 837 4104 843 4124
rect 847 4104 849 4124
rect 861 4104 863 4124
rect 867 4104 871 4124
rect 875 4104 877 4124
rect 915 4104 917 4124
rect 921 4104 925 4124
rect 937 4104 939 4124
rect 943 4104 949 4124
rect 953 4104 955 4124
rect 967 4104 971 4124
rect 975 4104 981 4124
rect 985 4104 987 4124
rect 999 4104 1001 4124
rect 1005 4104 1007 4144
rect 1051 4104 1053 4144
rect 1057 4104 1063 4144
rect 1067 4104 1069 4144
rect 1129 4104 1131 4144
rect 1135 4124 1148 4144
rect 1311 4124 1321 4144
rect 1135 4104 1139 4124
rect 1151 4104 1153 4124
rect 1157 4104 1163 4124
rect 1167 4104 1169 4124
rect 1181 4104 1183 4124
rect 1187 4104 1191 4124
rect 1195 4104 1197 4124
rect 1235 4104 1237 4124
rect 1241 4104 1245 4124
rect 1257 4104 1259 4124
rect 1263 4104 1269 4124
rect 1273 4104 1275 4124
rect 1287 4104 1291 4124
rect 1295 4104 1301 4124
rect 1305 4104 1307 4124
rect 1319 4104 1321 4124
rect 1325 4104 1327 4144
rect 1371 4104 1373 4144
rect 1377 4104 1383 4144
rect 1387 4104 1389 4144
rect 1449 4104 1451 4124
rect 1455 4104 1457 4124
rect 1523 4104 1525 4144
rect 1529 4104 1531 4144
rect 1543 4104 1545 4144
rect 1549 4132 1565 4144
rect 1549 4104 1551 4132
rect 1563 4104 1565 4132
rect 1569 4104 1571 4144
rect 1630 4104 1632 4124
rect 1636 4104 1640 4124
rect 1652 4104 1654 4144
rect 1658 4104 1662 4144
rect 1666 4104 1668 4144
rect 1731 4104 1733 4144
rect 1737 4104 1743 4144
rect 1747 4104 1749 4144
rect 1791 4104 1793 4144
rect 1797 4104 1803 4144
rect 1807 4104 1809 4144
rect 1869 4104 1871 4144
rect 1875 4124 1888 4144
rect 2051 4124 2061 4144
rect 1875 4104 1879 4124
rect 1891 4104 1893 4124
rect 1897 4104 1903 4124
rect 1907 4104 1909 4124
rect 1921 4104 1923 4124
rect 1927 4104 1931 4124
rect 1935 4104 1937 4124
rect 1975 4104 1977 4124
rect 1981 4104 1985 4124
rect 1997 4104 1999 4124
rect 2003 4104 2009 4124
rect 2013 4104 2015 4124
rect 2027 4104 2031 4124
rect 2035 4104 2041 4124
rect 2045 4104 2047 4124
rect 2059 4104 2061 4124
rect 2065 4104 2067 4144
rect 2111 4104 2113 4144
rect 2117 4104 2123 4144
rect 2127 4104 2129 4144
rect 2203 4104 2205 4144
rect 2209 4104 2211 4144
rect 2223 4104 2225 4144
rect 2229 4132 2245 4144
rect 2229 4104 2231 4132
rect 2243 4104 2245 4132
rect 2249 4104 2251 4144
rect 2293 4104 2295 4144
rect 2299 4124 2309 4144
rect 2472 4124 2485 4144
rect 2299 4104 2301 4124
rect 2313 4104 2315 4124
rect 2319 4104 2325 4124
rect 2329 4104 2333 4124
rect 2345 4104 2347 4124
rect 2351 4104 2357 4124
rect 2361 4104 2363 4124
rect 2375 4104 2379 4124
rect 2383 4104 2385 4124
rect 2423 4104 2425 4124
rect 2429 4104 2433 4124
rect 2437 4104 2439 4124
rect 2451 4104 2453 4124
rect 2457 4104 2463 4124
rect 2467 4104 2469 4124
rect 2481 4104 2485 4124
rect 2489 4104 2491 4144
rect 2543 4104 2545 4124
rect 2549 4104 2551 4124
rect 2563 4104 2565 4124
rect 2569 4104 2571 4124
rect 2609 4104 2611 4124
rect 2615 4104 2617 4124
rect 2669 4104 2671 4144
rect 2675 4132 2691 4144
rect 2675 4104 2677 4132
rect 2689 4104 2691 4132
rect 2695 4104 2697 4144
rect 2709 4104 2711 4144
rect 2715 4104 2717 4144
rect 2771 4104 2773 4144
rect 2777 4104 2783 4144
rect 2787 4104 2789 4144
rect 2863 4104 2865 4144
rect 2869 4104 2871 4144
rect 2883 4104 2885 4144
rect 2889 4132 2905 4144
rect 2889 4104 2891 4132
rect 2903 4104 2905 4132
rect 2909 4104 2911 4144
rect 2949 4104 2951 4124
rect 2955 4104 2957 4124
rect 3009 4104 3011 4124
rect 3015 4104 3017 4124
rect 3029 4104 3031 4124
rect 3035 4104 3037 4124
rect 3103 4104 3105 4124
rect 3109 4104 3111 4124
rect 3149 4104 3151 4144
rect 3155 4124 3168 4144
rect 3331 4124 3341 4144
rect 3155 4104 3159 4124
rect 3171 4104 3173 4124
rect 3177 4104 3183 4124
rect 3187 4104 3189 4124
rect 3201 4104 3203 4124
rect 3207 4104 3211 4124
rect 3215 4104 3217 4124
rect 3255 4104 3257 4124
rect 3261 4104 3265 4124
rect 3277 4104 3279 4124
rect 3283 4104 3289 4124
rect 3293 4104 3295 4124
rect 3307 4104 3311 4124
rect 3315 4104 3321 4124
rect 3325 4104 3327 4124
rect 3339 4104 3341 4124
rect 3345 4104 3347 4144
rect 3389 4104 3391 4144
rect 3395 4134 3411 4144
rect 3395 4104 3397 4134
rect 3409 4104 3411 4134
rect 3415 4104 3417 4144
rect 3429 4104 3431 4144
rect 3435 4116 3437 4144
rect 3449 4116 3451 4144
rect 3435 4104 3451 4116
rect 3455 4104 3457 4144
rect 3511 4104 3513 4144
rect 3517 4104 3523 4144
rect 3527 4104 3529 4144
rect 3589 4104 3591 4144
rect 3595 4104 3597 4144
rect 3609 4104 3611 4144
rect 3615 4104 3617 4144
rect 3629 4104 3631 4144
rect 3635 4104 3637 4144
rect 3649 4104 3651 4144
rect 3655 4104 3657 4144
rect 3669 4104 3671 4144
rect 3675 4104 3677 4144
rect 3689 4104 3691 4144
rect 3695 4104 3697 4144
rect 3709 4104 3711 4144
rect 3715 4104 3717 4144
rect 3729 4104 3731 4144
rect 3735 4104 3737 4144
rect 3791 4104 3793 4144
rect 3797 4104 3803 4144
rect 3807 4104 3809 4144
rect 3871 4104 3873 4144
rect 3877 4104 3883 4144
rect 3887 4104 3889 4144
rect 3971 4104 3973 4144
rect 3977 4104 3983 4144
rect 3987 4104 3989 4144
rect 4029 4104 4031 4124
rect 4035 4104 4037 4124
rect 4103 4104 4105 4144
rect 4109 4104 4111 4144
rect 4123 4104 4125 4144
rect 4129 4132 4145 4144
rect 4129 4104 4131 4132
rect 4143 4104 4145 4132
rect 4149 4104 4151 4144
rect 4189 4104 4191 4144
rect 4195 4132 4211 4144
rect 4195 4104 4197 4132
rect 4209 4104 4211 4132
rect 4215 4104 4217 4144
rect 4229 4104 4231 4144
rect 4235 4104 4237 4144
rect 4293 4104 4295 4144
rect 4299 4124 4309 4144
rect 4472 4124 4485 4144
rect 4299 4104 4301 4124
rect 4313 4104 4315 4124
rect 4319 4104 4325 4124
rect 4329 4104 4333 4124
rect 4345 4104 4347 4124
rect 4351 4104 4357 4124
rect 4361 4104 4363 4124
rect 4375 4104 4379 4124
rect 4383 4104 4385 4124
rect 4423 4104 4425 4124
rect 4429 4104 4433 4124
rect 4437 4104 4439 4124
rect 4451 4104 4453 4124
rect 4457 4104 4463 4124
rect 4467 4104 4469 4124
rect 4481 4104 4485 4124
rect 4489 4104 4491 4144
rect 4543 4104 4545 4144
rect 4549 4104 4551 4144
rect 4563 4104 4565 4144
rect 4569 4132 4585 4144
rect 4569 4104 4571 4132
rect 4583 4104 4585 4132
rect 4589 4104 4591 4144
rect 4633 4104 4635 4144
rect 4639 4124 4649 4144
rect 4812 4124 4825 4144
rect 4639 4104 4641 4124
rect 4653 4104 4655 4124
rect 4659 4104 4665 4124
rect 4669 4104 4673 4124
rect 4685 4104 4687 4124
rect 4691 4104 4697 4124
rect 4701 4104 4703 4124
rect 4715 4104 4719 4124
rect 4723 4104 4725 4124
rect 4763 4104 4765 4124
rect 4769 4104 4773 4124
rect 4777 4104 4779 4124
rect 4791 4104 4793 4124
rect 4797 4104 4803 4124
rect 4807 4104 4809 4124
rect 4821 4104 4825 4124
rect 4829 4104 4831 4144
rect 4883 4104 4885 4144
rect 4889 4104 4891 4144
rect 4950 4104 4952 4124
rect 4956 4104 4960 4124
rect 4972 4104 4974 4144
rect 4978 4104 4982 4144
rect 4986 4104 4988 4144
rect 5030 4104 5032 4164
rect 5036 4104 5040 4164
rect 5044 4104 5048 4164
rect 5052 4162 5066 4164
rect 5052 4104 5054 4162
rect 5143 4104 5145 4124
rect 5149 4104 5151 4124
rect 5189 4104 5191 4144
rect 5195 4132 5211 4144
rect 5195 4104 5197 4132
rect 5209 4104 5211 4132
rect 5215 4104 5217 4144
rect 5229 4104 5231 4144
rect 5235 4104 5237 4144
rect 5293 4104 5295 4144
rect 5299 4124 5309 4144
rect 5472 4124 5485 4144
rect 5299 4104 5301 4124
rect 5313 4104 5315 4124
rect 5319 4104 5325 4124
rect 5329 4104 5333 4124
rect 5345 4104 5347 4124
rect 5351 4104 5357 4124
rect 5361 4104 5363 4124
rect 5375 4104 5379 4124
rect 5383 4104 5385 4124
rect 5423 4104 5425 4124
rect 5429 4104 5433 4124
rect 5437 4104 5439 4124
rect 5451 4104 5453 4124
rect 5457 4104 5463 4124
rect 5467 4104 5469 4124
rect 5481 4104 5485 4124
rect 5489 4104 5491 4144
rect 5531 4104 5533 4144
rect 5537 4104 5543 4144
rect 5547 4104 5549 4144
rect 5609 4104 5611 4124
rect 5615 4104 5617 4124
rect 5669 4104 5671 4144
rect 5675 4132 5691 4144
rect 5675 4104 5677 4132
rect 5689 4104 5691 4132
rect 5695 4104 5697 4144
rect 5709 4104 5711 4144
rect 5715 4104 5717 4144
rect 5793 4104 5795 4144
rect 5799 4104 5801 4144
rect 5813 4104 5815 4144
rect 5819 4104 5825 4144
rect 5829 4104 5831 4144
rect 5870 4104 5872 4164
rect 5876 4104 5880 4164
rect 5884 4104 5888 4164
rect 5892 4162 5906 4164
rect 5892 4104 5894 4162
rect 5983 4104 5985 4144
rect 5989 4104 5991 4144
rect 6029 4104 6031 4144
rect 6035 4132 6051 4144
rect 6035 4104 6037 4132
rect 6049 4104 6051 4132
rect 6055 4104 6057 4144
rect 6069 4104 6071 4144
rect 6075 4104 6077 4144
rect 6129 4104 6131 4124
rect 6135 4104 6139 4124
rect 6151 4104 6153 4144
rect 6157 4104 6159 4144
rect 6211 4104 6213 4144
rect 6217 4104 6223 4144
rect 6227 4104 6229 4144
rect 6313 4104 6315 4144
rect 6319 4104 6321 4144
rect 6333 4104 6335 4144
rect 6339 4104 6345 4144
rect 6349 4104 6351 4144
rect 6391 4104 6393 4144
rect 6397 4104 6403 4144
rect 6407 4104 6409 4144
rect 6469 4104 6471 4124
rect 6475 4104 6477 4124
rect 6550 4104 6552 4124
rect 6556 4104 6560 4124
rect 6572 4104 6574 4144
rect 6578 4104 6582 4144
rect 6586 4104 6588 4144
rect 6630 4104 6632 4164
rect 6636 4104 6640 4164
rect 6644 4104 6648 4164
rect 6652 4162 6666 4164
rect 6652 4104 6654 4162
rect 41 4036 43 4076
rect 47 4036 49 4076
rect 61 4056 65 4076
rect 69 4056 71 4076
rect 109 4036 111 4076
rect 115 4056 119 4076
rect 131 4056 133 4076
rect 137 4056 143 4076
rect 147 4056 149 4076
rect 161 4056 163 4076
rect 167 4056 171 4076
rect 175 4056 177 4076
rect 215 4056 217 4076
rect 221 4056 225 4076
rect 237 4056 239 4076
rect 243 4056 249 4076
rect 253 4056 255 4076
rect 267 4056 271 4076
rect 275 4056 281 4076
rect 285 4056 287 4076
rect 299 4056 301 4076
rect 115 4036 128 4056
rect 291 4036 301 4056
rect 305 4036 307 4076
rect 351 4036 353 4076
rect 357 4036 363 4076
rect 367 4036 369 4076
rect 450 4056 452 4076
rect 456 4056 460 4076
rect 472 4036 474 4076
rect 478 4036 482 4076
rect 486 4036 488 4076
rect 551 4036 553 4076
rect 557 4036 563 4076
rect 567 4036 569 4076
rect 631 4036 633 4076
rect 637 4036 643 4076
rect 647 4036 649 4076
rect 701 4036 703 4076
rect 707 4036 709 4076
rect 721 4056 725 4076
rect 729 4056 731 4076
rect 769 4036 771 4076
rect 775 4056 779 4076
rect 791 4056 793 4076
rect 797 4056 803 4076
rect 807 4056 809 4076
rect 821 4056 823 4076
rect 827 4056 831 4076
rect 835 4056 837 4076
rect 875 4056 877 4076
rect 881 4056 885 4076
rect 897 4056 899 4076
rect 903 4056 909 4076
rect 913 4056 915 4076
rect 927 4056 931 4076
rect 935 4056 941 4076
rect 945 4056 947 4076
rect 959 4056 961 4076
rect 775 4036 788 4056
rect 951 4036 961 4056
rect 965 4036 967 4076
rect 1031 4036 1033 4076
rect 1037 4036 1043 4076
rect 1047 4036 1049 4076
rect 1091 4036 1093 4076
rect 1097 4036 1103 4076
rect 1107 4036 1109 4076
rect 1171 4036 1173 4076
rect 1177 4036 1183 4076
rect 1187 4036 1189 4076
rect 1270 4056 1272 4076
rect 1276 4056 1280 4076
rect 1292 4036 1294 4076
rect 1298 4036 1302 4076
rect 1306 4036 1308 4076
rect 1349 4036 1351 4076
rect 1355 4056 1359 4076
rect 1371 4056 1373 4076
rect 1377 4056 1383 4076
rect 1387 4056 1389 4076
rect 1401 4056 1403 4076
rect 1407 4056 1411 4076
rect 1415 4056 1417 4076
rect 1455 4056 1457 4076
rect 1461 4056 1465 4076
rect 1477 4056 1479 4076
rect 1483 4056 1489 4076
rect 1493 4056 1495 4076
rect 1507 4056 1511 4076
rect 1515 4056 1521 4076
rect 1525 4056 1527 4076
rect 1539 4056 1541 4076
rect 1355 4036 1368 4056
rect 1531 4036 1541 4056
rect 1545 4036 1547 4076
rect 1611 4036 1613 4076
rect 1617 4036 1623 4076
rect 1627 4036 1629 4076
rect 1669 4056 1671 4076
rect 1675 4056 1679 4076
rect 1691 4036 1693 4076
rect 1697 4036 1699 4076
rect 1751 4036 1753 4076
rect 1757 4036 1763 4076
rect 1767 4036 1769 4076
rect 1829 4036 1831 4076
rect 1835 4056 1839 4076
rect 1851 4056 1853 4076
rect 1857 4056 1863 4076
rect 1867 4056 1869 4076
rect 1881 4056 1883 4076
rect 1887 4056 1891 4076
rect 1895 4056 1897 4076
rect 1935 4056 1937 4076
rect 1941 4056 1945 4076
rect 1957 4056 1959 4076
rect 1963 4056 1969 4076
rect 1973 4056 1975 4076
rect 1987 4056 1991 4076
rect 1995 4056 2001 4076
rect 2005 4056 2007 4076
rect 2019 4056 2021 4076
rect 1835 4036 1848 4056
rect 2011 4036 2021 4056
rect 2025 4036 2027 4076
rect 2071 4036 2073 4076
rect 2077 4036 2083 4076
rect 2087 4036 2089 4076
rect 2163 4036 2165 4076
rect 2169 4036 2171 4076
rect 2183 4036 2185 4076
rect 2189 4048 2191 4076
rect 2203 4048 2205 4076
rect 2189 4036 2205 4048
rect 2209 4036 2211 4076
rect 2271 4036 2273 4076
rect 2277 4036 2283 4076
rect 2287 4036 2289 4076
rect 2331 4036 2333 4076
rect 2337 4036 2343 4076
rect 2347 4036 2349 4076
rect 2423 4056 2425 4076
rect 2429 4056 2431 4076
rect 2483 4036 2485 4076
rect 2489 4036 2491 4076
rect 2503 4036 2505 4076
rect 2509 4048 2511 4076
rect 2523 4048 2525 4076
rect 2509 4036 2525 4048
rect 2529 4036 2531 4076
rect 2569 4056 2571 4076
rect 2575 4056 2577 4076
rect 2589 4056 2591 4076
rect 2595 4056 2597 4076
rect 2663 4056 2665 4076
rect 2669 4056 2671 4076
rect 2683 4056 2685 4076
rect 2689 4056 2691 4076
rect 2729 4056 2731 4076
rect 2735 4056 2737 4076
rect 2803 4056 2805 4076
rect 2809 4056 2811 4076
rect 2871 4036 2873 4076
rect 2877 4036 2883 4076
rect 2887 4036 2889 4076
rect 2929 4056 2931 4076
rect 2935 4056 2937 4076
rect 2949 4056 2951 4076
rect 2955 4056 2957 4076
rect 3009 4036 3011 4076
rect 3015 4048 3017 4076
rect 3029 4048 3031 4076
rect 3015 4036 3031 4048
rect 3035 4036 3037 4076
rect 3049 4036 3051 4076
rect 3055 4036 3057 4076
rect 3109 4056 3111 4076
rect 3115 4056 3117 4076
rect 3169 4056 3171 4076
rect 3175 4056 3177 4076
rect 3189 4056 3191 4076
rect 3195 4056 3197 4076
rect 3271 4036 3273 4076
rect 3277 4036 3283 4076
rect 3287 4036 3289 4076
rect 3351 4036 3353 4076
rect 3357 4036 3363 4076
rect 3367 4036 3369 4076
rect 3413 4036 3415 4076
rect 3419 4056 3421 4076
rect 3433 4056 3435 4076
rect 3439 4056 3445 4076
rect 3449 4056 3453 4076
rect 3465 4056 3467 4076
rect 3471 4056 3477 4076
rect 3481 4056 3483 4076
rect 3495 4056 3499 4076
rect 3503 4056 3505 4076
rect 3543 4056 3545 4076
rect 3549 4056 3553 4076
rect 3557 4056 3559 4076
rect 3571 4056 3573 4076
rect 3577 4056 3583 4076
rect 3587 4056 3589 4076
rect 3601 4056 3605 4076
rect 3419 4036 3429 4056
rect 3592 4036 3605 4056
rect 3609 4036 3611 4076
rect 3663 4056 3665 4076
rect 3669 4056 3671 4076
rect 3713 4036 3715 4076
rect 3719 4056 3721 4076
rect 3733 4056 3735 4076
rect 3739 4056 3745 4076
rect 3749 4056 3753 4076
rect 3765 4056 3767 4076
rect 3771 4056 3777 4076
rect 3781 4056 3783 4076
rect 3795 4056 3799 4076
rect 3803 4056 3805 4076
rect 3843 4056 3845 4076
rect 3849 4056 3853 4076
rect 3857 4056 3859 4076
rect 3871 4056 3873 4076
rect 3877 4056 3883 4076
rect 3887 4056 3889 4076
rect 3901 4056 3905 4076
rect 3719 4036 3729 4056
rect 3892 4036 3905 4056
rect 3909 4036 3911 4076
rect 3986 4018 3988 4076
rect 3974 4016 3988 4018
rect 3992 4016 3996 4076
rect 4000 4016 4004 4076
rect 4008 4016 4010 4076
rect 4051 4036 4053 4076
rect 4057 4036 4063 4076
rect 4067 4036 4069 4076
rect 4143 4036 4145 4076
rect 4149 4036 4151 4076
rect 4163 4036 4165 4076
rect 4169 4048 4171 4076
rect 4183 4048 4185 4076
rect 4169 4036 4185 4048
rect 4189 4036 4191 4076
rect 4229 4056 4231 4076
rect 4235 4056 4237 4076
rect 4249 4056 4251 4076
rect 4255 4056 4257 4076
rect 4323 4056 4325 4076
rect 4329 4056 4331 4076
rect 4391 4036 4393 4076
rect 4397 4036 4403 4076
rect 4407 4036 4409 4076
rect 4463 4036 4465 4076
rect 4469 4036 4471 4076
rect 4483 4036 4485 4076
rect 4489 4048 4491 4076
rect 4503 4048 4505 4076
rect 4489 4036 4505 4048
rect 4509 4036 4511 4076
rect 4553 4036 4555 4076
rect 4559 4056 4561 4076
rect 4573 4056 4575 4076
rect 4579 4056 4585 4076
rect 4589 4056 4593 4076
rect 4605 4056 4607 4076
rect 4611 4056 4617 4076
rect 4621 4056 4623 4076
rect 4635 4056 4639 4076
rect 4643 4056 4645 4076
rect 4683 4056 4685 4076
rect 4689 4056 4693 4076
rect 4697 4056 4699 4076
rect 4711 4056 4713 4076
rect 4717 4056 4723 4076
rect 4727 4056 4729 4076
rect 4741 4056 4745 4076
rect 4559 4036 4569 4056
rect 4732 4036 4745 4056
rect 4749 4036 4751 4076
rect 4811 4036 4813 4076
rect 4817 4036 4823 4076
rect 4827 4036 4829 4076
rect 4883 4036 4885 4076
rect 4889 4036 4891 4076
rect 4903 4036 4905 4076
rect 4909 4048 4911 4076
rect 4923 4048 4925 4076
rect 4909 4036 4925 4048
rect 4929 4036 4931 4076
rect 4973 4036 4975 4076
rect 4979 4056 4981 4076
rect 4993 4056 4995 4076
rect 4999 4056 5005 4076
rect 5009 4056 5013 4076
rect 5025 4056 5027 4076
rect 5031 4056 5037 4076
rect 5041 4056 5043 4076
rect 5055 4056 5059 4076
rect 5063 4056 5065 4076
rect 5103 4056 5105 4076
rect 5109 4056 5113 4076
rect 5117 4056 5119 4076
rect 5131 4056 5133 4076
rect 5137 4056 5143 4076
rect 5147 4056 5149 4076
rect 5161 4056 5165 4076
rect 4979 4036 4989 4056
rect 5152 4036 5165 4056
rect 5169 4036 5171 4076
rect 5231 4036 5233 4076
rect 5237 4036 5243 4076
rect 5247 4036 5249 4076
rect 5303 4036 5305 4076
rect 5309 4036 5311 4076
rect 5323 4036 5325 4076
rect 5329 4048 5331 4076
rect 5343 4048 5345 4076
rect 5329 4036 5345 4048
rect 5349 4036 5351 4076
rect 5411 4036 5413 4076
rect 5417 4036 5423 4076
rect 5427 4036 5429 4076
rect 5469 4036 5471 4076
rect 5475 4048 5477 4076
rect 5489 4048 5491 4076
rect 5475 4036 5491 4048
rect 5495 4036 5497 4076
rect 5509 4036 5511 4076
rect 5515 4036 5517 4076
rect 5583 4056 5585 4076
rect 5589 4056 5591 4076
rect 5633 4036 5635 4076
rect 5639 4056 5641 4076
rect 5653 4056 5655 4076
rect 5659 4056 5665 4076
rect 5669 4056 5673 4076
rect 5685 4056 5687 4076
rect 5691 4056 5697 4076
rect 5701 4056 5703 4076
rect 5715 4056 5719 4076
rect 5723 4056 5725 4076
rect 5763 4056 5765 4076
rect 5769 4056 5773 4076
rect 5777 4056 5779 4076
rect 5791 4056 5793 4076
rect 5797 4056 5803 4076
rect 5807 4056 5809 4076
rect 5821 4056 5825 4076
rect 5639 4036 5649 4056
rect 5812 4036 5825 4056
rect 5829 4036 5831 4076
rect 5869 4056 5871 4076
rect 5875 4056 5877 4076
rect 5966 4018 5968 4076
rect 5954 4016 5968 4018
rect 5972 4016 5976 4076
rect 5980 4016 5984 4076
rect 5988 4016 5990 4076
rect 6029 4036 6031 4076
rect 6035 4056 6039 4076
rect 6051 4056 6053 4076
rect 6057 4056 6063 4076
rect 6067 4056 6069 4076
rect 6081 4056 6083 4076
rect 6087 4056 6091 4076
rect 6095 4056 6097 4076
rect 6135 4056 6137 4076
rect 6141 4056 6145 4076
rect 6157 4056 6159 4076
rect 6163 4056 6169 4076
rect 6173 4056 6175 4076
rect 6187 4056 6191 4076
rect 6195 4056 6201 4076
rect 6205 4056 6207 4076
rect 6219 4056 6221 4076
rect 6035 4036 6048 4056
rect 6211 4036 6221 4056
rect 6225 4036 6227 4076
rect 6269 4036 6271 4076
rect 6275 4056 6279 4076
rect 6291 4056 6293 4076
rect 6297 4056 6303 4076
rect 6307 4056 6309 4076
rect 6321 4056 6323 4076
rect 6327 4056 6331 4076
rect 6335 4056 6337 4076
rect 6375 4056 6377 4076
rect 6381 4056 6385 4076
rect 6397 4056 6399 4076
rect 6403 4056 6409 4076
rect 6413 4056 6415 4076
rect 6427 4056 6431 4076
rect 6435 4056 6441 4076
rect 6445 4056 6447 4076
rect 6459 4056 6461 4076
rect 6275 4036 6288 4056
rect 6451 4036 6461 4056
rect 6465 4036 6467 4076
rect 6509 4036 6511 4076
rect 6515 4056 6519 4076
rect 6531 4056 6533 4076
rect 6537 4056 6543 4076
rect 6547 4056 6549 4076
rect 6561 4056 6563 4076
rect 6567 4056 6571 4076
rect 6575 4056 6577 4076
rect 6615 4056 6617 4076
rect 6621 4056 6625 4076
rect 6637 4056 6639 4076
rect 6643 4056 6649 4076
rect 6653 4056 6655 4076
rect 6667 4056 6671 4076
rect 6675 4056 6681 4076
rect 6685 4056 6687 4076
rect 6699 4056 6701 4076
rect 6515 4036 6528 4056
rect 6691 4036 6701 4056
rect 6705 4036 6707 4076
rect 41 3624 43 3664
rect 47 3624 49 3664
rect 61 3624 65 3644
rect 69 3624 71 3644
rect 121 3624 123 3664
rect 127 3624 129 3664
rect 141 3624 145 3644
rect 149 3624 151 3644
rect 211 3624 213 3664
rect 217 3624 223 3664
rect 227 3624 229 3664
rect 269 3624 271 3664
rect 275 3644 288 3664
rect 451 3644 461 3664
rect 275 3624 279 3644
rect 291 3624 293 3644
rect 297 3624 303 3644
rect 307 3624 309 3644
rect 321 3624 323 3644
rect 327 3624 331 3644
rect 335 3624 337 3644
rect 375 3624 377 3644
rect 381 3624 385 3644
rect 397 3624 399 3644
rect 403 3624 409 3644
rect 413 3624 415 3644
rect 427 3624 431 3644
rect 435 3624 441 3644
rect 445 3624 447 3644
rect 459 3624 461 3644
rect 465 3624 467 3664
rect 530 3624 532 3644
rect 536 3624 540 3644
rect 552 3624 554 3664
rect 558 3624 562 3664
rect 566 3624 568 3664
rect 631 3624 633 3664
rect 637 3624 643 3664
rect 647 3624 649 3664
rect 691 3624 693 3664
rect 697 3624 703 3664
rect 707 3624 709 3664
rect 791 3624 793 3664
rect 797 3624 803 3664
rect 807 3624 809 3664
rect 849 3624 851 3664
rect 855 3644 868 3664
rect 1031 3644 1041 3664
rect 855 3624 859 3644
rect 871 3624 873 3644
rect 877 3624 883 3644
rect 887 3624 889 3644
rect 901 3624 903 3644
rect 907 3624 911 3644
rect 915 3624 917 3644
rect 955 3624 957 3644
rect 961 3624 965 3644
rect 977 3624 979 3644
rect 983 3624 989 3644
rect 993 3624 995 3644
rect 1007 3624 1011 3644
rect 1015 3624 1021 3644
rect 1025 3624 1027 3644
rect 1039 3624 1041 3644
rect 1045 3624 1047 3664
rect 1092 3624 1094 3664
rect 1098 3624 1102 3664
rect 1106 3624 1108 3664
rect 1120 3624 1124 3644
rect 1128 3624 1130 3644
rect 1211 3624 1213 3664
rect 1217 3624 1223 3664
rect 1227 3624 1229 3664
rect 1269 3624 1271 3644
rect 1275 3624 1279 3644
rect 1291 3624 1293 3664
rect 1297 3624 1299 3664
rect 1370 3624 1372 3644
rect 1376 3624 1380 3644
rect 1392 3624 1394 3664
rect 1398 3624 1402 3664
rect 1406 3624 1408 3664
rect 1471 3624 1473 3664
rect 1477 3624 1483 3664
rect 1487 3624 1489 3664
rect 1531 3624 1533 3664
rect 1537 3624 1543 3664
rect 1547 3624 1549 3664
rect 1609 3624 1611 3644
rect 1615 3624 1617 3644
rect 1629 3624 1631 3644
rect 1635 3624 1637 3644
rect 1689 3624 1691 3664
rect 1695 3644 1708 3664
rect 1871 3644 1881 3664
rect 1695 3624 1699 3644
rect 1711 3624 1713 3644
rect 1717 3624 1723 3644
rect 1727 3624 1729 3644
rect 1741 3624 1743 3644
rect 1747 3624 1751 3644
rect 1755 3624 1757 3644
rect 1795 3624 1797 3644
rect 1801 3624 1805 3644
rect 1817 3624 1819 3644
rect 1823 3624 1829 3644
rect 1833 3624 1835 3644
rect 1847 3624 1851 3644
rect 1855 3624 1861 3644
rect 1865 3624 1867 3644
rect 1879 3624 1881 3644
rect 1885 3624 1887 3664
rect 1951 3624 1953 3664
rect 1957 3624 1963 3664
rect 1967 3624 1969 3664
rect 2009 3624 2011 3644
rect 2015 3624 2017 3644
rect 2029 3624 2031 3644
rect 2035 3624 2037 3644
rect 2089 3624 2091 3644
rect 2095 3624 2097 3644
rect 2149 3624 2151 3664
rect 2155 3652 2171 3664
rect 2155 3624 2157 3652
rect 2169 3624 2171 3652
rect 2175 3624 2177 3664
rect 2189 3624 2191 3664
rect 2195 3624 2197 3664
rect 2263 3624 2265 3664
rect 2269 3624 2271 3664
rect 2283 3624 2285 3664
rect 2289 3652 2305 3664
rect 2289 3624 2291 3652
rect 2303 3624 2305 3652
rect 2309 3624 2311 3664
rect 2370 3624 2372 3644
rect 2376 3624 2380 3644
rect 2392 3624 2394 3664
rect 2398 3624 2402 3664
rect 2406 3624 2408 3664
rect 2449 3624 2451 3644
rect 2455 3624 2457 3644
rect 2523 3624 2525 3644
rect 2529 3624 2531 3644
rect 2569 3624 2571 3664
rect 2575 3652 2591 3664
rect 2575 3624 2577 3652
rect 2589 3624 2591 3652
rect 2595 3624 2597 3664
rect 2609 3624 2611 3664
rect 2615 3624 2617 3664
rect 2670 3624 2672 3684
rect 2676 3624 2680 3684
rect 2684 3624 2688 3684
rect 2692 3682 2706 3684
rect 2692 3624 2694 3682
rect 2783 3624 2785 3644
rect 2789 3624 2791 3644
rect 2851 3624 2853 3664
rect 2857 3624 2863 3664
rect 2867 3624 2869 3664
rect 2909 3624 2911 3664
rect 2915 3652 2931 3664
rect 2915 3624 2917 3652
rect 2929 3624 2931 3652
rect 2935 3624 2937 3664
rect 2949 3624 2951 3664
rect 2955 3624 2957 3664
rect 3009 3624 3011 3664
rect 3015 3652 3031 3664
rect 3015 3624 3017 3652
rect 3029 3624 3031 3652
rect 3035 3624 3037 3664
rect 3049 3624 3051 3664
rect 3055 3624 3057 3664
rect 3112 3624 3114 3664
rect 3118 3624 3122 3664
rect 3126 3624 3128 3664
rect 3140 3624 3144 3644
rect 3148 3624 3150 3644
rect 3244 3624 3246 3664
rect 3250 3624 3254 3664
rect 3258 3624 3260 3664
rect 3272 3624 3274 3664
rect 3278 3624 3282 3664
rect 3286 3624 3288 3664
rect 3351 3624 3353 3664
rect 3357 3624 3363 3664
rect 3367 3624 3369 3664
rect 3431 3624 3433 3664
rect 3437 3624 3443 3664
rect 3447 3624 3449 3664
rect 3493 3624 3495 3664
rect 3499 3644 3509 3664
rect 3672 3644 3685 3664
rect 3499 3624 3501 3644
rect 3513 3624 3515 3644
rect 3519 3624 3525 3644
rect 3529 3624 3533 3644
rect 3545 3624 3547 3644
rect 3551 3624 3557 3644
rect 3561 3624 3563 3644
rect 3575 3624 3579 3644
rect 3583 3624 3585 3644
rect 3623 3624 3625 3644
rect 3629 3624 3633 3644
rect 3637 3624 3639 3644
rect 3651 3624 3653 3644
rect 3657 3624 3663 3644
rect 3667 3624 3669 3644
rect 3681 3624 3685 3644
rect 3689 3624 3691 3664
rect 3751 3624 3753 3664
rect 3757 3624 3763 3664
rect 3767 3624 3769 3664
rect 3844 3624 3846 3664
rect 3850 3624 3854 3664
rect 3858 3624 3860 3664
rect 3872 3624 3874 3664
rect 3878 3624 3882 3664
rect 3886 3624 3888 3664
rect 3929 3624 3931 3644
rect 3935 3624 3937 3644
rect 3991 3624 3993 3664
rect 3997 3624 4003 3664
rect 4007 3624 4009 3664
rect 4069 3624 4071 3664
rect 4075 3652 4091 3664
rect 4075 3624 4077 3652
rect 4089 3624 4091 3652
rect 4095 3624 4097 3664
rect 4109 3624 4111 3664
rect 4115 3624 4117 3664
rect 4173 3624 4175 3664
rect 4179 3644 4189 3664
rect 4352 3644 4365 3664
rect 4179 3624 4181 3644
rect 4193 3624 4195 3644
rect 4199 3624 4205 3644
rect 4209 3624 4213 3644
rect 4225 3624 4227 3644
rect 4231 3624 4237 3644
rect 4241 3624 4243 3644
rect 4255 3624 4259 3644
rect 4263 3624 4265 3644
rect 4303 3624 4305 3644
rect 4309 3624 4313 3644
rect 4317 3624 4319 3644
rect 4331 3624 4333 3644
rect 4337 3624 4343 3644
rect 4347 3624 4349 3644
rect 4361 3624 4365 3644
rect 4369 3624 4371 3664
rect 4411 3624 4413 3664
rect 4417 3624 4423 3664
rect 4427 3624 4429 3664
rect 4511 3624 4513 3664
rect 4517 3624 4523 3664
rect 4527 3624 4529 3664
rect 4583 3624 4585 3664
rect 4589 3624 4591 3664
rect 4603 3624 4605 3664
rect 4609 3624 4611 3664
rect 4623 3624 4625 3664
rect 4629 3624 4631 3664
rect 4643 3624 4645 3664
rect 4649 3624 4651 3664
rect 4663 3624 4665 3664
rect 4669 3624 4671 3664
rect 4683 3624 4685 3664
rect 4689 3624 4691 3664
rect 4703 3624 4705 3664
rect 4709 3624 4711 3664
rect 4723 3624 4725 3664
rect 4729 3624 4731 3664
rect 4773 3624 4775 3664
rect 4779 3644 4789 3664
rect 4952 3644 4965 3664
rect 4779 3624 4781 3644
rect 4793 3624 4795 3644
rect 4799 3624 4805 3644
rect 4809 3624 4813 3644
rect 4825 3624 4827 3644
rect 4831 3624 4837 3644
rect 4841 3624 4843 3644
rect 4855 3624 4859 3644
rect 4863 3624 4865 3644
rect 4903 3624 4905 3644
rect 4909 3624 4913 3644
rect 4917 3624 4919 3644
rect 4931 3624 4933 3644
rect 4937 3624 4943 3644
rect 4947 3624 4949 3644
rect 4961 3624 4965 3644
rect 4969 3624 4971 3664
rect 5009 3624 5011 3664
rect 5015 3652 5031 3664
rect 5015 3624 5017 3652
rect 5029 3624 5031 3652
rect 5035 3624 5037 3664
rect 5049 3624 5051 3664
rect 5055 3624 5057 3664
rect 5131 3624 5133 3664
rect 5137 3624 5143 3664
rect 5147 3624 5149 3664
rect 5211 3624 5213 3664
rect 5217 3624 5223 3664
rect 5227 3624 5229 3664
rect 5283 3624 5285 3644
rect 5289 3624 5291 3644
rect 5329 3624 5331 3664
rect 5335 3624 5337 3664
rect 5349 3624 5351 3664
rect 5355 3624 5357 3664
rect 5369 3624 5371 3664
rect 5375 3624 5377 3664
rect 5389 3624 5391 3664
rect 5395 3624 5397 3664
rect 5409 3624 5411 3664
rect 5415 3624 5417 3664
rect 5429 3624 5431 3664
rect 5435 3624 5437 3664
rect 5449 3624 5451 3664
rect 5455 3624 5457 3664
rect 5469 3624 5471 3664
rect 5475 3624 5477 3664
rect 5529 3624 5531 3664
rect 5535 3644 5548 3664
rect 5711 3644 5721 3664
rect 5535 3624 5539 3644
rect 5551 3624 5553 3644
rect 5557 3624 5563 3644
rect 5567 3624 5569 3644
rect 5581 3624 5583 3644
rect 5587 3624 5591 3644
rect 5595 3624 5597 3644
rect 5635 3624 5637 3644
rect 5641 3624 5645 3644
rect 5657 3624 5659 3644
rect 5663 3624 5669 3644
rect 5673 3624 5675 3644
rect 5687 3624 5691 3644
rect 5695 3624 5701 3644
rect 5705 3624 5707 3644
rect 5719 3624 5721 3644
rect 5725 3624 5727 3664
rect 5783 3624 5785 3644
rect 5789 3624 5791 3644
rect 5831 3624 5833 3664
rect 5837 3624 5843 3664
rect 5847 3624 5849 3664
rect 5911 3624 5913 3664
rect 5917 3624 5923 3664
rect 5927 3624 5929 3664
rect 6003 3624 6005 3644
rect 6009 3624 6011 3644
rect 6049 3624 6051 3644
rect 6055 3624 6057 3644
rect 6069 3624 6071 3644
rect 6075 3624 6077 3644
rect 6143 3624 6145 3644
rect 6149 3624 6151 3644
rect 6163 3624 6165 3644
rect 6169 3624 6171 3644
rect 6212 3624 6214 3664
rect 6218 3624 6222 3664
rect 6226 3624 6228 3664
rect 6240 3624 6244 3644
rect 6248 3624 6250 3644
rect 6309 3624 6311 3664
rect 6315 3644 6328 3664
rect 6491 3644 6501 3664
rect 6315 3624 6319 3644
rect 6331 3624 6333 3644
rect 6337 3624 6343 3644
rect 6347 3624 6349 3644
rect 6361 3624 6363 3644
rect 6367 3624 6371 3644
rect 6375 3624 6377 3644
rect 6415 3624 6417 3644
rect 6421 3624 6425 3644
rect 6437 3624 6439 3644
rect 6443 3624 6449 3644
rect 6453 3624 6455 3644
rect 6467 3624 6471 3644
rect 6475 3624 6481 3644
rect 6485 3624 6487 3644
rect 6499 3624 6501 3644
rect 6505 3624 6507 3664
rect 6549 3624 6551 3664
rect 6555 3652 6571 3664
rect 6555 3624 6557 3652
rect 6569 3624 6571 3652
rect 6575 3624 6577 3664
rect 6589 3624 6591 3664
rect 6595 3624 6597 3664
rect 6651 3624 6653 3664
rect 6657 3624 6663 3664
rect 6667 3624 6669 3664
rect 41 3556 43 3596
rect 47 3556 49 3596
rect 61 3576 65 3596
rect 69 3576 71 3596
rect 109 3556 111 3596
rect 115 3576 119 3596
rect 131 3576 133 3596
rect 137 3576 143 3596
rect 147 3576 149 3596
rect 161 3576 163 3596
rect 167 3576 171 3596
rect 175 3576 177 3596
rect 215 3576 217 3596
rect 221 3576 225 3596
rect 237 3576 239 3596
rect 243 3576 249 3596
rect 253 3576 255 3596
rect 267 3576 271 3596
rect 275 3576 281 3596
rect 285 3576 287 3596
rect 299 3576 301 3596
rect 115 3556 128 3576
rect 291 3556 301 3576
rect 305 3556 307 3596
rect 351 3556 353 3596
rect 357 3556 363 3596
rect 367 3556 369 3596
rect 429 3576 431 3596
rect 435 3576 439 3596
rect 451 3556 453 3596
rect 457 3556 459 3596
rect 530 3576 532 3596
rect 536 3576 540 3596
rect 552 3556 554 3596
rect 558 3556 562 3596
rect 566 3556 568 3596
rect 631 3556 633 3596
rect 637 3556 643 3596
rect 647 3556 649 3596
rect 701 3556 703 3596
rect 707 3556 709 3596
rect 721 3576 725 3596
rect 729 3576 731 3596
rect 769 3576 771 3596
rect 775 3576 779 3596
rect 791 3556 793 3596
rect 797 3556 799 3596
rect 851 3556 853 3596
rect 857 3556 863 3596
rect 867 3556 869 3596
rect 941 3556 943 3596
rect 947 3556 949 3596
rect 961 3576 965 3596
rect 969 3576 971 3596
rect 1023 3576 1025 3596
rect 1029 3576 1031 3596
rect 1081 3556 1083 3596
rect 1087 3556 1089 3596
rect 1101 3576 1105 3596
rect 1109 3576 1111 3596
rect 1161 3556 1163 3596
rect 1167 3556 1169 3596
rect 1181 3576 1185 3596
rect 1189 3576 1191 3596
rect 1229 3556 1231 3596
rect 1235 3576 1239 3596
rect 1251 3576 1253 3596
rect 1257 3576 1263 3596
rect 1267 3576 1269 3596
rect 1281 3576 1283 3596
rect 1287 3576 1291 3596
rect 1295 3576 1297 3596
rect 1335 3576 1337 3596
rect 1341 3576 1345 3596
rect 1357 3576 1359 3596
rect 1363 3576 1369 3596
rect 1373 3576 1375 3596
rect 1387 3576 1391 3596
rect 1395 3576 1401 3596
rect 1405 3576 1407 3596
rect 1419 3576 1421 3596
rect 1235 3556 1248 3576
rect 1411 3556 1421 3576
rect 1425 3556 1427 3596
rect 1483 3576 1485 3596
rect 1489 3576 1491 3596
rect 1503 3576 1505 3596
rect 1509 3576 1511 3596
rect 1549 3556 1551 3596
rect 1555 3576 1559 3596
rect 1571 3576 1573 3596
rect 1577 3576 1583 3596
rect 1587 3576 1589 3596
rect 1601 3576 1603 3596
rect 1607 3576 1611 3596
rect 1615 3576 1617 3596
rect 1655 3576 1657 3596
rect 1661 3576 1665 3596
rect 1677 3576 1679 3596
rect 1683 3576 1689 3596
rect 1693 3576 1695 3596
rect 1707 3576 1711 3596
rect 1715 3576 1721 3596
rect 1725 3576 1727 3596
rect 1739 3576 1741 3596
rect 1555 3556 1568 3576
rect 1731 3556 1741 3576
rect 1745 3556 1747 3596
rect 1813 3556 1815 3596
rect 1819 3556 1821 3596
rect 1833 3556 1835 3596
rect 1839 3556 1845 3596
rect 1849 3556 1851 3596
rect 1903 3576 1905 3596
rect 1909 3576 1911 3596
rect 1963 3556 1965 3596
rect 1969 3556 1971 3596
rect 1983 3556 1985 3596
rect 1989 3568 1991 3596
rect 2003 3568 2005 3596
rect 1989 3556 2005 3568
rect 2009 3556 2011 3596
rect 2049 3576 2051 3596
rect 2055 3576 2057 3596
rect 2069 3576 2071 3596
rect 2075 3576 2077 3596
rect 2143 3576 2145 3596
rect 2149 3576 2151 3596
rect 2213 3556 2215 3596
rect 2219 3556 2221 3596
rect 2233 3556 2235 3596
rect 2239 3556 2245 3596
rect 2249 3556 2251 3596
rect 2303 3576 2305 3596
rect 2309 3576 2311 3596
rect 2323 3576 2325 3596
rect 2329 3576 2331 3596
rect 2369 3556 2371 3596
rect 2375 3576 2379 3596
rect 2391 3576 2393 3596
rect 2397 3576 2403 3596
rect 2407 3576 2409 3596
rect 2421 3576 2423 3596
rect 2427 3576 2431 3596
rect 2435 3576 2437 3596
rect 2475 3576 2477 3596
rect 2481 3576 2485 3596
rect 2497 3576 2499 3596
rect 2503 3576 2509 3596
rect 2513 3576 2515 3596
rect 2527 3576 2531 3596
rect 2535 3576 2541 3596
rect 2545 3576 2547 3596
rect 2559 3576 2561 3596
rect 2375 3556 2388 3576
rect 2551 3556 2561 3576
rect 2565 3556 2567 3596
rect 2609 3576 2611 3596
rect 2615 3576 2617 3596
rect 2629 3576 2631 3596
rect 2635 3576 2637 3596
rect 2689 3556 2691 3596
rect 2695 3568 2697 3596
rect 2709 3568 2711 3596
rect 2695 3556 2711 3568
rect 2715 3556 2717 3596
rect 2729 3556 2731 3596
rect 2735 3556 2737 3596
rect 2803 3576 2805 3596
rect 2809 3576 2811 3596
rect 2871 3556 2873 3596
rect 2877 3556 2883 3596
rect 2887 3556 2889 3596
rect 2929 3556 2931 3596
rect 2935 3568 2937 3596
rect 2949 3568 2951 3596
rect 2935 3556 2951 3568
rect 2955 3556 2957 3596
rect 2969 3556 2971 3596
rect 2975 3556 2977 3596
rect 3032 3556 3034 3596
rect 3038 3556 3042 3596
rect 3046 3556 3048 3596
rect 3060 3576 3064 3596
rect 3068 3576 3070 3596
rect 3129 3556 3131 3596
rect 3135 3556 3137 3596
rect 3224 3556 3226 3596
rect 3230 3556 3234 3596
rect 3238 3556 3240 3596
rect 3252 3556 3254 3596
rect 3258 3556 3262 3596
rect 3266 3556 3268 3596
rect 3323 3576 3325 3596
rect 3329 3576 3331 3596
rect 3369 3556 3371 3596
rect 3375 3576 3379 3596
rect 3391 3576 3393 3596
rect 3397 3576 3403 3596
rect 3407 3576 3409 3596
rect 3421 3576 3423 3596
rect 3427 3576 3431 3596
rect 3435 3576 3437 3596
rect 3475 3576 3477 3596
rect 3481 3576 3485 3596
rect 3497 3576 3499 3596
rect 3503 3576 3509 3596
rect 3513 3576 3515 3596
rect 3527 3576 3531 3596
rect 3535 3576 3541 3596
rect 3545 3576 3547 3596
rect 3559 3576 3561 3596
rect 3375 3556 3388 3576
rect 3551 3556 3561 3576
rect 3565 3556 3567 3596
rect 3644 3556 3646 3596
rect 3650 3556 3654 3596
rect 3658 3556 3660 3596
rect 3672 3556 3674 3596
rect 3678 3556 3682 3596
rect 3686 3556 3688 3596
rect 3729 3556 3731 3596
rect 3735 3576 3739 3596
rect 3751 3576 3753 3596
rect 3757 3576 3763 3596
rect 3767 3576 3769 3596
rect 3781 3576 3783 3596
rect 3787 3576 3791 3596
rect 3795 3576 3797 3596
rect 3835 3576 3837 3596
rect 3841 3576 3845 3596
rect 3857 3576 3859 3596
rect 3863 3576 3869 3596
rect 3873 3576 3875 3596
rect 3887 3576 3891 3596
rect 3895 3576 3901 3596
rect 3905 3576 3907 3596
rect 3919 3576 3921 3596
rect 3735 3556 3748 3576
rect 3911 3556 3921 3576
rect 3925 3556 3927 3596
rect 3983 3576 3985 3596
rect 3989 3576 3991 3596
rect 4029 3556 4031 3596
rect 4035 3576 4039 3596
rect 4051 3576 4053 3596
rect 4057 3576 4063 3596
rect 4067 3576 4069 3596
rect 4081 3576 4083 3596
rect 4087 3576 4091 3596
rect 4095 3576 4097 3596
rect 4135 3576 4137 3596
rect 4141 3576 4145 3596
rect 4157 3576 4159 3596
rect 4163 3576 4169 3596
rect 4173 3576 4175 3596
rect 4187 3576 4191 3596
rect 4195 3576 4201 3596
rect 4205 3576 4207 3596
rect 4219 3576 4221 3596
rect 4035 3556 4048 3576
rect 4211 3556 4221 3576
rect 4225 3556 4227 3596
rect 4283 3576 4285 3596
rect 4289 3576 4291 3596
rect 4343 3576 4345 3596
rect 4349 3576 4351 3596
rect 4391 3556 4393 3596
rect 4397 3556 4403 3596
rect 4407 3556 4409 3596
rect 4473 3556 4475 3596
rect 4479 3576 4481 3596
rect 4493 3576 4495 3596
rect 4499 3576 4505 3596
rect 4509 3576 4513 3596
rect 4525 3576 4527 3596
rect 4531 3576 4537 3596
rect 4541 3576 4543 3596
rect 4555 3576 4559 3596
rect 4563 3576 4565 3596
rect 4603 3576 4605 3596
rect 4609 3576 4613 3596
rect 4617 3576 4619 3596
rect 4631 3576 4633 3596
rect 4637 3576 4643 3596
rect 4647 3576 4649 3596
rect 4661 3576 4665 3596
rect 4479 3556 4489 3576
rect 4652 3556 4665 3576
rect 4669 3556 4671 3596
rect 4723 3576 4725 3596
rect 4729 3576 4731 3596
rect 4769 3556 4771 3596
rect 4775 3576 4779 3596
rect 4791 3576 4793 3596
rect 4797 3576 4803 3596
rect 4807 3576 4809 3596
rect 4821 3576 4823 3596
rect 4827 3576 4831 3596
rect 4835 3576 4837 3596
rect 4875 3576 4877 3596
rect 4881 3576 4885 3596
rect 4897 3576 4899 3596
rect 4903 3576 4909 3596
rect 4913 3576 4915 3596
rect 4927 3576 4931 3596
rect 4935 3576 4941 3596
rect 4945 3576 4947 3596
rect 4959 3576 4961 3596
rect 4775 3556 4788 3576
rect 4951 3556 4961 3576
rect 4965 3556 4967 3596
rect 5044 3556 5046 3596
rect 5050 3556 5054 3596
rect 5058 3556 5060 3596
rect 5072 3556 5074 3596
rect 5078 3556 5082 3596
rect 5086 3556 5088 3596
rect 5143 3576 5145 3596
rect 5149 3576 5151 3596
rect 5189 3556 5191 3596
rect 5195 3576 5199 3596
rect 5211 3576 5213 3596
rect 5217 3576 5223 3596
rect 5227 3576 5229 3596
rect 5241 3576 5243 3596
rect 5247 3576 5251 3596
rect 5255 3576 5257 3596
rect 5295 3576 5297 3596
rect 5301 3576 5305 3596
rect 5317 3576 5319 3596
rect 5323 3576 5329 3596
rect 5333 3576 5335 3596
rect 5347 3576 5351 3596
rect 5355 3576 5361 3596
rect 5365 3576 5367 3596
rect 5379 3576 5381 3596
rect 5195 3556 5208 3576
rect 5371 3556 5381 3576
rect 5385 3556 5387 3596
rect 5429 3556 5431 3596
rect 5435 3576 5439 3596
rect 5451 3576 5453 3596
rect 5457 3576 5463 3596
rect 5467 3576 5469 3596
rect 5481 3576 5483 3596
rect 5487 3576 5491 3596
rect 5495 3576 5497 3596
rect 5535 3576 5537 3596
rect 5541 3576 5545 3596
rect 5557 3576 5559 3596
rect 5563 3576 5569 3596
rect 5573 3576 5575 3596
rect 5587 3576 5591 3596
rect 5595 3576 5601 3596
rect 5605 3576 5607 3596
rect 5619 3576 5621 3596
rect 5435 3556 5448 3576
rect 5611 3556 5621 3576
rect 5625 3556 5627 3596
rect 5669 3556 5671 3596
rect 5675 3568 5677 3596
rect 5689 3568 5691 3596
rect 5675 3556 5691 3568
rect 5695 3556 5697 3596
rect 5709 3556 5711 3596
rect 5715 3556 5717 3596
rect 5769 3556 5771 3596
rect 5775 3568 5777 3596
rect 5789 3568 5791 3596
rect 5775 3556 5791 3568
rect 5795 3556 5797 3596
rect 5809 3556 5811 3596
rect 5815 3556 5817 3596
rect 5883 3576 5885 3596
rect 5889 3576 5891 3596
rect 5964 3556 5966 3596
rect 5970 3556 5974 3596
rect 5978 3556 5980 3596
rect 5992 3556 5994 3596
rect 5998 3556 6002 3596
rect 6006 3556 6008 3596
rect 6051 3556 6053 3596
rect 6057 3556 6063 3596
rect 6067 3556 6069 3596
rect 6143 3576 6145 3596
rect 6149 3576 6151 3596
rect 6209 3576 6211 3596
rect 6215 3576 6217 3596
rect 6229 3576 6231 3596
rect 6235 3576 6237 3596
rect 6249 3576 6251 3596
rect 6255 3576 6257 3596
rect 6383 3576 6385 3596
rect 6389 3576 6391 3596
rect 6429 3556 6431 3596
rect 6435 3576 6439 3596
rect 6451 3576 6453 3596
rect 6457 3576 6463 3596
rect 6467 3576 6469 3596
rect 6481 3576 6483 3596
rect 6487 3576 6491 3596
rect 6495 3576 6497 3596
rect 6535 3576 6537 3596
rect 6541 3576 6545 3596
rect 6557 3576 6559 3596
rect 6563 3576 6569 3596
rect 6573 3576 6575 3596
rect 6587 3576 6591 3596
rect 6595 3576 6601 3596
rect 6605 3576 6607 3596
rect 6619 3576 6621 3596
rect 6435 3556 6448 3576
rect 6611 3556 6621 3576
rect 6625 3556 6627 3596
rect 41 3144 43 3184
rect 47 3144 49 3184
rect 61 3144 65 3164
rect 69 3144 71 3164
rect 109 3144 111 3184
rect 115 3164 128 3184
rect 291 3164 301 3184
rect 115 3144 119 3164
rect 131 3144 133 3164
rect 137 3144 143 3164
rect 147 3144 149 3164
rect 161 3144 163 3164
rect 167 3144 171 3164
rect 175 3144 177 3164
rect 215 3144 217 3164
rect 221 3144 225 3164
rect 237 3144 239 3164
rect 243 3144 249 3164
rect 253 3144 255 3164
rect 267 3144 271 3164
rect 275 3144 281 3164
rect 285 3144 287 3164
rect 299 3144 301 3164
rect 305 3144 307 3184
rect 351 3144 353 3184
rect 357 3144 363 3184
rect 367 3144 369 3184
rect 450 3144 452 3164
rect 456 3144 460 3164
rect 472 3144 474 3184
rect 478 3144 482 3184
rect 486 3144 488 3184
rect 551 3144 553 3184
rect 557 3144 563 3184
rect 567 3144 569 3184
rect 609 3144 611 3164
rect 615 3144 617 3164
rect 670 3144 672 3204
rect 676 3144 680 3204
rect 684 3144 688 3204
rect 692 3202 706 3204
rect 692 3144 694 3202
rect 771 3144 773 3184
rect 777 3144 783 3184
rect 787 3144 789 3184
rect 863 3144 865 3184
rect 869 3144 871 3184
rect 883 3144 885 3184
rect 889 3172 905 3184
rect 889 3144 891 3172
rect 903 3144 905 3172
rect 909 3144 911 3184
rect 949 3144 951 3164
rect 955 3144 957 3164
rect 1009 3144 1011 3164
rect 1015 3144 1017 3164
rect 1029 3144 1031 3164
rect 1035 3144 1037 3164
rect 1089 3144 1091 3184
rect 1095 3172 1111 3184
rect 1095 3144 1097 3172
rect 1109 3144 1111 3172
rect 1115 3144 1117 3184
rect 1129 3144 1131 3184
rect 1135 3144 1137 3184
rect 1189 3144 1191 3184
rect 1195 3172 1211 3184
rect 1195 3144 1197 3172
rect 1209 3144 1211 3172
rect 1215 3144 1217 3184
rect 1229 3144 1231 3184
rect 1235 3144 1237 3184
rect 1291 3144 1293 3184
rect 1297 3144 1303 3184
rect 1307 3144 1309 3184
rect 1369 3144 1371 3184
rect 1375 3164 1388 3184
rect 1551 3164 1561 3184
rect 1375 3144 1379 3164
rect 1391 3144 1393 3164
rect 1397 3144 1403 3164
rect 1407 3144 1409 3164
rect 1421 3144 1423 3164
rect 1427 3144 1431 3164
rect 1435 3144 1437 3164
rect 1475 3144 1477 3164
rect 1481 3144 1485 3164
rect 1497 3144 1499 3164
rect 1503 3144 1509 3164
rect 1513 3144 1515 3164
rect 1527 3144 1531 3164
rect 1535 3144 1541 3164
rect 1545 3144 1547 3164
rect 1559 3144 1561 3164
rect 1565 3144 1567 3184
rect 1633 3144 1635 3184
rect 1639 3144 1641 3184
rect 1653 3144 1655 3184
rect 1659 3144 1665 3184
rect 1669 3144 1671 3184
rect 1834 3202 1848 3204
rect 1730 3144 1732 3164
rect 1736 3144 1740 3164
rect 1752 3144 1754 3184
rect 1758 3144 1762 3184
rect 1766 3144 1768 3184
rect 1846 3144 1848 3202
rect 1852 3144 1856 3204
rect 1860 3144 1864 3204
rect 1868 3144 1870 3204
rect 1912 3144 1914 3184
rect 1918 3144 1922 3184
rect 1926 3144 1928 3184
rect 1940 3144 1944 3164
rect 1948 3144 1950 3164
rect 2013 3144 2015 3184
rect 2019 3164 2029 3184
rect 2192 3164 2205 3184
rect 2019 3144 2021 3164
rect 2033 3144 2035 3164
rect 2039 3144 2045 3164
rect 2049 3144 2053 3164
rect 2065 3144 2067 3164
rect 2071 3144 2077 3164
rect 2081 3144 2083 3164
rect 2095 3144 2099 3164
rect 2103 3144 2105 3164
rect 2143 3144 2145 3164
rect 2149 3144 2153 3164
rect 2157 3144 2159 3164
rect 2171 3144 2173 3164
rect 2177 3144 2183 3164
rect 2187 3144 2189 3164
rect 2201 3144 2205 3164
rect 2209 3144 2211 3184
rect 2251 3144 2253 3184
rect 2257 3144 2263 3184
rect 2267 3144 2269 3184
rect 2329 3144 2331 3164
rect 2335 3144 2337 3164
rect 2349 3144 2351 3164
rect 2355 3144 2357 3164
rect 2423 3144 2425 3164
rect 2429 3144 2431 3164
rect 2443 3144 2445 3164
rect 2449 3144 2451 3164
rect 2503 3144 2505 3184
rect 2509 3144 2511 3184
rect 2523 3144 2525 3184
rect 2529 3172 2545 3184
rect 2529 3144 2531 3172
rect 2543 3144 2545 3172
rect 2549 3144 2551 3184
rect 2589 3144 2591 3164
rect 2595 3144 2597 3164
rect 2653 3144 2655 3184
rect 2659 3164 2669 3184
rect 2832 3164 2845 3184
rect 2659 3144 2661 3164
rect 2673 3144 2675 3164
rect 2679 3144 2685 3164
rect 2689 3144 2693 3164
rect 2705 3144 2707 3164
rect 2711 3144 2717 3164
rect 2721 3144 2723 3164
rect 2735 3144 2739 3164
rect 2743 3144 2745 3164
rect 2783 3144 2785 3164
rect 2789 3144 2793 3164
rect 2797 3144 2799 3164
rect 2811 3144 2813 3164
rect 2817 3144 2823 3164
rect 2827 3144 2829 3164
rect 2841 3144 2845 3164
rect 2849 3144 2851 3184
rect 2891 3144 2893 3184
rect 2897 3144 2903 3184
rect 2907 3144 2909 3184
rect 2991 3144 2993 3184
rect 2997 3144 3003 3184
rect 3007 3144 3009 3184
rect 3063 3144 3065 3184
rect 3069 3144 3071 3184
rect 3083 3144 3085 3184
rect 3089 3172 3105 3184
rect 3089 3144 3091 3172
rect 3103 3144 3105 3172
rect 3109 3144 3111 3184
rect 3171 3144 3173 3184
rect 3177 3144 3183 3184
rect 3187 3144 3189 3184
rect 3243 3144 3245 3164
rect 3249 3144 3251 3164
rect 3303 3144 3305 3184
rect 3309 3144 3311 3184
rect 3323 3144 3325 3184
rect 3329 3172 3345 3184
rect 3329 3144 3331 3172
rect 3343 3144 3345 3172
rect 3349 3144 3351 3184
rect 3389 3144 3391 3164
rect 3395 3144 3397 3164
rect 3463 3144 3465 3164
rect 3469 3144 3471 3164
rect 3483 3144 3485 3164
rect 3489 3144 3491 3164
rect 3550 3144 3552 3164
rect 3556 3144 3560 3164
rect 3572 3144 3574 3184
rect 3578 3144 3582 3184
rect 3586 3144 3588 3184
rect 3643 3144 3645 3164
rect 3649 3144 3651 3164
rect 3663 3144 3665 3164
rect 3669 3144 3671 3164
rect 3709 3144 3711 3184
rect 3715 3164 3728 3184
rect 3891 3164 3901 3184
rect 3715 3144 3719 3164
rect 3731 3144 3733 3164
rect 3737 3144 3743 3164
rect 3747 3144 3749 3164
rect 3761 3144 3763 3164
rect 3767 3144 3771 3164
rect 3775 3144 3777 3164
rect 3815 3144 3817 3164
rect 3821 3144 3825 3164
rect 3837 3144 3839 3164
rect 3843 3144 3849 3164
rect 3853 3144 3855 3164
rect 3867 3144 3871 3164
rect 3875 3144 3881 3164
rect 3885 3144 3887 3164
rect 3899 3144 3901 3164
rect 3905 3144 3907 3184
rect 3952 3144 3954 3184
rect 3958 3144 3962 3184
rect 3966 3144 3968 3184
rect 3980 3144 3982 3184
rect 3986 3144 3990 3184
rect 3994 3144 3996 3184
rect 4104 3144 4106 3184
rect 4110 3144 4114 3184
rect 4118 3144 4120 3184
rect 4132 3144 4134 3184
rect 4138 3144 4142 3184
rect 4146 3144 4148 3184
rect 4193 3144 4195 3184
rect 4199 3164 4209 3184
rect 4372 3164 4385 3184
rect 4199 3144 4201 3164
rect 4213 3144 4215 3164
rect 4219 3144 4225 3164
rect 4229 3144 4233 3164
rect 4245 3144 4247 3164
rect 4251 3144 4257 3164
rect 4261 3144 4263 3164
rect 4275 3144 4279 3164
rect 4283 3144 4285 3164
rect 4323 3144 4325 3164
rect 4329 3144 4333 3164
rect 4337 3144 4339 3164
rect 4351 3144 4353 3164
rect 4357 3144 4363 3164
rect 4367 3144 4369 3164
rect 4381 3144 4385 3164
rect 4389 3144 4391 3184
rect 4429 3144 4431 3164
rect 4435 3144 4437 3164
rect 4449 3144 4451 3164
rect 4455 3144 4457 3164
rect 4512 3144 4514 3184
rect 4518 3144 4522 3184
rect 4526 3144 4528 3184
rect 4540 3144 4542 3184
rect 4546 3144 4550 3184
rect 4554 3144 4556 3184
rect 4629 3144 4631 3164
rect 4635 3144 4637 3164
rect 4649 3144 4651 3164
rect 4655 3144 4657 3164
rect 4709 3144 4711 3164
rect 4715 3144 4717 3164
rect 4729 3144 4731 3164
rect 4735 3144 4737 3164
rect 4789 3144 4791 3164
rect 4795 3144 4797 3164
rect 4852 3144 4854 3184
rect 4858 3144 4862 3184
rect 4866 3144 4868 3184
rect 4880 3144 4882 3184
rect 4886 3144 4890 3184
rect 4894 3144 4896 3184
rect 4972 3144 4974 3184
rect 4978 3144 4982 3184
rect 4986 3144 4988 3184
rect 5000 3144 5004 3164
rect 5008 3144 5010 3164
rect 5069 3144 5071 3184
rect 5075 3164 5088 3184
rect 5251 3164 5261 3184
rect 5075 3144 5079 3164
rect 5091 3144 5093 3164
rect 5097 3144 5103 3164
rect 5107 3144 5109 3164
rect 5121 3144 5123 3164
rect 5127 3144 5131 3164
rect 5135 3144 5137 3164
rect 5175 3144 5177 3164
rect 5181 3144 5185 3164
rect 5197 3144 5199 3164
rect 5203 3144 5209 3164
rect 5213 3144 5215 3164
rect 5227 3144 5231 3164
rect 5235 3144 5241 3164
rect 5245 3144 5247 3164
rect 5259 3144 5261 3164
rect 5265 3144 5267 3184
rect 5379 3172 5391 3192
rect 5323 3144 5325 3164
rect 5329 3144 5331 3164
rect 5369 3152 5371 3172
rect 5375 3152 5377 3172
rect 5389 3152 5391 3172
rect 5395 3152 5401 3192
rect 5405 3184 5421 3192
rect 5405 3152 5407 3184
rect 5419 3152 5421 3184
rect 5425 3152 5431 3192
rect 5435 3152 5437 3192
rect 5503 3144 5505 3164
rect 5509 3144 5511 3164
rect 5553 3144 5555 3184
rect 5559 3164 5569 3184
rect 5732 3164 5745 3184
rect 5559 3144 5561 3164
rect 5573 3144 5575 3164
rect 5579 3144 5585 3164
rect 5589 3144 5593 3164
rect 5605 3144 5607 3164
rect 5611 3144 5617 3164
rect 5621 3144 5623 3164
rect 5635 3144 5639 3164
rect 5643 3144 5645 3164
rect 5683 3144 5685 3164
rect 5689 3144 5693 3164
rect 5697 3144 5699 3164
rect 5711 3144 5713 3164
rect 5717 3144 5723 3164
rect 5727 3144 5729 3164
rect 5741 3144 5745 3164
rect 5749 3144 5751 3184
rect 5803 3144 5805 3184
rect 5809 3144 5811 3184
rect 5823 3144 5825 3184
rect 5829 3172 5845 3184
rect 5829 3144 5831 3172
rect 5843 3144 5845 3172
rect 5849 3144 5851 3184
rect 5903 3144 5905 3164
rect 5909 3144 5911 3164
rect 5970 3144 5972 3164
rect 5976 3144 5980 3164
rect 5992 3144 5994 3184
rect 5998 3144 6002 3184
rect 6006 3144 6008 3184
rect 6049 3144 6051 3184
rect 6055 3172 6071 3184
rect 6055 3144 6057 3172
rect 6069 3144 6071 3172
rect 6075 3144 6077 3184
rect 6089 3144 6091 3184
rect 6095 3144 6097 3184
rect 6171 3144 6173 3184
rect 6177 3144 6183 3184
rect 6187 3144 6189 3184
rect 6250 3144 6252 3164
rect 6256 3144 6260 3164
rect 6272 3144 6274 3184
rect 6278 3144 6282 3184
rect 6286 3144 6288 3184
rect 6351 3144 6353 3184
rect 6357 3144 6363 3184
rect 6367 3144 6369 3184
rect 6409 3144 6411 3184
rect 6415 3172 6431 3184
rect 6415 3144 6417 3172
rect 6429 3144 6431 3172
rect 6435 3144 6437 3184
rect 6449 3144 6451 3184
rect 6455 3144 6457 3184
rect 6509 3144 6511 3184
rect 6515 3164 6528 3184
rect 6691 3164 6701 3184
rect 6515 3144 6519 3164
rect 6531 3144 6533 3164
rect 6537 3144 6543 3164
rect 6547 3144 6549 3164
rect 6561 3144 6563 3164
rect 6567 3144 6571 3164
rect 6575 3144 6577 3164
rect 6615 3144 6617 3164
rect 6621 3144 6625 3164
rect 6637 3144 6639 3164
rect 6643 3144 6649 3164
rect 6653 3144 6655 3164
rect 6667 3144 6671 3164
rect 6675 3144 6681 3164
rect 6685 3144 6687 3164
rect 6699 3144 6701 3164
rect 6705 3144 6707 3184
rect 29 3076 31 3116
rect 35 3076 37 3116
rect 49 3076 51 3116
rect 55 3076 57 3116
rect 69 3076 71 3116
rect 75 3076 77 3116
rect 89 3076 91 3116
rect 95 3076 97 3116
rect 109 3076 111 3116
rect 115 3076 117 3116
rect 129 3076 131 3116
rect 135 3076 137 3116
rect 149 3076 151 3116
rect 155 3076 157 3116
rect 169 3076 171 3116
rect 175 3076 177 3116
rect 241 3076 243 3116
rect 247 3076 249 3116
rect 261 3096 265 3116
rect 269 3096 271 3116
rect 313 3076 315 3116
rect 319 3096 321 3116
rect 333 3096 335 3116
rect 339 3096 345 3116
rect 349 3096 353 3116
rect 365 3096 367 3116
rect 371 3096 377 3116
rect 381 3096 383 3116
rect 395 3096 399 3116
rect 403 3096 405 3116
rect 443 3096 445 3116
rect 449 3096 453 3116
rect 457 3096 459 3116
rect 471 3096 473 3116
rect 477 3096 483 3116
rect 487 3096 489 3116
rect 501 3096 505 3116
rect 319 3076 329 3096
rect 492 3076 505 3096
rect 509 3076 511 3116
rect 571 3076 573 3116
rect 577 3076 583 3116
rect 587 3076 589 3116
rect 631 3076 633 3116
rect 637 3076 643 3116
rect 647 3076 649 3116
rect 723 3076 725 3116
rect 729 3076 731 3116
rect 743 3076 745 3116
rect 749 3088 751 3116
rect 763 3088 765 3116
rect 749 3076 765 3088
rect 769 3076 771 3116
rect 831 3076 833 3116
rect 837 3076 843 3116
rect 847 3076 849 3116
rect 911 3076 913 3116
rect 917 3076 923 3116
rect 927 3076 929 3116
rect 972 3076 974 3116
rect 978 3076 982 3116
rect 986 3076 988 3116
rect 1000 3096 1004 3116
rect 1008 3096 1010 3116
rect 1069 3076 1071 3116
rect 1075 3096 1079 3116
rect 1091 3096 1093 3116
rect 1097 3096 1103 3116
rect 1107 3096 1109 3116
rect 1121 3096 1123 3116
rect 1127 3096 1131 3116
rect 1135 3096 1137 3116
rect 1175 3096 1177 3116
rect 1181 3096 1185 3116
rect 1197 3096 1199 3116
rect 1203 3096 1209 3116
rect 1213 3096 1215 3116
rect 1227 3096 1231 3116
rect 1235 3096 1241 3116
rect 1245 3096 1247 3116
rect 1259 3096 1261 3116
rect 1075 3076 1088 3096
rect 1251 3076 1261 3096
rect 1265 3076 1267 3116
rect 1331 3076 1333 3116
rect 1337 3076 1343 3116
rect 1347 3076 1349 3116
rect 1389 3076 1391 3116
rect 1395 3096 1399 3116
rect 1411 3096 1413 3116
rect 1417 3096 1423 3116
rect 1427 3096 1429 3116
rect 1441 3096 1443 3116
rect 1447 3096 1451 3116
rect 1455 3096 1457 3116
rect 1495 3096 1497 3116
rect 1501 3096 1505 3116
rect 1517 3096 1519 3116
rect 1523 3096 1529 3116
rect 1533 3096 1535 3116
rect 1547 3096 1551 3116
rect 1555 3096 1561 3116
rect 1565 3096 1567 3116
rect 1579 3096 1581 3116
rect 1395 3076 1408 3096
rect 1571 3076 1581 3096
rect 1585 3076 1587 3116
rect 1643 3096 1645 3116
rect 1649 3096 1651 3116
rect 1703 3076 1705 3116
rect 1709 3076 1711 3116
rect 1723 3076 1725 3116
rect 1729 3088 1731 3116
rect 1743 3088 1745 3116
rect 1729 3076 1745 3088
rect 1749 3076 1751 3116
rect 1803 3096 1805 3116
rect 1809 3096 1811 3116
rect 1823 3096 1825 3116
rect 1829 3096 1831 3116
rect 1893 3076 1895 3116
rect 1899 3076 1901 3116
rect 1913 3076 1915 3116
rect 1919 3076 1925 3116
rect 1929 3076 1931 3116
rect 1969 3076 1971 3116
rect 1975 3088 1977 3116
rect 1989 3088 1991 3116
rect 1975 3076 1991 3088
rect 1995 3076 1997 3116
rect 2009 3076 2011 3116
rect 2015 3076 2017 3116
rect 2090 3096 2092 3116
rect 2096 3096 2100 3116
rect 2112 3076 2114 3116
rect 2118 3076 2122 3116
rect 2126 3076 2128 3116
rect 2171 3076 2173 3116
rect 2177 3076 2183 3116
rect 2187 3076 2189 3116
rect 2263 3096 2265 3116
rect 2269 3096 2271 3116
rect 2309 3076 2311 3116
rect 2315 3076 2321 3116
rect 2325 3076 2327 3116
rect 2339 3076 2341 3116
rect 2345 3076 2347 3116
rect 2413 3076 2415 3116
rect 2419 3096 2421 3116
rect 2433 3096 2435 3116
rect 2439 3096 2445 3116
rect 2449 3096 2453 3116
rect 2465 3096 2467 3116
rect 2471 3096 2477 3116
rect 2481 3096 2483 3116
rect 2495 3096 2499 3116
rect 2503 3096 2505 3116
rect 2543 3096 2545 3116
rect 2549 3096 2553 3116
rect 2557 3096 2559 3116
rect 2571 3096 2573 3116
rect 2577 3096 2583 3116
rect 2587 3096 2589 3116
rect 2601 3096 2605 3116
rect 2419 3076 2429 3096
rect 2592 3076 2605 3096
rect 2609 3076 2611 3116
rect 2649 3096 2651 3116
rect 2655 3096 2657 3116
rect 2709 3096 2711 3116
rect 2715 3096 2717 3116
rect 2729 3096 2731 3116
rect 2735 3096 2737 3116
rect 2803 3096 2805 3116
rect 2809 3096 2811 3116
rect 2863 3076 2865 3116
rect 2869 3076 2871 3116
rect 2883 3076 2885 3116
rect 2889 3088 2891 3116
rect 2903 3088 2905 3116
rect 2889 3076 2905 3088
rect 2909 3076 2911 3116
rect 2949 3076 2951 3116
rect 2955 3076 2957 3116
rect 3046 3058 3048 3116
rect 3034 3056 3048 3058
rect 3052 3056 3056 3116
rect 3060 3056 3064 3116
rect 3068 3056 3070 3116
rect 3131 3076 3133 3116
rect 3137 3076 3143 3116
rect 3147 3076 3149 3116
rect 3203 3076 3205 3116
rect 3209 3076 3211 3116
rect 3223 3076 3225 3116
rect 3229 3088 3231 3116
rect 3243 3088 3245 3116
rect 3229 3076 3245 3088
rect 3249 3076 3251 3116
rect 3291 3076 3293 3116
rect 3297 3076 3303 3116
rect 3307 3076 3309 3116
rect 3371 3076 3373 3116
rect 3377 3076 3383 3116
rect 3387 3076 3389 3116
rect 3449 3076 3451 3116
rect 3455 3088 3457 3116
rect 3469 3088 3471 3116
rect 3455 3076 3471 3088
rect 3475 3076 3477 3116
rect 3489 3076 3491 3116
rect 3495 3076 3497 3116
rect 3549 3076 3551 3116
rect 3555 3076 3561 3116
rect 3565 3076 3567 3116
rect 3579 3076 3581 3116
rect 3585 3076 3587 3116
rect 3684 3076 3686 3116
rect 3690 3076 3694 3116
rect 3698 3076 3700 3116
rect 3712 3076 3714 3116
rect 3718 3076 3722 3116
rect 3726 3076 3728 3116
rect 3783 3076 3785 3116
rect 3789 3076 3791 3116
rect 3803 3076 3805 3116
rect 3809 3076 3811 3116
rect 3853 3076 3855 3116
rect 3859 3096 3861 3116
rect 3873 3096 3875 3116
rect 3879 3096 3885 3116
rect 3889 3096 3893 3116
rect 3905 3096 3907 3116
rect 3911 3096 3917 3116
rect 3921 3096 3923 3116
rect 3935 3096 3939 3116
rect 3943 3096 3945 3116
rect 3983 3096 3985 3116
rect 3989 3096 3993 3116
rect 3997 3096 3999 3116
rect 4011 3096 4013 3116
rect 4017 3096 4023 3116
rect 4027 3096 4029 3116
rect 4041 3096 4045 3116
rect 3859 3076 3869 3096
rect 4032 3076 4045 3096
rect 4049 3076 4051 3116
rect 4089 3076 4091 3116
rect 4095 3088 4097 3116
rect 4109 3088 4111 3116
rect 4095 3076 4111 3088
rect 4115 3076 4117 3116
rect 4129 3076 4131 3116
rect 4135 3076 4137 3116
rect 4226 3058 4228 3116
rect 4214 3056 4228 3058
rect 4232 3056 4236 3116
rect 4240 3056 4244 3116
rect 4248 3056 4250 3116
rect 4293 3076 4295 3116
rect 4299 3096 4301 3116
rect 4313 3096 4315 3116
rect 4319 3096 4325 3116
rect 4329 3096 4333 3116
rect 4345 3096 4347 3116
rect 4351 3096 4357 3116
rect 4361 3096 4363 3116
rect 4375 3096 4379 3116
rect 4383 3096 4385 3116
rect 4423 3096 4425 3116
rect 4429 3096 4433 3116
rect 4437 3096 4439 3116
rect 4451 3096 4453 3116
rect 4457 3096 4463 3116
rect 4467 3096 4469 3116
rect 4481 3096 4485 3116
rect 4299 3076 4309 3096
rect 4472 3076 4485 3096
rect 4489 3076 4491 3116
rect 4543 3076 4545 3116
rect 4549 3104 4565 3116
rect 4549 3076 4551 3104
rect 4563 3076 4565 3104
rect 4569 3076 4571 3116
rect 4583 3076 4585 3116
rect 4589 3086 4591 3116
rect 4603 3086 4605 3116
rect 4589 3076 4605 3086
rect 4609 3076 4611 3116
rect 4663 3096 4665 3116
rect 4669 3096 4671 3116
rect 4723 3068 4725 3108
rect 4729 3068 4735 3108
rect 4739 3076 4741 3108
rect 4753 3076 4755 3108
rect 4739 3068 4755 3076
rect 4759 3068 4765 3108
rect 4769 3088 4771 3108
rect 4783 3088 4785 3108
rect 4789 3088 4791 3108
rect 4769 3068 4781 3088
rect 4832 3076 4834 3116
rect 4838 3076 4842 3116
rect 4846 3076 4848 3116
rect 4860 3076 4862 3116
rect 4866 3076 4870 3116
rect 4874 3076 4876 3116
rect 4963 3096 4965 3116
rect 4969 3096 4971 3116
rect 5012 3076 5014 3116
rect 5018 3076 5022 3116
rect 5026 3076 5028 3116
rect 5040 3076 5042 3116
rect 5046 3076 5050 3116
rect 5054 3076 5056 3116
rect 5129 3096 5131 3116
rect 5135 3096 5137 3116
rect 5189 3096 5191 3116
rect 5195 3096 5197 3116
rect 5209 3096 5211 3116
rect 5215 3096 5217 3116
rect 5273 3076 5275 3116
rect 5279 3096 5281 3116
rect 5293 3096 5295 3116
rect 5299 3096 5305 3116
rect 5309 3096 5313 3116
rect 5325 3096 5327 3116
rect 5331 3096 5337 3116
rect 5341 3096 5343 3116
rect 5355 3096 5359 3116
rect 5363 3096 5365 3116
rect 5403 3096 5405 3116
rect 5409 3096 5413 3116
rect 5417 3096 5419 3116
rect 5431 3096 5433 3116
rect 5437 3096 5443 3116
rect 5447 3096 5449 3116
rect 5461 3096 5465 3116
rect 5279 3076 5289 3096
rect 5452 3076 5465 3096
rect 5469 3076 5471 3116
rect 5523 3096 5525 3116
rect 5529 3096 5531 3116
rect 5543 3096 5545 3116
rect 5549 3096 5551 3116
rect 5589 3076 5591 3116
rect 5595 3088 5597 3116
rect 5609 3088 5611 3116
rect 5595 3076 5611 3088
rect 5615 3076 5617 3116
rect 5629 3076 5631 3116
rect 5635 3076 5637 3116
rect 5726 3058 5728 3116
rect 5714 3056 5728 3058
rect 5732 3056 5736 3116
rect 5740 3056 5744 3116
rect 5748 3056 5750 3116
rect 5803 3076 5805 3116
rect 5809 3104 5825 3116
rect 5809 3076 5811 3104
rect 5823 3076 5825 3104
rect 5829 3076 5831 3116
rect 5843 3076 5845 3116
rect 5849 3086 5851 3116
rect 5863 3086 5865 3116
rect 5849 3076 5865 3086
rect 5869 3076 5871 3116
rect 5909 3096 5911 3116
rect 5915 3096 5917 3116
rect 5969 3088 5971 3108
rect 5975 3088 5977 3108
rect 5989 3088 5991 3108
rect 5979 3068 5991 3088
rect 5995 3068 6001 3108
rect 6005 3076 6007 3108
rect 6019 3076 6021 3108
rect 6005 3068 6021 3076
rect 6025 3068 6031 3108
rect 6035 3068 6037 3108
rect 6110 3096 6112 3116
rect 6116 3096 6120 3116
rect 6132 3076 6134 3116
rect 6138 3076 6142 3116
rect 6146 3076 6148 3116
rect 6203 3096 6205 3116
rect 6209 3096 6211 3116
rect 6223 3096 6225 3116
rect 6229 3096 6231 3116
rect 6269 3096 6271 3116
rect 6275 3096 6277 3116
rect 6364 3076 6366 3116
rect 6370 3076 6374 3116
rect 6378 3076 6380 3116
rect 6392 3076 6394 3116
rect 6398 3076 6402 3116
rect 6406 3076 6408 3116
rect 6463 3096 6465 3116
rect 6469 3096 6471 3116
rect 6509 3096 6511 3116
rect 6515 3096 6517 3116
rect 6569 3076 6571 3116
rect 6575 3088 6577 3116
rect 6589 3088 6591 3116
rect 6575 3076 6591 3088
rect 6595 3076 6597 3116
rect 6609 3076 6611 3116
rect 6615 3076 6617 3116
rect 29 2664 31 2684
rect 35 2664 37 2684
rect 103 2664 105 2684
rect 109 2664 111 2684
rect 123 2664 125 2684
rect 129 2664 131 2684
rect 173 2664 175 2704
rect 179 2684 189 2704
rect 352 2684 365 2704
rect 179 2664 181 2684
rect 193 2664 195 2684
rect 199 2664 205 2684
rect 209 2664 213 2684
rect 225 2664 227 2684
rect 231 2664 237 2684
rect 241 2664 243 2684
rect 255 2664 259 2684
rect 263 2664 265 2684
rect 303 2664 305 2684
rect 309 2664 313 2684
rect 317 2664 319 2684
rect 331 2664 333 2684
rect 337 2664 343 2684
rect 347 2664 349 2684
rect 361 2664 365 2684
rect 369 2664 371 2704
rect 409 2664 411 2684
rect 415 2664 417 2684
rect 483 2664 485 2684
rect 489 2664 491 2684
rect 503 2664 505 2684
rect 509 2664 511 2684
rect 553 2664 555 2704
rect 559 2684 569 2704
rect 732 2684 745 2704
rect 559 2664 561 2684
rect 573 2664 575 2684
rect 579 2664 585 2684
rect 589 2664 593 2684
rect 605 2664 607 2684
rect 611 2664 617 2684
rect 621 2664 623 2684
rect 635 2664 639 2684
rect 643 2664 645 2684
rect 683 2664 685 2684
rect 689 2664 693 2684
rect 697 2664 699 2684
rect 711 2664 713 2684
rect 717 2664 723 2684
rect 727 2664 729 2684
rect 741 2664 745 2684
rect 749 2664 751 2704
rect 801 2664 803 2704
rect 807 2664 809 2704
rect 821 2664 825 2684
rect 829 2664 831 2684
rect 869 2664 871 2704
rect 875 2664 877 2704
rect 889 2664 891 2704
rect 895 2664 897 2704
rect 951 2664 953 2704
rect 957 2664 963 2704
rect 967 2664 969 2704
rect 1031 2664 1033 2704
rect 1037 2664 1043 2704
rect 1047 2664 1049 2704
rect 1109 2664 1111 2684
rect 1115 2664 1117 2684
rect 1172 2664 1174 2704
rect 1178 2664 1182 2704
rect 1186 2664 1188 2704
rect 1200 2664 1202 2704
rect 1206 2664 1210 2704
rect 1214 2664 1216 2704
rect 1310 2664 1312 2684
rect 1316 2664 1320 2684
rect 1332 2664 1334 2704
rect 1338 2664 1342 2704
rect 1346 2664 1348 2704
rect 1403 2664 1405 2684
rect 1409 2664 1411 2684
rect 1463 2664 1465 2704
rect 1469 2664 1471 2704
rect 1483 2664 1485 2704
rect 1489 2692 1505 2704
rect 1489 2664 1491 2692
rect 1503 2664 1505 2692
rect 1509 2664 1511 2704
rect 1549 2664 1551 2684
rect 1555 2664 1557 2684
rect 1569 2664 1571 2684
rect 1575 2664 1577 2684
rect 1631 2664 1633 2704
rect 1637 2664 1643 2704
rect 1647 2664 1649 2704
rect 1709 2664 1711 2684
rect 1715 2664 1717 2684
rect 1729 2664 1731 2684
rect 1735 2664 1737 2684
rect 1803 2664 1805 2704
rect 1809 2664 1811 2704
rect 1823 2664 1825 2704
rect 1829 2692 1845 2704
rect 1829 2664 1831 2692
rect 1843 2664 1845 2692
rect 1849 2664 1851 2704
rect 1919 2684 1931 2704
rect 1889 2664 1891 2684
rect 1895 2664 1897 2684
rect 1909 2664 1911 2684
rect 1915 2664 1917 2684
rect 1929 2664 1931 2684
rect 1935 2664 1937 2704
rect 1989 2664 1991 2704
rect 1995 2692 2011 2704
rect 1995 2664 1997 2692
rect 2009 2664 2011 2692
rect 2015 2664 2017 2704
rect 2029 2664 2031 2704
rect 2035 2664 2037 2704
rect 2110 2664 2112 2684
rect 2116 2664 2120 2684
rect 2132 2664 2134 2704
rect 2138 2664 2142 2704
rect 2146 2664 2148 2704
rect 2193 2664 2195 2704
rect 2199 2684 2209 2704
rect 2372 2684 2385 2704
rect 2199 2664 2201 2684
rect 2213 2664 2215 2684
rect 2219 2664 2225 2684
rect 2229 2664 2233 2684
rect 2245 2664 2247 2684
rect 2251 2664 2257 2684
rect 2261 2664 2263 2684
rect 2275 2664 2279 2684
rect 2283 2664 2285 2684
rect 2323 2664 2325 2684
rect 2329 2664 2333 2684
rect 2337 2664 2339 2684
rect 2351 2664 2353 2684
rect 2357 2664 2363 2684
rect 2367 2664 2369 2684
rect 2381 2664 2385 2684
rect 2389 2664 2391 2704
rect 2431 2664 2433 2704
rect 2437 2664 2443 2704
rect 2447 2664 2449 2704
rect 2509 2664 2511 2684
rect 2515 2664 2517 2684
rect 2583 2664 2585 2684
rect 2589 2664 2591 2684
rect 2633 2664 2635 2704
rect 2639 2684 2649 2704
rect 2812 2684 2825 2704
rect 2639 2664 2641 2684
rect 2653 2664 2655 2684
rect 2659 2664 2665 2684
rect 2669 2664 2673 2684
rect 2685 2664 2687 2684
rect 2691 2664 2697 2684
rect 2701 2664 2703 2684
rect 2715 2664 2719 2684
rect 2723 2664 2725 2684
rect 2763 2664 2765 2684
rect 2769 2664 2773 2684
rect 2777 2664 2779 2684
rect 2791 2664 2793 2684
rect 2797 2664 2803 2684
rect 2807 2664 2809 2684
rect 2821 2664 2825 2684
rect 2829 2664 2831 2704
rect 2869 2664 2871 2704
rect 2875 2692 2891 2704
rect 2875 2664 2877 2692
rect 2889 2664 2891 2692
rect 2895 2664 2897 2704
rect 2909 2664 2911 2704
rect 2915 2664 2917 2704
rect 2990 2664 2992 2684
rect 2996 2664 3000 2684
rect 3012 2664 3014 2704
rect 3018 2664 3022 2704
rect 3026 2664 3028 2704
rect 3069 2664 3071 2704
rect 3075 2684 3088 2704
rect 3251 2684 3261 2704
rect 3075 2664 3079 2684
rect 3091 2664 3093 2684
rect 3097 2664 3103 2684
rect 3107 2664 3109 2684
rect 3121 2664 3123 2684
rect 3127 2664 3131 2684
rect 3135 2664 3137 2684
rect 3175 2664 3177 2684
rect 3181 2664 3185 2684
rect 3197 2664 3199 2684
rect 3203 2664 3209 2684
rect 3213 2664 3215 2684
rect 3227 2664 3231 2684
rect 3235 2664 3241 2684
rect 3245 2664 3247 2684
rect 3259 2664 3261 2684
rect 3265 2664 3267 2704
rect 3309 2664 3311 2684
rect 3315 2664 3317 2684
rect 3369 2664 3371 2704
rect 3375 2694 3391 2704
rect 3375 2664 3377 2694
rect 3389 2664 3391 2694
rect 3395 2664 3397 2704
rect 3409 2664 3411 2704
rect 3415 2676 3417 2704
rect 3429 2676 3431 2704
rect 3415 2664 3431 2676
rect 3435 2664 3437 2704
rect 3489 2664 3491 2704
rect 3495 2692 3511 2704
rect 3495 2664 3497 2692
rect 3509 2664 3511 2692
rect 3515 2664 3517 2704
rect 3529 2664 3531 2704
rect 3535 2664 3537 2704
rect 3603 2664 3605 2704
rect 3609 2676 3611 2704
rect 3623 2676 3625 2704
rect 3609 2664 3625 2676
rect 3629 2664 3631 2704
rect 3643 2664 3645 2704
rect 3649 2694 3665 2704
rect 3649 2664 3651 2694
rect 3663 2664 3665 2694
rect 3669 2664 3671 2704
rect 3709 2664 3711 2704
rect 3715 2692 3731 2704
rect 3715 2664 3717 2692
rect 3729 2664 3731 2692
rect 3735 2664 3737 2704
rect 3749 2664 3751 2704
rect 3755 2664 3757 2704
rect 3823 2664 3825 2704
rect 3829 2676 3831 2704
rect 3843 2676 3845 2704
rect 3829 2664 3845 2676
rect 3849 2664 3851 2704
rect 3863 2664 3865 2704
rect 3869 2694 3885 2704
rect 3869 2664 3871 2694
rect 3883 2664 3885 2694
rect 3889 2664 3891 2704
rect 4374 2722 4388 2724
rect 3943 2664 3945 2684
rect 3949 2664 3951 2684
rect 3989 2664 3991 2684
rect 3995 2664 3997 2684
rect 4009 2664 4011 2684
rect 4015 2664 4017 2684
rect 4069 2664 4071 2684
rect 4075 2664 4077 2684
rect 4089 2664 4091 2684
rect 4095 2664 4097 2684
rect 4170 2664 4172 2684
rect 4176 2664 4180 2684
rect 4192 2664 4194 2704
rect 4198 2664 4202 2704
rect 4206 2664 4208 2704
rect 4249 2664 4251 2704
rect 4255 2692 4271 2704
rect 4255 2664 4257 2692
rect 4269 2664 4271 2692
rect 4275 2664 4277 2704
rect 4289 2664 4291 2704
rect 4295 2664 4297 2704
rect 4386 2664 4388 2722
rect 4392 2664 4396 2724
rect 4400 2664 4404 2724
rect 4408 2664 4410 2724
rect 4453 2664 4455 2704
rect 4459 2684 4469 2704
rect 4632 2684 4645 2704
rect 4459 2664 4461 2684
rect 4473 2664 4475 2684
rect 4479 2664 4485 2684
rect 4489 2664 4493 2684
rect 4505 2664 4507 2684
rect 4511 2664 4517 2684
rect 4521 2664 4523 2684
rect 4535 2664 4539 2684
rect 4543 2664 4545 2684
rect 4583 2664 4585 2684
rect 4589 2664 4593 2684
rect 4597 2664 4599 2684
rect 4611 2664 4613 2684
rect 4617 2664 4623 2684
rect 4627 2664 4629 2684
rect 4641 2664 4645 2684
rect 4649 2664 4651 2704
rect 4689 2664 4691 2684
rect 4695 2664 4697 2684
rect 4749 2664 4751 2684
rect 4755 2664 4757 2684
rect 4769 2664 4771 2684
rect 4775 2664 4777 2684
rect 4829 2664 4831 2704
rect 4835 2692 4851 2704
rect 4835 2664 4837 2692
rect 4849 2664 4851 2692
rect 4855 2664 4857 2704
rect 4869 2664 4871 2704
rect 4875 2664 4877 2704
rect 4943 2664 4945 2684
rect 4949 2664 4951 2684
rect 4963 2664 4965 2684
rect 4969 2664 4971 2684
rect 5023 2664 5025 2704
rect 5029 2676 5031 2704
rect 5043 2676 5045 2704
rect 5029 2664 5045 2676
rect 5049 2664 5051 2704
rect 5063 2664 5065 2704
rect 5069 2694 5085 2704
rect 5069 2664 5071 2694
rect 5083 2664 5085 2694
rect 5089 2664 5091 2704
rect 5132 2664 5134 2704
rect 5138 2664 5142 2704
rect 5146 2664 5148 2704
rect 5160 2664 5164 2684
rect 5168 2664 5170 2684
rect 5229 2664 5231 2684
rect 5235 2664 5239 2684
rect 5251 2664 5253 2704
rect 5257 2664 5259 2704
rect 5309 2664 5311 2704
rect 5315 2692 5331 2704
rect 5315 2664 5317 2692
rect 5329 2664 5331 2692
rect 5335 2664 5337 2704
rect 5349 2664 5351 2704
rect 5355 2664 5357 2704
rect 5423 2664 5425 2704
rect 5429 2676 5431 2704
rect 5443 2676 5445 2704
rect 5429 2664 5445 2676
rect 5449 2664 5451 2704
rect 5463 2664 5465 2704
rect 5469 2694 5485 2704
rect 5469 2664 5471 2694
rect 5483 2664 5485 2694
rect 5489 2664 5491 2704
rect 5543 2664 5545 2684
rect 5549 2664 5551 2684
rect 5593 2664 5595 2704
rect 5599 2684 5609 2704
rect 5772 2684 5785 2704
rect 5599 2664 5601 2684
rect 5613 2664 5615 2684
rect 5619 2664 5625 2684
rect 5629 2664 5633 2684
rect 5645 2664 5647 2684
rect 5651 2664 5657 2684
rect 5661 2664 5663 2684
rect 5675 2664 5679 2684
rect 5683 2664 5685 2684
rect 5723 2664 5725 2684
rect 5729 2664 5733 2684
rect 5737 2664 5739 2684
rect 5751 2664 5753 2684
rect 5757 2664 5763 2684
rect 5767 2664 5769 2684
rect 5781 2664 5785 2684
rect 5789 2664 5791 2704
rect 5839 2692 5851 2712
rect 5829 2672 5831 2692
rect 5835 2672 5837 2692
rect 5849 2672 5851 2692
rect 5855 2672 5861 2712
rect 5865 2704 5881 2712
rect 5865 2672 5867 2704
rect 5879 2672 5881 2704
rect 5885 2672 5891 2712
rect 5895 2672 5897 2712
rect 5959 2692 5971 2712
rect 5949 2672 5951 2692
rect 5955 2672 5957 2692
rect 5969 2672 5971 2692
rect 5975 2672 5981 2712
rect 5985 2704 6001 2712
rect 5985 2672 5987 2704
rect 5999 2672 6001 2704
rect 6005 2672 6011 2712
rect 6015 2672 6017 2712
rect 6079 2692 6091 2712
rect 6069 2672 6071 2692
rect 6075 2672 6077 2692
rect 6089 2672 6091 2692
rect 6095 2672 6101 2712
rect 6105 2704 6121 2712
rect 6105 2672 6107 2704
rect 6119 2672 6121 2704
rect 6125 2672 6131 2712
rect 6135 2672 6137 2712
rect 6213 2664 6215 2704
rect 6219 2664 6221 2704
rect 6233 2664 6235 2704
rect 6239 2664 6245 2704
rect 6249 2664 6251 2704
rect 6303 2664 6305 2704
rect 6309 2664 6311 2704
rect 6323 2664 6325 2704
rect 6329 2664 6331 2704
rect 6369 2664 6371 2704
rect 6375 2664 6381 2704
rect 6385 2664 6387 2704
rect 6399 2664 6401 2704
rect 6405 2664 6407 2704
rect 6469 2664 6471 2704
rect 6475 2684 6488 2704
rect 6651 2684 6661 2704
rect 6475 2664 6479 2684
rect 6491 2664 6493 2684
rect 6497 2664 6503 2684
rect 6507 2664 6509 2684
rect 6521 2664 6523 2684
rect 6527 2664 6531 2684
rect 6535 2664 6537 2684
rect 6575 2664 6577 2684
rect 6581 2664 6585 2684
rect 6597 2664 6599 2684
rect 6603 2664 6609 2684
rect 6613 2664 6615 2684
rect 6627 2664 6631 2684
rect 6635 2664 6641 2684
rect 6645 2664 6647 2684
rect 6659 2664 6661 2684
rect 6665 2664 6667 2704
rect 29 2596 31 2636
rect 35 2616 39 2636
rect 51 2616 53 2636
rect 57 2616 63 2636
rect 67 2616 69 2636
rect 81 2616 83 2636
rect 87 2616 91 2636
rect 95 2616 97 2636
rect 135 2616 137 2636
rect 141 2616 145 2636
rect 157 2616 159 2636
rect 163 2616 169 2636
rect 173 2616 175 2636
rect 187 2616 191 2636
rect 195 2616 201 2636
rect 205 2616 207 2636
rect 219 2616 221 2636
rect 35 2596 48 2616
rect 211 2596 221 2616
rect 225 2596 227 2636
rect 281 2596 283 2636
rect 287 2596 289 2636
rect 301 2616 305 2636
rect 309 2616 311 2636
rect 349 2596 351 2636
rect 355 2616 359 2636
rect 371 2616 373 2636
rect 377 2616 383 2636
rect 387 2616 389 2636
rect 401 2616 403 2636
rect 407 2616 411 2636
rect 415 2616 417 2636
rect 455 2616 457 2636
rect 461 2616 465 2636
rect 477 2616 479 2636
rect 483 2616 489 2636
rect 493 2616 495 2636
rect 507 2616 511 2636
rect 515 2616 521 2636
rect 525 2616 527 2636
rect 539 2616 541 2636
rect 355 2596 368 2616
rect 531 2596 541 2616
rect 545 2596 547 2636
rect 610 2616 612 2636
rect 616 2616 620 2636
rect 632 2596 634 2636
rect 638 2596 642 2636
rect 646 2596 648 2636
rect 691 2596 693 2636
rect 697 2596 703 2636
rect 707 2596 709 2636
rect 791 2596 793 2636
rect 797 2596 803 2636
rect 807 2596 809 2636
rect 863 2596 865 2636
rect 869 2596 871 2636
rect 883 2596 885 2636
rect 889 2596 891 2636
rect 903 2596 905 2636
rect 909 2596 911 2636
rect 923 2596 925 2636
rect 929 2596 931 2636
rect 943 2596 945 2636
rect 949 2596 951 2636
rect 963 2596 965 2636
rect 969 2596 971 2636
rect 983 2596 985 2636
rect 989 2596 991 2636
rect 1003 2596 1005 2636
rect 1009 2596 1011 2636
rect 1049 2596 1051 2636
rect 1055 2616 1059 2636
rect 1071 2616 1073 2636
rect 1077 2616 1083 2636
rect 1087 2616 1089 2636
rect 1101 2616 1103 2636
rect 1107 2616 1111 2636
rect 1115 2616 1117 2636
rect 1155 2616 1157 2636
rect 1161 2616 1165 2636
rect 1177 2616 1179 2636
rect 1183 2616 1189 2636
rect 1193 2616 1195 2636
rect 1207 2616 1211 2636
rect 1215 2616 1221 2636
rect 1225 2616 1227 2636
rect 1239 2616 1241 2636
rect 1055 2596 1068 2616
rect 1231 2596 1241 2616
rect 1245 2596 1247 2636
rect 1311 2596 1313 2636
rect 1317 2596 1323 2636
rect 1327 2596 1329 2636
rect 1369 2616 1371 2636
rect 1375 2616 1377 2636
rect 1389 2616 1391 2636
rect 1395 2616 1397 2636
rect 1449 2616 1451 2636
rect 1455 2616 1457 2636
rect 1523 2596 1525 2636
rect 1529 2596 1531 2636
rect 1543 2596 1545 2636
rect 1549 2608 1551 2636
rect 1563 2608 1565 2636
rect 1549 2596 1565 2608
rect 1569 2596 1571 2636
rect 1613 2596 1615 2636
rect 1619 2616 1621 2636
rect 1633 2616 1635 2636
rect 1639 2616 1645 2636
rect 1649 2616 1653 2636
rect 1665 2616 1667 2636
rect 1671 2616 1677 2636
rect 1681 2616 1683 2636
rect 1695 2616 1699 2636
rect 1703 2616 1705 2636
rect 1743 2616 1745 2636
rect 1749 2616 1753 2636
rect 1757 2616 1759 2636
rect 1771 2616 1773 2636
rect 1777 2616 1783 2636
rect 1787 2616 1789 2636
rect 1801 2616 1805 2636
rect 1619 2596 1629 2616
rect 1792 2596 1805 2616
rect 1809 2596 1811 2636
rect 1849 2616 1851 2636
rect 1855 2616 1857 2636
rect 1909 2616 1911 2636
rect 1915 2616 1917 2636
rect 1969 2596 1971 2636
rect 1975 2606 1977 2636
rect 1989 2606 1991 2636
rect 1975 2596 1991 2606
rect 1995 2596 1997 2636
rect 2009 2596 2011 2636
rect 2015 2624 2031 2636
rect 2015 2596 2017 2624
rect 2029 2596 2031 2624
rect 2035 2596 2037 2636
rect 2089 2616 2091 2636
rect 2095 2616 2097 2636
rect 2109 2616 2111 2636
rect 2115 2616 2117 2636
rect 2169 2608 2171 2628
rect 2175 2608 2177 2628
rect 2189 2608 2191 2628
rect 2179 2588 2191 2608
rect 2195 2588 2201 2628
rect 2205 2596 2207 2628
rect 2219 2596 2221 2628
rect 2205 2588 2221 2596
rect 2225 2588 2231 2628
rect 2235 2588 2237 2628
rect 2289 2608 2291 2628
rect 2295 2608 2297 2628
rect 2309 2608 2311 2628
rect 2299 2588 2311 2608
rect 2315 2588 2321 2628
rect 2325 2596 2327 2628
rect 2339 2596 2341 2628
rect 2325 2588 2341 2596
rect 2345 2588 2351 2628
rect 2355 2588 2357 2628
rect 2413 2596 2415 2636
rect 2419 2616 2421 2636
rect 2433 2616 2435 2636
rect 2439 2616 2445 2636
rect 2449 2616 2453 2636
rect 2465 2616 2467 2636
rect 2471 2616 2477 2636
rect 2481 2616 2483 2636
rect 2495 2616 2499 2636
rect 2503 2616 2505 2636
rect 2543 2616 2545 2636
rect 2549 2616 2553 2636
rect 2557 2616 2559 2636
rect 2571 2616 2573 2636
rect 2577 2616 2583 2636
rect 2587 2616 2589 2636
rect 2601 2616 2605 2636
rect 2419 2596 2429 2616
rect 2592 2596 2605 2616
rect 2609 2596 2611 2636
rect 2649 2608 2651 2628
rect 2655 2608 2657 2628
rect 2669 2608 2671 2628
rect 2659 2588 2671 2608
rect 2675 2588 2681 2628
rect 2685 2596 2687 2628
rect 2699 2596 2701 2628
rect 2685 2588 2701 2596
rect 2705 2588 2711 2628
rect 2715 2588 2717 2628
rect 2783 2616 2785 2636
rect 2789 2616 2791 2636
rect 2803 2616 2805 2636
rect 2809 2616 2811 2636
rect 2863 2588 2865 2628
rect 2869 2588 2875 2628
rect 2879 2596 2881 2628
rect 2893 2596 2895 2628
rect 2879 2588 2895 2596
rect 2899 2588 2905 2628
rect 2909 2608 2911 2628
rect 2923 2608 2925 2628
rect 2929 2608 2931 2628
rect 2909 2588 2921 2608
rect 2983 2596 2985 2636
rect 2989 2624 3005 2636
rect 2989 2596 2991 2624
rect 3003 2596 3005 2624
rect 3009 2596 3011 2636
rect 3023 2596 3025 2636
rect 3029 2606 3031 2636
rect 3043 2606 3045 2636
rect 3029 2596 3045 2606
rect 3049 2596 3051 2636
rect 3103 2616 3105 2636
rect 3109 2616 3111 2636
rect 3153 2596 3155 2636
rect 3159 2616 3161 2636
rect 3173 2616 3175 2636
rect 3179 2616 3185 2636
rect 3189 2616 3193 2636
rect 3205 2616 3207 2636
rect 3211 2616 3217 2636
rect 3221 2616 3223 2636
rect 3235 2616 3239 2636
rect 3243 2616 3245 2636
rect 3283 2616 3285 2636
rect 3289 2616 3293 2636
rect 3297 2616 3299 2636
rect 3311 2616 3313 2636
rect 3317 2616 3323 2636
rect 3327 2616 3329 2636
rect 3341 2616 3345 2636
rect 3159 2596 3169 2616
rect 3332 2596 3345 2616
rect 3349 2596 3351 2636
rect 3389 2616 3391 2636
rect 3395 2616 3397 2636
rect 3409 2616 3411 2636
rect 3415 2616 3417 2636
rect 3491 2596 3493 2636
rect 3497 2596 3503 2636
rect 3507 2596 3509 2636
rect 3549 2616 3551 2636
rect 3555 2616 3557 2636
rect 3610 2576 3612 2636
rect 3616 2576 3620 2636
rect 3624 2576 3628 2636
rect 3632 2578 3634 2636
rect 3632 2576 3646 2578
rect 3710 2576 3712 2636
rect 3716 2576 3720 2636
rect 3724 2576 3728 2636
rect 3732 2578 3734 2636
rect 3732 2576 3746 2578
rect 3846 2578 3848 2636
rect 3834 2576 3848 2578
rect 3852 2576 3856 2636
rect 3860 2576 3864 2636
rect 3868 2576 3870 2636
rect 3909 2596 3911 2636
rect 3915 2608 3917 2636
rect 3929 2608 3931 2636
rect 3915 2596 3931 2608
rect 3935 2596 3937 2636
rect 3949 2596 3951 2636
rect 3955 2596 3957 2636
rect 4012 2596 4014 2636
rect 4018 2596 4022 2636
rect 4026 2596 4028 2636
rect 4040 2616 4044 2636
rect 4048 2616 4050 2636
rect 4123 2616 4125 2636
rect 4129 2616 4131 2636
rect 4143 2616 4145 2636
rect 4149 2616 4151 2636
rect 4203 2596 4205 2636
rect 4209 2624 4225 2636
rect 4209 2596 4211 2624
rect 4223 2596 4225 2624
rect 4229 2596 4231 2636
rect 4243 2596 4245 2636
rect 4249 2606 4251 2636
rect 4263 2606 4265 2636
rect 4249 2596 4265 2606
rect 4269 2596 4271 2636
rect 4313 2596 4315 2636
rect 4319 2616 4321 2636
rect 4333 2616 4335 2636
rect 4339 2616 4345 2636
rect 4349 2616 4353 2636
rect 4365 2616 4367 2636
rect 4371 2616 4377 2636
rect 4381 2616 4383 2636
rect 4395 2616 4399 2636
rect 4403 2616 4405 2636
rect 4443 2616 4445 2636
rect 4449 2616 4453 2636
rect 4457 2616 4459 2636
rect 4471 2616 4473 2636
rect 4477 2616 4483 2636
rect 4487 2616 4489 2636
rect 4501 2616 4505 2636
rect 4319 2596 4329 2616
rect 4492 2596 4505 2616
rect 4509 2596 4511 2636
rect 4563 2616 4565 2636
rect 4569 2616 4571 2636
rect 4623 2596 4625 2636
rect 4629 2624 4645 2636
rect 4629 2596 4631 2624
rect 4643 2596 4645 2624
rect 4649 2596 4651 2636
rect 4663 2596 4665 2636
rect 4669 2606 4671 2636
rect 4683 2606 4685 2636
rect 4669 2596 4685 2606
rect 4689 2596 4691 2636
rect 4729 2608 4731 2628
rect 4735 2608 4737 2628
rect 4749 2608 4751 2628
rect 4739 2588 4751 2608
rect 4755 2588 4761 2628
rect 4765 2596 4767 2628
rect 4779 2596 4781 2628
rect 4765 2588 4781 2596
rect 4785 2588 4791 2628
rect 4795 2588 4797 2628
rect 4849 2596 4851 2636
rect 4855 2616 4859 2636
rect 4871 2616 4873 2636
rect 4877 2616 4883 2636
rect 4887 2616 4889 2636
rect 4901 2616 4903 2636
rect 4907 2616 4911 2636
rect 4915 2616 4917 2636
rect 4955 2616 4957 2636
rect 4961 2616 4965 2636
rect 4977 2616 4979 2636
rect 4983 2616 4989 2636
rect 4993 2616 4995 2636
rect 5007 2616 5011 2636
rect 5015 2616 5021 2636
rect 5025 2616 5027 2636
rect 5039 2616 5041 2636
rect 4855 2596 4868 2616
rect 5031 2596 5041 2616
rect 5045 2596 5047 2636
rect 5089 2616 5091 2636
rect 5095 2616 5097 2636
rect 5149 2596 5151 2636
rect 5155 2606 5157 2636
rect 5169 2606 5171 2636
rect 5155 2596 5171 2606
rect 5175 2596 5177 2636
rect 5189 2596 5191 2636
rect 5195 2624 5211 2636
rect 5195 2596 5197 2624
rect 5209 2596 5211 2624
rect 5215 2596 5217 2636
rect 5269 2596 5271 2636
rect 5275 2608 5277 2636
rect 5289 2608 5291 2636
rect 5275 2596 5291 2608
rect 5295 2596 5297 2636
rect 5309 2596 5311 2636
rect 5315 2596 5317 2636
rect 5369 2616 5371 2636
rect 5375 2616 5377 2636
rect 5389 2616 5391 2636
rect 5395 2616 5397 2636
rect 5463 2616 5465 2636
rect 5469 2616 5471 2636
rect 5483 2616 5485 2636
rect 5489 2616 5491 2636
rect 5529 2596 5531 2636
rect 5535 2596 5537 2636
rect 5549 2596 5551 2636
rect 5555 2596 5557 2636
rect 5569 2596 5571 2636
rect 5575 2596 5577 2636
rect 5589 2596 5591 2636
rect 5595 2596 5597 2636
rect 5609 2596 5611 2636
rect 5615 2596 5617 2636
rect 5629 2596 5631 2636
rect 5635 2596 5637 2636
rect 5649 2596 5651 2636
rect 5655 2596 5657 2636
rect 5669 2596 5671 2636
rect 5675 2596 5677 2636
rect 5743 2616 5745 2636
rect 5749 2616 5751 2636
rect 5763 2616 5765 2636
rect 5769 2616 5771 2636
rect 5809 2596 5811 2636
rect 5815 2608 5817 2636
rect 5829 2608 5831 2636
rect 5815 2596 5831 2608
rect 5835 2596 5837 2636
rect 5849 2596 5851 2636
rect 5855 2596 5857 2636
rect 5923 2596 5925 2636
rect 5929 2624 5945 2636
rect 5929 2596 5931 2624
rect 5943 2596 5945 2624
rect 5949 2596 5951 2636
rect 5963 2596 5965 2636
rect 5969 2606 5971 2636
rect 5983 2606 5985 2636
rect 5969 2596 5985 2606
rect 5989 2596 5991 2636
rect 6043 2616 6045 2636
rect 6049 2616 6051 2636
rect 6089 2596 6091 2636
rect 6095 2616 6099 2636
rect 6111 2616 6113 2636
rect 6117 2616 6123 2636
rect 6127 2616 6129 2636
rect 6141 2616 6143 2636
rect 6147 2616 6151 2636
rect 6155 2616 6157 2636
rect 6195 2616 6197 2636
rect 6201 2616 6205 2636
rect 6217 2616 6219 2636
rect 6223 2616 6229 2636
rect 6233 2616 6235 2636
rect 6247 2616 6251 2636
rect 6255 2616 6261 2636
rect 6265 2616 6267 2636
rect 6279 2616 6281 2636
rect 6095 2596 6108 2616
rect 6271 2596 6281 2616
rect 6285 2596 6287 2636
rect 6364 2596 6366 2636
rect 6370 2596 6374 2636
rect 6378 2596 6380 2636
rect 6392 2596 6394 2636
rect 6398 2596 6402 2636
rect 6406 2596 6408 2636
rect 6449 2596 6451 2636
rect 6455 2596 6457 2636
rect 6469 2596 6471 2636
rect 6475 2596 6477 2636
rect 6529 2616 6531 2636
rect 6535 2616 6537 2636
rect 6592 2596 6594 2636
rect 6598 2596 6602 2636
rect 6606 2596 6608 2636
rect 6620 2596 6622 2636
rect 6626 2596 6630 2636
rect 6634 2596 6636 2636
rect 33 2184 35 2224
rect 39 2204 49 2224
rect 212 2204 225 2224
rect 39 2184 41 2204
rect 53 2184 55 2204
rect 59 2184 65 2204
rect 69 2184 73 2204
rect 85 2184 87 2204
rect 91 2184 97 2204
rect 101 2184 103 2204
rect 115 2184 119 2204
rect 123 2184 125 2204
rect 163 2184 165 2204
rect 169 2184 173 2204
rect 177 2184 179 2204
rect 191 2184 193 2204
rect 197 2184 203 2204
rect 207 2184 209 2204
rect 221 2184 225 2204
rect 229 2184 231 2224
rect 281 2184 283 2224
rect 287 2184 289 2224
rect 301 2184 305 2204
rect 309 2184 311 2204
rect 363 2184 365 2224
rect 369 2184 371 2224
rect 423 2184 425 2204
rect 429 2184 431 2204
rect 483 2184 485 2204
rect 489 2184 491 2204
rect 503 2184 505 2204
rect 509 2184 511 2204
rect 549 2184 551 2224
rect 555 2212 571 2224
rect 555 2184 557 2212
rect 569 2184 571 2212
rect 575 2184 577 2224
rect 589 2184 591 2224
rect 595 2184 597 2224
rect 673 2184 675 2224
rect 679 2184 681 2224
rect 693 2184 695 2224
rect 699 2184 705 2224
rect 709 2184 711 2224
rect 750 2184 752 2244
rect 756 2184 760 2244
rect 764 2184 768 2244
rect 772 2242 786 2244
rect 772 2184 774 2242
rect 851 2184 853 2224
rect 857 2184 863 2224
rect 867 2184 869 2224
rect 929 2184 931 2224
rect 935 2204 948 2224
rect 1111 2204 1121 2224
rect 935 2184 939 2204
rect 951 2184 953 2204
rect 957 2184 963 2204
rect 967 2184 969 2204
rect 981 2184 983 2204
rect 987 2184 991 2204
rect 995 2184 997 2204
rect 1035 2184 1037 2204
rect 1041 2184 1045 2204
rect 1057 2184 1059 2204
rect 1063 2184 1069 2204
rect 1073 2184 1075 2204
rect 1087 2184 1091 2204
rect 1095 2184 1101 2204
rect 1105 2184 1107 2204
rect 1119 2184 1121 2204
rect 1125 2184 1127 2224
rect 1169 2184 1171 2204
rect 1175 2184 1177 2204
rect 1233 2184 1235 2224
rect 1239 2204 1249 2224
rect 1412 2204 1425 2224
rect 1239 2184 1241 2204
rect 1253 2184 1255 2204
rect 1259 2184 1265 2204
rect 1269 2184 1273 2204
rect 1285 2184 1287 2204
rect 1291 2184 1297 2204
rect 1301 2184 1303 2204
rect 1315 2184 1319 2204
rect 1323 2184 1325 2204
rect 1363 2184 1365 2204
rect 1369 2184 1373 2204
rect 1377 2184 1379 2204
rect 1391 2184 1393 2204
rect 1397 2184 1403 2204
rect 1407 2184 1409 2204
rect 1421 2184 1425 2204
rect 1429 2184 1431 2224
rect 1483 2184 1485 2204
rect 1489 2184 1491 2204
rect 1529 2184 1531 2224
rect 1535 2214 1551 2224
rect 1535 2184 1537 2214
rect 1549 2184 1551 2214
rect 1555 2184 1557 2224
rect 1569 2184 1571 2224
rect 1575 2196 1577 2224
rect 1589 2196 1591 2224
rect 1575 2184 1591 2196
rect 1595 2184 1597 2224
rect 1649 2184 1651 2224
rect 1655 2212 1671 2224
rect 1655 2184 1657 2212
rect 1669 2184 1671 2212
rect 1675 2184 1677 2224
rect 1689 2184 1691 2224
rect 1695 2184 1697 2224
rect 1763 2184 1765 2204
rect 1769 2184 1771 2204
rect 1783 2184 1785 2204
rect 1789 2184 1791 2204
rect 1843 2184 1845 2204
rect 1849 2184 1851 2204
rect 1863 2184 1865 2204
rect 1869 2184 1871 2204
rect 1923 2184 1925 2224
rect 1929 2196 1931 2224
rect 1943 2196 1945 2224
rect 1929 2184 1945 2196
rect 1949 2184 1951 2224
rect 1963 2184 1965 2224
rect 1969 2214 1985 2224
rect 1969 2184 1971 2214
rect 1983 2184 1985 2214
rect 1989 2184 1991 2224
rect 2043 2184 2045 2204
rect 2049 2184 2051 2204
rect 2093 2184 2095 2224
rect 2099 2204 2109 2224
rect 2272 2204 2285 2224
rect 2099 2184 2101 2204
rect 2113 2184 2115 2204
rect 2119 2184 2125 2204
rect 2129 2184 2133 2204
rect 2145 2184 2147 2204
rect 2151 2184 2157 2204
rect 2161 2184 2163 2204
rect 2175 2184 2179 2204
rect 2183 2184 2185 2204
rect 2223 2184 2225 2204
rect 2229 2184 2233 2204
rect 2237 2184 2239 2204
rect 2251 2184 2253 2204
rect 2257 2184 2263 2204
rect 2267 2184 2269 2204
rect 2281 2184 2285 2204
rect 2289 2184 2291 2224
rect 2534 2242 2548 2244
rect 2343 2184 2345 2204
rect 2349 2184 2351 2204
rect 2363 2184 2365 2204
rect 2369 2184 2371 2204
rect 2409 2184 2411 2224
rect 2415 2212 2431 2224
rect 2415 2184 2417 2212
rect 2429 2184 2431 2212
rect 2435 2184 2437 2224
rect 2449 2184 2451 2224
rect 2455 2184 2457 2224
rect 2546 2184 2548 2242
rect 2552 2184 2556 2244
rect 2560 2184 2564 2244
rect 2568 2184 2570 2244
rect 2630 2184 2632 2204
rect 2636 2184 2640 2204
rect 2652 2184 2654 2224
rect 2658 2184 2662 2224
rect 2666 2184 2668 2224
rect 2709 2184 2711 2224
rect 2715 2212 2731 2224
rect 2715 2184 2717 2212
rect 2729 2184 2731 2212
rect 2735 2184 2737 2224
rect 2749 2184 2751 2224
rect 2755 2184 2757 2224
rect 2823 2184 2825 2204
rect 2829 2184 2831 2204
rect 2843 2184 2845 2204
rect 2849 2184 2851 2204
rect 2889 2184 2891 2224
rect 2895 2204 2908 2224
rect 3071 2204 3081 2224
rect 2895 2184 2899 2204
rect 2911 2184 2913 2204
rect 2917 2184 2923 2204
rect 2927 2184 2929 2204
rect 2941 2184 2943 2204
rect 2947 2184 2951 2204
rect 2955 2184 2957 2204
rect 2995 2184 2997 2204
rect 3001 2184 3005 2204
rect 3017 2184 3019 2204
rect 3023 2184 3029 2204
rect 3033 2184 3035 2204
rect 3047 2184 3051 2204
rect 3055 2184 3061 2204
rect 3065 2184 3067 2204
rect 3079 2184 3081 2204
rect 3085 2184 3087 2224
rect 3129 2184 3131 2224
rect 3135 2212 3151 2224
rect 3135 2184 3137 2212
rect 3149 2184 3151 2212
rect 3155 2184 3157 2224
rect 3169 2184 3171 2224
rect 3175 2184 3177 2224
rect 3243 2184 3245 2224
rect 3249 2196 3251 2224
rect 3263 2196 3265 2224
rect 3249 2184 3265 2196
rect 3269 2184 3271 2224
rect 3283 2184 3285 2224
rect 3289 2214 3305 2224
rect 3289 2184 3291 2214
rect 3303 2184 3305 2214
rect 3309 2184 3311 2224
rect 3363 2184 3365 2204
rect 3369 2184 3371 2204
rect 3383 2184 3385 2204
rect 3389 2184 3391 2204
rect 3443 2184 3445 2204
rect 3449 2184 3451 2204
rect 3503 2184 3505 2204
rect 3509 2184 3511 2204
rect 3523 2184 3525 2204
rect 3529 2184 3531 2204
rect 3573 2184 3575 2224
rect 3579 2204 3589 2224
rect 3752 2204 3765 2224
rect 3579 2184 3581 2204
rect 3593 2184 3595 2204
rect 3599 2184 3605 2204
rect 3609 2184 3613 2204
rect 3625 2184 3627 2204
rect 3631 2184 3637 2204
rect 3641 2184 3643 2204
rect 3655 2184 3659 2204
rect 3663 2184 3665 2204
rect 3703 2184 3705 2204
rect 3709 2184 3713 2204
rect 3717 2184 3719 2204
rect 3731 2184 3733 2204
rect 3737 2184 3743 2204
rect 3747 2184 3749 2204
rect 3761 2184 3765 2204
rect 3769 2184 3771 2224
rect 3811 2184 3813 2224
rect 3817 2184 3823 2224
rect 3827 2184 3829 2224
rect 3890 2184 3892 2244
rect 3896 2184 3900 2244
rect 3904 2184 3908 2244
rect 3912 2242 3926 2244
rect 3912 2184 3914 2242
rect 3999 2212 4011 2232
rect 3989 2192 3991 2212
rect 3995 2192 3997 2212
rect 4009 2192 4011 2212
rect 4015 2192 4021 2232
rect 4025 2224 4041 2232
rect 4025 2192 4027 2224
rect 4039 2192 4041 2224
rect 4045 2192 4051 2232
rect 4055 2192 4057 2232
rect 4119 2212 4131 2232
rect 4109 2192 4111 2212
rect 4115 2192 4117 2212
rect 4129 2192 4131 2212
rect 4135 2192 4141 2232
rect 4145 2224 4161 2232
rect 4145 2192 4147 2224
rect 4159 2192 4161 2224
rect 4165 2192 4171 2232
rect 4175 2192 4177 2232
rect 4239 2212 4251 2232
rect 4229 2192 4231 2212
rect 4235 2192 4237 2212
rect 4249 2192 4251 2212
rect 4255 2192 4261 2232
rect 4265 2224 4281 2232
rect 4265 2192 4267 2224
rect 4279 2192 4281 2224
rect 4285 2192 4291 2232
rect 4295 2192 4297 2232
rect 4349 2184 4351 2204
rect 4355 2184 4359 2204
rect 4371 2184 4373 2224
rect 4377 2184 4379 2224
rect 4519 2212 4531 2232
rect 4443 2184 4445 2204
rect 4449 2184 4451 2204
rect 4463 2184 4465 2204
rect 4469 2184 4471 2204
rect 4509 2192 4511 2212
rect 4515 2192 4517 2212
rect 4529 2192 4531 2212
rect 4535 2192 4541 2232
rect 4545 2224 4561 2232
rect 4545 2192 4547 2224
rect 4559 2192 4561 2224
rect 4565 2192 4571 2232
rect 4575 2192 4577 2232
rect 4643 2192 4645 2232
rect 4649 2192 4655 2232
rect 4659 2224 4675 2232
rect 4659 2192 4661 2224
rect 4673 2192 4675 2224
rect 4679 2192 4685 2232
rect 4689 2212 4701 2232
rect 4759 2212 4771 2232
rect 4689 2192 4691 2212
rect 4703 2192 4705 2212
rect 4709 2192 4711 2212
rect 4749 2192 4751 2212
rect 4755 2192 4757 2212
rect 4769 2192 4771 2212
rect 4775 2192 4781 2232
rect 4785 2224 4801 2232
rect 4785 2192 4787 2224
rect 4799 2192 4801 2224
rect 4805 2192 4811 2232
rect 4815 2192 4817 2232
rect 4959 2212 4971 2232
rect 4869 2184 4871 2204
rect 4875 2184 4877 2204
rect 4889 2184 4891 2204
rect 4895 2184 4897 2204
rect 4949 2192 4951 2212
rect 4955 2192 4957 2212
rect 4969 2192 4971 2212
rect 4975 2192 4981 2232
rect 4985 2224 5001 2232
rect 4985 2192 4987 2224
rect 4999 2192 5001 2224
rect 5005 2192 5011 2232
rect 5015 2192 5017 2232
rect 5090 2184 5092 2204
rect 5096 2184 5100 2204
rect 5112 2184 5114 2224
rect 5118 2184 5122 2224
rect 5126 2184 5128 2224
rect 5169 2184 5171 2204
rect 5175 2184 5177 2204
rect 5229 2184 5231 2224
rect 5235 2214 5251 2224
rect 5235 2184 5237 2214
rect 5249 2184 5251 2214
rect 5255 2184 5257 2224
rect 5269 2184 5271 2224
rect 5275 2196 5277 2224
rect 5289 2196 5291 2224
rect 5275 2184 5291 2196
rect 5295 2184 5297 2224
rect 5363 2192 5365 2232
rect 5369 2192 5375 2232
rect 5379 2224 5395 2232
rect 5379 2192 5381 2224
rect 5393 2192 5395 2224
rect 5399 2192 5405 2232
rect 5409 2212 5421 2232
rect 5479 2212 5491 2232
rect 5409 2192 5411 2212
rect 5423 2192 5425 2212
rect 5429 2192 5431 2212
rect 5469 2192 5471 2212
rect 5475 2192 5477 2212
rect 5489 2192 5491 2212
rect 5495 2192 5501 2232
rect 5505 2224 5521 2232
rect 5505 2192 5507 2224
rect 5519 2192 5521 2224
rect 5525 2192 5531 2232
rect 5535 2192 5537 2232
rect 5734 2242 5748 2244
rect 5599 2212 5611 2232
rect 5589 2192 5591 2212
rect 5595 2192 5597 2212
rect 5609 2192 5611 2212
rect 5615 2192 5621 2232
rect 5625 2224 5641 2232
rect 5625 2192 5627 2224
rect 5639 2192 5641 2224
rect 5645 2192 5651 2232
rect 5655 2192 5657 2232
rect 5746 2184 5748 2242
rect 5752 2184 5756 2244
rect 5760 2184 5764 2244
rect 5768 2184 5770 2244
rect 5834 2242 5848 2244
rect 5846 2184 5848 2242
rect 5852 2184 5856 2244
rect 5860 2184 5864 2244
rect 5868 2184 5870 2244
rect 5923 2184 5925 2204
rect 5929 2184 5931 2204
rect 6004 2184 6006 2224
rect 6010 2184 6014 2224
rect 6018 2184 6020 2224
rect 6032 2184 6034 2224
rect 6038 2184 6042 2224
rect 6046 2184 6048 2224
rect 6103 2192 6105 2232
rect 6109 2192 6115 2232
rect 6119 2224 6135 2232
rect 6119 2192 6121 2224
rect 6133 2192 6135 2224
rect 6139 2192 6145 2232
rect 6149 2212 6161 2232
rect 6149 2192 6151 2212
rect 6163 2192 6165 2212
rect 6169 2192 6171 2212
rect 6223 2192 6225 2232
rect 6229 2192 6235 2232
rect 6239 2224 6255 2232
rect 6239 2192 6241 2224
rect 6253 2192 6255 2224
rect 6259 2192 6265 2232
rect 6269 2212 6281 2232
rect 6269 2192 6271 2212
rect 6283 2192 6285 2212
rect 6289 2192 6291 2212
rect 6329 2184 6331 2204
rect 6335 2184 6337 2204
rect 6389 2184 6391 2224
rect 6395 2212 6411 2224
rect 6395 2184 6397 2212
rect 6409 2184 6411 2212
rect 6415 2184 6417 2224
rect 6429 2184 6431 2224
rect 6435 2184 6437 2224
rect 6491 2184 6493 2224
rect 6497 2184 6503 2224
rect 6507 2184 6509 2224
rect 6572 2184 6574 2224
rect 6578 2184 6582 2224
rect 6586 2184 6588 2224
rect 6600 2184 6604 2204
rect 6608 2184 6610 2204
rect 6669 2184 6671 2204
rect 6675 2184 6677 2204
rect 43 2136 45 2156
rect 49 2136 51 2156
rect 63 2136 65 2156
rect 69 2136 71 2156
rect 131 2116 133 2156
rect 137 2116 143 2156
rect 147 2116 149 2156
rect 226 2098 228 2156
rect 214 2096 228 2098
rect 232 2096 236 2156
rect 240 2096 244 2156
rect 248 2096 250 2156
rect 326 2098 328 2156
rect 314 2096 328 2098
rect 332 2096 336 2156
rect 340 2096 344 2156
rect 348 2096 350 2156
rect 411 2116 413 2156
rect 417 2116 423 2156
rect 427 2116 429 2156
rect 470 2096 472 2156
rect 476 2096 480 2156
rect 484 2096 488 2156
rect 492 2098 494 2156
rect 583 2136 585 2156
rect 589 2136 591 2156
rect 603 2136 605 2156
rect 609 2136 611 2156
rect 492 2096 506 2098
rect 649 2116 651 2156
rect 655 2128 657 2156
rect 669 2128 671 2156
rect 655 2116 671 2128
rect 675 2116 677 2156
rect 689 2116 691 2156
rect 695 2116 697 2156
rect 750 2096 752 2156
rect 756 2096 760 2156
rect 764 2096 768 2156
rect 772 2098 774 2156
rect 849 2136 851 2156
rect 855 2136 857 2156
rect 869 2136 871 2156
rect 875 2136 877 2156
rect 772 2096 786 2098
rect 951 2116 953 2156
rect 957 2116 963 2156
rect 967 2116 969 2156
rect 1009 2128 1011 2148
rect 1015 2128 1017 2148
rect 1029 2128 1031 2148
rect 1019 2108 1031 2128
rect 1035 2108 1041 2148
rect 1045 2116 1047 2148
rect 1059 2116 1061 2148
rect 1045 2108 1061 2116
rect 1065 2108 1071 2148
rect 1075 2108 1077 2148
rect 1133 2116 1135 2156
rect 1139 2136 1141 2156
rect 1153 2136 1155 2156
rect 1159 2136 1165 2156
rect 1169 2136 1173 2156
rect 1185 2136 1187 2156
rect 1191 2136 1197 2156
rect 1201 2136 1203 2156
rect 1215 2136 1219 2156
rect 1223 2136 1225 2156
rect 1263 2136 1265 2156
rect 1269 2136 1273 2156
rect 1277 2136 1279 2156
rect 1291 2136 1293 2156
rect 1297 2136 1303 2156
rect 1307 2136 1309 2156
rect 1321 2136 1325 2156
rect 1139 2116 1149 2136
rect 1312 2116 1325 2136
rect 1329 2116 1331 2156
rect 1369 2136 1371 2156
rect 1375 2136 1377 2156
rect 1429 2116 1431 2156
rect 1435 2126 1437 2156
rect 1449 2126 1451 2156
rect 1435 2116 1451 2126
rect 1455 2116 1457 2156
rect 1469 2116 1471 2156
rect 1475 2144 1491 2156
rect 1475 2116 1477 2144
rect 1489 2116 1491 2144
rect 1495 2116 1497 2156
rect 1563 2116 1565 2156
rect 1569 2116 1571 2156
rect 1583 2116 1585 2156
rect 1589 2128 1591 2156
rect 1603 2128 1605 2156
rect 1589 2116 1605 2128
rect 1609 2116 1611 2156
rect 1663 2116 1665 2156
rect 1669 2116 1671 2156
rect 1683 2116 1685 2156
rect 1689 2128 1691 2156
rect 1703 2128 1705 2156
rect 1689 2116 1705 2128
rect 1709 2116 1711 2156
rect 1763 2136 1765 2156
rect 1769 2136 1771 2156
rect 1783 2136 1785 2156
rect 1789 2136 1791 2156
rect 1843 2116 1845 2156
rect 1849 2116 1851 2156
rect 1863 2116 1865 2156
rect 1869 2128 1871 2156
rect 1883 2128 1885 2156
rect 1869 2116 1885 2128
rect 1889 2116 1891 2156
rect 1943 2108 1945 2148
rect 1949 2108 1955 2148
rect 1959 2116 1961 2148
rect 1973 2116 1975 2148
rect 1959 2108 1975 2116
rect 1979 2108 1985 2148
rect 1989 2128 1991 2148
rect 2003 2128 2005 2148
rect 2009 2128 2011 2148
rect 1989 2108 2001 2128
rect 2063 2108 2065 2148
rect 2069 2108 2075 2148
rect 2079 2116 2081 2148
rect 2093 2116 2095 2148
rect 2079 2108 2095 2116
rect 2099 2108 2105 2148
rect 2109 2128 2111 2148
rect 2123 2128 2125 2148
rect 2129 2128 2131 2148
rect 2109 2108 2121 2128
rect 2173 2116 2175 2156
rect 2179 2136 2181 2156
rect 2193 2136 2195 2156
rect 2199 2136 2205 2156
rect 2209 2136 2213 2156
rect 2225 2136 2227 2156
rect 2231 2136 2237 2156
rect 2241 2136 2243 2156
rect 2255 2136 2259 2156
rect 2263 2136 2265 2156
rect 2303 2136 2305 2156
rect 2309 2136 2313 2156
rect 2317 2136 2319 2156
rect 2331 2136 2333 2156
rect 2337 2136 2343 2156
rect 2347 2136 2349 2156
rect 2361 2136 2365 2156
rect 2179 2116 2189 2136
rect 2352 2116 2365 2136
rect 2369 2116 2371 2156
rect 2423 2116 2425 2156
rect 2429 2116 2431 2156
rect 2443 2116 2445 2156
rect 2449 2128 2451 2156
rect 2463 2128 2465 2156
rect 2449 2116 2465 2128
rect 2469 2116 2471 2156
rect 2509 2136 2511 2156
rect 2515 2136 2517 2156
rect 2529 2136 2531 2156
rect 2535 2136 2537 2156
rect 2626 2098 2628 2156
rect 2614 2096 2628 2098
rect 2632 2096 2636 2156
rect 2640 2096 2644 2156
rect 2648 2096 2650 2156
rect 2689 2128 2691 2148
rect 2695 2128 2697 2148
rect 2709 2128 2711 2148
rect 2699 2108 2711 2128
rect 2715 2108 2721 2148
rect 2725 2116 2727 2148
rect 2739 2116 2741 2148
rect 2725 2108 2741 2116
rect 2745 2108 2751 2148
rect 2755 2108 2757 2148
rect 2823 2108 2825 2148
rect 2829 2108 2835 2148
rect 2839 2116 2841 2148
rect 2853 2116 2855 2148
rect 2839 2108 2855 2116
rect 2859 2108 2865 2148
rect 2869 2128 2871 2148
rect 2883 2128 2885 2148
rect 2889 2128 2891 2148
rect 2929 2136 2931 2156
rect 2935 2136 2937 2156
rect 2869 2108 2881 2128
rect 2989 2116 2991 2156
rect 2995 2126 2997 2156
rect 3009 2126 3011 2156
rect 2995 2116 3011 2126
rect 3015 2116 3017 2156
rect 3029 2116 3031 2156
rect 3035 2144 3051 2156
rect 3035 2116 3037 2144
rect 3049 2116 3051 2144
rect 3055 2116 3057 2156
rect 3130 2136 3132 2156
rect 3136 2136 3140 2156
rect 3152 2116 3154 2156
rect 3158 2116 3162 2156
rect 3166 2116 3168 2156
rect 3209 2136 3211 2156
rect 3215 2136 3217 2156
rect 3269 2116 3271 2156
rect 3275 2126 3277 2156
rect 3289 2126 3291 2156
rect 3275 2116 3291 2126
rect 3295 2116 3297 2156
rect 3309 2116 3311 2156
rect 3315 2144 3331 2156
rect 3315 2116 3317 2144
rect 3329 2116 3331 2144
rect 3335 2116 3337 2156
rect 3389 2136 3391 2156
rect 3395 2136 3397 2156
rect 3409 2136 3411 2156
rect 3415 2136 3417 2156
rect 3473 2116 3475 2156
rect 3479 2136 3481 2156
rect 3493 2136 3495 2156
rect 3499 2136 3505 2156
rect 3509 2136 3513 2156
rect 3525 2136 3527 2156
rect 3531 2136 3537 2156
rect 3541 2136 3543 2156
rect 3555 2136 3559 2156
rect 3563 2136 3565 2156
rect 3603 2136 3605 2156
rect 3609 2136 3613 2156
rect 3617 2136 3619 2156
rect 3631 2136 3633 2156
rect 3637 2136 3643 2156
rect 3647 2136 3649 2156
rect 3661 2136 3665 2156
rect 3479 2116 3489 2136
rect 3652 2116 3665 2136
rect 3669 2116 3671 2156
rect 3723 2136 3725 2156
rect 3729 2136 3731 2156
rect 3743 2136 3745 2156
rect 3749 2136 3751 2156
rect 3803 2116 3805 2156
rect 3809 2144 3825 2156
rect 3809 2116 3811 2144
rect 3823 2116 3825 2144
rect 3829 2116 3831 2156
rect 3843 2116 3845 2156
rect 3849 2126 3851 2156
rect 3863 2126 3865 2156
rect 3849 2116 3865 2126
rect 3869 2116 3871 2156
rect 3923 2136 3925 2156
rect 3929 2136 3931 2156
rect 3969 2116 3971 2156
rect 3975 2128 3977 2156
rect 3989 2128 3991 2156
rect 3975 2116 3991 2128
rect 3995 2116 3997 2156
rect 4009 2116 4011 2156
rect 4015 2116 4017 2156
rect 4071 2116 4073 2156
rect 4077 2116 4083 2156
rect 4087 2116 4089 2156
rect 4163 2136 4165 2156
rect 4169 2136 4171 2156
rect 4183 2136 4185 2156
rect 4189 2136 4191 2156
rect 4233 2116 4235 2156
rect 4239 2136 4241 2156
rect 4253 2136 4255 2156
rect 4259 2136 4265 2156
rect 4269 2136 4273 2156
rect 4285 2136 4287 2156
rect 4291 2136 4297 2156
rect 4301 2136 4303 2156
rect 4315 2136 4319 2156
rect 4323 2136 4325 2156
rect 4363 2136 4365 2156
rect 4369 2136 4373 2156
rect 4377 2136 4379 2156
rect 4391 2136 4393 2156
rect 4397 2136 4403 2156
rect 4407 2136 4409 2156
rect 4421 2136 4425 2156
rect 4239 2116 4249 2136
rect 4412 2116 4425 2136
rect 4429 2116 4431 2156
rect 4469 2136 4471 2156
rect 4475 2136 4477 2156
rect 4529 2116 4531 2156
rect 4535 2126 4537 2156
rect 4549 2126 4551 2156
rect 4535 2116 4551 2126
rect 4555 2116 4557 2156
rect 4569 2116 4571 2156
rect 4575 2144 4591 2156
rect 4575 2116 4577 2144
rect 4589 2116 4591 2144
rect 4595 2116 4597 2156
rect 4649 2136 4651 2156
rect 4655 2136 4657 2156
rect 4669 2136 4671 2156
rect 4675 2136 4677 2156
rect 4743 2116 4745 2156
rect 4749 2116 4751 2156
rect 4763 2116 4765 2156
rect 4769 2128 4771 2156
rect 4783 2128 4785 2156
rect 4769 2116 4785 2128
rect 4789 2116 4791 2156
rect 4843 2136 4845 2156
rect 4849 2136 4851 2156
rect 4863 2136 4865 2156
rect 4869 2136 4871 2156
rect 4909 2116 4911 2156
rect 4915 2126 4917 2156
rect 4929 2126 4931 2156
rect 4915 2116 4931 2126
rect 4935 2116 4937 2156
rect 4949 2116 4951 2156
rect 4955 2144 4971 2156
rect 4955 2116 4957 2144
rect 4969 2116 4971 2144
rect 4975 2116 4977 2156
rect 5051 2116 5053 2156
rect 5057 2116 5063 2156
rect 5067 2116 5069 2156
rect 5123 2136 5125 2156
rect 5129 2136 5131 2156
rect 5143 2136 5145 2156
rect 5149 2136 5151 2156
rect 5189 2136 5191 2156
rect 5195 2136 5197 2156
rect 5209 2136 5211 2156
rect 5215 2136 5217 2156
rect 5229 2136 5231 2156
rect 5219 2116 5231 2136
rect 5235 2116 5237 2156
rect 5303 2116 5305 2156
rect 5309 2144 5325 2156
rect 5309 2116 5311 2144
rect 5323 2116 5325 2144
rect 5329 2116 5331 2156
rect 5343 2116 5345 2156
rect 5349 2126 5351 2156
rect 5363 2126 5365 2156
rect 5349 2116 5365 2126
rect 5369 2116 5371 2156
rect 5409 2116 5411 2156
rect 5415 2126 5417 2156
rect 5429 2126 5431 2156
rect 5415 2116 5431 2126
rect 5435 2116 5437 2156
rect 5449 2116 5451 2156
rect 5455 2144 5471 2156
rect 5455 2116 5457 2144
rect 5469 2116 5471 2144
rect 5475 2116 5477 2156
rect 5543 2136 5545 2156
rect 5549 2136 5551 2156
rect 5563 2136 5565 2156
rect 5569 2136 5571 2156
rect 5623 2116 5625 2156
rect 5629 2144 5645 2156
rect 5629 2116 5631 2144
rect 5643 2116 5645 2144
rect 5649 2116 5651 2156
rect 5663 2116 5665 2156
rect 5669 2126 5671 2156
rect 5683 2126 5685 2156
rect 5669 2116 5685 2126
rect 5689 2116 5691 2156
rect 5743 2136 5745 2156
rect 5749 2136 5751 2156
rect 5791 2116 5793 2156
rect 5797 2116 5803 2156
rect 5807 2116 5809 2156
rect 5869 2116 5871 2156
rect 5875 2136 5879 2156
rect 5891 2136 5893 2156
rect 5897 2136 5903 2156
rect 5907 2136 5909 2156
rect 5921 2136 5923 2156
rect 5927 2136 5931 2156
rect 5935 2136 5937 2156
rect 5975 2136 5977 2156
rect 5981 2136 5985 2156
rect 5997 2136 5999 2156
rect 6003 2136 6009 2156
rect 6013 2136 6015 2156
rect 6027 2136 6031 2156
rect 6035 2136 6041 2156
rect 6045 2136 6047 2156
rect 6059 2136 6061 2156
rect 5875 2116 5888 2136
rect 6051 2116 6061 2136
rect 6065 2116 6067 2156
rect 6113 2116 6115 2156
rect 6119 2136 6121 2156
rect 6133 2136 6135 2156
rect 6139 2136 6145 2156
rect 6149 2136 6153 2156
rect 6165 2136 6167 2156
rect 6171 2136 6177 2156
rect 6181 2136 6183 2156
rect 6195 2136 6199 2156
rect 6203 2136 6205 2156
rect 6243 2136 6245 2156
rect 6249 2136 6253 2156
rect 6257 2136 6259 2156
rect 6271 2136 6273 2156
rect 6277 2136 6283 2156
rect 6287 2136 6289 2156
rect 6301 2136 6305 2156
rect 6119 2116 6129 2136
rect 6292 2116 6305 2136
rect 6309 2116 6311 2156
rect 6349 2128 6351 2148
rect 6355 2128 6357 2148
rect 6369 2128 6371 2148
rect 6359 2108 6371 2128
rect 6375 2108 6381 2148
rect 6385 2116 6387 2148
rect 6399 2116 6401 2148
rect 6385 2108 6401 2116
rect 6405 2108 6411 2148
rect 6415 2108 6417 2148
rect 6472 2116 6474 2156
rect 6478 2116 6482 2156
rect 6486 2116 6488 2156
rect 6500 2136 6504 2156
rect 6508 2136 6510 2156
rect 6569 2116 6571 2156
rect 6575 2128 6577 2156
rect 6589 2128 6591 2156
rect 6575 2116 6591 2128
rect 6595 2116 6597 2156
rect 6609 2116 6611 2156
rect 6615 2116 6617 2156
rect 43 1704 45 1724
rect 49 1704 51 1724
rect 89 1704 91 1744
rect 95 1724 108 1744
rect 271 1724 281 1744
rect 95 1704 99 1724
rect 111 1704 113 1724
rect 117 1704 123 1724
rect 127 1704 129 1724
rect 141 1704 143 1724
rect 147 1704 151 1724
rect 155 1704 157 1724
rect 195 1704 197 1724
rect 201 1704 205 1724
rect 217 1704 219 1724
rect 223 1704 229 1724
rect 233 1704 235 1724
rect 247 1704 251 1724
rect 255 1704 261 1724
rect 265 1704 267 1724
rect 279 1704 281 1724
rect 285 1704 287 1744
rect 329 1704 331 1724
rect 335 1704 337 1724
rect 349 1704 351 1724
rect 355 1704 357 1724
rect 423 1704 425 1724
rect 429 1704 431 1724
rect 443 1704 445 1724
rect 449 1704 451 1724
rect 503 1704 505 1724
rect 509 1704 511 1724
rect 563 1704 565 1744
rect 569 1704 571 1744
rect 583 1704 585 1744
rect 589 1732 605 1744
rect 589 1704 591 1732
rect 603 1704 605 1732
rect 609 1704 611 1744
rect 649 1704 651 1744
rect 655 1724 668 1744
rect 914 1762 928 1764
rect 831 1724 841 1744
rect 655 1704 659 1724
rect 671 1704 673 1724
rect 677 1704 683 1724
rect 687 1704 689 1724
rect 701 1704 703 1724
rect 707 1704 711 1724
rect 715 1704 717 1724
rect 755 1704 757 1724
rect 761 1704 765 1724
rect 777 1704 779 1724
rect 783 1704 789 1724
rect 793 1704 795 1724
rect 807 1704 811 1724
rect 815 1704 821 1724
rect 825 1704 827 1724
rect 839 1704 841 1724
rect 845 1704 847 1744
rect 926 1704 928 1762
rect 932 1704 936 1764
rect 940 1704 944 1764
rect 948 1704 950 1764
rect 989 1704 991 1744
rect 995 1704 1001 1744
rect 1005 1704 1007 1744
rect 1019 1704 1021 1744
rect 1025 1704 1027 1744
rect 1354 1762 1368 1764
rect 1089 1704 1091 1724
rect 1095 1704 1097 1724
rect 1149 1704 1151 1744
rect 1155 1732 1171 1744
rect 1155 1704 1157 1732
rect 1169 1704 1171 1732
rect 1175 1704 1177 1744
rect 1189 1704 1191 1744
rect 1195 1704 1197 1744
rect 1271 1704 1273 1744
rect 1277 1704 1283 1744
rect 1287 1704 1289 1744
rect 1366 1704 1368 1762
rect 1372 1704 1376 1764
rect 1380 1704 1384 1764
rect 1388 1704 1390 1764
rect 1429 1704 1431 1724
rect 1435 1704 1437 1724
rect 1493 1704 1495 1744
rect 1499 1724 1509 1744
rect 1672 1724 1685 1744
rect 1499 1704 1501 1724
rect 1513 1704 1515 1724
rect 1519 1704 1525 1724
rect 1529 1704 1533 1724
rect 1545 1704 1547 1724
rect 1551 1704 1557 1724
rect 1561 1704 1563 1724
rect 1575 1704 1579 1724
rect 1583 1704 1585 1724
rect 1623 1704 1625 1724
rect 1629 1704 1633 1724
rect 1637 1704 1639 1724
rect 1651 1704 1653 1724
rect 1657 1704 1663 1724
rect 1667 1704 1669 1724
rect 1681 1704 1685 1724
rect 1689 1704 1691 1744
rect 1729 1704 1731 1724
rect 1735 1704 1737 1724
rect 1789 1704 1791 1744
rect 1795 1734 1811 1744
rect 1795 1704 1797 1734
rect 1809 1704 1811 1734
rect 1815 1704 1817 1744
rect 1829 1704 1831 1744
rect 1835 1716 1837 1744
rect 1849 1716 1851 1744
rect 1835 1704 1851 1716
rect 1855 1704 1857 1744
rect 1909 1704 1911 1724
rect 1915 1704 1917 1724
rect 1929 1704 1931 1724
rect 1935 1704 1937 1724
rect 1989 1704 1991 1744
rect 1995 1732 2011 1744
rect 1995 1704 1997 1732
rect 2009 1704 2011 1732
rect 2015 1704 2017 1744
rect 2029 1704 2031 1744
rect 2035 1704 2037 1744
rect 2089 1704 2091 1744
rect 2095 1724 2108 1744
rect 2271 1724 2281 1744
rect 2095 1704 2099 1724
rect 2111 1704 2113 1724
rect 2117 1704 2123 1724
rect 2127 1704 2129 1724
rect 2141 1704 2143 1724
rect 2147 1704 2151 1724
rect 2155 1704 2157 1724
rect 2195 1704 2197 1724
rect 2201 1704 2205 1724
rect 2217 1704 2219 1724
rect 2223 1704 2229 1724
rect 2233 1704 2235 1724
rect 2247 1704 2251 1724
rect 2255 1704 2261 1724
rect 2265 1704 2267 1724
rect 2279 1704 2281 1724
rect 2285 1704 2287 1744
rect 2343 1704 2345 1744
rect 2349 1716 2351 1744
rect 2363 1716 2365 1744
rect 2349 1704 2365 1716
rect 2369 1704 2371 1744
rect 2383 1704 2385 1744
rect 2389 1734 2405 1744
rect 2389 1704 2391 1734
rect 2403 1704 2405 1734
rect 2409 1704 2411 1744
rect 2449 1704 2451 1724
rect 2455 1704 2457 1724
rect 2509 1704 2511 1724
rect 2515 1704 2517 1724
rect 2529 1704 2531 1724
rect 2535 1704 2537 1724
rect 2589 1704 2591 1744
rect 2595 1724 2608 1744
rect 2771 1724 2781 1744
rect 2595 1704 2599 1724
rect 2611 1704 2613 1724
rect 2617 1704 2623 1724
rect 2627 1704 2629 1724
rect 2641 1704 2643 1724
rect 2647 1704 2651 1724
rect 2655 1704 2657 1724
rect 2695 1704 2697 1724
rect 2701 1704 2705 1724
rect 2717 1704 2719 1724
rect 2723 1704 2729 1724
rect 2733 1704 2735 1724
rect 2747 1704 2751 1724
rect 2755 1704 2761 1724
rect 2765 1704 2767 1724
rect 2779 1704 2781 1724
rect 2785 1704 2787 1744
rect 2830 1704 2832 1764
rect 2836 1704 2840 1764
rect 2844 1704 2848 1764
rect 2852 1762 2866 1764
rect 2852 1704 2854 1762
rect 2943 1704 2945 1744
rect 2949 1704 2951 1744
rect 2963 1704 2965 1744
rect 2969 1732 2985 1744
rect 2969 1704 2971 1732
rect 2983 1704 2985 1732
rect 2989 1704 2991 1744
rect 3029 1704 3031 1724
rect 3035 1704 3037 1724
rect 3049 1704 3051 1724
rect 3055 1704 3057 1724
rect 3130 1704 3132 1724
rect 3136 1704 3140 1724
rect 3152 1704 3154 1744
rect 3158 1704 3162 1744
rect 3166 1704 3168 1744
rect 3230 1704 3232 1724
rect 3236 1704 3240 1724
rect 3252 1704 3254 1744
rect 3258 1704 3262 1744
rect 3266 1704 3268 1744
rect 3321 1704 3323 1744
rect 3327 1704 3329 1744
rect 3341 1704 3345 1724
rect 3349 1704 3351 1724
rect 3411 1704 3413 1744
rect 3417 1704 3423 1744
rect 3427 1704 3429 1744
rect 3469 1704 3471 1724
rect 3475 1704 3477 1724
rect 3489 1704 3491 1724
rect 3495 1704 3497 1724
rect 3551 1704 3553 1744
rect 3557 1704 3563 1744
rect 3567 1704 3569 1744
rect 3629 1704 3631 1744
rect 3635 1732 3651 1744
rect 3635 1704 3637 1732
rect 3649 1704 3651 1732
rect 3655 1704 3657 1744
rect 3669 1704 3671 1744
rect 3675 1704 3677 1744
rect 3751 1704 3753 1744
rect 3757 1704 3763 1744
rect 3767 1704 3769 1744
rect 3823 1704 3825 1724
rect 3829 1704 3831 1724
rect 3871 1704 3873 1744
rect 3877 1704 3883 1744
rect 3887 1704 3889 1744
rect 3949 1704 3951 1724
rect 3955 1704 3957 1724
rect 3969 1704 3971 1724
rect 3975 1704 3977 1724
rect 4029 1704 4031 1744
rect 4035 1734 4051 1744
rect 4035 1704 4037 1734
rect 4049 1704 4051 1734
rect 4055 1704 4057 1744
rect 4069 1704 4071 1744
rect 4075 1716 4077 1744
rect 4089 1716 4091 1744
rect 4075 1704 4091 1716
rect 4095 1704 4097 1744
rect 4163 1704 4165 1724
rect 4169 1704 4171 1724
rect 4183 1704 4185 1724
rect 4189 1704 4191 1724
rect 4229 1704 4231 1744
rect 4235 1732 4251 1744
rect 4235 1704 4237 1732
rect 4249 1704 4251 1732
rect 4255 1704 4257 1744
rect 4269 1704 4271 1744
rect 4275 1704 4277 1744
rect 4329 1704 4331 1744
rect 4335 1704 4337 1744
rect 4349 1704 4351 1744
rect 4355 1704 4357 1744
rect 4409 1704 4411 1744
rect 4415 1732 4431 1744
rect 4415 1704 4417 1732
rect 4429 1704 4431 1732
rect 4435 1704 4437 1744
rect 4449 1704 4451 1744
rect 4455 1704 4457 1744
rect 4523 1704 4525 1724
rect 4529 1704 4531 1724
rect 4543 1704 4545 1724
rect 4549 1704 4551 1724
rect 4603 1704 4605 1744
rect 4609 1716 4611 1744
rect 4623 1716 4625 1744
rect 4609 1704 4625 1716
rect 4629 1704 4631 1744
rect 4643 1704 4645 1744
rect 4649 1734 4665 1744
rect 4649 1704 4651 1734
rect 4663 1704 4665 1734
rect 4669 1704 4671 1744
rect 4723 1704 4725 1724
rect 4729 1704 4731 1724
rect 4769 1704 4771 1744
rect 4775 1724 4788 1744
rect 4951 1724 4961 1744
rect 4775 1704 4779 1724
rect 4791 1704 4793 1724
rect 4797 1704 4803 1724
rect 4807 1704 4809 1724
rect 4821 1704 4823 1724
rect 4827 1704 4831 1724
rect 4835 1704 4837 1724
rect 4875 1704 4877 1724
rect 4881 1704 4885 1724
rect 4897 1704 4899 1724
rect 4903 1704 4909 1724
rect 4913 1704 4915 1724
rect 4927 1704 4931 1724
rect 4935 1704 4941 1724
rect 4945 1704 4947 1724
rect 4959 1704 4961 1724
rect 4965 1704 4967 1744
rect 5012 1704 5014 1744
rect 5018 1704 5022 1744
rect 5026 1704 5028 1744
rect 5040 1704 5044 1724
rect 5048 1704 5050 1724
rect 5109 1704 5111 1724
rect 5115 1704 5117 1724
rect 5129 1704 5131 1724
rect 5135 1704 5137 1724
rect 5189 1704 5191 1744
rect 5195 1732 5211 1744
rect 5195 1704 5197 1732
rect 5209 1704 5211 1732
rect 5215 1704 5217 1744
rect 5229 1704 5231 1744
rect 5235 1704 5237 1744
rect 5290 1704 5292 1764
rect 5296 1704 5300 1764
rect 5304 1704 5308 1764
rect 5312 1762 5326 1764
rect 5312 1704 5314 1762
rect 5389 1704 5391 1724
rect 5395 1704 5399 1724
rect 5411 1704 5413 1744
rect 5417 1704 5419 1744
rect 5483 1704 5485 1724
rect 5489 1704 5491 1724
rect 5543 1704 5545 1744
rect 5549 1704 5551 1744
rect 5603 1704 5605 1744
rect 5609 1704 5611 1744
rect 5623 1704 5625 1744
rect 5629 1732 5645 1744
rect 5629 1704 5631 1732
rect 5643 1704 5645 1732
rect 5649 1704 5651 1744
rect 5691 1704 5693 1744
rect 5697 1704 5703 1744
rect 5707 1704 5709 1744
rect 5804 1704 5806 1744
rect 5810 1704 5814 1744
rect 5818 1704 5820 1744
rect 5832 1704 5834 1744
rect 5838 1704 5842 1744
rect 5846 1704 5848 1744
rect 5889 1704 5891 1724
rect 5895 1704 5899 1724
rect 5911 1704 5913 1744
rect 5917 1704 5919 1744
rect 5983 1704 5985 1744
rect 5989 1704 5991 1744
rect 6003 1704 6005 1744
rect 6009 1732 6025 1744
rect 6009 1704 6011 1732
rect 6023 1704 6025 1732
rect 6029 1704 6031 1744
rect 6083 1704 6085 1744
rect 6089 1716 6091 1744
rect 6103 1716 6105 1744
rect 6089 1704 6105 1716
rect 6109 1704 6111 1744
rect 6123 1704 6125 1744
rect 6129 1734 6145 1744
rect 6129 1704 6131 1734
rect 6143 1704 6145 1734
rect 6149 1704 6151 1744
rect 6199 1732 6211 1752
rect 6189 1712 6191 1732
rect 6195 1712 6197 1732
rect 6209 1712 6211 1732
rect 6215 1712 6221 1752
rect 6225 1744 6241 1752
rect 6225 1712 6227 1744
rect 6239 1712 6241 1744
rect 6245 1712 6251 1752
rect 6255 1712 6257 1752
rect 6319 1732 6331 1752
rect 6309 1712 6311 1732
rect 6315 1712 6317 1732
rect 6329 1712 6331 1732
rect 6335 1712 6341 1752
rect 6345 1744 6361 1752
rect 6345 1712 6347 1744
rect 6359 1712 6361 1744
rect 6365 1712 6371 1752
rect 6375 1712 6377 1752
rect 6429 1704 6431 1724
rect 6435 1704 6437 1724
rect 6489 1704 6491 1744
rect 6495 1732 6511 1744
rect 6495 1704 6497 1732
rect 6509 1704 6511 1732
rect 6515 1704 6517 1744
rect 6529 1704 6531 1744
rect 6535 1704 6537 1744
rect 6611 1704 6613 1744
rect 6617 1704 6623 1744
rect 6627 1704 6629 1744
rect 43 1656 45 1676
rect 49 1656 51 1676
rect 63 1656 65 1676
rect 69 1656 71 1676
rect 123 1636 125 1676
rect 129 1636 131 1676
rect 143 1636 145 1676
rect 149 1636 151 1676
rect 163 1636 165 1676
rect 169 1636 171 1676
rect 183 1636 185 1676
rect 189 1636 191 1676
rect 203 1636 205 1676
rect 209 1636 211 1676
rect 223 1636 225 1676
rect 229 1636 231 1676
rect 243 1636 245 1676
rect 249 1636 251 1676
rect 263 1636 265 1676
rect 269 1636 271 1676
rect 313 1636 315 1676
rect 319 1656 321 1676
rect 333 1656 335 1676
rect 339 1656 345 1676
rect 349 1656 353 1676
rect 365 1656 367 1676
rect 371 1656 377 1676
rect 381 1656 383 1676
rect 395 1656 399 1676
rect 403 1656 405 1676
rect 443 1656 445 1676
rect 449 1656 453 1676
rect 457 1656 459 1676
rect 471 1656 473 1676
rect 477 1656 483 1676
rect 487 1656 489 1676
rect 501 1656 505 1676
rect 319 1636 329 1656
rect 492 1636 505 1656
rect 509 1636 511 1676
rect 563 1656 565 1676
rect 569 1656 571 1676
rect 610 1616 612 1676
rect 616 1616 620 1676
rect 624 1616 628 1676
rect 632 1618 634 1676
rect 712 1636 714 1676
rect 718 1636 722 1676
rect 726 1636 728 1676
rect 740 1656 744 1676
rect 748 1656 750 1676
rect 632 1616 646 1618
rect 813 1636 815 1676
rect 819 1656 821 1676
rect 833 1656 835 1676
rect 839 1656 845 1676
rect 849 1656 853 1676
rect 865 1656 867 1676
rect 871 1656 877 1676
rect 881 1656 883 1676
rect 895 1656 899 1676
rect 903 1656 905 1676
rect 943 1656 945 1676
rect 949 1656 953 1676
rect 957 1656 959 1676
rect 971 1656 973 1676
rect 977 1656 983 1676
rect 987 1656 989 1676
rect 1001 1656 1005 1676
rect 819 1636 829 1656
rect 992 1636 1005 1656
rect 1009 1636 1011 1676
rect 1063 1656 1065 1676
rect 1069 1656 1071 1676
rect 1109 1636 1111 1676
rect 1115 1646 1117 1676
rect 1129 1646 1131 1676
rect 1115 1636 1131 1646
rect 1135 1636 1137 1676
rect 1149 1636 1151 1676
rect 1155 1664 1171 1676
rect 1155 1636 1157 1664
rect 1169 1636 1171 1664
rect 1175 1636 1177 1676
rect 1243 1636 1245 1676
rect 1249 1636 1251 1676
rect 1263 1636 1265 1676
rect 1269 1648 1271 1676
rect 1283 1648 1285 1676
rect 1269 1636 1285 1648
rect 1289 1636 1291 1676
rect 1343 1656 1345 1676
rect 1349 1656 1351 1676
rect 1363 1656 1365 1676
rect 1369 1656 1371 1676
rect 1423 1628 1425 1668
rect 1429 1628 1435 1668
rect 1439 1636 1441 1668
rect 1453 1636 1455 1668
rect 1439 1628 1455 1636
rect 1459 1628 1465 1668
rect 1469 1648 1471 1668
rect 1483 1648 1485 1668
rect 1489 1648 1491 1668
rect 1469 1628 1481 1648
rect 1543 1628 1545 1668
rect 1549 1628 1555 1668
rect 1559 1636 1561 1668
rect 1573 1636 1575 1668
rect 1559 1628 1575 1636
rect 1579 1628 1585 1668
rect 1589 1648 1591 1668
rect 1603 1648 1605 1668
rect 1609 1648 1611 1668
rect 1589 1628 1601 1648
rect 1663 1628 1665 1668
rect 1669 1628 1675 1668
rect 1679 1636 1681 1668
rect 1693 1636 1695 1668
rect 1679 1628 1695 1636
rect 1699 1628 1705 1668
rect 1709 1648 1711 1668
rect 1723 1648 1725 1668
rect 1729 1648 1731 1668
rect 1709 1628 1721 1648
rect 1769 1636 1771 1676
rect 1775 1656 1779 1676
rect 1791 1656 1793 1676
rect 1797 1656 1803 1676
rect 1807 1656 1809 1676
rect 1821 1656 1823 1676
rect 1827 1656 1831 1676
rect 1835 1656 1837 1676
rect 1875 1656 1877 1676
rect 1881 1656 1885 1676
rect 1897 1656 1899 1676
rect 1903 1656 1909 1676
rect 1913 1656 1915 1676
rect 1927 1656 1931 1676
rect 1935 1656 1941 1676
rect 1945 1656 1947 1676
rect 1959 1656 1961 1676
rect 1775 1636 1788 1656
rect 1951 1636 1961 1656
rect 1965 1636 1967 1676
rect 2009 1648 2011 1668
rect 2015 1648 2017 1668
rect 2029 1648 2031 1668
rect 2019 1628 2031 1648
rect 2035 1628 2041 1668
rect 2045 1636 2047 1668
rect 2059 1636 2061 1668
rect 2045 1628 2061 1636
rect 2065 1628 2071 1668
rect 2075 1628 2077 1668
rect 2129 1656 2131 1676
rect 2135 1656 2137 1676
rect 2189 1636 2191 1676
rect 2195 1646 2197 1676
rect 2209 1646 2211 1676
rect 2195 1636 2211 1646
rect 2215 1636 2217 1676
rect 2229 1636 2231 1676
rect 2235 1664 2251 1676
rect 2235 1636 2237 1664
rect 2249 1636 2251 1664
rect 2255 1636 2257 1676
rect 2309 1656 2311 1676
rect 2315 1656 2317 1676
rect 2329 1656 2331 1676
rect 2335 1656 2337 1676
rect 2403 1636 2405 1676
rect 2409 1636 2411 1676
rect 2423 1636 2425 1676
rect 2429 1648 2431 1676
rect 2443 1648 2445 1676
rect 2429 1636 2445 1648
rect 2449 1636 2451 1676
rect 2501 1636 2503 1676
rect 2507 1636 2509 1676
rect 2521 1656 2525 1676
rect 2529 1656 2531 1676
rect 2569 1656 2571 1676
rect 2575 1656 2577 1676
rect 2589 1656 2591 1676
rect 2595 1656 2597 1676
rect 2671 1636 2673 1676
rect 2677 1636 2683 1676
rect 2687 1636 2689 1676
rect 2731 1636 2733 1676
rect 2737 1636 2743 1676
rect 2747 1636 2749 1676
rect 2823 1628 2825 1668
rect 2829 1628 2835 1668
rect 2839 1636 2841 1668
rect 2853 1636 2855 1668
rect 2839 1628 2855 1636
rect 2859 1628 2865 1668
rect 2869 1648 2871 1668
rect 2883 1648 2885 1668
rect 2889 1648 2891 1668
rect 2869 1628 2881 1648
rect 2966 1618 2968 1676
rect 2954 1616 2968 1618
rect 2972 1616 2976 1676
rect 2980 1616 2984 1676
rect 2988 1616 2990 1676
rect 3043 1636 3045 1676
rect 3049 1636 3051 1676
rect 3093 1636 3095 1676
rect 3099 1656 3101 1676
rect 3113 1656 3115 1676
rect 3119 1656 3125 1676
rect 3129 1656 3133 1676
rect 3145 1656 3147 1676
rect 3151 1656 3157 1676
rect 3161 1656 3163 1676
rect 3175 1656 3179 1676
rect 3183 1656 3185 1676
rect 3223 1656 3225 1676
rect 3229 1656 3233 1676
rect 3237 1656 3239 1676
rect 3251 1656 3253 1676
rect 3257 1656 3263 1676
rect 3267 1656 3269 1676
rect 3281 1656 3285 1676
rect 3099 1636 3109 1656
rect 3272 1636 3285 1656
rect 3289 1636 3291 1676
rect 3351 1636 3353 1676
rect 3357 1636 3363 1676
rect 3367 1636 3369 1676
rect 3423 1636 3425 1676
rect 3429 1636 3431 1676
rect 3443 1636 3445 1676
rect 3449 1648 3451 1676
rect 3463 1648 3465 1676
rect 3449 1636 3465 1648
rect 3469 1636 3471 1676
rect 3512 1636 3514 1676
rect 3518 1636 3522 1676
rect 3526 1636 3528 1676
rect 3540 1636 3542 1676
rect 3546 1636 3550 1676
rect 3554 1636 3556 1676
rect 3643 1636 3645 1676
rect 3649 1636 3651 1676
rect 3663 1636 3665 1676
rect 3669 1648 3671 1676
rect 3683 1648 3685 1676
rect 3669 1636 3685 1648
rect 3689 1636 3691 1676
rect 3743 1656 3745 1676
rect 3749 1656 3751 1676
rect 3803 1656 3805 1676
rect 3809 1656 3811 1676
rect 3823 1656 3825 1676
rect 3829 1656 3831 1676
rect 3883 1636 3885 1676
rect 3889 1664 3905 1676
rect 3889 1636 3891 1664
rect 3903 1636 3905 1664
rect 3909 1636 3911 1676
rect 3923 1636 3925 1676
rect 3929 1646 3931 1676
rect 3943 1646 3945 1676
rect 3929 1636 3945 1646
rect 3949 1636 3951 1676
rect 4003 1656 4005 1676
rect 4009 1656 4011 1676
rect 4053 1636 4055 1676
rect 4059 1656 4061 1676
rect 4073 1656 4075 1676
rect 4079 1656 4085 1676
rect 4089 1656 4093 1676
rect 4105 1656 4107 1676
rect 4111 1656 4117 1676
rect 4121 1656 4123 1676
rect 4135 1656 4139 1676
rect 4143 1656 4145 1676
rect 4183 1656 4185 1676
rect 4189 1656 4193 1676
rect 4197 1656 4199 1676
rect 4211 1656 4213 1676
rect 4217 1656 4223 1676
rect 4227 1656 4229 1676
rect 4241 1656 4245 1676
rect 4059 1636 4069 1656
rect 4232 1636 4245 1656
rect 4249 1636 4251 1676
rect 4303 1628 4305 1668
rect 4309 1628 4315 1668
rect 4319 1636 4321 1668
rect 4333 1636 4335 1668
rect 4319 1628 4335 1636
rect 4339 1628 4345 1668
rect 4349 1648 4351 1668
rect 4363 1648 4365 1668
rect 4369 1648 4371 1668
rect 4349 1628 4361 1648
rect 4423 1628 4425 1668
rect 4429 1628 4435 1668
rect 4439 1636 4441 1668
rect 4453 1636 4455 1668
rect 4439 1628 4455 1636
rect 4459 1628 4465 1668
rect 4469 1648 4471 1668
rect 4483 1648 4485 1668
rect 4489 1648 4491 1668
rect 4529 1648 4531 1668
rect 4535 1648 4537 1668
rect 4549 1648 4551 1668
rect 4469 1628 4481 1648
rect 4539 1628 4551 1648
rect 4555 1628 4561 1668
rect 4565 1636 4567 1668
rect 4579 1636 4581 1668
rect 4565 1628 4581 1636
rect 4585 1628 4591 1668
rect 4595 1628 4597 1668
rect 4649 1648 4651 1668
rect 4655 1648 4657 1668
rect 4669 1648 4671 1668
rect 4659 1628 4671 1648
rect 4675 1628 4681 1668
rect 4685 1636 4687 1668
rect 4699 1636 4701 1668
rect 4685 1628 4701 1636
rect 4705 1628 4711 1668
rect 4715 1628 4717 1668
rect 4769 1648 4771 1668
rect 4775 1648 4777 1668
rect 4789 1648 4791 1668
rect 4779 1628 4791 1648
rect 4795 1628 4801 1668
rect 4805 1636 4807 1668
rect 4819 1636 4821 1668
rect 4805 1628 4821 1636
rect 4825 1628 4831 1668
rect 4835 1628 4837 1668
rect 4889 1648 4891 1668
rect 4895 1648 4897 1668
rect 4909 1648 4911 1668
rect 4899 1628 4911 1648
rect 4915 1628 4921 1668
rect 4925 1636 4927 1668
rect 4939 1636 4941 1668
rect 4925 1628 4941 1636
rect 4945 1628 4951 1668
rect 4955 1628 4957 1668
rect 5009 1636 5011 1676
rect 5015 1656 5019 1676
rect 5031 1656 5033 1676
rect 5037 1656 5043 1676
rect 5047 1656 5049 1676
rect 5061 1656 5063 1676
rect 5067 1656 5071 1676
rect 5075 1656 5077 1676
rect 5115 1656 5117 1676
rect 5121 1656 5125 1676
rect 5137 1656 5139 1676
rect 5143 1656 5149 1676
rect 5153 1656 5155 1676
rect 5167 1656 5171 1676
rect 5175 1656 5181 1676
rect 5185 1656 5187 1676
rect 5199 1656 5201 1676
rect 5015 1636 5028 1656
rect 5191 1636 5201 1656
rect 5205 1636 5207 1676
rect 5249 1636 5251 1676
rect 5255 1656 5259 1676
rect 5271 1656 5273 1676
rect 5277 1656 5283 1676
rect 5287 1656 5289 1676
rect 5301 1656 5303 1676
rect 5307 1656 5311 1676
rect 5315 1656 5317 1676
rect 5355 1656 5357 1676
rect 5361 1656 5365 1676
rect 5377 1656 5379 1676
rect 5383 1656 5389 1676
rect 5393 1656 5395 1676
rect 5407 1656 5411 1676
rect 5415 1656 5421 1676
rect 5425 1656 5427 1676
rect 5439 1656 5441 1676
rect 5255 1636 5268 1656
rect 5431 1636 5441 1656
rect 5445 1636 5447 1676
rect 5492 1636 5494 1676
rect 5498 1636 5502 1676
rect 5506 1636 5508 1676
rect 5520 1636 5522 1676
rect 5526 1636 5530 1676
rect 5534 1636 5536 1676
rect 5609 1648 5611 1668
rect 5615 1648 5617 1668
rect 5629 1648 5631 1668
rect 5619 1628 5631 1648
rect 5635 1628 5641 1668
rect 5645 1636 5647 1668
rect 5659 1636 5661 1668
rect 5645 1628 5661 1636
rect 5665 1628 5671 1668
rect 5675 1628 5677 1668
rect 5743 1636 5745 1676
rect 5749 1636 5751 1676
rect 5763 1636 5765 1676
rect 5769 1648 5771 1676
rect 5783 1648 5785 1676
rect 5769 1636 5785 1648
rect 5789 1636 5791 1676
rect 5843 1656 5845 1676
rect 5849 1656 5851 1676
rect 5863 1656 5865 1676
rect 5869 1656 5871 1676
rect 5931 1636 5933 1676
rect 5937 1636 5943 1676
rect 5947 1636 5949 1676
rect 6003 1636 6005 1676
rect 6009 1636 6011 1676
rect 6023 1636 6025 1676
rect 6029 1648 6031 1676
rect 6043 1648 6045 1676
rect 6029 1636 6045 1648
rect 6049 1636 6051 1676
rect 6103 1656 6105 1676
rect 6109 1656 6111 1676
rect 6123 1656 6125 1676
rect 6129 1656 6131 1676
rect 6183 1636 6185 1676
rect 6189 1664 6205 1676
rect 6189 1636 6191 1664
rect 6203 1636 6205 1664
rect 6209 1636 6211 1676
rect 6223 1636 6225 1676
rect 6229 1646 6231 1676
rect 6243 1646 6245 1676
rect 6229 1636 6245 1646
rect 6249 1636 6251 1676
rect 6303 1628 6305 1668
rect 6309 1628 6315 1668
rect 6319 1636 6321 1668
rect 6333 1636 6335 1668
rect 6319 1628 6335 1636
rect 6339 1628 6345 1668
rect 6349 1648 6351 1668
rect 6363 1648 6365 1668
rect 6369 1648 6371 1668
rect 6409 1656 6411 1676
rect 6415 1656 6417 1676
rect 6349 1628 6361 1648
rect 6469 1636 6471 1676
rect 6475 1656 6479 1676
rect 6491 1656 6493 1676
rect 6497 1656 6503 1676
rect 6507 1656 6509 1676
rect 6521 1656 6523 1676
rect 6527 1656 6531 1676
rect 6535 1656 6537 1676
rect 6575 1656 6577 1676
rect 6581 1656 6585 1676
rect 6597 1656 6599 1676
rect 6603 1656 6609 1676
rect 6613 1656 6615 1676
rect 6627 1656 6631 1676
rect 6635 1656 6641 1676
rect 6645 1656 6647 1676
rect 6659 1656 6661 1676
rect 6475 1636 6488 1656
rect 6651 1636 6661 1656
rect 6665 1636 6667 1676
rect 29 1224 31 1264
rect 35 1224 41 1264
rect 45 1224 47 1264
rect 59 1224 61 1264
rect 65 1224 67 1264
rect 129 1224 131 1244
rect 135 1224 137 1244
rect 149 1224 151 1244
rect 155 1224 157 1244
rect 223 1224 225 1264
rect 229 1224 231 1264
rect 243 1224 245 1264
rect 249 1252 265 1264
rect 249 1224 251 1252
rect 263 1224 265 1252
rect 269 1224 271 1264
rect 323 1224 325 1244
rect 329 1224 331 1244
rect 343 1224 345 1244
rect 349 1224 351 1244
rect 389 1224 391 1244
rect 395 1224 397 1244
rect 449 1224 451 1244
rect 455 1224 457 1244
rect 531 1224 533 1264
rect 537 1224 543 1264
rect 547 1224 549 1264
rect 592 1224 594 1264
rect 598 1224 602 1264
rect 606 1224 608 1264
rect 620 1224 624 1244
rect 628 1224 630 1244
rect 693 1224 695 1264
rect 699 1244 709 1264
rect 872 1244 885 1264
rect 699 1224 701 1244
rect 713 1224 715 1244
rect 719 1224 725 1244
rect 729 1224 733 1244
rect 745 1224 747 1244
rect 751 1224 757 1244
rect 761 1224 763 1244
rect 775 1224 779 1244
rect 783 1224 785 1244
rect 823 1224 825 1244
rect 829 1224 833 1244
rect 837 1224 839 1244
rect 851 1224 853 1244
rect 857 1224 863 1244
rect 867 1224 869 1244
rect 881 1224 885 1244
rect 889 1224 891 1264
rect 951 1224 953 1264
rect 957 1224 963 1264
rect 967 1224 969 1264
rect 1010 1224 1012 1284
rect 1016 1224 1020 1284
rect 1024 1224 1028 1284
rect 1032 1282 1046 1284
rect 1032 1224 1034 1282
rect 1109 1224 1111 1244
rect 1115 1224 1117 1244
rect 1129 1224 1131 1244
rect 1135 1224 1137 1244
rect 1193 1224 1195 1264
rect 1199 1244 1209 1264
rect 1372 1244 1385 1264
rect 1199 1224 1201 1244
rect 1213 1224 1215 1244
rect 1219 1224 1225 1244
rect 1229 1224 1233 1244
rect 1245 1224 1247 1244
rect 1251 1224 1257 1244
rect 1261 1224 1263 1244
rect 1275 1224 1279 1244
rect 1283 1224 1285 1244
rect 1323 1224 1325 1244
rect 1329 1224 1333 1244
rect 1337 1224 1339 1244
rect 1351 1224 1353 1244
rect 1357 1224 1363 1244
rect 1367 1224 1369 1244
rect 1381 1224 1385 1244
rect 1389 1224 1391 1264
rect 1443 1224 1445 1264
rect 1449 1224 1451 1264
rect 1463 1224 1465 1264
rect 1469 1224 1471 1264
rect 1483 1224 1485 1264
rect 1489 1224 1491 1264
rect 1503 1224 1505 1264
rect 1509 1224 1511 1264
rect 1523 1224 1525 1264
rect 1529 1224 1531 1264
rect 1543 1224 1545 1264
rect 1549 1224 1551 1264
rect 1563 1224 1565 1264
rect 1569 1224 1571 1264
rect 1583 1224 1585 1264
rect 1589 1224 1591 1264
rect 1643 1232 1645 1272
rect 1649 1232 1655 1272
rect 1659 1264 1675 1272
rect 1659 1232 1661 1264
rect 1673 1232 1675 1264
rect 1679 1232 1685 1272
rect 1689 1252 1701 1272
rect 1689 1232 1691 1252
rect 1703 1232 1705 1252
rect 1709 1232 1711 1252
rect 1763 1224 1765 1244
rect 1769 1224 1771 1244
rect 1783 1224 1785 1244
rect 1789 1224 1791 1244
rect 1843 1224 1845 1264
rect 1849 1236 1851 1264
rect 1863 1236 1865 1264
rect 1849 1224 1865 1236
rect 1869 1224 1871 1264
rect 1883 1224 1885 1264
rect 1889 1254 1905 1264
rect 1889 1224 1891 1254
rect 1903 1224 1905 1254
rect 1909 1224 1911 1264
rect 1963 1224 1965 1264
rect 1969 1224 1971 1264
rect 1983 1224 1985 1264
rect 1989 1252 2005 1264
rect 1989 1224 1991 1252
rect 2003 1224 2005 1252
rect 2009 1224 2011 1264
rect 2049 1224 2051 1244
rect 2055 1224 2057 1244
rect 2109 1224 2111 1264
rect 2115 1252 2131 1264
rect 2115 1224 2117 1252
rect 2129 1224 2131 1252
rect 2135 1224 2137 1264
rect 2149 1224 2151 1264
rect 2155 1224 2157 1264
rect 2211 1224 2213 1264
rect 2217 1224 2223 1264
rect 2227 1224 2229 1264
rect 2299 1252 2311 1272
rect 2289 1232 2291 1252
rect 2295 1232 2297 1252
rect 2309 1232 2311 1252
rect 2315 1232 2321 1272
rect 2325 1264 2341 1272
rect 2325 1232 2327 1264
rect 2339 1232 2341 1264
rect 2345 1232 2351 1272
rect 2355 1232 2357 1272
rect 2423 1232 2425 1272
rect 2429 1232 2435 1272
rect 2439 1264 2455 1272
rect 2439 1232 2441 1264
rect 2453 1232 2455 1264
rect 2459 1232 2465 1272
rect 2469 1252 2481 1272
rect 2469 1232 2471 1252
rect 2483 1232 2485 1252
rect 2489 1232 2491 1252
rect 2564 1224 2566 1264
rect 2570 1224 2574 1264
rect 2578 1224 2580 1264
rect 2592 1224 2594 1264
rect 2598 1224 2602 1264
rect 2606 1224 2608 1264
rect 2652 1224 2654 1264
rect 2658 1224 2662 1264
rect 2666 1224 2668 1264
rect 2680 1224 2682 1264
rect 2686 1224 2690 1264
rect 2694 1224 2696 1264
rect 2804 1224 2806 1264
rect 2810 1224 2814 1264
rect 2818 1224 2820 1264
rect 2832 1224 2834 1264
rect 2838 1224 2842 1264
rect 2846 1224 2848 1264
rect 2889 1224 2891 1244
rect 2895 1224 2899 1244
rect 2911 1224 2913 1264
rect 2917 1224 2919 1264
rect 3004 1224 3006 1264
rect 3010 1224 3014 1264
rect 3018 1224 3020 1264
rect 3032 1224 3034 1264
rect 3038 1224 3042 1264
rect 3046 1224 3048 1264
rect 3103 1224 3105 1244
rect 3109 1224 3111 1244
rect 3163 1232 3165 1272
rect 3169 1232 3175 1272
rect 3179 1264 3195 1272
rect 3179 1232 3181 1264
rect 3193 1232 3195 1264
rect 3199 1232 3205 1272
rect 3209 1252 3221 1272
rect 3209 1232 3211 1252
rect 3223 1232 3225 1252
rect 3229 1232 3231 1252
rect 3273 1224 3275 1264
rect 3279 1244 3289 1264
rect 3452 1244 3465 1264
rect 3279 1224 3281 1244
rect 3293 1224 3295 1244
rect 3299 1224 3305 1244
rect 3309 1224 3313 1244
rect 3325 1224 3327 1244
rect 3331 1224 3337 1244
rect 3341 1224 3343 1244
rect 3355 1224 3359 1244
rect 3363 1224 3365 1244
rect 3403 1224 3405 1244
rect 3409 1224 3413 1244
rect 3417 1224 3419 1244
rect 3431 1224 3433 1244
rect 3437 1224 3443 1244
rect 3447 1224 3449 1244
rect 3461 1224 3465 1244
rect 3469 1224 3471 1264
rect 3523 1224 3525 1244
rect 3529 1224 3531 1244
rect 3543 1224 3545 1244
rect 3549 1224 3551 1244
rect 3603 1224 3605 1264
rect 3609 1236 3611 1264
rect 3623 1236 3625 1264
rect 3609 1224 3625 1236
rect 3629 1224 3631 1264
rect 3643 1224 3645 1264
rect 3649 1254 3665 1264
rect 3649 1224 3651 1254
rect 3663 1224 3665 1254
rect 3669 1224 3671 1264
rect 3723 1224 3725 1264
rect 3729 1224 3731 1264
rect 3743 1224 3745 1264
rect 3749 1252 3765 1264
rect 3749 1224 3751 1252
rect 3763 1224 3765 1252
rect 3769 1224 3771 1264
rect 3823 1224 3825 1244
rect 3829 1224 3831 1244
rect 3869 1224 3871 1264
rect 3875 1244 3888 1264
rect 4051 1244 4061 1264
rect 3875 1224 3879 1244
rect 3891 1224 3893 1244
rect 3897 1224 3903 1244
rect 3907 1224 3909 1244
rect 3921 1224 3923 1244
rect 3927 1224 3931 1244
rect 3935 1224 3937 1244
rect 3975 1224 3977 1244
rect 3981 1224 3985 1244
rect 3997 1224 3999 1244
rect 4003 1224 4009 1244
rect 4013 1224 4015 1244
rect 4027 1224 4031 1244
rect 4035 1224 4041 1244
rect 4045 1224 4047 1244
rect 4059 1224 4061 1244
rect 4065 1224 4067 1264
rect 4109 1224 4111 1264
rect 4115 1244 4128 1264
rect 4291 1244 4301 1264
rect 4115 1224 4119 1244
rect 4131 1224 4133 1244
rect 4137 1224 4143 1244
rect 4147 1224 4149 1244
rect 4161 1224 4163 1244
rect 4167 1224 4171 1244
rect 4175 1224 4177 1244
rect 4215 1224 4217 1244
rect 4221 1224 4225 1244
rect 4237 1224 4239 1244
rect 4243 1224 4249 1244
rect 4253 1224 4255 1244
rect 4267 1224 4271 1244
rect 4275 1224 4281 1244
rect 4285 1224 4287 1244
rect 4299 1224 4301 1244
rect 4305 1224 4307 1264
rect 4363 1224 4365 1244
rect 4369 1224 4371 1244
rect 4412 1224 4414 1264
rect 4418 1224 4422 1264
rect 4426 1224 4428 1264
rect 4440 1224 4442 1264
rect 4446 1224 4450 1264
rect 4454 1224 4456 1264
rect 4539 1252 4551 1272
rect 4529 1232 4531 1252
rect 4535 1232 4537 1252
rect 4549 1232 4551 1252
rect 4555 1232 4561 1272
rect 4565 1264 4581 1272
rect 4565 1232 4567 1264
rect 4579 1232 4581 1264
rect 4585 1232 4591 1272
rect 4595 1232 4597 1272
rect 4684 1224 4686 1264
rect 4690 1224 4694 1264
rect 4698 1224 4700 1264
rect 4712 1224 4714 1264
rect 4718 1224 4722 1264
rect 4726 1224 4728 1264
rect 4781 1224 4783 1264
rect 4787 1224 4789 1264
rect 4801 1224 4805 1244
rect 4809 1224 4811 1244
rect 4871 1224 4873 1264
rect 4877 1224 4883 1264
rect 4887 1224 4889 1264
rect 4951 1224 4953 1264
rect 4957 1224 4963 1264
rect 4967 1224 4969 1264
rect 5023 1224 5025 1264
rect 5029 1236 5031 1264
rect 5043 1236 5045 1264
rect 5029 1224 5045 1236
rect 5049 1224 5051 1264
rect 5063 1224 5065 1264
rect 5069 1254 5085 1264
rect 5069 1224 5071 1254
rect 5083 1224 5085 1254
rect 5089 1224 5091 1264
rect 5143 1224 5145 1264
rect 5149 1236 5151 1264
rect 5163 1236 5165 1264
rect 5149 1224 5165 1236
rect 5169 1224 5171 1264
rect 5183 1224 5185 1264
rect 5189 1254 5205 1264
rect 5189 1224 5191 1254
rect 5203 1224 5205 1254
rect 5209 1224 5211 1264
rect 5249 1224 5251 1264
rect 5255 1224 5257 1264
rect 5331 1224 5333 1264
rect 5337 1224 5343 1264
rect 5347 1224 5349 1264
rect 5389 1224 5391 1264
rect 5395 1254 5411 1264
rect 5395 1224 5397 1254
rect 5409 1224 5411 1254
rect 5415 1224 5417 1264
rect 5429 1224 5431 1264
rect 5435 1236 5437 1264
rect 5449 1236 5451 1264
rect 5435 1224 5451 1236
rect 5455 1224 5457 1264
rect 5530 1224 5532 1244
rect 5536 1224 5540 1244
rect 5552 1224 5554 1264
rect 5558 1224 5562 1264
rect 5566 1224 5568 1264
rect 5609 1224 5611 1264
rect 5615 1224 5617 1264
rect 5679 1252 5691 1272
rect 5669 1232 5671 1252
rect 5675 1232 5677 1252
rect 5689 1232 5691 1252
rect 5695 1232 5701 1272
rect 5705 1264 5721 1272
rect 5705 1232 5707 1264
rect 5719 1232 5721 1264
rect 5725 1232 5731 1272
rect 5735 1232 5737 1272
rect 5811 1224 5813 1264
rect 5817 1224 5823 1264
rect 5827 1224 5829 1264
rect 5883 1224 5885 1264
rect 5889 1224 5891 1264
rect 5903 1224 5905 1264
rect 5909 1252 5925 1264
rect 5909 1224 5911 1252
rect 5923 1224 5925 1252
rect 5929 1224 5931 1264
rect 5983 1224 5985 1244
rect 5989 1224 5991 1244
rect 6029 1224 6031 1264
rect 6035 1252 6051 1264
rect 6035 1224 6037 1252
rect 6049 1224 6051 1252
rect 6055 1224 6057 1264
rect 6069 1224 6071 1264
rect 6075 1224 6077 1264
rect 6129 1224 6131 1264
rect 6135 1254 6151 1264
rect 6135 1224 6137 1254
rect 6149 1224 6151 1254
rect 6155 1224 6157 1264
rect 6169 1224 6171 1264
rect 6175 1236 6177 1264
rect 6189 1236 6191 1264
rect 6175 1224 6191 1236
rect 6195 1224 6197 1264
rect 6249 1224 6251 1264
rect 6255 1244 6268 1264
rect 6431 1244 6441 1264
rect 6255 1224 6259 1244
rect 6271 1224 6273 1244
rect 6277 1224 6283 1244
rect 6287 1224 6289 1244
rect 6301 1224 6303 1244
rect 6307 1224 6311 1244
rect 6315 1224 6317 1244
rect 6355 1224 6357 1244
rect 6361 1224 6365 1244
rect 6377 1224 6379 1244
rect 6383 1224 6389 1244
rect 6393 1224 6395 1244
rect 6407 1224 6411 1244
rect 6415 1224 6421 1244
rect 6425 1224 6427 1244
rect 6439 1224 6441 1244
rect 6445 1224 6447 1264
rect 6489 1224 6491 1264
rect 6495 1244 6508 1264
rect 6671 1244 6681 1264
rect 6495 1224 6499 1244
rect 6511 1224 6513 1244
rect 6517 1224 6523 1244
rect 6527 1224 6529 1244
rect 6541 1224 6543 1244
rect 6547 1224 6551 1244
rect 6555 1224 6557 1244
rect 6595 1224 6597 1244
rect 6601 1224 6605 1244
rect 6617 1224 6619 1244
rect 6623 1224 6629 1244
rect 6633 1224 6635 1244
rect 6647 1224 6651 1244
rect 6655 1224 6661 1244
rect 6665 1224 6667 1244
rect 6679 1224 6681 1244
rect 6685 1224 6687 1264
rect 29 1156 31 1196
rect 35 1176 39 1196
rect 51 1176 53 1196
rect 57 1176 63 1196
rect 67 1176 69 1196
rect 81 1176 83 1196
rect 87 1176 91 1196
rect 95 1176 97 1196
rect 135 1176 137 1196
rect 141 1176 145 1196
rect 157 1176 159 1196
rect 163 1176 169 1196
rect 173 1176 175 1196
rect 187 1176 191 1196
rect 195 1176 201 1196
rect 205 1176 207 1196
rect 219 1176 221 1196
rect 35 1156 48 1176
rect 211 1156 221 1176
rect 225 1156 227 1196
rect 283 1176 285 1196
rect 289 1176 291 1196
rect 329 1156 331 1196
rect 335 1176 339 1196
rect 351 1176 353 1196
rect 357 1176 363 1196
rect 367 1176 369 1196
rect 381 1176 383 1196
rect 387 1176 391 1196
rect 395 1176 397 1196
rect 435 1176 437 1196
rect 441 1176 445 1196
rect 457 1176 459 1196
rect 463 1176 469 1196
rect 473 1176 475 1196
rect 487 1176 491 1196
rect 495 1176 501 1196
rect 505 1176 507 1196
rect 519 1176 521 1196
rect 335 1156 348 1176
rect 511 1156 521 1176
rect 525 1156 527 1196
rect 569 1176 571 1196
rect 575 1176 577 1196
rect 630 1136 632 1196
rect 636 1136 640 1196
rect 644 1136 648 1196
rect 652 1138 654 1196
rect 729 1176 731 1196
rect 735 1176 737 1196
rect 749 1176 751 1196
rect 755 1176 757 1196
rect 652 1136 666 1138
rect 810 1136 812 1196
rect 816 1136 820 1196
rect 824 1136 828 1196
rect 832 1138 834 1196
rect 911 1156 913 1196
rect 917 1156 923 1196
rect 927 1156 929 1196
rect 989 1176 991 1196
rect 995 1176 997 1196
rect 832 1136 846 1138
rect 1053 1156 1055 1196
rect 1059 1176 1061 1196
rect 1073 1176 1075 1196
rect 1079 1176 1085 1196
rect 1089 1176 1093 1196
rect 1105 1176 1107 1196
rect 1111 1176 1117 1196
rect 1121 1176 1123 1196
rect 1135 1176 1139 1196
rect 1143 1176 1145 1196
rect 1183 1176 1185 1196
rect 1189 1176 1193 1196
rect 1197 1176 1199 1196
rect 1211 1176 1213 1196
rect 1217 1176 1223 1196
rect 1227 1176 1229 1196
rect 1241 1176 1245 1196
rect 1059 1156 1069 1176
rect 1232 1156 1245 1176
rect 1249 1156 1251 1196
rect 1289 1156 1291 1196
rect 1295 1156 1297 1196
rect 1309 1156 1311 1196
rect 1315 1156 1317 1196
rect 1329 1156 1331 1196
rect 1335 1156 1337 1196
rect 1349 1156 1351 1196
rect 1355 1156 1357 1196
rect 1369 1156 1371 1196
rect 1375 1156 1377 1196
rect 1389 1156 1391 1196
rect 1395 1156 1397 1196
rect 1409 1156 1411 1196
rect 1415 1156 1417 1196
rect 1429 1156 1431 1196
rect 1435 1156 1437 1196
rect 1493 1156 1495 1196
rect 1499 1176 1501 1196
rect 1513 1176 1515 1196
rect 1519 1176 1525 1196
rect 1529 1176 1533 1196
rect 1545 1176 1547 1196
rect 1551 1176 1557 1196
rect 1561 1176 1563 1196
rect 1575 1176 1579 1196
rect 1583 1176 1585 1196
rect 1623 1176 1625 1196
rect 1629 1176 1633 1196
rect 1637 1176 1639 1196
rect 1651 1176 1653 1196
rect 1657 1176 1663 1196
rect 1667 1176 1669 1196
rect 1681 1176 1685 1196
rect 1499 1156 1509 1176
rect 1672 1156 1685 1176
rect 1689 1156 1691 1196
rect 1743 1176 1745 1196
rect 1749 1176 1751 1196
rect 1763 1176 1765 1196
rect 1769 1176 1771 1196
rect 1823 1156 1825 1196
rect 1829 1184 1845 1196
rect 1829 1156 1831 1184
rect 1843 1156 1845 1184
rect 1849 1156 1851 1196
rect 1863 1156 1865 1196
rect 1869 1166 1871 1196
rect 1883 1166 1885 1196
rect 1869 1156 1885 1166
rect 1889 1156 1891 1196
rect 1943 1156 1945 1196
rect 1949 1156 1951 1196
rect 1963 1156 1965 1196
rect 1969 1168 1971 1196
rect 1983 1168 1985 1196
rect 1969 1156 1985 1168
rect 1989 1156 1991 1196
rect 2043 1156 2045 1196
rect 2049 1156 2051 1196
rect 2063 1156 2065 1196
rect 2069 1168 2071 1196
rect 2083 1168 2085 1196
rect 2069 1156 2085 1168
rect 2089 1156 2091 1196
rect 2143 1176 2145 1196
rect 2149 1176 2151 1196
rect 2163 1176 2165 1196
rect 2169 1176 2171 1196
rect 2223 1156 2225 1196
rect 2229 1184 2245 1196
rect 2229 1156 2231 1184
rect 2243 1156 2245 1184
rect 2249 1156 2251 1196
rect 2263 1156 2265 1196
rect 2269 1166 2271 1196
rect 2283 1166 2285 1196
rect 2269 1156 2285 1166
rect 2289 1156 2291 1196
rect 2333 1156 2335 1196
rect 2339 1176 2341 1196
rect 2353 1176 2355 1196
rect 2359 1176 2365 1196
rect 2369 1176 2373 1196
rect 2385 1176 2387 1196
rect 2391 1176 2397 1196
rect 2401 1176 2403 1196
rect 2415 1176 2419 1196
rect 2423 1176 2425 1196
rect 2463 1176 2465 1196
rect 2469 1176 2473 1196
rect 2477 1176 2479 1196
rect 2491 1176 2493 1196
rect 2497 1176 2503 1196
rect 2507 1176 2509 1196
rect 2521 1176 2525 1196
rect 2339 1156 2349 1176
rect 2512 1156 2525 1176
rect 2529 1156 2531 1196
rect 2583 1176 2585 1196
rect 2589 1176 2591 1196
rect 2629 1156 2631 1196
rect 2635 1168 2637 1196
rect 2649 1168 2651 1196
rect 2635 1156 2651 1168
rect 2655 1156 2657 1196
rect 2669 1156 2671 1196
rect 2675 1156 2677 1196
rect 2741 1156 2743 1196
rect 2747 1156 2749 1196
rect 2761 1176 2765 1196
rect 2769 1176 2771 1196
rect 2809 1176 2811 1196
rect 2815 1176 2817 1196
rect 2904 1156 2906 1196
rect 2910 1156 2914 1196
rect 2918 1156 2920 1196
rect 2932 1156 2934 1196
rect 2938 1156 2942 1196
rect 2946 1156 2948 1196
rect 2993 1156 2995 1196
rect 2999 1176 3001 1196
rect 3013 1176 3015 1196
rect 3019 1176 3025 1196
rect 3029 1176 3033 1196
rect 3045 1176 3047 1196
rect 3051 1176 3057 1196
rect 3061 1176 3063 1196
rect 3075 1176 3079 1196
rect 3083 1176 3085 1196
rect 3123 1176 3125 1196
rect 3129 1176 3133 1196
rect 3137 1176 3139 1196
rect 3151 1176 3153 1196
rect 3157 1176 3163 1196
rect 3167 1176 3169 1196
rect 3181 1176 3185 1196
rect 2999 1156 3009 1176
rect 3172 1156 3185 1176
rect 3189 1156 3191 1196
rect 3231 1156 3233 1196
rect 3237 1156 3243 1196
rect 3247 1156 3249 1196
rect 3323 1148 3325 1188
rect 3329 1148 3335 1188
rect 3339 1156 3341 1188
rect 3353 1156 3355 1188
rect 3339 1148 3355 1156
rect 3359 1148 3365 1188
rect 3369 1168 3371 1188
rect 3383 1168 3385 1188
rect 3389 1168 3391 1188
rect 3429 1168 3431 1188
rect 3435 1168 3437 1188
rect 3449 1168 3451 1188
rect 3369 1148 3381 1168
rect 3439 1148 3451 1168
rect 3455 1148 3461 1188
rect 3465 1156 3467 1188
rect 3479 1156 3481 1188
rect 3465 1148 3481 1156
rect 3485 1148 3491 1188
rect 3495 1148 3497 1188
rect 3561 1156 3563 1196
rect 3567 1156 3569 1196
rect 3581 1176 3585 1196
rect 3589 1176 3591 1196
rect 3633 1156 3635 1196
rect 3639 1176 3641 1196
rect 3653 1176 3655 1196
rect 3659 1176 3665 1196
rect 3669 1176 3673 1196
rect 3685 1176 3687 1196
rect 3691 1176 3697 1196
rect 3701 1176 3703 1196
rect 3715 1176 3719 1196
rect 3723 1176 3725 1196
rect 3763 1176 3765 1196
rect 3769 1176 3773 1196
rect 3777 1176 3779 1196
rect 3791 1176 3793 1196
rect 3797 1176 3803 1196
rect 3807 1176 3809 1196
rect 3821 1176 3825 1196
rect 3639 1156 3649 1176
rect 3812 1156 3825 1176
rect 3829 1156 3831 1196
rect 3869 1168 3871 1188
rect 3875 1168 3877 1188
rect 3889 1168 3891 1188
rect 3879 1148 3891 1168
rect 3895 1148 3901 1188
rect 3905 1156 3907 1188
rect 3919 1156 3921 1188
rect 3905 1148 3921 1156
rect 3925 1148 3931 1188
rect 3935 1148 3937 1188
rect 4003 1148 4005 1188
rect 4009 1148 4015 1188
rect 4019 1156 4021 1188
rect 4033 1156 4035 1188
rect 4019 1148 4035 1156
rect 4039 1148 4045 1188
rect 4049 1168 4051 1188
rect 4063 1168 4065 1188
rect 4069 1168 4071 1188
rect 4109 1176 4111 1196
rect 4115 1176 4117 1196
rect 4049 1148 4061 1168
rect 4169 1156 4171 1196
rect 4175 1166 4177 1196
rect 4189 1166 4191 1196
rect 4175 1156 4191 1166
rect 4195 1156 4197 1196
rect 4209 1156 4211 1196
rect 4215 1184 4231 1196
rect 4215 1156 4217 1184
rect 4229 1156 4231 1184
rect 4235 1156 4237 1196
rect 4289 1176 4291 1196
rect 4295 1176 4297 1196
rect 4309 1176 4311 1196
rect 4315 1176 4317 1196
rect 4383 1156 4385 1196
rect 4389 1156 4391 1196
rect 4403 1156 4405 1196
rect 4409 1168 4411 1196
rect 4423 1168 4425 1196
rect 4409 1156 4425 1168
rect 4429 1156 4431 1196
rect 4490 1176 4492 1196
rect 4496 1176 4500 1196
rect 4512 1156 4514 1196
rect 4518 1156 4522 1196
rect 4526 1156 4528 1196
rect 4573 1156 4575 1196
rect 4579 1176 4581 1196
rect 4593 1176 4595 1196
rect 4599 1176 4605 1196
rect 4609 1176 4613 1196
rect 4625 1176 4627 1196
rect 4631 1176 4637 1196
rect 4641 1176 4643 1196
rect 4655 1176 4659 1196
rect 4663 1176 4665 1196
rect 4703 1176 4705 1196
rect 4709 1176 4713 1196
rect 4717 1176 4719 1196
rect 4731 1176 4733 1196
rect 4737 1176 4743 1196
rect 4747 1176 4749 1196
rect 4761 1176 4765 1196
rect 4579 1156 4589 1176
rect 4752 1156 4765 1176
rect 4769 1156 4771 1196
rect 4809 1156 4811 1196
rect 4815 1166 4817 1196
rect 4829 1166 4831 1196
rect 4815 1156 4831 1166
rect 4835 1156 4837 1196
rect 4849 1156 4851 1196
rect 4855 1184 4871 1196
rect 4855 1156 4857 1184
rect 4869 1156 4871 1184
rect 4875 1156 4877 1196
rect 4943 1176 4945 1196
rect 4949 1176 4951 1196
rect 4963 1176 4965 1196
rect 4969 1176 4971 1196
rect 5023 1156 5025 1196
rect 5029 1156 5031 1196
rect 5043 1156 5045 1196
rect 5049 1168 5051 1196
rect 5063 1168 5065 1196
rect 5049 1156 5065 1168
rect 5069 1156 5071 1196
rect 5123 1176 5125 1196
rect 5129 1176 5131 1196
rect 5143 1176 5145 1196
rect 5149 1176 5151 1196
rect 5189 1176 5191 1196
rect 5195 1176 5197 1196
rect 5209 1176 5211 1196
rect 5215 1176 5217 1196
rect 5269 1176 5271 1196
rect 5275 1176 5277 1196
rect 5289 1176 5291 1196
rect 5295 1176 5297 1196
rect 5361 1156 5363 1196
rect 5367 1156 5369 1196
rect 5381 1176 5385 1196
rect 5389 1176 5391 1196
rect 5429 1176 5431 1196
rect 5435 1176 5437 1196
rect 5449 1176 5451 1196
rect 5455 1176 5457 1196
rect 5509 1176 5511 1196
rect 5515 1176 5517 1196
rect 5529 1176 5531 1196
rect 5535 1176 5537 1196
rect 5592 1156 5594 1196
rect 5598 1156 5602 1196
rect 5606 1156 5608 1196
rect 5620 1176 5624 1196
rect 5628 1176 5630 1196
rect 5689 1176 5691 1196
rect 5695 1176 5697 1196
rect 5709 1176 5711 1196
rect 5715 1176 5717 1196
rect 5729 1176 5731 1196
rect 5719 1156 5731 1176
rect 5735 1156 5737 1196
rect 5803 1176 5805 1196
rect 5809 1176 5811 1196
rect 5823 1176 5825 1196
rect 5829 1176 5831 1196
rect 5869 1156 5871 1196
rect 5875 1168 5877 1196
rect 5889 1168 5891 1196
rect 5875 1156 5891 1168
rect 5895 1156 5897 1196
rect 5909 1156 5911 1196
rect 5915 1156 5917 1196
rect 6006 1138 6008 1196
rect 5994 1136 6008 1138
rect 6012 1136 6016 1196
rect 6020 1136 6024 1196
rect 6028 1136 6030 1196
rect 6069 1156 6071 1196
rect 6075 1168 6077 1196
rect 6089 1168 6091 1196
rect 6075 1156 6091 1168
rect 6095 1156 6097 1196
rect 6109 1156 6111 1196
rect 6115 1156 6117 1196
rect 6183 1176 6185 1196
rect 6189 1176 6191 1196
rect 6203 1176 6205 1196
rect 6209 1176 6211 1196
rect 6249 1176 6251 1196
rect 6255 1176 6257 1196
rect 6269 1176 6271 1196
rect 6275 1176 6277 1196
rect 6329 1156 6331 1196
rect 6335 1176 6339 1196
rect 6351 1176 6353 1196
rect 6357 1176 6363 1196
rect 6367 1176 6369 1196
rect 6381 1176 6383 1196
rect 6387 1176 6391 1196
rect 6395 1176 6397 1196
rect 6435 1176 6437 1196
rect 6441 1176 6445 1196
rect 6457 1176 6459 1196
rect 6463 1176 6469 1196
rect 6473 1176 6475 1196
rect 6487 1176 6491 1196
rect 6495 1176 6501 1196
rect 6505 1176 6507 1196
rect 6519 1176 6521 1196
rect 6335 1156 6348 1176
rect 6511 1156 6521 1176
rect 6525 1156 6527 1196
rect 6569 1156 6571 1196
rect 6575 1166 6577 1196
rect 6589 1166 6591 1196
rect 6575 1156 6591 1166
rect 6595 1156 6597 1196
rect 6609 1156 6611 1196
rect 6615 1184 6631 1196
rect 6615 1156 6617 1184
rect 6629 1156 6631 1184
rect 6635 1156 6637 1196
rect 59 764 71 784
rect 29 744 31 764
rect 35 744 37 764
rect 49 744 51 764
rect 55 744 57 764
rect 69 744 71 764
rect 75 744 77 784
rect 151 744 153 784
rect 157 744 163 784
rect 167 744 169 784
rect 209 744 211 784
rect 215 764 228 784
rect 391 764 401 784
rect 215 744 219 764
rect 231 744 233 764
rect 237 744 243 764
rect 247 744 249 764
rect 261 744 263 764
rect 267 744 271 764
rect 275 744 277 764
rect 315 744 317 764
rect 321 744 325 764
rect 337 744 339 764
rect 343 744 349 764
rect 353 744 355 764
rect 367 744 371 764
rect 375 744 381 764
rect 385 744 387 764
rect 399 744 401 764
rect 405 744 407 784
rect 463 744 465 764
rect 469 744 471 764
rect 523 744 525 764
rect 529 744 531 764
rect 543 744 545 764
rect 549 744 551 764
rect 589 744 591 764
rect 595 744 597 764
rect 609 744 611 764
rect 615 744 617 764
rect 671 744 673 784
rect 677 744 683 784
rect 687 744 689 784
rect 750 744 752 804
rect 756 744 760 804
rect 764 744 768 804
rect 772 802 786 804
rect 772 744 774 802
rect 849 744 851 784
rect 855 774 871 784
rect 855 744 857 774
rect 869 744 871 774
rect 875 744 877 784
rect 889 744 891 784
rect 895 756 897 784
rect 909 756 911 784
rect 895 744 911 756
rect 915 744 917 784
rect 969 744 971 784
rect 975 772 991 784
rect 975 744 977 772
rect 989 744 991 772
rect 995 744 997 784
rect 1009 744 1011 784
rect 1015 744 1017 784
rect 1069 744 1071 784
rect 1075 772 1091 784
rect 1075 744 1077 772
rect 1089 744 1091 772
rect 1095 744 1097 784
rect 1109 744 1111 784
rect 1115 744 1117 784
rect 1243 744 1245 764
rect 1249 744 1251 764
rect 1263 744 1265 764
rect 1269 744 1271 764
rect 1283 744 1285 764
rect 1289 744 1291 764
rect 1349 744 1351 784
rect 1355 772 1371 784
rect 1355 744 1357 772
rect 1369 744 1371 772
rect 1375 744 1377 784
rect 1389 744 1391 784
rect 1395 744 1397 784
rect 1463 744 1465 764
rect 1469 744 1471 764
rect 1513 744 1515 784
rect 1519 764 1529 784
rect 1692 764 1705 784
rect 1519 744 1521 764
rect 1533 744 1535 764
rect 1539 744 1545 764
rect 1549 744 1553 764
rect 1565 744 1567 764
rect 1571 744 1577 764
rect 1581 744 1583 764
rect 1595 744 1599 764
rect 1603 744 1605 764
rect 1643 744 1645 764
rect 1649 744 1653 764
rect 1657 744 1659 764
rect 1671 744 1673 764
rect 1677 744 1683 764
rect 1687 744 1689 764
rect 1701 744 1705 764
rect 1709 744 1711 784
rect 1819 772 1831 792
rect 1749 744 1751 764
rect 1755 744 1757 764
rect 1809 752 1811 772
rect 1815 752 1817 772
rect 1829 752 1831 772
rect 1835 752 1841 792
rect 1845 784 1861 792
rect 1845 752 1847 784
rect 1859 752 1861 784
rect 1865 752 1871 792
rect 1875 752 1877 792
rect 1929 744 1931 784
rect 1935 772 1951 784
rect 1935 744 1937 772
rect 1949 744 1951 772
rect 1955 744 1957 784
rect 1969 744 1971 784
rect 1975 744 1977 784
rect 2031 744 2033 784
rect 2037 744 2043 784
rect 2047 744 2049 784
rect 2109 744 2111 784
rect 2115 764 2128 784
rect 2291 764 2301 784
rect 2115 744 2119 764
rect 2131 744 2133 764
rect 2137 744 2143 764
rect 2147 744 2149 764
rect 2161 744 2163 764
rect 2167 744 2171 764
rect 2175 744 2177 764
rect 2215 744 2217 764
rect 2221 744 2225 764
rect 2237 744 2239 764
rect 2243 744 2249 764
rect 2253 744 2255 764
rect 2267 744 2271 764
rect 2275 744 2281 764
rect 2285 744 2287 764
rect 2299 744 2301 764
rect 2305 744 2307 784
rect 2349 744 2351 764
rect 2355 744 2357 764
rect 2409 744 2411 784
rect 2415 774 2431 784
rect 2415 744 2417 774
rect 2429 744 2431 774
rect 2435 744 2437 784
rect 2449 744 2451 784
rect 2455 756 2457 784
rect 2469 756 2471 784
rect 2455 744 2471 756
rect 2475 744 2477 784
rect 2529 744 2531 764
rect 2535 744 2537 764
rect 2549 744 2551 764
rect 2555 744 2557 764
rect 2623 744 2625 784
rect 2629 744 2631 784
rect 2643 744 2645 784
rect 2649 772 2665 784
rect 2649 744 2651 772
rect 2663 744 2665 772
rect 2669 744 2671 784
rect 2723 744 2725 784
rect 2729 744 2731 784
rect 2743 744 2745 784
rect 2749 744 2751 784
rect 2763 744 2765 784
rect 2769 744 2771 784
rect 2783 744 2785 784
rect 2789 744 2791 784
rect 2803 744 2805 784
rect 2809 744 2811 784
rect 2823 744 2825 784
rect 2829 744 2831 784
rect 2843 744 2845 784
rect 2849 744 2851 784
rect 2863 744 2865 784
rect 2869 744 2871 784
rect 2912 744 2914 784
rect 2918 744 2922 784
rect 2926 744 2928 784
rect 2940 744 2944 764
rect 2948 744 2950 764
rect 3030 744 3032 764
rect 3036 744 3040 764
rect 3052 744 3054 784
rect 3058 744 3062 784
rect 3066 744 3068 784
rect 3123 752 3125 792
rect 3129 752 3135 792
rect 3139 784 3155 792
rect 3139 752 3141 784
rect 3153 752 3155 784
rect 3159 752 3165 792
rect 3169 772 3181 792
rect 3169 752 3171 772
rect 3183 752 3185 772
rect 3189 752 3191 772
rect 3243 752 3245 792
rect 3249 752 3255 792
rect 3259 784 3275 792
rect 3259 752 3261 784
rect 3273 752 3275 784
rect 3279 752 3285 792
rect 3289 772 3301 792
rect 3289 752 3291 772
rect 3303 752 3305 772
rect 3309 752 3311 772
rect 3363 744 3365 784
rect 3369 744 3371 784
rect 3383 744 3385 784
rect 3389 772 3405 784
rect 3389 744 3391 772
rect 3403 744 3405 772
rect 3409 744 3411 784
rect 3451 744 3453 784
rect 3457 744 3463 784
rect 3467 744 3469 784
rect 3539 772 3551 792
rect 3529 752 3531 772
rect 3535 752 3537 772
rect 3549 752 3551 772
rect 3555 752 3561 792
rect 3565 784 3581 792
rect 3565 752 3567 784
rect 3579 752 3581 784
rect 3585 752 3591 792
rect 3595 752 3597 792
rect 3663 744 3665 764
rect 3669 744 3671 764
rect 3723 752 3725 792
rect 3729 752 3735 792
rect 3739 784 3755 792
rect 3739 752 3741 784
rect 3753 752 3755 784
rect 3759 752 3765 792
rect 3769 772 3781 792
rect 3769 752 3771 772
rect 3783 752 3785 772
rect 3789 752 3791 772
rect 3833 744 3835 784
rect 3839 764 3849 784
rect 4012 764 4025 784
rect 3839 744 3841 764
rect 3853 744 3855 764
rect 3859 744 3865 764
rect 3869 744 3873 764
rect 3885 744 3887 764
rect 3891 744 3897 764
rect 3901 744 3903 764
rect 3915 744 3919 764
rect 3923 744 3925 764
rect 3963 744 3965 764
rect 3969 744 3973 764
rect 3977 744 3979 764
rect 3991 744 3993 764
rect 3997 744 4003 764
rect 4007 744 4009 764
rect 4021 744 4025 764
rect 4029 744 4031 784
rect 4079 772 4091 792
rect 4069 752 4071 772
rect 4075 752 4077 772
rect 4089 752 4091 772
rect 4095 752 4101 792
rect 4105 784 4121 792
rect 4105 752 4107 784
rect 4119 752 4121 784
rect 4125 752 4131 792
rect 4135 752 4137 792
rect 4192 744 4194 784
rect 4198 744 4202 784
rect 4206 744 4208 784
rect 4414 802 4428 804
rect 4220 744 4224 764
rect 4228 744 4230 764
rect 4289 744 4291 784
rect 4295 772 4311 784
rect 4295 744 4297 772
rect 4309 744 4311 772
rect 4315 744 4317 784
rect 4329 744 4331 784
rect 4335 744 4337 784
rect 4426 744 4428 802
rect 4432 744 4436 804
rect 4440 744 4444 804
rect 4448 744 4450 804
rect 4489 744 4491 764
rect 4495 744 4497 764
rect 4549 744 4551 784
rect 4555 772 4571 784
rect 4555 744 4557 772
rect 4569 744 4571 772
rect 4575 744 4577 784
rect 4589 744 4591 784
rect 4595 744 4597 784
rect 4651 744 4653 784
rect 4657 744 4663 784
rect 4667 744 4669 784
rect 4743 744 4745 764
rect 4749 744 4751 764
rect 4789 744 4791 784
rect 4795 772 4811 784
rect 4795 744 4797 772
rect 4809 744 4811 772
rect 4815 744 4817 784
rect 4829 744 4831 784
rect 4835 744 4837 784
rect 4891 744 4893 784
rect 4897 744 4903 784
rect 4907 744 4909 784
rect 4979 772 4991 792
rect 4969 752 4971 772
rect 4975 752 4977 772
rect 4989 752 4991 772
rect 4995 752 5001 792
rect 5005 784 5021 792
rect 5005 752 5007 784
rect 5019 752 5021 784
rect 5025 752 5031 792
rect 5035 752 5037 792
rect 5103 752 5105 792
rect 5109 752 5115 792
rect 5119 784 5135 792
rect 5119 752 5121 784
rect 5133 752 5135 784
rect 5139 752 5145 792
rect 5149 772 5161 792
rect 5149 752 5151 772
rect 5163 752 5165 772
rect 5169 752 5171 772
rect 5209 744 5211 784
rect 5215 744 5217 784
rect 5229 744 5231 784
rect 5235 744 5237 784
rect 5249 744 5251 784
rect 5255 744 5257 784
rect 5269 744 5271 784
rect 5275 744 5277 784
rect 5289 744 5291 784
rect 5295 744 5297 784
rect 5309 744 5311 784
rect 5315 744 5317 784
rect 5329 744 5331 784
rect 5335 744 5337 784
rect 5349 744 5351 784
rect 5355 744 5357 784
rect 5412 744 5414 784
rect 5418 744 5422 784
rect 5426 744 5428 784
rect 5874 802 5888 804
rect 5440 744 5444 764
rect 5448 744 5450 764
rect 5523 744 5525 764
rect 5529 744 5531 764
rect 5569 744 5571 784
rect 5575 772 5591 784
rect 5575 744 5577 772
rect 5589 744 5591 772
rect 5595 744 5597 784
rect 5609 744 5611 784
rect 5615 744 5617 784
rect 5671 744 5673 784
rect 5677 744 5683 784
rect 5687 744 5689 784
rect 5749 744 5751 784
rect 5755 772 5771 784
rect 5755 744 5757 772
rect 5769 744 5771 772
rect 5775 744 5777 784
rect 5789 744 5791 784
rect 5795 744 5797 784
rect 5886 744 5888 802
rect 5892 744 5896 804
rect 5900 744 5904 804
rect 5908 744 5910 804
rect 5953 744 5955 784
rect 5959 764 5969 784
rect 6132 764 6145 784
rect 5959 744 5961 764
rect 5973 744 5975 764
rect 5979 744 5985 764
rect 5989 744 5993 764
rect 6005 744 6007 764
rect 6011 744 6017 764
rect 6021 744 6023 764
rect 6035 744 6039 764
rect 6043 744 6045 764
rect 6083 744 6085 764
rect 6089 744 6093 764
rect 6097 744 6099 764
rect 6111 744 6113 764
rect 6117 744 6123 764
rect 6127 744 6129 764
rect 6141 744 6145 764
rect 6149 744 6151 784
rect 6189 744 6191 784
rect 6195 772 6211 784
rect 6195 744 6197 772
rect 6209 744 6211 772
rect 6215 744 6217 784
rect 6229 744 6231 784
rect 6235 744 6237 784
rect 6289 744 6291 784
rect 6295 772 6311 784
rect 6295 744 6297 772
rect 6309 744 6311 772
rect 6315 744 6317 784
rect 6329 744 6331 784
rect 6335 744 6337 784
rect 6411 744 6413 784
rect 6417 744 6423 784
rect 6427 744 6429 784
rect 6473 744 6475 784
rect 6479 764 6489 784
rect 6652 764 6665 784
rect 6479 744 6481 764
rect 6493 744 6495 764
rect 6499 744 6505 764
rect 6509 744 6513 764
rect 6525 744 6527 764
rect 6531 744 6537 764
rect 6541 744 6543 764
rect 6555 744 6559 764
rect 6563 744 6565 764
rect 6603 744 6605 764
rect 6609 744 6613 764
rect 6617 744 6619 764
rect 6631 744 6633 764
rect 6637 744 6643 764
rect 6647 744 6649 764
rect 6661 744 6665 764
rect 6669 744 6671 784
rect 29 696 31 716
rect 35 696 37 716
rect 91 676 93 716
rect 97 676 103 716
rect 107 676 109 716
rect 172 676 174 716
rect 178 676 182 716
rect 186 676 188 716
rect 200 696 204 716
rect 208 696 210 716
rect 269 696 271 716
rect 275 696 277 716
rect 350 696 352 716
rect 356 696 360 716
rect 372 676 374 716
rect 378 676 382 716
rect 386 676 388 716
rect 430 656 432 716
rect 436 656 440 716
rect 444 656 448 716
rect 452 658 454 716
rect 551 676 553 716
rect 557 676 563 716
rect 567 676 569 716
rect 452 656 466 658
rect 646 658 648 716
rect 634 656 648 658
rect 652 656 656 716
rect 660 656 664 716
rect 668 656 670 716
rect 709 696 711 716
rect 715 696 717 716
rect 769 696 771 716
rect 775 696 777 716
rect 843 696 845 716
rect 849 696 851 716
rect 863 696 865 716
rect 869 696 871 716
rect 983 696 985 716
rect 989 696 991 716
rect 1003 696 1005 716
rect 1009 696 1011 716
rect 1023 696 1025 716
rect 1029 696 1031 716
rect 1093 676 1095 716
rect 1099 696 1101 716
rect 1113 696 1115 716
rect 1119 696 1125 716
rect 1129 696 1133 716
rect 1145 696 1147 716
rect 1151 696 1157 716
rect 1161 696 1163 716
rect 1175 696 1179 716
rect 1183 696 1185 716
rect 1223 696 1225 716
rect 1229 696 1233 716
rect 1237 696 1239 716
rect 1251 696 1253 716
rect 1257 696 1263 716
rect 1267 696 1269 716
rect 1281 696 1285 716
rect 1099 676 1109 696
rect 1272 676 1285 696
rect 1289 676 1291 716
rect 1329 696 1331 716
rect 1335 696 1339 716
rect 1351 676 1353 716
rect 1357 676 1359 716
rect 1411 676 1413 716
rect 1417 676 1423 716
rect 1427 676 1429 716
rect 1493 676 1495 716
rect 1499 696 1501 716
rect 1513 696 1515 716
rect 1519 696 1525 716
rect 1529 696 1533 716
rect 1545 696 1547 716
rect 1551 696 1557 716
rect 1561 696 1563 716
rect 1575 696 1579 716
rect 1583 696 1585 716
rect 1623 696 1625 716
rect 1629 696 1633 716
rect 1637 696 1639 716
rect 1651 696 1653 716
rect 1657 696 1663 716
rect 1667 696 1669 716
rect 1681 696 1685 716
rect 1499 676 1509 696
rect 1672 676 1685 696
rect 1689 676 1691 716
rect 1733 676 1735 716
rect 1739 696 1741 716
rect 1753 696 1755 716
rect 1759 696 1765 716
rect 1769 696 1773 716
rect 1785 696 1787 716
rect 1791 696 1797 716
rect 1801 696 1803 716
rect 1815 696 1819 716
rect 1823 696 1825 716
rect 1863 696 1865 716
rect 1869 696 1873 716
rect 1877 696 1879 716
rect 1891 696 1893 716
rect 1897 696 1903 716
rect 1907 696 1909 716
rect 1921 696 1925 716
rect 1739 676 1749 696
rect 1912 676 1925 696
rect 1929 676 1931 716
rect 1973 676 1975 716
rect 1979 696 1981 716
rect 1993 696 1995 716
rect 1999 696 2005 716
rect 2009 696 2013 716
rect 2025 696 2027 716
rect 2031 696 2037 716
rect 2041 696 2043 716
rect 2055 696 2059 716
rect 2063 696 2065 716
rect 2103 696 2105 716
rect 2109 696 2113 716
rect 2117 696 2119 716
rect 2131 696 2133 716
rect 2137 696 2143 716
rect 2147 696 2149 716
rect 2161 696 2165 716
rect 1979 676 1989 696
rect 2152 676 2165 696
rect 2169 676 2171 716
rect 2213 676 2215 716
rect 2219 696 2221 716
rect 2233 696 2235 716
rect 2239 696 2245 716
rect 2249 696 2253 716
rect 2265 696 2267 716
rect 2271 696 2277 716
rect 2281 696 2283 716
rect 2295 696 2299 716
rect 2303 696 2305 716
rect 2343 696 2345 716
rect 2349 696 2353 716
rect 2357 696 2359 716
rect 2371 696 2373 716
rect 2377 696 2383 716
rect 2387 696 2389 716
rect 2401 696 2405 716
rect 2219 676 2229 696
rect 2392 676 2405 696
rect 2409 676 2411 716
rect 2449 676 2451 716
rect 2455 696 2459 716
rect 2471 696 2473 716
rect 2477 696 2483 716
rect 2487 696 2489 716
rect 2501 696 2503 716
rect 2507 696 2511 716
rect 2515 696 2517 716
rect 2555 696 2557 716
rect 2561 696 2565 716
rect 2577 696 2579 716
rect 2583 696 2589 716
rect 2593 696 2595 716
rect 2607 696 2611 716
rect 2615 696 2621 716
rect 2625 696 2627 716
rect 2639 696 2641 716
rect 2455 676 2468 696
rect 2631 676 2641 696
rect 2645 676 2647 716
rect 2724 676 2726 716
rect 2730 676 2734 716
rect 2738 676 2740 716
rect 2752 676 2754 716
rect 2758 676 2762 716
rect 2766 676 2768 716
rect 2823 696 2825 716
rect 2829 696 2831 716
rect 2890 696 2892 716
rect 2896 696 2900 716
rect 2912 676 2914 716
rect 2918 676 2922 716
rect 2926 676 2928 716
rect 2969 696 2971 716
rect 2975 696 2977 716
rect 3029 676 3031 716
rect 3035 688 3037 716
rect 3049 688 3051 716
rect 3035 676 3051 688
rect 3055 676 3057 716
rect 3069 676 3071 716
rect 3075 676 3077 716
rect 3131 676 3133 716
rect 3137 676 3143 716
rect 3147 676 3149 716
rect 3210 656 3212 716
rect 3216 656 3220 716
rect 3224 656 3228 716
rect 3232 658 3234 716
rect 3309 696 3311 716
rect 3315 696 3317 716
rect 3232 656 3246 658
rect 3369 676 3371 716
rect 3375 688 3377 716
rect 3389 688 3391 716
rect 3375 676 3391 688
rect 3395 676 3397 716
rect 3409 676 3411 716
rect 3415 676 3417 716
rect 3471 676 3473 716
rect 3477 676 3483 716
rect 3487 676 3489 716
rect 3552 676 3554 716
rect 3558 676 3562 716
rect 3566 676 3568 716
rect 3580 696 3584 716
rect 3588 696 3590 716
rect 3649 696 3651 716
rect 3655 696 3657 716
rect 3669 696 3671 716
rect 3675 696 3677 716
rect 3729 676 3731 716
rect 3735 688 3737 716
rect 3749 688 3751 716
rect 3735 676 3751 688
rect 3755 676 3757 716
rect 3769 676 3771 716
rect 3775 676 3777 716
rect 3866 658 3868 716
rect 3854 656 3868 658
rect 3872 656 3876 716
rect 3880 656 3884 716
rect 3888 656 3890 716
rect 3929 676 3931 716
rect 3935 696 3939 716
rect 3951 696 3953 716
rect 3957 696 3963 716
rect 3967 696 3969 716
rect 3981 696 3983 716
rect 3987 696 3991 716
rect 3995 696 3997 716
rect 4035 696 4037 716
rect 4041 696 4045 716
rect 4057 696 4059 716
rect 4063 696 4069 716
rect 4073 696 4075 716
rect 4087 696 4091 716
rect 4095 696 4101 716
rect 4105 696 4107 716
rect 4119 696 4121 716
rect 3935 676 3948 696
rect 4111 676 4121 696
rect 4125 676 4127 716
rect 4183 696 4185 716
rect 4189 696 4191 716
rect 4203 696 4205 716
rect 4209 696 4211 716
rect 4249 676 4251 716
rect 4255 696 4259 716
rect 4271 696 4273 716
rect 4277 696 4283 716
rect 4287 696 4289 716
rect 4301 696 4303 716
rect 4307 696 4311 716
rect 4315 696 4317 716
rect 4355 696 4357 716
rect 4361 696 4365 716
rect 4377 696 4379 716
rect 4383 696 4389 716
rect 4393 696 4395 716
rect 4407 696 4411 716
rect 4415 696 4421 716
rect 4425 696 4427 716
rect 4439 696 4441 716
rect 4255 676 4268 696
rect 4431 676 4441 696
rect 4445 676 4447 716
rect 4489 696 4491 716
rect 4495 696 4497 716
rect 4552 676 4554 716
rect 4558 676 4562 716
rect 4566 676 4568 716
rect 4580 676 4582 716
rect 4586 676 4590 716
rect 4594 676 4596 716
rect 4690 696 4692 716
rect 4696 696 4700 716
rect 4712 676 4714 716
rect 4718 676 4722 716
rect 4726 676 4728 716
rect 4783 676 4785 716
rect 4789 676 4791 716
rect 4803 676 4805 716
rect 4809 688 4811 716
rect 4823 688 4825 716
rect 4809 676 4825 688
rect 4829 676 4831 716
rect 4871 676 4873 716
rect 4877 676 4883 716
rect 4887 676 4889 716
rect 4963 696 4965 716
rect 4969 696 4971 716
rect 5023 668 5025 708
rect 5029 668 5035 708
rect 5039 676 5041 708
rect 5053 676 5055 708
rect 5039 668 5055 676
rect 5059 668 5065 708
rect 5069 688 5071 708
rect 5083 688 5085 708
rect 5089 688 5091 708
rect 5069 668 5081 688
rect 5130 656 5132 716
rect 5136 656 5140 716
rect 5144 656 5148 716
rect 5152 658 5154 716
rect 5229 676 5231 716
rect 5235 696 5239 716
rect 5251 696 5253 716
rect 5257 696 5263 716
rect 5267 696 5269 716
rect 5281 696 5283 716
rect 5287 696 5291 716
rect 5295 696 5297 716
rect 5335 696 5337 716
rect 5341 696 5345 716
rect 5357 696 5359 716
rect 5363 696 5369 716
rect 5373 696 5375 716
rect 5387 696 5391 716
rect 5395 696 5401 716
rect 5405 696 5407 716
rect 5419 696 5421 716
rect 5235 676 5248 696
rect 5152 656 5166 658
rect 5411 676 5421 696
rect 5425 676 5427 716
rect 5469 676 5471 716
rect 5475 676 5477 716
rect 5529 688 5531 708
rect 5535 688 5537 708
rect 5549 688 5551 708
rect 5539 668 5551 688
rect 5555 668 5561 708
rect 5565 676 5567 708
rect 5579 676 5581 708
rect 5565 668 5581 676
rect 5585 668 5591 708
rect 5595 668 5597 708
rect 5663 696 5665 716
rect 5669 696 5671 716
rect 5683 696 5685 716
rect 5689 696 5691 716
rect 5743 696 5745 716
rect 5749 696 5751 716
rect 5763 696 5765 716
rect 5769 696 5771 716
rect 5823 696 5825 716
rect 5829 696 5831 716
rect 5843 696 5845 716
rect 5849 696 5851 716
rect 5889 696 5891 716
rect 5895 696 5897 716
rect 5909 696 5911 716
rect 5915 696 5917 716
rect 5983 696 5985 716
rect 5989 696 5991 716
rect 6003 696 6005 716
rect 6009 696 6011 716
rect 6049 676 6051 716
rect 6055 688 6057 716
rect 6069 688 6071 716
rect 6055 676 6071 688
rect 6075 676 6077 716
rect 6089 676 6091 716
rect 6095 676 6097 716
rect 6149 676 6151 716
rect 6155 688 6157 716
rect 6169 688 6171 716
rect 6155 676 6171 688
rect 6175 676 6177 716
rect 6189 676 6191 716
rect 6195 676 6197 716
rect 6271 676 6273 716
rect 6277 676 6283 716
rect 6287 676 6289 716
rect 6333 676 6335 716
rect 6339 696 6341 716
rect 6353 696 6355 716
rect 6359 696 6365 716
rect 6369 696 6373 716
rect 6385 696 6387 716
rect 6391 696 6397 716
rect 6401 696 6403 716
rect 6415 696 6419 716
rect 6423 696 6425 716
rect 6463 696 6465 716
rect 6469 696 6473 716
rect 6477 696 6479 716
rect 6491 696 6493 716
rect 6497 696 6503 716
rect 6507 696 6509 716
rect 6521 696 6525 716
rect 6339 676 6349 696
rect 6512 676 6525 696
rect 6529 676 6531 716
rect 6569 696 6571 716
rect 6575 696 6577 716
rect 6629 696 6631 716
rect 6635 696 6637 716
rect 29 264 31 304
rect 35 284 48 304
rect 211 284 221 304
rect 35 264 39 284
rect 51 264 53 284
rect 57 264 63 284
rect 67 264 69 284
rect 81 264 83 284
rect 87 264 91 284
rect 95 264 97 284
rect 135 264 137 284
rect 141 264 145 284
rect 157 264 159 284
rect 163 264 169 284
rect 173 264 175 284
rect 187 264 191 284
rect 195 264 201 284
rect 205 264 207 284
rect 219 264 221 284
rect 225 264 227 304
rect 273 264 275 304
rect 279 284 289 304
rect 452 284 465 304
rect 279 264 281 284
rect 293 264 295 284
rect 299 264 305 284
rect 309 264 313 284
rect 325 264 327 284
rect 331 264 337 284
rect 341 264 343 284
rect 355 264 359 284
rect 363 264 365 284
rect 403 264 405 284
rect 409 264 413 284
rect 417 264 419 284
rect 431 264 433 284
rect 437 264 443 284
rect 447 264 449 284
rect 461 264 465 284
rect 469 264 471 304
rect 510 264 512 324
rect 516 264 520 324
rect 524 264 528 324
rect 532 322 546 324
rect 532 264 534 322
rect 609 264 611 284
rect 615 264 617 284
rect 629 264 631 284
rect 635 264 637 284
rect 703 264 705 284
rect 709 264 711 284
rect 723 264 725 284
rect 729 264 731 284
rect 771 264 773 304
rect 777 264 783 304
rect 787 264 789 304
rect 863 264 865 284
rect 869 264 871 284
rect 913 264 915 304
rect 919 284 929 304
rect 1092 284 1105 304
rect 919 264 921 284
rect 933 264 935 284
rect 939 264 945 284
rect 949 264 953 284
rect 965 264 967 284
rect 971 264 977 284
rect 981 264 983 284
rect 995 264 999 284
rect 1003 264 1005 284
rect 1043 264 1045 284
rect 1049 264 1053 284
rect 1057 264 1059 284
rect 1071 264 1073 284
rect 1077 264 1083 284
rect 1087 264 1089 284
rect 1101 264 1105 284
rect 1109 264 1111 304
rect 1161 264 1163 304
rect 1167 264 1169 304
rect 1181 264 1185 284
rect 1189 264 1191 284
rect 1229 264 1231 284
rect 1235 264 1239 284
rect 1251 264 1253 304
rect 1257 264 1259 304
rect 1309 264 1311 284
rect 1315 264 1319 284
rect 1331 264 1333 304
rect 1337 264 1339 304
rect 1403 264 1405 284
rect 1409 264 1411 284
rect 1449 264 1451 304
rect 1455 292 1471 304
rect 1455 264 1457 292
rect 1469 264 1471 292
rect 1475 264 1477 304
rect 1489 264 1491 304
rect 1495 264 1497 304
rect 1563 264 1565 284
rect 1569 264 1571 284
rect 1609 264 1611 304
rect 1615 292 1631 304
rect 1615 264 1617 292
rect 1629 264 1631 292
rect 1635 264 1637 304
rect 1649 264 1651 304
rect 1655 264 1657 304
rect 1713 264 1715 304
rect 1719 284 1729 304
rect 1892 284 1905 304
rect 1719 264 1721 284
rect 1733 264 1735 284
rect 1739 264 1745 284
rect 1749 264 1753 284
rect 1765 264 1767 284
rect 1771 264 1777 284
rect 1781 264 1783 284
rect 1795 264 1799 284
rect 1803 264 1805 284
rect 1843 264 1845 284
rect 1849 264 1853 284
rect 1857 264 1859 284
rect 1871 264 1873 284
rect 1877 264 1883 284
rect 1887 264 1889 284
rect 1901 264 1905 284
rect 1909 264 1911 304
rect 1963 264 1965 284
rect 1969 264 1971 284
rect 2023 264 2025 284
rect 2029 264 2031 284
rect 2069 264 2071 304
rect 2075 292 2091 304
rect 2075 264 2077 292
rect 2089 264 2091 292
rect 2095 264 2097 304
rect 2109 264 2111 304
rect 2115 264 2117 304
rect 2169 264 2171 284
rect 2175 264 2177 284
rect 2229 264 2231 304
rect 2235 294 2251 304
rect 2235 264 2237 294
rect 2249 264 2251 294
rect 2255 264 2257 304
rect 2269 264 2271 304
rect 2275 276 2277 304
rect 2289 276 2291 304
rect 2275 264 2291 276
rect 2295 264 2297 304
rect 2363 264 2365 304
rect 2369 264 2371 304
rect 2383 264 2385 304
rect 2389 292 2405 304
rect 2389 264 2391 292
rect 2403 264 2405 292
rect 2409 264 2411 304
rect 2449 264 2451 284
rect 2455 264 2457 284
rect 2469 264 2471 284
rect 2475 264 2477 284
rect 2533 264 2535 304
rect 2539 284 2549 304
rect 2712 284 2725 304
rect 2539 264 2541 284
rect 2553 264 2555 284
rect 2559 264 2565 284
rect 2569 264 2573 284
rect 2585 264 2587 284
rect 2591 264 2597 284
rect 2601 264 2603 284
rect 2615 264 2619 284
rect 2623 264 2625 284
rect 2663 264 2665 284
rect 2669 264 2673 284
rect 2677 264 2679 284
rect 2691 264 2693 284
rect 2697 264 2703 284
rect 2707 264 2709 284
rect 2721 264 2725 284
rect 2729 264 2731 304
rect 2783 264 2785 304
rect 2789 264 2791 304
rect 2803 264 2805 304
rect 2809 292 2825 304
rect 2809 264 2811 292
rect 2823 264 2825 292
rect 2829 264 2831 304
rect 2869 264 2871 284
rect 2875 264 2877 284
rect 2889 264 2891 284
rect 2895 264 2897 284
rect 2953 264 2955 304
rect 2959 284 2969 304
rect 3132 284 3145 304
rect 2959 264 2961 284
rect 2973 264 2975 284
rect 2979 264 2985 284
rect 2989 264 2993 284
rect 3005 264 3007 284
rect 3011 264 3017 284
rect 3021 264 3023 284
rect 3035 264 3039 284
rect 3043 264 3045 284
rect 3083 264 3085 284
rect 3089 264 3093 284
rect 3097 264 3099 284
rect 3111 264 3113 284
rect 3117 264 3123 284
rect 3127 264 3129 284
rect 3141 264 3145 284
rect 3149 264 3151 304
rect 3191 264 3193 304
rect 3197 264 3203 304
rect 3207 264 3209 304
rect 3283 264 3285 304
rect 3289 264 3291 304
rect 3303 264 3305 304
rect 3309 292 3325 304
rect 3309 264 3311 292
rect 3323 264 3325 292
rect 3329 264 3331 304
rect 3369 264 3371 284
rect 3375 264 3377 284
rect 3389 264 3391 284
rect 3395 264 3397 284
rect 3470 264 3472 284
rect 3476 264 3480 284
rect 3492 264 3494 304
rect 3498 264 3502 304
rect 3506 264 3508 304
rect 3549 264 3551 304
rect 3555 292 3571 304
rect 3555 264 3557 292
rect 3569 264 3571 292
rect 3575 264 3577 304
rect 3589 264 3591 304
rect 3595 264 3597 304
rect 3649 264 3651 284
rect 3655 264 3657 284
rect 3669 264 3671 284
rect 3675 264 3677 284
rect 3732 264 3734 304
rect 3738 264 3742 304
rect 3746 264 3748 304
rect 4034 322 4048 324
rect 3760 264 3764 284
rect 3768 264 3770 284
rect 3843 264 3845 284
rect 3849 264 3851 284
rect 3863 264 3865 284
rect 3869 264 3871 284
rect 3909 264 3911 304
rect 3915 292 3931 304
rect 3915 264 3917 292
rect 3929 264 3931 292
rect 3935 264 3937 304
rect 3949 264 3951 304
rect 3955 264 3957 304
rect 4046 264 4048 322
rect 4052 264 4056 324
rect 4060 264 4064 324
rect 4068 264 4070 324
rect 4109 264 4111 284
rect 4115 264 4117 284
rect 4129 264 4131 284
rect 4135 264 4137 284
rect 4189 264 4191 304
rect 4195 284 4208 304
rect 4371 284 4381 304
rect 4195 264 4199 284
rect 4211 264 4213 284
rect 4217 264 4223 284
rect 4227 264 4229 284
rect 4241 264 4243 284
rect 4247 264 4251 284
rect 4255 264 4257 284
rect 4295 264 4297 284
rect 4301 264 4305 284
rect 4317 264 4319 284
rect 4323 264 4329 284
rect 4333 264 4335 284
rect 4347 264 4351 284
rect 4355 264 4361 284
rect 4365 264 4367 284
rect 4379 264 4381 284
rect 4385 264 4387 304
rect 4429 264 4431 284
rect 4435 264 4437 284
rect 4449 264 4451 284
rect 4455 264 4457 284
rect 4523 264 4525 304
rect 4529 264 4531 304
rect 4543 264 4545 304
rect 4549 292 4565 304
rect 4549 264 4551 292
rect 4563 264 4565 292
rect 4569 264 4571 304
rect 4609 264 4611 284
rect 4615 264 4617 284
rect 4629 264 4631 284
rect 4635 264 4637 284
rect 4703 264 4705 304
rect 4709 276 4711 304
rect 4723 276 4725 304
rect 4709 264 4725 276
rect 4729 264 4731 304
rect 4743 264 4745 304
rect 4749 294 4765 304
rect 4749 264 4751 294
rect 4763 264 4765 294
rect 4769 264 4771 304
rect 4823 264 4825 284
rect 4829 264 4831 284
rect 4873 264 4875 304
rect 4879 284 4889 304
rect 5052 284 5065 304
rect 4879 264 4881 284
rect 4893 264 4895 284
rect 4899 264 4905 284
rect 4909 264 4913 284
rect 4925 264 4927 284
rect 4931 264 4937 284
rect 4941 264 4943 284
rect 4955 264 4959 284
rect 4963 264 4965 284
rect 5003 264 5005 284
rect 5009 264 5013 284
rect 5017 264 5019 284
rect 5031 264 5033 284
rect 5037 264 5043 284
rect 5047 264 5049 284
rect 5061 264 5065 284
rect 5069 264 5071 304
rect 5130 264 5132 284
rect 5136 264 5140 284
rect 5152 264 5154 304
rect 5158 264 5162 304
rect 5166 264 5168 304
rect 5209 264 5211 284
rect 5215 264 5217 284
rect 5229 264 5231 284
rect 5235 264 5237 284
rect 5303 264 5305 304
rect 5309 264 5311 304
rect 5323 264 5325 304
rect 5329 292 5345 304
rect 5329 264 5331 292
rect 5343 264 5345 292
rect 5349 264 5351 304
rect 5389 264 5391 284
rect 5395 264 5397 284
rect 5409 264 5411 284
rect 5415 264 5417 284
rect 5472 264 5474 304
rect 5478 264 5482 304
rect 5486 264 5488 304
rect 5500 264 5504 284
rect 5508 264 5510 284
rect 5570 264 5572 324
rect 5576 264 5580 324
rect 5584 264 5588 324
rect 5592 322 5606 324
rect 5592 264 5594 322
rect 5669 264 5671 304
rect 5675 292 5691 304
rect 5675 264 5677 292
rect 5689 264 5691 292
rect 5695 264 5697 304
rect 5709 264 5711 304
rect 5715 264 5717 304
rect 5791 264 5793 304
rect 5797 264 5803 304
rect 5807 264 5809 304
rect 5863 264 5865 304
rect 5869 264 5871 304
rect 5883 264 5885 304
rect 5889 292 5905 304
rect 5889 264 5891 292
rect 5903 264 5905 292
rect 5909 264 5911 304
rect 5949 264 5951 304
rect 5955 292 5971 304
rect 5955 264 5957 292
rect 5969 264 5971 292
rect 5975 264 5977 304
rect 5989 264 5991 304
rect 5995 264 5997 304
rect 6049 264 6051 304
rect 6055 292 6071 304
rect 6055 264 6057 292
rect 6069 264 6071 292
rect 6075 264 6077 304
rect 6089 264 6091 304
rect 6095 264 6097 304
rect 6163 264 6165 284
rect 6169 264 6171 284
rect 6183 264 6185 284
rect 6189 264 6191 284
rect 6243 264 6245 284
rect 6249 264 6251 284
rect 6263 264 6265 284
rect 6269 264 6271 284
rect 6323 264 6325 304
rect 6329 276 6331 304
rect 6343 276 6345 304
rect 6329 264 6345 276
rect 6349 264 6351 304
rect 6363 264 6365 304
rect 6369 294 6385 304
rect 6369 264 6371 294
rect 6383 264 6385 294
rect 6389 264 6391 304
rect 6433 264 6435 304
rect 6439 284 6449 304
rect 6612 284 6625 304
rect 6439 264 6441 284
rect 6453 264 6455 284
rect 6459 264 6465 284
rect 6469 264 6473 284
rect 6485 264 6487 284
rect 6491 264 6497 284
rect 6501 264 6503 284
rect 6515 264 6519 284
rect 6523 264 6525 284
rect 6563 264 6565 284
rect 6569 264 6573 284
rect 6577 264 6579 284
rect 6591 264 6593 284
rect 6597 264 6603 284
rect 6607 264 6609 284
rect 6621 264 6625 284
rect 6629 264 6631 304
rect 29 196 31 236
rect 35 216 39 236
rect 51 216 53 236
rect 57 216 63 236
rect 67 216 69 236
rect 81 216 83 236
rect 87 216 91 236
rect 95 216 97 236
rect 135 216 137 236
rect 141 216 145 236
rect 157 216 159 236
rect 163 216 169 236
rect 173 216 175 236
rect 187 216 191 236
rect 195 216 201 236
rect 205 216 207 236
rect 219 216 221 236
rect 35 196 48 216
rect 211 196 221 216
rect 225 196 227 236
rect 269 196 271 236
rect 275 216 279 236
rect 291 216 293 236
rect 297 216 303 236
rect 307 216 309 236
rect 321 216 323 236
rect 327 216 331 236
rect 335 216 337 236
rect 375 216 377 236
rect 381 216 385 236
rect 397 216 399 236
rect 403 216 409 236
rect 413 216 415 236
rect 427 216 431 236
rect 435 216 441 236
rect 445 216 447 236
rect 459 216 461 236
rect 275 196 288 216
rect 451 196 461 216
rect 465 196 467 236
rect 521 196 523 236
rect 527 196 529 236
rect 541 216 545 236
rect 549 216 551 236
rect 589 216 591 236
rect 595 216 599 236
rect 611 196 613 236
rect 617 196 619 236
rect 681 196 683 236
rect 687 196 689 236
rect 701 216 705 236
rect 709 216 711 236
rect 749 196 751 236
rect 755 216 759 236
rect 771 216 773 236
rect 777 216 783 236
rect 787 216 789 236
rect 801 216 803 236
rect 807 216 811 236
rect 815 216 817 236
rect 855 216 857 236
rect 861 216 865 236
rect 877 216 879 236
rect 883 216 889 236
rect 893 216 895 236
rect 907 216 911 236
rect 915 216 921 236
rect 925 216 927 236
rect 939 216 941 236
rect 755 196 768 216
rect 931 196 941 216
rect 945 196 947 236
rect 989 216 991 236
rect 995 216 999 236
rect 1011 196 1013 236
rect 1017 196 1019 236
rect 1091 196 1093 236
rect 1097 196 1103 236
rect 1107 196 1109 236
rect 1163 196 1165 236
rect 1169 196 1171 236
rect 1183 196 1185 236
rect 1189 208 1191 236
rect 1203 208 1205 236
rect 1189 196 1205 208
rect 1209 196 1211 236
rect 1253 196 1255 236
rect 1259 216 1261 236
rect 1273 216 1275 236
rect 1279 216 1285 236
rect 1289 216 1293 236
rect 1305 216 1307 236
rect 1311 216 1317 236
rect 1321 216 1323 236
rect 1335 216 1339 236
rect 1343 216 1345 236
rect 1383 216 1385 236
rect 1389 216 1393 236
rect 1397 216 1399 236
rect 1411 216 1413 236
rect 1417 216 1423 236
rect 1427 216 1429 236
rect 1441 216 1445 236
rect 1259 196 1269 216
rect 1432 196 1445 216
rect 1449 196 1451 236
rect 1503 216 1505 236
rect 1509 216 1511 236
rect 1551 196 1553 236
rect 1557 196 1563 236
rect 1567 196 1569 236
rect 1643 196 1645 236
rect 1649 196 1651 236
rect 1663 196 1665 236
rect 1669 208 1671 236
rect 1683 208 1685 236
rect 1669 196 1685 208
rect 1689 196 1691 236
rect 1729 216 1731 236
rect 1735 216 1737 236
rect 1791 196 1793 236
rect 1797 196 1803 236
rect 1807 196 1809 236
rect 1871 196 1873 236
rect 1877 196 1883 236
rect 1887 196 1889 236
rect 1951 196 1953 236
rect 1957 196 1963 236
rect 1967 196 1969 236
rect 2043 196 2045 236
rect 2049 196 2051 236
rect 2063 196 2065 236
rect 2069 208 2071 236
rect 2083 208 2085 236
rect 2069 196 2085 208
rect 2089 196 2091 236
rect 2133 196 2135 236
rect 2139 216 2141 236
rect 2153 216 2155 236
rect 2159 216 2165 236
rect 2169 216 2173 236
rect 2185 216 2187 236
rect 2191 216 2197 236
rect 2201 216 2203 236
rect 2215 216 2219 236
rect 2223 216 2225 236
rect 2263 216 2265 236
rect 2269 216 2273 236
rect 2277 216 2279 236
rect 2291 216 2293 236
rect 2297 216 2303 236
rect 2307 216 2309 236
rect 2321 216 2325 236
rect 2139 196 2149 216
rect 2312 196 2325 216
rect 2329 196 2331 236
rect 2371 196 2373 236
rect 2377 196 2383 236
rect 2387 196 2389 236
rect 2471 196 2473 236
rect 2477 196 2483 236
rect 2487 196 2489 236
rect 2543 196 2545 236
rect 2549 196 2551 236
rect 2563 196 2565 236
rect 2569 208 2571 236
rect 2583 208 2585 236
rect 2569 196 2585 208
rect 2589 196 2591 236
rect 2643 216 2645 236
rect 2649 216 2651 236
rect 2693 196 2695 236
rect 2699 216 2701 236
rect 2713 216 2715 236
rect 2719 216 2725 236
rect 2729 216 2733 236
rect 2745 216 2747 236
rect 2751 216 2757 236
rect 2761 216 2763 236
rect 2775 216 2779 236
rect 2783 216 2785 236
rect 2823 216 2825 236
rect 2829 216 2833 236
rect 2837 216 2839 236
rect 2851 216 2853 236
rect 2857 216 2863 236
rect 2867 216 2869 236
rect 2881 216 2885 236
rect 2699 196 2709 216
rect 2872 196 2885 216
rect 2889 196 2891 236
rect 2943 196 2945 236
rect 2949 196 2951 236
rect 2963 196 2965 236
rect 2969 208 2971 236
rect 2983 208 2985 236
rect 2969 196 2985 208
rect 2989 196 2991 236
rect 3043 216 3045 236
rect 3049 216 3051 236
rect 3063 216 3065 236
rect 3069 216 3071 236
rect 3123 196 3125 236
rect 3129 224 3145 236
rect 3129 196 3131 224
rect 3143 196 3145 224
rect 3149 196 3151 236
rect 3163 196 3165 236
rect 3169 206 3171 236
rect 3183 206 3185 236
rect 3169 196 3185 206
rect 3189 196 3191 236
rect 3243 216 3245 236
rect 3249 216 3251 236
rect 3289 196 3291 236
rect 3295 216 3299 236
rect 3311 216 3313 236
rect 3317 216 3323 236
rect 3327 216 3329 236
rect 3341 216 3343 236
rect 3347 216 3351 236
rect 3355 216 3357 236
rect 3395 216 3397 236
rect 3401 216 3405 236
rect 3417 216 3419 236
rect 3423 216 3429 236
rect 3433 216 3435 236
rect 3447 216 3451 236
rect 3455 216 3461 236
rect 3465 216 3467 236
rect 3479 216 3481 236
rect 3295 196 3308 216
rect 3471 196 3481 216
rect 3485 196 3487 236
rect 3551 196 3553 236
rect 3557 196 3563 236
rect 3567 196 3569 236
rect 3623 196 3625 236
rect 3629 196 3631 236
rect 3643 196 3645 236
rect 3649 208 3651 236
rect 3663 208 3665 236
rect 3649 196 3665 208
rect 3669 196 3671 236
rect 3709 196 3711 236
rect 3715 208 3717 236
rect 3729 208 3731 236
rect 3715 196 3731 208
rect 3735 196 3737 236
rect 3749 196 3751 236
rect 3755 196 3757 236
rect 3809 196 3811 236
rect 3815 216 3819 236
rect 3831 216 3833 236
rect 3837 216 3843 236
rect 3847 216 3849 236
rect 3861 216 3863 236
rect 3867 216 3871 236
rect 3875 216 3877 236
rect 3915 216 3917 236
rect 3921 216 3925 236
rect 3937 216 3939 236
rect 3943 216 3949 236
rect 3953 216 3955 236
rect 3967 216 3971 236
rect 3975 216 3981 236
rect 3985 216 3987 236
rect 3999 216 4001 236
rect 3815 196 3828 216
rect 3991 196 4001 216
rect 4005 196 4007 236
rect 4049 196 4051 236
rect 4055 208 4057 236
rect 4069 208 4071 236
rect 4055 196 4071 208
rect 4075 196 4077 236
rect 4089 196 4091 236
rect 4095 196 4097 236
rect 4149 196 4151 236
rect 4155 208 4157 236
rect 4169 208 4171 236
rect 4155 196 4171 208
rect 4175 196 4177 236
rect 4189 196 4191 236
rect 4195 196 4197 236
rect 4251 196 4253 236
rect 4257 196 4263 236
rect 4267 196 4269 236
rect 4329 196 4331 236
rect 4335 216 4339 236
rect 4351 216 4353 236
rect 4357 216 4363 236
rect 4367 216 4369 236
rect 4381 216 4383 236
rect 4387 216 4391 236
rect 4395 216 4397 236
rect 4435 216 4437 236
rect 4441 216 4445 236
rect 4457 216 4459 236
rect 4463 216 4469 236
rect 4473 216 4475 236
rect 4487 216 4491 236
rect 4495 216 4501 236
rect 4505 216 4507 236
rect 4519 216 4521 236
rect 4335 196 4348 216
rect 4511 196 4521 216
rect 4525 196 4527 236
rect 4569 196 4571 236
rect 4575 208 4577 236
rect 4589 208 4591 236
rect 4575 196 4591 208
rect 4595 196 4597 236
rect 4609 196 4611 236
rect 4615 196 4617 236
rect 4669 196 4671 236
rect 4675 208 4677 236
rect 4689 208 4691 236
rect 4675 196 4691 208
rect 4695 196 4697 236
rect 4709 196 4711 236
rect 4715 196 4717 236
rect 4771 196 4773 236
rect 4777 196 4783 236
rect 4787 196 4789 236
rect 4849 196 4851 236
rect 4855 216 4859 236
rect 4871 216 4873 236
rect 4877 216 4883 236
rect 4887 216 4889 236
rect 4901 216 4903 236
rect 4907 216 4911 236
rect 4915 216 4917 236
rect 4955 216 4957 236
rect 4961 216 4965 236
rect 4977 216 4979 236
rect 4983 216 4989 236
rect 4993 216 4995 236
rect 5007 216 5011 236
rect 5015 216 5021 236
rect 5025 216 5027 236
rect 5039 216 5041 236
rect 4855 196 4868 216
rect 5031 196 5041 216
rect 5045 196 5047 236
rect 5103 196 5105 236
rect 5109 196 5111 236
rect 5123 196 5125 236
rect 5129 208 5131 236
rect 5143 208 5145 236
rect 5129 196 5145 208
rect 5149 196 5151 236
rect 5189 196 5191 236
rect 5195 208 5197 236
rect 5209 208 5211 236
rect 5195 196 5211 208
rect 5215 196 5217 236
rect 5229 196 5231 236
rect 5235 196 5237 236
rect 5291 196 5293 236
rect 5297 196 5303 236
rect 5307 196 5309 236
rect 5369 196 5371 236
rect 5375 216 5379 236
rect 5391 216 5393 236
rect 5397 216 5403 236
rect 5407 216 5409 236
rect 5421 216 5423 236
rect 5427 216 5431 236
rect 5435 216 5437 236
rect 5475 216 5477 236
rect 5481 216 5485 236
rect 5497 216 5499 236
rect 5503 216 5509 236
rect 5513 216 5515 236
rect 5527 216 5531 236
rect 5535 216 5541 236
rect 5545 216 5547 236
rect 5559 216 5561 236
rect 5375 196 5388 216
rect 5551 196 5561 216
rect 5565 196 5567 236
rect 5609 196 5611 236
rect 5615 216 5619 236
rect 5631 216 5633 236
rect 5637 216 5643 236
rect 5647 216 5649 236
rect 5661 216 5663 236
rect 5667 216 5671 236
rect 5675 216 5677 236
rect 5715 216 5717 236
rect 5721 216 5725 236
rect 5737 216 5739 236
rect 5743 216 5749 236
rect 5753 216 5755 236
rect 5767 216 5771 236
rect 5775 216 5781 236
rect 5785 216 5787 236
rect 5799 216 5801 236
rect 5615 196 5628 216
rect 5791 196 5801 216
rect 5805 196 5807 236
rect 5849 196 5851 236
rect 5855 216 5859 236
rect 5871 216 5873 236
rect 5877 216 5883 236
rect 5887 216 5889 236
rect 5901 216 5903 236
rect 5907 216 5911 236
rect 5915 216 5917 236
rect 5955 216 5957 236
rect 5961 216 5965 236
rect 5977 216 5979 236
rect 5983 216 5989 236
rect 5993 216 5995 236
rect 6007 216 6011 236
rect 6015 216 6021 236
rect 6025 216 6027 236
rect 6039 216 6041 236
rect 5855 196 5868 216
rect 6031 196 6041 216
rect 6045 196 6047 236
rect 6103 196 6105 236
rect 6109 196 6111 236
rect 6149 196 6151 236
rect 6155 208 6157 236
rect 6169 208 6171 236
rect 6155 196 6171 208
rect 6175 196 6177 236
rect 6189 196 6191 236
rect 6195 196 6197 236
rect 6263 196 6265 236
rect 6269 224 6285 236
rect 6269 196 6271 224
rect 6283 196 6285 224
rect 6289 196 6291 236
rect 6303 196 6305 236
rect 6309 206 6311 236
rect 6323 206 6325 236
rect 6309 196 6325 206
rect 6329 196 6331 236
rect 6383 216 6385 236
rect 6389 216 6391 236
rect 6429 196 6431 236
rect 6435 216 6439 236
rect 6451 216 6453 236
rect 6457 216 6463 236
rect 6467 216 6469 236
rect 6481 216 6483 236
rect 6487 216 6491 236
rect 6495 216 6497 236
rect 6535 216 6537 236
rect 6541 216 6545 236
rect 6557 216 6559 236
rect 6563 216 6569 236
rect 6573 216 6575 236
rect 6587 216 6591 236
rect 6595 216 6601 236
rect 6605 216 6607 236
rect 6619 216 6621 236
rect 6435 196 6448 216
rect 6611 196 6621 216
rect 6625 196 6627 236
<< pdiffusion >>
rect 33 6264 35 6344
rect 39 6304 48 6344
rect 39 6264 41 6304
rect 53 6264 55 6304
rect 59 6264 69 6304
rect 73 6264 75 6304
rect 87 6264 89 6304
rect 93 6264 101 6304
rect 105 6264 107 6304
rect 119 6264 121 6304
rect 125 6264 127 6304
rect 165 6264 167 6304
rect 171 6264 175 6304
rect 179 6284 190 6304
rect 216 6284 225 6344
rect 179 6264 181 6284
rect 193 6264 195 6284
rect 199 6264 203 6284
rect 207 6264 211 6284
rect 223 6264 225 6284
rect 229 6264 231 6344
rect 288 6264 290 6304
rect 294 6264 298 6304
rect 310 6264 312 6344
rect 316 6264 320 6344
rect 324 6264 326 6344
rect 369 6264 371 6304
rect 375 6264 377 6304
rect 389 6264 391 6304
rect 395 6264 397 6304
rect 463 6264 465 6304
rect 469 6264 471 6304
rect 483 6264 485 6304
rect 489 6264 491 6304
rect 529 6264 531 6304
rect 535 6264 537 6304
rect 549 6264 551 6304
rect 555 6264 557 6304
rect 609 6264 611 6344
rect 615 6284 624 6344
rect 792 6304 801 6344
rect 650 6284 661 6304
rect 615 6264 617 6284
rect 629 6264 633 6284
rect 637 6264 641 6284
rect 645 6264 647 6284
rect 659 6264 661 6284
rect 665 6264 669 6304
rect 673 6264 675 6304
rect 713 6264 715 6304
rect 719 6264 721 6304
rect 733 6264 735 6304
rect 739 6264 747 6304
rect 751 6264 753 6304
rect 765 6264 767 6304
rect 771 6264 781 6304
rect 785 6264 787 6304
rect 799 6264 801 6304
rect 805 6264 807 6344
rect 897 6342 911 6344
rect 849 6264 851 6304
rect 855 6264 857 6304
rect 909 6264 911 6342
rect 915 6330 931 6344
rect 915 6264 917 6330
rect 929 6264 931 6330
rect 935 6342 951 6344
rect 935 6264 937 6342
rect 949 6264 951 6342
rect 955 6276 957 6344
rect 969 6276 971 6344
rect 955 6264 971 6276
rect 975 6264 977 6344
rect 1043 6264 1045 6304
rect 1049 6264 1051 6304
rect 1089 6264 1091 6344
rect 1095 6284 1104 6344
rect 1272 6304 1281 6344
rect 1130 6284 1141 6304
rect 1095 6264 1097 6284
rect 1109 6264 1113 6284
rect 1117 6264 1121 6284
rect 1125 6264 1127 6284
rect 1139 6264 1141 6284
rect 1145 6264 1149 6304
rect 1153 6264 1155 6304
rect 1193 6264 1195 6304
rect 1199 6264 1201 6304
rect 1213 6264 1215 6304
rect 1219 6264 1227 6304
rect 1231 6264 1233 6304
rect 1245 6264 1247 6304
rect 1251 6264 1261 6304
rect 1265 6264 1267 6304
rect 1279 6264 1281 6304
rect 1285 6264 1287 6344
rect 1329 6264 1331 6344
rect 1335 6264 1341 6344
rect 1345 6264 1347 6344
rect 1369 6264 1371 6344
rect 1375 6264 1381 6344
rect 1385 6264 1387 6344
rect 1468 6264 1470 6304
rect 1474 6264 1478 6304
rect 1490 6264 1492 6344
rect 1496 6264 1500 6344
rect 1504 6264 1506 6344
rect 1559 6264 1561 6344
rect 1565 6264 1567 6344
rect 1579 6264 1583 6304
rect 1587 6264 1591 6304
rect 1603 6264 1605 6304
rect 1609 6264 1611 6304
rect 1663 6264 1665 6304
rect 1669 6264 1671 6304
rect 1709 6264 1711 6344
rect 1715 6284 1724 6344
rect 1892 6304 1901 6344
rect 1750 6284 1761 6304
rect 1715 6264 1717 6284
rect 1729 6264 1733 6284
rect 1737 6264 1741 6284
rect 1745 6264 1747 6284
rect 1759 6264 1761 6284
rect 1765 6264 1769 6304
rect 1773 6264 1775 6304
rect 1813 6264 1815 6304
rect 1819 6264 1821 6304
rect 1833 6264 1835 6304
rect 1839 6264 1847 6304
rect 1851 6264 1853 6304
rect 1865 6264 1867 6304
rect 1871 6264 1881 6304
rect 1885 6264 1887 6304
rect 1899 6264 1901 6304
rect 1905 6264 1907 6344
rect 1954 6264 1956 6344
rect 1960 6264 1964 6344
rect 1968 6264 1970 6344
rect 1982 6264 1986 6304
rect 1990 6264 1992 6304
rect 2049 6264 2051 6304
rect 2055 6264 2057 6304
rect 2069 6264 2071 6304
rect 2075 6264 2077 6304
rect 2148 6264 2150 6304
rect 2154 6264 2158 6304
rect 2170 6264 2172 6344
rect 2176 6264 2180 6344
rect 2184 6264 2186 6344
rect 2243 6264 2245 6344
rect 2249 6264 2251 6344
rect 2263 6264 2265 6344
rect 2269 6332 2285 6344
rect 2269 6264 2271 6332
rect 2283 6264 2285 6332
rect 2289 6336 2303 6344
rect 2289 6264 2291 6336
rect 2343 6264 2345 6304
rect 2349 6264 2351 6304
rect 2363 6264 2365 6304
rect 2369 6264 2371 6304
rect 2435 6264 2437 6344
rect 2441 6264 2445 6344
rect 2449 6264 2451 6344
rect 2489 6264 2491 6344
rect 2495 6264 2499 6344
rect 2503 6264 2505 6344
rect 2569 6264 2571 6304
rect 2575 6264 2577 6304
rect 2589 6264 2591 6304
rect 2595 6264 2597 6304
rect 2663 6264 2665 6304
rect 2669 6300 2685 6304
rect 2669 6264 2671 6300
rect 2683 6264 2685 6300
rect 2689 6264 2691 6304
rect 2703 6264 2705 6304
rect 2709 6264 2711 6304
rect 2749 6264 2751 6304
rect 2755 6264 2757 6304
rect 2769 6264 2771 6304
rect 2775 6264 2777 6304
rect 2843 6264 2845 6304
rect 2849 6300 2865 6304
rect 2849 6264 2851 6300
rect 2863 6264 2865 6300
rect 2869 6264 2871 6304
rect 2883 6264 2885 6304
rect 2889 6264 2891 6304
rect 2948 6264 2950 6304
rect 2954 6264 2958 6304
rect 2970 6264 2972 6344
rect 2976 6264 2980 6344
rect 2984 6264 2986 6344
rect 3048 6264 3050 6304
rect 3054 6264 3058 6304
rect 3070 6264 3072 6344
rect 3076 6264 3080 6344
rect 3084 6264 3086 6344
rect 3237 6336 3251 6344
rect 3143 6264 3145 6304
rect 3149 6264 3151 6304
rect 3203 6264 3205 6304
rect 3209 6264 3211 6304
rect 3249 6264 3251 6336
rect 3255 6332 3271 6344
rect 3255 6264 3257 6332
rect 3269 6264 3271 6332
rect 3275 6264 3277 6344
rect 3289 6264 3291 6344
rect 3295 6264 3297 6344
rect 3354 6264 3356 6344
rect 3360 6264 3364 6344
rect 3368 6264 3370 6344
rect 3382 6264 3386 6304
rect 3390 6264 3392 6304
rect 3463 6264 3465 6344
rect 3469 6264 3471 6344
rect 3483 6264 3485 6344
rect 3489 6332 3505 6344
rect 3489 6264 3491 6332
rect 3503 6264 3505 6332
rect 3509 6336 3523 6344
rect 3509 6264 3511 6336
rect 3563 6264 3565 6344
rect 3569 6264 3571 6344
rect 3583 6264 3585 6344
rect 3589 6332 3605 6344
rect 3589 6264 3591 6332
rect 3603 6264 3605 6332
rect 3609 6336 3623 6344
rect 3609 6264 3611 6336
rect 3649 6264 3651 6304
rect 3655 6264 3657 6304
rect 3669 6264 3671 6304
rect 3675 6300 3691 6304
rect 3675 6264 3677 6300
rect 3689 6264 3691 6300
rect 3695 6264 3697 6304
rect 3768 6264 3770 6304
rect 3774 6264 3778 6304
rect 3790 6264 3792 6344
rect 3796 6264 3800 6344
rect 3804 6264 3806 6344
rect 3854 6264 3856 6344
rect 3860 6264 3864 6344
rect 3868 6264 3870 6344
rect 3882 6264 3886 6304
rect 3890 6264 3892 6304
rect 3949 6264 3951 6304
rect 3955 6264 3957 6304
rect 4009 6264 4011 6304
rect 4015 6264 4017 6304
rect 4029 6264 4031 6304
rect 4035 6264 4037 6304
rect 4099 6264 4101 6344
rect 4105 6264 4107 6344
rect 4617 6336 4631 6344
rect 4119 6264 4123 6304
rect 4127 6264 4131 6304
rect 4143 6264 4145 6304
rect 4149 6264 4151 6304
rect 4189 6264 4191 6304
rect 4195 6264 4197 6304
rect 4209 6264 4211 6304
rect 4215 6264 4217 6304
rect 4283 6264 4285 6304
rect 4289 6300 4305 6304
rect 4289 6264 4291 6300
rect 4303 6264 4305 6300
rect 4309 6264 4311 6304
rect 4323 6264 4325 6304
rect 4329 6264 4331 6304
rect 4383 6264 4385 6304
rect 4389 6300 4405 6304
rect 4389 6264 4391 6300
rect 4403 6264 4405 6300
rect 4409 6264 4411 6304
rect 4423 6264 4425 6304
rect 4429 6264 4431 6304
rect 4483 6264 4485 6304
rect 4489 6300 4505 6304
rect 4489 6264 4491 6300
rect 4503 6264 4505 6300
rect 4509 6264 4511 6304
rect 4523 6264 4525 6304
rect 4529 6264 4531 6304
rect 4569 6264 4571 6304
rect 4575 6264 4577 6304
rect 4629 6264 4631 6336
rect 4635 6332 4651 6344
rect 4635 6264 4637 6332
rect 4649 6264 4651 6332
rect 4655 6264 4657 6344
rect 4669 6264 4671 6344
rect 4675 6264 4677 6344
rect 4717 6336 4731 6344
rect 4729 6264 4731 6336
rect 4735 6332 4751 6344
rect 4735 6264 4737 6332
rect 4749 6264 4751 6332
rect 4755 6264 4757 6344
rect 4769 6264 4771 6344
rect 4775 6264 4777 6344
rect 4834 6264 4836 6344
rect 4840 6264 4844 6344
rect 4848 6264 4850 6344
rect 4862 6264 4866 6304
rect 4870 6264 4872 6304
rect 4948 6264 4950 6304
rect 4954 6264 4958 6304
rect 4970 6264 4972 6344
rect 4976 6264 4980 6344
rect 4984 6264 4986 6344
rect 5034 6264 5036 6344
rect 5040 6264 5044 6344
rect 5048 6264 5050 6344
rect 5417 6336 5431 6344
rect 5062 6264 5066 6304
rect 5070 6264 5072 6304
rect 5143 6264 5145 6304
rect 5149 6300 5165 6304
rect 5149 6264 5151 6300
rect 5163 6264 5165 6300
rect 5169 6264 5171 6304
rect 5183 6264 5185 6304
rect 5189 6264 5191 6304
rect 5243 6264 5245 6304
rect 5249 6300 5265 6304
rect 5249 6264 5251 6300
rect 5263 6264 5265 6300
rect 5269 6264 5271 6304
rect 5283 6264 5285 6304
rect 5289 6264 5291 6304
rect 5343 6264 5345 6304
rect 5349 6300 5365 6304
rect 5349 6264 5351 6300
rect 5363 6264 5365 6300
rect 5369 6264 5371 6304
rect 5383 6264 5385 6304
rect 5389 6264 5391 6304
rect 5429 6264 5431 6336
rect 5435 6332 5451 6344
rect 5435 6264 5437 6332
rect 5449 6264 5451 6332
rect 5455 6264 5457 6344
rect 5469 6264 5471 6344
rect 5475 6264 5477 6344
rect 5543 6264 5545 6344
rect 5549 6264 5551 6344
rect 5563 6264 5565 6344
rect 5569 6332 5585 6344
rect 5569 6264 5571 6332
rect 5583 6264 5585 6332
rect 5589 6336 5603 6344
rect 5589 6264 5591 6336
rect 5677 6336 5691 6344
rect 5643 6264 5645 6304
rect 5649 6264 5651 6304
rect 5689 6264 5691 6336
rect 5695 6332 5711 6344
rect 5695 6264 5697 6332
rect 5709 6264 5711 6332
rect 5715 6264 5717 6344
rect 5729 6264 5731 6344
rect 5735 6264 5737 6344
rect 5789 6264 5791 6304
rect 5795 6264 5797 6304
rect 5809 6264 5811 6304
rect 5815 6300 5831 6304
rect 5815 6264 5817 6300
rect 5829 6264 5831 6300
rect 5835 6264 5837 6304
rect 5903 6264 5905 6344
rect 5909 6264 5911 6344
rect 5923 6264 5925 6344
rect 5929 6332 5945 6344
rect 5929 6264 5931 6332
rect 5943 6264 5945 6332
rect 5949 6336 5963 6344
rect 5949 6264 5951 6336
rect 6003 6264 6005 6304
rect 6009 6264 6011 6304
rect 6063 6264 6065 6344
rect 6069 6264 6071 6344
rect 6083 6264 6085 6344
rect 6089 6332 6105 6344
rect 6089 6264 6091 6332
rect 6103 6264 6105 6332
rect 6109 6336 6123 6344
rect 6109 6264 6111 6336
rect 6168 6264 6170 6304
rect 6174 6264 6178 6304
rect 6190 6264 6192 6344
rect 6196 6264 6200 6344
rect 6204 6264 6206 6344
rect 6263 6264 6265 6344
rect 6269 6264 6271 6344
rect 6283 6264 6285 6344
rect 6289 6332 6305 6344
rect 6289 6264 6291 6332
rect 6303 6264 6305 6332
rect 6309 6336 6323 6344
rect 6309 6264 6311 6336
rect 6597 6342 6611 6344
rect 6349 6264 6351 6304
rect 6355 6264 6357 6304
rect 6369 6264 6371 6304
rect 6375 6300 6391 6304
rect 6375 6264 6377 6300
rect 6389 6264 6391 6300
rect 6395 6264 6397 6304
rect 6463 6264 6465 6304
rect 6469 6300 6485 6304
rect 6469 6264 6471 6300
rect 6483 6264 6485 6300
rect 6489 6264 6491 6304
rect 6503 6264 6505 6304
rect 6509 6264 6511 6304
rect 6549 6264 6551 6304
rect 6555 6264 6557 6304
rect 6609 6264 6611 6342
rect 6615 6330 6631 6344
rect 6615 6264 6617 6330
rect 6629 6264 6631 6330
rect 6635 6342 6651 6344
rect 6635 6264 6637 6342
rect 6649 6264 6651 6342
rect 6655 6276 6657 6344
rect 6669 6276 6671 6344
rect 6655 6264 6671 6276
rect 6675 6264 6677 6344
rect 29 6156 31 6236
rect 35 6216 37 6236
rect 49 6216 53 6236
rect 57 6216 61 6236
rect 65 6216 67 6236
rect 79 6216 81 6236
rect 35 6156 44 6216
rect 70 6196 81 6216
rect 85 6196 89 6236
rect 93 6196 95 6236
rect 133 6196 135 6236
rect 139 6196 141 6236
rect 153 6196 155 6236
rect 159 6196 167 6236
rect 171 6196 173 6236
rect 185 6196 187 6236
rect 191 6196 201 6236
rect 205 6196 207 6236
rect 219 6196 221 6236
rect 212 6156 221 6196
rect 225 6156 227 6236
rect 283 6156 285 6236
rect 289 6156 291 6236
rect 303 6156 305 6236
rect 309 6168 311 6236
rect 323 6168 325 6236
rect 309 6156 325 6168
rect 329 6164 331 6236
rect 383 6196 385 6236
rect 389 6196 391 6236
rect 403 6196 405 6236
rect 409 6196 411 6236
rect 329 6156 343 6164
rect 449 6156 451 6236
rect 455 6156 459 6236
rect 463 6156 465 6236
rect 543 6196 545 6236
rect 549 6196 551 6236
rect 563 6196 565 6236
rect 569 6196 571 6236
rect 614 6156 616 6236
rect 620 6156 624 6236
rect 628 6156 630 6236
rect 642 6196 646 6236
rect 650 6196 652 6236
rect 728 6196 730 6236
rect 734 6196 738 6236
rect 750 6156 752 6236
rect 756 6156 760 6236
rect 764 6156 766 6236
rect 809 6156 811 6236
rect 815 6156 819 6236
rect 823 6156 825 6236
rect 903 6156 905 6236
rect 909 6156 911 6236
rect 923 6156 925 6236
rect 929 6168 931 6236
rect 943 6168 945 6236
rect 929 6156 945 6168
rect 949 6164 951 6236
rect 949 6156 963 6164
rect 989 6156 991 6236
rect 995 6156 1001 6236
rect 1005 6157 1007 6236
rect 1019 6157 1021 6236
rect 1005 6156 1021 6157
rect 1025 6157 1027 6236
rect 1103 6196 1105 6236
rect 1109 6196 1111 6236
rect 1025 6156 1039 6157
rect 1149 6156 1151 6236
rect 1155 6156 1159 6236
rect 1163 6156 1165 6236
rect 1248 6196 1250 6236
rect 1254 6196 1258 6236
rect 1270 6156 1272 6236
rect 1276 6156 1280 6236
rect 1284 6156 1286 6236
rect 1343 6196 1345 6236
rect 1349 6196 1351 6236
rect 1403 6196 1405 6236
rect 1409 6196 1411 6236
rect 1449 6156 1451 6236
rect 1455 6156 1459 6236
rect 1463 6156 1465 6236
rect 1529 6156 1531 6236
rect 1535 6156 1539 6236
rect 1543 6156 1545 6236
rect 1609 6196 1611 6236
rect 1615 6196 1617 6236
rect 1669 6156 1671 6236
rect 1675 6156 1679 6236
rect 1683 6156 1685 6236
rect 1749 6156 1751 6236
rect 1755 6156 1759 6236
rect 1763 6156 1765 6236
rect 1834 6156 1836 6236
rect 1840 6156 1844 6236
rect 1848 6156 1850 6236
rect 1862 6196 1866 6236
rect 1870 6196 1872 6236
rect 1929 6196 1931 6236
rect 1935 6196 1937 6236
rect 2003 6156 2005 6236
rect 2009 6156 2011 6236
rect 2023 6156 2025 6236
rect 2029 6168 2031 6236
rect 2043 6168 2045 6236
rect 2029 6156 2045 6168
rect 2049 6164 2051 6236
rect 2089 6196 2091 6236
rect 2095 6196 2097 6236
rect 2168 6196 2170 6236
rect 2174 6196 2178 6236
rect 2049 6156 2063 6164
rect 2190 6156 2192 6236
rect 2196 6156 2200 6236
rect 2204 6156 2206 6236
rect 2249 6196 2251 6236
rect 2255 6196 2257 6236
rect 2328 6196 2330 6236
rect 2334 6196 2338 6236
rect 2350 6156 2352 6236
rect 2356 6156 2360 6236
rect 2364 6156 2366 6236
rect 2423 6196 2425 6236
rect 2429 6200 2431 6236
rect 2443 6200 2445 6236
rect 2429 6196 2445 6200
rect 2449 6196 2451 6236
rect 2463 6196 2465 6236
rect 2469 6196 2471 6236
rect 2523 6156 2525 6236
rect 2529 6156 2531 6236
rect 2543 6156 2545 6236
rect 2549 6168 2551 6236
rect 2563 6168 2565 6236
rect 2549 6156 2565 6168
rect 2569 6164 2571 6236
rect 2569 6156 2583 6164
rect 2635 6156 2637 6236
rect 2641 6156 2645 6236
rect 2649 6156 2651 6236
rect 2703 6196 2705 6236
rect 2709 6200 2711 6236
rect 2723 6200 2725 6236
rect 2709 6196 2725 6200
rect 2729 6196 2731 6236
rect 2743 6196 2745 6236
rect 2749 6196 2751 6236
rect 2803 6156 2805 6236
rect 2809 6224 2825 6236
rect 2809 6156 2811 6224
rect 2823 6156 2825 6224
rect 2829 6158 2831 6236
rect 2843 6158 2845 6236
rect 2829 6156 2845 6158
rect 2849 6170 2851 6236
rect 2863 6170 2865 6236
rect 2849 6156 2865 6170
rect 2869 6158 2871 6236
rect 2923 6196 2925 6236
rect 2929 6196 2931 6236
rect 2969 6196 2971 6236
rect 2975 6196 2977 6236
rect 2989 6196 2991 6236
rect 2995 6200 2997 6236
rect 3009 6200 3011 6236
rect 2995 6196 3011 6200
rect 3015 6196 3017 6236
rect 2869 6156 2883 6158
rect 3083 6156 3085 6236
rect 3089 6156 3091 6236
rect 3103 6156 3105 6236
rect 3109 6168 3111 6236
rect 3123 6168 3125 6236
rect 3109 6156 3125 6168
rect 3129 6164 3131 6236
rect 3183 6196 3185 6236
rect 3189 6200 3191 6236
rect 3203 6200 3205 6236
rect 3189 6196 3205 6200
rect 3209 6196 3211 6236
rect 3223 6196 3225 6236
rect 3229 6196 3231 6236
rect 3129 6156 3143 6164
rect 3283 6156 3285 6236
rect 3289 6156 3291 6236
rect 3303 6156 3305 6236
rect 3309 6168 3311 6236
rect 3323 6168 3325 6236
rect 3309 6156 3325 6168
rect 3329 6164 3331 6236
rect 3383 6196 3385 6236
rect 3389 6196 3391 6236
rect 3443 6196 3445 6236
rect 3449 6200 3451 6236
rect 3463 6200 3465 6236
rect 3449 6196 3465 6200
rect 3469 6196 3471 6236
rect 3483 6196 3485 6236
rect 3489 6196 3491 6236
rect 3529 6196 3531 6236
rect 3535 6196 3537 6236
rect 3549 6196 3551 6236
rect 3555 6200 3557 6236
rect 3569 6200 3571 6236
rect 3555 6196 3571 6200
rect 3575 6196 3577 6236
rect 3629 6196 3631 6236
rect 3635 6196 3637 6236
rect 3329 6156 3343 6164
rect 3689 6164 3691 6236
rect 3677 6156 3691 6164
rect 3695 6168 3697 6236
rect 3709 6168 3711 6236
rect 3695 6156 3711 6168
rect 3715 6156 3717 6236
rect 3729 6156 3731 6236
rect 3735 6156 3737 6236
rect 3803 6196 3805 6236
rect 3809 6196 3811 6236
rect 3823 6196 3825 6236
rect 3829 6196 3831 6236
rect 3869 6196 3871 6236
rect 3875 6196 3877 6236
rect 3889 6196 3891 6236
rect 3895 6196 3897 6236
rect 3968 6196 3970 6236
rect 3974 6196 3978 6236
rect 3990 6156 3992 6236
rect 3996 6156 4000 6236
rect 4004 6156 4006 6236
rect 4054 6156 4056 6236
rect 4060 6156 4064 6236
rect 4068 6156 4070 6236
rect 4082 6196 4086 6236
rect 4090 6196 4092 6236
rect 4175 6156 4177 6236
rect 4181 6156 4185 6236
rect 4189 6156 4191 6236
rect 4229 6196 4231 6236
rect 4235 6196 4237 6236
rect 4303 6196 4305 6236
rect 4309 6196 4311 6236
rect 4323 6196 4325 6236
rect 4329 6196 4331 6236
rect 4369 6196 4371 6236
rect 4375 6196 4377 6236
rect 4389 6196 4393 6236
rect 4397 6196 4401 6236
rect 4413 6156 4415 6236
rect 4419 6156 4421 6236
rect 4488 6196 4490 6236
rect 4494 6196 4498 6236
rect 4510 6156 4512 6236
rect 4516 6156 4520 6236
rect 4524 6156 4526 6236
rect 4583 6156 4585 6236
rect 4589 6156 4591 6236
rect 4603 6156 4605 6236
rect 4609 6168 4611 6236
rect 4623 6168 4625 6236
rect 4609 6156 4625 6168
rect 4629 6164 4631 6236
rect 4669 6196 4671 6236
rect 4675 6196 4677 6236
rect 4689 6196 4691 6236
rect 4695 6200 4697 6236
rect 4709 6200 4711 6236
rect 4695 6196 4711 6200
rect 4715 6196 4717 6236
rect 4629 6156 4643 6164
rect 4783 6156 4785 6236
rect 4789 6156 4791 6236
rect 4803 6156 4805 6236
rect 4809 6168 4811 6236
rect 4823 6168 4825 6236
rect 4809 6156 4825 6168
rect 4829 6164 4831 6236
rect 4883 6196 4885 6236
rect 4889 6200 4891 6236
rect 4903 6200 4905 6236
rect 4889 6196 4905 6200
rect 4909 6196 4911 6236
rect 4923 6196 4925 6236
rect 4929 6196 4931 6236
rect 4969 6196 4971 6236
rect 4975 6196 4977 6236
rect 4989 6196 4991 6236
rect 4995 6200 4997 6236
rect 5009 6200 5011 6236
rect 4995 6196 5011 6200
rect 5015 6196 5017 6236
rect 5088 6196 5090 6236
rect 5094 6196 5098 6236
rect 4829 6156 4843 6164
rect 5110 6156 5112 6236
rect 5116 6156 5120 6236
rect 5124 6156 5126 6236
rect 5183 6196 5185 6236
rect 5189 6196 5191 6236
rect 5203 6196 5205 6236
rect 5209 6196 5211 6236
rect 5249 6196 5251 6236
rect 5255 6196 5257 6236
rect 5269 6196 5273 6236
rect 5277 6196 5281 6236
rect 5293 6156 5295 6236
rect 5299 6156 5301 6236
rect 5354 6156 5356 6236
rect 5360 6156 5364 6236
rect 5368 6156 5370 6236
rect 5382 6196 5386 6236
rect 5390 6196 5392 6236
rect 5463 6156 5465 6236
rect 5469 6156 5471 6236
rect 5483 6156 5485 6236
rect 5489 6168 5491 6236
rect 5503 6168 5505 6236
rect 5489 6156 5505 6168
rect 5509 6164 5511 6236
rect 5563 6196 5565 6236
rect 5569 6200 5571 6236
rect 5583 6200 5585 6236
rect 5569 6196 5585 6200
rect 5589 6196 5591 6236
rect 5603 6196 5605 6236
rect 5609 6196 5611 6236
rect 5649 6196 5651 6236
rect 5655 6196 5657 6236
rect 5669 6196 5671 6236
rect 5675 6200 5677 6236
rect 5689 6200 5691 6236
rect 5675 6196 5691 6200
rect 5695 6196 5697 6236
rect 5509 6156 5523 6164
rect 5763 6156 5765 6236
rect 5769 6156 5771 6236
rect 5783 6156 5785 6236
rect 5789 6168 5791 6236
rect 5803 6168 5805 6236
rect 5789 6156 5805 6168
rect 5809 6164 5811 6236
rect 5849 6196 5851 6236
rect 5855 6196 5857 6236
rect 5869 6196 5871 6236
rect 5875 6200 5877 6236
rect 5889 6200 5891 6236
rect 5875 6196 5891 6200
rect 5895 6196 5897 6236
rect 5809 6156 5823 6164
rect 5954 6156 5956 6236
rect 5960 6156 5964 6236
rect 5968 6156 5970 6236
rect 5982 6196 5986 6236
rect 5990 6196 5992 6236
rect 6054 6156 6056 6236
rect 6060 6156 6064 6236
rect 6068 6156 6070 6236
rect 6082 6196 6086 6236
rect 6090 6196 6092 6236
rect 6149 6196 6151 6236
rect 6155 6196 6157 6236
rect 6169 6196 6171 6236
rect 6175 6200 6177 6236
rect 6189 6200 6191 6236
rect 6175 6196 6191 6200
rect 6195 6196 6197 6236
rect 6249 6196 6251 6236
rect 6255 6196 6257 6236
rect 6269 6196 6271 6236
rect 6275 6200 6277 6236
rect 6289 6200 6291 6236
rect 6275 6196 6291 6200
rect 6295 6196 6297 6236
rect 6363 6196 6365 6236
rect 6369 6200 6371 6236
rect 6383 6200 6385 6236
rect 6369 6196 6385 6200
rect 6389 6196 6391 6236
rect 6403 6196 6405 6236
rect 6409 6196 6411 6236
rect 6463 6156 6465 6236
rect 6469 6156 6471 6236
rect 6483 6156 6485 6236
rect 6489 6168 6491 6236
rect 6503 6168 6505 6236
rect 6489 6156 6505 6168
rect 6509 6164 6511 6236
rect 6549 6196 6551 6236
rect 6555 6196 6557 6236
rect 6609 6196 6611 6236
rect 6615 6196 6617 6236
rect 6509 6156 6523 6164
rect 41 5784 43 5864
rect 47 5784 49 5864
rect 61 5784 65 5824
rect 69 5784 71 5824
rect 109 5784 111 5824
rect 115 5784 117 5824
rect 129 5784 131 5824
rect 135 5784 137 5824
rect 189 5784 191 5824
rect 195 5784 197 5824
rect 209 5784 211 5824
rect 215 5784 217 5824
rect 283 5784 285 5864
rect 289 5784 291 5864
rect 303 5784 305 5864
rect 309 5852 325 5864
rect 309 5784 311 5852
rect 323 5784 325 5852
rect 329 5856 343 5864
rect 329 5784 331 5856
rect 383 5784 385 5824
rect 389 5784 391 5824
rect 403 5784 405 5824
rect 409 5784 411 5824
rect 449 5784 451 5824
rect 455 5784 457 5824
rect 535 5784 537 5864
rect 541 5784 545 5864
rect 549 5784 551 5864
rect 589 5784 591 5864
rect 595 5784 599 5864
rect 603 5784 605 5864
rect 674 5784 676 5864
rect 680 5784 684 5864
rect 688 5784 690 5864
rect 702 5784 706 5824
rect 710 5784 712 5824
rect 783 5784 785 5824
rect 789 5784 791 5824
rect 829 5784 831 5864
rect 835 5784 839 5864
rect 843 5784 845 5864
rect 923 5784 925 5824
rect 929 5784 931 5824
rect 943 5784 945 5824
rect 949 5784 951 5824
rect 1008 5784 1010 5824
rect 1014 5784 1018 5824
rect 1030 5784 1032 5864
rect 1036 5784 1040 5864
rect 1044 5784 1046 5864
rect 1089 5784 1091 5864
rect 1095 5784 1099 5864
rect 1103 5784 1105 5864
rect 1183 5784 1185 5824
rect 1189 5784 1191 5824
rect 1229 5784 1231 5864
rect 1235 5804 1244 5864
rect 1412 5824 1421 5864
rect 1270 5804 1281 5824
rect 1235 5784 1237 5804
rect 1249 5784 1253 5804
rect 1257 5784 1261 5804
rect 1265 5784 1267 5804
rect 1279 5784 1281 5804
rect 1285 5784 1289 5824
rect 1293 5784 1295 5824
rect 1333 5784 1335 5824
rect 1339 5784 1341 5824
rect 1353 5784 1355 5824
rect 1359 5784 1367 5824
rect 1371 5784 1373 5824
rect 1385 5784 1387 5824
rect 1391 5784 1401 5824
rect 1405 5784 1407 5824
rect 1419 5784 1421 5824
rect 1425 5784 1427 5864
rect 1469 5784 1471 5824
rect 1475 5784 1477 5824
rect 1489 5784 1491 5824
rect 1495 5784 1497 5824
rect 1563 5784 1565 5824
rect 1569 5820 1585 5824
rect 1569 5784 1571 5820
rect 1583 5784 1585 5820
rect 1589 5784 1591 5824
rect 1603 5784 1605 5824
rect 1609 5784 1611 5824
rect 1668 5784 1670 5824
rect 1674 5784 1678 5824
rect 1690 5784 1692 5864
rect 1696 5784 1700 5864
rect 1704 5784 1706 5864
rect 1775 5784 1777 5864
rect 1781 5784 1785 5864
rect 1789 5784 1791 5864
rect 1843 5784 1845 5824
rect 1849 5820 1865 5824
rect 1849 5784 1851 5820
rect 1863 5784 1865 5820
rect 1869 5784 1871 5824
rect 1883 5784 1885 5824
rect 1889 5784 1891 5824
rect 1929 5784 1931 5824
rect 1935 5784 1937 5824
rect 2008 5784 2010 5824
rect 2014 5784 2018 5824
rect 2030 5784 2032 5864
rect 2036 5784 2040 5864
rect 2044 5784 2046 5864
rect 2089 5784 2091 5824
rect 2095 5784 2097 5824
rect 2109 5784 2111 5824
rect 2115 5820 2131 5824
rect 2115 5784 2117 5820
rect 2129 5784 2131 5820
rect 2135 5784 2137 5824
rect 2203 5784 2205 5864
rect 2209 5784 2211 5864
rect 2223 5784 2225 5864
rect 2229 5852 2245 5864
rect 2229 5784 2231 5852
rect 2243 5784 2245 5852
rect 2249 5856 2263 5864
rect 2249 5784 2251 5856
rect 2294 5784 2296 5864
rect 2300 5784 2304 5864
rect 2308 5784 2310 5864
rect 2322 5784 2326 5824
rect 2330 5784 2332 5824
rect 2403 5784 2405 5824
rect 2409 5784 2411 5824
rect 2423 5784 2425 5824
rect 2429 5784 2431 5824
rect 2483 5784 2485 5824
rect 2489 5820 2505 5824
rect 2489 5784 2491 5820
rect 2503 5784 2505 5820
rect 2509 5784 2511 5824
rect 2523 5784 2525 5824
rect 2529 5784 2531 5824
rect 2583 5784 2585 5864
rect 2589 5784 2591 5864
rect 2603 5784 2605 5864
rect 2609 5852 2625 5864
rect 2609 5784 2611 5852
rect 2623 5784 2625 5852
rect 2629 5856 2643 5864
rect 2629 5784 2631 5856
rect 2669 5784 2671 5824
rect 2675 5784 2677 5824
rect 2689 5784 2691 5824
rect 2695 5784 2697 5824
rect 2763 5784 2765 5824
rect 2769 5820 2785 5824
rect 2769 5784 2771 5820
rect 2783 5784 2785 5820
rect 2789 5784 2791 5824
rect 2803 5784 2805 5824
rect 2809 5784 2811 5824
rect 2863 5784 2865 5824
rect 2869 5820 2885 5824
rect 2869 5784 2871 5820
rect 2883 5784 2885 5820
rect 2889 5784 2891 5824
rect 2903 5784 2905 5824
rect 2909 5784 2911 5824
rect 2963 5784 2965 5824
rect 2969 5820 2985 5824
rect 2969 5784 2971 5820
rect 2983 5784 2985 5820
rect 2989 5784 2991 5824
rect 3003 5784 3005 5824
rect 3009 5784 3011 5824
rect 3063 5784 3065 5824
rect 3069 5820 3085 5824
rect 3069 5784 3071 5820
rect 3083 5784 3085 5820
rect 3089 5784 3091 5824
rect 3103 5784 3105 5824
rect 3109 5784 3111 5824
rect 3149 5784 3151 5824
rect 3155 5784 3157 5824
rect 3169 5784 3171 5824
rect 3175 5820 3191 5824
rect 3175 5784 3177 5820
rect 3189 5784 3191 5820
rect 3195 5784 3197 5824
rect 3268 5784 3270 5824
rect 3274 5784 3278 5824
rect 3290 5784 3292 5864
rect 3296 5784 3300 5864
rect 3304 5784 3306 5864
rect 3354 5784 3356 5864
rect 3360 5784 3364 5864
rect 3368 5784 3370 5864
rect 3382 5784 3386 5824
rect 3390 5784 3392 5824
rect 3463 5784 3465 5864
rect 3469 5784 3471 5864
rect 3483 5784 3485 5864
rect 3489 5852 3505 5864
rect 3489 5784 3491 5852
rect 3503 5784 3505 5852
rect 3509 5856 3523 5864
rect 3509 5784 3511 5856
rect 3568 5784 3570 5824
rect 3574 5784 3578 5824
rect 3590 5784 3592 5864
rect 3596 5784 3600 5864
rect 3604 5784 3606 5864
rect 3737 5856 3751 5864
rect 3663 5784 3665 5824
rect 3669 5820 3685 5824
rect 3669 5784 3671 5820
rect 3683 5784 3685 5820
rect 3689 5784 3691 5824
rect 3703 5784 3705 5824
rect 3709 5784 3711 5824
rect 3749 5784 3751 5856
rect 3755 5852 3771 5864
rect 3755 5784 3757 5852
rect 3769 5784 3771 5852
rect 3775 5784 3777 5864
rect 3789 5784 3791 5864
rect 3795 5784 3797 5864
rect 3863 5784 3865 5824
rect 3869 5820 3885 5824
rect 3869 5784 3871 5820
rect 3883 5784 3885 5820
rect 3889 5784 3891 5824
rect 3903 5784 3905 5824
rect 3909 5784 3911 5824
rect 3963 5784 3965 5864
rect 3969 5784 3971 5864
rect 3983 5784 3985 5864
rect 3989 5852 4005 5864
rect 3989 5784 3991 5852
rect 4003 5784 4005 5852
rect 4009 5856 4023 5864
rect 4009 5784 4011 5856
rect 4063 5784 4065 5824
rect 4069 5820 4085 5824
rect 4069 5784 4071 5820
rect 4083 5784 4085 5820
rect 4089 5784 4091 5824
rect 4103 5784 4105 5824
rect 4109 5784 4111 5824
rect 4163 5784 4165 5864
rect 4169 5784 4171 5864
rect 4183 5784 4185 5864
rect 4189 5852 4205 5864
rect 4189 5784 4191 5852
rect 4203 5784 4205 5852
rect 4209 5856 4223 5864
rect 4209 5784 4211 5856
rect 4249 5784 4251 5824
rect 4255 5784 4257 5824
rect 4269 5784 4271 5824
rect 4275 5820 4291 5824
rect 4275 5784 4277 5820
rect 4289 5784 4291 5820
rect 4295 5784 4297 5824
rect 4349 5784 4351 5824
rect 4355 5784 4357 5824
rect 4369 5784 4371 5824
rect 4375 5784 4377 5824
rect 4448 5784 4450 5824
rect 4454 5784 4458 5824
rect 4470 5784 4472 5864
rect 4476 5784 4480 5864
rect 4484 5784 4486 5864
rect 4555 5784 4557 5864
rect 4561 5784 4565 5864
rect 4569 5784 4571 5864
rect 4609 5784 4611 5824
rect 4615 5784 4617 5824
rect 4629 5784 4633 5824
rect 4637 5784 4641 5824
rect 4653 5784 4655 5864
rect 4659 5784 4661 5864
rect 4723 5784 4725 5864
rect 4729 5784 4731 5864
rect 4743 5784 4745 5864
rect 4749 5852 4765 5864
rect 4749 5784 4751 5852
rect 4763 5784 4765 5852
rect 4769 5856 4783 5864
rect 4769 5784 4771 5856
rect 5037 5856 5051 5864
rect 4809 5784 4811 5824
rect 4815 5784 4817 5824
rect 4829 5784 4831 5824
rect 4835 5784 4837 5824
rect 4903 5784 4905 5824
rect 4909 5784 4911 5824
rect 4963 5784 4965 5824
rect 4969 5820 4985 5824
rect 4969 5784 4971 5820
rect 4983 5784 4985 5820
rect 4989 5784 4991 5824
rect 5003 5784 5005 5824
rect 5009 5784 5011 5824
rect 5049 5784 5051 5856
rect 5055 5852 5071 5864
rect 5055 5784 5057 5852
rect 5069 5784 5071 5852
rect 5075 5784 5077 5864
rect 5089 5784 5091 5864
rect 5095 5784 5097 5864
rect 5154 5784 5156 5864
rect 5160 5784 5164 5864
rect 5168 5784 5170 5864
rect 5182 5784 5186 5824
rect 5190 5784 5192 5824
rect 5254 5784 5256 5864
rect 5260 5784 5264 5864
rect 5268 5784 5270 5864
rect 5337 5862 5351 5864
rect 5282 5784 5286 5824
rect 5290 5784 5292 5824
rect 5349 5784 5351 5862
rect 5355 5850 5371 5864
rect 5355 5784 5357 5850
rect 5369 5784 5371 5850
rect 5375 5862 5391 5864
rect 5375 5784 5377 5862
rect 5389 5784 5391 5862
rect 5395 5796 5397 5864
rect 5409 5796 5411 5864
rect 5395 5784 5411 5796
rect 5415 5784 5417 5864
rect 5697 5856 5711 5864
rect 5483 5784 5485 5824
rect 5489 5784 5491 5824
rect 5503 5784 5505 5824
rect 5509 5784 5511 5824
rect 5549 5784 5551 5824
rect 5555 5784 5557 5824
rect 5623 5784 5625 5824
rect 5629 5820 5645 5824
rect 5629 5784 5631 5820
rect 5643 5784 5645 5820
rect 5649 5784 5651 5824
rect 5663 5784 5665 5824
rect 5669 5784 5671 5824
rect 5709 5784 5711 5856
rect 5715 5852 5731 5864
rect 5715 5784 5717 5852
rect 5729 5784 5731 5852
rect 5735 5784 5737 5864
rect 5749 5784 5751 5864
rect 5755 5784 5757 5864
rect 5828 5784 5830 5824
rect 5834 5784 5838 5824
rect 5850 5784 5852 5864
rect 5856 5784 5860 5864
rect 5864 5784 5866 5864
rect 5914 5784 5916 5864
rect 5920 5784 5924 5864
rect 5928 5784 5930 5864
rect 5942 5784 5946 5824
rect 5950 5784 5952 5824
rect 6028 5784 6030 5824
rect 6034 5784 6038 5824
rect 6050 5784 6052 5864
rect 6056 5784 6060 5864
rect 6064 5784 6066 5864
rect 6097 5862 6111 5864
rect 6109 5784 6111 5862
rect 6115 5850 6131 5864
rect 6115 5784 6117 5850
rect 6129 5784 6131 5850
rect 6135 5862 6151 5864
rect 6135 5784 6137 5862
rect 6149 5784 6151 5862
rect 6155 5796 6157 5864
rect 6169 5796 6171 5864
rect 6155 5784 6171 5796
rect 6175 5784 6177 5864
rect 6243 5784 6245 5824
rect 6249 5784 6251 5824
rect 6263 5784 6265 5824
rect 6269 5784 6271 5824
rect 6309 5784 6311 5824
rect 6315 5784 6317 5824
rect 6329 5784 6333 5824
rect 6337 5784 6341 5824
rect 6353 5784 6355 5864
rect 6359 5784 6361 5864
rect 6414 5784 6416 5864
rect 6420 5784 6424 5864
rect 6428 5784 6430 5864
rect 6442 5784 6446 5824
rect 6450 5784 6452 5824
rect 6509 5784 6511 5824
rect 6515 5784 6517 5824
rect 6529 5784 6531 5824
rect 6535 5820 6551 5824
rect 6535 5784 6537 5820
rect 6549 5784 6551 5820
rect 6555 5784 6557 5824
rect 6609 5784 6611 5824
rect 6615 5784 6617 5824
rect 6629 5784 6631 5824
rect 6635 5784 6637 5824
rect 41 5676 43 5756
rect 47 5676 49 5756
rect 61 5716 65 5756
rect 69 5716 71 5756
rect 121 5676 123 5756
rect 127 5676 129 5756
rect 141 5716 145 5756
rect 149 5716 151 5756
rect 189 5676 191 5756
rect 195 5736 197 5756
rect 209 5736 213 5756
rect 217 5736 221 5756
rect 225 5736 227 5756
rect 239 5736 241 5756
rect 195 5676 204 5736
rect 230 5716 241 5736
rect 245 5716 249 5756
rect 253 5716 255 5756
rect 293 5716 295 5756
rect 299 5716 301 5756
rect 313 5716 315 5756
rect 319 5716 327 5756
rect 331 5716 333 5756
rect 345 5716 347 5756
rect 351 5716 361 5756
rect 365 5716 367 5756
rect 379 5716 381 5756
rect 372 5676 381 5716
rect 385 5676 387 5756
rect 455 5676 457 5756
rect 461 5676 465 5756
rect 469 5676 471 5756
rect 509 5684 511 5756
rect 497 5676 511 5684
rect 515 5688 517 5756
rect 529 5688 531 5756
rect 515 5676 531 5688
rect 535 5676 537 5756
rect 549 5676 551 5756
rect 555 5676 557 5756
rect 609 5716 611 5756
rect 615 5716 617 5756
rect 629 5716 631 5756
rect 635 5716 637 5756
rect 689 5716 691 5756
rect 695 5716 697 5756
rect 709 5716 713 5756
rect 717 5716 721 5756
rect 733 5676 735 5756
rect 739 5676 741 5756
rect 789 5716 791 5756
rect 795 5716 797 5756
rect 809 5716 811 5756
rect 815 5716 817 5756
rect 869 5716 871 5756
rect 875 5716 877 5756
rect 889 5716 891 5756
rect 895 5716 897 5756
rect 949 5676 951 5756
rect 955 5676 959 5756
rect 963 5676 965 5756
rect 1029 5716 1031 5756
rect 1035 5716 1037 5756
rect 1089 5676 1091 5756
rect 1095 5676 1101 5756
rect 1105 5677 1107 5756
rect 1119 5677 1121 5756
rect 1105 5676 1121 5677
rect 1125 5677 1127 5756
rect 1125 5676 1139 5677
rect 1189 5676 1191 5756
rect 1195 5676 1199 5756
rect 1203 5676 1205 5756
rect 1269 5716 1271 5756
rect 1275 5716 1277 5756
rect 1329 5676 1331 5756
rect 1335 5676 1339 5756
rect 1343 5676 1345 5756
rect 1409 5716 1411 5756
rect 1415 5716 1417 5756
rect 1469 5676 1471 5756
rect 1475 5736 1477 5756
rect 1489 5736 1493 5756
rect 1497 5736 1501 5756
rect 1505 5736 1507 5756
rect 1519 5736 1521 5756
rect 1475 5676 1484 5736
rect 1510 5716 1521 5736
rect 1525 5716 1529 5756
rect 1533 5716 1535 5756
rect 1573 5716 1575 5756
rect 1579 5716 1581 5756
rect 1593 5716 1595 5756
rect 1599 5716 1607 5756
rect 1611 5716 1613 5756
rect 1625 5716 1627 5756
rect 1631 5716 1641 5756
rect 1645 5716 1647 5756
rect 1659 5716 1661 5756
rect 1652 5676 1661 5716
rect 1665 5676 1667 5756
rect 1709 5676 1711 5756
rect 1715 5676 1721 5756
rect 1725 5676 1727 5756
rect 1749 5676 1751 5756
rect 1755 5676 1761 5756
rect 1765 5676 1767 5756
rect 1848 5716 1850 5756
rect 1854 5716 1858 5756
rect 1870 5676 1872 5756
rect 1876 5676 1880 5756
rect 1884 5676 1886 5756
rect 1943 5716 1945 5756
rect 1949 5716 1951 5756
rect 1963 5716 1965 5756
rect 1969 5716 1971 5756
rect 2009 5716 2011 5756
rect 2015 5716 2017 5756
rect 2083 5676 2085 5756
rect 2089 5676 2091 5756
rect 2103 5676 2105 5756
rect 2109 5688 2111 5756
rect 2123 5688 2125 5756
rect 2109 5676 2125 5688
rect 2129 5684 2131 5756
rect 2129 5676 2143 5684
rect 2169 5676 2171 5756
rect 2175 5676 2179 5756
rect 2183 5676 2185 5756
rect 2249 5716 2251 5756
rect 2255 5716 2257 5756
rect 2269 5716 2271 5756
rect 2275 5716 2277 5756
rect 2339 5688 2341 5748
rect 2345 5744 2361 5748
rect 2345 5692 2347 5744
rect 2359 5692 2361 5744
rect 2345 5688 2361 5692
rect 2365 5688 2367 5748
rect 2403 5698 2405 5756
rect 2391 5696 2405 5698
rect 2409 5744 2425 5756
rect 2409 5696 2411 5744
rect 2423 5696 2425 5744
rect 2429 5696 2431 5756
rect 2443 5696 2445 5756
rect 2449 5696 2451 5756
rect 2463 5696 2465 5756
rect 2469 5696 2471 5756
rect 2523 5716 2525 5756
rect 2529 5716 2531 5756
rect 2543 5716 2545 5756
rect 2549 5716 2551 5756
rect 2603 5716 2605 5756
rect 2609 5720 2611 5756
rect 2623 5720 2625 5756
rect 2609 5716 2625 5720
rect 2629 5716 2631 5756
rect 2643 5716 2645 5756
rect 2649 5716 2651 5756
rect 2703 5716 2705 5756
rect 2709 5720 2711 5756
rect 2723 5720 2725 5756
rect 2709 5716 2725 5720
rect 2729 5716 2731 5756
rect 2743 5716 2745 5756
rect 2749 5716 2751 5756
rect 2789 5716 2791 5756
rect 2795 5716 2797 5756
rect 2809 5716 2811 5756
rect 2815 5716 2817 5756
rect 2874 5676 2876 5756
rect 2880 5676 2884 5756
rect 2888 5676 2890 5756
rect 2902 5716 2906 5756
rect 2910 5716 2912 5756
rect 2983 5716 2985 5756
rect 2989 5720 2991 5756
rect 3003 5720 3005 5756
rect 2989 5716 3005 5720
rect 3009 5716 3011 5756
rect 3023 5716 3025 5756
rect 3029 5716 3031 5756
rect 3069 5684 3071 5756
rect 3057 5676 3071 5684
rect 3075 5688 3077 5756
rect 3089 5688 3091 5756
rect 3075 5676 3091 5688
rect 3095 5676 3097 5756
rect 3109 5676 3111 5756
rect 3115 5676 3117 5756
rect 3188 5716 3190 5756
rect 3194 5716 3198 5756
rect 3210 5676 3212 5756
rect 3216 5676 3220 5756
rect 3224 5676 3226 5756
rect 3283 5716 3285 5756
rect 3289 5716 3291 5756
rect 3329 5716 3331 5756
rect 3335 5716 3337 5756
rect 3349 5716 3351 5756
rect 3355 5720 3357 5756
rect 3369 5720 3371 5756
rect 3355 5716 3371 5720
rect 3375 5716 3377 5756
rect 3443 5716 3445 5756
rect 3449 5720 3451 5756
rect 3463 5720 3465 5756
rect 3449 5716 3465 5720
rect 3469 5716 3471 5756
rect 3483 5716 3485 5756
rect 3489 5716 3491 5756
rect 3543 5716 3545 5756
rect 3549 5720 3551 5756
rect 3563 5720 3565 5756
rect 3549 5716 3565 5720
rect 3569 5716 3571 5756
rect 3583 5716 3585 5756
rect 3589 5716 3591 5756
rect 3643 5716 3645 5756
rect 3649 5716 3651 5756
rect 3708 5716 3710 5756
rect 3714 5716 3718 5756
rect 3730 5676 3732 5756
rect 3736 5676 3740 5756
rect 3744 5676 3746 5756
rect 3815 5676 3817 5756
rect 3821 5676 3825 5756
rect 3829 5676 3831 5756
rect 3874 5676 3876 5756
rect 3880 5676 3884 5756
rect 3888 5676 3890 5756
rect 3902 5716 3906 5756
rect 3910 5716 3912 5756
rect 3983 5716 3985 5756
rect 3989 5716 3991 5756
rect 4043 5676 4045 5756
rect 4049 5744 4065 5756
rect 4049 5676 4051 5744
rect 4063 5676 4065 5744
rect 4069 5678 4071 5756
rect 4083 5678 4085 5756
rect 4069 5676 4085 5678
rect 4089 5690 4091 5756
rect 4103 5690 4105 5756
rect 4089 5676 4105 5690
rect 4109 5678 4111 5756
rect 4168 5716 4170 5756
rect 4174 5716 4178 5756
rect 4109 5676 4123 5678
rect 4190 5676 4192 5756
rect 4196 5676 4200 5756
rect 4204 5676 4206 5756
rect 4263 5716 4265 5756
rect 4269 5720 4271 5756
rect 4283 5720 4285 5756
rect 4269 5716 4285 5720
rect 4289 5716 4291 5756
rect 4303 5716 4305 5756
rect 4309 5716 4311 5756
rect 4349 5716 4351 5756
rect 4355 5716 4357 5756
rect 4428 5716 4430 5756
rect 4434 5716 4438 5756
rect 4450 5676 4452 5756
rect 4456 5676 4460 5756
rect 4464 5676 4466 5756
rect 4519 5676 4521 5756
rect 4525 5676 4527 5756
rect 4539 5716 4543 5756
rect 4547 5716 4551 5756
rect 4563 5716 4565 5756
rect 4569 5716 4571 5756
rect 4609 5716 4611 5756
rect 4615 5716 4617 5756
rect 4629 5716 4631 5756
rect 4635 5716 4637 5756
rect 4708 5716 4710 5756
rect 4714 5716 4718 5756
rect 4730 5676 4732 5756
rect 4736 5676 4740 5756
rect 4744 5676 4746 5756
rect 4794 5676 4796 5756
rect 4800 5676 4804 5756
rect 4808 5676 4810 5756
rect 4822 5716 4826 5756
rect 4830 5716 4832 5756
rect 4903 5716 4905 5756
rect 4909 5720 4911 5756
rect 4923 5720 4925 5756
rect 4909 5716 4925 5720
rect 4929 5716 4931 5756
rect 4943 5716 4945 5756
rect 4949 5716 4951 5756
rect 4989 5684 4991 5756
rect 4977 5676 4991 5684
rect 4995 5688 4997 5756
rect 5009 5688 5011 5756
rect 4995 5676 5011 5688
rect 5015 5676 5017 5756
rect 5029 5676 5031 5756
rect 5035 5676 5037 5756
rect 5094 5676 5096 5756
rect 5100 5676 5104 5756
rect 5108 5676 5110 5756
rect 5122 5716 5126 5756
rect 5130 5716 5132 5756
rect 5189 5716 5191 5756
rect 5195 5716 5197 5756
rect 5209 5716 5211 5756
rect 5215 5720 5217 5756
rect 5229 5720 5231 5756
rect 5215 5716 5231 5720
rect 5235 5716 5237 5756
rect 5289 5716 5291 5756
rect 5295 5716 5297 5756
rect 5309 5716 5311 5756
rect 5315 5716 5317 5756
rect 5369 5716 5371 5756
rect 5375 5716 5377 5756
rect 5389 5716 5391 5756
rect 5395 5720 5397 5756
rect 5409 5720 5411 5756
rect 5395 5716 5411 5720
rect 5415 5716 5417 5756
rect 5469 5684 5471 5756
rect 5457 5676 5471 5684
rect 5475 5688 5477 5756
rect 5489 5688 5491 5756
rect 5475 5676 5491 5688
rect 5495 5676 5497 5756
rect 5509 5676 5511 5756
rect 5515 5676 5517 5756
rect 5569 5716 5571 5756
rect 5575 5716 5577 5756
rect 5589 5716 5591 5756
rect 5595 5716 5597 5756
rect 5663 5716 5665 5756
rect 5669 5716 5671 5756
rect 5683 5716 5685 5756
rect 5689 5716 5691 5756
rect 5729 5678 5731 5756
rect 5717 5676 5731 5678
rect 5735 5690 5737 5756
rect 5749 5690 5751 5756
rect 5735 5676 5751 5690
rect 5755 5678 5757 5756
rect 5769 5678 5771 5756
rect 5755 5676 5771 5678
rect 5775 5744 5791 5756
rect 5775 5676 5777 5744
rect 5789 5676 5791 5744
rect 5795 5676 5797 5756
rect 5868 5716 5870 5756
rect 5874 5716 5878 5756
rect 5890 5676 5892 5756
rect 5896 5676 5900 5756
rect 5904 5676 5906 5756
rect 5949 5716 5951 5756
rect 5955 5716 5957 5756
rect 6009 5678 6011 5756
rect 5997 5676 6011 5678
rect 6015 5690 6017 5756
rect 6029 5690 6031 5756
rect 6015 5676 6031 5690
rect 6035 5678 6037 5756
rect 6049 5678 6051 5756
rect 6035 5676 6051 5678
rect 6055 5744 6071 5756
rect 6055 5676 6057 5744
rect 6069 5676 6071 5744
rect 6075 5676 6077 5756
rect 6129 5716 6131 5756
rect 6135 5716 6137 5756
rect 6149 5716 6151 5756
rect 6155 5720 6157 5756
rect 6169 5720 6171 5756
rect 6155 5716 6171 5720
rect 6175 5716 6177 5756
rect 6243 5716 6245 5756
rect 6249 5716 6251 5756
rect 6289 5684 6291 5756
rect 6277 5676 6291 5684
rect 6295 5688 6297 5756
rect 6309 5688 6311 5756
rect 6295 5676 6311 5688
rect 6315 5676 6317 5756
rect 6329 5676 6331 5756
rect 6335 5676 6337 5756
rect 6389 5716 6391 5756
rect 6395 5716 6397 5756
rect 6409 5716 6411 5756
rect 6415 5720 6417 5756
rect 6429 5720 6431 5756
rect 6415 5716 6431 5720
rect 6435 5716 6437 5756
rect 6489 5716 6491 5756
rect 6495 5716 6497 5756
rect 6509 5716 6511 5756
rect 6515 5720 6517 5756
rect 6529 5720 6531 5756
rect 6515 5716 6531 5720
rect 6535 5716 6537 5756
rect 6589 5716 6591 5756
rect 6595 5716 6597 5756
rect 6609 5716 6611 5756
rect 6615 5720 6617 5756
rect 6629 5720 6631 5756
rect 6615 5716 6631 5720
rect 6635 5716 6637 5756
rect 29 5304 31 5384
rect 35 5324 44 5384
rect 212 5344 221 5384
rect 70 5324 81 5344
rect 35 5304 37 5324
rect 49 5304 53 5324
rect 57 5304 61 5324
rect 65 5304 67 5324
rect 79 5304 81 5324
rect 85 5304 89 5344
rect 93 5304 95 5344
rect 133 5304 135 5344
rect 139 5304 141 5344
rect 153 5304 155 5344
rect 159 5304 167 5344
rect 171 5304 173 5344
rect 185 5304 187 5344
rect 191 5304 201 5344
rect 205 5304 207 5344
rect 219 5304 221 5344
rect 225 5304 227 5384
rect 269 5304 271 5344
rect 275 5304 277 5344
rect 289 5304 291 5344
rect 295 5304 297 5344
rect 363 5304 365 5384
rect 369 5304 371 5384
rect 383 5304 385 5384
rect 389 5372 405 5384
rect 389 5304 391 5372
rect 403 5304 405 5372
rect 409 5376 423 5384
rect 409 5304 411 5376
rect 463 5304 465 5344
rect 469 5304 471 5344
rect 483 5304 485 5344
rect 489 5304 491 5344
rect 539 5304 541 5384
rect 545 5304 547 5384
rect 559 5304 563 5344
rect 567 5304 571 5344
rect 583 5304 585 5344
rect 589 5304 591 5344
rect 629 5304 631 5384
rect 635 5304 639 5384
rect 643 5304 645 5384
rect 709 5304 711 5384
rect 715 5304 719 5384
rect 723 5304 725 5384
rect 997 5376 1011 5384
rect 789 5304 791 5344
rect 795 5304 797 5344
rect 809 5304 811 5344
rect 815 5304 817 5344
rect 869 5304 871 5344
rect 875 5304 877 5344
rect 889 5304 891 5344
rect 895 5304 897 5344
rect 949 5304 951 5344
rect 955 5304 957 5344
rect 1009 5304 1011 5376
rect 1015 5372 1031 5384
rect 1015 5304 1017 5372
rect 1029 5304 1031 5372
rect 1035 5304 1037 5384
rect 1049 5304 1051 5384
rect 1055 5304 1057 5384
rect 1123 5304 1125 5384
rect 1129 5316 1131 5384
rect 1143 5316 1145 5384
rect 1129 5304 1145 5316
rect 1149 5382 1165 5384
rect 1149 5304 1151 5382
rect 1163 5304 1165 5382
rect 1169 5370 1185 5384
rect 1169 5304 1171 5370
rect 1183 5304 1185 5370
rect 1189 5382 1203 5384
rect 1189 5304 1191 5382
rect 1229 5304 1231 5384
rect 1235 5324 1244 5384
rect 1412 5344 1421 5384
rect 1270 5324 1281 5344
rect 1235 5304 1237 5324
rect 1249 5304 1253 5324
rect 1257 5304 1261 5324
rect 1265 5304 1267 5324
rect 1279 5304 1281 5324
rect 1285 5304 1289 5344
rect 1293 5304 1295 5344
rect 1333 5304 1335 5344
rect 1339 5304 1341 5344
rect 1353 5304 1355 5344
rect 1359 5304 1367 5344
rect 1371 5304 1373 5344
rect 1385 5304 1387 5344
rect 1391 5304 1401 5344
rect 1405 5304 1407 5344
rect 1419 5304 1421 5344
rect 1425 5304 1427 5384
rect 1483 5304 1485 5344
rect 1489 5340 1505 5344
rect 1489 5304 1491 5340
rect 1503 5304 1505 5340
rect 1509 5304 1511 5344
rect 1523 5304 1525 5344
rect 1529 5304 1531 5344
rect 1583 5304 1585 5344
rect 1589 5340 1605 5344
rect 1589 5304 1591 5340
rect 1603 5304 1605 5340
rect 1609 5304 1611 5344
rect 1623 5304 1625 5344
rect 1629 5304 1631 5344
rect 1683 5304 1685 5344
rect 1689 5304 1691 5344
rect 1748 5304 1750 5344
rect 1754 5304 1758 5344
rect 1770 5304 1772 5384
rect 1776 5304 1780 5384
rect 1784 5304 1786 5384
rect 1839 5304 1841 5384
rect 1845 5304 1847 5384
rect 1859 5304 1863 5344
rect 1867 5304 1871 5344
rect 1883 5304 1885 5344
rect 1889 5304 1891 5344
rect 1943 5304 1945 5344
rect 1949 5304 1951 5344
rect 1963 5304 1965 5344
rect 1969 5304 1971 5344
rect 2028 5304 2030 5344
rect 2034 5304 2038 5344
rect 2050 5304 2052 5384
rect 2056 5304 2060 5384
rect 2064 5304 2066 5384
rect 2109 5304 2111 5344
rect 2115 5304 2117 5344
rect 2129 5304 2131 5344
rect 2135 5304 2137 5344
rect 2203 5304 2205 5344
rect 2209 5304 2211 5344
rect 2268 5304 2270 5344
rect 2274 5304 2278 5344
rect 2290 5304 2292 5384
rect 2296 5304 2300 5384
rect 2304 5304 2306 5384
rect 2349 5304 2351 5384
rect 2355 5304 2359 5384
rect 2363 5304 2365 5384
rect 2443 5304 2445 5344
rect 2449 5304 2451 5344
rect 2503 5304 2505 5384
rect 2509 5304 2511 5384
rect 2523 5304 2525 5384
rect 2529 5372 2545 5384
rect 2529 5304 2531 5372
rect 2543 5304 2545 5372
rect 2549 5376 2563 5384
rect 2549 5304 2551 5376
rect 2594 5304 2596 5384
rect 2600 5304 2604 5384
rect 2608 5304 2610 5384
rect 2622 5304 2626 5344
rect 2630 5304 2632 5344
rect 2689 5304 2691 5344
rect 2695 5304 2697 5344
rect 2709 5304 2711 5344
rect 2715 5304 2717 5344
rect 2783 5304 2785 5344
rect 2789 5340 2805 5344
rect 2789 5304 2791 5340
rect 2803 5304 2805 5340
rect 2809 5304 2811 5344
rect 2823 5304 2825 5344
rect 2829 5304 2831 5344
rect 2883 5304 2885 5344
rect 2889 5304 2891 5344
rect 2903 5304 2905 5344
rect 2909 5304 2911 5344
rect 2975 5304 2977 5384
rect 2981 5304 2985 5384
rect 2989 5304 2991 5384
rect 3034 5304 3036 5384
rect 3040 5304 3044 5384
rect 3048 5304 3050 5384
rect 3062 5304 3066 5344
rect 3070 5304 3072 5344
rect 3143 5304 3145 5344
rect 3149 5304 3151 5344
rect 3163 5304 3165 5344
rect 3169 5304 3171 5344
rect 3214 5304 3216 5384
rect 3220 5304 3224 5384
rect 3228 5304 3230 5384
rect 3242 5304 3246 5344
rect 3250 5304 3252 5344
rect 3319 5304 3321 5384
rect 3325 5304 3327 5384
rect 3339 5304 3343 5344
rect 3347 5304 3351 5344
rect 3363 5304 3365 5344
rect 3369 5304 3371 5344
rect 3409 5304 3411 5384
rect 3415 5304 3419 5384
rect 3423 5304 3425 5384
rect 3489 5304 3491 5384
rect 3495 5304 3501 5384
rect 3505 5383 3521 5384
rect 3505 5304 3507 5383
rect 3519 5304 3521 5383
rect 3525 5383 3539 5384
rect 3525 5304 3527 5383
rect 3594 5304 3596 5384
rect 3600 5304 3604 5384
rect 3608 5304 3610 5384
rect 3622 5304 3626 5344
rect 3630 5304 3632 5344
rect 3715 5304 3717 5384
rect 3721 5304 3725 5384
rect 3729 5304 3731 5384
rect 3769 5304 3771 5384
rect 3775 5304 3781 5384
rect 3785 5304 3787 5384
rect 3809 5304 3811 5384
rect 3815 5304 3821 5384
rect 3825 5304 3827 5384
rect 3915 5304 3917 5384
rect 3921 5304 3925 5384
rect 3929 5304 3931 5384
rect 3974 5304 3976 5384
rect 3980 5304 3984 5384
rect 3988 5304 3990 5384
rect 4002 5304 4006 5344
rect 4010 5304 4012 5344
rect 4083 5304 4085 5344
rect 4089 5340 4105 5344
rect 4089 5304 4091 5340
rect 4103 5304 4105 5340
rect 4109 5304 4111 5344
rect 4123 5304 4125 5344
rect 4129 5304 4131 5344
rect 4183 5304 4185 5344
rect 4189 5304 4191 5344
rect 4203 5304 4205 5344
rect 4209 5304 4211 5344
rect 4249 5304 4251 5344
rect 4255 5304 4257 5344
rect 4328 5304 4330 5344
rect 4334 5304 4338 5344
rect 4350 5304 4352 5384
rect 4356 5304 4360 5384
rect 4364 5304 4366 5384
rect 4423 5304 4425 5344
rect 4429 5304 4431 5344
rect 4443 5304 4445 5344
rect 4449 5304 4451 5344
rect 4489 5304 4491 5344
rect 4495 5304 4497 5344
rect 4509 5304 4511 5344
rect 4515 5304 4517 5344
rect 4588 5304 4590 5344
rect 4594 5304 4598 5344
rect 4610 5304 4612 5384
rect 4616 5304 4620 5384
rect 4624 5304 4626 5384
rect 4688 5304 4690 5344
rect 4694 5304 4698 5344
rect 4710 5304 4712 5384
rect 4716 5304 4720 5384
rect 4724 5304 4726 5384
rect 4779 5304 4781 5384
rect 4785 5304 4787 5384
rect 4799 5304 4803 5344
rect 4807 5304 4811 5344
rect 4823 5304 4825 5344
rect 4829 5304 4831 5344
rect 4888 5304 4890 5344
rect 4894 5304 4898 5344
rect 4910 5304 4912 5384
rect 4916 5304 4920 5384
rect 4924 5304 4926 5384
rect 4983 5304 4985 5344
rect 4989 5304 4991 5344
rect 5003 5304 5005 5344
rect 5009 5304 5011 5344
rect 5059 5304 5061 5384
rect 5065 5304 5067 5384
rect 5079 5304 5083 5344
rect 5087 5304 5091 5344
rect 5103 5304 5105 5344
rect 5109 5304 5111 5344
rect 5149 5304 5151 5344
rect 5155 5304 5157 5344
rect 5169 5304 5171 5344
rect 5175 5304 5177 5344
rect 5234 5304 5236 5384
rect 5240 5304 5244 5384
rect 5248 5304 5250 5384
rect 5262 5304 5266 5344
rect 5270 5304 5272 5344
rect 5339 5304 5341 5384
rect 5345 5304 5347 5384
rect 5359 5304 5363 5344
rect 5367 5304 5371 5344
rect 5383 5304 5385 5344
rect 5389 5304 5391 5344
rect 5434 5304 5436 5384
rect 5440 5304 5444 5384
rect 5448 5304 5450 5384
rect 5462 5304 5466 5344
rect 5470 5304 5472 5344
rect 5529 5304 5531 5344
rect 5535 5304 5537 5344
rect 5549 5304 5551 5344
rect 5555 5304 5557 5344
rect 5609 5304 5611 5344
rect 5615 5304 5617 5344
rect 5629 5304 5631 5344
rect 5635 5340 5651 5344
rect 5635 5304 5637 5340
rect 5649 5304 5651 5340
rect 5655 5304 5657 5344
rect 5719 5304 5721 5384
rect 5725 5304 5727 5384
rect 5739 5304 5743 5344
rect 5747 5304 5751 5344
rect 5763 5304 5765 5344
rect 5769 5304 5771 5344
rect 5823 5304 5825 5384
rect 5829 5316 5831 5384
rect 5843 5316 5845 5384
rect 5829 5304 5845 5316
rect 5849 5382 5865 5384
rect 5849 5304 5851 5382
rect 5863 5304 5865 5382
rect 5869 5370 5885 5384
rect 5869 5304 5871 5370
rect 5883 5304 5885 5370
rect 5889 5382 5903 5384
rect 5889 5304 5891 5382
rect 6097 5376 6111 5384
rect 5929 5304 5931 5344
rect 5935 5304 5937 5344
rect 5949 5304 5951 5344
rect 5955 5304 5957 5344
rect 6009 5304 6011 5344
rect 6015 5304 6017 5344
rect 6029 5304 6031 5344
rect 6035 5340 6051 5344
rect 6035 5304 6037 5340
rect 6049 5304 6051 5340
rect 6055 5304 6057 5344
rect 6109 5304 6111 5376
rect 6115 5372 6131 5384
rect 6115 5304 6117 5372
rect 6129 5304 6131 5372
rect 6135 5304 6137 5384
rect 6149 5304 6151 5384
rect 6155 5304 6157 5384
rect 6228 5304 6230 5344
rect 6234 5304 6238 5344
rect 6250 5304 6252 5384
rect 6256 5304 6260 5384
rect 6264 5304 6266 5384
rect 6314 5304 6316 5384
rect 6320 5304 6324 5384
rect 6328 5304 6330 5384
rect 6342 5304 6346 5344
rect 6350 5304 6352 5344
rect 6428 5304 6430 5344
rect 6434 5304 6438 5344
rect 6450 5304 6452 5384
rect 6456 5304 6460 5384
rect 6464 5304 6466 5384
rect 6523 5304 6525 5344
rect 6529 5340 6545 5344
rect 6529 5304 6531 5340
rect 6543 5304 6545 5340
rect 6549 5304 6551 5344
rect 6563 5304 6565 5344
rect 6569 5304 6571 5344
rect 6623 5304 6625 5384
rect 6629 5304 6631 5384
rect 6643 5304 6645 5384
rect 6649 5372 6665 5384
rect 6649 5304 6651 5372
rect 6663 5304 6665 5372
rect 6669 5376 6683 5384
rect 6669 5304 6671 5376
rect 41 5196 43 5276
rect 47 5196 49 5276
rect 61 5236 65 5276
rect 69 5236 71 5276
rect 109 5196 111 5276
rect 115 5256 117 5276
rect 129 5256 133 5276
rect 137 5256 141 5276
rect 145 5256 147 5276
rect 159 5256 161 5276
rect 115 5196 124 5256
rect 150 5236 161 5256
rect 165 5236 169 5276
rect 173 5236 175 5276
rect 213 5236 215 5276
rect 219 5236 221 5276
rect 233 5236 235 5276
rect 239 5236 247 5276
rect 251 5236 253 5276
rect 265 5236 267 5276
rect 271 5236 281 5276
rect 285 5236 287 5276
rect 299 5236 301 5276
rect 292 5196 301 5236
rect 305 5196 307 5276
rect 349 5236 351 5276
rect 355 5236 357 5276
rect 369 5236 371 5276
rect 375 5236 377 5276
rect 443 5196 445 5276
rect 449 5196 451 5276
rect 463 5196 465 5276
rect 469 5208 471 5276
rect 483 5208 485 5276
rect 469 5196 485 5208
rect 489 5204 491 5276
rect 543 5236 545 5276
rect 549 5236 551 5276
rect 563 5236 565 5276
rect 569 5236 571 5276
rect 489 5196 503 5204
rect 613 5196 615 5276
rect 619 5236 621 5276
rect 633 5236 635 5276
rect 639 5236 649 5276
rect 653 5236 655 5276
rect 667 5236 669 5276
rect 673 5236 681 5276
rect 685 5236 687 5276
rect 699 5236 701 5276
rect 705 5236 707 5276
rect 745 5236 747 5276
rect 751 5236 755 5276
rect 759 5256 761 5276
rect 773 5256 775 5276
rect 779 5256 783 5276
rect 787 5256 791 5276
rect 803 5256 805 5276
rect 759 5236 770 5256
rect 619 5196 628 5236
rect 796 5196 805 5256
rect 809 5196 811 5276
rect 849 5236 851 5276
rect 855 5236 857 5276
rect 869 5236 871 5276
rect 875 5236 877 5276
rect 948 5236 950 5276
rect 954 5236 958 5276
rect 970 5196 972 5276
rect 976 5196 980 5276
rect 984 5196 986 5276
rect 1048 5236 1050 5276
rect 1054 5236 1058 5276
rect 1070 5196 1072 5276
rect 1076 5196 1080 5276
rect 1084 5196 1086 5276
rect 1139 5196 1141 5276
rect 1145 5196 1147 5276
rect 1159 5236 1163 5276
rect 1167 5236 1171 5276
rect 1183 5236 1185 5276
rect 1189 5236 1191 5276
rect 1229 5196 1231 5276
rect 1235 5256 1237 5276
rect 1249 5256 1253 5276
rect 1257 5256 1261 5276
rect 1265 5256 1267 5276
rect 1279 5256 1281 5276
rect 1235 5196 1244 5256
rect 1270 5236 1281 5256
rect 1285 5236 1289 5276
rect 1293 5236 1295 5276
rect 1333 5236 1335 5276
rect 1339 5236 1341 5276
rect 1353 5236 1355 5276
rect 1359 5236 1367 5276
rect 1371 5236 1373 5276
rect 1385 5236 1387 5276
rect 1391 5236 1401 5276
rect 1405 5236 1407 5276
rect 1419 5236 1421 5276
rect 1412 5196 1421 5236
rect 1425 5196 1427 5276
rect 1483 5236 1485 5276
rect 1489 5236 1491 5276
rect 1503 5236 1505 5276
rect 1509 5236 1511 5276
rect 1549 5236 1551 5276
rect 1555 5236 1557 5276
rect 1569 5236 1571 5276
rect 1575 5236 1577 5276
rect 1629 5196 1631 5276
rect 1635 5256 1637 5276
rect 1649 5256 1653 5276
rect 1657 5256 1661 5276
rect 1665 5256 1667 5276
rect 1679 5256 1681 5276
rect 1635 5196 1644 5256
rect 1670 5236 1681 5256
rect 1685 5236 1689 5276
rect 1693 5236 1695 5276
rect 1733 5236 1735 5276
rect 1739 5236 1741 5276
rect 1753 5236 1755 5276
rect 1759 5236 1767 5276
rect 1771 5236 1773 5276
rect 1785 5236 1787 5276
rect 1791 5236 1801 5276
rect 1805 5236 1807 5276
rect 1819 5236 1821 5276
rect 1812 5196 1821 5236
rect 1825 5196 1827 5276
rect 1883 5196 1885 5276
rect 1889 5264 1905 5276
rect 1889 5196 1891 5264
rect 1903 5196 1905 5264
rect 1909 5198 1911 5276
rect 1923 5198 1925 5276
rect 1909 5196 1925 5198
rect 1929 5210 1931 5276
rect 1943 5210 1945 5276
rect 1929 5196 1945 5210
rect 1949 5198 1951 5276
rect 1989 5236 1991 5276
rect 1995 5236 1997 5276
rect 1949 5196 1963 5198
rect 2059 5196 2061 5276
rect 2065 5196 2067 5276
rect 2079 5236 2083 5276
rect 2087 5236 2091 5276
rect 2103 5236 2105 5276
rect 2109 5236 2111 5276
rect 2149 5236 2151 5276
rect 2155 5236 2157 5276
rect 2169 5236 2171 5276
rect 2175 5236 2177 5276
rect 2253 5197 2255 5276
rect 2241 5196 2255 5197
rect 2259 5197 2261 5276
rect 2273 5197 2275 5276
rect 2259 5196 2275 5197
rect 2279 5196 2285 5276
rect 2289 5196 2291 5276
rect 2343 5236 2345 5276
rect 2349 5236 2351 5276
rect 2363 5236 2365 5276
rect 2369 5236 2371 5276
rect 2423 5236 2425 5276
rect 2429 5240 2431 5276
rect 2443 5240 2445 5276
rect 2429 5236 2445 5240
rect 2449 5236 2451 5276
rect 2463 5236 2465 5276
rect 2469 5236 2471 5276
rect 2535 5196 2537 5276
rect 2541 5196 2545 5276
rect 2549 5196 2551 5276
rect 2589 5236 2591 5276
rect 2595 5236 2597 5276
rect 2659 5196 2661 5276
rect 2665 5196 2667 5276
rect 2679 5236 2683 5276
rect 2687 5236 2691 5276
rect 2703 5236 2705 5276
rect 2709 5236 2711 5276
rect 2749 5196 2751 5276
rect 2755 5196 2759 5276
rect 2763 5196 2765 5276
rect 2843 5236 2845 5276
rect 2849 5236 2851 5276
rect 2863 5236 2865 5276
rect 2869 5236 2871 5276
rect 2923 5236 2925 5276
rect 2929 5236 2931 5276
rect 2943 5236 2945 5276
rect 2949 5236 2951 5276
rect 2989 5196 2991 5276
rect 2995 5196 3001 5276
rect 3005 5197 3007 5276
rect 3019 5197 3021 5276
rect 3005 5196 3021 5197
rect 3025 5197 3027 5276
rect 3025 5196 3039 5197
rect 3099 5196 3101 5276
rect 3105 5196 3107 5276
rect 3119 5236 3123 5276
rect 3127 5236 3131 5276
rect 3143 5236 3145 5276
rect 3149 5236 3151 5276
rect 3189 5236 3191 5276
rect 3195 5236 3197 5276
rect 3209 5236 3211 5276
rect 3215 5236 3217 5276
rect 3283 5236 3285 5276
rect 3289 5240 3291 5276
rect 3303 5240 3305 5276
rect 3289 5236 3305 5240
rect 3309 5236 3311 5276
rect 3323 5236 3325 5276
rect 3329 5236 3331 5276
rect 3383 5236 3385 5276
rect 3389 5236 3391 5276
rect 3443 5196 3445 5276
rect 3449 5196 3451 5276
rect 3463 5196 3465 5276
rect 3469 5208 3471 5276
rect 3483 5208 3485 5276
rect 3469 5196 3485 5208
rect 3489 5204 3491 5276
rect 3489 5196 3503 5204
rect 3555 5196 3557 5276
rect 3561 5196 3565 5276
rect 3569 5196 3571 5276
rect 3614 5196 3616 5276
rect 3620 5196 3624 5276
rect 3628 5196 3630 5276
rect 3642 5236 3646 5276
rect 3650 5236 3652 5276
rect 3728 5236 3730 5276
rect 3734 5236 3738 5276
rect 3750 5196 3752 5276
rect 3756 5196 3760 5276
rect 3764 5196 3766 5276
rect 3809 5196 3811 5276
rect 3815 5196 3819 5276
rect 3823 5196 3825 5276
rect 3889 5236 3891 5276
rect 3895 5236 3897 5276
rect 3909 5236 3911 5276
rect 3915 5236 3917 5276
rect 3983 5236 3985 5276
rect 3989 5236 3991 5276
rect 4003 5236 4005 5276
rect 4009 5236 4011 5276
rect 4054 5196 4056 5276
rect 4060 5196 4064 5276
rect 4068 5196 4070 5276
rect 4082 5236 4086 5276
rect 4090 5236 4092 5276
rect 4163 5236 4165 5276
rect 4169 5236 4171 5276
rect 4183 5236 4185 5276
rect 4189 5236 4191 5276
rect 4239 5196 4241 5276
rect 4245 5196 4247 5276
rect 4259 5236 4263 5276
rect 4267 5236 4271 5276
rect 4283 5236 4285 5276
rect 4289 5236 4291 5276
rect 4343 5236 4345 5276
rect 4349 5236 4351 5276
rect 4363 5236 4365 5276
rect 4369 5236 4371 5276
rect 4428 5236 4430 5276
rect 4434 5236 4438 5276
rect 4450 5196 4452 5276
rect 4456 5196 4460 5276
rect 4464 5196 4466 5276
rect 4528 5236 4530 5276
rect 4534 5236 4538 5276
rect 4550 5196 4552 5276
rect 4556 5196 4560 5276
rect 4564 5196 4566 5276
rect 4609 5236 4611 5276
rect 4615 5236 4617 5276
rect 4629 5236 4631 5276
rect 4635 5236 4637 5276
rect 4689 5236 4691 5276
rect 4695 5236 4697 5276
rect 4709 5236 4711 5276
rect 4715 5236 4717 5276
rect 4769 5236 4771 5276
rect 4775 5236 4777 5276
rect 4843 5236 4845 5276
rect 4849 5240 4851 5276
rect 4863 5240 4865 5276
rect 4849 5236 4865 5240
rect 4869 5236 4871 5276
rect 4883 5236 4885 5276
rect 4889 5236 4891 5276
rect 4934 5196 4936 5276
rect 4940 5196 4944 5276
rect 4948 5196 4950 5276
rect 4962 5236 4966 5276
rect 4970 5236 4972 5276
rect 5029 5196 5031 5276
rect 5035 5196 5037 5276
rect 5089 5236 5091 5276
rect 5095 5236 5097 5276
rect 5109 5236 5111 5276
rect 5115 5236 5117 5276
rect 5157 5274 5171 5276
rect 5169 5196 5171 5274
rect 5175 5196 5177 5276
rect 5189 5196 5191 5276
rect 5195 5196 5197 5276
rect 5249 5236 5251 5276
rect 5255 5236 5257 5276
rect 5269 5236 5271 5276
rect 5275 5236 5277 5276
rect 5334 5196 5336 5276
rect 5340 5196 5344 5276
rect 5348 5196 5350 5276
rect 5362 5236 5366 5276
rect 5370 5236 5372 5276
rect 5429 5236 5431 5276
rect 5435 5236 5437 5276
rect 5449 5236 5451 5276
rect 5455 5240 5457 5276
rect 5469 5240 5471 5276
rect 5455 5236 5471 5240
rect 5475 5236 5477 5276
rect 5529 5236 5531 5276
rect 5535 5236 5537 5276
rect 5549 5236 5551 5276
rect 5555 5240 5557 5276
rect 5569 5240 5571 5276
rect 5555 5236 5571 5240
rect 5575 5236 5577 5276
rect 5629 5236 5631 5276
rect 5635 5236 5637 5276
rect 5689 5236 5691 5276
rect 5695 5236 5697 5276
rect 5709 5236 5711 5276
rect 5715 5240 5717 5276
rect 5729 5240 5731 5276
rect 5715 5236 5731 5240
rect 5735 5236 5737 5276
rect 5794 5196 5796 5276
rect 5800 5196 5804 5276
rect 5808 5196 5810 5276
rect 5822 5236 5826 5276
rect 5830 5236 5832 5276
rect 5903 5236 5905 5276
rect 5909 5236 5911 5276
rect 5923 5236 5925 5276
rect 5929 5236 5931 5276
rect 5969 5236 5971 5276
rect 5975 5236 5977 5276
rect 5989 5236 5991 5276
rect 5995 5240 5997 5276
rect 6009 5240 6011 5276
rect 5995 5236 6011 5240
rect 6015 5236 6017 5276
rect 6069 5236 6071 5276
rect 6075 5236 6077 5276
rect 6089 5236 6091 5276
rect 6095 5236 6097 5276
rect 6163 5196 6165 5276
rect 6169 5196 6171 5276
rect 6183 5196 6185 5276
rect 6189 5208 6191 5276
rect 6203 5208 6205 5276
rect 6189 5196 6205 5208
rect 6209 5204 6211 5276
rect 6263 5236 6265 5276
rect 6269 5236 6271 5276
rect 6323 5236 6325 5276
rect 6329 5240 6331 5276
rect 6343 5240 6345 5276
rect 6329 5236 6345 5240
rect 6349 5236 6351 5276
rect 6363 5236 6365 5276
rect 6369 5236 6371 5276
rect 6423 5236 6425 5276
rect 6429 5240 6431 5276
rect 6443 5240 6445 5276
rect 6429 5236 6445 5240
rect 6449 5236 6451 5276
rect 6463 5236 6465 5276
rect 6469 5236 6471 5276
rect 6509 5236 6511 5276
rect 6515 5236 6517 5276
rect 6583 5236 6585 5276
rect 6589 5240 6591 5276
rect 6603 5240 6605 5276
rect 6589 5236 6605 5240
rect 6609 5236 6611 5276
rect 6623 5236 6625 5276
rect 6629 5236 6631 5276
rect 6669 5236 6671 5276
rect 6675 5236 6677 5276
rect 6689 5236 6691 5276
rect 6695 5236 6697 5276
rect 6209 5196 6223 5204
rect 41 4824 43 4904
rect 47 4824 49 4904
rect 61 4824 65 4864
rect 69 4824 71 4864
rect 121 4824 123 4904
rect 127 4824 129 4904
rect 141 4824 145 4864
rect 149 4824 151 4864
rect 203 4824 205 4864
rect 209 4824 211 4864
rect 223 4824 225 4864
rect 229 4824 231 4864
rect 269 4824 271 4904
rect 275 4844 284 4904
rect 452 4864 461 4904
rect 310 4844 321 4864
rect 275 4824 277 4844
rect 289 4824 293 4844
rect 297 4824 301 4844
rect 305 4824 307 4844
rect 319 4824 321 4844
rect 325 4824 329 4864
rect 333 4824 335 4864
rect 373 4824 375 4864
rect 379 4824 381 4864
rect 393 4824 395 4864
rect 399 4824 407 4864
rect 411 4824 413 4864
rect 425 4824 427 4864
rect 431 4824 441 4864
rect 445 4824 447 4864
rect 459 4824 461 4864
rect 465 4824 467 4904
rect 523 4824 525 4904
rect 529 4824 531 4904
rect 543 4824 545 4904
rect 549 4892 565 4904
rect 549 4824 551 4892
rect 563 4824 565 4892
rect 569 4896 583 4904
rect 569 4824 571 4896
rect 623 4824 625 4864
rect 629 4824 631 4864
rect 643 4824 645 4864
rect 649 4824 651 4864
rect 689 4824 691 4864
rect 695 4824 697 4864
rect 709 4824 711 4864
rect 715 4824 717 4864
rect 783 4824 785 4864
rect 789 4824 791 4864
rect 803 4824 805 4864
rect 809 4824 811 4864
rect 849 4824 851 4904
rect 855 4844 864 4904
rect 1032 4864 1041 4904
rect 890 4844 901 4864
rect 855 4824 857 4844
rect 869 4824 873 4844
rect 877 4824 881 4844
rect 885 4824 887 4844
rect 899 4824 901 4844
rect 905 4824 909 4864
rect 913 4824 915 4864
rect 953 4824 955 4864
rect 959 4824 961 4864
rect 973 4824 975 4864
rect 979 4824 987 4864
rect 991 4824 993 4864
rect 1005 4824 1007 4864
rect 1011 4824 1021 4864
rect 1025 4824 1027 4864
rect 1039 4824 1041 4864
rect 1045 4824 1047 4904
rect 1101 4824 1103 4904
rect 1107 4824 1109 4904
rect 1121 4824 1125 4864
rect 1129 4824 1131 4864
rect 1183 4824 1185 4904
rect 1189 4824 1191 4904
rect 1203 4824 1205 4904
rect 1209 4892 1225 4904
rect 1209 4824 1211 4892
rect 1223 4824 1225 4892
rect 1229 4896 1243 4904
rect 1229 4824 1231 4896
rect 1283 4824 1285 4864
rect 1289 4824 1291 4864
rect 1303 4824 1305 4864
rect 1309 4824 1311 4864
rect 1361 4824 1363 4904
rect 1367 4824 1369 4904
rect 1381 4824 1385 4864
rect 1389 4824 1391 4864
rect 1429 4824 1431 4864
rect 1435 4824 1437 4864
rect 1449 4824 1451 4864
rect 1455 4824 1457 4864
rect 1523 4824 1525 4864
rect 1529 4824 1531 4864
rect 1543 4824 1545 4864
rect 1549 4824 1551 4864
rect 1608 4824 1610 4864
rect 1614 4824 1618 4864
rect 1630 4824 1632 4904
rect 1636 4824 1640 4904
rect 1644 4824 1646 4904
rect 1703 4824 1705 4864
rect 1709 4824 1711 4864
rect 1723 4824 1725 4864
rect 1729 4824 1731 4864
rect 1788 4824 1790 4864
rect 1794 4824 1798 4864
rect 1810 4824 1812 4904
rect 1816 4824 1820 4904
rect 1824 4824 1826 4904
rect 1869 4824 1871 4864
rect 1875 4824 1877 4864
rect 1889 4824 1891 4864
rect 1895 4824 1897 4864
rect 1968 4824 1970 4864
rect 1974 4824 1978 4864
rect 1990 4824 1992 4904
rect 1996 4824 2000 4904
rect 2004 4824 2006 4904
rect 2068 4824 2070 4864
rect 2074 4824 2078 4864
rect 2090 4824 2092 4904
rect 2096 4824 2100 4904
rect 2104 4824 2106 4904
rect 2159 4824 2161 4904
rect 2165 4824 2167 4904
rect 2179 4824 2183 4864
rect 2187 4824 2191 4864
rect 2203 4824 2205 4864
rect 2209 4824 2211 4864
rect 2249 4824 2251 4864
rect 2255 4824 2257 4864
rect 2335 4824 2337 4904
rect 2341 4824 2345 4904
rect 2349 4824 2351 4904
rect 2401 4903 2415 4904
rect 2413 4824 2415 4903
rect 2419 4903 2435 4904
rect 2419 4824 2421 4903
rect 2433 4824 2435 4903
rect 2439 4824 2445 4904
rect 2449 4824 2451 4904
rect 2503 4824 2505 4864
rect 2509 4824 2511 4864
rect 2523 4824 2525 4864
rect 2529 4824 2531 4864
rect 2588 4824 2590 4864
rect 2594 4824 2598 4864
rect 2610 4824 2612 4904
rect 2616 4824 2620 4904
rect 2624 4824 2626 4904
rect 2688 4824 2690 4864
rect 2694 4824 2698 4864
rect 2710 4824 2712 4904
rect 2716 4824 2720 4904
rect 2724 4824 2726 4904
rect 2783 4824 2785 4864
rect 2789 4824 2791 4864
rect 2834 4824 2836 4904
rect 2840 4824 2844 4904
rect 2848 4824 2850 4904
rect 2862 4824 2866 4864
rect 2870 4824 2872 4864
rect 2948 4824 2950 4864
rect 2954 4824 2958 4864
rect 2970 4824 2972 4904
rect 2976 4824 2980 4904
rect 2984 4824 2986 4904
rect 3048 4824 3050 4864
rect 3054 4824 3058 4864
rect 3070 4824 3072 4904
rect 3076 4824 3080 4904
rect 3084 4824 3086 4904
rect 3155 4824 3157 4904
rect 3161 4824 3165 4904
rect 3169 4824 3171 4904
rect 3223 4824 3225 4904
rect 3229 4824 3231 4904
rect 3283 4824 3285 4864
rect 3289 4824 3291 4864
rect 3303 4824 3305 4864
rect 3309 4824 3311 4864
rect 3368 4824 3370 4864
rect 3374 4824 3378 4864
rect 3390 4824 3392 4904
rect 3396 4824 3400 4904
rect 3404 4824 3406 4904
rect 3453 4824 3455 4904
rect 3459 4864 3468 4904
rect 3459 4824 3461 4864
rect 3473 4824 3475 4864
rect 3479 4824 3489 4864
rect 3493 4824 3495 4864
rect 3507 4824 3509 4864
rect 3513 4824 3521 4864
rect 3525 4824 3527 4864
rect 3539 4824 3541 4864
rect 3545 4824 3547 4864
rect 3585 4824 3587 4864
rect 3591 4824 3595 4864
rect 3599 4844 3610 4864
rect 3636 4844 3645 4904
rect 3599 4824 3601 4844
rect 3613 4824 3615 4844
rect 3619 4824 3623 4844
rect 3627 4824 3631 4844
rect 3643 4824 3645 4844
rect 3649 4824 3651 4904
rect 3694 4824 3696 4904
rect 3700 4824 3704 4904
rect 3708 4824 3710 4904
rect 3722 4824 3726 4864
rect 3730 4824 3732 4864
rect 3803 4824 3805 4904
rect 3809 4824 3811 4904
rect 3823 4824 3825 4904
rect 3829 4892 3845 4904
rect 3829 4824 3831 4892
rect 3843 4824 3845 4892
rect 3849 4896 3863 4904
rect 3849 4824 3851 4896
rect 3903 4824 3905 4864
rect 3909 4860 3925 4864
rect 3909 4824 3911 4860
rect 3923 4824 3925 4860
rect 3929 4824 3931 4864
rect 3943 4824 3945 4864
rect 3949 4824 3951 4864
rect 4003 4824 4005 4904
rect 4009 4824 4011 4904
rect 4023 4824 4025 4904
rect 4029 4892 4045 4904
rect 4029 4824 4031 4892
rect 4043 4824 4045 4892
rect 4049 4896 4063 4904
rect 4049 4824 4051 4896
rect 4103 4824 4105 4904
rect 4109 4824 4111 4904
rect 4159 4824 4161 4904
rect 4165 4824 4167 4904
rect 4179 4824 4183 4864
rect 4187 4824 4191 4864
rect 4203 4824 4205 4864
rect 4209 4824 4211 4864
rect 4263 4824 4265 4864
rect 4269 4824 4271 4864
rect 4283 4824 4285 4864
rect 4289 4824 4291 4864
rect 4329 4824 4331 4864
rect 4335 4824 4337 4864
rect 4349 4824 4353 4864
rect 4357 4824 4361 4864
rect 4373 4824 4375 4904
rect 4379 4824 4381 4904
rect 4448 4824 4450 4864
rect 4454 4824 4458 4864
rect 4470 4824 4472 4904
rect 4476 4824 4480 4904
rect 4484 4824 4486 4904
rect 4529 4824 4531 4864
rect 4535 4824 4537 4864
rect 4549 4824 4551 4864
rect 4555 4860 4571 4864
rect 4555 4824 4557 4860
rect 4569 4824 4571 4860
rect 4575 4824 4577 4864
rect 4634 4824 4636 4904
rect 4640 4824 4644 4904
rect 4648 4824 4650 4904
rect 4662 4824 4666 4864
rect 4670 4824 4672 4864
rect 4743 4824 4745 4864
rect 4749 4824 4751 4864
rect 4763 4824 4765 4864
rect 4769 4824 4771 4864
rect 4819 4824 4821 4904
rect 4825 4824 4827 4904
rect 4839 4824 4843 4864
rect 4847 4824 4851 4864
rect 4863 4824 4865 4864
rect 4869 4824 4871 4864
rect 4923 4824 4925 4864
rect 4929 4824 4931 4864
rect 4943 4824 4945 4864
rect 4949 4824 4951 4864
rect 4989 4824 4991 4864
rect 4995 4824 4997 4864
rect 5009 4824 5011 4864
rect 5015 4824 5017 4864
rect 5069 4824 5071 4864
rect 5075 4824 5077 4864
rect 5089 4824 5093 4864
rect 5097 4824 5101 4864
rect 5113 4824 5115 4904
rect 5119 4824 5121 4904
rect 5183 4824 5185 4864
rect 5189 4824 5191 4864
rect 5203 4824 5205 4864
rect 5209 4824 5211 4864
rect 5259 4824 5261 4904
rect 5265 4824 5267 4904
rect 5279 4824 5283 4864
rect 5287 4824 5291 4864
rect 5303 4824 5305 4864
rect 5309 4824 5311 4864
rect 5349 4824 5351 4864
rect 5355 4824 5357 4864
rect 5369 4824 5373 4864
rect 5377 4824 5381 4864
rect 5393 4824 5395 4904
rect 5399 4824 5401 4904
rect 5463 4824 5465 4904
rect 5469 4836 5471 4904
rect 5483 4836 5485 4904
rect 5469 4824 5485 4836
rect 5489 4902 5505 4904
rect 5489 4824 5491 4902
rect 5503 4824 5505 4902
rect 5509 4890 5525 4904
rect 5509 4824 5511 4890
rect 5523 4824 5525 4890
rect 5529 4902 5543 4904
rect 5529 4824 5531 4902
rect 5583 4824 5585 4864
rect 5589 4824 5591 4864
rect 5603 4824 5605 4864
rect 5609 4824 5611 4864
rect 5649 4824 5651 4864
rect 5655 4824 5657 4864
rect 5669 4824 5671 4864
rect 5675 4860 5691 4864
rect 5675 4824 5677 4860
rect 5689 4824 5691 4860
rect 5695 4824 5697 4864
rect 5763 4824 5765 4904
rect 5769 4824 5771 4904
rect 5783 4824 5785 4904
rect 5789 4892 5805 4904
rect 5789 4824 5791 4892
rect 5803 4824 5805 4892
rect 5809 4896 5823 4904
rect 5809 4824 5811 4896
rect 6017 4902 6031 4904
rect 5863 4824 5865 4864
rect 5869 4860 5885 4864
rect 5869 4824 5871 4860
rect 5883 4824 5885 4860
rect 5889 4824 5891 4864
rect 5903 4824 5905 4864
rect 5909 4824 5911 4864
rect 5963 4824 5965 4864
rect 5969 4824 5971 4864
rect 5983 4824 5985 4864
rect 5989 4824 5991 4864
rect 6029 4824 6031 4902
rect 6035 4890 6051 4904
rect 6035 4824 6037 4890
rect 6049 4824 6051 4890
rect 6055 4902 6071 4904
rect 6055 4824 6057 4902
rect 6069 4824 6071 4902
rect 6075 4836 6077 4904
rect 6089 4836 6091 4904
rect 6075 4824 6091 4836
rect 6095 4824 6097 4904
rect 6163 4824 6165 4864
rect 6169 4860 6185 4864
rect 6169 4824 6171 4860
rect 6183 4824 6185 4860
rect 6189 4824 6191 4864
rect 6203 4824 6205 4864
rect 6209 4824 6211 4864
rect 6254 4824 6256 4904
rect 6260 4824 6264 4904
rect 6268 4824 6270 4904
rect 6282 4824 6286 4864
rect 6290 4824 6292 4864
rect 6363 4824 6365 4864
rect 6369 4860 6385 4864
rect 6369 4824 6371 4860
rect 6383 4824 6385 4860
rect 6389 4824 6391 4864
rect 6403 4824 6405 4864
rect 6409 4824 6411 4864
rect 6463 4824 6465 4864
rect 6469 4860 6485 4864
rect 6469 4824 6471 4860
rect 6483 4824 6485 4860
rect 6489 4824 6491 4864
rect 6503 4824 6505 4864
rect 6509 4824 6511 4864
rect 6549 4824 6551 4864
rect 6555 4824 6557 4864
rect 6569 4824 6571 4864
rect 6575 4824 6577 4864
rect 6643 4824 6645 4864
rect 6649 4824 6651 4864
rect 29 4716 31 4796
rect 35 4716 37 4796
rect 49 4716 51 4796
rect 55 4716 57 4796
rect 69 4716 71 4796
rect 75 4716 77 4796
rect 89 4716 91 4796
rect 95 4716 97 4796
rect 109 4716 111 4796
rect 115 4716 117 4796
rect 129 4716 131 4796
rect 135 4716 137 4796
rect 149 4716 151 4796
rect 155 4716 157 4796
rect 169 4716 171 4796
rect 175 4716 177 4796
rect 255 4716 257 4796
rect 261 4716 265 4796
rect 269 4716 271 4796
rect 323 4756 325 4796
rect 329 4756 331 4796
rect 383 4716 385 4796
rect 389 4716 391 4796
rect 403 4716 405 4796
rect 409 4728 411 4796
rect 423 4728 425 4796
rect 409 4716 425 4728
rect 429 4724 431 4796
rect 483 4756 485 4796
rect 489 4756 491 4796
rect 429 4716 443 4724
rect 555 4716 557 4796
rect 561 4716 565 4796
rect 569 4716 571 4796
rect 619 4716 621 4796
rect 625 4716 627 4796
rect 639 4756 643 4796
rect 647 4756 651 4796
rect 663 4756 665 4796
rect 669 4756 671 4796
rect 709 4716 711 4796
rect 715 4716 719 4796
rect 723 4716 725 4796
rect 801 4716 803 4796
rect 807 4716 809 4796
rect 821 4756 825 4796
rect 829 4756 831 4796
rect 883 4756 885 4796
rect 889 4756 891 4796
rect 903 4756 905 4796
rect 909 4756 911 4796
rect 949 4716 951 4796
rect 955 4776 957 4796
rect 969 4776 973 4796
rect 977 4776 981 4796
rect 985 4776 987 4796
rect 999 4776 1001 4796
rect 955 4716 964 4776
rect 990 4756 1001 4776
rect 1005 4756 1009 4796
rect 1013 4756 1015 4796
rect 1053 4756 1055 4796
rect 1059 4756 1061 4796
rect 1073 4756 1075 4796
rect 1079 4756 1087 4796
rect 1091 4756 1093 4796
rect 1105 4756 1107 4796
rect 1111 4756 1121 4796
rect 1125 4756 1127 4796
rect 1139 4756 1141 4796
rect 1132 4716 1141 4756
rect 1145 4716 1147 4796
rect 1208 4756 1210 4796
rect 1214 4756 1218 4796
rect 1230 4716 1232 4796
rect 1236 4716 1240 4796
rect 1244 4716 1246 4796
rect 1303 4756 1305 4796
rect 1309 4756 1311 4796
rect 1323 4756 1325 4796
rect 1329 4756 1331 4796
rect 1369 4756 1371 4796
rect 1375 4756 1377 4796
rect 1389 4756 1391 4796
rect 1395 4756 1397 4796
rect 1468 4756 1470 4796
rect 1474 4756 1478 4796
rect 1490 4716 1492 4796
rect 1496 4716 1500 4796
rect 1504 4716 1506 4796
rect 1549 4716 1551 4796
rect 1555 4716 1559 4796
rect 1563 4716 1565 4796
rect 1629 4716 1631 4796
rect 1635 4716 1639 4796
rect 1643 4716 1645 4796
rect 1709 4756 1711 4796
rect 1715 4756 1717 4796
rect 1769 4716 1771 4796
rect 1775 4716 1779 4796
rect 1783 4716 1785 4796
rect 1854 4716 1856 4796
rect 1860 4716 1864 4796
rect 1868 4716 1870 4796
rect 1882 4756 1886 4796
rect 1890 4756 1892 4796
rect 1949 4716 1951 4796
rect 1955 4776 1957 4796
rect 1969 4776 1973 4796
rect 1977 4776 1981 4796
rect 1985 4776 1987 4796
rect 1999 4776 2001 4796
rect 1955 4716 1964 4776
rect 1990 4756 2001 4776
rect 2005 4756 2009 4796
rect 2013 4756 2015 4796
rect 2053 4756 2055 4796
rect 2059 4756 2061 4796
rect 2073 4756 2075 4796
rect 2079 4756 2087 4796
rect 2091 4756 2093 4796
rect 2105 4756 2107 4796
rect 2111 4756 2121 4796
rect 2125 4756 2127 4796
rect 2139 4756 2141 4796
rect 2132 4716 2141 4756
rect 2145 4716 2147 4796
rect 2203 4756 2205 4796
rect 2209 4756 2211 4796
rect 2223 4756 2225 4796
rect 2229 4756 2231 4796
rect 2293 4717 2295 4796
rect 2281 4716 2295 4717
rect 2299 4717 2301 4796
rect 2313 4717 2315 4796
rect 2299 4716 2315 4717
rect 2319 4716 2325 4796
rect 2329 4716 2331 4796
rect 2369 4756 2371 4796
rect 2375 4756 2377 4796
rect 2389 4756 2391 4796
rect 2395 4756 2397 4796
rect 2449 4716 2451 4796
rect 2455 4716 2459 4796
rect 2463 4716 2465 4796
rect 2529 4724 2531 4796
rect 2517 4716 2531 4724
rect 2535 4728 2537 4796
rect 2549 4728 2551 4796
rect 2535 4716 2551 4728
rect 2555 4716 2557 4796
rect 2569 4716 2571 4796
rect 2575 4716 2577 4796
rect 2643 4756 2645 4796
rect 2649 4756 2651 4796
rect 2689 4716 2691 4796
rect 2695 4776 2697 4796
rect 2709 4776 2713 4796
rect 2717 4776 2721 4796
rect 2725 4776 2727 4796
rect 2739 4776 2741 4796
rect 2695 4716 2704 4776
rect 2730 4756 2741 4776
rect 2745 4756 2749 4796
rect 2753 4756 2755 4796
rect 2793 4756 2795 4796
rect 2799 4756 2801 4796
rect 2813 4756 2815 4796
rect 2819 4756 2827 4796
rect 2831 4756 2833 4796
rect 2845 4756 2847 4796
rect 2851 4756 2861 4796
rect 2865 4756 2867 4796
rect 2879 4756 2881 4796
rect 2872 4716 2881 4756
rect 2885 4716 2887 4796
rect 2934 4716 2936 4796
rect 2940 4716 2944 4796
rect 2948 4716 2950 4796
rect 2962 4756 2966 4796
rect 2970 4756 2972 4796
rect 3029 4716 3031 4796
rect 3035 4776 3037 4796
rect 3049 4776 3053 4796
rect 3057 4776 3061 4796
rect 3065 4776 3067 4796
rect 3079 4776 3081 4796
rect 3035 4716 3044 4776
rect 3070 4756 3081 4776
rect 3085 4756 3089 4796
rect 3093 4756 3095 4796
rect 3133 4756 3135 4796
rect 3139 4756 3141 4796
rect 3153 4756 3155 4796
rect 3159 4756 3167 4796
rect 3171 4756 3173 4796
rect 3185 4756 3187 4796
rect 3191 4756 3201 4796
rect 3205 4756 3207 4796
rect 3219 4756 3221 4796
rect 3212 4716 3221 4756
rect 3225 4716 3227 4796
rect 3269 4716 3271 4796
rect 3275 4776 3277 4796
rect 3289 4776 3293 4796
rect 3297 4776 3301 4796
rect 3305 4776 3307 4796
rect 3319 4776 3321 4796
rect 3275 4716 3284 4776
rect 3310 4756 3321 4776
rect 3325 4756 3329 4796
rect 3333 4756 3335 4796
rect 3373 4756 3375 4796
rect 3379 4756 3381 4796
rect 3393 4756 3395 4796
rect 3399 4756 3407 4796
rect 3411 4756 3413 4796
rect 3425 4756 3427 4796
rect 3431 4756 3441 4796
rect 3445 4756 3447 4796
rect 3459 4756 3461 4796
rect 3452 4716 3461 4756
rect 3465 4716 3467 4796
rect 3528 4756 3530 4796
rect 3534 4756 3538 4796
rect 3550 4716 3552 4796
rect 3556 4716 3560 4796
rect 3564 4716 3566 4796
rect 3623 4716 3625 4796
rect 3629 4716 3631 4796
rect 3683 4756 3685 4796
rect 3689 4756 3691 4796
rect 3703 4756 3705 4796
rect 3709 4756 3711 4796
rect 3768 4756 3770 4796
rect 3774 4756 3778 4796
rect 3790 4716 3792 4796
rect 3796 4716 3800 4796
rect 3804 4716 3806 4796
rect 3853 4716 3855 4796
rect 3859 4756 3861 4796
rect 3873 4756 3875 4796
rect 3879 4756 3889 4796
rect 3893 4756 3895 4796
rect 3907 4756 3909 4796
rect 3913 4756 3921 4796
rect 3925 4756 3927 4796
rect 3939 4756 3941 4796
rect 3945 4756 3947 4796
rect 3985 4756 3987 4796
rect 3991 4756 3995 4796
rect 3999 4776 4001 4796
rect 4013 4776 4015 4796
rect 4019 4776 4023 4796
rect 4027 4776 4031 4796
rect 4043 4776 4045 4796
rect 3999 4756 4010 4776
rect 3859 4716 3868 4756
rect 4036 4716 4045 4776
rect 4049 4716 4051 4796
rect 4103 4716 4105 4796
rect 4109 4716 4111 4796
rect 4163 4756 4165 4796
rect 4169 4756 4171 4796
rect 4183 4756 4185 4796
rect 4189 4756 4191 4796
rect 4229 4716 4231 4796
rect 4235 4776 4237 4796
rect 4249 4776 4253 4796
rect 4257 4776 4261 4796
rect 4265 4776 4267 4796
rect 4279 4776 4281 4796
rect 4235 4716 4244 4776
rect 4270 4756 4281 4776
rect 4285 4756 4289 4796
rect 4293 4756 4295 4796
rect 4333 4756 4335 4796
rect 4339 4756 4341 4796
rect 4353 4756 4355 4796
rect 4359 4756 4367 4796
rect 4371 4756 4373 4796
rect 4385 4756 4387 4796
rect 4391 4756 4401 4796
rect 4405 4756 4407 4796
rect 4419 4756 4421 4796
rect 4412 4716 4421 4756
rect 4425 4716 4427 4796
rect 4483 4756 4485 4796
rect 4489 4760 4491 4796
rect 4503 4760 4505 4796
rect 4489 4756 4505 4760
rect 4509 4756 4511 4796
rect 4523 4756 4525 4796
rect 4529 4756 4531 4796
rect 4569 4756 4571 4796
rect 4575 4756 4577 4796
rect 4629 4716 4631 4796
rect 4635 4716 4637 4796
rect 4703 4756 4705 4796
rect 4709 4756 4711 4796
rect 4754 4716 4756 4796
rect 4760 4716 4764 4796
rect 4768 4716 4770 4796
rect 4782 4756 4786 4796
rect 4790 4756 4792 4796
rect 4849 4716 4851 4796
rect 4855 4716 4859 4796
rect 4863 4716 4865 4796
rect 4929 4756 4931 4796
rect 4935 4756 4937 4796
rect 4949 4756 4951 4796
rect 4955 4756 4957 4796
rect 5009 4756 5011 4796
rect 5015 4756 5017 4796
rect 5029 4756 5031 4796
rect 5035 4756 5037 4796
rect 5103 4756 5105 4796
rect 5109 4756 5111 4796
rect 5123 4756 5125 4796
rect 5129 4756 5131 4796
rect 5174 4716 5176 4796
rect 5180 4716 5184 4796
rect 5188 4716 5190 4796
rect 5202 4756 5206 4796
rect 5210 4756 5212 4796
rect 5293 4716 5295 4796
rect 5299 4716 5305 4796
rect 5309 4716 5311 4796
rect 5333 4716 5335 4796
rect 5339 4716 5345 4796
rect 5349 4716 5351 4796
rect 5389 4756 5391 4796
rect 5395 4756 5397 4796
rect 5409 4756 5411 4796
rect 5415 4756 5417 4796
rect 5483 4756 5485 4796
rect 5489 4756 5491 4796
rect 5503 4756 5505 4796
rect 5509 4756 5511 4796
rect 5549 4756 5551 4796
rect 5555 4756 5557 4796
rect 5569 4756 5571 4796
rect 5575 4760 5577 4796
rect 5589 4760 5591 4796
rect 5575 4756 5591 4760
rect 5595 4756 5597 4796
rect 5663 4756 5665 4796
rect 5669 4756 5671 4796
rect 5683 4756 5685 4796
rect 5689 4756 5691 4796
rect 5729 4756 5731 4796
rect 5735 4756 5737 4796
rect 5749 4756 5751 4796
rect 5755 4760 5757 4796
rect 5769 4760 5771 4796
rect 5755 4756 5771 4760
rect 5775 4756 5777 4796
rect 5843 4756 5845 4796
rect 5849 4756 5851 4796
rect 5889 4756 5891 4796
rect 5895 4756 5897 4796
rect 5909 4756 5911 4796
rect 5915 4760 5917 4796
rect 5929 4760 5931 4796
rect 5915 4756 5931 4760
rect 5935 4756 5937 4796
rect 5999 4716 6001 4796
rect 6005 4716 6007 4796
rect 6019 4756 6023 4796
rect 6027 4756 6031 4796
rect 6043 4756 6045 4796
rect 6049 4756 6051 4796
rect 6094 4716 6096 4796
rect 6100 4716 6104 4796
rect 6108 4716 6110 4796
rect 6122 4756 6126 4796
rect 6130 4756 6132 4796
rect 6203 4756 6205 4796
rect 6209 4756 6211 4796
rect 6223 4756 6225 4796
rect 6229 4756 6231 4796
rect 6269 4724 6271 4796
rect 6257 4716 6271 4724
rect 6275 4728 6277 4796
rect 6289 4728 6291 4796
rect 6275 4716 6291 4728
rect 6295 4716 6297 4796
rect 6309 4716 6311 4796
rect 6315 4716 6317 4796
rect 6369 4756 6371 4796
rect 6375 4756 6377 4796
rect 6389 4756 6391 4796
rect 6395 4760 6397 4796
rect 6409 4760 6411 4796
rect 6395 4756 6411 4760
rect 6415 4756 6417 4796
rect 6479 4716 6481 4796
rect 6485 4716 6487 4796
rect 6499 4756 6503 4796
rect 6507 4756 6511 4796
rect 6523 4756 6525 4796
rect 6529 4756 6531 4796
rect 6583 4756 6585 4796
rect 6589 4760 6591 4796
rect 6603 4760 6605 4796
rect 6589 4756 6605 4760
rect 6609 4756 6611 4796
rect 6623 4756 6625 4796
rect 6629 4756 6631 4796
rect 43 4344 45 4384
rect 49 4344 51 4384
rect 115 4344 117 4424
rect 121 4344 125 4424
rect 129 4344 131 4424
rect 183 4344 185 4384
rect 189 4344 191 4384
rect 234 4344 236 4424
rect 240 4344 244 4424
rect 248 4344 250 4424
rect 262 4344 266 4384
rect 270 4344 272 4384
rect 355 4344 357 4424
rect 361 4344 365 4424
rect 369 4344 371 4424
rect 414 4344 416 4424
rect 420 4344 424 4424
rect 428 4344 430 4424
rect 442 4344 446 4384
rect 450 4344 452 4384
rect 509 4344 511 4424
rect 515 4344 521 4424
rect 525 4423 541 4424
rect 525 4344 527 4423
rect 539 4344 541 4423
rect 545 4423 559 4424
rect 545 4344 547 4423
rect 597 4416 611 4424
rect 609 4344 611 4416
rect 615 4412 631 4424
rect 615 4344 617 4412
rect 629 4344 631 4412
rect 635 4344 637 4424
rect 649 4344 651 4424
rect 655 4344 657 4424
rect 723 4344 725 4384
rect 729 4344 731 4384
rect 769 4344 771 4424
rect 775 4344 779 4424
rect 783 4344 785 4424
rect 849 4344 851 4384
rect 855 4344 857 4384
rect 909 4344 911 4424
rect 915 4344 919 4424
rect 923 4344 925 4424
rect 989 4344 991 4384
rect 995 4344 997 4384
rect 1049 4344 1051 4424
rect 1055 4344 1057 4424
rect 1069 4344 1071 4424
rect 1075 4344 1077 4424
rect 1089 4344 1091 4424
rect 1095 4344 1097 4424
rect 1109 4344 1111 4424
rect 1115 4344 1117 4424
rect 1129 4344 1131 4424
rect 1135 4344 1137 4424
rect 1149 4344 1151 4424
rect 1155 4344 1157 4424
rect 1169 4344 1171 4424
rect 1175 4344 1177 4424
rect 1189 4344 1191 4424
rect 1195 4344 1197 4424
rect 1249 4344 1251 4384
rect 1255 4344 1259 4384
rect 1271 4344 1273 4424
rect 1277 4344 1279 4424
rect 1343 4344 1345 4384
rect 1349 4344 1351 4384
rect 1415 4344 1417 4424
rect 1421 4344 1425 4424
rect 1429 4344 1431 4424
rect 1483 4344 1485 4384
rect 1489 4344 1491 4384
rect 1503 4344 1505 4384
rect 1509 4344 1511 4384
rect 1549 4344 1551 4384
rect 1555 4344 1557 4384
rect 1569 4344 1571 4384
rect 1575 4344 1577 4384
rect 1643 4344 1645 4424
rect 1649 4344 1651 4424
rect 1663 4344 1665 4424
rect 1669 4344 1671 4424
rect 1683 4344 1685 4424
rect 1689 4344 1691 4424
rect 1703 4344 1705 4424
rect 1709 4344 1711 4424
rect 1753 4344 1755 4424
rect 1759 4384 1768 4424
rect 1759 4344 1761 4384
rect 1773 4344 1775 4384
rect 1779 4344 1789 4384
rect 1793 4344 1795 4384
rect 1807 4344 1809 4384
rect 1813 4344 1821 4384
rect 1825 4344 1827 4384
rect 1839 4344 1841 4384
rect 1845 4344 1847 4384
rect 1885 4344 1887 4384
rect 1891 4344 1895 4384
rect 1899 4364 1910 4384
rect 1936 4364 1945 4424
rect 1899 4344 1901 4364
rect 1913 4344 1915 4364
rect 1919 4344 1923 4364
rect 1927 4344 1931 4364
rect 1943 4344 1945 4364
rect 1949 4344 1951 4424
rect 1989 4344 1991 4384
rect 1995 4344 1997 4384
rect 2009 4344 2011 4384
rect 2015 4344 2017 4384
rect 2069 4344 2071 4424
rect 2075 4364 2084 4424
rect 2252 4384 2261 4424
rect 2110 4364 2121 4384
rect 2075 4344 2077 4364
rect 2089 4344 2093 4364
rect 2097 4344 2101 4364
rect 2105 4344 2107 4364
rect 2119 4344 2121 4364
rect 2125 4344 2129 4384
rect 2133 4344 2135 4384
rect 2173 4344 2175 4384
rect 2179 4344 2181 4384
rect 2193 4344 2195 4384
rect 2199 4344 2207 4384
rect 2211 4344 2213 4384
rect 2225 4344 2227 4384
rect 2231 4344 2241 4384
rect 2245 4344 2247 4384
rect 2259 4344 2261 4384
rect 2265 4344 2267 4424
rect 2309 4344 2311 4384
rect 2315 4344 2317 4384
rect 2369 4344 2371 4424
rect 2375 4344 2379 4424
rect 2383 4344 2385 4424
rect 2449 4344 2451 4424
rect 2455 4344 2459 4424
rect 2463 4344 2465 4424
rect 2529 4344 2531 4384
rect 2535 4344 2537 4384
rect 2589 4344 2591 4424
rect 2595 4364 2604 4424
rect 2772 4384 2781 4424
rect 2630 4364 2641 4384
rect 2595 4344 2597 4364
rect 2609 4344 2613 4364
rect 2617 4344 2621 4364
rect 2625 4344 2627 4364
rect 2639 4344 2641 4364
rect 2645 4344 2649 4384
rect 2653 4344 2655 4384
rect 2693 4344 2695 4384
rect 2699 4344 2701 4384
rect 2713 4344 2715 4384
rect 2719 4344 2727 4384
rect 2731 4344 2733 4384
rect 2745 4344 2747 4384
rect 2751 4344 2761 4384
rect 2765 4344 2767 4384
rect 2779 4344 2781 4384
rect 2785 4344 2787 4424
rect 2834 4344 2836 4424
rect 2840 4344 2844 4424
rect 2848 4344 2850 4424
rect 2862 4344 2866 4384
rect 2870 4344 2872 4384
rect 2929 4344 2931 4384
rect 2935 4344 2937 4384
rect 2949 4344 2951 4384
rect 2955 4344 2957 4384
rect 3023 4344 3025 4384
rect 3029 4344 3031 4384
rect 3074 4344 3076 4424
rect 3080 4344 3084 4424
rect 3088 4344 3090 4424
rect 3102 4344 3106 4384
rect 3110 4344 3112 4384
rect 3169 4344 3171 4424
rect 3175 4364 3184 4424
rect 3352 4384 3361 4424
rect 3210 4364 3221 4384
rect 3175 4344 3177 4364
rect 3189 4344 3193 4364
rect 3197 4344 3201 4364
rect 3205 4344 3207 4364
rect 3219 4344 3221 4364
rect 3225 4344 3229 4384
rect 3233 4344 3235 4384
rect 3273 4344 3275 4384
rect 3279 4344 3281 4384
rect 3293 4344 3295 4384
rect 3299 4344 3307 4384
rect 3311 4344 3313 4384
rect 3325 4344 3327 4384
rect 3331 4344 3341 4384
rect 3345 4344 3347 4384
rect 3359 4344 3361 4384
rect 3365 4344 3367 4424
rect 3414 4344 3416 4424
rect 3420 4344 3424 4424
rect 3428 4344 3430 4424
rect 3442 4344 3446 4384
rect 3450 4344 3452 4384
rect 3528 4344 3530 4384
rect 3534 4344 3538 4384
rect 3550 4344 3552 4424
rect 3556 4344 3560 4424
rect 3564 4344 3566 4424
rect 3613 4344 3615 4424
rect 3619 4384 3628 4424
rect 3619 4344 3621 4384
rect 3633 4344 3635 4384
rect 3639 4344 3649 4384
rect 3653 4344 3655 4384
rect 3667 4344 3669 4384
rect 3673 4344 3681 4384
rect 3685 4344 3687 4384
rect 3699 4344 3701 4384
rect 3705 4344 3707 4384
rect 3745 4344 3747 4384
rect 3751 4344 3755 4384
rect 3759 4364 3770 4384
rect 3796 4364 3805 4424
rect 3759 4344 3761 4364
rect 3773 4344 3775 4364
rect 3779 4344 3783 4364
rect 3787 4344 3791 4364
rect 3803 4344 3805 4364
rect 3809 4344 3811 4424
rect 3854 4344 3856 4424
rect 3860 4344 3864 4424
rect 3868 4344 3870 4424
rect 3882 4344 3886 4384
rect 3890 4344 3892 4384
rect 3953 4344 3955 4424
rect 3959 4384 3968 4424
rect 3959 4344 3961 4384
rect 3973 4344 3975 4384
rect 3979 4344 3989 4384
rect 3993 4344 3995 4384
rect 4007 4344 4009 4384
rect 4013 4344 4021 4384
rect 4025 4344 4027 4384
rect 4039 4344 4041 4384
rect 4045 4344 4047 4384
rect 4085 4344 4087 4384
rect 4091 4344 4095 4384
rect 4099 4364 4110 4384
rect 4136 4364 4145 4424
rect 4099 4344 4101 4364
rect 4113 4344 4115 4364
rect 4119 4344 4123 4364
rect 4127 4344 4131 4364
rect 4143 4344 4145 4364
rect 4149 4344 4151 4424
rect 4203 4344 4205 4384
rect 4209 4380 4225 4384
rect 4209 4344 4211 4380
rect 4223 4344 4225 4380
rect 4229 4344 4231 4384
rect 4243 4344 4245 4384
rect 4249 4344 4251 4384
rect 4294 4344 4296 4424
rect 4300 4344 4304 4424
rect 4308 4344 4310 4424
rect 4322 4344 4326 4384
rect 4330 4344 4332 4384
rect 4415 4344 4417 4424
rect 4421 4344 4425 4424
rect 4429 4344 4431 4424
rect 4483 4344 4485 4424
rect 4489 4344 4491 4424
rect 4503 4344 4505 4424
rect 4509 4412 4525 4424
rect 4509 4344 4511 4412
rect 4523 4344 4525 4412
rect 4529 4416 4543 4424
rect 4529 4344 4531 4416
rect 4569 4344 4571 4384
rect 4575 4344 4577 4384
rect 4589 4344 4591 4384
rect 4595 4380 4611 4384
rect 4595 4344 4597 4380
rect 4609 4344 4611 4380
rect 4615 4344 4617 4384
rect 4683 4344 4685 4384
rect 4689 4344 4691 4384
rect 4734 4344 4736 4424
rect 4740 4344 4744 4424
rect 4748 4344 4750 4424
rect 4841 4423 4855 4424
rect 4762 4344 4766 4384
rect 4770 4344 4772 4384
rect 4853 4344 4855 4423
rect 4859 4423 4875 4424
rect 4859 4344 4861 4423
rect 4873 4344 4875 4423
rect 4879 4344 4885 4424
rect 4889 4344 4891 4424
rect 4943 4344 4945 4384
rect 4949 4344 4951 4384
rect 4963 4344 4965 4384
rect 4969 4344 4971 4384
rect 5023 4344 5025 4384
rect 5029 4380 5045 4384
rect 5029 4344 5031 4380
rect 5043 4344 5045 4380
rect 5049 4344 5051 4384
rect 5063 4344 5065 4384
rect 5069 4344 5071 4384
rect 5114 4344 5116 4424
rect 5120 4344 5124 4424
rect 5128 4344 5130 4424
rect 5221 4423 5235 4424
rect 5142 4344 5146 4384
rect 5150 4344 5152 4384
rect 5233 4344 5235 4423
rect 5239 4423 5255 4424
rect 5239 4344 5241 4423
rect 5253 4344 5255 4423
rect 5259 4344 5265 4424
rect 5269 4344 5271 4424
rect 5314 4344 5316 4424
rect 5320 4344 5324 4424
rect 5328 4344 5330 4424
rect 5342 4344 5346 4384
rect 5350 4344 5352 4384
rect 5409 4344 5411 4384
rect 5415 4344 5417 4384
rect 5483 4344 5485 4384
rect 5489 4380 5505 4384
rect 5489 4344 5491 4380
rect 5503 4344 5505 4380
rect 5509 4344 5511 4384
rect 5523 4344 5525 4384
rect 5529 4344 5531 4384
rect 5569 4344 5571 4384
rect 5575 4344 5577 4384
rect 5589 4344 5591 4384
rect 5595 4344 5597 4384
rect 5654 4344 5656 4424
rect 5660 4344 5664 4424
rect 5668 4344 5670 4424
rect 5682 4344 5686 4384
rect 5690 4344 5692 4384
rect 5763 4344 5765 4384
rect 5769 4344 5771 4384
rect 5783 4344 5785 4384
rect 5789 4344 5791 4384
rect 5843 4344 5845 4384
rect 5849 4380 5865 4384
rect 5849 4344 5851 4380
rect 5863 4344 5865 4380
rect 5869 4344 5871 4384
rect 5883 4344 5885 4384
rect 5889 4344 5891 4384
rect 5948 4344 5950 4384
rect 5954 4344 5958 4384
rect 5970 4344 5972 4424
rect 5976 4344 5980 4424
rect 5984 4344 5986 4424
rect 6029 4344 6031 4384
rect 6035 4344 6037 4384
rect 6103 4344 6105 4384
rect 6109 4344 6111 4384
rect 6149 4344 6151 4384
rect 6155 4344 6157 4384
rect 6169 4344 6171 4384
rect 6175 4380 6191 4384
rect 6175 4344 6177 4380
rect 6189 4344 6191 4380
rect 6195 4344 6197 4384
rect 6268 4344 6270 4384
rect 6274 4344 6278 4384
rect 6290 4344 6292 4424
rect 6296 4344 6300 4424
rect 6304 4344 6306 4424
rect 6349 4344 6351 4384
rect 6355 4344 6357 4384
rect 6369 4344 6371 4384
rect 6375 4380 6391 4384
rect 6375 4344 6377 4380
rect 6389 4344 6391 4380
rect 6395 4344 6397 4384
rect 6449 4344 6451 4384
rect 6455 4344 6457 4384
rect 6469 4344 6471 4384
rect 6475 4380 6491 4384
rect 6475 4344 6477 4380
rect 6489 4344 6491 4380
rect 6495 4344 6497 4384
rect 6554 4344 6556 4424
rect 6560 4344 6564 4424
rect 6568 4344 6570 4424
rect 6582 4344 6586 4384
rect 6590 4344 6592 4384
rect 6649 4344 6651 4384
rect 6655 4344 6657 4384
rect 41 4236 43 4316
rect 47 4236 49 4316
rect 61 4276 65 4316
rect 69 4276 71 4316
rect 128 4276 130 4316
rect 134 4276 138 4316
rect 150 4236 152 4316
rect 156 4236 160 4316
rect 164 4236 166 4316
rect 214 4236 216 4316
rect 220 4236 224 4316
rect 228 4236 230 4316
rect 242 4276 246 4316
rect 250 4276 252 4316
rect 313 4236 315 4316
rect 319 4276 321 4316
rect 333 4276 335 4316
rect 339 4276 349 4316
rect 353 4276 355 4316
rect 367 4276 369 4316
rect 373 4276 381 4316
rect 385 4276 387 4316
rect 399 4276 401 4316
rect 405 4276 407 4316
rect 445 4276 447 4316
rect 451 4276 455 4316
rect 459 4296 461 4316
rect 473 4296 475 4316
rect 479 4296 483 4316
rect 487 4296 491 4316
rect 503 4296 505 4316
rect 459 4276 470 4296
rect 319 4236 328 4276
rect 496 4236 505 4296
rect 509 4236 511 4316
rect 549 4276 551 4316
rect 555 4276 557 4316
rect 569 4276 571 4316
rect 575 4276 577 4316
rect 643 4236 645 4316
rect 649 4304 665 4316
rect 649 4236 651 4304
rect 663 4236 665 4304
rect 669 4238 671 4316
rect 683 4238 685 4316
rect 669 4236 685 4238
rect 689 4250 691 4316
rect 703 4250 705 4316
rect 689 4236 705 4250
rect 709 4238 711 4316
rect 763 4276 765 4316
rect 769 4276 771 4316
rect 709 4236 723 4238
rect 809 4236 811 4316
rect 815 4296 817 4316
rect 829 4296 833 4316
rect 837 4296 841 4316
rect 845 4296 847 4316
rect 859 4296 861 4316
rect 815 4236 824 4296
rect 850 4276 861 4296
rect 865 4276 869 4316
rect 873 4276 875 4316
rect 913 4276 915 4316
rect 919 4276 921 4316
rect 933 4276 935 4316
rect 939 4276 947 4316
rect 951 4276 953 4316
rect 965 4276 967 4316
rect 971 4276 981 4316
rect 985 4276 987 4316
rect 999 4276 1001 4316
rect 992 4236 1001 4276
rect 1005 4236 1007 4316
rect 1049 4276 1051 4316
rect 1055 4276 1057 4316
rect 1069 4276 1071 4316
rect 1075 4276 1077 4316
rect 1129 4236 1131 4316
rect 1135 4296 1137 4316
rect 1149 4296 1153 4316
rect 1157 4296 1161 4316
rect 1165 4296 1167 4316
rect 1179 4296 1181 4316
rect 1135 4236 1144 4296
rect 1170 4276 1181 4296
rect 1185 4276 1189 4316
rect 1193 4276 1195 4316
rect 1233 4276 1235 4316
rect 1239 4276 1241 4316
rect 1253 4276 1255 4316
rect 1259 4276 1267 4316
rect 1271 4276 1273 4316
rect 1285 4276 1287 4316
rect 1291 4276 1301 4316
rect 1305 4276 1307 4316
rect 1319 4276 1321 4316
rect 1312 4236 1321 4276
rect 1325 4236 1327 4316
rect 1369 4276 1371 4316
rect 1375 4276 1377 4316
rect 1389 4276 1391 4316
rect 1395 4276 1397 4316
rect 1449 4276 1451 4316
rect 1455 4276 1457 4316
rect 1528 4276 1530 4316
rect 1534 4276 1538 4316
rect 1550 4236 1552 4316
rect 1556 4236 1560 4316
rect 1564 4236 1566 4316
rect 1623 4236 1625 4316
rect 1629 4236 1631 4316
rect 1643 4236 1645 4316
rect 1649 4248 1651 4316
rect 1663 4248 1665 4316
rect 1649 4236 1665 4248
rect 1669 4244 1671 4316
rect 1723 4276 1725 4316
rect 1729 4276 1731 4316
rect 1743 4276 1745 4316
rect 1749 4276 1751 4316
rect 1789 4276 1791 4316
rect 1795 4276 1797 4316
rect 1809 4276 1811 4316
rect 1815 4276 1817 4316
rect 1669 4236 1683 4244
rect 1869 4236 1871 4316
rect 1875 4296 1877 4316
rect 1889 4296 1893 4316
rect 1897 4296 1901 4316
rect 1905 4296 1907 4316
rect 1919 4296 1921 4316
rect 1875 4236 1884 4296
rect 1910 4276 1921 4296
rect 1925 4276 1929 4316
rect 1933 4276 1935 4316
rect 1973 4276 1975 4316
rect 1979 4276 1981 4316
rect 1993 4276 1995 4316
rect 1999 4276 2007 4316
rect 2011 4276 2013 4316
rect 2025 4276 2027 4316
rect 2031 4276 2041 4316
rect 2045 4276 2047 4316
rect 2059 4276 2061 4316
rect 2052 4236 2061 4276
rect 2065 4236 2067 4316
rect 2109 4276 2111 4316
rect 2115 4276 2117 4316
rect 2129 4276 2131 4316
rect 2135 4276 2137 4316
rect 2208 4276 2210 4316
rect 2214 4276 2218 4316
rect 2230 4236 2232 4316
rect 2236 4236 2240 4316
rect 2244 4236 2246 4316
rect 2293 4236 2295 4316
rect 2299 4276 2301 4316
rect 2313 4276 2315 4316
rect 2319 4276 2329 4316
rect 2333 4276 2335 4316
rect 2347 4276 2349 4316
rect 2353 4276 2361 4316
rect 2365 4276 2367 4316
rect 2379 4276 2381 4316
rect 2385 4276 2387 4316
rect 2425 4276 2427 4316
rect 2431 4276 2435 4316
rect 2439 4296 2441 4316
rect 2453 4296 2455 4316
rect 2459 4296 2463 4316
rect 2467 4296 2471 4316
rect 2483 4296 2485 4316
rect 2439 4276 2450 4296
rect 2299 4236 2308 4276
rect 2476 4236 2485 4296
rect 2489 4236 2491 4316
rect 2555 4236 2557 4316
rect 2561 4236 2565 4316
rect 2569 4236 2571 4316
rect 2609 4276 2611 4316
rect 2615 4276 2617 4316
rect 2674 4236 2676 4316
rect 2680 4236 2684 4316
rect 2688 4236 2690 4316
rect 2702 4276 2706 4316
rect 2710 4276 2712 4316
rect 2769 4276 2771 4316
rect 2775 4276 2777 4316
rect 2789 4276 2791 4316
rect 2795 4276 2797 4316
rect 2868 4276 2870 4316
rect 2874 4276 2878 4316
rect 2890 4236 2892 4316
rect 2896 4236 2900 4316
rect 2904 4236 2906 4316
rect 2949 4276 2951 4316
rect 2955 4276 2957 4316
rect 3009 4236 3011 4316
rect 3015 4236 3019 4316
rect 3023 4236 3025 4316
rect 3103 4276 3105 4316
rect 3109 4276 3111 4316
rect 3149 4236 3151 4316
rect 3155 4296 3157 4316
rect 3169 4296 3173 4316
rect 3177 4296 3181 4316
rect 3185 4296 3187 4316
rect 3199 4296 3201 4316
rect 3155 4236 3164 4296
rect 3190 4276 3201 4296
rect 3205 4276 3209 4316
rect 3213 4276 3215 4316
rect 3253 4276 3255 4316
rect 3259 4276 3261 4316
rect 3273 4276 3275 4316
rect 3279 4276 3287 4316
rect 3291 4276 3293 4316
rect 3305 4276 3307 4316
rect 3311 4276 3321 4316
rect 3325 4276 3327 4316
rect 3339 4276 3341 4316
rect 3332 4236 3341 4276
rect 3345 4236 3347 4316
rect 3389 4236 3391 4316
rect 3395 4236 3401 4316
rect 3405 4236 3407 4316
rect 3429 4236 3431 4316
rect 3435 4236 3441 4316
rect 3445 4236 3447 4316
rect 3509 4276 3511 4316
rect 3515 4276 3517 4316
rect 3529 4276 3531 4316
rect 3535 4276 3537 4316
rect 3589 4236 3591 4316
rect 3595 4236 3597 4316
rect 3609 4236 3611 4316
rect 3615 4236 3617 4316
rect 3629 4236 3631 4316
rect 3635 4236 3637 4316
rect 3649 4236 3651 4316
rect 3655 4236 3657 4316
rect 3669 4236 3671 4316
rect 3675 4236 3677 4316
rect 3689 4236 3691 4316
rect 3695 4236 3697 4316
rect 3709 4236 3711 4316
rect 3715 4236 3717 4316
rect 3729 4236 3731 4316
rect 3735 4236 3737 4316
rect 3789 4276 3791 4316
rect 3795 4276 3797 4316
rect 3809 4276 3811 4316
rect 3815 4276 3817 4316
rect 3869 4276 3871 4316
rect 3875 4276 3877 4316
rect 3889 4276 3891 4316
rect 3895 4276 3897 4316
rect 3963 4276 3965 4316
rect 3969 4276 3971 4316
rect 3983 4276 3985 4316
rect 3989 4276 3991 4316
rect 4029 4276 4031 4316
rect 4035 4276 4037 4316
rect 4108 4276 4110 4316
rect 4114 4276 4118 4316
rect 4130 4236 4132 4316
rect 4136 4236 4140 4316
rect 4144 4236 4146 4316
rect 4194 4236 4196 4316
rect 4200 4236 4204 4316
rect 4208 4236 4210 4316
rect 4222 4276 4226 4316
rect 4230 4276 4232 4316
rect 4293 4236 4295 4316
rect 4299 4276 4301 4316
rect 4313 4276 4315 4316
rect 4319 4276 4329 4316
rect 4333 4276 4335 4316
rect 4347 4276 4349 4316
rect 4353 4276 4361 4316
rect 4365 4276 4367 4316
rect 4379 4276 4381 4316
rect 4385 4276 4387 4316
rect 4425 4276 4427 4316
rect 4431 4276 4435 4316
rect 4439 4296 4441 4316
rect 4453 4296 4455 4316
rect 4459 4296 4463 4316
rect 4467 4296 4471 4316
rect 4483 4296 4485 4316
rect 4439 4276 4450 4296
rect 4299 4236 4308 4276
rect 4476 4236 4485 4296
rect 4489 4236 4491 4316
rect 4548 4276 4550 4316
rect 4554 4276 4558 4316
rect 4570 4236 4572 4316
rect 4576 4236 4580 4316
rect 4584 4236 4586 4316
rect 4633 4236 4635 4316
rect 4639 4276 4641 4316
rect 4653 4276 4655 4316
rect 4659 4276 4669 4316
rect 4673 4276 4675 4316
rect 4687 4276 4689 4316
rect 4693 4276 4701 4316
rect 4705 4276 4707 4316
rect 4719 4276 4721 4316
rect 4725 4276 4727 4316
rect 4765 4276 4767 4316
rect 4771 4276 4775 4316
rect 4779 4296 4781 4316
rect 4793 4296 4795 4316
rect 4799 4296 4803 4316
rect 4807 4296 4811 4316
rect 4823 4296 4825 4316
rect 4779 4276 4790 4296
rect 4639 4236 4648 4276
rect 4816 4236 4825 4296
rect 4829 4236 4831 4316
rect 4883 4236 4885 4316
rect 4889 4236 4891 4316
rect 4943 4236 4945 4316
rect 4949 4236 4951 4316
rect 4963 4236 4965 4316
rect 4969 4248 4971 4316
rect 4983 4248 4985 4316
rect 4969 4236 4985 4248
rect 4989 4244 4991 4316
rect 5029 4276 5031 4316
rect 5035 4276 5037 4316
rect 5049 4276 5051 4316
rect 5055 4280 5057 4316
rect 5069 4280 5071 4316
rect 5055 4276 5071 4280
rect 5075 4276 5077 4316
rect 5143 4276 5145 4316
rect 5149 4276 5151 4316
rect 4989 4236 5003 4244
rect 5194 4236 5196 4316
rect 5200 4236 5204 4316
rect 5208 4236 5210 4316
rect 5222 4276 5226 4316
rect 5230 4276 5232 4316
rect 5293 4236 5295 4316
rect 5299 4276 5301 4316
rect 5313 4276 5315 4316
rect 5319 4276 5329 4316
rect 5333 4276 5335 4316
rect 5347 4276 5349 4316
rect 5353 4276 5361 4316
rect 5365 4276 5367 4316
rect 5379 4276 5381 4316
rect 5385 4276 5387 4316
rect 5425 4276 5427 4316
rect 5431 4276 5435 4316
rect 5439 4296 5441 4316
rect 5453 4296 5455 4316
rect 5459 4296 5463 4316
rect 5467 4296 5471 4316
rect 5483 4296 5485 4316
rect 5439 4276 5450 4296
rect 5299 4236 5308 4276
rect 5476 4236 5485 4296
rect 5489 4236 5491 4316
rect 5529 4276 5531 4316
rect 5535 4276 5537 4316
rect 5549 4276 5551 4316
rect 5555 4276 5557 4316
rect 5609 4276 5611 4316
rect 5615 4276 5617 4316
rect 5674 4236 5676 4316
rect 5680 4236 5684 4316
rect 5688 4236 5690 4316
rect 5702 4276 5706 4316
rect 5710 4276 5712 4316
rect 5779 4236 5781 4316
rect 5785 4236 5787 4316
rect 5799 4276 5803 4316
rect 5807 4276 5811 4316
rect 5823 4276 5825 4316
rect 5829 4276 5831 4316
rect 5869 4276 5871 4316
rect 5875 4276 5877 4316
rect 5889 4276 5891 4316
rect 5895 4280 5897 4316
rect 5909 4280 5911 4316
rect 5895 4276 5911 4280
rect 5915 4276 5917 4316
rect 5983 4236 5985 4316
rect 5989 4236 5991 4316
rect 6034 4236 6036 4316
rect 6040 4236 6044 4316
rect 6048 4236 6050 4316
rect 6062 4276 6066 4316
rect 6070 4276 6072 4316
rect 6129 4276 6131 4316
rect 6135 4276 6139 4316
rect 6151 4236 6153 4316
rect 6157 4236 6159 4316
rect 6209 4276 6211 4316
rect 6215 4276 6217 4316
rect 6229 4276 6231 4316
rect 6235 4276 6237 4316
rect 6299 4236 6301 4316
rect 6305 4236 6307 4316
rect 6319 4276 6323 4316
rect 6327 4276 6331 4316
rect 6343 4276 6345 4316
rect 6349 4276 6351 4316
rect 6389 4276 6391 4316
rect 6395 4276 6397 4316
rect 6409 4276 6411 4316
rect 6415 4276 6417 4316
rect 6469 4276 6471 4316
rect 6475 4276 6477 4316
rect 6543 4236 6545 4316
rect 6549 4236 6551 4316
rect 6563 4236 6565 4316
rect 6569 4248 6571 4316
rect 6583 4248 6585 4316
rect 6569 4236 6585 4248
rect 6589 4244 6591 4316
rect 6629 4276 6631 4316
rect 6635 4276 6637 4316
rect 6649 4276 6651 4316
rect 6655 4280 6657 4316
rect 6669 4280 6671 4316
rect 6655 4276 6671 4280
rect 6675 4276 6677 4316
rect 6589 4236 6603 4244
rect 41 3864 43 3944
rect 47 3864 49 3944
rect 61 3864 65 3904
rect 69 3864 71 3904
rect 109 3864 111 3944
rect 115 3884 124 3944
rect 292 3904 301 3944
rect 150 3884 161 3904
rect 115 3864 117 3884
rect 129 3864 133 3884
rect 137 3864 141 3884
rect 145 3864 147 3884
rect 159 3864 161 3884
rect 165 3864 169 3904
rect 173 3864 175 3904
rect 213 3864 215 3904
rect 219 3864 221 3904
rect 233 3864 235 3904
rect 239 3864 247 3904
rect 251 3864 253 3904
rect 265 3864 267 3904
rect 271 3864 281 3904
rect 285 3864 287 3904
rect 299 3864 301 3904
rect 305 3864 307 3944
rect 349 3864 351 3904
rect 355 3864 357 3904
rect 369 3864 371 3904
rect 375 3864 377 3904
rect 443 3864 445 3944
rect 449 3864 451 3944
rect 463 3864 465 3944
rect 469 3932 485 3944
rect 469 3864 471 3932
rect 483 3864 485 3932
rect 489 3936 503 3944
rect 489 3864 491 3936
rect 543 3864 545 3904
rect 549 3864 551 3904
rect 563 3864 565 3904
rect 569 3864 571 3904
rect 623 3864 625 3904
rect 629 3864 631 3904
rect 643 3864 645 3904
rect 649 3864 651 3904
rect 701 3864 703 3944
rect 707 3864 709 3944
rect 721 3864 725 3904
rect 729 3864 731 3904
rect 769 3864 771 3944
rect 775 3884 784 3944
rect 952 3904 961 3944
rect 810 3884 821 3904
rect 775 3864 777 3884
rect 789 3864 793 3884
rect 797 3864 801 3884
rect 805 3864 807 3884
rect 819 3864 821 3884
rect 825 3864 829 3904
rect 833 3864 835 3904
rect 873 3864 875 3904
rect 879 3864 881 3904
rect 893 3864 895 3904
rect 899 3864 907 3904
rect 911 3864 913 3904
rect 925 3864 927 3904
rect 931 3864 941 3904
rect 945 3864 947 3904
rect 959 3864 961 3904
rect 965 3864 967 3944
rect 1023 3864 1025 3904
rect 1029 3864 1031 3904
rect 1043 3864 1045 3904
rect 1049 3864 1051 3904
rect 1089 3864 1091 3904
rect 1095 3864 1097 3904
rect 1109 3864 1111 3904
rect 1115 3864 1117 3904
rect 1169 3864 1171 3904
rect 1175 3864 1177 3904
rect 1189 3864 1191 3904
rect 1195 3864 1197 3904
rect 1263 3864 1265 3944
rect 1269 3864 1271 3944
rect 1283 3864 1285 3944
rect 1289 3932 1305 3944
rect 1289 3864 1291 3932
rect 1303 3864 1305 3932
rect 1309 3936 1323 3944
rect 1309 3864 1311 3936
rect 1349 3864 1351 3944
rect 1355 3884 1364 3944
rect 1532 3904 1541 3944
rect 1390 3884 1401 3904
rect 1355 3864 1357 3884
rect 1369 3864 1373 3884
rect 1377 3864 1381 3884
rect 1385 3864 1387 3884
rect 1399 3864 1401 3884
rect 1405 3864 1409 3904
rect 1413 3864 1415 3904
rect 1453 3864 1455 3904
rect 1459 3864 1461 3904
rect 1473 3864 1475 3904
rect 1479 3864 1487 3904
rect 1491 3864 1493 3904
rect 1505 3864 1507 3904
rect 1511 3864 1521 3904
rect 1525 3864 1527 3904
rect 1539 3864 1541 3904
rect 1545 3864 1547 3944
rect 1603 3864 1605 3904
rect 1609 3864 1611 3904
rect 1623 3864 1625 3904
rect 1629 3864 1631 3904
rect 1669 3864 1671 3904
rect 1675 3864 1679 3904
rect 1691 3864 1693 3944
rect 1697 3864 1699 3944
rect 1749 3864 1751 3904
rect 1755 3864 1757 3904
rect 1769 3864 1771 3904
rect 1775 3864 1777 3904
rect 1829 3864 1831 3944
rect 1835 3884 1844 3944
rect 2012 3904 2021 3944
rect 1870 3884 1881 3904
rect 1835 3864 1837 3884
rect 1849 3864 1853 3884
rect 1857 3864 1861 3884
rect 1865 3864 1867 3884
rect 1879 3864 1881 3884
rect 1885 3864 1889 3904
rect 1893 3864 1895 3904
rect 1933 3864 1935 3904
rect 1939 3864 1941 3904
rect 1953 3864 1955 3904
rect 1959 3864 1967 3904
rect 1971 3864 1973 3904
rect 1985 3864 1987 3904
rect 1991 3864 2001 3904
rect 2005 3864 2007 3904
rect 2019 3864 2021 3904
rect 2025 3864 2027 3944
rect 2069 3864 2071 3904
rect 2075 3864 2077 3904
rect 2089 3864 2091 3904
rect 2095 3864 2097 3904
rect 2168 3864 2170 3904
rect 2174 3864 2178 3904
rect 2190 3864 2192 3944
rect 2196 3864 2200 3944
rect 2204 3864 2206 3944
rect 2263 3864 2265 3904
rect 2269 3864 2271 3904
rect 2283 3864 2285 3904
rect 2289 3864 2291 3904
rect 2329 3864 2331 3904
rect 2335 3864 2337 3904
rect 2349 3864 2351 3904
rect 2355 3864 2357 3904
rect 2423 3864 2425 3904
rect 2429 3864 2431 3904
rect 2488 3864 2490 3904
rect 2494 3864 2498 3904
rect 2510 3864 2512 3944
rect 2516 3864 2520 3944
rect 2524 3864 2526 3944
rect 2569 3864 2571 3944
rect 2575 3864 2579 3944
rect 2583 3864 2585 3944
rect 2675 3864 2677 3944
rect 2681 3864 2685 3944
rect 2689 3864 2691 3944
rect 2729 3864 2731 3904
rect 2735 3864 2737 3904
rect 2803 3864 2805 3904
rect 2809 3864 2811 3904
rect 2863 3864 2865 3904
rect 2869 3864 2871 3904
rect 2883 3864 2885 3904
rect 2889 3864 2891 3904
rect 2929 3864 2931 3944
rect 2935 3864 2939 3944
rect 2943 3864 2945 3944
rect 3014 3864 3016 3944
rect 3020 3864 3024 3944
rect 3028 3864 3030 3944
rect 3042 3864 3046 3904
rect 3050 3864 3052 3904
rect 3109 3864 3111 3904
rect 3115 3864 3117 3904
rect 3169 3864 3171 3944
rect 3175 3864 3179 3944
rect 3183 3864 3185 3944
rect 3263 3864 3265 3904
rect 3269 3864 3271 3904
rect 3283 3864 3285 3904
rect 3289 3864 3291 3904
rect 3343 3864 3345 3904
rect 3349 3864 3351 3904
rect 3363 3864 3365 3904
rect 3369 3864 3371 3904
rect 3413 3864 3415 3944
rect 3419 3904 3428 3944
rect 3419 3864 3421 3904
rect 3433 3864 3435 3904
rect 3439 3864 3449 3904
rect 3453 3864 3455 3904
rect 3467 3864 3469 3904
rect 3473 3864 3481 3904
rect 3485 3864 3487 3904
rect 3499 3864 3501 3904
rect 3505 3864 3507 3904
rect 3545 3864 3547 3904
rect 3551 3864 3555 3904
rect 3559 3884 3570 3904
rect 3596 3884 3605 3944
rect 3559 3864 3561 3884
rect 3573 3864 3575 3884
rect 3579 3864 3583 3884
rect 3587 3864 3591 3884
rect 3603 3864 3605 3884
rect 3609 3864 3611 3944
rect 3663 3864 3665 3904
rect 3669 3864 3671 3904
rect 3713 3864 3715 3944
rect 3719 3904 3728 3944
rect 3719 3864 3721 3904
rect 3733 3864 3735 3904
rect 3739 3864 3749 3904
rect 3753 3864 3755 3904
rect 3767 3864 3769 3904
rect 3773 3864 3781 3904
rect 3785 3864 3787 3904
rect 3799 3864 3801 3904
rect 3805 3864 3807 3904
rect 3845 3864 3847 3904
rect 3851 3864 3855 3904
rect 3859 3884 3870 3904
rect 3896 3884 3905 3944
rect 3859 3864 3861 3884
rect 3873 3864 3875 3884
rect 3879 3864 3883 3884
rect 3887 3864 3891 3884
rect 3903 3864 3905 3884
rect 3909 3864 3911 3944
rect 3963 3864 3965 3904
rect 3969 3900 3985 3904
rect 3969 3864 3971 3900
rect 3983 3864 3985 3900
rect 3989 3864 3991 3904
rect 4003 3864 4005 3904
rect 4009 3864 4011 3904
rect 4049 3864 4051 3904
rect 4055 3864 4057 3904
rect 4069 3864 4071 3904
rect 4075 3864 4077 3904
rect 4148 3864 4150 3904
rect 4154 3864 4158 3904
rect 4170 3864 4172 3944
rect 4176 3864 4180 3944
rect 4184 3864 4186 3944
rect 4229 3864 4231 3944
rect 4235 3864 4239 3944
rect 4243 3864 4245 3944
rect 4323 3864 4325 3904
rect 4329 3864 4331 3904
rect 4383 3864 4385 3904
rect 4389 3864 4391 3904
rect 4403 3864 4405 3904
rect 4409 3864 4411 3904
rect 4468 3864 4470 3904
rect 4474 3864 4478 3904
rect 4490 3864 4492 3944
rect 4496 3864 4500 3944
rect 4504 3864 4506 3944
rect 4553 3864 4555 3944
rect 4559 3904 4568 3944
rect 4559 3864 4561 3904
rect 4573 3864 4575 3904
rect 4579 3864 4589 3904
rect 4593 3864 4595 3904
rect 4607 3864 4609 3904
rect 4613 3864 4621 3904
rect 4625 3864 4627 3904
rect 4639 3864 4641 3904
rect 4645 3864 4647 3904
rect 4685 3864 4687 3904
rect 4691 3864 4695 3904
rect 4699 3884 4710 3904
rect 4736 3884 4745 3944
rect 4699 3864 4701 3884
rect 4713 3864 4715 3884
rect 4719 3864 4723 3884
rect 4727 3864 4731 3884
rect 4743 3864 4745 3884
rect 4749 3864 4751 3944
rect 4803 3864 4805 3904
rect 4809 3864 4811 3904
rect 4823 3864 4825 3904
rect 4829 3864 4831 3904
rect 4888 3864 4890 3904
rect 4894 3864 4898 3904
rect 4910 3864 4912 3944
rect 4916 3864 4920 3944
rect 4924 3864 4926 3944
rect 4973 3864 4975 3944
rect 4979 3904 4988 3944
rect 4979 3864 4981 3904
rect 4993 3864 4995 3904
rect 4999 3864 5009 3904
rect 5013 3864 5015 3904
rect 5027 3864 5029 3904
rect 5033 3864 5041 3904
rect 5045 3864 5047 3904
rect 5059 3864 5061 3904
rect 5065 3864 5067 3904
rect 5105 3864 5107 3904
rect 5111 3864 5115 3904
rect 5119 3884 5130 3904
rect 5156 3884 5165 3944
rect 5119 3864 5121 3884
rect 5133 3864 5135 3884
rect 5139 3864 5143 3884
rect 5147 3864 5151 3884
rect 5163 3864 5165 3884
rect 5169 3864 5171 3944
rect 5223 3864 5225 3904
rect 5229 3864 5231 3904
rect 5243 3864 5245 3904
rect 5249 3864 5251 3904
rect 5308 3864 5310 3904
rect 5314 3864 5318 3904
rect 5330 3864 5332 3944
rect 5336 3864 5340 3944
rect 5344 3864 5346 3944
rect 5403 3864 5405 3904
rect 5409 3864 5411 3904
rect 5423 3864 5425 3904
rect 5429 3864 5431 3904
rect 5474 3864 5476 3944
rect 5480 3864 5484 3944
rect 5488 3864 5490 3944
rect 5502 3864 5506 3904
rect 5510 3864 5512 3904
rect 5583 3864 5585 3904
rect 5589 3864 5591 3904
rect 5633 3864 5635 3944
rect 5639 3904 5648 3944
rect 5639 3864 5641 3904
rect 5653 3864 5655 3904
rect 5659 3864 5669 3904
rect 5673 3864 5675 3904
rect 5687 3864 5689 3904
rect 5693 3864 5701 3904
rect 5705 3864 5707 3904
rect 5719 3864 5721 3904
rect 5725 3864 5727 3904
rect 5765 3864 5767 3904
rect 5771 3864 5775 3904
rect 5779 3884 5790 3904
rect 5816 3884 5825 3944
rect 5779 3864 5781 3884
rect 5793 3864 5795 3884
rect 5799 3864 5803 3884
rect 5807 3864 5811 3884
rect 5823 3864 5825 3884
rect 5829 3864 5831 3944
rect 5869 3864 5871 3904
rect 5875 3864 5877 3904
rect 5943 3864 5945 3904
rect 5949 3900 5965 3904
rect 5949 3864 5951 3900
rect 5963 3864 5965 3900
rect 5969 3864 5971 3904
rect 5983 3864 5985 3904
rect 5989 3864 5991 3904
rect 6029 3864 6031 3944
rect 6035 3884 6044 3944
rect 6212 3904 6221 3944
rect 6070 3884 6081 3904
rect 6035 3864 6037 3884
rect 6049 3864 6053 3884
rect 6057 3864 6061 3884
rect 6065 3864 6067 3884
rect 6079 3864 6081 3884
rect 6085 3864 6089 3904
rect 6093 3864 6095 3904
rect 6133 3864 6135 3904
rect 6139 3864 6141 3904
rect 6153 3864 6155 3904
rect 6159 3864 6167 3904
rect 6171 3864 6173 3904
rect 6185 3864 6187 3904
rect 6191 3864 6201 3904
rect 6205 3864 6207 3904
rect 6219 3864 6221 3904
rect 6225 3864 6227 3944
rect 6269 3864 6271 3944
rect 6275 3884 6284 3944
rect 6452 3904 6461 3944
rect 6310 3884 6321 3904
rect 6275 3864 6277 3884
rect 6289 3864 6293 3884
rect 6297 3864 6301 3884
rect 6305 3864 6307 3884
rect 6319 3864 6321 3884
rect 6325 3864 6329 3904
rect 6333 3864 6335 3904
rect 6373 3864 6375 3904
rect 6379 3864 6381 3904
rect 6393 3864 6395 3904
rect 6399 3864 6407 3904
rect 6411 3864 6413 3904
rect 6425 3864 6427 3904
rect 6431 3864 6441 3904
rect 6445 3864 6447 3904
rect 6459 3864 6461 3904
rect 6465 3864 6467 3944
rect 6509 3864 6511 3944
rect 6515 3884 6524 3944
rect 6692 3904 6701 3944
rect 6550 3884 6561 3904
rect 6515 3864 6517 3884
rect 6529 3864 6533 3884
rect 6537 3864 6541 3884
rect 6545 3864 6547 3884
rect 6559 3864 6561 3884
rect 6565 3864 6569 3904
rect 6573 3864 6575 3904
rect 6613 3864 6615 3904
rect 6619 3864 6621 3904
rect 6633 3864 6635 3904
rect 6639 3864 6647 3904
rect 6651 3864 6653 3904
rect 6665 3864 6667 3904
rect 6671 3864 6681 3904
rect 6685 3864 6687 3904
rect 6699 3864 6701 3904
rect 6705 3864 6707 3944
rect 41 3756 43 3836
rect 47 3756 49 3836
rect 61 3796 65 3836
rect 69 3796 71 3836
rect 121 3756 123 3836
rect 127 3756 129 3836
rect 141 3796 145 3836
rect 149 3796 151 3836
rect 203 3796 205 3836
rect 209 3796 211 3836
rect 223 3796 225 3836
rect 229 3796 231 3836
rect 269 3756 271 3836
rect 275 3816 277 3836
rect 289 3816 293 3836
rect 297 3816 301 3836
rect 305 3816 307 3836
rect 319 3816 321 3836
rect 275 3756 284 3816
rect 310 3796 321 3816
rect 325 3796 329 3836
rect 333 3796 335 3836
rect 373 3796 375 3836
rect 379 3796 381 3836
rect 393 3796 395 3836
rect 399 3796 407 3836
rect 411 3796 413 3836
rect 425 3796 427 3836
rect 431 3796 441 3836
rect 445 3796 447 3836
rect 459 3796 461 3836
rect 452 3756 461 3796
rect 465 3756 467 3836
rect 523 3756 525 3836
rect 529 3756 531 3836
rect 543 3756 545 3836
rect 549 3768 551 3836
rect 563 3768 565 3836
rect 549 3756 565 3768
rect 569 3764 571 3836
rect 623 3796 625 3836
rect 629 3796 631 3836
rect 643 3796 645 3836
rect 649 3796 651 3836
rect 689 3796 691 3836
rect 695 3796 697 3836
rect 709 3796 711 3836
rect 715 3796 717 3836
rect 783 3796 785 3836
rect 789 3796 791 3836
rect 803 3796 805 3836
rect 809 3796 811 3836
rect 569 3756 583 3764
rect 849 3756 851 3836
rect 855 3816 857 3836
rect 869 3816 873 3836
rect 877 3816 881 3836
rect 885 3816 887 3836
rect 899 3816 901 3836
rect 855 3756 864 3816
rect 890 3796 901 3816
rect 905 3796 909 3836
rect 913 3796 915 3836
rect 953 3796 955 3836
rect 959 3796 961 3836
rect 973 3796 975 3836
rect 979 3796 987 3836
rect 991 3796 993 3836
rect 1005 3796 1007 3836
rect 1011 3796 1021 3836
rect 1025 3796 1027 3836
rect 1039 3796 1041 3836
rect 1032 3756 1041 3796
rect 1045 3756 1047 3836
rect 1089 3764 1091 3836
rect 1077 3756 1091 3764
rect 1095 3768 1097 3836
rect 1109 3768 1111 3836
rect 1095 3756 1111 3768
rect 1115 3756 1117 3836
rect 1129 3756 1131 3836
rect 1135 3756 1137 3836
rect 1203 3796 1205 3836
rect 1209 3796 1211 3836
rect 1223 3796 1225 3836
rect 1229 3796 1231 3836
rect 1269 3796 1271 3836
rect 1275 3796 1279 3836
rect 1291 3756 1293 3836
rect 1297 3756 1299 3836
rect 1363 3756 1365 3836
rect 1369 3756 1371 3836
rect 1383 3756 1385 3836
rect 1389 3768 1391 3836
rect 1403 3768 1405 3836
rect 1389 3756 1405 3768
rect 1409 3764 1411 3836
rect 1463 3796 1465 3836
rect 1469 3796 1471 3836
rect 1483 3796 1485 3836
rect 1489 3796 1491 3836
rect 1529 3796 1531 3836
rect 1535 3796 1537 3836
rect 1549 3796 1551 3836
rect 1555 3796 1557 3836
rect 1409 3756 1423 3764
rect 1609 3756 1611 3836
rect 1615 3756 1619 3836
rect 1623 3756 1625 3836
rect 1689 3756 1691 3836
rect 1695 3816 1697 3836
rect 1709 3816 1713 3836
rect 1717 3816 1721 3836
rect 1725 3816 1727 3836
rect 1739 3816 1741 3836
rect 1695 3756 1704 3816
rect 1730 3796 1741 3816
rect 1745 3796 1749 3836
rect 1753 3796 1755 3836
rect 1793 3796 1795 3836
rect 1799 3796 1801 3836
rect 1813 3796 1815 3836
rect 1819 3796 1827 3836
rect 1831 3796 1833 3836
rect 1845 3796 1847 3836
rect 1851 3796 1861 3836
rect 1865 3796 1867 3836
rect 1879 3796 1881 3836
rect 1872 3756 1881 3796
rect 1885 3756 1887 3836
rect 1943 3796 1945 3836
rect 1949 3796 1951 3836
rect 1963 3796 1965 3836
rect 1969 3796 1971 3836
rect 2009 3756 2011 3836
rect 2015 3756 2019 3836
rect 2023 3756 2025 3836
rect 2089 3796 2091 3836
rect 2095 3796 2097 3836
rect 2154 3756 2156 3836
rect 2160 3756 2164 3836
rect 2168 3756 2170 3836
rect 2182 3796 2186 3836
rect 2190 3796 2192 3836
rect 2268 3796 2270 3836
rect 2274 3796 2278 3836
rect 2290 3756 2292 3836
rect 2296 3756 2300 3836
rect 2304 3756 2306 3836
rect 2363 3756 2365 3836
rect 2369 3756 2371 3836
rect 2383 3756 2385 3836
rect 2389 3768 2391 3836
rect 2403 3768 2405 3836
rect 2389 3756 2405 3768
rect 2409 3764 2411 3836
rect 2449 3796 2451 3836
rect 2455 3796 2457 3836
rect 2523 3796 2525 3836
rect 2529 3796 2531 3836
rect 2409 3756 2423 3764
rect 2574 3756 2576 3836
rect 2580 3756 2584 3836
rect 2588 3756 2590 3836
rect 2602 3796 2606 3836
rect 2610 3796 2612 3836
rect 2669 3796 2671 3836
rect 2675 3796 2677 3836
rect 2689 3796 2691 3836
rect 2695 3800 2697 3836
rect 2709 3800 2711 3836
rect 2695 3796 2711 3800
rect 2715 3796 2717 3836
rect 2783 3796 2785 3836
rect 2789 3796 2791 3836
rect 2843 3796 2845 3836
rect 2849 3796 2851 3836
rect 2863 3796 2865 3836
rect 2869 3796 2871 3836
rect 2914 3756 2916 3836
rect 2920 3756 2924 3836
rect 2928 3756 2930 3836
rect 2942 3796 2946 3836
rect 2950 3796 2952 3836
rect 3014 3756 3016 3836
rect 3020 3756 3024 3836
rect 3028 3756 3030 3836
rect 3042 3796 3046 3836
rect 3050 3796 3052 3836
rect 3109 3764 3111 3836
rect 3097 3756 3111 3764
rect 3115 3768 3117 3836
rect 3129 3768 3131 3836
rect 3115 3756 3131 3768
rect 3135 3756 3137 3836
rect 3149 3756 3151 3836
rect 3155 3756 3157 3836
rect 3223 3756 3225 3836
rect 3229 3824 3245 3836
rect 3229 3756 3231 3824
rect 3243 3756 3245 3824
rect 3249 3758 3251 3836
rect 3263 3758 3265 3836
rect 3249 3756 3265 3758
rect 3269 3770 3271 3836
rect 3283 3770 3285 3836
rect 3269 3756 3285 3770
rect 3289 3758 3291 3836
rect 3343 3796 3345 3836
rect 3349 3796 3351 3836
rect 3363 3796 3365 3836
rect 3369 3796 3371 3836
rect 3423 3796 3425 3836
rect 3429 3796 3431 3836
rect 3443 3796 3445 3836
rect 3449 3796 3451 3836
rect 3289 3756 3303 3758
rect 3493 3756 3495 3836
rect 3499 3796 3501 3836
rect 3513 3796 3515 3836
rect 3519 3796 3529 3836
rect 3533 3796 3535 3836
rect 3547 3796 3549 3836
rect 3553 3796 3561 3836
rect 3565 3796 3567 3836
rect 3579 3796 3581 3836
rect 3585 3796 3587 3836
rect 3625 3796 3627 3836
rect 3631 3796 3635 3836
rect 3639 3816 3641 3836
rect 3653 3816 3655 3836
rect 3659 3816 3663 3836
rect 3667 3816 3671 3836
rect 3683 3816 3685 3836
rect 3639 3796 3650 3816
rect 3499 3756 3508 3796
rect 3676 3756 3685 3816
rect 3689 3756 3691 3836
rect 3743 3796 3745 3836
rect 3749 3796 3751 3836
rect 3763 3796 3765 3836
rect 3769 3796 3771 3836
rect 3823 3756 3825 3836
rect 3829 3824 3845 3836
rect 3829 3756 3831 3824
rect 3843 3756 3845 3824
rect 3849 3758 3851 3836
rect 3863 3758 3865 3836
rect 3849 3756 3865 3758
rect 3869 3770 3871 3836
rect 3883 3770 3885 3836
rect 3869 3756 3885 3770
rect 3889 3758 3891 3836
rect 3929 3796 3931 3836
rect 3935 3796 3937 3836
rect 3989 3796 3991 3836
rect 3995 3796 3997 3836
rect 4009 3796 4011 3836
rect 4015 3796 4017 3836
rect 3889 3756 3903 3758
rect 4074 3756 4076 3836
rect 4080 3756 4084 3836
rect 4088 3756 4090 3836
rect 4102 3796 4106 3836
rect 4110 3796 4112 3836
rect 4173 3756 4175 3836
rect 4179 3796 4181 3836
rect 4193 3796 4195 3836
rect 4199 3796 4209 3836
rect 4213 3796 4215 3836
rect 4227 3796 4229 3836
rect 4233 3796 4241 3836
rect 4245 3796 4247 3836
rect 4259 3796 4261 3836
rect 4265 3796 4267 3836
rect 4305 3796 4307 3836
rect 4311 3796 4315 3836
rect 4319 3816 4321 3836
rect 4333 3816 4335 3836
rect 4339 3816 4343 3836
rect 4347 3816 4351 3836
rect 4363 3816 4365 3836
rect 4319 3796 4330 3816
rect 4179 3756 4188 3796
rect 4356 3756 4365 3816
rect 4369 3756 4371 3836
rect 4409 3796 4411 3836
rect 4415 3796 4417 3836
rect 4429 3796 4431 3836
rect 4435 3796 4437 3836
rect 4503 3796 4505 3836
rect 4509 3796 4511 3836
rect 4523 3796 4525 3836
rect 4529 3796 4531 3836
rect 4583 3756 4585 3836
rect 4589 3756 4591 3836
rect 4603 3756 4605 3836
rect 4609 3756 4611 3836
rect 4623 3756 4625 3836
rect 4629 3756 4631 3836
rect 4643 3756 4645 3836
rect 4649 3756 4651 3836
rect 4663 3756 4665 3836
rect 4669 3756 4671 3836
rect 4683 3756 4685 3836
rect 4689 3756 4691 3836
rect 4703 3756 4705 3836
rect 4709 3756 4711 3836
rect 4723 3756 4725 3836
rect 4729 3756 4731 3836
rect 4773 3756 4775 3836
rect 4779 3796 4781 3836
rect 4793 3796 4795 3836
rect 4799 3796 4809 3836
rect 4813 3796 4815 3836
rect 4827 3796 4829 3836
rect 4833 3796 4841 3836
rect 4845 3796 4847 3836
rect 4859 3796 4861 3836
rect 4865 3796 4867 3836
rect 4905 3796 4907 3836
rect 4911 3796 4915 3836
rect 4919 3816 4921 3836
rect 4933 3816 4935 3836
rect 4939 3816 4943 3836
rect 4947 3816 4951 3836
rect 4963 3816 4965 3836
rect 4919 3796 4930 3816
rect 4779 3756 4788 3796
rect 4956 3756 4965 3816
rect 4969 3756 4971 3836
rect 5014 3756 5016 3836
rect 5020 3756 5024 3836
rect 5028 3756 5030 3836
rect 5042 3796 5046 3836
rect 5050 3796 5052 3836
rect 5123 3796 5125 3836
rect 5129 3796 5131 3836
rect 5143 3796 5145 3836
rect 5149 3796 5151 3836
rect 5203 3796 5205 3836
rect 5209 3796 5211 3836
rect 5223 3796 5225 3836
rect 5229 3796 5231 3836
rect 5283 3796 5285 3836
rect 5289 3796 5291 3836
rect 5329 3756 5331 3836
rect 5335 3756 5337 3836
rect 5349 3756 5351 3836
rect 5355 3756 5357 3836
rect 5369 3756 5371 3836
rect 5375 3756 5377 3836
rect 5389 3756 5391 3836
rect 5395 3756 5397 3836
rect 5409 3756 5411 3836
rect 5415 3756 5417 3836
rect 5429 3756 5431 3836
rect 5435 3756 5437 3836
rect 5449 3756 5451 3836
rect 5455 3756 5457 3836
rect 5469 3756 5471 3836
rect 5475 3756 5477 3836
rect 5529 3756 5531 3836
rect 5535 3816 5537 3836
rect 5549 3816 5553 3836
rect 5557 3816 5561 3836
rect 5565 3816 5567 3836
rect 5579 3816 5581 3836
rect 5535 3756 5544 3816
rect 5570 3796 5581 3816
rect 5585 3796 5589 3836
rect 5593 3796 5595 3836
rect 5633 3796 5635 3836
rect 5639 3796 5641 3836
rect 5653 3796 5655 3836
rect 5659 3796 5667 3836
rect 5671 3796 5673 3836
rect 5685 3796 5687 3836
rect 5691 3796 5701 3836
rect 5705 3796 5707 3836
rect 5719 3796 5721 3836
rect 5712 3756 5721 3796
rect 5725 3756 5727 3836
rect 5783 3796 5785 3836
rect 5789 3796 5791 3836
rect 5829 3796 5831 3836
rect 5835 3796 5837 3836
rect 5849 3796 5851 3836
rect 5855 3796 5857 3836
rect 5909 3796 5911 3836
rect 5915 3796 5917 3836
rect 5929 3796 5931 3836
rect 5935 3796 5937 3836
rect 6003 3796 6005 3836
rect 6009 3796 6011 3836
rect 6049 3756 6051 3836
rect 6055 3756 6059 3836
rect 6063 3756 6065 3836
rect 6155 3756 6157 3836
rect 6161 3756 6165 3836
rect 6169 3756 6171 3836
rect 6209 3764 6211 3836
rect 6197 3756 6211 3764
rect 6215 3768 6217 3836
rect 6229 3768 6231 3836
rect 6215 3756 6231 3768
rect 6235 3756 6237 3836
rect 6249 3756 6251 3836
rect 6255 3756 6257 3836
rect 6309 3756 6311 3836
rect 6315 3816 6317 3836
rect 6329 3816 6333 3836
rect 6337 3816 6341 3836
rect 6345 3816 6347 3836
rect 6359 3816 6361 3836
rect 6315 3756 6324 3816
rect 6350 3796 6361 3816
rect 6365 3796 6369 3836
rect 6373 3796 6375 3836
rect 6413 3796 6415 3836
rect 6419 3796 6421 3836
rect 6433 3796 6435 3836
rect 6439 3796 6447 3836
rect 6451 3796 6453 3836
rect 6465 3796 6467 3836
rect 6471 3796 6481 3836
rect 6485 3796 6487 3836
rect 6499 3796 6501 3836
rect 6492 3756 6501 3796
rect 6505 3756 6507 3836
rect 6554 3756 6556 3836
rect 6560 3756 6564 3836
rect 6568 3756 6570 3836
rect 6582 3796 6586 3836
rect 6590 3796 6592 3836
rect 6649 3796 6651 3836
rect 6655 3796 6657 3836
rect 6669 3796 6671 3836
rect 6675 3796 6677 3836
rect 41 3384 43 3464
rect 47 3384 49 3464
rect 61 3384 65 3424
rect 69 3384 71 3424
rect 109 3384 111 3464
rect 115 3404 124 3464
rect 292 3424 301 3464
rect 150 3404 161 3424
rect 115 3384 117 3404
rect 129 3384 133 3404
rect 137 3384 141 3404
rect 145 3384 147 3404
rect 159 3384 161 3404
rect 165 3384 169 3424
rect 173 3384 175 3424
rect 213 3384 215 3424
rect 219 3384 221 3424
rect 233 3384 235 3424
rect 239 3384 247 3424
rect 251 3384 253 3424
rect 265 3384 267 3424
rect 271 3384 281 3424
rect 285 3384 287 3424
rect 299 3384 301 3424
rect 305 3384 307 3464
rect 349 3384 351 3424
rect 355 3384 357 3424
rect 369 3384 371 3424
rect 375 3384 377 3424
rect 429 3384 431 3424
rect 435 3384 439 3424
rect 451 3384 453 3464
rect 457 3384 459 3464
rect 523 3384 525 3464
rect 529 3384 531 3464
rect 543 3384 545 3464
rect 549 3452 565 3464
rect 549 3384 551 3452
rect 563 3384 565 3452
rect 569 3456 583 3464
rect 569 3384 571 3456
rect 623 3384 625 3424
rect 629 3384 631 3424
rect 643 3384 645 3424
rect 649 3384 651 3424
rect 701 3384 703 3464
rect 707 3384 709 3464
rect 721 3384 725 3424
rect 729 3384 731 3424
rect 769 3384 771 3424
rect 775 3384 779 3424
rect 791 3384 793 3464
rect 797 3384 799 3464
rect 849 3384 851 3424
rect 855 3384 857 3424
rect 869 3384 871 3424
rect 875 3384 877 3424
rect 941 3384 943 3464
rect 947 3384 949 3464
rect 961 3384 965 3424
rect 969 3384 971 3424
rect 1023 3384 1025 3424
rect 1029 3384 1031 3424
rect 1081 3384 1083 3464
rect 1087 3384 1089 3464
rect 1101 3384 1105 3424
rect 1109 3384 1111 3424
rect 1161 3384 1163 3464
rect 1167 3384 1169 3464
rect 1181 3384 1185 3424
rect 1189 3384 1191 3424
rect 1229 3384 1231 3464
rect 1235 3404 1244 3464
rect 1412 3424 1421 3464
rect 1270 3404 1281 3424
rect 1235 3384 1237 3404
rect 1249 3384 1253 3404
rect 1257 3384 1261 3404
rect 1265 3384 1267 3404
rect 1279 3384 1281 3404
rect 1285 3384 1289 3424
rect 1293 3384 1295 3424
rect 1333 3384 1335 3424
rect 1339 3384 1341 3424
rect 1353 3384 1355 3424
rect 1359 3384 1367 3424
rect 1371 3384 1373 3424
rect 1385 3384 1387 3424
rect 1391 3384 1401 3424
rect 1405 3384 1407 3424
rect 1419 3384 1421 3424
rect 1425 3384 1427 3464
rect 1495 3384 1497 3464
rect 1501 3384 1505 3464
rect 1509 3384 1511 3464
rect 1549 3384 1551 3464
rect 1555 3404 1564 3464
rect 1732 3424 1741 3464
rect 1590 3404 1601 3424
rect 1555 3384 1557 3404
rect 1569 3384 1573 3404
rect 1577 3384 1581 3404
rect 1585 3384 1587 3404
rect 1599 3384 1601 3404
rect 1605 3384 1609 3424
rect 1613 3384 1615 3424
rect 1653 3384 1655 3424
rect 1659 3384 1661 3424
rect 1673 3384 1675 3424
rect 1679 3384 1687 3424
rect 1691 3384 1693 3424
rect 1705 3384 1707 3424
rect 1711 3384 1721 3424
rect 1725 3384 1727 3424
rect 1739 3384 1741 3424
rect 1745 3384 1747 3464
rect 1799 3384 1801 3464
rect 1805 3384 1807 3464
rect 1819 3384 1823 3424
rect 1827 3384 1831 3424
rect 1843 3384 1845 3424
rect 1849 3384 1851 3424
rect 1903 3384 1905 3424
rect 1909 3384 1911 3424
rect 1968 3384 1970 3424
rect 1974 3384 1978 3424
rect 1990 3384 1992 3464
rect 1996 3384 2000 3464
rect 2004 3384 2006 3464
rect 2049 3384 2051 3464
rect 2055 3384 2059 3464
rect 2063 3384 2065 3464
rect 2143 3384 2145 3424
rect 2149 3384 2151 3424
rect 2199 3384 2201 3464
rect 2205 3384 2207 3464
rect 2219 3384 2223 3424
rect 2227 3384 2231 3424
rect 2243 3384 2245 3424
rect 2249 3384 2251 3424
rect 2315 3384 2317 3464
rect 2321 3384 2325 3464
rect 2329 3384 2331 3464
rect 2369 3384 2371 3464
rect 2375 3404 2384 3464
rect 2552 3424 2561 3464
rect 2410 3404 2421 3424
rect 2375 3384 2377 3404
rect 2389 3384 2393 3404
rect 2397 3384 2401 3404
rect 2405 3384 2407 3404
rect 2419 3384 2421 3404
rect 2425 3384 2429 3424
rect 2433 3384 2435 3424
rect 2473 3384 2475 3424
rect 2479 3384 2481 3424
rect 2493 3384 2495 3424
rect 2499 3384 2507 3424
rect 2511 3384 2513 3424
rect 2525 3384 2527 3424
rect 2531 3384 2541 3424
rect 2545 3384 2547 3424
rect 2559 3384 2561 3424
rect 2565 3384 2567 3464
rect 2609 3384 2611 3464
rect 2615 3384 2619 3464
rect 2623 3384 2625 3464
rect 2694 3384 2696 3464
rect 2700 3384 2704 3464
rect 2708 3384 2710 3464
rect 2722 3384 2726 3424
rect 2730 3384 2732 3424
rect 2803 3384 2805 3424
rect 2809 3384 2811 3424
rect 2863 3384 2865 3424
rect 2869 3384 2871 3424
rect 2883 3384 2885 3424
rect 2889 3384 2891 3424
rect 2934 3384 2936 3464
rect 2940 3384 2944 3464
rect 2948 3384 2950 3464
rect 3017 3456 3031 3464
rect 2962 3384 2966 3424
rect 2970 3384 2972 3424
rect 3029 3384 3031 3456
rect 3035 3452 3051 3464
rect 3035 3384 3037 3452
rect 3049 3384 3051 3452
rect 3055 3384 3057 3464
rect 3069 3384 3071 3464
rect 3075 3384 3077 3464
rect 3129 3384 3131 3464
rect 3135 3384 3137 3464
rect 3203 3384 3205 3464
rect 3209 3396 3211 3464
rect 3223 3396 3225 3464
rect 3209 3384 3225 3396
rect 3229 3462 3245 3464
rect 3229 3384 3231 3462
rect 3243 3384 3245 3462
rect 3249 3450 3265 3464
rect 3249 3384 3251 3450
rect 3263 3384 3265 3450
rect 3269 3462 3283 3464
rect 3269 3384 3271 3462
rect 3323 3384 3325 3424
rect 3329 3384 3331 3424
rect 3369 3384 3371 3464
rect 3375 3404 3384 3464
rect 3552 3424 3561 3464
rect 3410 3404 3421 3424
rect 3375 3384 3377 3404
rect 3389 3384 3393 3404
rect 3397 3384 3401 3404
rect 3405 3384 3407 3404
rect 3419 3384 3421 3404
rect 3425 3384 3429 3424
rect 3433 3384 3435 3424
rect 3473 3384 3475 3424
rect 3479 3384 3481 3424
rect 3493 3384 3495 3424
rect 3499 3384 3507 3424
rect 3511 3384 3513 3424
rect 3525 3384 3527 3424
rect 3531 3384 3541 3424
rect 3545 3384 3547 3424
rect 3559 3384 3561 3424
rect 3565 3384 3567 3464
rect 3623 3384 3625 3464
rect 3629 3396 3631 3464
rect 3643 3396 3645 3464
rect 3629 3384 3645 3396
rect 3649 3462 3665 3464
rect 3649 3384 3651 3462
rect 3663 3384 3665 3462
rect 3669 3450 3685 3464
rect 3669 3384 3671 3450
rect 3683 3384 3685 3450
rect 3689 3462 3703 3464
rect 3689 3384 3691 3462
rect 3729 3384 3731 3464
rect 3735 3404 3744 3464
rect 3912 3424 3921 3464
rect 3770 3404 3781 3424
rect 3735 3384 3737 3404
rect 3749 3384 3753 3404
rect 3757 3384 3761 3404
rect 3765 3384 3767 3404
rect 3779 3384 3781 3404
rect 3785 3384 3789 3424
rect 3793 3384 3795 3424
rect 3833 3384 3835 3424
rect 3839 3384 3841 3424
rect 3853 3384 3855 3424
rect 3859 3384 3867 3424
rect 3871 3384 3873 3424
rect 3885 3384 3887 3424
rect 3891 3384 3901 3424
rect 3905 3384 3907 3424
rect 3919 3384 3921 3424
rect 3925 3384 3927 3464
rect 3983 3384 3985 3424
rect 3989 3384 3991 3424
rect 4029 3384 4031 3464
rect 4035 3404 4044 3464
rect 4212 3424 4221 3464
rect 4070 3404 4081 3424
rect 4035 3384 4037 3404
rect 4049 3384 4053 3404
rect 4057 3384 4061 3404
rect 4065 3384 4067 3404
rect 4079 3384 4081 3404
rect 4085 3384 4089 3424
rect 4093 3384 4095 3424
rect 4133 3384 4135 3424
rect 4139 3384 4141 3424
rect 4153 3384 4155 3424
rect 4159 3384 4167 3424
rect 4171 3384 4173 3424
rect 4185 3384 4187 3424
rect 4191 3384 4201 3424
rect 4205 3384 4207 3424
rect 4219 3384 4221 3424
rect 4225 3384 4227 3464
rect 4283 3384 4285 3424
rect 4289 3384 4291 3424
rect 4343 3384 4345 3424
rect 4349 3384 4351 3424
rect 4389 3384 4391 3424
rect 4395 3384 4397 3424
rect 4409 3384 4411 3424
rect 4415 3384 4417 3424
rect 4473 3384 4475 3464
rect 4479 3424 4488 3464
rect 4479 3384 4481 3424
rect 4493 3384 4495 3424
rect 4499 3384 4509 3424
rect 4513 3384 4515 3424
rect 4527 3384 4529 3424
rect 4533 3384 4541 3424
rect 4545 3384 4547 3424
rect 4559 3384 4561 3424
rect 4565 3384 4567 3424
rect 4605 3384 4607 3424
rect 4611 3384 4615 3424
rect 4619 3404 4630 3424
rect 4656 3404 4665 3464
rect 4619 3384 4621 3404
rect 4633 3384 4635 3404
rect 4639 3384 4643 3404
rect 4647 3384 4651 3404
rect 4663 3384 4665 3404
rect 4669 3384 4671 3464
rect 4723 3384 4725 3424
rect 4729 3384 4731 3424
rect 4769 3384 4771 3464
rect 4775 3404 4784 3464
rect 4952 3424 4961 3464
rect 4810 3404 4821 3424
rect 4775 3384 4777 3404
rect 4789 3384 4793 3404
rect 4797 3384 4801 3404
rect 4805 3384 4807 3404
rect 4819 3384 4821 3404
rect 4825 3384 4829 3424
rect 4833 3384 4835 3424
rect 4873 3384 4875 3424
rect 4879 3384 4881 3424
rect 4893 3384 4895 3424
rect 4899 3384 4907 3424
rect 4911 3384 4913 3424
rect 4925 3384 4927 3424
rect 4931 3384 4941 3424
rect 4945 3384 4947 3424
rect 4959 3384 4961 3424
rect 4965 3384 4967 3464
rect 5023 3384 5025 3464
rect 5029 3396 5031 3464
rect 5043 3396 5045 3464
rect 5029 3384 5045 3396
rect 5049 3462 5065 3464
rect 5049 3384 5051 3462
rect 5063 3384 5065 3462
rect 5069 3450 5085 3464
rect 5069 3384 5071 3450
rect 5083 3384 5085 3450
rect 5089 3462 5103 3464
rect 5089 3384 5091 3462
rect 5143 3384 5145 3424
rect 5149 3384 5151 3424
rect 5189 3384 5191 3464
rect 5195 3404 5204 3464
rect 5372 3424 5381 3464
rect 5230 3404 5241 3424
rect 5195 3384 5197 3404
rect 5209 3384 5213 3404
rect 5217 3384 5221 3404
rect 5225 3384 5227 3404
rect 5239 3384 5241 3404
rect 5245 3384 5249 3424
rect 5253 3384 5255 3424
rect 5293 3384 5295 3424
rect 5299 3384 5301 3424
rect 5313 3384 5315 3424
rect 5319 3384 5327 3424
rect 5331 3384 5333 3424
rect 5345 3384 5347 3424
rect 5351 3384 5361 3424
rect 5365 3384 5367 3424
rect 5379 3384 5381 3424
rect 5385 3384 5387 3464
rect 5429 3384 5431 3464
rect 5435 3404 5444 3464
rect 5612 3424 5621 3464
rect 5470 3404 5481 3424
rect 5435 3384 5437 3404
rect 5449 3384 5453 3404
rect 5457 3384 5461 3404
rect 5465 3384 5467 3404
rect 5479 3384 5481 3404
rect 5485 3384 5489 3424
rect 5493 3384 5495 3424
rect 5533 3384 5535 3424
rect 5539 3384 5541 3424
rect 5553 3384 5555 3424
rect 5559 3384 5567 3424
rect 5571 3384 5573 3424
rect 5585 3384 5587 3424
rect 5591 3384 5601 3424
rect 5605 3384 5607 3424
rect 5619 3384 5621 3424
rect 5625 3384 5627 3464
rect 5674 3384 5676 3464
rect 5680 3384 5684 3464
rect 5688 3384 5690 3464
rect 5702 3384 5706 3424
rect 5710 3384 5712 3424
rect 5774 3384 5776 3464
rect 5780 3384 5784 3464
rect 5788 3384 5790 3464
rect 5802 3384 5806 3424
rect 5810 3384 5812 3424
rect 5883 3384 5885 3424
rect 5889 3384 5891 3424
rect 5943 3384 5945 3464
rect 5949 3396 5951 3464
rect 5963 3396 5965 3464
rect 5949 3384 5965 3396
rect 5969 3462 5985 3464
rect 5969 3384 5971 3462
rect 5983 3384 5985 3462
rect 5989 3450 6005 3464
rect 5989 3384 5991 3450
rect 6003 3384 6005 3450
rect 6009 3462 6023 3464
rect 6009 3384 6011 3462
rect 6049 3384 6051 3424
rect 6055 3384 6057 3424
rect 6069 3384 6071 3424
rect 6075 3384 6077 3424
rect 6143 3384 6145 3424
rect 6149 3384 6151 3424
rect 6189 3384 6191 3444
rect 6195 3384 6197 3444
rect 6209 3384 6211 3444
rect 6215 3384 6217 3444
rect 6229 3384 6231 3444
rect 6235 3396 6237 3444
rect 6249 3396 6251 3444
rect 6235 3384 6251 3396
rect 6255 3442 6269 3444
rect 6255 3384 6257 3442
rect 6293 3392 6295 3452
rect 6299 3448 6315 3452
rect 6299 3396 6301 3448
rect 6313 3396 6315 3448
rect 6299 3392 6315 3396
rect 6319 3392 6321 3452
rect 6383 3384 6385 3424
rect 6389 3384 6391 3424
rect 6429 3384 6431 3464
rect 6435 3404 6444 3464
rect 6612 3424 6621 3464
rect 6470 3404 6481 3424
rect 6435 3384 6437 3404
rect 6449 3384 6453 3404
rect 6457 3384 6461 3404
rect 6465 3384 6467 3404
rect 6479 3384 6481 3404
rect 6485 3384 6489 3424
rect 6493 3384 6495 3424
rect 6533 3384 6535 3424
rect 6539 3384 6541 3424
rect 6553 3384 6555 3424
rect 6559 3384 6567 3424
rect 6571 3384 6573 3424
rect 6585 3384 6587 3424
rect 6591 3384 6601 3424
rect 6605 3384 6607 3424
rect 6619 3384 6621 3424
rect 6625 3384 6627 3464
rect 41 3276 43 3356
rect 47 3276 49 3356
rect 61 3316 65 3356
rect 69 3316 71 3356
rect 109 3276 111 3356
rect 115 3336 117 3356
rect 129 3336 133 3356
rect 137 3336 141 3356
rect 145 3336 147 3356
rect 159 3336 161 3356
rect 115 3276 124 3336
rect 150 3316 161 3336
rect 165 3316 169 3356
rect 173 3316 175 3356
rect 213 3316 215 3356
rect 219 3316 221 3356
rect 233 3316 235 3356
rect 239 3316 247 3356
rect 251 3316 253 3356
rect 265 3316 267 3356
rect 271 3316 281 3356
rect 285 3316 287 3356
rect 299 3316 301 3356
rect 292 3276 301 3316
rect 305 3276 307 3356
rect 349 3316 351 3356
rect 355 3316 357 3356
rect 369 3316 371 3356
rect 375 3316 377 3356
rect 443 3276 445 3356
rect 449 3276 451 3356
rect 463 3276 465 3356
rect 469 3288 471 3356
rect 483 3288 485 3356
rect 469 3276 485 3288
rect 489 3284 491 3356
rect 543 3316 545 3356
rect 549 3316 551 3356
rect 563 3316 565 3356
rect 569 3316 571 3356
rect 609 3316 611 3356
rect 615 3316 617 3356
rect 669 3316 671 3356
rect 675 3316 677 3356
rect 689 3316 691 3356
rect 695 3320 697 3356
rect 709 3320 711 3356
rect 695 3316 711 3320
rect 715 3316 717 3356
rect 769 3316 771 3356
rect 775 3316 777 3356
rect 789 3316 791 3356
rect 795 3316 797 3356
rect 868 3316 870 3356
rect 874 3316 878 3356
rect 489 3276 503 3284
rect 890 3276 892 3356
rect 896 3276 900 3356
rect 904 3276 906 3356
rect 949 3316 951 3356
rect 955 3316 957 3356
rect 1009 3276 1011 3356
rect 1015 3276 1019 3356
rect 1023 3276 1025 3356
rect 1094 3276 1096 3356
rect 1100 3276 1104 3356
rect 1108 3276 1110 3356
rect 1122 3316 1126 3356
rect 1130 3316 1132 3356
rect 1194 3276 1196 3356
rect 1200 3276 1204 3356
rect 1208 3276 1210 3356
rect 1222 3316 1226 3356
rect 1230 3316 1232 3356
rect 1289 3316 1291 3356
rect 1295 3316 1297 3356
rect 1309 3316 1311 3356
rect 1315 3316 1317 3356
rect 1369 3276 1371 3356
rect 1375 3336 1377 3356
rect 1389 3336 1393 3356
rect 1397 3336 1401 3356
rect 1405 3336 1407 3356
rect 1419 3336 1421 3356
rect 1375 3276 1384 3336
rect 1410 3316 1421 3336
rect 1425 3316 1429 3356
rect 1433 3316 1435 3356
rect 1473 3316 1475 3356
rect 1479 3316 1481 3356
rect 1493 3316 1495 3356
rect 1499 3316 1507 3356
rect 1511 3316 1513 3356
rect 1525 3316 1527 3356
rect 1531 3316 1541 3356
rect 1545 3316 1547 3356
rect 1559 3316 1561 3356
rect 1552 3276 1561 3316
rect 1565 3276 1567 3356
rect 1619 3276 1621 3356
rect 1625 3276 1627 3356
rect 1639 3316 1643 3356
rect 1647 3316 1651 3356
rect 1663 3316 1665 3356
rect 1669 3316 1671 3356
rect 1723 3276 1725 3356
rect 1729 3276 1731 3356
rect 1743 3276 1745 3356
rect 1749 3288 1751 3356
rect 1763 3288 1765 3356
rect 1749 3276 1765 3288
rect 1769 3284 1771 3356
rect 1823 3316 1825 3356
rect 1829 3320 1831 3356
rect 1843 3320 1845 3356
rect 1829 3316 1845 3320
rect 1849 3316 1851 3356
rect 1863 3316 1865 3356
rect 1869 3316 1871 3356
rect 1769 3276 1783 3284
rect 1909 3284 1911 3356
rect 1897 3276 1911 3284
rect 1915 3288 1917 3356
rect 1929 3288 1931 3356
rect 1915 3276 1931 3288
rect 1935 3276 1937 3356
rect 1949 3276 1951 3356
rect 1955 3276 1957 3356
rect 2013 3276 2015 3356
rect 2019 3316 2021 3356
rect 2033 3316 2035 3356
rect 2039 3316 2049 3356
rect 2053 3316 2055 3356
rect 2067 3316 2069 3356
rect 2073 3316 2081 3356
rect 2085 3316 2087 3356
rect 2099 3316 2101 3356
rect 2105 3316 2107 3356
rect 2145 3316 2147 3356
rect 2151 3316 2155 3356
rect 2159 3336 2161 3356
rect 2173 3336 2175 3356
rect 2179 3336 2183 3356
rect 2187 3336 2191 3356
rect 2203 3336 2205 3356
rect 2159 3316 2170 3336
rect 2019 3276 2028 3316
rect 2196 3276 2205 3336
rect 2209 3276 2211 3356
rect 2249 3316 2251 3356
rect 2255 3316 2257 3356
rect 2269 3316 2271 3356
rect 2275 3316 2277 3356
rect 2329 3276 2331 3356
rect 2335 3276 2339 3356
rect 2343 3276 2345 3356
rect 2435 3276 2437 3356
rect 2441 3276 2445 3356
rect 2449 3276 2451 3356
rect 2508 3316 2510 3356
rect 2514 3316 2518 3356
rect 2530 3276 2532 3356
rect 2536 3276 2540 3356
rect 2544 3276 2546 3356
rect 2589 3316 2591 3356
rect 2595 3316 2597 3356
rect 2653 3276 2655 3356
rect 2659 3316 2661 3356
rect 2673 3316 2675 3356
rect 2679 3316 2689 3356
rect 2693 3316 2695 3356
rect 2707 3316 2709 3356
rect 2713 3316 2721 3356
rect 2725 3316 2727 3356
rect 2739 3316 2741 3356
rect 2745 3316 2747 3356
rect 2785 3316 2787 3356
rect 2791 3316 2795 3356
rect 2799 3336 2801 3356
rect 2813 3336 2815 3356
rect 2819 3336 2823 3356
rect 2827 3336 2831 3356
rect 2843 3336 2845 3356
rect 2799 3316 2810 3336
rect 2659 3276 2668 3316
rect 2836 3276 2845 3336
rect 2849 3276 2851 3356
rect 2889 3316 2891 3356
rect 2895 3316 2897 3356
rect 2909 3316 2911 3356
rect 2915 3316 2917 3356
rect 2983 3316 2985 3356
rect 2989 3316 2991 3356
rect 3003 3316 3005 3356
rect 3009 3316 3011 3356
rect 3068 3316 3070 3356
rect 3074 3316 3078 3356
rect 3090 3276 3092 3356
rect 3096 3276 3100 3356
rect 3104 3276 3106 3356
rect 3163 3316 3165 3356
rect 3169 3316 3171 3356
rect 3183 3316 3185 3356
rect 3189 3316 3191 3356
rect 3243 3316 3245 3356
rect 3249 3316 3251 3356
rect 3308 3316 3310 3356
rect 3314 3316 3318 3356
rect 3330 3276 3332 3356
rect 3336 3276 3340 3356
rect 3344 3276 3346 3356
rect 3389 3316 3391 3356
rect 3395 3316 3397 3356
rect 3475 3276 3477 3356
rect 3481 3276 3485 3356
rect 3489 3276 3491 3356
rect 3543 3276 3545 3356
rect 3549 3276 3551 3356
rect 3563 3276 3565 3356
rect 3569 3288 3571 3356
rect 3583 3288 3585 3356
rect 3569 3276 3585 3288
rect 3589 3284 3591 3356
rect 3589 3276 3603 3284
rect 3655 3276 3657 3356
rect 3661 3276 3665 3356
rect 3669 3276 3671 3356
rect 3709 3276 3711 3356
rect 3715 3336 3717 3356
rect 3729 3336 3733 3356
rect 3737 3336 3741 3356
rect 3745 3336 3747 3356
rect 3759 3336 3761 3356
rect 3715 3276 3724 3336
rect 3750 3316 3761 3336
rect 3765 3316 3769 3356
rect 3773 3316 3775 3356
rect 3813 3316 3815 3356
rect 3819 3316 3821 3356
rect 3833 3316 3835 3356
rect 3839 3316 3847 3356
rect 3851 3316 3853 3356
rect 3865 3316 3867 3356
rect 3871 3316 3881 3356
rect 3885 3316 3887 3356
rect 3899 3316 3901 3356
rect 3892 3276 3901 3316
rect 3905 3276 3907 3356
rect 3949 3278 3951 3356
rect 3937 3276 3951 3278
rect 3955 3290 3957 3356
rect 3969 3290 3971 3356
rect 3955 3276 3971 3290
rect 3975 3278 3977 3356
rect 3989 3278 3991 3356
rect 3975 3276 3991 3278
rect 3995 3344 4011 3356
rect 3995 3276 3997 3344
rect 4009 3276 4011 3344
rect 4015 3276 4017 3356
rect 4083 3276 4085 3356
rect 4089 3344 4105 3356
rect 4089 3276 4091 3344
rect 4103 3276 4105 3344
rect 4109 3278 4111 3356
rect 4123 3278 4125 3356
rect 4109 3276 4125 3278
rect 4129 3290 4131 3356
rect 4143 3290 4145 3356
rect 4129 3276 4145 3290
rect 4149 3278 4151 3356
rect 4149 3276 4163 3278
rect 4193 3276 4195 3356
rect 4199 3316 4201 3356
rect 4213 3316 4215 3356
rect 4219 3316 4229 3356
rect 4233 3316 4235 3356
rect 4247 3316 4249 3356
rect 4253 3316 4261 3356
rect 4265 3316 4267 3356
rect 4279 3316 4281 3356
rect 4285 3316 4287 3356
rect 4325 3316 4327 3356
rect 4331 3316 4335 3356
rect 4339 3336 4341 3356
rect 4353 3336 4355 3356
rect 4359 3336 4363 3356
rect 4367 3336 4371 3356
rect 4383 3336 4385 3356
rect 4339 3316 4350 3336
rect 4199 3276 4208 3316
rect 4376 3276 4385 3336
rect 4389 3276 4391 3356
rect 4429 3276 4431 3356
rect 4435 3276 4439 3356
rect 4443 3276 4445 3356
rect 4509 3278 4511 3356
rect 4497 3276 4511 3278
rect 4515 3290 4517 3356
rect 4529 3290 4531 3356
rect 4515 3276 4531 3290
rect 4535 3278 4537 3356
rect 4549 3278 4551 3356
rect 4535 3276 4551 3278
rect 4555 3344 4571 3356
rect 4555 3276 4557 3344
rect 4569 3276 4571 3344
rect 4575 3276 4577 3356
rect 4629 3276 4631 3356
rect 4635 3276 4639 3356
rect 4643 3276 4645 3356
rect 4709 3276 4711 3356
rect 4715 3276 4719 3356
rect 4723 3276 4725 3356
rect 4789 3316 4791 3356
rect 4795 3316 4797 3356
rect 4849 3278 4851 3356
rect 4837 3276 4851 3278
rect 4855 3290 4857 3356
rect 4869 3290 4871 3356
rect 4855 3276 4871 3290
rect 4875 3278 4877 3356
rect 4889 3278 4891 3356
rect 4875 3276 4891 3278
rect 4895 3344 4911 3356
rect 4895 3276 4897 3344
rect 4909 3276 4911 3344
rect 4915 3276 4917 3356
rect 4969 3284 4971 3356
rect 4957 3276 4971 3284
rect 4975 3288 4977 3356
rect 4989 3288 4991 3356
rect 4975 3276 4991 3288
rect 4995 3276 4997 3356
rect 5009 3276 5011 3356
rect 5015 3276 5017 3356
rect 5069 3276 5071 3356
rect 5075 3336 5077 3356
rect 5089 3336 5093 3356
rect 5097 3336 5101 3356
rect 5105 3336 5107 3356
rect 5119 3336 5121 3356
rect 5075 3276 5084 3336
rect 5110 3316 5121 3336
rect 5125 3316 5129 3356
rect 5133 3316 5135 3356
rect 5173 3316 5175 3356
rect 5179 3316 5181 3356
rect 5193 3316 5195 3356
rect 5199 3316 5207 3356
rect 5211 3316 5213 3356
rect 5225 3316 5227 3356
rect 5231 3316 5241 3356
rect 5245 3316 5247 3356
rect 5259 3316 5261 3356
rect 5252 3276 5261 3316
rect 5265 3276 5267 3356
rect 5323 3316 5325 3356
rect 5329 3316 5331 3356
rect 5412 3348 5421 3356
rect 5369 3308 5371 3348
rect 5375 3308 5377 3348
rect 5389 3308 5391 3348
rect 5381 3268 5391 3308
rect 5395 3268 5401 3348
rect 5405 3284 5407 3348
rect 5419 3284 5421 3348
rect 5405 3276 5421 3284
rect 5425 3276 5431 3356
rect 5435 3276 5437 3356
rect 5503 3316 5505 3356
rect 5509 3316 5511 3356
rect 5405 3268 5413 3276
rect 5553 3276 5555 3356
rect 5559 3316 5561 3356
rect 5573 3316 5575 3356
rect 5579 3316 5589 3356
rect 5593 3316 5595 3356
rect 5607 3316 5609 3356
rect 5613 3316 5621 3356
rect 5625 3316 5627 3356
rect 5639 3316 5641 3356
rect 5645 3316 5647 3356
rect 5685 3316 5687 3356
rect 5691 3316 5695 3356
rect 5699 3336 5701 3356
rect 5713 3336 5715 3356
rect 5719 3336 5723 3356
rect 5727 3336 5731 3356
rect 5743 3336 5745 3356
rect 5699 3316 5710 3336
rect 5559 3276 5568 3316
rect 5736 3276 5745 3336
rect 5749 3276 5751 3356
rect 5808 3316 5810 3356
rect 5814 3316 5818 3356
rect 5830 3276 5832 3356
rect 5836 3276 5840 3356
rect 5844 3276 5846 3356
rect 5903 3316 5905 3356
rect 5909 3316 5911 3356
rect 5963 3276 5965 3356
rect 5969 3276 5971 3356
rect 5983 3276 5985 3356
rect 5989 3288 5991 3356
rect 6003 3288 6005 3356
rect 5989 3276 6005 3288
rect 6009 3284 6011 3356
rect 6009 3276 6023 3284
rect 6054 3276 6056 3356
rect 6060 3276 6064 3356
rect 6068 3276 6070 3356
rect 6082 3316 6086 3356
rect 6090 3316 6092 3356
rect 6163 3316 6165 3356
rect 6169 3316 6171 3356
rect 6183 3316 6185 3356
rect 6189 3316 6191 3356
rect 6243 3276 6245 3356
rect 6249 3276 6251 3356
rect 6263 3276 6265 3356
rect 6269 3288 6271 3356
rect 6283 3288 6285 3356
rect 6269 3276 6285 3288
rect 6289 3284 6291 3356
rect 6343 3316 6345 3356
rect 6349 3316 6351 3356
rect 6363 3316 6365 3356
rect 6369 3316 6371 3356
rect 6289 3276 6303 3284
rect 6414 3276 6416 3356
rect 6420 3276 6424 3356
rect 6428 3276 6430 3356
rect 6442 3316 6446 3356
rect 6450 3316 6452 3356
rect 6509 3276 6511 3356
rect 6515 3336 6517 3356
rect 6529 3336 6533 3356
rect 6537 3336 6541 3356
rect 6545 3336 6547 3356
rect 6559 3336 6561 3356
rect 6515 3276 6524 3336
rect 6550 3316 6561 3336
rect 6565 3316 6569 3356
rect 6573 3316 6575 3356
rect 6613 3316 6615 3356
rect 6619 3316 6621 3356
rect 6633 3316 6635 3356
rect 6639 3316 6647 3356
rect 6651 3316 6653 3356
rect 6665 3316 6667 3356
rect 6671 3316 6681 3356
rect 6685 3316 6687 3356
rect 6699 3316 6701 3356
rect 6692 3276 6701 3316
rect 6705 3276 6707 3356
rect 29 2904 31 2984
rect 35 2904 37 2984
rect 49 2904 51 2984
rect 55 2904 57 2984
rect 69 2904 71 2984
rect 75 2904 77 2984
rect 89 2904 91 2984
rect 95 2904 97 2984
rect 109 2904 111 2984
rect 115 2904 117 2984
rect 129 2904 131 2984
rect 135 2904 137 2984
rect 149 2904 151 2984
rect 155 2904 157 2984
rect 169 2904 171 2984
rect 175 2904 177 2984
rect 241 2904 243 2984
rect 247 2904 249 2984
rect 261 2904 265 2944
rect 269 2904 271 2944
rect 313 2904 315 2984
rect 319 2944 328 2984
rect 319 2904 321 2944
rect 333 2904 335 2944
rect 339 2904 349 2944
rect 353 2904 355 2944
rect 367 2904 369 2944
rect 373 2904 381 2944
rect 385 2904 387 2944
rect 399 2904 401 2944
rect 405 2904 407 2944
rect 445 2904 447 2944
rect 451 2904 455 2944
rect 459 2924 470 2944
rect 496 2924 505 2984
rect 459 2904 461 2924
rect 473 2904 475 2924
rect 479 2904 483 2924
rect 487 2904 491 2924
rect 503 2904 505 2924
rect 509 2904 511 2984
rect 563 2904 565 2944
rect 569 2904 571 2944
rect 583 2904 585 2944
rect 589 2904 591 2944
rect 629 2904 631 2944
rect 635 2904 637 2944
rect 649 2904 651 2944
rect 655 2904 657 2944
rect 728 2904 730 2944
rect 734 2904 738 2944
rect 750 2904 752 2984
rect 756 2904 760 2984
rect 764 2904 766 2984
rect 957 2976 971 2984
rect 823 2904 825 2944
rect 829 2904 831 2944
rect 843 2904 845 2944
rect 849 2904 851 2944
rect 903 2904 905 2944
rect 909 2904 911 2944
rect 923 2904 925 2944
rect 929 2904 931 2944
rect 969 2904 971 2976
rect 975 2972 991 2984
rect 975 2904 977 2972
rect 989 2904 991 2972
rect 995 2904 997 2984
rect 1009 2904 1011 2984
rect 1015 2904 1017 2984
rect 1069 2904 1071 2984
rect 1075 2924 1084 2984
rect 1252 2944 1261 2984
rect 1110 2924 1121 2944
rect 1075 2904 1077 2924
rect 1089 2904 1093 2924
rect 1097 2904 1101 2924
rect 1105 2904 1107 2924
rect 1119 2904 1121 2924
rect 1125 2904 1129 2944
rect 1133 2904 1135 2944
rect 1173 2904 1175 2944
rect 1179 2904 1181 2944
rect 1193 2904 1195 2944
rect 1199 2904 1207 2944
rect 1211 2904 1213 2944
rect 1225 2904 1227 2944
rect 1231 2904 1241 2944
rect 1245 2904 1247 2944
rect 1259 2904 1261 2944
rect 1265 2904 1267 2984
rect 1323 2904 1325 2944
rect 1329 2904 1331 2944
rect 1343 2904 1345 2944
rect 1349 2904 1351 2944
rect 1389 2904 1391 2984
rect 1395 2924 1404 2984
rect 1572 2944 1581 2984
rect 1430 2924 1441 2944
rect 1395 2904 1397 2924
rect 1409 2904 1413 2924
rect 1417 2904 1421 2924
rect 1425 2904 1427 2924
rect 1439 2904 1441 2924
rect 1445 2904 1449 2944
rect 1453 2904 1455 2944
rect 1493 2904 1495 2944
rect 1499 2904 1501 2944
rect 1513 2904 1515 2944
rect 1519 2904 1527 2944
rect 1531 2904 1533 2944
rect 1545 2904 1547 2944
rect 1551 2904 1561 2944
rect 1565 2904 1567 2944
rect 1579 2904 1581 2944
rect 1585 2904 1587 2984
rect 1643 2904 1645 2944
rect 1649 2904 1651 2944
rect 1708 2904 1710 2944
rect 1714 2904 1718 2944
rect 1730 2904 1732 2984
rect 1736 2904 1740 2984
rect 1744 2904 1746 2984
rect 1815 2904 1817 2984
rect 1821 2904 1825 2984
rect 1829 2904 1831 2984
rect 1879 2904 1881 2984
rect 1885 2904 1887 2984
rect 1899 2904 1903 2944
rect 1907 2904 1911 2944
rect 1923 2904 1925 2944
rect 1929 2904 1931 2944
rect 1974 2904 1976 2984
rect 1980 2904 1984 2984
rect 1988 2904 1990 2984
rect 2002 2904 2006 2944
rect 2010 2904 2012 2944
rect 2083 2904 2085 2984
rect 2089 2904 2091 2984
rect 2103 2904 2105 2984
rect 2109 2972 2125 2984
rect 2109 2904 2111 2972
rect 2123 2904 2125 2972
rect 2129 2976 2143 2984
rect 2129 2904 2131 2976
rect 2169 2904 2171 2944
rect 2175 2904 2177 2944
rect 2189 2904 2191 2944
rect 2195 2904 2197 2944
rect 2263 2904 2265 2944
rect 2269 2904 2271 2944
rect 2309 2904 2311 2944
rect 2315 2904 2317 2944
rect 2329 2904 2333 2944
rect 2337 2904 2341 2944
rect 2353 2904 2355 2984
rect 2359 2904 2361 2984
rect 2413 2904 2415 2984
rect 2419 2944 2428 2984
rect 2419 2904 2421 2944
rect 2433 2904 2435 2944
rect 2439 2904 2449 2944
rect 2453 2904 2455 2944
rect 2467 2904 2469 2944
rect 2473 2904 2481 2944
rect 2485 2904 2487 2944
rect 2499 2904 2501 2944
rect 2505 2904 2507 2944
rect 2545 2904 2547 2944
rect 2551 2904 2555 2944
rect 2559 2924 2570 2944
rect 2596 2924 2605 2984
rect 2559 2904 2561 2924
rect 2573 2904 2575 2924
rect 2579 2904 2583 2924
rect 2587 2904 2591 2924
rect 2603 2904 2605 2924
rect 2609 2904 2611 2984
rect 2649 2904 2651 2944
rect 2655 2904 2657 2944
rect 2709 2904 2711 2984
rect 2715 2904 2719 2984
rect 2723 2904 2725 2984
rect 2803 2904 2805 2944
rect 2809 2904 2811 2944
rect 2868 2904 2870 2944
rect 2874 2904 2878 2944
rect 2890 2904 2892 2984
rect 2896 2904 2900 2984
rect 2904 2904 2906 2984
rect 2949 2904 2951 2984
rect 2955 2904 2957 2984
rect 3023 2904 3025 2944
rect 3029 2940 3045 2944
rect 3029 2904 3031 2940
rect 3043 2904 3045 2940
rect 3049 2904 3051 2944
rect 3063 2904 3065 2944
rect 3069 2904 3071 2944
rect 3123 2904 3125 2944
rect 3129 2904 3131 2944
rect 3143 2904 3145 2944
rect 3149 2904 3151 2944
rect 3208 2904 3210 2944
rect 3214 2904 3218 2944
rect 3230 2904 3232 2984
rect 3236 2904 3240 2984
rect 3244 2904 3246 2984
rect 3289 2904 3291 2944
rect 3295 2904 3297 2944
rect 3309 2904 3311 2944
rect 3315 2904 3317 2944
rect 3369 2904 3371 2944
rect 3375 2904 3377 2944
rect 3389 2904 3391 2944
rect 3395 2904 3397 2944
rect 3454 2904 3456 2984
rect 3460 2904 3464 2984
rect 3468 2904 3470 2984
rect 3482 2904 3486 2944
rect 3490 2904 3492 2944
rect 3549 2904 3551 2944
rect 3555 2904 3557 2944
rect 3569 2904 3573 2944
rect 3577 2904 3581 2944
rect 3593 2904 3595 2984
rect 3599 2904 3601 2984
rect 3663 2904 3665 2984
rect 3669 2916 3671 2984
rect 3683 2916 3685 2984
rect 3669 2904 3685 2916
rect 3689 2982 3705 2984
rect 3689 2904 3691 2982
rect 3703 2904 3705 2982
rect 3709 2970 3725 2984
rect 3709 2904 3711 2970
rect 3723 2904 3725 2970
rect 3729 2982 3743 2984
rect 3729 2904 3731 2982
rect 3783 2904 3785 2984
rect 3789 2904 3791 2984
rect 3803 2904 3805 2984
rect 3809 2906 3811 2984
rect 3809 2904 3823 2906
rect 3853 2904 3855 2984
rect 3859 2944 3868 2984
rect 3859 2904 3861 2944
rect 3873 2904 3875 2944
rect 3879 2904 3889 2944
rect 3893 2904 3895 2944
rect 3907 2904 3909 2944
rect 3913 2904 3921 2944
rect 3925 2904 3927 2944
rect 3939 2904 3941 2944
rect 3945 2904 3947 2944
rect 3985 2904 3987 2944
rect 3991 2904 3995 2944
rect 3999 2924 4010 2944
rect 4036 2924 4045 2984
rect 3999 2904 4001 2924
rect 4013 2904 4015 2924
rect 4019 2904 4023 2924
rect 4027 2904 4031 2924
rect 4043 2904 4045 2924
rect 4049 2904 4051 2984
rect 4094 2904 4096 2984
rect 4100 2904 4104 2984
rect 4108 2904 4110 2984
rect 4122 2904 4126 2944
rect 4130 2904 4132 2944
rect 4203 2904 4205 2944
rect 4209 2940 4225 2944
rect 4209 2904 4211 2940
rect 4223 2904 4225 2940
rect 4229 2904 4231 2944
rect 4243 2904 4245 2944
rect 4249 2904 4251 2944
rect 4293 2904 4295 2984
rect 4299 2944 4308 2984
rect 4299 2904 4301 2944
rect 4313 2904 4315 2944
rect 4319 2904 4329 2944
rect 4333 2904 4335 2944
rect 4347 2904 4349 2944
rect 4353 2904 4361 2944
rect 4365 2904 4367 2944
rect 4379 2904 4381 2944
rect 4385 2904 4387 2944
rect 4425 2904 4427 2944
rect 4431 2904 4435 2944
rect 4439 2924 4450 2944
rect 4476 2924 4485 2984
rect 4439 2904 4441 2924
rect 4453 2904 4455 2924
rect 4459 2904 4463 2924
rect 4467 2904 4471 2924
rect 4483 2904 4485 2924
rect 4489 2904 4491 2984
rect 4553 2904 4555 2984
rect 4559 2904 4565 2984
rect 4569 2904 4571 2984
rect 4593 2904 4595 2984
rect 4599 2904 4605 2984
rect 4609 2904 4611 2984
rect 4747 2984 4755 2992
rect 4663 2904 4665 2944
rect 4669 2904 4671 2944
rect 4723 2904 4725 2984
rect 4729 2904 4735 2984
rect 4739 2976 4755 2984
rect 4739 2912 4741 2976
rect 4753 2912 4755 2976
rect 4759 2912 4765 2992
rect 4769 2952 4779 2992
rect 4817 2982 4831 2984
rect 4769 2912 4771 2952
rect 4783 2912 4785 2952
rect 4789 2912 4791 2952
rect 4739 2904 4748 2912
rect 4829 2904 4831 2982
rect 4835 2970 4851 2984
rect 4835 2904 4837 2970
rect 4849 2904 4851 2970
rect 4855 2982 4871 2984
rect 4855 2904 4857 2982
rect 4869 2904 4871 2982
rect 4875 2916 4877 2984
rect 4889 2916 4891 2984
rect 4875 2904 4891 2916
rect 4895 2904 4897 2984
rect 4997 2982 5011 2984
rect 4963 2904 4965 2944
rect 4969 2904 4971 2944
rect 5009 2904 5011 2982
rect 5015 2970 5031 2984
rect 5015 2904 5017 2970
rect 5029 2904 5031 2970
rect 5035 2982 5051 2984
rect 5035 2904 5037 2982
rect 5049 2904 5051 2982
rect 5055 2916 5057 2984
rect 5069 2916 5071 2984
rect 5055 2904 5071 2916
rect 5075 2904 5077 2984
rect 5129 2904 5131 2944
rect 5135 2904 5137 2944
rect 5189 2904 5191 2984
rect 5195 2904 5199 2984
rect 5203 2904 5205 2984
rect 5273 2904 5275 2984
rect 5279 2944 5288 2984
rect 5279 2904 5281 2944
rect 5293 2904 5295 2944
rect 5299 2904 5309 2944
rect 5313 2904 5315 2944
rect 5327 2904 5329 2944
rect 5333 2904 5341 2944
rect 5345 2904 5347 2944
rect 5359 2904 5361 2944
rect 5365 2904 5367 2944
rect 5405 2904 5407 2944
rect 5411 2904 5415 2944
rect 5419 2924 5430 2944
rect 5456 2924 5465 2984
rect 5419 2904 5421 2924
rect 5433 2904 5435 2924
rect 5439 2904 5443 2924
rect 5447 2904 5451 2924
rect 5463 2904 5465 2924
rect 5469 2904 5471 2984
rect 5535 2904 5537 2984
rect 5541 2904 5545 2984
rect 5549 2904 5551 2984
rect 5594 2904 5596 2984
rect 5600 2904 5604 2984
rect 5608 2904 5610 2984
rect 5622 2904 5626 2944
rect 5630 2904 5632 2944
rect 5703 2904 5705 2944
rect 5709 2940 5725 2944
rect 5709 2904 5711 2940
rect 5723 2904 5725 2940
rect 5729 2904 5731 2944
rect 5743 2904 5745 2944
rect 5749 2904 5751 2944
rect 5813 2904 5815 2984
rect 5819 2904 5825 2984
rect 5829 2904 5831 2984
rect 5853 2904 5855 2984
rect 5859 2904 5865 2984
rect 5869 2904 5871 2984
rect 5981 2952 5991 2992
rect 5909 2904 5911 2944
rect 5915 2904 5917 2944
rect 5969 2912 5971 2952
rect 5975 2912 5977 2952
rect 5989 2912 5991 2952
rect 5995 2912 6001 2992
rect 6005 2984 6013 2992
rect 6005 2976 6021 2984
rect 6005 2912 6007 2976
rect 6019 2912 6021 2976
rect 6012 2904 6021 2912
rect 6025 2904 6031 2984
rect 6035 2904 6037 2984
rect 6103 2904 6105 2984
rect 6109 2904 6111 2984
rect 6123 2904 6125 2984
rect 6129 2972 6145 2984
rect 6129 2904 6131 2972
rect 6143 2904 6145 2972
rect 6149 2976 6163 2984
rect 6149 2904 6151 2976
rect 6215 2904 6217 2984
rect 6221 2904 6225 2984
rect 6229 2904 6231 2984
rect 6269 2904 6271 2944
rect 6275 2904 6277 2944
rect 6343 2904 6345 2984
rect 6349 2916 6351 2984
rect 6363 2916 6365 2984
rect 6349 2904 6365 2916
rect 6369 2982 6385 2984
rect 6369 2904 6371 2982
rect 6383 2904 6385 2982
rect 6389 2970 6405 2984
rect 6389 2904 6391 2970
rect 6403 2904 6405 2970
rect 6409 2982 6423 2984
rect 6409 2904 6411 2982
rect 6463 2904 6465 2944
rect 6469 2904 6471 2944
rect 6509 2904 6511 2944
rect 6515 2904 6517 2944
rect 6574 2904 6576 2984
rect 6580 2904 6584 2984
rect 6588 2904 6590 2984
rect 6602 2904 6606 2944
rect 6610 2904 6612 2944
rect 29 2836 31 2876
rect 35 2836 37 2876
rect 115 2796 117 2876
rect 121 2796 125 2876
rect 129 2796 131 2876
rect 173 2796 175 2876
rect 179 2836 181 2876
rect 193 2836 195 2876
rect 199 2836 209 2876
rect 213 2836 215 2876
rect 227 2836 229 2876
rect 233 2836 241 2876
rect 245 2836 247 2876
rect 259 2836 261 2876
rect 265 2836 267 2876
rect 305 2836 307 2876
rect 311 2836 315 2876
rect 319 2856 321 2876
rect 333 2856 335 2876
rect 339 2856 343 2876
rect 347 2856 351 2876
rect 363 2856 365 2876
rect 319 2836 330 2856
rect 179 2796 188 2836
rect 356 2796 365 2856
rect 369 2796 371 2876
rect 409 2836 411 2876
rect 415 2836 417 2876
rect 495 2796 497 2876
rect 501 2796 505 2876
rect 509 2796 511 2876
rect 553 2796 555 2876
rect 559 2836 561 2876
rect 573 2836 575 2876
rect 579 2836 589 2876
rect 593 2836 595 2876
rect 607 2836 609 2876
rect 613 2836 621 2876
rect 625 2836 627 2876
rect 639 2836 641 2876
rect 645 2836 647 2876
rect 685 2836 687 2876
rect 691 2836 695 2876
rect 699 2856 701 2876
rect 713 2856 715 2876
rect 719 2856 723 2876
rect 727 2856 731 2876
rect 743 2856 745 2876
rect 699 2836 710 2856
rect 559 2796 568 2836
rect 736 2796 745 2856
rect 749 2796 751 2876
rect 801 2796 803 2876
rect 807 2796 809 2876
rect 821 2836 825 2876
rect 829 2836 831 2876
rect 857 2874 871 2876
rect 869 2796 871 2874
rect 875 2796 877 2876
rect 889 2796 891 2876
rect 895 2796 897 2876
rect 949 2836 951 2876
rect 955 2836 957 2876
rect 969 2836 971 2876
rect 975 2836 977 2876
rect 1029 2836 1031 2876
rect 1035 2836 1037 2876
rect 1049 2836 1051 2876
rect 1055 2836 1057 2876
rect 1109 2836 1111 2876
rect 1115 2836 1117 2876
rect 1169 2798 1171 2876
rect 1157 2796 1171 2798
rect 1175 2810 1177 2876
rect 1189 2810 1191 2876
rect 1175 2796 1191 2810
rect 1195 2798 1197 2876
rect 1209 2798 1211 2876
rect 1195 2796 1211 2798
rect 1215 2864 1231 2876
rect 1215 2796 1217 2864
rect 1229 2796 1231 2864
rect 1235 2796 1237 2876
rect 1303 2796 1305 2876
rect 1309 2796 1311 2876
rect 1323 2796 1325 2876
rect 1329 2808 1331 2876
rect 1343 2808 1345 2876
rect 1329 2796 1345 2808
rect 1349 2804 1351 2876
rect 1403 2836 1405 2876
rect 1409 2836 1411 2876
rect 1468 2836 1470 2876
rect 1474 2836 1478 2876
rect 1349 2796 1363 2804
rect 1490 2796 1492 2876
rect 1496 2796 1500 2876
rect 1504 2796 1506 2876
rect 1549 2796 1551 2876
rect 1555 2796 1559 2876
rect 1563 2796 1565 2876
rect 1629 2836 1631 2876
rect 1635 2836 1637 2876
rect 1649 2836 1651 2876
rect 1655 2836 1657 2876
rect 1709 2796 1711 2876
rect 1715 2796 1719 2876
rect 1723 2796 1725 2876
rect 1808 2836 1810 2876
rect 1814 2836 1818 2876
rect 1830 2796 1832 2876
rect 1836 2796 1840 2876
rect 1844 2796 1846 2876
rect 1889 2796 1891 2876
rect 1895 2796 1901 2876
rect 1905 2797 1907 2876
rect 1919 2797 1921 2876
rect 1905 2796 1921 2797
rect 1925 2797 1927 2876
rect 1925 2796 1939 2797
rect 1994 2796 1996 2876
rect 2000 2796 2004 2876
rect 2008 2796 2010 2876
rect 2022 2836 2026 2876
rect 2030 2836 2032 2876
rect 2103 2796 2105 2876
rect 2109 2796 2111 2876
rect 2123 2796 2125 2876
rect 2129 2808 2131 2876
rect 2143 2808 2145 2876
rect 2129 2796 2145 2808
rect 2149 2804 2151 2876
rect 2149 2796 2163 2804
rect 2193 2796 2195 2876
rect 2199 2836 2201 2876
rect 2213 2836 2215 2876
rect 2219 2836 2229 2876
rect 2233 2836 2235 2876
rect 2247 2836 2249 2876
rect 2253 2836 2261 2876
rect 2265 2836 2267 2876
rect 2279 2836 2281 2876
rect 2285 2836 2287 2876
rect 2325 2836 2327 2876
rect 2331 2836 2335 2876
rect 2339 2856 2341 2876
rect 2353 2856 2355 2876
rect 2359 2856 2363 2876
rect 2367 2856 2371 2876
rect 2383 2856 2385 2876
rect 2339 2836 2350 2856
rect 2199 2796 2208 2836
rect 2376 2796 2385 2856
rect 2389 2796 2391 2876
rect 2429 2836 2431 2876
rect 2435 2836 2437 2876
rect 2449 2836 2451 2876
rect 2455 2836 2457 2876
rect 2509 2836 2511 2876
rect 2515 2836 2517 2876
rect 2583 2836 2585 2876
rect 2589 2836 2591 2876
rect 2633 2796 2635 2876
rect 2639 2836 2641 2876
rect 2653 2836 2655 2876
rect 2659 2836 2669 2876
rect 2673 2836 2675 2876
rect 2687 2836 2689 2876
rect 2693 2836 2701 2876
rect 2705 2836 2707 2876
rect 2719 2836 2721 2876
rect 2725 2836 2727 2876
rect 2765 2836 2767 2876
rect 2771 2836 2775 2876
rect 2779 2856 2781 2876
rect 2793 2856 2795 2876
rect 2799 2856 2803 2876
rect 2807 2856 2811 2876
rect 2823 2856 2825 2876
rect 2779 2836 2790 2856
rect 2639 2796 2648 2836
rect 2816 2796 2825 2856
rect 2829 2796 2831 2876
rect 2874 2796 2876 2876
rect 2880 2796 2884 2876
rect 2888 2796 2890 2876
rect 2902 2836 2906 2876
rect 2910 2836 2912 2876
rect 2983 2796 2985 2876
rect 2989 2796 2991 2876
rect 3003 2796 3005 2876
rect 3009 2808 3011 2876
rect 3023 2808 3025 2876
rect 3009 2796 3025 2808
rect 3029 2804 3031 2876
rect 3029 2796 3043 2804
rect 3069 2796 3071 2876
rect 3075 2856 3077 2876
rect 3089 2856 3093 2876
rect 3097 2856 3101 2876
rect 3105 2856 3107 2876
rect 3119 2856 3121 2876
rect 3075 2796 3084 2856
rect 3110 2836 3121 2856
rect 3125 2836 3129 2876
rect 3133 2836 3135 2876
rect 3173 2836 3175 2876
rect 3179 2836 3181 2876
rect 3193 2836 3195 2876
rect 3199 2836 3207 2876
rect 3211 2836 3213 2876
rect 3225 2836 3227 2876
rect 3231 2836 3241 2876
rect 3245 2836 3247 2876
rect 3259 2836 3261 2876
rect 3252 2796 3261 2836
rect 3265 2796 3267 2876
rect 3309 2836 3311 2876
rect 3315 2836 3317 2876
rect 3369 2796 3371 2876
rect 3375 2796 3381 2876
rect 3385 2796 3387 2876
rect 3409 2796 3411 2876
rect 3415 2796 3421 2876
rect 3425 2796 3427 2876
rect 3494 2796 3496 2876
rect 3500 2796 3504 2876
rect 3508 2796 3510 2876
rect 3522 2836 3526 2876
rect 3530 2836 3532 2876
rect 3613 2796 3615 2876
rect 3619 2796 3625 2876
rect 3629 2796 3631 2876
rect 3653 2796 3655 2876
rect 3659 2796 3665 2876
rect 3669 2796 3671 2876
rect 3714 2796 3716 2876
rect 3720 2796 3724 2876
rect 3728 2796 3730 2876
rect 3742 2836 3746 2876
rect 3750 2836 3752 2876
rect 3833 2796 3835 2876
rect 3839 2796 3845 2876
rect 3849 2796 3851 2876
rect 3873 2796 3875 2876
rect 3879 2796 3885 2876
rect 3889 2796 3891 2876
rect 3943 2836 3945 2876
rect 3949 2836 3951 2876
rect 3989 2796 3991 2876
rect 3995 2796 3999 2876
rect 4003 2796 4005 2876
rect 4069 2796 4071 2876
rect 4075 2796 4079 2876
rect 4083 2796 4085 2876
rect 4163 2796 4165 2876
rect 4169 2796 4171 2876
rect 4183 2796 4185 2876
rect 4189 2808 4191 2876
rect 4203 2808 4205 2876
rect 4189 2796 4205 2808
rect 4209 2804 4211 2876
rect 4209 2796 4223 2804
rect 4254 2796 4256 2876
rect 4260 2796 4264 2876
rect 4268 2796 4270 2876
rect 4282 2836 4286 2876
rect 4290 2836 4292 2876
rect 4363 2836 4365 2876
rect 4369 2840 4371 2876
rect 4383 2840 4385 2876
rect 4369 2836 4385 2840
rect 4389 2836 4391 2876
rect 4403 2836 4405 2876
rect 4409 2836 4411 2876
rect 4453 2796 4455 2876
rect 4459 2836 4461 2876
rect 4473 2836 4475 2876
rect 4479 2836 4489 2876
rect 4493 2836 4495 2876
rect 4507 2836 4509 2876
rect 4513 2836 4521 2876
rect 4525 2836 4527 2876
rect 4539 2836 4541 2876
rect 4545 2836 4547 2876
rect 4585 2836 4587 2876
rect 4591 2836 4595 2876
rect 4599 2856 4601 2876
rect 4613 2856 4615 2876
rect 4619 2856 4623 2876
rect 4627 2856 4631 2876
rect 4643 2856 4645 2876
rect 4599 2836 4610 2856
rect 4459 2796 4468 2836
rect 4636 2796 4645 2856
rect 4649 2796 4651 2876
rect 4689 2836 4691 2876
rect 4695 2836 4697 2876
rect 4749 2796 4751 2876
rect 4755 2796 4759 2876
rect 4763 2796 4765 2876
rect 4834 2796 4836 2876
rect 4840 2796 4844 2876
rect 4848 2796 4850 2876
rect 4862 2836 4866 2876
rect 4870 2836 4872 2876
rect 4955 2796 4957 2876
rect 4961 2796 4965 2876
rect 4969 2796 4971 2876
rect 5033 2796 5035 2876
rect 5039 2796 5045 2876
rect 5049 2796 5051 2876
rect 5073 2796 5075 2876
rect 5079 2796 5085 2876
rect 5089 2796 5091 2876
rect 5129 2804 5131 2876
rect 5117 2796 5131 2804
rect 5135 2808 5137 2876
rect 5149 2808 5151 2876
rect 5135 2796 5151 2808
rect 5155 2796 5157 2876
rect 5169 2796 5171 2876
rect 5175 2796 5177 2876
rect 5229 2836 5231 2876
rect 5235 2836 5239 2876
rect 5251 2796 5253 2876
rect 5257 2796 5259 2876
rect 5314 2796 5316 2876
rect 5320 2796 5324 2876
rect 5328 2796 5330 2876
rect 5342 2836 5346 2876
rect 5350 2836 5352 2876
rect 5433 2796 5435 2876
rect 5439 2796 5445 2876
rect 5449 2796 5451 2876
rect 5473 2796 5475 2876
rect 5479 2796 5485 2876
rect 5489 2796 5491 2876
rect 5543 2836 5545 2876
rect 5549 2836 5551 2876
rect 5593 2796 5595 2876
rect 5599 2836 5601 2876
rect 5613 2836 5615 2876
rect 5619 2836 5629 2876
rect 5633 2836 5635 2876
rect 5647 2836 5649 2876
rect 5653 2836 5661 2876
rect 5665 2836 5667 2876
rect 5679 2836 5681 2876
rect 5685 2836 5687 2876
rect 5725 2836 5727 2876
rect 5731 2836 5735 2876
rect 5739 2856 5741 2876
rect 5753 2856 5755 2876
rect 5759 2856 5763 2876
rect 5767 2856 5771 2876
rect 5783 2856 5785 2876
rect 5739 2836 5750 2856
rect 5599 2796 5608 2836
rect 5776 2796 5785 2856
rect 5789 2796 5791 2876
rect 5872 2868 5881 2876
rect 5829 2828 5831 2868
rect 5835 2828 5837 2868
rect 5849 2828 5851 2868
rect 5841 2788 5851 2828
rect 5855 2788 5861 2868
rect 5865 2804 5867 2868
rect 5879 2804 5881 2868
rect 5865 2796 5881 2804
rect 5885 2796 5891 2876
rect 5895 2796 5897 2876
rect 5992 2868 6001 2876
rect 5949 2828 5951 2868
rect 5955 2828 5957 2868
rect 5969 2828 5971 2868
rect 5865 2788 5873 2796
rect 5961 2788 5971 2828
rect 5975 2788 5981 2868
rect 5985 2804 5987 2868
rect 5999 2804 6001 2868
rect 5985 2796 6001 2804
rect 6005 2796 6011 2876
rect 6015 2796 6017 2876
rect 6112 2868 6121 2876
rect 6069 2828 6071 2868
rect 6075 2828 6077 2868
rect 6089 2828 6091 2868
rect 5985 2788 5993 2796
rect 6081 2788 6091 2828
rect 6095 2788 6101 2868
rect 6105 2804 6107 2868
rect 6119 2804 6121 2868
rect 6105 2796 6121 2804
rect 6125 2796 6131 2876
rect 6135 2796 6137 2876
rect 6199 2796 6201 2876
rect 6205 2796 6207 2876
rect 6219 2836 6223 2876
rect 6227 2836 6231 2876
rect 6243 2836 6245 2876
rect 6249 2836 6251 2876
rect 6105 2788 6113 2796
rect 6303 2796 6305 2876
rect 6309 2796 6311 2876
rect 6323 2796 6325 2876
rect 6329 2874 6343 2876
rect 6329 2796 6331 2874
rect 6369 2836 6371 2876
rect 6375 2836 6377 2876
rect 6389 2836 6393 2876
rect 6397 2836 6401 2876
rect 6413 2796 6415 2876
rect 6419 2796 6421 2876
rect 6469 2796 6471 2876
rect 6475 2856 6477 2876
rect 6489 2856 6493 2876
rect 6497 2856 6501 2876
rect 6505 2856 6507 2876
rect 6519 2856 6521 2876
rect 6475 2796 6484 2856
rect 6510 2836 6521 2856
rect 6525 2836 6529 2876
rect 6533 2836 6535 2876
rect 6573 2836 6575 2876
rect 6579 2836 6581 2876
rect 6593 2836 6595 2876
rect 6599 2836 6607 2876
rect 6611 2836 6613 2876
rect 6625 2836 6627 2876
rect 6631 2836 6641 2876
rect 6645 2836 6647 2876
rect 6659 2836 6661 2876
rect 6652 2796 6661 2836
rect 6665 2796 6667 2876
rect 29 2424 31 2504
rect 35 2444 44 2504
rect 212 2464 221 2504
rect 70 2444 81 2464
rect 35 2424 37 2444
rect 49 2424 53 2444
rect 57 2424 61 2444
rect 65 2424 67 2444
rect 79 2424 81 2444
rect 85 2424 89 2464
rect 93 2424 95 2464
rect 133 2424 135 2464
rect 139 2424 141 2464
rect 153 2424 155 2464
rect 159 2424 167 2464
rect 171 2424 173 2464
rect 185 2424 187 2464
rect 191 2424 201 2464
rect 205 2424 207 2464
rect 219 2424 221 2464
rect 225 2424 227 2504
rect 281 2424 283 2504
rect 287 2424 289 2504
rect 301 2424 305 2464
rect 309 2424 311 2464
rect 349 2424 351 2504
rect 355 2444 364 2504
rect 532 2464 541 2504
rect 390 2444 401 2464
rect 355 2424 357 2444
rect 369 2424 373 2444
rect 377 2424 381 2444
rect 385 2424 387 2444
rect 399 2424 401 2444
rect 405 2424 409 2464
rect 413 2424 415 2464
rect 453 2424 455 2464
rect 459 2424 461 2464
rect 473 2424 475 2464
rect 479 2424 487 2464
rect 491 2424 493 2464
rect 505 2424 507 2464
rect 511 2424 521 2464
rect 525 2424 527 2464
rect 539 2424 541 2464
rect 545 2424 547 2504
rect 603 2424 605 2504
rect 609 2424 611 2504
rect 623 2424 625 2504
rect 629 2492 645 2504
rect 629 2424 631 2492
rect 643 2424 645 2492
rect 649 2496 663 2504
rect 649 2424 651 2496
rect 689 2424 691 2464
rect 695 2424 697 2464
rect 709 2424 711 2464
rect 715 2424 717 2464
rect 783 2424 785 2464
rect 789 2424 791 2464
rect 803 2424 805 2464
rect 809 2424 811 2464
rect 863 2424 865 2504
rect 869 2424 871 2504
rect 883 2424 885 2504
rect 889 2424 891 2504
rect 903 2424 905 2504
rect 909 2424 911 2504
rect 923 2424 925 2504
rect 929 2424 931 2504
rect 943 2424 945 2504
rect 949 2424 951 2504
rect 963 2424 965 2504
rect 969 2424 971 2504
rect 983 2424 985 2504
rect 989 2424 991 2504
rect 1003 2424 1005 2504
rect 1009 2424 1011 2504
rect 1049 2424 1051 2504
rect 1055 2444 1064 2504
rect 1232 2464 1241 2504
rect 1090 2444 1101 2464
rect 1055 2424 1057 2444
rect 1069 2424 1073 2444
rect 1077 2424 1081 2444
rect 1085 2424 1087 2444
rect 1099 2424 1101 2444
rect 1105 2424 1109 2464
rect 1113 2424 1115 2464
rect 1153 2424 1155 2464
rect 1159 2424 1161 2464
rect 1173 2424 1175 2464
rect 1179 2424 1187 2464
rect 1191 2424 1193 2464
rect 1205 2424 1207 2464
rect 1211 2424 1221 2464
rect 1225 2424 1227 2464
rect 1239 2424 1241 2464
rect 1245 2424 1247 2504
rect 1303 2424 1305 2464
rect 1309 2424 1311 2464
rect 1323 2424 1325 2464
rect 1329 2424 1331 2464
rect 1369 2424 1371 2504
rect 1375 2424 1379 2504
rect 1383 2424 1385 2504
rect 1449 2424 1451 2464
rect 1455 2424 1457 2464
rect 1528 2424 1530 2464
rect 1534 2424 1538 2464
rect 1550 2424 1552 2504
rect 1556 2424 1560 2504
rect 1564 2424 1566 2504
rect 1613 2424 1615 2504
rect 1619 2464 1628 2504
rect 1619 2424 1621 2464
rect 1633 2424 1635 2464
rect 1639 2424 1649 2464
rect 1653 2424 1655 2464
rect 1667 2424 1669 2464
rect 1673 2424 1681 2464
rect 1685 2424 1687 2464
rect 1699 2424 1701 2464
rect 1705 2424 1707 2464
rect 1745 2424 1747 2464
rect 1751 2424 1755 2464
rect 1759 2444 1770 2464
rect 1796 2444 1805 2504
rect 1759 2424 1761 2444
rect 1773 2424 1775 2444
rect 1779 2424 1783 2444
rect 1787 2424 1791 2444
rect 1803 2424 1805 2444
rect 1809 2424 1811 2504
rect 1849 2424 1851 2464
rect 1855 2424 1857 2464
rect 1909 2424 1911 2464
rect 1915 2424 1917 2464
rect 1969 2424 1971 2504
rect 1975 2424 1981 2504
rect 1985 2424 1987 2504
rect 2009 2424 2011 2504
rect 2015 2424 2021 2504
rect 2025 2424 2027 2504
rect 2089 2424 2091 2504
rect 2095 2424 2099 2504
rect 2103 2424 2105 2504
rect 2181 2472 2191 2512
rect 2169 2432 2171 2472
rect 2175 2432 2177 2472
rect 2189 2432 2191 2472
rect 2195 2432 2201 2512
rect 2205 2504 2213 2512
rect 2205 2496 2221 2504
rect 2205 2432 2207 2496
rect 2219 2432 2221 2496
rect 2212 2424 2221 2432
rect 2225 2424 2231 2504
rect 2235 2424 2237 2504
rect 2301 2472 2311 2512
rect 2289 2432 2291 2472
rect 2295 2432 2297 2472
rect 2309 2432 2311 2472
rect 2315 2432 2321 2512
rect 2325 2504 2333 2512
rect 2325 2496 2341 2504
rect 2325 2432 2327 2496
rect 2339 2432 2341 2496
rect 2332 2424 2341 2432
rect 2345 2424 2351 2504
rect 2355 2424 2357 2504
rect 2413 2424 2415 2504
rect 2419 2464 2428 2504
rect 2419 2424 2421 2464
rect 2433 2424 2435 2464
rect 2439 2424 2449 2464
rect 2453 2424 2455 2464
rect 2467 2424 2469 2464
rect 2473 2424 2481 2464
rect 2485 2424 2487 2464
rect 2499 2424 2501 2464
rect 2505 2424 2507 2464
rect 2545 2424 2547 2464
rect 2551 2424 2555 2464
rect 2559 2444 2570 2464
rect 2596 2444 2605 2504
rect 2559 2424 2561 2444
rect 2573 2424 2575 2444
rect 2579 2424 2583 2444
rect 2587 2424 2591 2444
rect 2603 2424 2605 2444
rect 2609 2424 2611 2504
rect 2661 2472 2671 2512
rect 2649 2432 2651 2472
rect 2655 2432 2657 2472
rect 2669 2432 2671 2472
rect 2675 2432 2681 2512
rect 2685 2504 2693 2512
rect 2887 2504 2895 2512
rect 2685 2496 2701 2504
rect 2685 2432 2687 2496
rect 2699 2432 2701 2496
rect 2692 2424 2701 2432
rect 2705 2424 2711 2504
rect 2715 2424 2717 2504
rect 2795 2424 2797 2504
rect 2801 2424 2805 2504
rect 2809 2424 2811 2504
rect 2863 2424 2865 2504
rect 2869 2424 2875 2504
rect 2879 2496 2895 2504
rect 2879 2432 2881 2496
rect 2893 2432 2895 2496
rect 2899 2432 2905 2512
rect 2909 2472 2919 2512
rect 2909 2432 2911 2472
rect 2923 2432 2925 2472
rect 2929 2432 2931 2472
rect 2879 2424 2888 2432
rect 2993 2424 2995 2504
rect 2999 2424 3005 2504
rect 3009 2424 3011 2504
rect 3033 2424 3035 2504
rect 3039 2424 3045 2504
rect 3049 2424 3051 2504
rect 3103 2424 3105 2464
rect 3109 2424 3111 2464
rect 3153 2424 3155 2504
rect 3159 2464 3168 2504
rect 3159 2424 3161 2464
rect 3173 2424 3175 2464
rect 3179 2424 3189 2464
rect 3193 2424 3195 2464
rect 3207 2424 3209 2464
rect 3213 2424 3221 2464
rect 3225 2424 3227 2464
rect 3239 2424 3241 2464
rect 3245 2424 3247 2464
rect 3285 2424 3287 2464
rect 3291 2424 3295 2464
rect 3299 2444 3310 2464
rect 3336 2444 3345 2504
rect 3299 2424 3301 2444
rect 3313 2424 3315 2444
rect 3319 2424 3323 2444
rect 3327 2424 3331 2444
rect 3343 2424 3345 2444
rect 3349 2424 3351 2504
rect 3389 2424 3391 2504
rect 3395 2424 3399 2504
rect 3403 2424 3405 2504
rect 3483 2424 3485 2464
rect 3489 2424 3491 2464
rect 3503 2424 3505 2464
rect 3509 2424 3511 2464
rect 3549 2424 3551 2464
rect 3555 2424 3557 2464
rect 3609 2424 3611 2464
rect 3615 2424 3617 2464
rect 3629 2424 3631 2464
rect 3635 2460 3651 2464
rect 3635 2424 3637 2460
rect 3649 2424 3651 2460
rect 3655 2424 3657 2464
rect 3709 2424 3711 2464
rect 3715 2424 3717 2464
rect 3729 2424 3731 2464
rect 3735 2460 3751 2464
rect 3735 2424 3737 2460
rect 3749 2424 3751 2460
rect 3755 2424 3757 2464
rect 3823 2424 3825 2464
rect 3829 2460 3845 2464
rect 3829 2424 3831 2460
rect 3843 2424 3845 2460
rect 3849 2424 3851 2464
rect 3863 2424 3865 2464
rect 3869 2424 3871 2464
rect 3914 2424 3916 2504
rect 3920 2424 3924 2504
rect 3928 2424 3930 2504
rect 3997 2496 4011 2504
rect 3942 2424 3946 2464
rect 3950 2424 3952 2464
rect 4009 2424 4011 2496
rect 4015 2492 4031 2504
rect 4015 2424 4017 2492
rect 4029 2424 4031 2492
rect 4035 2424 4037 2504
rect 4049 2424 4051 2504
rect 4055 2424 4057 2504
rect 4135 2424 4137 2504
rect 4141 2424 4145 2504
rect 4149 2424 4151 2504
rect 4213 2424 4215 2504
rect 4219 2424 4225 2504
rect 4229 2424 4231 2504
rect 4253 2424 4255 2504
rect 4259 2424 4265 2504
rect 4269 2424 4271 2504
rect 4313 2424 4315 2504
rect 4319 2464 4328 2504
rect 4319 2424 4321 2464
rect 4333 2424 4335 2464
rect 4339 2424 4349 2464
rect 4353 2424 4355 2464
rect 4367 2424 4369 2464
rect 4373 2424 4381 2464
rect 4385 2424 4387 2464
rect 4399 2424 4401 2464
rect 4405 2424 4407 2464
rect 4445 2424 4447 2464
rect 4451 2424 4455 2464
rect 4459 2444 4470 2464
rect 4496 2444 4505 2504
rect 4459 2424 4461 2444
rect 4473 2424 4475 2444
rect 4479 2424 4483 2444
rect 4487 2424 4491 2444
rect 4503 2424 4505 2444
rect 4509 2424 4511 2504
rect 4563 2424 4565 2464
rect 4569 2424 4571 2464
rect 4633 2424 4635 2504
rect 4639 2424 4645 2504
rect 4649 2424 4651 2504
rect 4673 2424 4675 2504
rect 4679 2424 4685 2504
rect 4689 2424 4691 2504
rect 4741 2472 4751 2512
rect 4729 2432 4731 2472
rect 4735 2432 4737 2472
rect 4749 2432 4751 2472
rect 4755 2432 4761 2512
rect 4765 2504 4773 2512
rect 4765 2496 4781 2504
rect 4765 2432 4767 2496
rect 4779 2432 4781 2496
rect 4772 2424 4781 2432
rect 4785 2424 4791 2504
rect 4795 2424 4797 2504
rect 4849 2424 4851 2504
rect 4855 2444 4864 2504
rect 5032 2464 5041 2504
rect 4890 2444 4901 2464
rect 4855 2424 4857 2444
rect 4869 2424 4873 2444
rect 4877 2424 4881 2444
rect 4885 2424 4887 2444
rect 4899 2424 4901 2444
rect 4905 2424 4909 2464
rect 4913 2424 4915 2464
rect 4953 2424 4955 2464
rect 4959 2424 4961 2464
rect 4973 2424 4975 2464
rect 4979 2424 4987 2464
rect 4991 2424 4993 2464
rect 5005 2424 5007 2464
rect 5011 2424 5021 2464
rect 5025 2424 5027 2464
rect 5039 2424 5041 2464
rect 5045 2424 5047 2504
rect 5089 2424 5091 2464
rect 5095 2424 5097 2464
rect 5149 2424 5151 2504
rect 5155 2424 5161 2504
rect 5165 2424 5167 2504
rect 5189 2424 5191 2504
rect 5195 2424 5201 2504
rect 5205 2424 5207 2504
rect 5274 2424 5276 2504
rect 5280 2424 5284 2504
rect 5288 2424 5290 2504
rect 5302 2424 5306 2464
rect 5310 2424 5312 2464
rect 5369 2424 5371 2504
rect 5375 2424 5379 2504
rect 5383 2424 5385 2504
rect 5475 2424 5477 2504
rect 5481 2424 5485 2504
rect 5489 2424 5491 2504
rect 5529 2424 5531 2504
rect 5535 2424 5537 2504
rect 5549 2424 5551 2504
rect 5555 2424 5557 2504
rect 5569 2424 5571 2504
rect 5575 2424 5577 2504
rect 5589 2424 5591 2504
rect 5595 2424 5597 2504
rect 5609 2424 5611 2504
rect 5615 2424 5617 2504
rect 5629 2424 5631 2504
rect 5635 2424 5637 2504
rect 5649 2424 5651 2504
rect 5655 2424 5657 2504
rect 5669 2424 5671 2504
rect 5675 2424 5677 2504
rect 5755 2424 5757 2504
rect 5761 2424 5765 2504
rect 5769 2424 5771 2504
rect 5814 2424 5816 2504
rect 5820 2424 5824 2504
rect 5828 2424 5830 2504
rect 5842 2424 5846 2464
rect 5850 2424 5852 2464
rect 5933 2424 5935 2504
rect 5939 2424 5945 2504
rect 5949 2424 5951 2504
rect 5973 2424 5975 2504
rect 5979 2424 5985 2504
rect 5989 2424 5991 2504
rect 6043 2424 6045 2464
rect 6049 2424 6051 2464
rect 6089 2424 6091 2504
rect 6095 2444 6104 2504
rect 6272 2464 6281 2504
rect 6130 2444 6141 2464
rect 6095 2424 6097 2444
rect 6109 2424 6113 2444
rect 6117 2424 6121 2444
rect 6125 2424 6127 2444
rect 6139 2424 6141 2444
rect 6145 2424 6149 2464
rect 6153 2424 6155 2464
rect 6193 2424 6195 2464
rect 6199 2424 6201 2464
rect 6213 2424 6215 2464
rect 6219 2424 6227 2464
rect 6231 2424 6233 2464
rect 6245 2424 6247 2464
rect 6251 2424 6261 2464
rect 6265 2424 6267 2464
rect 6279 2424 6281 2464
rect 6285 2424 6287 2504
rect 6343 2424 6345 2504
rect 6349 2436 6351 2504
rect 6363 2436 6365 2504
rect 6349 2424 6365 2436
rect 6369 2502 6385 2504
rect 6369 2424 6371 2502
rect 6383 2424 6385 2502
rect 6389 2490 6405 2504
rect 6389 2424 6391 2490
rect 6403 2424 6405 2490
rect 6409 2502 6423 2504
rect 6409 2424 6411 2502
rect 6449 2426 6451 2504
rect 6437 2424 6451 2426
rect 6455 2424 6457 2504
rect 6469 2424 6471 2504
rect 6475 2424 6477 2504
rect 6577 2502 6591 2504
rect 6529 2424 6531 2464
rect 6535 2424 6537 2464
rect 6589 2424 6591 2502
rect 6595 2490 6611 2504
rect 6595 2424 6597 2490
rect 6609 2424 6611 2490
rect 6615 2502 6631 2504
rect 6615 2424 6617 2502
rect 6629 2424 6631 2502
rect 6635 2436 6637 2504
rect 6649 2436 6651 2504
rect 6635 2424 6651 2436
rect 6655 2424 6657 2504
rect 33 2316 35 2396
rect 39 2356 41 2396
rect 53 2356 55 2396
rect 59 2356 69 2396
rect 73 2356 75 2396
rect 87 2356 89 2396
rect 93 2356 101 2396
rect 105 2356 107 2396
rect 119 2356 121 2396
rect 125 2356 127 2396
rect 165 2356 167 2396
rect 171 2356 175 2396
rect 179 2376 181 2396
rect 193 2376 195 2396
rect 199 2376 203 2396
rect 207 2376 211 2396
rect 223 2376 225 2396
rect 179 2356 190 2376
rect 39 2316 48 2356
rect 216 2316 225 2376
rect 229 2316 231 2396
rect 281 2316 283 2396
rect 287 2316 289 2396
rect 301 2356 305 2396
rect 309 2356 311 2396
rect 363 2316 365 2396
rect 369 2316 371 2396
rect 423 2356 425 2396
rect 429 2356 431 2396
rect 495 2316 497 2396
rect 501 2316 505 2396
rect 509 2316 511 2396
rect 554 2316 556 2396
rect 560 2316 564 2396
rect 568 2316 570 2396
rect 582 2356 586 2396
rect 590 2356 592 2396
rect 659 2316 661 2396
rect 665 2316 667 2396
rect 679 2356 683 2396
rect 687 2356 691 2396
rect 703 2356 705 2396
rect 709 2356 711 2396
rect 749 2356 751 2396
rect 755 2356 757 2396
rect 769 2356 771 2396
rect 775 2360 777 2396
rect 789 2360 791 2396
rect 775 2356 791 2360
rect 795 2356 797 2396
rect 849 2356 851 2396
rect 855 2356 857 2396
rect 869 2356 871 2396
rect 875 2356 877 2396
rect 929 2316 931 2396
rect 935 2376 937 2396
rect 949 2376 953 2396
rect 957 2376 961 2396
rect 965 2376 967 2396
rect 979 2376 981 2396
rect 935 2316 944 2376
rect 970 2356 981 2376
rect 985 2356 989 2396
rect 993 2356 995 2396
rect 1033 2356 1035 2396
rect 1039 2356 1041 2396
rect 1053 2356 1055 2396
rect 1059 2356 1067 2396
rect 1071 2356 1073 2396
rect 1085 2356 1087 2396
rect 1091 2356 1101 2396
rect 1105 2356 1107 2396
rect 1119 2356 1121 2396
rect 1112 2316 1121 2356
rect 1125 2316 1127 2396
rect 1169 2356 1171 2396
rect 1175 2356 1177 2396
rect 1233 2316 1235 2396
rect 1239 2356 1241 2396
rect 1253 2356 1255 2396
rect 1259 2356 1269 2396
rect 1273 2356 1275 2396
rect 1287 2356 1289 2396
rect 1293 2356 1301 2396
rect 1305 2356 1307 2396
rect 1319 2356 1321 2396
rect 1325 2356 1327 2396
rect 1365 2356 1367 2396
rect 1371 2356 1375 2396
rect 1379 2376 1381 2396
rect 1393 2376 1395 2396
rect 1399 2376 1403 2396
rect 1407 2376 1411 2396
rect 1423 2376 1425 2396
rect 1379 2356 1390 2376
rect 1239 2316 1248 2356
rect 1416 2316 1425 2376
rect 1429 2316 1431 2396
rect 1483 2356 1485 2396
rect 1489 2356 1491 2396
rect 1529 2316 1531 2396
rect 1535 2316 1541 2396
rect 1545 2316 1547 2396
rect 1569 2316 1571 2396
rect 1575 2316 1581 2396
rect 1585 2316 1587 2396
rect 1654 2316 1656 2396
rect 1660 2316 1664 2396
rect 1668 2316 1670 2396
rect 1682 2356 1686 2396
rect 1690 2356 1692 2396
rect 1775 2316 1777 2396
rect 1781 2316 1785 2396
rect 1789 2316 1791 2396
rect 1855 2316 1857 2396
rect 1861 2316 1865 2396
rect 1869 2316 1871 2396
rect 1933 2316 1935 2396
rect 1939 2316 1945 2396
rect 1949 2316 1951 2396
rect 1973 2316 1975 2396
rect 1979 2316 1985 2396
rect 1989 2316 1991 2396
rect 2043 2356 2045 2396
rect 2049 2356 2051 2396
rect 2093 2316 2095 2396
rect 2099 2356 2101 2396
rect 2113 2356 2115 2396
rect 2119 2356 2129 2396
rect 2133 2356 2135 2396
rect 2147 2356 2149 2396
rect 2153 2356 2161 2396
rect 2165 2356 2167 2396
rect 2179 2356 2181 2396
rect 2185 2356 2187 2396
rect 2225 2356 2227 2396
rect 2231 2356 2235 2396
rect 2239 2376 2241 2396
rect 2253 2376 2255 2396
rect 2259 2376 2263 2396
rect 2267 2376 2271 2396
rect 2283 2376 2285 2396
rect 2239 2356 2250 2376
rect 2099 2316 2108 2356
rect 2276 2316 2285 2376
rect 2289 2316 2291 2396
rect 2355 2316 2357 2396
rect 2361 2316 2365 2396
rect 2369 2316 2371 2396
rect 2414 2316 2416 2396
rect 2420 2316 2424 2396
rect 2428 2316 2430 2396
rect 2442 2356 2446 2396
rect 2450 2356 2452 2396
rect 2523 2356 2525 2396
rect 2529 2360 2531 2396
rect 2543 2360 2545 2396
rect 2529 2356 2545 2360
rect 2549 2356 2551 2396
rect 2563 2356 2565 2396
rect 2569 2356 2571 2396
rect 2623 2316 2625 2396
rect 2629 2316 2631 2396
rect 2643 2316 2645 2396
rect 2649 2328 2651 2396
rect 2663 2328 2665 2396
rect 2649 2316 2665 2328
rect 2669 2324 2671 2396
rect 2669 2316 2683 2324
rect 2714 2316 2716 2396
rect 2720 2316 2724 2396
rect 2728 2316 2730 2396
rect 2742 2356 2746 2396
rect 2750 2356 2752 2396
rect 2835 2316 2837 2396
rect 2841 2316 2845 2396
rect 2849 2316 2851 2396
rect 2889 2316 2891 2396
rect 2895 2376 2897 2396
rect 2909 2376 2913 2396
rect 2917 2376 2921 2396
rect 2925 2376 2927 2396
rect 2939 2376 2941 2396
rect 2895 2316 2904 2376
rect 2930 2356 2941 2376
rect 2945 2356 2949 2396
rect 2953 2356 2955 2396
rect 2993 2356 2995 2396
rect 2999 2356 3001 2396
rect 3013 2356 3015 2396
rect 3019 2356 3027 2396
rect 3031 2356 3033 2396
rect 3045 2356 3047 2396
rect 3051 2356 3061 2396
rect 3065 2356 3067 2396
rect 3079 2356 3081 2396
rect 3072 2316 3081 2356
rect 3085 2316 3087 2396
rect 3134 2316 3136 2396
rect 3140 2316 3144 2396
rect 3148 2316 3150 2396
rect 3162 2356 3166 2396
rect 3170 2356 3172 2396
rect 3253 2316 3255 2396
rect 3259 2316 3265 2396
rect 3269 2316 3271 2396
rect 3293 2316 3295 2396
rect 3299 2316 3305 2396
rect 3309 2316 3311 2396
rect 3375 2316 3377 2396
rect 3381 2316 3385 2396
rect 3389 2316 3391 2396
rect 3443 2356 3445 2396
rect 3449 2356 3451 2396
rect 3515 2316 3517 2396
rect 3521 2316 3525 2396
rect 3529 2316 3531 2396
rect 3573 2316 3575 2396
rect 3579 2356 3581 2396
rect 3593 2356 3595 2396
rect 3599 2356 3609 2396
rect 3613 2356 3615 2396
rect 3627 2356 3629 2396
rect 3633 2356 3641 2396
rect 3645 2356 3647 2396
rect 3659 2356 3661 2396
rect 3665 2356 3667 2396
rect 3705 2356 3707 2396
rect 3711 2356 3715 2396
rect 3719 2376 3721 2396
rect 3733 2376 3735 2396
rect 3739 2376 3743 2396
rect 3747 2376 3751 2396
rect 3763 2376 3765 2396
rect 3719 2356 3730 2376
rect 3579 2316 3588 2356
rect 3756 2316 3765 2376
rect 3769 2316 3771 2396
rect 3809 2356 3811 2396
rect 3815 2356 3817 2396
rect 3829 2356 3831 2396
rect 3835 2356 3837 2396
rect 3889 2356 3891 2396
rect 3895 2356 3897 2396
rect 3909 2356 3911 2396
rect 3915 2360 3917 2396
rect 3929 2360 3931 2396
rect 3915 2356 3931 2360
rect 3935 2356 3937 2396
rect 4032 2388 4041 2396
rect 3989 2348 3991 2388
rect 3995 2348 3997 2388
rect 4009 2348 4011 2388
rect 4001 2308 4011 2348
rect 4015 2308 4021 2388
rect 4025 2324 4027 2388
rect 4039 2324 4041 2388
rect 4025 2316 4041 2324
rect 4045 2316 4051 2396
rect 4055 2316 4057 2396
rect 4152 2388 4161 2396
rect 4109 2348 4111 2388
rect 4115 2348 4117 2388
rect 4129 2348 4131 2388
rect 4025 2308 4033 2316
rect 4121 2308 4131 2348
rect 4135 2308 4141 2388
rect 4145 2324 4147 2388
rect 4159 2324 4161 2388
rect 4145 2316 4161 2324
rect 4165 2316 4171 2396
rect 4175 2316 4177 2396
rect 4272 2388 4281 2396
rect 4229 2348 4231 2388
rect 4235 2348 4237 2388
rect 4249 2348 4251 2388
rect 4145 2308 4153 2316
rect 4241 2308 4251 2348
rect 4255 2308 4261 2388
rect 4265 2324 4267 2388
rect 4279 2324 4281 2388
rect 4265 2316 4281 2324
rect 4285 2316 4291 2396
rect 4295 2316 4297 2396
rect 4349 2356 4351 2396
rect 4355 2356 4359 2396
rect 4265 2308 4273 2316
rect 4371 2316 4373 2396
rect 4377 2316 4379 2396
rect 4455 2316 4457 2396
rect 4461 2316 4465 2396
rect 4469 2316 4471 2396
rect 4552 2388 4561 2396
rect 4509 2348 4511 2388
rect 4515 2348 4517 2388
rect 4529 2348 4531 2388
rect 4521 2308 4531 2348
rect 4535 2308 4541 2388
rect 4545 2324 4547 2388
rect 4559 2324 4561 2388
rect 4545 2316 4561 2324
rect 4565 2316 4571 2396
rect 4575 2316 4577 2396
rect 4643 2316 4645 2396
rect 4649 2316 4655 2396
rect 4659 2388 4668 2396
rect 4792 2388 4801 2396
rect 4659 2324 4661 2388
rect 4673 2324 4675 2388
rect 4659 2316 4675 2324
rect 4545 2308 4553 2316
rect 4667 2308 4675 2316
rect 4679 2308 4685 2388
rect 4689 2348 4691 2388
rect 4703 2348 4705 2388
rect 4709 2348 4711 2388
rect 4749 2348 4751 2388
rect 4755 2348 4757 2388
rect 4769 2348 4771 2388
rect 4689 2308 4699 2348
rect 4761 2308 4771 2348
rect 4775 2308 4781 2388
rect 4785 2324 4787 2388
rect 4799 2324 4801 2388
rect 4785 2316 4801 2324
rect 4805 2316 4811 2396
rect 4815 2316 4817 2396
rect 4869 2316 4871 2396
rect 4875 2316 4879 2396
rect 4883 2316 4885 2396
rect 4992 2388 5001 2396
rect 4949 2348 4951 2388
rect 4955 2348 4957 2388
rect 4969 2348 4971 2388
rect 4785 2308 4793 2316
rect 4961 2308 4971 2348
rect 4975 2308 4981 2388
rect 4985 2324 4987 2388
rect 4999 2324 5001 2388
rect 4985 2316 5001 2324
rect 5005 2316 5011 2396
rect 5015 2316 5017 2396
rect 5083 2316 5085 2396
rect 5089 2316 5091 2396
rect 5103 2316 5105 2396
rect 5109 2328 5111 2396
rect 5123 2328 5125 2396
rect 5109 2316 5125 2328
rect 5129 2324 5131 2396
rect 5169 2356 5171 2396
rect 5175 2356 5177 2396
rect 5129 2316 5143 2324
rect 4985 2308 4993 2316
rect 5229 2316 5231 2396
rect 5235 2316 5241 2396
rect 5245 2316 5247 2396
rect 5269 2316 5271 2396
rect 5275 2316 5281 2396
rect 5285 2316 5287 2396
rect 5363 2316 5365 2396
rect 5369 2316 5375 2396
rect 5379 2388 5388 2396
rect 5512 2388 5521 2396
rect 5379 2324 5381 2388
rect 5393 2324 5395 2388
rect 5379 2316 5395 2324
rect 5387 2308 5395 2316
rect 5399 2308 5405 2388
rect 5409 2348 5411 2388
rect 5423 2348 5425 2388
rect 5429 2348 5431 2388
rect 5469 2348 5471 2388
rect 5475 2348 5477 2388
rect 5489 2348 5491 2388
rect 5409 2308 5419 2348
rect 5481 2308 5491 2348
rect 5495 2308 5501 2388
rect 5505 2324 5507 2388
rect 5519 2324 5521 2388
rect 5505 2316 5521 2324
rect 5525 2316 5531 2396
rect 5535 2316 5537 2396
rect 5632 2388 5641 2396
rect 5589 2348 5591 2388
rect 5595 2348 5597 2388
rect 5609 2348 5611 2388
rect 5505 2308 5513 2316
rect 5601 2308 5611 2348
rect 5615 2308 5621 2388
rect 5625 2324 5627 2388
rect 5639 2324 5641 2388
rect 5625 2316 5641 2324
rect 5645 2316 5651 2396
rect 5655 2316 5657 2396
rect 5723 2356 5725 2396
rect 5729 2360 5731 2396
rect 5743 2360 5745 2396
rect 5729 2356 5745 2360
rect 5749 2356 5751 2396
rect 5763 2356 5765 2396
rect 5769 2356 5771 2396
rect 5823 2356 5825 2396
rect 5829 2360 5831 2396
rect 5843 2360 5845 2396
rect 5829 2356 5845 2360
rect 5849 2356 5851 2396
rect 5863 2356 5865 2396
rect 5869 2356 5871 2396
rect 5923 2356 5925 2396
rect 5929 2356 5931 2396
rect 5625 2308 5633 2316
rect 5983 2316 5985 2396
rect 5989 2384 6005 2396
rect 5989 2316 5991 2384
rect 6003 2316 6005 2384
rect 6009 2318 6011 2396
rect 6023 2318 6025 2396
rect 6009 2316 6025 2318
rect 6029 2330 6031 2396
rect 6043 2330 6045 2396
rect 6029 2316 6045 2330
rect 6049 2318 6051 2396
rect 6049 2316 6063 2318
rect 6103 2316 6105 2396
rect 6109 2316 6115 2396
rect 6119 2388 6128 2396
rect 6119 2324 6121 2388
rect 6133 2324 6135 2388
rect 6119 2316 6135 2324
rect 6127 2308 6135 2316
rect 6139 2308 6145 2388
rect 6149 2348 6151 2388
rect 6163 2348 6165 2388
rect 6169 2348 6171 2388
rect 6149 2308 6159 2348
rect 6223 2316 6225 2396
rect 6229 2316 6235 2396
rect 6239 2388 6248 2396
rect 6239 2324 6241 2388
rect 6253 2324 6255 2388
rect 6239 2316 6255 2324
rect 6247 2308 6255 2316
rect 6259 2308 6265 2388
rect 6269 2348 6271 2388
rect 6283 2348 6285 2388
rect 6289 2348 6291 2388
rect 6329 2356 6331 2396
rect 6335 2356 6337 2396
rect 6269 2308 6279 2348
rect 6394 2316 6396 2396
rect 6400 2316 6404 2396
rect 6408 2316 6410 2396
rect 6422 2356 6426 2396
rect 6430 2356 6432 2396
rect 6489 2356 6491 2396
rect 6495 2356 6497 2396
rect 6509 2356 6511 2396
rect 6515 2356 6517 2396
rect 6569 2324 6571 2396
rect 6557 2316 6571 2324
rect 6575 2328 6577 2396
rect 6589 2328 6591 2396
rect 6575 2316 6591 2328
rect 6595 2316 6597 2396
rect 6609 2316 6611 2396
rect 6615 2316 6617 2396
rect 6669 2356 6671 2396
rect 6675 2356 6677 2396
rect 55 1944 57 2024
rect 61 1944 65 2024
rect 69 1944 71 2024
rect 123 1944 125 1984
rect 129 1944 131 1984
rect 143 1944 145 1984
rect 149 1944 151 1984
rect 203 1944 205 1984
rect 209 1980 225 1984
rect 209 1944 211 1980
rect 223 1944 225 1980
rect 229 1944 231 1984
rect 243 1944 245 1984
rect 249 1944 251 1984
rect 303 1944 305 1984
rect 309 1980 325 1984
rect 309 1944 311 1980
rect 323 1944 325 1980
rect 329 1944 331 1984
rect 343 1944 345 1984
rect 349 1944 351 1984
rect 403 1944 405 1984
rect 409 1944 411 1984
rect 423 1944 425 1984
rect 429 1944 431 1984
rect 469 1944 471 1984
rect 475 1944 477 1984
rect 489 1944 491 1984
rect 495 1980 511 1984
rect 495 1944 497 1980
rect 509 1944 511 1980
rect 515 1944 517 1984
rect 595 1944 597 2024
rect 601 1944 605 2024
rect 609 1944 611 2024
rect 654 1944 656 2024
rect 660 1944 664 2024
rect 668 1944 670 2024
rect 682 1944 686 1984
rect 690 1944 692 1984
rect 749 1944 751 1984
rect 755 1944 757 1984
rect 769 1944 771 1984
rect 775 1980 791 1984
rect 775 1944 777 1980
rect 789 1944 791 1980
rect 795 1944 797 1984
rect 849 1944 851 2024
rect 855 1944 859 2024
rect 863 1944 865 2024
rect 1021 1992 1031 2032
rect 943 1944 945 1984
rect 949 1944 951 1984
rect 963 1944 965 1984
rect 969 1944 971 1984
rect 1009 1952 1011 1992
rect 1015 1952 1017 1992
rect 1029 1952 1031 1992
rect 1035 1952 1041 2032
rect 1045 2024 1053 2032
rect 1045 2016 1061 2024
rect 1045 1952 1047 2016
rect 1059 1952 1061 2016
rect 1052 1944 1061 1952
rect 1065 1944 1071 2024
rect 1075 1944 1077 2024
rect 1133 1944 1135 2024
rect 1139 1984 1148 2024
rect 1139 1944 1141 1984
rect 1153 1944 1155 1984
rect 1159 1944 1169 1984
rect 1173 1944 1175 1984
rect 1187 1944 1189 1984
rect 1193 1944 1201 1984
rect 1205 1944 1207 1984
rect 1219 1944 1221 1984
rect 1225 1944 1227 1984
rect 1265 1944 1267 1984
rect 1271 1944 1275 1984
rect 1279 1964 1290 1984
rect 1316 1964 1325 2024
rect 1279 1944 1281 1964
rect 1293 1944 1295 1964
rect 1299 1944 1303 1964
rect 1307 1944 1311 1964
rect 1323 1944 1325 1964
rect 1329 1944 1331 2024
rect 1369 1944 1371 1984
rect 1375 1944 1377 1984
rect 1429 1944 1431 2024
rect 1435 1944 1441 2024
rect 1445 1944 1447 2024
rect 1469 1944 1471 2024
rect 1475 1944 1481 2024
rect 1485 1944 1487 2024
rect 1568 1944 1570 1984
rect 1574 1944 1578 1984
rect 1590 1944 1592 2024
rect 1596 1944 1600 2024
rect 1604 1944 1606 2024
rect 1668 1944 1670 1984
rect 1674 1944 1678 1984
rect 1690 1944 1692 2024
rect 1696 1944 1700 2024
rect 1704 1944 1706 2024
rect 1775 1944 1777 2024
rect 1781 1944 1785 2024
rect 1789 1944 1791 2024
rect 1967 2024 1975 2032
rect 1848 1944 1850 1984
rect 1854 1944 1858 1984
rect 1870 1944 1872 2024
rect 1876 1944 1880 2024
rect 1884 1944 1886 2024
rect 1943 1944 1945 2024
rect 1949 1944 1955 2024
rect 1959 2016 1975 2024
rect 1959 1952 1961 2016
rect 1973 1952 1975 2016
rect 1979 1952 1985 2032
rect 1989 1992 1999 2032
rect 2087 2024 2095 2032
rect 1989 1952 1991 1992
rect 2003 1952 2005 1992
rect 2009 1952 2011 1992
rect 1959 1944 1968 1952
rect 2063 1944 2065 2024
rect 2069 1944 2075 2024
rect 2079 2016 2095 2024
rect 2079 1952 2081 2016
rect 2093 1952 2095 2016
rect 2099 1952 2105 2032
rect 2109 1992 2119 2032
rect 2109 1952 2111 1992
rect 2123 1952 2125 1992
rect 2129 1952 2131 1992
rect 2079 1944 2088 1952
rect 2173 1944 2175 2024
rect 2179 1984 2188 2024
rect 2179 1944 2181 1984
rect 2193 1944 2195 1984
rect 2199 1944 2209 1984
rect 2213 1944 2215 1984
rect 2227 1944 2229 1984
rect 2233 1944 2241 1984
rect 2245 1944 2247 1984
rect 2259 1944 2261 1984
rect 2265 1944 2267 1984
rect 2305 1944 2307 1984
rect 2311 1944 2315 1984
rect 2319 1964 2330 1984
rect 2356 1964 2365 2024
rect 2319 1944 2321 1964
rect 2333 1944 2335 1964
rect 2339 1944 2343 1964
rect 2347 1944 2351 1964
rect 2363 1944 2365 1964
rect 2369 1944 2371 2024
rect 2428 1944 2430 1984
rect 2434 1944 2438 1984
rect 2450 1944 2452 2024
rect 2456 1944 2460 2024
rect 2464 1944 2466 2024
rect 2509 1944 2511 2024
rect 2515 1944 2519 2024
rect 2523 1944 2525 2024
rect 2701 1992 2711 2032
rect 2603 1944 2605 1984
rect 2609 1980 2625 1984
rect 2609 1944 2611 1980
rect 2623 1944 2625 1980
rect 2629 1944 2631 1984
rect 2643 1944 2645 1984
rect 2649 1944 2651 1984
rect 2689 1952 2691 1992
rect 2695 1952 2697 1992
rect 2709 1952 2711 1992
rect 2715 1952 2721 2032
rect 2725 2024 2733 2032
rect 2847 2024 2855 2032
rect 2725 2016 2741 2024
rect 2725 1952 2727 2016
rect 2739 1952 2741 2016
rect 2732 1944 2741 1952
rect 2745 1944 2751 2024
rect 2755 1944 2757 2024
rect 2823 1944 2825 2024
rect 2829 1944 2835 2024
rect 2839 2016 2855 2024
rect 2839 1952 2841 2016
rect 2853 1952 2855 2016
rect 2859 1952 2865 2032
rect 2869 1992 2879 2032
rect 2869 1952 2871 1992
rect 2883 1952 2885 1992
rect 2889 1952 2891 1992
rect 2839 1944 2848 1952
rect 2929 1944 2931 1984
rect 2935 1944 2937 1984
rect 2989 1944 2991 2024
rect 2995 1944 3001 2024
rect 3005 1944 3007 2024
rect 3029 1944 3031 2024
rect 3035 1944 3041 2024
rect 3045 1944 3047 2024
rect 3123 1944 3125 2024
rect 3129 1944 3131 2024
rect 3143 1944 3145 2024
rect 3149 2012 3165 2024
rect 3149 1944 3151 2012
rect 3163 1944 3165 2012
rect 3169 2016 3183 2024
rect 3169 1944 3171 2016
rect 3209 1944 3211 1984
rect 3215 1944 3217 1984
rect 3269 1944 3271 2024
rect 3275 1944 3281 2024
rect 3285 1944 3287 2024
rect 3309 1944 3311 2024
rect 3315 1944 3321 2024
rect 3325 1944 3327 2024
rect 3389 1944 3391 2024
rect 3395 1944 3399 2024
rect 3403 1944 3405 2024
rect 3473 1944 3475 2024
rect 3479 1984 3488 2024
rect 3479 1944 3481 1984
rect 3493 1944 3495 1984
rect 3499 1944 3509 1984
rect 3513 1944 3515 1984
rect 3527 1944 3529 1984
rect 3533 1944 3541 1984
rect 3545 1944 3547 1984
rect 3559 1944 3561 1984
rect 3565 1944 3567 1984
rect 3605 1944 3607 1984
rect 3611 1944 3615 1984
rect 3619 1964 3630 1984
rect 3656 1964 3665 2024
rect 3619 1944 3621 1964
rect 3633 1944 3635 1964
rect 3639 1944 3643 1964
rect 3647 1944 3651 1964
rect 3663 1944 3665 1964
rect 3669 1944 3671 2024
rect 3735 1944 3737 2024
rect 3741 1944 3745 2024
rect 3749 1944 3751 2024
rect 3813 1944 3815 2024
rect 3819 1944 3825 2024
rect 3829 1944 3831 2024
rect 3853 1944 3855 2024
rect 3859 1944 3865 2024
rect 3869 1944 3871 2024
rect 3923 1944 3925 1984
rect 3929 1944 3931 1984
rect 3974 1944 3976 2024
rect 3980 1944 3984 2024
rect 3988 1944 3990 2024
rect 4002 1944 4006 1984
rect 4010 1944 4012 1984
rect 4069 1944 4071 1984
rect 4075 1944 4077 1984
rect 4089 1944 4091 1984
rect 4095 1944 4097 1984
rect 4175 1944 4177 2024
rect 4181 1944 4185 2024
rect 4189 1944 4191 2024
rect 4233 1944 4235 2024
rect 4239 1984 4248 2024
rect 4239 1944 4241 1984
rect 4253 1944 4255 1984
rect 4259 1944 4269 1984
rect 4273 1944 4275 1984
rect 4287 1944 4289 1984
rect 4293 1944 4301 1984
rect 4305 1944 4307 1984
rect 4319 1944 4321 1984
rect 4325 1944 4327 1984
rect 4365 1944 4367 1984
rect 4371 1944 4375 1984
rect 4379 1964 4390 1984
rect 4416 1964 4425 2024
rect 4379 1944 4381 1964
rect 4393 1944 4395 1964
rect 4399 1944 4403 1964
rect 4407 1944 4411 1964
rect 4423 1944 4425 1964
rect 4429 1944 4431 2024
rect 4469 1944 4471 1984
rect 4475 1944 4477 1984
rect 4529 1944 4531 2024
rect 4535 1944 4541 2024
rect 4545 1944 4547 2024
rect 4569 1944 4571 2024
rect 4575 1944 4581 2024
rect 4585 1944 4587 2024
rect 4649 1944 4651 2024
rect 4655 1944 4659 2024
rect 4663 1944 4665 2024
rect 4748 1944 4750 1984
rect 4754 1944 4758 1984
rect 4770 1944 4772 2024
rect 4776 1944 4780 2024
rect 4784 1944 4786 2024
rect 4855 1944 4857 2024
rect 4861 1944 4865 2024
rect 4869 1944 4871 2024
rect 4909 1944 4911 2024
rect 4915 1944 4921 2024
rect 4925 1944 4927 2024
rect 4949 1944 4951 2024
rect 4955 1944 4961 2024
rect 4965 1944 4967 2024
rect 5043 1944 5045 1984
rect 5049 1944 5051 1984
rect 5063 1944 5065 1984
rect 5069 1944 5071 1984
rect 5135 1944 5137 2024
rect 5141 1944 5145 2024
rect 5149 1944 5151 2024
rect 5189 1944 5191 2024
rect 5195 1944 5201 2024
rect 5205 2023 5221 2024
rect 5205 1944 5207 2023
rect 5219 1944 5221 2023
rect 5225 2023 5239 2024
rect 5225 1944 5227 2023
rect 5313 1944 5315 2024
rect 5319 1944 5325 2024
rect 5329 1944 5331 2024
rect 5353 1944 5355 2024
rect 5359 1944 5365 2024
rect 5369 1944 5371 2024
rect 5409 1944 5411 2024
rect 5415 1944 5421 2024
rect 5425 1944 5427 2024
rect 5449 1944 5451 2024
rect 5455 1944 5461 2024
rect 5465 1944 5467 2024
rect 5555 1944 5557 2024
rect 5561 1944 5565 2024
rect 5569 1944 5571 2024
rect 5633 1944 5635 2024
rect 5639 1944 5645 2024
rect 5649 1944 5651 2024
rect 5673 1944 5675 2024
rect 5679 1944 5685 2024
rect 5689 1944 5691 2024
rect 5743 1944 5745 1984
rect 5749 1944 5751 1984
rect 5789 1944 5791 1984
rect 5795 1944 5797 1984
rect 5809 1944 5811 1984
rect 5815 1944 5817 1984
rect 5869 1944 5871 2024
rect 5875 1964 5884 2024
rect 6052 1984 6061 2024
rect 5910 1964 5921 1984
rect 5875 1944 5877 1964
rect 5889 1944 5893 1964
rect 5897 1944 5901 1964
rect 5905 1944 5907 1964
rect 5919 1944 5921 1964
rect 5925 1944 5929 1984
rect 5933 1944 5935 1984
rect 5973 1944 5975 1984
rect 5979 1944 5981 1984
rect 5993 1944 5995 1984
rect 5999 1944 6007 1984
rect 6011 1944 6013 1984
rect 6025 1944 6027 1984
rect 6031 1944 6041 1984
rect 6045 1944 6047 1984
rect 6059 1944 6061 1984
rect 6065 1944 6067 2024
rect 6113 1944 6115 2024
rect 6119 1984 6128 2024
rect 6119 1944 6121 1984
rect 6133 1944 6135 1984
rect 6139 1944 6149 1984
rect 6153 1944 6155 1984
rect 6167 1944 6169 1984
rect 6173 1944 6181 1984
rect 6185 1944 6187 1984
rect 6199 1944 6201 1984
rect 6205 1944 6207 1984
rect 6245 1944 6247 1984
rect 6251 1944 6255 1984
rect 6259 1964 6270 1984
rect 6296 1964 6305 2024
rect 6259 1944 6261 1964
rect 6273 1944 6275 1964
rect 6279 1944 6283 1964
rect 6287 1944 6291 1964
rect 6303 1944 6305 1964
rect 6309 1944 6311 2024
rect 6361 1992 6371 2032
rect 6349 1952 6351 1992
rect 6355 1952 6357 1992
rect 6369 1952 6371 1992
rect 6375 1952 6381 2032
rect 6385 2024 6393 2032
rect 6385 2016 6401 2024
rect 6385 1952 6387 2016
rect 6399 1952 6401 2016
rect 6392 1944 6401 1952
rect 6405 1944 6411 2024
rect 6415 1944 6417 2024
rect 6457 2016 6471 2024
rect 6469 1944 6471 2016
rect 6475 2012 6491 2024
rect 6475 1944 6477 2012
rect 6489 1944 6491 2012
rect 6495 1944 6497 2024
rect 6509 1944 6511 2024
rect 6515 1944 6517 2024
rect 6574 1944 6576 2024
rect 6580 1944 6584 2024
rect 6588 1944 6590 2024
rect 6602 1944 6606 1984
rect 6610 1944 6612 1984
rect 43 1876 45 1916
rect 49 1876 51 1916
rect 89 1836 91 1916
rect 95 1896 97 1916
rect 109 1896 113 1916
rect 117 1896 121 1916
rect 125 1896 127 1916
rect 139 1896 141 1916
rect 95 1836 104 1896
rect 130 1876 141 1896
rect 145 1876 149 1916
rect 153 1876 155 1916
rect 193 1876 195 1916
rect 199 1876 201 1916
rect 213 1876 215 1916
rect 219 1876 227 1916
rect 231 1876 233 1916
rect 245 1876 247 1916
rect 251 1876 261 1916
rect 265 1876 267 1916
rect 279 1876 281 1916
rect 272 1836 281 1876
rect 285 1836 287 1916
rect 329 1836 331 1916
rect 335 1836 339 1916
rect 343 1836 345 1916
rect 435 1836 437 1916
rect 441 1836 445 1916
rect 449 1836 451 1916
rect 503 1876 505 1916
rect 509 1876 511 1916
rect 568 1876 570 1916
rect 574 1876 578 1916
rect 590 1836 592 1916
rect 596 1836 600 1916
rect 604 1836 606 1916
rect 649 1836 651 1916
rect 655 1896 657 1916
rect 669 1896 673 1916
rect 677 1896 681 1916
rect 685 1896 687 1916
rect 699 1896 701 1916
rect 655 1836 664 1896
rect 690 1876 701 1896
rect 705 1876 709 1916
rect 713 1876 715 1916
rect 753 1876 755 1916
rect 759 1876 761 1916
rect 773 1876 775 1916
rect 779 1876 787 1916
rect 791 1876 793 1916
rect 805 1876 807 1916
rect 811 1876 821 1916
rect 825 1876 827 1916
rect 839 1876 841 1916
rect 832 1836 841 1876
rect 845 1836 847 1916
rect 903 1876 905 1916
rect 909 1880 911 1916
rect 923 1880 925 1916
rect 909 1876 925 1880
rect 929 1876 931 1916
rect 943 1876 945 1916
rect 949 1876 951 1916
rect 989 1876 991 1916
rect 995 1876 997 1916
rect 1009 1876 1013 1916
rect 1017 1876 1021 1916
rect 1033 1836 1035 1916
rect 1039 1836 1041 1916
rect 1089 1876 1091 1916
rect 1095 1876 1097 1916
rect 1154 1836 1156 1916
rect 1160 1836 1164 1916
rect 1168 1836 1170 1916
rect 1182 1876 1186 1916
rect 1190 1876 1192 1916
rect 1263 1876 1265 1916
rect 1269 1876 1271 1916
rect 1283 1876 1285 1916
rect 1289 1876 1291 1916
rect 1343 1876 1345 1916
rect 1349 1880 1351 1916
rect 1363 1880 1365 1916
rect 1349 1876 1365 1880
rect 1369 1876 1371 1916
rect 1383 1876 1385 1916
rect 1389 1876 1391 1916
rect 1429 1876 1431 1916
rect 1435 1876 1437 1916
rect 1493 1836 1495 1916
rect 1499 1876 1501 1916
rect 1513 1876 1515 1916
rect 1519 1876 1529 1916
rect 1533 1876 1535 1916
rect 1547 1876 1549 1916
rect 1553 1876 1561 1916
rect 1565 1876 1567 1916
rect 1579 1876 1581 1916
rect 1585 1876 1587 1916
rect 1625 1876 1627 1916
rect 1631 1876 1635 1916
rect 1639 1896 1641 1916
rect 1653 1896 1655 1916
rect 1659 1896 1663 1916
rect 1667 1896 1671 1916
rect 1683 1896 1685 1916
rect 1639 1876 1650 1896
rect 1499 1836 1508 1876
rect 1676 1836 1685 1896
rect 1689 1836 1691 1916
rect 1729 1876 1731 1916
rect 1735 1876 1737 1916
rect 1789 1836 1791 1916
rect 1795 1836 1801 1916
rect 1805 1836 1807 1916
rect 1829 1836 1831 1916
rect 1835 1836 1841 1916
rect 1845 1836 1847 1916
rect 1909 1836 1911 1916
rect 1915 1836 1919 1916
rect 1923 1836 1925 1916
rect 1994 1836 1996 1916
rect 2000 1836 2004 1916
rect 2008 1836 2010 1916
rect 2022 1876 2026 1916
rect 2030 1876 2032 1916
rect 2089 1836 2091 1916
rect 2095 1896 2097 1916
rect 2109 1896 2113 1916
rect 2117 1896 2121 1916
rect 2125 1896 2127 1916
rect 2139 1896 2141 1916
rect 2095 1836 2104 1896
rect 2130 1876 2141 1896
rect 2145 1876 2149 1916
rect 2153 1876 2155 1916
rect 2193 1876 2195 1916
rect 2199 1876 2201 1916
rect 2213 1876 2215 1916
rect 2219 1876 2227 1916
rect 2231 1876 2233 1916
rect 2245 1876 2247 1916
rect 2251 1876 2261 1916
rect 2265 1876 2267 1916
rect 2279 1876 2281 1916
rect 2272 1836 2281 1876
rect 2285 1836 2287 1916
rect 2353 1836 2355 1916
rect 2359 1836 2365 1916
rect 2369 1836 2371 1916
rect 2393 1836 2395 1916
rect 2399 1836 2405 1916
rect 2409 1836 2411 1916
rect 2449 1876 2451 1916
rect 2455 1876 2457 1916
rect 2509 1836 2511 1916
rect 2515 1836 2519 1916
rect 2523 1836 2525 1916
rect 2589 1836 2591 1916
rect 2595 1896 2597 1916
rect 2609 1896 2613 1916
rect 2617 1896 2621 1916
rect 2625 1896 2627 1916
rect 2639 1896 2641 1916
rect 2595 1836 2604 1896
rect 2630 1876 2641 1896
rect 2645 1876 2649 1916
rect 2653 1876 2655 1916
rect 2693 1876 2695 1916
rect 2699 1876 2701 1916
rect 2713 1876 2715 1916
rect 2719 1876 2727 1916
rect 2731 1876 2733 1916
rect 2745 1876 2747 1916
rect 2751 1876 2761 1916
rect 2765 1876 2767 1916
rect 2779 1876 2781 1916
rect 2772 1836 2781 1876
rect 2785 1836 2787 1916
rect 2829 1876 2831 1916
rect 2835 1876 2837 1916
rect 2849 1876 2851 1916
rect 2855 1880 2857 1916
rect 2869 1880 2871 1916
rect 2855 1876 2871 1880
rect 2875 1876 2877 1916
rect 2948 1876 2950 1916
rect 2954 1876 2958 1916
rect 2970 1836 2972 1916
rect 2976 1836 2980 1916
rect 2984 1836 2986 1916
rect 3029 1836 3031 1916
rect 3035 1836 3039 1916
rect 3043 1836 3045 1916
rect 3123 1836 3125 1916
rect 3129 1836 3131 1916
rect 3143 1836 3145 1916
rect 3149 1848 3151 1916
rect 3163 1848 3165 1916
rect 3149 1836 3165 1848
rect 3169 1844 3171 1916
rect 3169 1836 3183 1844
rect 3223 1836 3225 1916
rect 3229 1836 3231 1916
rect 3243 1836 3245 1916
rect 3249 1848 3251 1916
rect 3263 1848 3265 1916
rect 3249 1836 3265 1848
rect 3269 1844 3271 1916
rect 3269 1836 3283 1844
rect 3321 1836 3323 1916
rect 3327 1836 3329 1916
rect 3341 1876 3345 1916
rect 3349 1876 3351 1916
rect 3403 1876 3405 1916
rect 3409 1876 3411 1916
rect 3423 1876 3425 1916
rect 3429 1876 3431 1916
rect 3469 1836 3471 1916
rect 3475 1836 3479 1916
rect 3483 1836 3485 1916
rect 3549 1876 3551 1916
rect 3555 1876 3557 1916
rect 3569 1876 3571 1916
rect 3575 1876 3577 1916
rect 3634 1836 3636 1916
rect 3640 1836 3644 1916
rect 3648 1836 3650 1916
rect 3662 1876 3666 1916
rect 3670 1876 3672 1916
rect 3743 1876 3745 1916
rect 3749 1876 3751 1916
rect 3763 1876 3765 1916
rect 3769 1876 3771 1916
rect 3823 1876 3825 1916
rect 3829 1876 3831 1916
rect 3869 1876 3871 1916
rect 3875 1876 3877 1916
rect 3889 1876 3891 1916
rect 3895 1876 3897 1916
rect 3949 1836 3951 1916
rect 3955 1836 3959 1916
rect 3963 1836 3965 1916
rect 4029 1836 4031 1916
rect 4035 1836 4041 1916
rect 4045 1836 4047 1916
rect 4069 1836 4071 1916
rect 4075 1836 4081 1916
rect 4085 1836 4087 1916
rect 4175 1836 4177 1916
rect 4181 1836 4185 1916
rect 4189 1836 4191 1916
rect 4234 1836 4236 1916
rect 4240 1836 4244 1916
rect 4248 1836 4250 1916
rect 4262 1876 4266 1916
rect 4270 1876 4272 1916
rect 4317 1914 4331 1916
rect 4329 1836 4331 1914
rect 4335 1836 4337 1916
rect 4349 1836 4351 1916
rect 4355 1836 4357 1916
rect 4414 1836 4416 1916
rect 4420 1836 4424 1916
rect 4428 1836 4430 1916
rect 4442 1876 4446 1916
rect 4450 1876 4452 1916
rect 4535 1836 4537 1916
rect 4541 1836 4545 1916
rect 4549 1836 4551 1916
rect 4613 1836 4615 1916
rect 4619 1836 4625 1916
rect 4629 1836 4631 1916
rect 4653 1836 4655 1916
rect 4659 1836 4665 1916
rect 4669 1836 4671 1916
rect 4723 1876 4725 1916
rect 4729 1876 4731 1916
rect 4769 1836 4771 1916
rect 4775 1896 4777 1916
rect 4789 1896 4793 1916
rect 4797 1896 4801 1916
rect 4805 1896 4807 1916
rect 4819 1896 4821 1916
rect 4775 1836 4784 1896
rect 4810 1876 4821 1896
rect 4825 1876 4829 1916
rect 4833 1876 4835 1916
rect 4873 1876 4875 1916
rect 4879 1876 4881 1916
rect 4893 1876 4895 1916
rect 4899 1876 4907 1916
rect 4911 1876 4913 1916
rect 4925 1876 4927 1916
rect 4931 1876 4941 1916
rect 4945 1876 4947 1916
rect 4959 1876 4961 1916
rect 4952 1836 4961 1876
rect 4965 1836 4967 1916
rect 5009 1844 5011 1916
rect 4997 1836 5011 1844
rect 5015 1848 5017 1916
rect 5029 1848 5031 1916
rect 5015 1836 5031 1848
rect 5035 1836 5037 1916
rect 5049 1836 5051 1916
rect 5055 1836 5057 1916
rect 5109 1836 5111 1916
rect 5115 1836 5119 1916
rect 5123 1836 5125 1916
rect 5194 1836 5196 1916
rect 5200 1836 5204 1916
rect 5208 1836 5210 1916
rect 5222 1876 5226 1916
rect 5230 1876 5232 1916
rect 5289 1876 5291 1916
rect 5295 1876 5297 1916
rect 5309 1876 5311 1916
rect 5315 1880 5317 1916
rect 5329 1880 5331 1916
rect 5315 1876 5331 1880
rect 5335 1876 5337 1916
rect 5389 1876 5391 1916
rect 5395 1876 5399 1916
rect 5411 1836 5413 1916
rect 5417 1836 5419 1916
rect 5483 1876 5485 1916
rect 5489 1876 5491 1916
rect 5543 1836 5545 1916
rect 5549 1836 5551 1916
rect 5608 1876 5610 1916
rect 5614 1876 5618 1916
rect 5630 1836 5632 1916
rect 5636 1836 5640 1916
rect 5644 1836 5646 1916
rect 5689 1876 5691 1916
rect 5695 1876 5697 1916
rect 5709 1876 5711 1916
rect 5715 1876 5717 1916
rect 5783 1836 5785 1916
rect 5789 1904 5805 1916
rect 5789 1836 5791 1904
rect 5803 1836 5805 1904
rect 5809 1838 5811 1916
rect 5823 1838 5825 1916
rect 5809 1836 5825 1838
rect 5829 1850 5831 1916
rect 5843 1850 5845 1916
rect 5829 1836 5845 1850
rect 5849 1838 5851 1916
rect 5889 1876 5891 1916
rect 5895 1876 5899 1916
rect 5849 1836 5863 1838
rect 5911 1836 5913 1916
rect 5917 1836 5919 1916
rect 5988 1876 5990 1916
rect 5994 1876 5998 1916
rect 6010 1836 6012 1916
rect 6016 1836 6020 1916
rect 6024 1836 6026 1916
rect 6093 1836 6095 1916
rect 6099 1836 6105 1916
rect 6109 1836 6111 1916
rect 6133 1836 6135 1916
rect 6139 1836 6145 1916
rect 6149 1836 6151 1916
rect 6232 1908 6241 1916
rect 6189 1868 6191 1908
rect 6195 1868 6197 1908
rect 6209 1868 6211 1908
rect 6201 1828 6211 1868
rect 6215 1828 6221 1908
rect 6225 1844 6227 1908
rect 6239 1844 6241 1908
rect 6225 1836 6241 1844
rect 6245 1836 6251 1916
rect 6255 1836 6257 1916
rect 6352 1908 6361 1916
rect 6309 1868 6311 1908
rect 6315 1868 6317 1908
rect 6329 1868 6331 1908
rect 6225 1828 6233 1836
rect 6321 1828 6331 1868
rect 6335 1828 6341 1908
rect 6345 1844 6347 1908
rect 6359 1844 6361 1908
rect 6345 1836 6361 1844
rect 6365 1836 6371 1916
rect 6375 1836 6377 1916
rect 6429 1876 6431 1916
rect 6435 1876 6437 1916
rect 6345 1828 6353 1836
rect 6494 1836 6496 1916
rect 6500 1836 6504 1916
rect 6508 1836 6510 1916
rect 6522 1876 6526 1916
rect 6530 1876 6532 1916
rect 6603 1876 6605 1916
rect 6609 1876 6611 1916
rect 6623 1876 6625 1916
rect 6629 1876 6631 1916
rect 55 1464 57 1544
rect 61 1464 65 1544
rect 69 1464 71 1544
rect 123 1464 125 1544
rect 129 1464 131 1544
rect 143 1464 145 1544
rect 149 1464 151 1544
rect 163 1464 165 1544
rect 169 1464 171 1544
rect 183 1464 185 1544
rect 189 1464 191 1544
rect 203 1464 205 1544
rect 209 1464 211 1544
rect 223 1464 225 1544
rect 229 1464 231 1544
rect 243 1464 245 1544
rect 249 1464 251 1544
rect 263 1464 265 1544
rect 269 1464 271 1544
rect 313 1464 315 1544
rect 319 1504 328 1544
rect 319 1464 321 1504
rect 333 1464 335 1504
rect 339 1464 349 1504
rect 353 1464 355 1504
rect 367 1464 369 1504
rect 373 1464 381 1504
rect 385 1464 387 1504
rect 399 1464 401 1504
rect 405 1464 407 1504
rect 445 1464 447 1504
rect 451 1464 455 1504
rect 459 1484 470 1504
rect 496 1484 505 1544
rect 459 1464 461 1484
rect 473 1464 475 1484
rect 479 1464 483 1484
rect 487 1464 491 1484
rect 503 1464 505 1484
rect 509 1464 511 1544
rect 697 1536 711 1544
rect 563 1464 565 1504
rect 569 1464 571 1504
rect 609 1464 611 1504
rect 615 1464 617 1504
rect 629 1464 631 1504
rect 635 1500 651 1504
rect 635 1464 637 1500
rect 649 1464 651 1500
rect 655 1464 657 1504
rect 709 1464 711 1536
rect 715 1532 731 1544
rect 715 1464 717 1532
rect 729 1464 731 1532
rect 735 1464 737 1544
rect 749 1464 751 1544
rect 755 1464 757 1544
rect 813 1464 815 1544
rect 819 1504 828 1544
rect 819 1464 821 1504
rect 833 1464 835 1504
rect 839 1464 849 1504
rect 853 1464 855 1504
rect 867 1464 869 1504
rect 873 1464 881 1504
rect 885 1464 887 1504
rect 899 1464 901 1504
rect 905 1464 907 1504
rect 945 1464 947 1504
rect 951 1464 955 1504
rect 959 1484 970 1504
rect 996 1484 1005 1544
rect 959 1464 961 1484
rect 973 1464 975 1484
rect 979 1464 983 1484
rect 987 1464 991 1484
rect 1003 1464 1005 1484
rect 1009 1464 1011 1544
rect 1063 1464 1065 1504
rect 1069 1464 1071 1504
rect 1109 1464 1111 1544
rect 1115 1464 1121 1544
rect 1125 1464 1127 1544
rect 1149 1464 1151 1544
rect 1155 1464 1161 1544
rect 1165 1464 1167 1544
rect 1447 1544 1455 1552
rect 1248 1464 1250 1504
rect 1254 1464 1258 1504
rect 1270 1464 1272 1544
rect 1276 1464 1280 1544
rect 1284 1464 1286 1544
rect 1355 1464 1357 1544
rect 1361 1464 1365 1544
rect 1369 1464 1371 1544
rect 1423 1464 1425 1544
rect 1429 1464 1435 1544
rect 1439 1536 1455 1544
rect 1439 1472 1441 1536
rect 1453 1472 1455 1536
rect 1459 1472 1465 1552
rect 1469 1512 1479 1552
rect 1567 1544 1575 1552
rect 1469 1472 1471 1512
rect 1483 1472 1485 1512
rect 1489 1472 1491 1512
rect 1439 1464 1448 1472
rect 1543 1464 1545 1544
rect 1549 1464 1555 1544
rect 1559 1536 1575 1544
rect 1559 1472 1561 1536
rect 1573 1472 1575 1536
rect 1579 1472 1585 1552
rect 1589 1512 1599 1552
rect 1687 1544 1695 1552
rect 1589 1472 1591 1512
rect 1603 1472 1605 1512
rect 1609 1472 1611 1512
rect 1559 1464 1568 1472
rect 1663 1464 1665 1544
rect 1669 1464 1675 1544
rect 1679 1536 1695 1544
rect 1679 1472 1681 1536
rect 1693 1472 1695 1536
rect 1699 1472 1705 1552
rect 1709 1512 1719 1552
rect 1709 1472 1711 1512
rect 1723 1472 1725 1512
rect 1729 1472 1731 1512
rect 1679 1464 1688 1472
rect 1769 1464 1771 1544
rect 1775 1484 1784 1544
rect 1952 1504 1961 1544
rect 1810 1484 1821 1504
rect 1775 1464 1777 1484
rect 1789 1464 1793 1484
rect 1797 1464 1801 1484
rect 1805 1464 1807 1484
rect 1819 1464 1821 1484
rect 1825 1464 1829 1504
rect 1833 1464 1835 1504
rect 1873 1464 1875 1504
rect 1879 1464 1881 1504
rect 1893 1464 1895 1504
rect 1899 1464 1907 1504
rect 1911 1464 1913 1504
rect 1925 1464 1927 1504
rect 1931 1464 1941 1504
rect 1945 1464 1947 1504
rect 1959 1464 1961 1504
rect 1965 1464 1967 1544
rect 2021 1512 2031 1552
rect 2009 1472 2011 1512
rect 2015 1472 2017 1512
rect 2029 1472 2031 1512
rect 2035 1472 2041 1552
rect 2045 1544 2053 1552
rect 2045 1536 2061 1544
rect 2045 1472 2047 1536
rect 2059 1472 2061 1536
rect 2052 1464 2061 1472
rect 2065 1464 2071 1544
rect 2075 1464 2077 1544
rect 2129 1464 2131 1504
rect 2135 1464 2137 1504
rect 2189 1464 2191 1544
rect 2195 1464 2201 1544
rect 2205 1464 2207 1544
rect 2229 1464 2231 1544
rect 2235 1464 2241 1544
rect 2245 1464 2247 1544
rect 2309 1464 2311 1544
rect 2315 1464 2319 1544
rect 2323 1464 2325 1544
rect 2408 1464 2410 1504
rect 2414 1464 2418 1504
rect 2430 1464 2432 1544
rect 2436 1464 2440 1544
rect 2444 1464 2446 1544
rect 2501 1464 2503 1544
rect 2507 1464 2509 1544
rect 2521 1464 2525 1504
rect 2529 1464 2531 1504
rect 2569 1464 2571 1544
rect 2575 1464 2579 1544
rect 2583 1464 2585 1544
rect 2847 1544 2855 1552
rect 2663 1464 2665 1504
rect 2669 1464 2671 1504
rect 2683 1464 2685 1504
rect 2689 1464 2691 1504
rect 2729 1464 2731 1504
rect 2735 1464 2737 1504
rect 2749 1464 2751 1504
rect 2755 1464 2757 1504
rect 2823 1464 2825 1544
rect 2829 1464 2835 1544
rect 2839 1536 2855 1544
rect 2839 1472 2841 1536
rect 2853 1472 2855 1536
rect 2859 1472 2865 1552
rect 2869 1512 2879 1552
rect 2869 1472 2871 1512
rect 2883 1472 2885 1512
rect 2889 1472 2891 1512
rect 2839 1464 2848 1472
rect 2943 1464 2945 1504
rect 2949 1500 2965 1504
rect 2949 1464 2951 1500
rect 2963 1464 2965 1500
rect 2969 1464 2971 1504
rect 2983 1464 2985 1504
rect 2989 1464 2991 1504
rect 3043 1464 3045 1544
rect 3049 1464 3051 1544
rect 3093 1464 3095 1544
rect 3099 1504 3108 1544
rect 3099 1464 3101 1504
rect 3113 1464 3115 1504
rect 3119 1464 3129 1504
rect 3133 1464 3135 1504
rect 3147 1464 3149 1504
rect 3153 1464 3161 1504
rect 3165 1464 3167 1504
rect 3179 1464 3181 1504
rect 3185 1464 3187 1504
rect 3225 1464 3227 1504
rect 3231 1464 3235 1504
rect 3239 1484 3250 1504
rect 3276 1484 3285 1544
rect 3239 1464 3241 1484
rect 3253 1464 3255 1484
rect 3259 1464 3263 1484
rect 3267 1464 3271 1484
rect 3283 1464 3285 1484
rect 3289 1464 3291 1544
rect 3343 1464 3345 1504
rect 3349 1464 3351 1504
rect 3363 1464 3365 1504
rect 3369 1464 3371 1504
rect 3428 1464 3430 1504
rect 3434 1464 3438 1504
rect 3450 1464 3452 1544
rect 3456 1464 3460 1544
rect 3464 1464 3466 1544
rect 3497 1542 3511 1544
rect 3509 1464 3511 1542
rect 3515 1530 3531 1544
rect 3515 1464 3517 1530
rect 3529 1464 3531 1530
rect 3535 1542 3551 1544
rect 3535 1464 3537 1542
rect 3549 1464 3551 1542
rect 3555 1476 3557 1544
rect 3569 1476 3571 1544
rect 3555 1464 3571 1476
rect 3575 1464 3577 1544
rect 3648 1464 3650 1504
rect 3654 1464 3658 1504
rect 3670 1464 3672 1544
rect 3676 1464 3680 1544
rect 3684 1464 3686 1544
rect 3743 1464 3745 1504
rect 3749 1464 3751 1504
rect 3815 1464 3817 1544
rect 3821 1464 3825 1544
rect 3829 1464 3831 1544
rect 3893 1464 3895 1544
rect 3899 1464 3905 1544
rect 3909 1464 3911 1544
rect 3933 1464 3935 1544
rect 3939 1464 3945 1544
rect 3949 1464 3951 1544
rect 4003 1464 4005 1504
rect 4009 1464 4011 1504
rect 4053 1464 4055 1544
rect 4059 1504 4068 1544
rect 4327 1544 4335 1552
rect 4059 1464 4061 1504
rect 4073 1464 4075 1504
rect 4079 1464 4089 1504
rect 4093 1464 4095 1504
rect 4107 1464 4109 1504
rect 4113 1464 4121 1504
rect 4125 1464 4127 1504
rect 4139 1464 4141 1504
rect 4145 1464 4147 1504
rect 4185 1464 4187 1504
rect 4191 1464 4195 1504
rect 4199 1484 4210 1504
rect 4236 1484 4245 1544
rect 4199 1464 4201 1484
rect 4213 1464 4215 1484
rect 4219 1464 4223 1484
rect 4227 1464 4231 1484
rect 4243 1464 4245 1484
rect 4249 1464 4251 1544
rect 4303 1464 4305 1544
rect 4309 1464 4315 1544
rect 4319 1536 4335 1544
rect 4319 1472 4321 1536
rect 4333 1472 4335 1536
rect 4339 1472 4345 1552
rect 4349 1512 4359 1552
rect 4447 1544 4455 1552
rect 4349 1472 4351 1512
rect 4363 1472 4365 1512
rect 4369 1472 4371 1512
rect 4319 1464 4328 1472
rect 4423 1464 4425 1544
rect 4429 1464 4435 1544
rect 4439 1536 4455 1544
rect 4439 1472 4441 1536
rect 4453 1472 4455 1536
rect 4459 1472 4465 1552
rect 4469 1512 4479 1552
rect 4541 1512 4551 1552
rect 4469 1472 4471 1512
rect 4483 1472 4485 1512
rect 4489 1472 4491 1512
rect 4529 1472 4531 1512
rect 4535 1472 4537 1512
rect 4549 1472 4551 1512
rect 4555 1472 4561 1552
rect 4565 1544 4573 1552
rect 4565 1536 4581 1544
rect 4565 1472 4567 1536
rect 4579 1472 4581 1536
rect 4439 1464 4448 1472
rect 4572 1464 4581 1472
rect 4585 1464 4591 1544
rect 4595 1464 4597 1544
rect 4661 1512 4671 1552
rect 4649 1472 4651 1512
rect 4655 1472 4657 1512
rect 4669 1472 4671 1512
rect 4675 1472 4681 1552
rect 4685 1544 4693 1552
rect 4685 1536 4701 1544
rect 4685 1472 4687 1536
rect 4699 1472 4701 1536
rect 4692 1464 4701 1472
rect 4705 1464 4711 1544
rect 4715 1464 4717 1544
rect 4781 1512 4791 1552
rect 4769 1472 4771 1512
rect 4775 1472 4777 1512
rect 4789 1472 4791 1512
rect 4795 1472 4801 1552
rect 4805 1544 4813 1552
rect 4805 1536 4821 1544
rect 4805 1472 4807 1536
rect 4819 1472 4821 1536
rect 4812 1464 4821 1472
rect 4825 1464 4831 1544
rect 4835 1464 4837 1544
rect 4901 1512 4911 1552
rect 4889 1472 4891 1512
rect 4895 1472 4897 1512
rect 4909 1472 4911 1512
rect 4915 1472 4921 1552
rect 4925 1544 4933 1552
rect 4925 1536 4941 1544
rect 4925 1472 4927 1536
rect 4939 1472 4941 1536
rect 4932 1464 4941 1472
rect 4945 1464 4951 1544
rect 4955 1464 4957 1544
rect 5009 1464 5011 1544
rect 5015 1484 5024 1544
rect 5192 1504 5201 1544
rect 5050 1484 5061 1504
rect 5015 1464 5017 1484
rect 5029 1464 5033 1484
rect 5037 1464 5041 1484
rect 5045 1464 5047 1484
rect 5059 1464 5061 1484
rect 5065 1464 5069 1504
rect 5073 1464 5075 1504
rect 5113 1464 5115 1504
rect 5119 1464 5121 1504
rect 5133 1464 5135 1504
rect 5139 1464 5147 1504
rect 5151 1464 5153 1504
rect 5165 1464 5167 1504
rect 5171 1464 5181 1504
rect 5185 1464 5187 1504
rect 5199 1464 5201 1504
rect 5205 1464 5207 1544
rect 5249 1464 5251 1544
rect 5255 1484 5264 1544
rect 5432 1504 5441 1544
rect 5290 1484 5301 1504
rect 5255 1464 5257 1484
rect 5269 1464 5273 1484
rect 5277 1464 5281 1484
rect 5285 1464 5287 1484
rect 5299 1464 5301 1484
rect 5305 1464 5309 1504
rect 5313 1464 5315 1504
rect 5353 1464 5355 1504
rect 5359 1464 5361 1504
rect 5373 1464 5375 1504
rect 5379 1464 5387 1504
rect 5391 1464 5393 1504
rect 5405 1464 5407 1504
rect 5411 1464 5421 1504
rect 5425 1464 5427 1504
rect 5439 1464 5441 1504
rect 5445 1464 5447 1544
rect 5477 1542 5491 1544
rect 5489 1464 5491 1542
rect 5495 1530 5511 1544
rect 5495 1464 5497 1530
rect 5509 1464 5511 1530
rect 5515 1542 5531 1544
rect 5515 1464 5517 1542
rect 5529 1464 5531 1542
rect 5535 1476 5537 1544
rect 5549 1476 5551 1544
rect 5535 1464 5551 1476
rect 5555 1464 5557 1544
rect 5621 1512 5631 1552
rect 5609 1472 5611 1512
rect 5615 1472 5617 1512
rect 5629 1472 5631 1512
rect 5635 1472 5641 1552
rect 5645 1544 5653 1552
rect 5645 1536 5661 1544
rect 5645 1472 5647 1536
rect 5659 1472 5661 1536
rect 5652 1464 5661 1472
rect 5665 1464 5671 1544
rect 5675 1464 5677 1544
rect 5748 1464 5750 1504
rect 5754 1464 5758 1504
rect 5770 1464 5772 1544
rect 5776 1464 5780 1544
rect 5784 1464 5786 1544
rect 5855 1464 5857 1544
rect 5861 1464 5865 1544
rect 5869 1464 5871 1544
rect 6327 1544 6335 1552
rect 5923 1464 5925 1504
rect 5929 1464 5931 1504
rect 5943 1464 5945 1504
rect 5949 1464 5951 1504
rect 6008 1464 6010 1504
rect 6014 1464 6018 1504
rect 6030 1464 6032 1544
rect 6036 1464 6040 1544
rect 6044 1464 6046 1544
rect 6115 1464 6117 1544
rect 6121 1464 6125 1544
rect 6129 1464 6131 1544
rect 6193 1464 6195 1544
rect 6199 1464 6205 1544
rect 6209 1464 6211 1544
rect 6233 1464 6235 1544
rect 6239 1464 6245 1544
rect 6249 1464 6251 1544
rect 6303 1464 6305 1544
rect 6309 1464 6315 1544
rect 6319 1536 6335 1544
rect 6319 1472 6321 1536
rect 6333 1472 6335 1536
rect 6339 1472 6345 1552
rect 6349 1512 6359 1552
rect 6349 1472 6351 1512
rect 6363 1472 6365 1512
rect 6369 1472 6371 1512
rect 6319 1464 6328 1472
rect 6409 1464 6411 1504
rect 6415 1464 6417 1504
rect 6469 1464 6471 1544
rect 6475 1484 6484 1544
rect 6652 1504 6661 1544
rect 6510 1484 6521 1504
rect 6475 1464 6477 1484
rect 6489 1464 6493 1484
rect 6497 1464 6501 1484
rect 6505 1464 6507 1484
rect 6519 1464 6521 1484
rect 6525 1464 6529 1504
rect 6533 1464 6535 1504
rect 6573 1464 6575 1504
rect 6579 1464 6581 1504
rect 6593 1464 6595 1504
rect 6599 1464 6607 1504
rect 6611 1464 6613 1504
rect 6625 1464 6627 1504
rect 6631 1464 6641 1504
rect 6645 1464 6647 1504
rect 6659 1464 6661 1504
rect 6665 1464 6667 1544
rect 29 1396 31 1436
rect 35 1396 37 1436
rect 49 1396 53 1436
rect 57 1396 61 1436
rect 73 1356 75 1436
rect 79 1356 81 1436
rect 129 1356 131 1436
rect 135 1356 139 1436
rect 143 1356 145 1436
rect 228 1396 230 1436
rect 234 1396 238 1436
rect 250 1356 252 1436
rect 256 1356 260 1436
rect 264 1356 266 1436
rect 335 1356 337 1436
rect 341 1356 345 1436
rect 349 1356 351 1436
rect 389 1396 391 1436
rect 395 1396 397 1436
rect 449 1396 451 1436
rect 455 1396 457 1436
rect 523 1396 525 1436
rect 529 1396 531 1436
rect 543 1396 545 1436
rect 549 1396 551 1436
rect 589 1364 591 1436
rect 577 1356 591 1364
rect 595 1368 597 1436
rect 609 1368 611 1436
rect 595 1356 611 1368
rect 615 1356 617 1436
rect 629 1356 631 1436
rect 635 1356 637 1436
rect 693 1356 695 1436
rect 699 1396 701 1436
rect 713 1396 715 1436
rect 719 1396 729 1436
rect 733 1396 735 1436
rect 747 1396 749 1436
rect 753 1396 761 1436
rect 765 1396 767 1436
rect 779 1396 781 1436
rect 785 1396 787 1436
rect 825 1396 827 1436
rect 831 1396 835 1436
rect 839 1416 841 1436
rect 853 1416 855 1436
rect 859 1416 863 1436
rect 867 1416 871 1436
rect 883 1416 885 1436
rect 839 1396 850 1416
rect 699 1356 708 1396
rect 876 1356 885 1416
rect 889 1356 891 1436
rect 943 1396 945 1436
rect 949 1396 951 1436
rect 963 1396 965 1436
rect 969 1396 971 1436
rect 1009 1396 1011 1436
rect 1015 1396 1017 1436
rect 1029 1396 1031 1436
rect 1035 1400 1037 1436
rect 1049 1400 1051 1436
rect 1035 1396 1051 1400
rect 1055 1396 1057 1436
rect 1109 1356 1111 1436
rect 1115 1356 1119 1436
rect 1123 1356 1125 1436
rect 1193 1356 1195 1436
rect 1199 1396 1201 1436
rect 1213 1396 1215 1436
rect 1219 1396 1229 1436
rect 1233 1396 1235 1436
rect 1247 1396 1249 1436
rect 1253 1396 1261 1436
rect 1265 1396 1267 1436
rect 1279 1396 1281 1436
rect 1285 1396 1287 1436
rect 1325 1396 1327 1436
rect 1331 1396 1335 1436
rect 1339 1416 1341 1436
rect 1353 1416 1355 1436
rect 1359 1416 1363 1436
rect 1367 1416 1371 1436
rect 1383 1416 1385 1436
rect 1339 1396 1350 1416
rect 1199 1356 1208 1396
rect 1376 1356 1385 1416
rect 1389 1356 1391 1436
rect 1443 1356 1445 1436
rect 1449 1356 1451 1436
rect 1463 1356 1465 1436
rect 1469 1356 1471 1436
rect 1483 1356 1485 1436
rect 1489 1356 1491 1436
rect 1503 1356 1505 1436
rect 1509 1356 1511 1436
rect 1523 1356 1525 1436
rect 1529 1356 1531 1436
rect 1543 1356 1545 1436
rect 1549 1356 1551 1436
rect 1563 1356 1565 1436
rect 1569 1356 1571 1436
rect 1583 1356 1585 1436
rect 1589 1356 1591 1436
rect 1643 1356 1645 1436
rect 1649 1356 1655 1436
rect 1659 1428 1668 1436
rect 1659 1364 1661 1428
rect 1673 1364 1675 1428
rect 1659 1356 1675 1364
rect 1667 1348 1675 1356
rect 1679 1348 1685 1428
rect 1689 1388 1691 1428
rect 1703 1388 1705 1428
rect 1709 1388 1711 1428
rect 1689 1348 1699 1388
rect 1775 1356 1777 1436
rect 1781 1356 1785 1436
rect 1789 1356 1791 1436
rect 1853 1356 1855 1436
rect 1859 1356 1865 1436
rect 1869 1356 1871 1436
rect 1893 1356 1895 1436
rect 1899 1356 1905 1436
rect 1909 1356 1911 1436
rect 1968 1396 1970 1436
rect 1974 1396 1978 1436
rect 1990 1356 1992 1436
rect 1996 1356 2000 1436
rect 2004 1356 2006 1436
rect 2049 1396 2051 1436
rect 2055 1396 2057 1436
rect 2114 1356 2116 1436
rect 2120 1356 2124 1436
rect 2128 1356 2130 1436
rect 2142 1396 2146 1436
rect 2150 1396 2152 1436
rect 2209 1396 2211 1436
rect 2215 1396 2217 1436
rect 2229 1396 2231 1436
rect 2235 1396 2237 1436
rect 2332 1428 2341 1436
rect 2289 1388 2291 1428
rect 2295 1388 2297 1428
rect 2309 1388 2311 1428
rect 2301 1348 2311 1388
rect 2315 1348 2321 1428
rect 2325 1364 2327 1428
rect 2339 1364 2341 1428
rect 2325 1356 2341 1364
rect 2345 1356 2351 1436
rect 2355 1356 2357 1436
rect 2423 1356 2425 1436
rect 2429 1356 2435 1436
rect 2439 1428 2448 1436
rect 2439 1364 2441 1428
rect 2453 1364 2455 1428
rect 2439 1356 2455 1364
rect 2325 1348 2333 1356
rect 2447 1348 2455 1356
rect 2459 1348 2465 1428
rect 2469 1388 2471 1428
rect 2483 1388 2485 1428
rect 2489 1388 2491 1428
rect 2469 1348 2479 1388
rect 2543 1356 2545 1436
rect 2549 1424 2565 1436
rect 2549 1356 2551 1424
rect 2563 1356 2565 1424
rect 2569 1358 2571 1436
rect 2583 1358 2585 1436
rect 2569 1356 2585 1358
rect 2589 1370 2591 1436
rect 2603 1370 2605 1436
rect 2589 1356 2605 1370
rect 2609 1358 2611 1436
rect 2609 1356 2623 1358
rect 2649 1358 2651 1436
rect 2637 1356 2651 1358
rect 2655 1370 2657 1436
rect 2669 1370 2671 1436
rect 2655 1356 2671 1370
rect 2675 1358 2677 1436
rect 2689 1358 2691 1436
rect 2675 1356 2691 1358
rect 2695 1424 2711 1436
rect 2695 1356 2697 1424
rect 2709 1356 2711 1424
rect 2715 1356 2717 1436
rect 2783 1356 2785 1436
rect 2789 1424 2805 1436
rect 2789 1356 2791 1424
rect 2803 1356 2805 1424
rect 2809 1358 2811 1436
rect 2823 1358 2825 1436
rect 2809 1356 2825 1358
rect 2829 1370 2831 1436
rect 2843 1370 2845 1436
rect 2829 1356 2845 1370
rect 2849 1358 2851 1436
rect 2889 1396 2891 1436
rect 2895 1396 2899 1436
rect 2849 1356 2863 1358
rect 2911 1356 2913 1436
rect 2917 1356 2919 1436
rect 2983 1356 2985 1436
rect 2989 1424 3005 1436
rect 2989 1356 2991 1424
rect 3003 1356 3005 1424
rect 3009 1358 3011 1436
rect 3023 1358 3025 1436
rect 3009 1356 3025 1358
rect 3029 1370 3031 1436
rect 3043 1370 3045 1436
rect 3029 1356 3045 1370
rect 3049 1358 3051 1436
rect 3103 1396 3105 1436
rect 3109 1396 3111 1436
rect 3049 1356 3063 1358
rect 3163 1356 3165 1436
rect 3169 1356 3175 1436
rect 3179 1428 3188 1436
rect 3179 1364 3181 1428
rect 3193 1364 3195 1428
rect 3179 1356 3195 1364
rect 3187 1348 3195 1356
rect 3199 1348 3205 1428
rect 3209 1388 3211 1428
rect 3223 1388 3225 1428
rect 3229 1388 3231 1428
rect 3209 1348 3219 1388
rect 3273 1356 3275 1436
rect 3279 1396 3281 1436
rect 3293 1396 3295 1436
rect 3299 1396 3309 1436
rect 3313 1396 3315 1436
rect 3327 1396 3329 1436
rect 3333 1396 3341 1436
rect 3345 1396 3347 1436
rect 3359 1396 3361 1436
rect 3365 1396 3367 1436
rect 3405 1396 3407 1436
rect 3411 1396 3415 1436
rect 3419 1416 3421 1436
rect 3433 1416 3435 1436
rect 3439 1416 3443 1436
rect 3447 1416 3451 1436
rect 3463 1416 3465 1436
rect 3419 1396 3430 1416
rect 3279 1356 3288 1396
rect 3456 1356 3465 1416
rect 3469 1356 3471 1436
rect 3535 1356 3537 1436
rect 3541 1356 3545 1436
rect 3549 1356 3551 1436
rect 3613 1356 3615 1436
rect 3619 1356 3625 1436
rect 3629 1356 3631 1436
rect 3653 1356 3655 1436
rect 3659 1356 3665 1436
rect 3669 1356 3671 1436
rect 3728 1396 3730 1436
rect 3734 1396 3738 1436
rect 3750 1356 3752 1436
rect 3756 1356 3760 1436
rect 3764 1356 3766 1436
rect 3823 1396 3825 1436
rect 3829 1396 3831 1436
rect 3869 1356 3871 1436
rect 3875 1416 3877 1436
rect 3889 1416 3893 1436
rect 3897 1416 3901 1436
rect 3905 1416 3907 1436
rect 3919 1416 3921 1436
rect 3875 1356 3884 1416
rect 3910 1396 3921 1416
rect 3925 1396 3929 1436
rect 3933 1396 3935 1436
rect 3973 1396 3975 1436
rect 3979 1396 3981 1436
rect 3993 1396 3995 1436
rect 3999 1396 4007 1436
rect 4011 1396 4013 1436
rect 4025 1396 4027 1436
rect 4031 1396 4041 1436
rect 4045 1396 4047 1436
rect 4059 1396 4061 1436
rect 4052 1356 4061 1396
rect 4065 1356 4067 1436
rect 4109 1356 4111 1436
rect 4115 1416 4117 1436
rect 4129 1416 4133 1436
rect 4137 1416 4141 1436
rect 4145 1416 4147 1436
rect 4159 1416 4161 1436
rect 4115 1356 4124 1416
rect 4150 1396 4161 1416
rect 4165 1396 4169 1436
rect 4173 1396 4175 1436
rect 4213 1396 4215 1436
rect 4219 1396 4221 1436
rect 4233 1396 4235 1436
rect 4239 1396 4247 1436
rect 4251 1396 4253 1436
rect 4265 1396 4267 1436
rect 4271 1396 4281 1436
rect 4285 1396 4287 1436
rect 4299 1396 4301 1436
rect 4292 1356 4301 1396
rect 4305 1356 4307 1436
rect 4363 1396 4365 1436
rect 4369 1396 4371 1436
rect 4409 1358 4411 1436
rect 4397 1356 4411 1358
rect 4415 1370 4417 1436
rect 4429 1370 4431 1436
rect 4415 1356 4431 1370
rect 4435 1358 4437 1436
rect 4449 1358 4451 1436
rect 4435 1356 4451 1358
rect 4455 1424 4471 1436
rect 4455 1356 4457 1424
rect 4469 1356 4471 1424
rect 4475 1356 4477 1436
rect 4572 1428 4581 1436
rect 4529 1388 4531 1428
rect 4535 1388 4537 1428
rect 4549 1388 4551 1428
rect 4541 1348 4551 1388
rect 4555 1348 4561 1428
rect 4565 1364 4567 1428
rect 4579 1364 4581 1428
rect 4565 1356 4581 1364
rect 4585 1356 4591 1436
rect 4595 1356 4597 1436
rect 4663 1356 4665 1436
rect 4669 1424 4685 1436
rect 4669 1356 4671 1424
rect 4683 1356 4685 1424
rect 4689 1358 4691 1436
rect 4703 1358 4705 1436
rect 4689 1356 4705 1358
rect 4709 1370 4711 1436
rect 4723 1370 4725 1436
rect 4709 1356 4725 1370
rect 4729 1358 4731 1436
rect 4729 1356 4743 1358
rect 4781 1356 4783 1436
rect 4787 1356 4789 1436
rect 4801 1396 4805 1436
rect 4809 1396 4811 1436
rect 4863 1396 4865 1436
rect 4869 1396 4871 1436
rect 4883 1396 4885 1436
rect 4889 1396 4891 1436
rect 4943 1396 4945 1436
rect 4949 1396 4951 1436
rect 4963 1396 4965 1436
rect 4969 1396 4971 1436
rect 4565 1348 4573 1356
rect 5033 1356 5035 1436
rect 5039 1356 5045 1436
rect 5049 1356 5051 1436
rect 5073 1356 5075 1436
rect 5079 1356 5085 1436
rect 5089 1356 5091 1436
rect 5153 1356 5155 1436
rect 5159 1356 5165 1436
rect 5169 1356 5171 1436
rect 5193 1356 5195 1436
rect 5199 1356 5205 1436
rect 5209 1356 5211 1436
rect 5249 1356 5251 1436
rect 5255 1356 5257 1436
rect 5323 1396 5325 1436
rect 5329 1396 5331 1436
rect 5343 1396 5345 1436
rect 5349 1396 5351 1436
rect 5389 1356 5391 1436
rect 5395 1356 5401 1436
rect 5405 1356 5407 1436
rect 5429 1356 5431 1436
rect 5435 1356 5441 1436
rect 5445 1356 5447 1436
rect 5523 1356 5525 1436
rect 5529 1356 5531 1436
rect 5543 1356 5545 1436
rect 5549 1368 5551 1436
rect 5563 1368 5565 1436
rect 5549 1356 5565 1368
rect 5569 1364 5571 1436
rect 5569 1356 5583 1364
rect 5609 1356 5611 1436
rect 5615 1356 5617 1436
rect 5712 1428 5721 1436
rect 5669 1388 5671 1428
rect 5675 1388 5677 1428
rect 5689 1388 5691 1428
rect 5681 1348 5691 1388
rect 5695 1348 5701 1428
rect 5705 1364 5707 1428
rect 5719 1364 5721 1428
rect 5705 1356 5721 1364
rect 5725 1356 5731 1436
rect 5735 1356 5737 1436
rect 5803 1396 5805 1436
rect 5809 1396 5811 1436
rect 5823 1396 5825 1436
rect 5829 1396 5831 1436
rect 5888 1396 5890 1436
rect 5894 1396 5898 1436
rect 5705 1348 5713 1356
rect 5910 1356 5912 1436
rect 5916 1356 5920 1436
rect 5924 1356 5926 1436
rect 5983 1396 5985 1436
rect 5989 1396 5991 1436
rect 6034 1356 6036 1436
rect 6040 1356 6044 1436
rect 6048 1356 6050 1436
rect 6062 1396 6066 1436
rect 6070 1396 6072 1436
rect 6129 1356 6131 1436
rect 6135 1356 6141 1436
rect 6145 1356 6147 1436
rect 6169 1356 6171 1436
rect 6175 1356 6181 1436
rect 6185 1356 6187 1436
rect 6249 1356 6251 1436
rect 6255 1416 6257 1436
rect 6269 1416 6273 1436
rect 6277 1416 6281 1436
rect 6285 1416 6287 1436
rect 6299 1416 6301 1436
rect 6255 1356 6264 1416
rect 6290 1396 6301 1416
rect 6305 1396 6309 1436
rect 6313 1396 6315 1436
rect 6353 1396 6355 1436
rect 6359 1396 6361 1436
rect 6373 1396 6375 1436
rect 6379 1396 6387 1436
rect 6391 1396 6393 1436
rect 6405 1396 6407 1436
rect 6411 1396 6421 1436
rect 6425 1396 6427 1436
rect 6439 1396 6441 1436
rect 6432 1356 6441 1396
rect 6445 1356 6447 1436
rect 6489 1356 6491 1436
rect 6495 1416 6497 1436
rect 6509 1416 6513 1436
rect 6517 1416 6521 1436
rect 6525 1416 6527 1436
rect 6539 1416 6541 1436
rect 6495 1356 6504 1416
rect 6530 1396 6541 1416
rect 6545 1396 6549 1436
rect 6553 1396 6555 1436
rect 6593 1396 6595 1436
rect 6599 1396 6601 1436
rect 6613 1396 6615 1436
rect 6619 1396 6627 1436
rect 6631 1396 6633 1436
rect 6645 1396 6647 1436
rect 6651 1396 6661 1436
rect 6665 1396 6667 1436
rect 6679 1396 6681 1436
rect 6672 1356 6681 1396
rect 6685 1356 6687 1436
rect 29 984 31 1064
rect 35 1004 44 1064
rect 212 1024 221 1064
rect 70 1004 81 1024
rect 35 984 37 1004
rect 49 984 53 1004
rect 57 984 61 1004
rect 65 984 67 1004
rect 79 984 81 1004
rect 85 984 89 1024
rect 93 984 95 1024
rect 133 984 135 1024
rect 139 984 141 1024
rect 153 984 155 1024
rect 159 984 167 1024
rect 171 984 173 1024
rect 185 984 187 1024
rect 191 984 201 1024
rect 205 984 207 1024
rect 219 984 221 1024
rect 225 984 227 1064
rect 283 984 285 1024
rect 289 984 291 1024
rect 329 984 331 1064
rect 335 1004 344 1064
rect 512 1024 521 1064
rect 370 1004 381 1024
rect 335 984 337 1004
rect 349 984 353 1004
rect 357 984 361 1004
rect 365 984 367 1004
rect 379 984 381 1004
rect 385 984 389 1024
rect 393 984 395 1024
rect 433 984 435 1024
rect 439 984 441 1024
rect 453 984 455 1024
rect 459 984 467 1024
rect 471 984 473 1024
rect 485 984 487 1024
rect 491 984 501 1024
rect 505 984 507 1024
rect 519 984 521 1024
rect 525 984 527 1064
rect 569 984 571 1024
rect 575 984 577 1024
rect 629 984 631 1024
rect 635 984 637 1024
rect 649 984 651 1024
rect 655 1020 671 1024
rect 655 984 657 1020
rect 669 984 671 1020
rect 675 984 677 1024
rect 729 984 731 1064
rect 735 984 739 1064
rect 743 984 745 1064
rect 809 984 811 1024
rect 815 984 817 1024
rect 829 984 831 1024
rect 835 1020 851 1024
rect 835 984 837 1020
rect 849 984 851 1020
rect 855 984 857 1024
rect 909 984 911 1024
rect 915 984 917 1024
rect 929 984 931 1024
rect 935 984 937 1024
rect 989 984 991 1024
rect 995 984 997 1024
rect 1053 984 1055 1064
rect 1059 1024 1068 1064
rect 1059 984 1061 1024
rect 1073 984 1075 1024
rect 1079 984 1089 1024
rect 1093 984 1095 1024
rect 1107 984 1109 1024
rect 1113 984 1121 1024
rect 1125 984 1127 1024
rect 1139 984 1141 1024
rect 1145 984 1147 1024
rect 1185 984 1187 1024
rect 1191 984 1195 1024
rect 1199 1004 1210 1024
rect 1236 1004 1245 1064
rect 1199 984 1201 1004
rect 1213 984 1215 1004
rect 1219 984 1223 1004
rect 1227 984 1231 1004
rect 1243 984 1245 1004
rect 1249 984 1251 1064
rect 1289 984 1291 1064
rect 1295 984 1297 1064
rect 1309 984 1311 1064
rect 1315 984 1317 1064
rect 1329 984 1331 1064
rect 1335 984 1337 1064
rect 1349 984 1351 1064
rect 1355 984 1357 1064
rect 1369 984 1371 1064
rect 1375 984 1377 1064
rect 1389 984 1391 1064
rect 1395 984 1397 1064
rect 1409 984 1411 1064
rect 1415 984 1417 1064
rect 1429 984 1431 1064
rect 1435 984 1437 1064
rect 1493 984 1495 1064
rect 1499 1024 1508 1064
rect 1499 984 1501 1024
rect 1513 984 1515 1024
rect 1519 984 1529 1024
rect 1533 984 1535 1024
rect 1547 984 1549 1024
rect 1553 984 1561 1024
rect 1565 984 1567 1024
rect 1579 984 1581 1024
rect 1585 984 1587 1024
rect 1625 984 1627 1024
rect 1631 984 1635 1024
rect 1639 1004 1650 1024
rect 1676 1004 1685 1064
rect 1639 984 1641 1004
rect 1653 984 1655 1004
rect 1659 984 1663 1004
rect 1667 984 1671 1004
rect 1683 984 1685 1004
rect 1689 984 1691 1064
rect 1755 984 1757 1064
rect 1761 984 1765 1064
rect 1769 984 1771 1064
rect 1833 984 1835 1064
rect 1839 984 1845 1064
rect 1849 984 1851 1064
rect 1873 984 1875 1064
rect 1879 984 1885 1064
rect 1889 984 1891 1064
rect 1948 984 1950 1024
rect 1954 984 1958 1024
rect 1970 984 1972 1064
rect 1976 984 1980 1064
rect 1984 984 1986 1064
rect 2048 984 2050 1024
rect 2054 984 2058 1024
rect 2070 984 2072 1064
rect 2076 984 2080 1064
rect 2084 984 2086 1064
rect 2155 984 2157 1064
rect 2161 984 2165 1064
rect 2169 984 2171 1064
rect 2233 984 2235 1064
rect 2239 984 2245 1064
rect 2249 984 2251 1064
rect 2273 984 2275 1064
rect 2279 984 2285 1064
rect 2289 984 2291 1064
rect 2333 984 2335 1064
rect 2339 1024 2348 1064
rect 2339 984 2341 1024
rect 2353 984 2355 1024
rect 2359 984 2369 1024
rect 2373 984 2375 1024
rect 2387 984 2389 1024
rect 2393 984 2401 1024
rect 2405 984 2407 1024
rect 2419 984 2421 1024
rect 2425 984 2427 1024
rect 2465 984 2467 1024
rect 2471 984 2475 1024
rect 2479 1004 2490 1024
rect 2516 1004 2525 1064
rect 2479 984 2481 1004
rect 2493 984 2495 1004
rect 2499 984 2503 1004
rect 2507 984 2511 1004
rect 2523 984 2525 1004
rect 2529 984 2531 1064
rect 2583 984 2585 1024
rect 2589 984 2591 1024
rect 2634 984 2636 1064
rect 2640 984 2644 1064
rect 2648 984 2650 1064
rect 2662 984 2666 1024
rect 2670 984 2672 1024
rect 2741 984 2743 1064
rect 2747 984 2749 1064
rect 2761 984 2765 1024
rect 2769 984 2771 1024
rect 2809 984 2811 1024
rect 2815 984 2817 1024
rect 2883 984 2885 1064
rect 2889 996 2891 1064
rect 2903 996 2905 1064
rect 2889 984 2905 996
rect 2909 1062 2925 1064
rect 2909 984 2911 1062
rect 2923 984 2925 1062
rect 2929 1050 2945 1064
rect 2929 984 2931 1050
rect 2943 984 2945 1050
rect 2949 1062 2963 1064
rect 2949 984 2951 1062
rect 2993 984 2995 1064
rect 2999 1024 3008 1064
rect 2999 984 3001 1024
rect 3013 984 3015 1024
rect 3019 984 3029 1024
rect 3033 984 3035 1024
rect 3047 984 3049 1024
rect 3053 984 3061 1024
rect 3065 984 3067 1024
rect 3079 984 3081 1024
rect 3085 984 3087 1024
rect 3125 984 3127 1024
rect 3131 984 3135 1024
rect 3139 1004 3150 1024
rect 3176 1004 3185 1064
rect 3139 984 3141 1004
rect 3153 984 3155 1004
rect 3159 984 3163 1004
rect 3167 984 3171 1004
rect 3183 984 3185 1004
rect 3189 984 3191 1064
rect 3347 1064 3355 1072
rect 3229 984 3231 1024
rect 3235 984 3237 1024
rect 3249 984 3251 1024
rect 3255 984 3257 1024
rect 3323 984 3325 1064
rect 3329 984 3335 1064
rect 3339 1056 3355 1064
rect 3339 992 3341 1056
rect 3353 992 3355 1056
rect 3359 992 3365 1072
rect 3369 1032 3379 1072
rect 3441 1032 3451 1072
rect 3369 992 3371 1032
rect 3383 992 3385 1032
rect 3389 992 3391 1032
rect 3429 992 3431 1032
rect 3435 992 3437 1032
rect 3449 992 3451 1032
rect 3455 992 3461 1072
rect 3465 1064 3473 1072
rect 3465 1056 3481 1064
rect 3465 992 3467 1056
rect 3479 992 3481 1056
rect 3339 984 3348 992
rect 3472 984 3481 992
rect 3485 984 3491 1064
rect 3495 984 3497 1064
rect 3561 984 3563 1064
rect 3567 984 3569 1064
rect 3581 984 3585 1024
rect 3589 984 3591 1024
rect 3633 984 3635 1064
rect 3639 1024 3648 1064
rect 3639 984 3641 1024
rect 3653 984 3655 1024
rect 3659 984 3669 1024
rect 3673 984 3675 1024
rect 3687 984 3689 1024
rect 3693 984 3701 1024
rect 3705 984 3707 1024
rect 3719 984 3721 1024
rect 3725 984 3727 1024
rect 3765 984 3767 1024
rect 3771 984 3775 1024
rect 3779 1004 3790 1024
rect 3816 1004 3825 1064
rect 3779 984 3781 1004
rect 3793 984 3795 1004
rect 3799 984 3803 1004
rect 3807 984 3811 1004
rect 3823 984 3825 1004
rect 3829 984 3831 1064
rect 3881 1032 3891 1072
rect 3869 992 3871 1032
rect 3875 992 3877 1032
rect 3889 992 3891 1032
rect 3895 992 3901 1072
rect 3905 1064 3913 1072
rect 4027 1064 4035 1072
rect 3905 1056 3921 1064
rect 3905 992 3907 1056
rect 3919 992 3921 1056
rect 3912 984 3921 992
rect 3925 984 3931 1064
rect 3935 984 3937 1064
rect 4003 984 4005 1064
rect 4009 984 4015 1064
rect 4019 1056 4035 1064
rect 4019 992 4021 1056
rect 4033 992 4035 1056
rect 4039 992 4045 1072
rect 4049 1032 4059 1072
rect 4049 992 4051 1032
rect 4063 992 4065 1032
rect 4069 992 4071 1032
rect 4019 984 4028 992
rect 4109 984 4111 1024
rect 4115 984 4117 1024
rect 4169 984 4171 1064
rect 4175 984 4181 1064
rect 4185 984 4187 1064
rect 4209 984 4211 1064
rect 4215 984 4221 1064
rect 4225 984 4227 1064
rect 4289 984 4291 1064
rect 4295 984 4299 1064
rect 4303 984 4305 1064
rect 4388 984 4390 1024
rect 4394 984 4398 1024
rect 4410 984 4412 1064
rect 4416 984 4420 1064
rect 4424 984 4426 1064
rect 4483 984 4485 1064
rect 4489 984 4491 1064
rect 4503 984 4505 1064
rect 4509 1052 4525 1064
rect 4509 984 4511 1052
rect 4523 984 4525 1052
rect 4529 1056 4543 1064
rect 4529 984 4531 1056
rect 4573 984 4575 1064
rect 4579 1024 4588 1064
rect 4579 984 4581 1024
rect 4593 984 4595 1024
rect 4599 984 4609 1024
rect 4613 984 4615 1024
rect 4627 984 4629 1024
rect 4633 984 4641 1024
rect 4645 984 4647 1024
rect 4659 984 4661 1024
rect 4665 984 4667 1024
rect 4705 984 4707 1024
rect 4711 984 4715 1024
rect 4719 1004 4730 1024
rect 4756 1004 4765 1064
rect 4719 984 4721 1004
rect 4733 984 4735 1004
rect 4739 984 4743 1004
rect 4747 984 4751 1004
rect 4763 984 4765 1004
rect 4769 984 4771 1064
rect 4809 984 4811 1064
rect 4815 984 4821 1064
rect 4825 984 4827 1064
rect 4849 984 4851 1064
rect 4855 984 4861 1064
rect 4865 984 4867 1064
rect 4955 984 4957 1064
rect 4961 984 4965 1064
rect 4969 984 4971 1064
rect 5028 984 5030 1024
rect 5034 984 5038 1024
rect 5050 984 5052 1064
rect 5056 984 5060 1064
rect 5064 984 5066 1064
rect 5135 984 5137 1064
rect 5141 984 5145 1064
rect 5149 984 5151 1064
rect 5189 984 5191 1064
rect 5195 984 5199 1064
rect 5203 984 5205 1064
rect 5269 984 5271 1064
rect 5275 984 5279 1064
rect 5283 984 5285 1064
rect 5361 984 5363 1064
rect 5367 984 5369 1064
rect 5381 984 5385 1024
rect 5389 984 5391 1024
rect 5429 984 5431 1064
rect 5435 984 5439 1064
rect 5443 984 5445 1064
rect 5509 984 5511 1064
rect 5515 984 5519 1064
rect 5523 984 5525 1064
rect 5577 1056 5591 1064
rect 5589 984 5591 1056
rect 5595 1052 5611 1064
rect 5595 984 5597 1052
rect 5609 984 5611 1052
rect 5615 984 5617 1064
rect 5629 984 5631 1064
rect 5635 984 5637 1064
rect 5689 984 5691 1064
rect 5695 984 5701 1064
rect 5705 1063 5721 1064
rect 5705 984 5707 1063
rect 5719 984 5721 1063
rect 5725 1063 5739 1064
rect 5725 984 5727 1063
rect 5815 984 5817 1064
rect 5821 984 5825 1064
rect 5829 984 5831 1064
rect 5874 984 5876 1064
rect 5880 984 5884 1064
rect 5888 984 5890 1064
rect 5902 984 5906 1024
rect 5910 984 5912 1024
rect 5983 984 5985 1024
rect 5989 1020 6005 1024
rect 5989 984 5991 1020
rect 6003 984 6005 1020
rect 6009 984 6011 1024
rect 6023 984 6025 1024
rect 6029 984 6031 1024
rect 6074 984 6076 1064
rect 6080 984 6084 1064
rect 6088 984 6090 1064
rect 6102 984 6106 1024
rect 6110 984 6112 1024
rect 6195 984 6197 1064
rect 6201 984 6205 1064
rect 6209 984 6211 1064
rect 6249 984 6251 1064
rect 6255 984 6259 1064
rect 6263 984 6265 1064
rect 6329 984 6331 1064
rect 6335 1004 6344 1064
rect 6512 1024 6521 1064
rect 6370 1004 6381 1024
rect 6335 984 6337 1004
rect 6349 984 6353 1004
rect 6357 984 6361 1004
rect 6365 984 6367 1004
rect 6379 984 6381 1004
rect 6385 984 6389 1024
rect 6393 984 6395 1024
rect 6433 984 6435 1024
rect 6439 984 6441 1024
rect 6453 984 6455 1024
rect 6459 984 6467 1024
rect 6471 984 6473 1024
rect 6485 984 6487 1024
rect 6491 984 6501 1024
rect 6505 984 6507 1024
rect 6519 984 6521 1024
rect 6525 984 6527 1064
rect 6569 984 6571 1064
rect 6575 984 6581 1064
rect 6585 984 6587 1064
rect 6609 984 6611 1064
rect 6615 984 6621 1064
rect 6625 984 6627 1064
rect 29 876 31 956
rect 35 876 41 956
rect 45 877 47 956
rect 59 877 61 956
rect 45 876 61 877
rect 65 877 67 956
rect 143 916 145 956
rect 149 916 151 956
rect 163 916 165 956
rect 169 916 171 956
rect 65 876 79 877
rect 209 876 211 956
rect 215 936 217 956
rect 229 936 233 956
rect 237 936 241 956
rect 245 936 247 956
rect 259 936 261 956
rect 215 876 224 936
rect 250 916 261 936
rect 265 916 269 956
rect 273 916 275 956
rect 313 916 315 956
rect 319 916 321 956
rect 333 916 335 956
rect 339 916 347 956
rect 351 916 353 956
rect 365 916 367 956
rect 371 916 381 956
rect 385 916 387 956
rect 399 916 401 956
rect 392 876 401 916
rect 405 876 407 956
rect 463 916 465 956
rect 469 916 471 956
rect 535 876 537 956
rect 541 876 545 956
rect 549 876 551 956
rect 589 876 591 956
rect 595 876 599 956
rect 603 876 605 956
rect 669 916 671 956
rect 675 916 677 956
rect 689 916 691 956
rect 695 916 697 956
rect 749 916 751 956
rect 755 916 757 956
rect 769 916 771 956
rect 775 920 777 956
rect 789 920 791 956
rect 775 916 791 920
rect 795 916 797 956
rect 849 876 851 956
rect 855 876 861 956
rect 865 876 867 956
rect 889 876 891 956
rect 895 876 901 956
rect 905 876 907 956
rect 974 876 976 956
rect 980 876 984 956
rect 988 876 990 956
rect 1002 916 1006 956
rect 1010 916 1012 956
rect 1074 876 1076 956
rect 1080 876 1084 956
rect 1088 876 1090 956
rect 1102 916 1106 956
rect 1110 916 1112 956
rect 1179 888 1181 948
rect 1185 944 1201 948
rect 1185 892 1187 944
rect 1199 892 1201 944
rect 1185 888 1201 892
rect 1205 888 1207 948
rect 1243 898 1245 956
rect 1231 896 1245 898
rect 1249 944 1265 956
rect 1249 896 1251 944
rect 1263 896 1265 944
rect 1269 896 1271 956
rect 1283 896 1285 956
rect 1289 896 1291 956
rect 1303 896 1305 956
rect 1309 896 1311 956
rect 1354 876 1356 956
rect 1360 876 1364 956
rect 1368 876 1370 956
rect 1382 916 1386 956
rect 1390 916 1392 956
rect 1463 916 1465 956
rect 1469 916 1471 956
rect 1513 876 1515 956
rect 1519 916 1521 956
rect 1533 916 1535 956
rect 1539 916 1549 956
rect 1553 916 1555 956
rect 1567 916 1569 956
rect 1573 916 1581 956
rect 1585 916 1587 956
rect 1599 916 1601 956
rect 1605 916 1607 956
rect 1645 916 1647 956
rect 1651 916 1655 956
rect 1659 936 1661 956
rect 1673 936 1675 956
rect 1679 936 1683 956
rect 1687 936 1691 956
rect 1703 936 1705 956
rect 1659 916 1670 936
rect 1519 876 1528 916
rect 1696 876 1705 936
rect 1709 876 1711 956
rect 1749 916 1751 956
rect 1755 916 1757 956
rect 1852 948 1861 956
rect 1809 908 1811 948
rect 1815 908 1817 948
rect 1829 908 1831 948
rect 1821 868 1831 908
rect 1835 868 1841 948
rect 1845 884 1847 948
rect 1859 884 1861 948
rect 1845 876 1861 884
rect 1865 876 1871 956
rect 1875 876 1877 956
rect 1934 876 1936 956
rect 1940 876 1944 956
rect 1948 876 1950 956
rect 1962 916 1966 956
rect 1970 916 1972 956
rect 2029 916 2031 956
rect 2035 916 2037 956
rect 2049 916 2051 956
rect 2055 916 2057 956
rect 1845 868 1853 876
rect 2109 876 2111 956
rect 2115 936 2117 956
rect 2129 936 2133 956
rect 2137 936 2141 956
rect 2145 936 2147 956
rect 2159 936 2161 956
rect 2115 876 2124 936
rect 2150 916 2161 936
rect 2165 916 2169 956
rect 2173 916 2175 956
rect 2213 916 2215 956
rect 2219 916 2221 956
rect 2233 916 2235 956
rect 2239 916 2247 956
rect 2251 916 2253 956
rect 2265 916 2267 956
rect 2271 916 2281 956
rect 2285 916 2287 956
rect 2299 916 2301 956
rect 2292 876 2301 916
rect 2305 876 2307 956
rect 2349 916 2351 956
rect 2355 916 2357 956
rect 2409 876 2411 956
rect 2415 876 2421 956
rect 2425 876 2427 956
rect 2449 876 2451 956
rect 2455 876 2461 956
rect 2465 876 2467 956
rect 2529 876 2531 956
rect 2535 876 2539 956
rect 2543 876 2545 956
rect 2628 916 2630 956
rect 2634 916 2638 956
rect 2650 876 2652 956
rect 2656 876 2660 956
rect 2664 876 2666 956
rect 2723 876 2725 956
rect 2729 876 2731 956
rect 2743 876 2745 956
rect 2749 876 2751 956
rect 2763 876 2765 956
rect 2769 876 2771 956
rect 2783 876 2785 956
rect 2789 876 2791 956
rect 2803 876 2805 956
rect 2809 876 2811 956
rect 2823 876 2825 956
rect 2829 876 2831 956
rect 2843 876 2845 956
rect 2849 876 2851 956
rect 2863 876 2865 956
rect 2869 876 2871 956
rect 2909 884 2911 956
rect 2897 876 2911 884
rect 2915 888 2917 956
rect 2929 888 2931 956
rect 2915 876 2931 888
rect 2935 876 2937 956
rect 2949 876 2951 956
rect 2955 876 2957 956
rect 3023 876 3025 956
rect 3029 876 3031 956
rect 3043 876 3045 956
rect 3049 888 3051 956
rect 3063 888 3065 956
rect 3049 876 3065 888
rect 3069 884 3071 956
rect 3069 876 3083 884
rect 3123 876 3125 956
rect 3129 876 3135 956
rect 3139 948 3148 956
rect 3139 884 3141 948
rect 3153 884 3155 948
rect 3139 876 3155 884
rect 3147 868 3155 876
rect 3159 868 3165 948
rect 3169 908 3171 948
rect 3183 908 3185 948
rect 3189 908 3191 948
rect 3169 868 3179 908
rect 3243 876 3245 956
rect 3249 876 3255 956
rect 3259 948 3268 956
rect 3259 884 3261 948
rect 3273 884 3275 948
rect 3259 876 3275 884
rect 3267 868 3275 876
rect 3279 868 3285 948
rect 3289 908 3291 948
rect 3303 908 3305 948
rect 3309 908 3311 948
rect 3368 916 3370 956
rect 3374 916 3378 956
rect 3289 868 3299 908
rect 3390 876 3392 956
rect 3396 876 3400 956
rect 3404 876 3406 956
rect 3449 916 3451 956
rect 3455 916 3457 956
rect 3469 916 3471 956
rect 3475 916 3477 956
rect 3572 948 3581 956
rect 3529 908 3531 948
rect 3535 908 3537 948
rect 3549 908 3551 948
rect 3541 868 3551 908
rect 3555 868 3561 948
rect 3565 884 3567 948
rect 3579 884 3581 948
rect 3565 876 3581 884
rect 3585 876 3591 956
rect 3595 876 3597 956
rect 3663 916 3665 956
rect 3669 916 3671 956
rect 3565 868 3573 876
rect 3723 876 3725 956
rect 3729 876 3735 956
rect 3739 948 3748 956
rect 3739 884 3741 948
rect 3753 884 3755 948
rect 3739 876 3755 884
rect 3747 868 3755 876
rect 3759 868 3765 948
rect 3769 908 3771 948
rect 3783 908 3785 948
rect 3789 908 3791 948
rect 3769 868 3779 908
rect 3833 876 3835 956
rect 3839 916 3841 956
rect 3853 916 3855 956
rect 3859 916 3869 956
rect 3873 916 3875 956
rect 3887 916 3889 956
rect 3893 916 3901 956
rect 3905 916 3907 956
rect 3919 916 3921 956
rect 3925 916 3927 956
rect 3965 916 3967 956
rect 3971 916 3975 956
rect 3979 936 3981 956
rect 3993 936 3995 956
rect 3999 936 4003 956
rect 4007 936 4011 956
rect 4023 936 4025 956
rect 3979 916 3990 936
rect 3839 876 3848 916
rect 4016 876 4025 936
rect 4029 876 4031 956
rect 4112 948 4121 956
rect 4069 908 4071 948
rect 4075 908 4077 948
rect 4089 908 4091 948
rect 4081 868 4091 908
rect 4095 868 4101 948
rect 4105 884 4107 948
rect 4119 884 4121 948
rect 4105 876 4121 884
rect 4125 876 4131 956
rect 4135 876 4137 956
rect 4189 884 4191 956
rect 4177 876 4191 884
rect 4195 888 4197 956
rect 4209 888 4211 956
rect 4195 876 4211 888
rect 4215 876 4217 956
rect 4229 876 4231 956
rect 4235 876 4237 956
rect 4294 876 4296 956
rect 4300 876 4304 956
rect 4308 876 4310 956
rect 4322 916 4326 956
rect 4330 916 4332 956
rect 4403 916 4405 956
rect 4409 920 4411 956
rect 4423 920 4425 956
rect 4409 916 4425 920
rect 4429 916 4431 956
rect 4443 916 4445 956
rect 4449 916 4451 956
rect 4489 916 4491 956
rect 4495 916 4497 956
rect 4105 868 4113 876
rect 4554 876 4556 956
rect 4560 876 4564 956
rect 4568 876 4570 956
rect 4582 916 4586 956
rect 4590 916 4592 956
rect 4649 916 4651 956
rect 4655 916 4657 956
rect 4669 916 4671 956
rect 4675 916 4677 956
rect 4743 916 4745 956
rect 4749 916 4751 956
rect 4794 876 4796 956
rect 4800 876 4804 956
rect 4808 876 4810 956
rect 4822 916 4826 956
rect 4830 916 4832 956
rect 4889 916 4891 956
rect 4895 916 4897 956
rect 4909 916 4911 956
rect 4915 916 4917 956
rect 5012 948 5021 956
rect 4969 908 4971 948
rect 4975 908 4977 948
rect 4989 908 4991 948
rect 4981 868 4991 908
rect 4995 868 5001 948
rect 5005 884 5007 948
rect 5019 884 5021 948
rect 5005 876 5021 884
rect 5025 876 5031 956
rect 5035 876 5037 956
rect 5103 876 5105 956
rect 5109 876 5115 956
rect 5119 948 5128 956
rect 5119 884 5121 948
rect 5133 884 5135 948
rect 5119 876 5135 884
rect 5005 868 5013 876
rect 5127 868 5135 876
rect 5139 868 5145 948
rect 5149 908 5151 948
rect 5163 908 5165 948
rect 5169 908 5171 948
rect 5149 868 5159 908
rect 5209 876 5211 956
rect 5215 876 5217 956
rect 5229 876 5231 956
rect 5235 876 5237 956
rect 5249 876 5251 956
rect 5255 876 5257 956
rect 5269 876 5271 956
rect 5275 876 5277 956
rect 5289 876 5291 956
rect 5295 876 5297 956
rect 5309 876 5311 956
rect 5315 876 5317 956
rect 5329 876 5331 956
rect 5335 876 5337 956
rect 5349 876 5351 956
rect 5355 876 5357 956
rect 5409 884 5411 956
rect 5397 876 5411 884
rect 5415 888 5417 956
rect 5429 888 5431 956
rect 5415 876 5431 888
rect 5435 876 5437 956
rect 5449 876 5451 956
rect 5455 876 5457 956
rect 5523 916 5525 956
rect 5529 916 5531 956
rect 5574 876 5576 956
rect 5580 876 5584 956
rect 5588 876 5590 956
rect 5602 916 5606 956
rect 5610 916 5612 956
rect 5669 916 5671 956
rect 5675 916 5677 956
rect 5689 916 5691 956
rect 5695 916 5697 956
rect 5754 876 5756 956
rect 5760 876 5764 956
rect 5768 876 5770 956
rect 5782 916 5786 956
rect 5790 916 5792 956
rect 5863 916 5865 956
rect 5869 920 5871 956
rect 5883 920 5885 956
rect 5869 916 5885 920
rect 5889 916 5891 956
rect 5903 916 5905 956
rect 5909 916 5911 956
rect 5953 876 5955 956
rect 5959 916 5961 956
rect 5973 916 5975 956
rect 5979 916 5989 956
rect 5993 916 5995 956
rect 6007 916 6009 956
rect 6013 916 6021 956
rect 6025 916 6027 956
rect 6039 916 6041 956
rect 6045 916 6047 956
rect 6085 916 6087 956
rect 6091 916 6095 956
rect 6099 936 6101 956
rect 6113 936 6115 956
rect 6119 936 6123 956
rect 6127 936 6131 956
rect 6143 936 6145 956
rect 6099 916 6110 936
rect 5959 876 5968 916
rect 6136 876 6145 936
rect 6149 876 6151 956
rect 6194 876 6196 956
rect 6200 876 6204 956
rect 6208 876 6210 956
rect 6222 916 6226 956
rect 6230 916 6232 956
rect 6294 876 6296 956
rect 6300 876 6304 956
rect 6308 876 6310 956
rect 6322 916 6326 956
rect 6330 916 6332 956
rect 6403 916 6405 956
rect 6409 916 6411 956
rect 6423 916 6425 956
rect 6429 916 6431 956
rect 6473 876 6475 956
rect 6479 916 6481 956
rect 6493 916 6495 956
rect 6499 916 6509 956
rect 6513 916 6515 956
rect 6527 916 6529 956
rect 6533 916 6541 956
rect 6545 916 6547 956
rect 6559 916 6561 956
rect 6565 916 6567 956
rect 6605 916 6607 956
rect 6611 916 6615 956
rect 6619 936 6621 956
rect 6633 936 6635 956
rect 6639 936 6643 956
rect 6647 936 6651 956
rect 6663 936 6665 956
rect 6619 916 6630 936
rect 6479 876 6488 916
rect 6656 876 6665 936
rect 6669 876 6671 956
rect 157 576 171 584
rect 29 504 31 544
rect 35 504 37 544
rect 89 504 91 544
rect 95 504 97 544
rect 109 504 111 544
rect 115 504 117 544
rect 169 504 171 576
rect 175 572 191 584
rect 175 504 177 572
rect 189 504 191 572
rect 195 504 197 584
rect 209 504 211 584
rect 215 504 217 584
rect 269 504 271 544
rect 275 504 277 544
rect 343 504 345 584
rect 349 504 351 584
rect 363 504 365 584
rect 369 572 385 584
rect 369 504 371 572
rect 383 504 385 572
rect 389 576 403 584
rect 389 504 391 576
rect 429 504 431 544
rect 435 504 437 544
rect 449 504 451 544
rect 455 540 471 544
rect 455 504 457 540
rect 469 504 471 540
rect 475 504 477 544
rect 543 504 545 544
rect 549 504 551 544
rect 563 504 565 544
rect 569 504 571 544
rect 623 504 625 544
rect 629 540 645 544
rect 629 504 631 540
rect 643 504 645 540
rect 649 504 651 544
rect 663 504 665 544
rect 669 504 671 544
rect 709 504 711 544
rect 715 504 717 544
rect 769 504 771 544
rect 775 504 777 544
rect 855 504 857 584
rect 861 504 865 584
rect 869 504 871 584
rect 919 512 921 572
rect 925 568 941 572
rect 925 516 927 568
rect 939 516 941 568
rect 925 512 941 516
rect 945 512 947 572
rect 971 562 985 564
rect 983 504 985 562
rect 989 516 991 564
rect 1003 516 1005 564
rect 989 504 1005 516
rect 1009 504 1011 564
rect 1023 504 1025 564
rect 1029 504 1031 564
rect 1043 504 1045 564
rect 1049 504 1051 564
rect 1093 504 1095 584
rect 1099 544 1108 584
rect 1099 504 1101 544
rect 1113 504 1115 544
rect 1119 504 1129 544
rect 1133 504 1135 544
rect 1147 504 1149 544
rect 1153 504 1161 544
rect 1165 504 1167 544
rect 1179 504 1181 544
rect 1185 504 1187 544
rect 1225 504 1227 544
rect 1231 504 1235 544
rect 1239 524 1250 544
rect 1276 524 1285 584
rect 1239 504 1241 524
rect 1253 504 1255 524
rect 1259 504 1263 524
rect 1267 504 1271 524
rect 1283 504 1285 524
rect 1289 504 1291 584
rect 1329 504 1331 544
rect 1335 504 1339 544
rect 1351 504 1353 584
rect 1357 504 1359 584
rect 1409 504 1411 544
rect 1415 504 1417 544
rect 1429 504 1431 544
rect 1435 504 1437 544
rect 1493 504 1495 584
rect 1499 544 1508 584
rect 1499 504 1501 544
rect 1513 504 1515 544
rect 1519 504 1529 544
rect 1533 504 1535 544
rect 1547 504 1549 544
rect 1553 504 1561 544
rect 1565 504 1567 544
rect 1579 504 1581 544
rect 1585 504 1587 544
rect 1625 504 1627 544
rect 1631 504 1635 544
rect 1639 524 1650 544
rect 1676 524 1685 584
rect 1639 504 1641 524
rect 1653 504 1655 524
rect 1659 504 1663 524
rect 1667 504 1671 524
rect 1683 504 1685 524
rect 1689 504 1691 584
rect 1733 504 1735 584
rect 1739 544 1748 584
rect 1739 504 1741 544
rect 1753 504 1755 544
rect 1759 504 1769 544
rect 1773 504 1775 544
rect 1787 504 1789 544
rect 1793 504 1801 544
rect 1805 504 1807 544
rect 1819 504 1821 544
rect 1825 504 1827 544
rect 1865 504 1867 544
rect 1871 504 1875 544
rect 1879 524 1890 544
rect 1916 524 1925 584
rect 1879 504 1881 524
rect 1893 504 1895 524
rect 1899 504 1903 524
rect 1907 504 1911 524
rect 1923 504 1925 524
rect 1929 504 1931 584
rect 1973 504 1975 584
rect 1979 544 1988 584
rect 1979 504 1981 544
rect 1993 504 1995 544
rect 1999 504 2009 544
rect 2013 504 2015 544
rect 2027 504 2029 544
rect 2033 504 2041 544
rect 2045 504 2047 544
rect 2059 504 2061 544
rect 2065 504 2067 544
rect 2105 504 2107 544
rect 2111 504 2115 544
rect 2119 524 2130 544
rect 2156 524 2165 584
rect 2119 504 2121 524
rect 2133 504 2135 524
rect 2139 504 2143 524
rect 2147 504 2151 524
rect 2163 504 2165 524
rect 2169 504 2171 584
rect 2213 504 2215 584
rect 2219 544 2228 584
rect 2219 504 2221 544
rect 2233 504 2235 544
rect 2239 504 2249 544
rect 2253 504 2255 544
rect 2267 504 2269 544
rect 2273 504 2281 544
rect 2285 504 2287 544
rect 2299 504 2301 544
rect 2305 504 2307 544
rect 2345 504 2347 544
rect 2351 504 2355 544
rect 2359 524 2370 544
rect 2396 524 2405 584
rect 2359 504 2361 524
rect 2373 504 2375 524
rect 2379 504 2383 524
rect 2387 504 2391 524
rect 2403 504 2405 524
rect 2409 504 2411 584
rect 2449 504 2451 584
rect 2455 524 2464 584
rect 2632 544 2641 584
rect 2490 524 2501 544
rect 2455 504 2457 524
rect 2469 504 2473 524
rect 2477 504 2481 524
rect 2485 504 2487 524
rect 2499 504 2501 524
rect 2505 504 2509 544
rect 2513 504 2515 544
rect 2553 504 2555 544
rect 2559 504 2561 544
rect 2573 504 2575 544
rect 2579 504 2587 544
rect 2591 504 2593 544
rect 2605 504 2607 544
rect 2611 504 2621 544
rect 2625 504 2627 544
rect 2639 504 2641 544
rect 2645 504 2647 584
rect 2703 504 2705 584
rect 2709 516 2711 584
rect 2723 516 2725 584
rect 2709 504 2725 516
rect 2729 582 2745 584
rect 2729 504 2731 582
rect 2743 504 2745 582
rect 2749 570 2765 584
rect 2749 504 2751 570
rect 2763 504 2765 570
rect 2769 582 2783 584
rect 2769 504 2771 582
rect 2823 504 2825 544
rect 2829 504 2831 544
rect 2883 504 2885 584
rect 2889 504 2891 584
rect 2903 504 2905 584
rect 2909 572 2925 584
rect 2909 504 2911 572
rect 2923 504 2925 572
rect 2929 576 2943 584
rect 2929 504 2931 576
rect 2969 504 2971 544
rect 2975 504 2977 544
rect 3034 504 3036 584
rect 3040 504 3044 584
rect 3048 504 3050 584
rect 3062 504 3066 544
rect 3070 504 3072 544
rect 3129 504 3131 544
rect 3135 504 3137 544
rect 3149 504 3151 544
rect 3155 504 3157 544
rect 3209 504 3211 544
rect 3215 504 3217 544
rect 3229 504 3231 544
rect 3235 540 3251 544
rect 3235 504 3237 540
rect 3249 504 3251 540
rect 3255 504 3257 544
rect 3309 504 3311 544
rect 3315 504 3317 544
rect 3374 504 3376 584
rect 3380 504 3384 584
rect 3388 504 3390 584
rect 3537 576 3551 584
rect 3402 504 3406 544
rect 3410 504 3412 544
rect 3469 504 3471 544
rect 3475 504 3477 544
rect 3489 504 3491 544
rect 3495 504 3497 544
rect 3549 504 3551 576
rect 3555 572 3571 584
rect 3555 504 3557 572
rect 3569 504 3571 572
rect 3575 504 3577 584
rect 3589 504 3591 584
rect 3595 504 3597 584
rect 3649 504 3651 584
rect 3655 504 3659 584
rect 3663 504 3665 584
rect 3734 504 3736 584
rect 3740 504 3744 584
rect 3748 504 3750 584
rect 3762 504 3766 544
rect 3770 504 3772 544
rect 3843 504 3845 544
rect 3849 540 3865 544
rect 3849 504 3851 540
rect 3863 504 3865 540
rect 3869 504 3871 544
rect 3883 504 3885 544
rect 3889 504 3891 544
rect 3929 504 3931 584
rect 3935 524 3944 584
rect 4112 544 4121 584
rect 3970 524 3981 544
rect 3935 504 3937 524
rect 3949 504 3953 524
rect 3957 504 3961 524
rect 3965 504 3967 524
rect 3979 504 3981 524
rect 3985 504 3989 544
rect 3993 504 3995 544
rect 4033 504 4035 544
rect 4039 504 4041 544
rect 4053 504 4055 544
rect 4059 504 4067 544
rect 4071 504 4073 544
rect 4085 504 4087 544
rect 4091 504 4101 544
rect 4105 504 4107 544
rect 4119 504 4121 544
rect 4125 504 4127 584
rect 4195 504 4197 584
rect 4201 504 4205 584
rect 4209 504 4211 584
rect 4249 504 4251 584
rect 4255 524 4264 584
rect 4432 544 4441 584
rect 4290 524 4301 544
rect 4255 504 4257 524
rect 4269 504 4273 524
rect 4277 504 4281 524
rect 4285 504 4287 524
rect 4299 504 4301 524
rect 4305 504 4309 544
rect 4313 504 4315 544
rect 4353 504 4355 544
rect 4359 504 4361 544
rect 4373 504 4375 544
rect 4379 504 4387 544
rect 4391 504 4393 544
rect 4405 504 4407 544
rect 4411 504 4421 544
rect 4425 504 4427 544
rect 4439 504 4441 544
rect 4445 504 4447 584
rect 4537 582 4551 584
rect 4489 504 4491 544
rect 4495 504 4497 544
rect 4549 504 4551 582
rect 4555 570 4571 584
rect 4555 504 4557 570
rect 4569 504 4571 570
rect 4575 582 4591 584
rect 4575 504 4577 582
rect 4589 504 4591 582
rect 4595 516 4597 584
rect 4609 516 4611 584
rect 4595 504 4611 516
rect 4615 504 4617 584
rect 4683 504 4685 584
rect 4689 504 4691 584
rect 4703 504 4705 584
rect 4709 572 4725 584
rect 4709 504 4711 572
rect 4723 504 4725 572
rect 4729 576 4743 584
rect 4729 504 4731 576
rect 4788 504 4790 544
rect 4794 504 4798 544
rect 4810 504 4812 584
rect 4816 504 4820 584
rect 4824 504 4826 584
rect 5047 584 5055 592
rect 4869 504 4871 544
rect 4875 504 4877 544
rect 4889 504 4891 544
rect 4895 504 4897 544
rect 4963 504 4965 544
rect 4969 504 4971 544
rect 5023 504 5025 584
rect 5029 504 5035 584
rect 5039 576 5055 584
rect 5039 512 5041 576
rect 5053 512 5055 576
rect 5059 512 5065 592
rect 5069 552 5079 592
rect 5069 512 5071 552
rect 5083 512 5085 552
rect 5089 512 5091 552
rect 5039 504 5048 512
rect 5129 504 5131 544
rect 5135 504 5137 544
rect 5149 504 5151 544
rect 5155 540 5171 544
rect 5155 504 5157 540
rect 5169 504 5171 540
rect 5175 504 5177 544
rect 5229 504 5231 584
rect 5235 524 5244 584
rect 5412 544 5421 584
rect 5270 524 5281 544
rect 5235 504 5237 524
rect 5249 504 5253 524
rect 5257 504 5261 524
rect 5265 504 5267 524
rect 5279 504 5281 524
rect 5285 504 5289 544
rect 5293 504 5295 544
rect 5333 504 5335 544
rect 5339 504 5341 544
rect 5353 504 5355 544
rect 5359 504 5367 544
rect 5371 504 5373 544
rect 5385 504 5387 544
rect 5391 504 5401 544
rect 5405 504 5407 544
rect 5419 504 5421 544
rect 5425 504 5427 584
rect 5469 504 5471 584
rect 5475 504 5477 584
rect 5541 552 5551 592
rect 5529 512 5531 552
rect 5535 512 5537 552
rect 5549 512 5551 552
rect 5555 512 5561 592
rect 5565 584 5573 592
rect 5565 576 5581 584
rect 5565 512 5567 576
rect 5579 512 5581 576
rect 5572 504 5581 512
rect 5585 504 5591 584
rect 5595 504 5597 584
rect 5675 504 5677 584
rect 5681 504 5685 584
rect 5689 504 5691 584
rect 5755 504 5757 584
rect 5761 504 5765 584
rect 5769 504 5771 584
rect 5835 504 5837 584
rect 5841 504 5845 584
rect 5849 504 5851 584
rect 5889 504 5891 584
rect 5895 504 5899 584
rect 5903 504 5905 584
rect 5995 504 5997 584
rect 6001 504 6005 584
rect 6009 504 6011 584
rect 6054 504 6056 584
rect 6060 504 6064 584
rect 6068 504 6070 584
rect 6082 504 6086 544
rect 6090 504 6092 544
rect 6154 504 6156 584
rect 6160 504 6164 584
rect 6168 504 6170 584
rect 6182 504 6186 544
rect 6190 504 6192 544
rect 6263 504 6265 544
rect 6269 504 6271 544
rect 6283 504 6285 544
rect 6289 504 6291 544
rect 6333 504 6335 584
rect 6339 544 6348 584
rect 6339 504 6341 544
rect 6353 504 6355 544
rect 6359 504 6369 544
rect 6373 504 6375 544
rect 6387 504 6389 544
rect 6393 504 6401 544
rect 6405 504 6407 544
rect 6419 504 6421 544
rect 6425 504 6427 544
rect 6465 504 6467 544
rect 6471 504 6475 544
rect 6479 524 6490 544
rect 6516 524 6525 584
rect 6479 504 6481 524
rect 6493 504 6495 524
rect 6499 504 6503 524
rect 6507 504 6511 524
rect 6523 504 6525 524
rect 6529 504 6531 584
rect 6569 504 6571 544
rect 6575 504 6577 544
rect 6629 504 6631 544
rect 6635 504 6637 544
rect 29 396 31 476
rect 35 456 37 476
rect 49 456 53 476
rect 57 456 61 476
rect 65 456 67 476
rect 79 456 81 476
rect 35 396 44 456
rect 70 436 81 456
rect 85 436 89 476
rect 93 436 95 476
rect 133 436 135 476
rect 139 436 141 476
rect 153 436 155 476
rect 159 436 167 476
rect 171 436 173 476
rect 185 436 187 476
rect 191 436 201 476
rect 205 436 207 476
rect 219 436 221 476
rect 212 396 221 436
rect 225 396 227 476
rect 273 396 275 476
rect 279 436 281 476
rect 293 436 295 476
rect 299 436 309 476
rect 313 436 315 476
rect 327 436 329 476
rect 333 436 341 476
rect 345 436 347 476
rect 359 436 361 476
rect 365 436 367 476
rect 405 436 407 476
rect 411 436 415 476
rect 419 456 421 476
rect 433 456 435 476
rect 439 456 443 476
rect 447 456 451 476
rect 463 456 465 476
rect 419 436 430 456
rect 279 396 288 436
rect 456 396 465 456
rect 469 396 471 476
rect 509 436 511 476
rect 515 436 517 476
rect 529 436 531 476
rect 535 440 537 476
rect 549 440 551 476
rect 535 436 551 440
rect 555 436 557 476
rect 609 396 611 476
rect 615 396 619 476
rect 623 396 625 476
rect 715 396 717 476
rect 721 396 725 476
rect 729 396 731 476
rect 769 436 771 476
rect 775 436 777 476
rect 789 436 791 476
rect 795 436 797 476
rect 863 436 865 476
rect 869 436 871 476
rect 913 396 915 476
rect 919 436 921 476
rect 933 436 935 476
rect 939 436 949 476
rect 953 436 955 476
rect 967 436 969 476
rect 973 436 981 476
rect 985 436 987 476
rect 999 436 1001 476
rect 1005 436 1007 476
rect 1045 436 1047 476
rect 1051 436 1055 476
rect 1059 456 1061 476
rect 1073 456 1075 476
rect 1079 456 1083 476
rect 1087 456 1091 476
rect 1103 456 1105 476
rect 1059 436 1070 456
rect 919 396 928 436
rect 1096 396 1105 456
rect 1109 396 1111 476
rect 1161 396 1163 476
rect 1167 396 1169 476
rect 1181 436 1185 476
rect 1189 436 1191 476
rect 1229 436 1231 476
rect 1235 436 1239 476
rect 1251 396 1253 476
rect 1257 396 1259 476
rect 1309 436 1311 476
rect 1315 436 1319 476
rect 1331 396 1333 476
rect 1337 396 1339 476
rect 1403 436 1405 476
rect 1409 436 1411 476
rect 1454 396 1456 476
rect 1460 396 1464 476
rect 1468 396 1470 476
rect 1482 436 1486 476
rect 1490 436 1492 476
rect 1563 436 1565 476
rect 1569 436 1571 476
rect 1614 396 1616 476
rect 1620 396 1624 476
rect 1628 396 1630 476
rect 1642 436 1646 476
rect 1650 436 1652 476
rect 1713 396 1715 476
rect 1719 436 1721 476
rect 1733 436 1735 476
rect 1739 436 1749 476
rect 1753 436 1755 476
rect 1767 436 1769 476
rect 1773 436 1781 476
rect 1785 436 1787 476
rect 1799 436 1801 476
rect 1805 436 1807 476
rect 1845 436 1847 476
rect 1851 436 1855 476
rect 1859 456 1861 476
rect 1873 456 1875 476
rect 1879 456 1883 476
rect 1887 456 1891 476
rect 1903 456 1905 476
rect 1859 436 1870 456
rect 1719 396 1728 436
rect 1896 396 1905 456
rect 1909 396 1911 476
rect 1963 436 1965 476
rect 1969 436 1971 476
rect 2023 436 2025 476
rect 2029 436 2031 476
rect 2074 396 2076 476
rect 2080 396 2084 476
rect 2088 396 2090 476
rect 2102 436 2106 476
rect 2110 436 2112 476
rect 2169 436 2171 476
rect 2175 436 2177 476
rect 2229 396 2231 476
rect 2235 396 2241 476
rect 2245 396 2247 476
rect 2269 396 2271 476
rect 2275 396 2281 476
rect 2285 396 2287 476
rect 2368 436 2370 476
rect 2374 436 2378 476
rect 2390 396 2392 476
rect 2396 396 2400 476
rect 2404 396 2406 476
rect 2449 396 2451 476
rect 2455 396 2459 476
rect 2463 396 2465 476
rect 2533 396 2535 476
rect 2539 436 2541 476
rect 2553 436 2555 476
rect 2559 436 2569 476
rect 2573 436 2575 476
rect 2587 436 2589 476
rect 2593 436 2601 476
rect 2605 436 2607 476
rect 2619 436 2621 476
rect 2625 436 2627 476
rect 2665 436 2667 476
rect 2671 436 2675 476
rect 2679 456 2681 476
rect 2693 456 2695 476
rect 2699 456 2703 476
rect 2707 456 2711 476
rect 2723 456 2725 476
rect 2679 436 2690 456
rect 2539 396 2548 436
rect 2716 396 2725 456
rect 2729 396 2731 476
rect 2788 436 2790 476
rect 2794 436 2798 476
rect 2810 396 2812 476
rect 2816 396 2820 476
rect 2824 396 2826 476
rect 2869 396 2871 476
rect 2875 396 2879 476
rect 2883 396 2885 476
rect 2953 396 2955 476
rect 2959 436 2961 476
rect 2973 436 2975 476
rect 2979 436 2989 476
rect 2993 436 2995 476
rect 3007 436 3009 476
rect 3013 436 3021 476
rect 3025 436 3027 476
rect 3039 436 3041 476
rect 3045 436 3047 476
rect 3085 436 3087 476
rect 3091 436 3095 476
rect 3099 456 3101 476
rect 3113 456 3115 476
rect 3119 456 3123 476
rect 3127 456 3131 476
rect 3143 456 3145 476
rect 3099 436 3110 456
rect 2959 396 2968 436
rect 3136 396 3145 456
rect 3149 396 3151 476
rect 3189 436 3191 476
rect 3195 436 3197 476
rect 3209 436 3211 476
rect 3215 436 3217 476
rect 3288 436 3290 476
rect 3294 436 3298 476
rect 3310 396 3312 476
rect 3316 396 3320 476
rect 3324 396 3326 476
rect 3369 396 3371 476
rect 3375 396 3379 476
rect 3383 396 3385 476
rect 3463 396 3465 476
rect 3469 396 3471 476
rect 3483 396 3485 476
rect 3489 408 3491 476
rect 3503 408 3505 476
rect 3489 396 3505 408
rect 3509 404 3511 476
rect 3509 396 3523 404
rect 3554 396 3556 476
rect 3560 396 3564 476
rect 3568 396 3570 476
rect 3582 436 3586 476
rect 3590 436 3592 476
rect 3649 396 3651 476
rect 3655 396 3659 476
rect 3663 396 3665 476
rect 3729 404 3731 476
rect 3717 396 3731 404
rect 3735 408 3737 476
rect 3749 408 3751 476
rect 3735 396 3751 408
rect 3755 396 3757 476
rect 3769 396 3771 476
rect 3775 396 3777 476
rect 3855 396 3857 476
rect 3861 396 3865 476
rect 3869 396 3871 476
rect 3914 396 3916 476
rect 3920 396 3924 476
rect 3928 396 3930 476
rect 3942 436 3946 476
rect 3950 436 3952 476
rect 4023 436 4025 476
rect 4029 440 4031 476
rect 4043 440 4045 476
rect 4029 436 4045 440
rect 4049 436 4051 476
rect 4063 436 4065 476
rect 4069 436 4071 476
rect 4109 396 4111 476
rect 4115 396 4119 476
rect 4123 396 4125 476
rect 4189 396 4191 476
rect 4195 456 4197 476
rect 4209 456 4213 476
rect 4217 456 4221 476
rect 4225 456 4227 476
rect 4239 456 4241 476
rect 4195 396 4204 456
rect 4230 436 4241 456
rect 4245 436 4249 476
rect 4253 436 4255 476
rect 4293 436 4295 476
rect 4299 436 4301 476
rect 4313 436 4315 476
rect 4319 436 4327 476
rect 4331 436 4333 476
rect 4345 436 4347 476
rect 4351 436 4361 476
rect 4365 436 4367 476
rect 4379 436 4381 476
rect 4372 396 4381 436
rect 4385 396 4387 476
rect 4429 396 4431 476
rect 4435 396 4439 476
rect 4443 396 4445 476
rect 4528 436 4530 476
rect 4534 436 4538 476
rect 4550 396 4552 476
rect 4556 396 4560 476
rect 4564 396 4566 476
rect 4609 396 4611 476
rect 4615 396 4619 476
rect 4623 396 4625 476
rect 4713 396 4715 476
rect 4719 396 4725 476
rect 4729 396 4731 476
rect 4753 396 4755 476
rect 4759 396 4765 476
rect 4769 396 4771 476
rect 4823 436 4825 476
rect 4829 436 4831 476
rect 4873 396 4875 476
rect 4879 436 4881 476
rect 4893 436 4895 476
rect 4899 436 4909 476
rect 4913 436 4915 476
rect 4927 436 4929 476
rect 4933 436 4941 476
rect 4945 436 4947 476
rect 4959 436 4961 476
rect 4965 436 4967 476
rect 5005 436 5007 476
rect 5011 436 5015 476
rect 5019 456 5021 476
rect 5033 456 5035 476
rect 5039 456 5043 476
rect 5047 456 5051 476
rect 5063 456 5065 476
rect 5019 436 5030 456
rect 4879 396 4888 436
rect 5056 396 5065 456
rect 5069 396 5071 476
rect 5123 396 5125 476
rect 5129 396 5131 476
rect 5143 396 5145 476
rect 5149 408 5151 476
rect 5163 408 5165 476
rect 5149 396 5165 408
rect 5169 404 5171 476
rect 5169 396 5183 404
rect 5209 396 5211 476
rect 5215 396 5219 476
rect 5223 396 5225 476
rect 5308 436 5310 476
rect 5314 436 5318 476
rect 5330 396 5332 476
rect 5336 396 5340 476
rect 5344 396 5346 476
rect 5389 396 5391 476
rect 5395 396 5399 476
rect 5403 396 5405 476
rect 5469 404 5471 476
rect 5457 396 5471 404
rect 5475 408 5477 476
rect 5489 408 5491 476
rect 5475 396 5491 408
rect 5495 396 5497 476
rect 5509 396 5511 476
rect 5515 396 5517 476
rect 5569 436 5571 476
rect 5575 436 5577 476
rect 5589 436 5591 476
rect 5595 440 5597 476
rect 5609 440 5611 476
rect 5595 436 5611 440
rect 5615 436 5617 476
rect 5674 396 5676 476
rect 5680 396 5684 476
rect 5688 396 5690 476
rect 5702 436 5706 476
rect 5710 436 5712 476
rect 5783 436 5785 476
rect 5789 436 5791 476
rect 5803 436 5805 476
rect 5809 436 5811 476
rect 5868 436 5870 476
rect 5874 436 5878 476
rect 5890 396 5892 476
rect 5896 396 5900 476
rect 5904 396 5906 476
rect 5954 396 5956 476
rect 5960 396 5964 476
rect 5968 396 5970 476
rect 5982 436 5986 476
rect 5990 436 5992 476
rect 6054 396 6056 476
rect 6060 396 6064 476
rect 6068 396 6070 476
rect 6082 436 6086 476
rect 6090 436 6092 476
rect 6175 396 6177 476
rect 6181 396 6185 476
rect 6189 396 6191 476
rect 6255 396 6257 476
rect 6261 396 6265 476
rect 6269 396 6271 476
rect 6333 396 6335 476
rect 6339 396 6345 476
rect 6349 396 6351 476
rect 6373 396 6375 476
rect 6379 396 6385 476
rect 6389 396 6391 476
rect 6433 396 6435 476
rect 6439 436 6441 476
rect 6453 436 6455 476
rect 6459 436 6469 476
rect 6473 436 6475 476
rect 6487 436 6489 476
rect 6493 436 6501 476
rect 6505 436 6507 476
rect 6519 436 6521 476
rect 6525 436 6527 476
rect 6565 436 6567 476
rect 6571 436 6575 476
rect 6579 456 6581 476
rect 6593 456 6595 476
rect 6599 456 6603 476
rect 6607 456 6611 476
rect 6623 456 6625 476
rect 6579 436 6590 456
rect 6439 396 6448 436
rect 6616 396 6625 456
rect 6629 396 6631 476
rect 29 24 31 104
rect 35 44 44 104
rect 212 64 221 104
rect 70 44 81 64
rect 35 24 37 44
rect 49 24 53 44
rect 57 24 61 44
rect 65 24 67 44
rect 79 24 81 44
rect 85 24 89 64
rect 93 24 95 64
rect 133 24 135 64
rect 139 24 141 64
rect 153 24 155 64
rect 159 24 167 64
rect 171 24 173 64
rect 185 24 187 64
rect 191 24 201 64
rect 205 24 207 64
rect 219 24 221 64
rect 225 24 227 104
rect 269 24 271 104
rect 275 44 284 104
rect 452 64 461 104
rect 310 44 321 64
rect 275 24 277 44
rect 289 24 293 44
rect 297 24 301 44
rect 305 24 307 44
rect 319 24 321 44
rect 325 24 329 64
rect 333 24 335 64
rect 373 24 375 64
rect 379 24 381 64
rect 393 24 395 64
rect 399 24 407 64
rect 411 24 413 64
rect 425 24 427 64
rect 431 24 441 64
rect 445 24 447 64
rect 459 24 461 64
rect 465 24 467 104
rect 521 24 523 104
rect 527 24 529 104
rect 541 24 545 64
rect 549 24 551 64
rect 589 24 591 64
rect 595 24 599 64
rect 611 24 613 104
rect 617 24 619 104
rect 681 24 683 104
rect 687 24 689 104
rect 701 24 705 64
rect 709 24 711 64
rect 749 24 751 104
rect 755 44 764 104
rect 932 64 941 104
rect 790 44 801 64
rect 755 24 757 44
rect 769 24 773 44
rect 777 24 781 44
rect 785 24 787 44
rect 799 24 801 44
rect 805 24 809 64
rect 813 24 815 64
rect 853 24 855 64
rect 859 24 861 64
rect 873 24 875 64
rect 879 24 887 64
rect 891 24 893 64
rect 905 24 907 64
rect 911 24 921 64
rect 925 24 927 64
rect 939 24 941 64
rect 945 24 947 104
rect 989 24 991 64
rect 995 24 999 64
rect 1011 24 1013 104
rect 1017 24 1019 104
rect 1083 24 1085 64
rect 1089 24 1091 64
rect 1103 24 1105 64
rect 1109 24 1111 64
rect 1168 24 1170 64
rect 1174 24 1178 64
rect 1190 24 1192 104
rect 1196 24 1200 104
rect 1204 24 1206 104
rect 1253 24 1255 104
rect 1259 64 1268 104
rect 1259 24 1261 64
rect 1273 24 1275 64
rect 1279 24 1289 64
rect 1293 24 1295 64
rect 1307 24 1309 64
rect 1313 24 1321 64
rect 1325 24 1327 64
rect 1339 24 1341 64
rect 1345 24 1347 64
rect 1385 24 1387 64
rect 1391 24 1395 64
rect 1399 44 1410 64
rect 1436 44 1445 104
rect 1399 24 1401 44
rect 1413 24 1415 44
rect 1419 24 1423 44
rect 1427 24 1431 44
rect 1443 24 1445 44
rect 1449 24 1451 104
rect 1503 24 1505 64
rect 1509 24 1511 64
rect 1549 24 1551 64
rect 1555 24 1557 64
rect 1569 24 1571 64
rect 1575 24 1577 64
rect 1648 24 1650 64
rect 1654 24 1658 64
rect 1670 24 1672 104
rect 1676 24 1680 104
rect 1684 24 1686 104
rect 1729 24 1731 64
rect 1735 24 1737 64
rect 1789 24 1791 64
rect 1795 24 1797 64
rect 1809 24 1811 64
rect 1815 24 1817 64
rect 1869 24 1871 64
rect 1875 24 1877 64
rect 1889 24 1891 64
rect 1895 24 1897 64
rect 1949 24 1951 64
rect 1955 24 1957 64
rect 1969 24 1971 64
rect 1975 24 1977 64
rect 2048 24 2050 64
rect 2054 24 2058 64
rect 2070 24 2072 104
rect 2076 24 2080 104
rect 2084 24 2086 104
rect 2133 24 2135 104
rect 2139 64 2148 104
rect 2139 24 2141 64
rect 2153 24 2155 64
rect 2159 24 2169 64
rect 2173 24 2175 64
rect 2187 24 2189 64
rect 2193 24 2201 64
rect 2205 24 2207 64
rect 2219 24 2221 64
rect 2225 24 2227 64
rect 2265 24 2267 64
rect 2271 24 2275 64
rect 2279 44 2290 64
rect 2316 44 2325 104
rect 2279 24 2281 44
rect 2293 24 2295 44
rect 2299 24 2303 44
rect 2307 24 2311 44
rect 2323 24 2325 44
rect 2329 24 2331 104
rect 2369 24 2371 64
rect 2375 24 2377 64
rect 2389 24 2391 64
rect 2395 24 2397 64
rect 2463 24 2465 64
rect 2469 24 2471 64
rect 2483 24 2485 64
rect 2489 24 2491 64
rect 2548 24 2550 64
rect 2554 24 2558 64
rect 2570 24 2572 104
rect 2576 24 2580 104
rect 2584 24 2586 104
rect 2643 24 2645 64
rect 2649 24 2651 64
rect 2693 24 2695 104
rect 2699 64 2708 104
rect 2699 24 2701 64
rect 2713 24 2715 64
rect 2719 24 2729 64
rect 2733 24 2735 64
rect 2747 24 2749 64
rect 2753 24 2761 64
rect 2765 24 2767 64
rect 2779 24 2781 64
rect 2785 24 2787 64
rect 2825 24 2827 64
rect 2831 24 2835 64
rect 2839 44 2850 64
rect 2876 44 2885 104
rect 2839 24 2841 44
rect 2853 24 2855 44
rect 2859 24 2863 44
rect 2867 24 2871 44
rect 2883 24 2885 44
rect 2889 24 2891 104
rect 2948 24 2950 64
rect 2954 24 2958 64
rect 2970 24 2972 104
rect 2976 24 2980 104
rect 2984 24 2986 104
rect 3055 24 3057 104
rect 3061 24 3065 104
rect 3069 24 3071 104
rect 3133 24 3135 104
rect 3139 24 3145 104
rect 3149 24 3151 104
rect 3173 24 3175 104
rect 3179 24 3185 104
rect 3189 24 3191 104
rect 3243 24 3245 64
rect 3249 24 3251 64
rect 3289 24 3291 104
rect 3295 44 3304 104
rect 3472 64 3481 104
rect 3330 44 3341 64
rect 3295 24 3297 44
rect 3309 24 3313 44
rect 3317 24 3321 44
rect 3325 24 3327 44
rect 3339 24 3341 44
rect 3345 24 3349 64
rect 3353 24 3355 64
rect 3393 24 3395 64
rect 3399 24 3401 64
rect 3413 24 3415 64
rect 3419 24 3427 64
rect 3431 24 3433 64
rect 3445 24 3447 64
rect 3451 24 3461 64
rect 3465 24 3467 64
rect 3479 24 3481 64
rect 3485 24 3487 104
rect 3543 24 3545 64
rect 3549 24 3551 64
rect 3563 24 3565 64
rect 3569 24 3571 64
rect 3628 24 3630 64
rect 3634 24 3638 64
rect 3650 24 3652 104
rect 3656 24 3660 104
rect 3664 24 3666 104
rect 3714 24 3716 104
rect 3720 24 3724 104
rect 3728 24 3730 104
rect 3742 24 3746 64
rect 3750 24 3752 64
rect 3809 24 3811 104
rect 3815 44 3824 104
rect 3992 64 4001 104
rect 3850 44 3861 64
rect 3815 24 3817 44
rect 3829 24 3833 44
rect 3837 24 3841 44
rect 3845 24 3847 44
rect 3859 24 3861 44
rect 3865 24 3869 64
rect 3873 24 3875 64
rect 3913 24 3915 64
rect 3919 24 3921 64
rect 3933 24 3935 64
rect 3939 24 3947 64
rect 3951 24 3953 64
rect 3965 24 3967 64
rect 3971 24 3981 64
rect 3985 24 3987 64
rect 3999 24 4001 64
rect 4005 24 4007 104
rect 4054 24 4056 104
rect 4060 24 4064 104
rect 4068 24 4070 104
rect 4082 24 4086 64
rect 4090 24 4092 64
rect 4154 24 4156 104
rect 4160 24 4164 104
rect 4168 24 4170 104
rect 4182 24 4186 64
rect 4190 24 4192 64
rect 4249 24 4251 64
rect 4255 24 4257 64
rect 4269 24 4271 64
rect 4275 24 4277 64
rect 4329 24 4331 104
rect 4335 44 4344 104
rect 4512 64 4521 104
rect 4370 44 4381 64
rect 4335 24 4337 44
rect 4349 24 4353 44
rect 4357 24 4361 44
rect 4365 24 4367 44
rect 4379 24 4381 44
rect 4385 24 4389 64
rect 4393 24 4395 64
rect 4433 24 4435 64
rect 4439 24 4441 64
rect 4453 24 4455 64
rect 4459 24 4467 64
rect 4471 24 4473 64
rect 4485 24 4487 64
rect 4491 24 4501 64
rect 4505 24 4507 64
rect 4519 24 4521 64
rect 4525 24 4527 104
rect 4574 24 4576 104
rect 4580 24 4584 104
rect 4588 24 4590 104
rect 4602 24 4606 64
rect 4610 24 4612 64
rect 4674 24 4676 104
rect 4680 24 4684 104
rect 4688 24 4690 104
rect 4702 24 4706 64
rect 4710 24 4712 64
rect 4769 24 4771 64
rect 4775 24 4777 64
rect 4789 24 4791 64
rect 4795 24 4797 64
rect 4849 24 4851 104
rect 4855 44 4864 104
rect 5032 64 5041 104
rect 4890 44 4901 64
rect 4855 24 4857 44
rect 4869 24 4873 44
rect 4877 24 4881 44
rect 4885 24 4887 44
rect 4899 24 4901 44
rect 4905 24 4909 64
rect 4913 24 4915 64
rect 4953 24 4955 64
rect 4959 24 4961 64
rect 4973 24 4975 64
rect 4979 24 4987 64
rect 4991 24 4993 64
rect 5005 24 5007 64
rect 5011 24 5021 64
rect 5025 24 5027 64
rect 5039 24 5041 64
rect 5045 24 5047 104
rect 5108 24 5110 64
rect 5114 24 5118 64
rect 5130 24 5132 104
rect 5136 24 5140 104
rect 5144 24 5146 104
rect 5194 24 5196 104
rect 5200 24 5204 104
rect 5208 24 5210 104
rect 5222 24 5226 64
rect 5230 24 5232 64
rect 5289 24 5291 64
rect 5295 24 5297 64
rect 5309 24 5311 64
rect 5315 24 5317 64
rect 5369 24 5371 104
rect 5375 44 5384 104
rect 5552 64 5561 104
rect 5410 44 5421 64
rect 5375 24 5377 44
rect 5389 24 5393 44
rect 5397 24 5401 44
rect 5405 24 5407 44
rect 5419 24 5421 44
rect 5425 24 5429 64
rect 5433 24 5435 64
rect 5473 24 5475 64
rect 5479 24 5481 64
rect 5493 24 5495 64
rect 5499 24 5507 64
rect 5511 24 5513 64
rect 5525 24 5527 64
rect 5531 24 5541 64
rect 5545 24 5547 64
rect 5559 24 5561 64
rect 5565 24 5567 104
rect 5609 24 5611 104
rect 5615 44 5624 104
rect 5792 64 5801 104
rect 5650 44 5661 64
rect 5615 24 5617 44
rect 5629 24 5633 44
rect 5637 24 5641 44
rect 5645 24 5647 44
rect 5659 24 5661 44
rect 5665 24 5669 64
rect 5673 24 5675 64
rect 5713 24 5715 64
rect 5719 24 5721 64
rect 5733 24 5735 64
rect 5739 24 5747 64
rect 5751 24 5753 64
rect 5765 24 5767 64
rect 5771 24 5781 64
rect 5785 24 5787 64
rect 5799 24 5801 64
rect 5805 24 5807 104
rect 5849 24 5851 104
rect 5855 44 5864 104
rect 6032 64 6041 104
rect 5890 44 5901 64
rect 5855 24 5857 44
rect 5869 24 5873 44
rect 5877 24 5881 44
rect 5885 24 5887 44
rect 5899 24 5901 44
rect 5905 24 5909 64
rect 5913 24 5915 64
rect 5953 24 5955 64
rect 5959 24 5961 64
rect 5973 24 5975 64
rect 5979 24 5987 64
rect 5991 24 5993 64
rect 6005 24 6007 64
rect 6011 24 6021 64
rect 6025 24 6027 64
rect 6039 24 6041 64
rect 6045 24 6047 104
rect 6103 24 6105 104
rect 6109 24 6111 104
rect 6154 24 6156 104
rect 6160 24 6164 104
rect 6168 24 6170 104
rect 6182 24 6186 64
rect 6190 24 6192 64
rect 6273 24 6275 104
rect 6279 24 6285 104
rect 6289 24 6291 104
rect 6313 24 6315 104
rect 6319 24 6325 104
rect 6329 24 6331 104
rect 6383 24 6385 64
rect 6389 24 6391 64
rect 6429 24 6431 104
rect 6435 44 6444 104
rect 6612 64 6621 104
rect 6470 44 6481 64
rect 6435 24 6437 44
rect 6449 24 6453 44
rect 6457 24 6461 44
rect 6465 24 6467 44
rect 6479 24 6481 44
rect 6485 24 6489 64
rect 6493 24 6495 64
rect 6533 24 6535 64
rect 6539 24 6541 64
rect 6553 24 6555 64
rect 6559 24 6567 64
rect 6571 24 6573 64
rect 6585 24 6587 64
rect 6591 24 6601 64
rect 6605 24 6607 64
rect 6619 24 6621 64
rect 6625 24 6627 104
<< ndcontact >>
rect 21 6436 33 6476
rect 41 6456 53 6476
rect 73 6456 85 6476
rect 103 6456 115 6476
rect 125 6456 137 6476
rect 151 6456 163 6476
rect 179 6456 191 6476
rect 209 6456 221 6476
rect 231 6436 243 6476
rect 271 6436 283 6476
rect 291 6436 303 6476
rect 311 6448 323 6476
rect 331 6436 343 6476
rect 359 6436 371 6476
rect 389 6436 401 6476
rect 459 6436 471 6476
rect 489 6436 501 6476
rect 519 6436 531 6476
rect 549 6436 561 6476
rect 597 6436 609 6476
rect 619 6456 631 6476
rect 649 6456 661 6476
rect 677 6456 689 6476
rect 703 6456 715 6476
rect 725 6456 737 6476
rect 755 6456 767 6476
rect 787 6456 799 6476
rect 807 6436 819 6476
rect 837 6456 849 6476
rect 857 6456 869 6476
rect 900 6436 912 6476
rect 928 6436 940 6476
rect 956 6436 968 6476
rect 1031 6456 1043 6476
rect 1051 6456 1063 6476
rect 1077 6436 1089 6476
rect 1099 6456 1111 6476
rect 1129 6456 1141 6476
rect 1157 6456 1169 6476
rect 1183 6456 1195 6476
rect 1205 6456 1217 6476
rect 1235 6456 1247 6476
rect 1267 6456 1279 6476
rect 1287 6436 1299 6476
rect 1317 6436 1329 6476
rect 1337 6446 1349 6476
rect 1357 6436 1369 6476
rect 1377 6436 1389 6464
rect 1397 6436 1409 6476
rect 1451 6436 1463 6476
rect 1471 6436 1483 6476
rect 1491 6448 1503 6476
rect 1511 6436 1523 6476
rect 1561 6436 1573 6476
rect 1581 6436 1593 6476
rect 1611 6436 1623 6476
rect 1651 6456 1663 6476
rect 1671 6456 1683 6476
rect 1697 6436 1709 6476
rect 1719 6456 1731 6476
rect 1749 6456 1761 6476
rect 1777 6456 1789 6476
rect 1803 6456 1815 6476
rect 1825 6456 1837 6476
rect 1855 6456 1867 6476
rect 1887 6456 1899 6476
rect 1907 6436 1919 6476
rect 1937 6436 1949 6476
rect 1957 6448 1969 6476
rect 1977 6436 1989 6476
rect 1997 6436 2009 6476
rect 2039 6436 2051 6476
rect 2069 6436 2081 6476
rect 2131 6436 2143 6476
rect 2151 6436 2163 6476
rect 2171 6448 2183 6476
rect 2191 6436 2203 6476
rect 2238 6456 2250 6476
rect 2260 6436 2272 6476
rect 2288 6436 2300 6476
rect 2339 6436 2351 6476
rect 2369 6436 2381 6476
rect 2411 6456 2423 6476
rect 2431 6456 2443 6476
rect 2451 6456 2463 6476
rect 2477 6456 2489 6476
rect 2497 6456 2509 6476
rect 2517 6456 2529 6476
rect 2559 6436 2571 6476
rect 2589 6436 2601 6476
rect 2674 6418 2686 6476
rect 2710 6416 2722 6476
rect 2739 6436 2751 6476
rect 2769 6436 2781 6476
rect 2854 6418 2866 6476
rect 2890 6416 2902 6476
rect 2931 6436 2943 6476
rect 2951 6436 2963 6476
rect 2971 6448 2983 6476
rect 2991 6436 3003 6476
rect 3031 6436 3043 6476
rect 3051 6436 3063 6476
rect 3071 6448 3083 6476
rect 3091 6436 3103 6476
rect 3131 6456 3143 6476
rect 3151 6456 3163 6476
rect 3191 6456 3203 6476
rect 3211 6456 3223 6476
rect 3240 6436 3252 6476
rect 3268 6436 3280 6476
rect 3290 6456 3302 6476
rect 3337 6436 3349 6476
rect 3357 6448 3369 6476
rect 3377 6436 3389 6476
rect 3397 6436 3409 6476
rect 3458 6456 3470 6476
rect 3480 6436 3492 6476
rect 3508 6436 3520 6476
rect 3558 6456 3570 6476
rect 3580 6436 3592 6476
rect 3608 6436 3620 6476
rect 3638 6416 3650 6476
rect 3674 6418 3686 6476
rect 3751 6436 3763 6476
rect 3771 6436 3783 6476
rect 3791 6448 3803 6476
rect 3811 6436 3823 6476
rect 3837 6436 3849 6476
rect 3857 6448 3869 6476
rect 3877 6436 3889 6476
rect 3897 6436 3909 6476
rect 3937 6456 3949 6476
rect 3957 6456 3969 6476
rect 3999 6436 4011 6476
rect 4029 6436 4041 6476
rect 4101 6436 4113 6476
rect 4121 6436 4133 6476
rect 4151 6436 4163 6476
rect 4179 6436 4191 6476
rect 4209 6436 4221 6476
rect 4294 6418 4306 6476
rect 4330 6416 4342 6476
rect 4394 6418 4406 6476
rect 4430 6416 4442 6476
rect 4494 6418 4506 6476
rect 4530 6416 4542 6476
rect 4557 6456 4569 6476
rect 4577 6456 4589 6476
rect 4620 6436 4632 6476
rect 4648 6436 4660 6476
rect 4670 6456 4682 6476
rect 4720 6436 4732 6476
rect 4748 6436 4760 6476
rect 4770 6456 4782 6476
rect 4817 6436 4829 6476
rect 4837 6448 4849 6476
rect 4857 6436 4869 6476
rect 4877 6436 4889 6476
rect 4931 6436 4943 6476
rect 4951 6436 4963 6476
rect 4971 6448 4983 6476
rect 4991 6436 5003 6476
rect 5017 6436 5029 6476
rect 5037 6448 5049 6476
rect 5057 6436 5069 6476
rect 5077 6436 5089 6476
rect 5154 6418 5166 6476
rect 5190 6416 5202 6476
rect 5254 6418 5266 6476
rect 5290 6416 5302 6476
rect 5354 6418 5366 6476
rect 5390 6416 5402 6476
rect 5420 6436 5432 6476
rect 5448 6436 5460 6476
rect 5470 6456 5482 6476
rect 5538 6456 5550 6476
rect 5560 6436 5572 6476
rect 5588 6436 5600 6476
rect 5631 6456 5643 6476
rect 5651 6456 5663 6476
rect 5680 6436 5692 6476
rect 5708 6436 5720 6476
rect 5730 6456 5742 6476
rect 5778 6416 5790 6476
rect 5814 6418 5826 6476
rect 5898 6456 5910 6476
rect 5920 6436 5932 6476
rect 5948 6436 5960 6476
rect 5991 6456 6003 6476
rect 6011 6456 6023 6476
rect 6058 6456 6070 6476
rect 6080 6436 6092 6476
rect 6108 6436 6120 6476
rect 6151 6436 6163 6476
rect 6171 6436 6183 6476
rect 6191 6448 6203 6476
rect 6211 6436 6223 6476
rect 6258 6456 6270 6476
rect 6280 6436 6292 6476
rect 6308 6436 6320 6476
rect 6338 6416 6350 6476
rect 6374 6418 6386 6476
rect 6474 6418 6486 6476
rect 6510 6416 6522 6476
rect 6537 6456 6549 6476
rect 6557 6456 6569 6476
rect 6600 6436 6612 6476
rect 6628 6436 6640 6476
rect 6656 6436 6668 6476
rect 17 6024 29 6064
rect 39 6024 51 6044
rect 69 6024 81 6044
rect 97 6024 109 6044
rect 123 6024 135 6044
rect 145 6024 157 6044
rect 175 6024 187 6044
rect 207 6024 219 6044
rect 227 6024 239 6064
rect 278 6024 290 6044
rect 300 6024 312 6064
rect 328 6024 340 6064
rect 379 6024 391 6064
rect 409 6024 421 6064
rect 437 6024 449 6044
rect 457 6024 469 6044
rect 477 6024 489 6044
rect 539 6024 551 6064
rect 569 6024 581 6064
rect 597 6024 609 6064
rect 617 6024 629 6052
rect 637 6024 649 6064
rect 657 6024 669 6064
rect 711 6024 723 6064
rect 731 6024 743 6064
rect 751 6024 763 6052
rect 771 6024 783 6064
rect 797 6024 809 6044
rect 817 6024 829 6044
rect 837 6024 849 6044
rect 898 6024 910 6044
rect 920 6024 932 6064
rect 948 6024 960 6064
rect 977 6024 989 6044
rect 997 6024 1009 6044
rect 1017 6024 1029 6044
rect 1037 6024 1049 6064
rect 1091 6024 1103 6044
rect 1111 6024 1123 6044
rect 1137 6024 1149 6044
rect 1157 6024 1169 6044
rect 1177 6024 1189 6044
rect 1231 6024 1243 6064
rect 1251 6024 1263 6064
rect 1271 6024 1283 6052
rect 1291 6024 1303 6064
rect 1331 6024 1343 6044
rect 1351 6024 1363 6044
rect 1391 6024 1403 6044
rect 1411 6024 1423 6044
rect 1437 6024 1449 6044
rect 1457 6024 1469 6044
rect 1477 6024 1489 6044
rect 1517 6024 1529 6044
rect 1537 6024 1549 6044
rect 1557 6024 1569 6044
rect 1597 6024 1609 6044
rect 1617 6024 1629 6044
rect 1657 6024 1669 6044
rect 1677 6024 1689 6044
rect 1697 6024 1709 6044
rect 1737 6024 1749 6044
rect 1757 6024 1769 6044
rect 1777 6024 1789 6044
rect 1817 6024 1829 6064
rect 1837 6024 1849 6052
rect 1857 6024 1869 6064
rect 1877 6024 1889 6064
rect 1917 6024 1929 6044
rect 1937 6024 1949 6044
rect 1998 6024 2010 6044
rect 2020 6024 2032 6064
rect 2048 6024 2060 6064
rect 2077 6024 2089 6044
rect 2097 6024 2109 6044
rect 2151 6024 2163 6064
rect 2171 6024 2183 6064
rect 2191 6024 2203 6052
rect 2211 6024 2223 6064
rect 2237 6024 2249 6044
rect 2257 6024 2269 6044
rect 2311 6024 2323 6064
rect 2331 6024 2343 6064
rect 2351 6024 2363 6052
rect 2371 6024 2383 6064
rect 2434 6024 2446 6082
rect 2470 6024 2482 6084
rect 2518 6024 2530 6044
rect 2540 6024 2552 6064
rect 2568 6024 2580 6064
rect 2611 6024 2623 6044
rect 2631 6024 2643 6044
rect 2651 6024 2663 6044
rect 2714 6024 2726 6082
rect 2750 6024 2762 6084
rect 2812 6024 2824 6064
rect 2840 6024 2852 6064
rect 2868 6024 2880 6064
rect 2911 6024 2923 6044
rect 2931 6024 2943 6044
rect 2958 6024 2970 6084
rect 2994 6024 3006 6082
rect 3078 6024 3090 6044
rect 3100 6024 3112 6064
rect 3128 6024 3140 6064
rect 3194 6024 3206 6082
rect 3230 6024 3242 6084
rect 3278 6024 3290 6044
rect 3300 6024 3312 6064
rect 3328 6024 3340 6064
rect 3371 6024 3383 6044
rect 3391 6024 3403 6044
rect 3454 6024 3466 6082
rect 3490 6024 3502 6084
rect 3518 6024 3530 6084
rect 3554 6024 3566 6082
rect 3617 6024 3629 6044
rect 3637 6024 3649 6044
rect 3680 6024 3692 6064
rect 3708 6024 3720 6064
rect 3730 6024 3742 6044
rect 3799 6024 3811 6064
rect 3829 6024 3841 6064
rect 3859 6024 3871 6064
rect 3889 6024 3901 6064
rect 3951 6024 3963 6064
rect 3971 6024 3983 6064
rect 3991 6024 4003 6052
rect 4011 6024 4023 6064
rect 4037 6024 4049 6064
rect 4057 6024 4069 6052
rect 4077 6024 4089 6064
rect 4097 6024 4109 6064
rect 4151 6024 4163 6044
rect 4171 6024 4183 6044
rect 4191 6024 4203 6044
rect 4217 6024 4229 6044
rect 4237 6024 4249 6044
rect 4299 6024 4311 6064
rect 4329 6024 4341 6064
rect 4357 6024 4369 6064
rect 4387 6024 4399 6064
rect 4407 6024 4419 6064
rect 4471 6024 4483 6064
rect 4491 6024 4503 6064
rect 4511 6024 4523 6052
rect 4531 6024 4543 6064
rect 4578 6024 4590 6044
rect 4600 6024 4612 6064
rect 4628 6024 4640 6064
rect 4658 6024 4670 6084
rect 4694 6024 4706 6082
rect 4778 6024 4790 6044
rect 4800 6024 4812 6064
rect 4828 6024 4840 6064
rect 4894 6024 4906 6082
rect 4930 6024 4942 6084
rect 4958 6024 4970 6084
rect 4994 6024 5006 6082
rect 5071 6024 5083 6064
rect 5091 6024 5103 6064
rect 5111 6024 5123 6052
rect 5131 6024 5143 6064
rect 5179 6024 5191 6064
rect 5209 6024 5221 6064
rect 5237 6024 5249 6064
rect 5267 6024 5279 6064
rect 5287 6024 5299 6064
rect 5337 6024 5349 6064
rect 5357 6024 5369 6052
rect 5377 6024 5389 6064
rect 5397 6024 5409 6064
rect 5458 6024 5470 6044
rect 5480 6024 5492 6064
rect 5508 6024 5520 6064
rect 5574 6024 5586 6082
rect 5610 6024 5622 6084
rect 5638 6024 5650 6084
rect 5674 6024 5686 6082
rect 5758 6024 5770 6044
rect 5780 6024 5792 6064
rect 5808 6024 5820 6064
rect 5838 6024 5850 6084
rect 5874 6024 5886 6082
rect 5937 6024 5949 6064
rect 5957 6024 5969 6052
rect 5977 6024 5989 6064
rect 5997 6024 6009 6064
rect 6037 6024 6049 6064
rect 6057 6024 6069 6052
rect 6077 6024 6089 6064
rect 6097 6024 6109 6064
rect 6138 6024 6150 6084
rect 6174 6024 6186 6082
rect 6238 6024 6250 6084
rect 6274 6024 6286 6082
rect 6374 6024 6386 6082
rect 6410 6024 6422 6084
rect 6458 6024 6470 6044
rect 6480 6024 6492 6064
rect 6508 6024 6520 6064
rect 6537 6024 6549 6044
rect 6557 6024 6569 6044
rect 6597 6024 6609 6044
rect 6617 6024 6629 6044
rect 29 5956 41 5996
rect 49 5956 61 5996
rect 71 5976 83 5996
rect 99 5956 111 5996
rect 129 5956 141 5996
rect 179 5956 191 5996
rect 209 5956 221 5996
rect 278 5976 290 5996
rect 300 5956 312 5996
rect 328 5956 340 5996
rect 379 5956 391 5996
rect 409 5956 421 5996
rect 437 5976 449 5996
rect 457 5976 469 5996
rect 511 5976 523 5996
rect 531 5976 543 5996
rect 551 5976 563 5996
rect 577 5976 589 5996
rect 597 5976 609 5996
rect 617 5976 629 5996
rect 657 5956 669 5996
rect 677 5968 689 5996
rect 697 5956 709 5996
rect 717 5956 729 5996
rect 771 5976 783 5996
rect 791 5976 803 5996
rect 817 5976 829 5996
rect 837 5976 849 5996
rect 857 5976 869 5996
rect 919 5956 931 5996
rect 949 5956 961 5996
rect 991 5956 1003 5996
rect 1011 5956 1023 5996
rect 1031 5968 1043 5996
rect 1051 5956 1063 5996
rect 1077 5976 1089 5996
rect 1097 5976 1109 5996
rect 1117 5976 1129 5996
rect 1171 5976 1183 5996
rect 1191 5976 1203 5996
rect 1217 5956 1229 5996
rect 1239 5976 1251 5996
rect 1269 5976 1281 5996
rect 1297 5976 1309 5996
rect 1323 5976 1335 5996
rect 1345 5976 1357 5996
rect 1375 5976 1387 5996
rect 1407 5976 1419 5996
rect 1427 5956 1439 5996
rect 1459 5956 1471 5996
rect 1489 5956 1501 5996
rect 1574 5938 1586 5996
rect 1610 5936 1622 5996
rect 1651 5956 1663 5996
rect 1671 5956 1683 5996
rect 1691 5968 1703 5996
rect 1711 5956 1723 5996
rect 1751 5976 1763 5996
rect 1771 5976 1783 5996
rect 1791 5976 1803 5996
rect 1854 5938 1866 5996
rect 1890 5936 1902 5996
rect 1917 5976 1929 5996
rect 1937 5976 1949 5996
rect 1991 5956 2003 5996
rect 2011 5956 2023 5996
rect 2031 5968 2043 5996
rect 2051 5956 2063 5996
rect 2078 5936 2090 5996
rect 2114 5938 2126 5996
rect 2198 5976 2210 5996
rect 2220 5956 2232 5996
rect 2248 5956 2260 5996
rect 2277 5956 2289 5996
rect 2297 5968 2309 5996
rect 2317 5956 2329 5996
rect 2337 5956 2349 5996
rect 2399 5956 2411 5996
rect 2429 5956 2441 5996
rect 2494 5938 2506 5996
rect 2530 5936 2542 5996
rect 2578 5976 2590 5996
rect 2600 5956 2612 5996
rect 2628 5956 2640 5996
rect 2659 5956 2671 5996
rect 2689 5956 2701 5996
rect 2774 5938 2786 5996
rect 2810 5936 2822 5996
rect 2874 5938 2886 5996
rect 2910 5936 2922 5996
rect 2974 5938 2986 5996
rect 3010 5936 3022 5996
rect 3074 5938 3086 5996
rect 3110 5936 3122 5996
rect 3138 5936 3150 5996
rect 3174 5938 3186 5996
rect 3251 5956 3263 5996
rect 3271 5956 3283 5996
rect 3291 5968 3303 5996
rect 3311 5956 3323 5996
rect 3337 5956 3349 5996
rect 3357 5968 3369 5996
rect 3377 5956 3389 5996
rect 3397 5956 3409 5996
rect 3458 5976 3470 5996
rect 3480 5956 3492 5996
rect 3508 5956 3520 5996
rect 3551 5956 3563 5996
rect 3571 5956 3583 5996
rect 3591 5968 3603 5996
rect 3611 5956 3623 5996
rect 3674 5938 3686 5996
rect 3710 5936 3722 5996
rect 3740 5956 3752 5996
rect 3768 5956 3780 5996
rect 3790 5976 3802 5996
rect 3874 5938 3886 5996
rect 3910 5936 3922 5996
rect 3958 5976 3970 5996
rect 3980 5956 3992 5996
rect 4008 5956 4020 5996
rect 4074 5938 4086 5996
rect 4110 5936 4122 5996
rect 4158 5976 4170 5996
rect 4180 5956 4192 5996
rect 4208 5956 4220 5996
rect 4238 5936 4250 5996
rect 4274 5938 4286 5996
rect 4339 5956 4351 5996
rect 4369 5956 4381 5996
rect 4431 5956 4443 5996
rect 4451 5956 4463 5996
rect 4471 5968 4483 5996
rect 4491 5956 4503 5996
rect 4531 5976 4543 5996
rect 4551 5976 4563 5996
rect 4571 5976 4583 5996
rect 4597 5956 4609 5996
rect 4627 5956 4639 5996
rect 4647 5956 4659 5996
rect 4718 5976 4730 5996
rect 4740 5956 4752 5996
rect 4768 5956 4780 5996
rect 4799 5956 4811 5996
rect 4829 5956 4841 5996
rect 4891 5976 4903 5996
rect 4911 5976 4923 5996
rect 4974 5938 4986 5996
rect 5010 5936 5022 5996
rect 5040 5956 5052 5996
rect 5068 5956 5080 5996
rect 5090 5976 5102 5996
rect 5137 5956 5149 5996
rect 5157 5968 5169 5996
rect 5177 5956 5189 5996
rect 5197 5956 5209 5996
rect 5237 5956 5249 5996
rect 5257 5968 5269 5996
rect 5277 5956 5289 5996
rect 5297 5956 5309 5996
rect 5340 5956 5352 5996
rect 5368 5956 5380 5996
rect 5396 5956 5408 5996
rect 5479 5956 5491 5996
rect 5509 5956 5521 5996
rect 5537 5976 5549 5996
rect 5557 5976 5569 5996
rect 5634 5938 5646 5996
rect 5670 5936 5682 5996
rect 5700 5956 5712 5996
rect 5728 5956 5740 5996
rect 5750 5976 5762 5996
rect 5811 5956 5823 5996
rect 5831 5956 5843 5996
rect 5851 5968 5863 5996
rect 5871 5956 5883 5996
rect 5897 5956 5909 5996
rect 5917 5968 5929 5996
rect 5937 5956 5949 5996
rect 5957 5956 5969 5996
rect 6011 5956 6023 5996
rect 6031 5956 6043 5996
rect 6051 5968 6063 5996
rect 6071 5956 6083 5996
rect 6100 5956 6112 5996
rect 6128 5956 6140 5996
rect 6156 5956 6168 5996
rect 6239 5956 6251 5996
rect 6269 5956 6281 5996
rect 6297 5956 6309 5996
rect 6327 5956 6339 5996
rect 6347 5956 6359 5996
rect 6397 5956 6409 5996
rect 6417 5968 6429 5996
rect 6437 5956 6449 5996
rect 6457 5956 6469 5996
rect 6498 5936 6510 5996
rect 6534 5938 6546 5996
rect 6599 5956 6611 5996
rect 6629 5956 6641 5996
rect 29 5544 41 5584
rect 49 5544 61 5584
rect 71 5544 83 5564
rect 109 5544 121 5584
rect 129 5544 141 5584
rect 151 5544 163 5564
rect 177 5544 189 5584
rect 199 5544 211 5564
rect 229 5544 241 5564
rect 257 5544 269 5564
rect 283 5544 295 5564
rect 305 5544 317 5564
rect 335 5544 347 5564
rect 367 5544 379 5564
rect 387 5544 399 5584
rect 431 5544 443 5564
rect 451 5544 463 5564
rect 471 5544 483 5564
rect 500 5544 512 5584
rect 528 5544 540 5584
rect 550 5544 562 5564
rect 599 5544 611 5584
rect 629 5544 641 5584
rect 677 5544 689 5584
rect 707 5544 719 5584
rect 727 5544 739 5584
rect 779 5544 791 5584
rect 809 5544 821 5584
rect 859 5544 871 5584
rect 889 5544 901 5584
rect 937 5544 949 5564
rect 957 5544 969 5564
rect 977 5544 989 5564
rect 1017 5544 1029 5564
rect 1037 5544 1049 5564
rect 1077 5544 1089 5564
rect 1097 5544 1109 5564
rect 1117 5544 1129 5564
rect 1137 5544 1149 5584
rect 1177 5544 1189 5564
rect 1197 5544 1209 5564
rect 1217 5544 1229 5564
rect 1257 5544 1269 5564
rect 1277 5544 1289 5564
rect 1317 5544 1329 5564
rect 1337 5544 1349 5564
rect 1357 5544 1369 5564
rect 1397 5544 1409 5564
rect 1417 5544 1429 5564
rect 1457 5544 1469 5584
rect 1479 5544 1491 5564
rect 1509 5544 1521 5564
rect 1537 5544 1549 5564
rect 1563 5544 1575 5564
rect 1585 5544 1597 5564
rect 1615 5544 1627 5564
rect 1647 5544 1659 5564
rect 1667 5544 1679 5584
rect 1697 5544 1709 5584
rect 1717 5544 1729 5574
rect 1737 5544 1749 5584
rect 1757 5556 1769 5584
rect 1777 5544 1789 5584
rect 1831 5544 1843 5584
rect 1851 5544 1863 5584
rect 1871 5544 1883 5572
rect 1891 5544 1903 5584
rect 1939 5544 1951 5584
rect 1969 5544 1981 5584
rect 1997 5544 2009 5564
rect 2017 5544 2029 5564
rect 2078 5544 2090 5564
rect 2100 5544 2112 5584
rect 2128 5544 2140 5584
rect 2157 5544 2169 5564
rect 2177 5544 2189 5564
rect 2197 5544 2209 5564
rect 2239 5544 2251 5584
rect 2269 5544 2281 5584
rect 2391 5544 2403 5564
rect 2411 5544 2423 5564
rect 2431 5544 2443 5564
rect 2451 5544 2465 5564
rect 2519 5544 2531 5584
rect 2549 5544 2561 5584
rect 2614 5544 2626 5602
rect 2650 5544 2662 5604
rect 2714 5544 2726 5602
rect 2750 5544 2762 5604
rect 2779 5544 2791 5584
rect 2809 5544 2821 5584
rect 2857 5544 2869 5584
rect 2877 5544 2889 5572
rect 2897 5544 2909 5584
rect 2917 5544 2929 5584
rect 2994 5544 3006 5602
rect 3030 5544 3042 5604
rect 3060 5544 3072 5584
rect 3088 5544 3100 5584
rect 3110 5544 3122 5564
rect 3171 5544 3183 5584
rect 3191 5544 3203 5584
rect 3211 5544 3223 5572
rect 3231 5544 3243 5584
rect 3271 5544 3283 5564
rect 3291 5544 3303 5564
rect 3318 5544 3330 5604
rect 3354 5544 3366 5602
rect 3454 5544 3466 5602
rect 3490 5544 3502 5604
rect 3554 5544 3566 5602
rect 3590 5544 3602 5604
rect 3631 5544 3643 5564
rect 3651 5544 3663 5564
rect 3691 5544 3703 5584
rect 3711 5544 3723 5584
rect 3731 5544 3743 5572
rect 3751 5544 3763 5584
rect 3791 5544 3803 5564
rect 3811 5544 3823 5564
rect 3831 5544 3843 5564
rect 3857 5544 3869 5584
rect 3877 5544 3889 5572
rect 3897 5544 3909 5584
rect 3917 5544 3929 5584
rect 3971 5544 3983 5564
rect 3991 5544 4003 5564
rect 4052 5544 4064 5584
rect 4080 5544 4092 5584
rect 4108 5544 4120 5584
rect 4151 5544 4163 5584
rect 4171 5544 4183 5584
rect 4191 5544 4203 5572
rect 4211 5544 4223 5584
rect 4274 5544 4286 5602
rect 4310 5544 4322 5604
rect 4337 5544 4349 5564
rect 4357 5544 4369 5564
rect 4411 5544 4423 5584
rect 4431 5544 4443 5584
rect 4451 5544 4463 5572
rect 4471 5544 4483 5584
rect 4521 5544 4533 5584
rect 4541 5544 4553 5584
rect 4571 5544 4583 5584
rect 4599 5544 4611 5584
rect 4629 5544 4641 5584
rect 4691 5544 4703 5584
rect 4711 5544 4723 5584
rect 4731 5544 4743 5572
rect 4751 5544 4763 5584
rect 4777 5544 4789 5584
rect 4797 5544 4809 5572
rect 4817 5544 4829 5584
rect 4837 5544 4849 5584
rect 4914 5544 4926 5602
rect 4950 5544 4962 5604
rect 4980 5544 4992 5584
rect 5008 5544 5020 5584
rect 5030 5544 5042 5564
rect 5077 5544 5089 5584
rect 5097 5544 5109 5572
rect 5117 5544 5129 5584
rect 5137 5544 5149 5584
rect 5178 5544 5190 5604
rect 5214 5544 5226 5602
rect 5279 5544 5291 5584
rect 5309 5544 5321 5584
rect 5358 5544 5370 5604
rect 5394 5544 5406 5602
rect 5460 5544 5472 5584
rect 5488 5544 5500 5584
rect 5510 5544 5522 5564
rect 5559 5544 5571 5584
rect 5589 5544 5601 5584
rect 5659 5544 5671 5584
rect 5689 5544 5701 5584
rect 5720 5544 5732 5584
rect 5748 5544 5760 5584
rect 5776 5544 5788 5584
rect 5851 5544 5863 5584
rect 5871 5544 5883 5584
rect 5891 5544 5903 5572
rect 5911 5544 5923 5584
rect 5937 5544 5949 5564
rect 5957 5544 5969 5564
rect 6000 5544 6012 5584
rect 6028 5544 6040 5584
rect 6056 5544 6068 5584
rect 6118 5544 6130 5604
rect 6154 5544 6166 5602
rect 6231 5544 6243 5564
rect 6251 5544 6263 5564
rect 6280 5544 6292 5584
rect 6308 5544 6320 5584
rect 6330 5544 6342 5564
rect 6378 5544 6390 5604
rect 6414 5544 6426 5602
rect 6478 5544 6490 5604
rect 6514 5544 6526 5602
rect 6578 5544 6590 5604
rect 6614 5544 6626 5602
rect 17 5476 29 5516
rect 39 5496 51 5516
rect 69 5496 81 5516
rect 97 5496 109 5516
rect 123 5496 135 5516
rect 145 5496 157 5516
rect 175 5496 187 5516
rect 207 5496 219 5516
rect 227 5476 239 5516
rect 259 5476 271 5516
rect 289 5476 301 5516
rect 358 5496 370 5516
rect 380 5476 392 5516
rect 408 5476 420 5516
rect 459 5476 471 5516
rect 489 5476 501 5516
rect 541 5476 553 5516
rect 561 5476 573 5516
rect 591 5476 603 5516
rect 617 5496 629 5516
rect 637 5496 649 5516
rect 657 5496 669 5516
rect 697 5496 709 5516
rect 717 5496 729 5516
rect 737 5496 749 5516
rect 779 5476 791 5516
rect 809 5476 821 5516
rect 859 5476 871 5516
rect 889 5476 901 5516
rect 937 5496 949 5516
rect 957 5496 969 5516
rect 1000 5476 1012 5516
rect 1028 5476 1040 5516
rect 1050 5496 1062 5516
rect 1132 5476 1144 5516
rect 1160 5476 1172 5516
rect 1188 5476 1200 5516
rect 1217 5476 1229 5516
rect 1239 5496 1251 5516
rect 1269 5496 1281 5516
rect 1297 5496 1309 5516
rect 1323 5496 1335 5516
rect 1345 5496 1357 5516
rect 1375 5496 1387 5516
rect 1407 5496 1419 5516
rect 1427 5476 1439 5516
rect 1494 5458 1506 5516
rect 1530 5456 1542 5516
rect 1594 5458 1606 5516
rect 1630 5456 1642 5516
rect 1671 5496 1683 5516
rect 1691 5496 1703 5516
rect 1731 5476 1743 5516
rect 1751 5476 1763 5516
rect 1771 5488 1783 5516
rect 1791 5476 1803 5516
rect 1841 5476 1853 5516
rect 1861 5476 1873 5516
rect 1891 5476 1903 5516
rect 1939 5476 1951 5516
rect 1969 5476 1981 5516
rect 2011 5476 2023 5516
rect 2031 5476 2043 5516
rect 2051 5488 2063 5516
rect 2071 5476 2083 5516
rect 2099 5476 2111 5516
rect 2129 5476 2141 5516
rect 2191 5496 2203 5516
rect 2211 5496 2223 5516
rect 2251 5476 2263 5516
rect 2271 5476 2283 5516
rect 2291 5488 2303 5516
rect 2311 5476 2323 5516
rect 2337 5496 2349 5516
rect 2357 5496 2369 5516
rect 2377 5496 2389 5516
rect 2431 5496 2443 5516
rect 2451 5496 2463 5516
rect 2498 5496 2510 5516
rect 2520 5476 2532 5516
rect 2548 5476 2560 5516
rect 2577 5476 2589 5516
rect 2597 5488 2609 5516
rect 2617 5476 2629 5516
rect 2637 5476 2649 5516
rect 2679 5476 2691 5516
rect 2709 5476 2721 5516
rect 2794 5458 2806 5516
rect 2830 5456 2842 5516
rect 2879 5476 2891 5516
rect 2909 5476 2921 5516
rect 2951 5496 2963 5516
rect 2971 5496 2983 5516
rect 2991 5496 3003 5516
rect 3017 5476 3029 5516
rect 3037 5488 3049 5516
rect 3057 5476 3069 5516
rect 3077 5476 3089 5516
rect 3139 5476 3151 5516
rect 3169 5476 3181 5516
rect 3197 5476 3209 5516
rect 3217 5488 3229 5516
rect 3237 5476 3249 5516
rect 3257 5476 3269 5516
rect 3321 5476 3333 5516
rect 3341 5476 3353 5516
rect 3371 5476 3383 5516
rect 3397 5496 3409 5516
rect 3417 5496 3429 5516
rect 3437 5496 3449 5516
rect 3477 5496 3489 5516
rect 3497 5496 3509 5516
rect 3517 5496 3529 5516
rect 3537 5476 3549 5516
rect 3577 5476 3589 5516
rect 3597 5488 3609 5516
rect 3617 5476 3629 5516
rect 3637 5476 3649 5516
rect 3691 5496 3703 5516
rect 3711 5496 3723 5516
rect 3731 5496 3743 5516
rect 3757 5476 3769 5516
rect 3777 5486 3789 5516
rect 3797 5476 3809 5516
rect 3817 5476 3829 5504
rect 3837 5476 3849 5516
rect 3891 5496 3903 5516
rect 3911 5496 3923 5516
rect 3931 5496 3943 5516
rect 3957 5476 3969 5516
rect 3977 5488 3989 5516
rect 3997 5476 4009 5516
rect 4017 5476 4029 5516
rect 4094 5458 4106 5516
rect 4130 5456 4142 5516
rect 4179 5476 4191 5516
rect 4209 5476 4221 5516
rect 4237 5496 4249 5516
rect 4257 5496 4269 5516
rect 4311 5476 4323 5516
rect 4331 5476 4343 5516
rect 4351 5488 4363 5516
rect 4371 5476 4383 5516
rect 4419 5476 4431 5516
rect 4449 5476 4461 5516
rect 4479 5476 4491 5516
rect 4509 5476 4521 5516
rect 4571 5476 4583 5516
rect 4591 5476 4603 5516
rect 4611 5488 4623 5516
rect 4631 5476 4643 5516
rect 4671 5476 4683 5516
rect 4691 5476 4703 5516
rect 4711 5488 4723 5516
rect 4731 5476 4743 5516
rect 4781 5476 4793 5516
rect 4801 5476 4813 5516
rect 4831 5476 4843 5516
rect 4871 5476 4883 5516
rect 4891 5476 4903 5516
rect 4911 5488 4923 5516
rect 4931 5476 4943 5516
rect 4979 5476 4991 5516
rect 5009 5476 5021 5516
rect 5061 5476 5073 5516
rect 5081 5476 5093 5516
rect 5111 5476 5123 5516
rect 5139 5476 5151 5516
rect 5169 5476 5181 5516
rect 5217 5476 5229 5516
rect 5237 5488 5249 5516
rect 5257 5476 5269 5516
rect 5277 5476 5289 5516
rect 5341 5476 5353 5516
rect 5361 5476 5373 5516
rect 5391 5476 5403 5516
rect 5417 5476 5429 5516
rect 5437 5488 5449 5516
rect 5457 5476 5469 5516
rect 5477 5476 5489 5516
rect 5519 5476 5531 5516
rect 5549 5476 5561 5516
rect 5598 5456 5610 5516
rect 5634 5458 5646 5516
rect 5721 5476 5733 5516
rect 5741 5476 5753 5516
rect 5771 5476 5783 5516
rect 5832 5476 5844 5516
rect 5860 5476 5872 5516
rect 5888 5476 5900 5516
rect 5919 5476 5931 5516
rect 5949 5476 5961 5516
rect 5998 5456 6010 5516
rect 6034 5458 6046 5516
rect 6100 5476 6112 5516
rect 6128 5476 6140 5516
rect 6150 5496 6162 5516
rect 6211 5476 6223 5516
rect 6231 5476 6243 5516
rect 6251 5488 6263 5516
rect 6271 5476 6283 5516
rect 6297 5476 6309 5516
rect 6317 5488 6329 5516
rect 6337 5476 6349 5516
rect 6357 5476 6369 5516
rect 6411 5476 6423 5516
rect 6431 5476 6443 5516
rect 6451 5488 6463 5516
rect 6471 5476 6483 5516
rect 6534 5458 6546 5516
rect 6570 5456 6582 5516
rect 6618 5496 6630 5516
rect 6640 5476 6652 5516
rect 6668 5476 6680 5516
rect 29 5064 41 5104
rect 49 5064 61 5104
rect 71 5064 83 5084
rect 97 5064 109 5104
rect 119 5064 131 5084
rect 149 5064 161 5084
rect 177 5064 189 5084
rect 203 5064 215 5084
rect 225 5064 237 5084
rect 255 5064 267 5084
rect 287 5064 299 5084
rect 307 5064 319 5104
rect 339 5064 351 5104
rect 369 5064 381 5104
rect 438 5064 450 5084
rect 460 5064 472 5104
rect 488 5064 500 5104
rect 539 5064 551 5104
rect 569 5064 581 5104
rect 601 5064 613 5104
rect 621 5064 633 5084
rect 653 5064 665 5084
rect 683 5064 695 5084
rect 705 5064 717 5084
rect 731 5064 743 5084
rect 759 5064 771 5084
rect 789 5064 801 5084
rect 811 5064 823 5104
rect 839 5064 851 5104
rect 869 5064 881 5104
rect 931 5064 943 5104
rect 951 5064 963 5104
rect 971 5064 983 5092
rect 991 5064 1003 5104
rect 1031 5064 1043 5104
rect 1051 5064 1063 5104
rect 1071 5064 1083 5092
rect 1091 5064 1103 5104
rect 1141 5064 1153 5104
rect 1161 5064 1173 5104
rect 1191 5064 1203 5104
rect 1217 5064 1229 5104
rect 1239 5064 1251 5084
rect 1269 5064 1281 5084
rect 1297 5064 1309 5084
rect 1323 5064 1335 5084
rect 1345 5064 1357 5084
rect 1375 5064 1387 5084
rect 1407 5064 1419 5084
rect 1427 5064 1439 5104
rect 1479 5064 1491 5104
rect 1509 5064 1521 5104
rect 1539 5064 1551 5104
rect 1569 5064 1581 5104
rect 1617 5064 1629 5104
rect 1639 5064 1651 5084
rect 1669 5064 1681 5084
rect 1697 5064 1709 5084
rect 1723 5064 1735 5084
rect 1745 5064 1757 5084
rect 1775 5064 1787 5084
rect 1807 5064 1819 5084
rect 1827 5064 1839 5104
rect 1892 5064 1904 5104
rect 1920 5064 1932 5104
rect 1948 5064 1960 5104
rect 1977 5064 1989 5084
rect 1997 5064 2009 5084
rect 2061 5064 2073 5104
rect 2081 5064 2093 5104
rect 2111 5064 2123 5104
rect 2139 5064 2151 5104
rect 2169 5064 2181 5104
rect 2231 5064 2243 5104
rect 2251 5064 2263 5084
rect 2271 5064 2283 5084
rect 2291 5064 2303 5084
rect 2339 5064 2351 5104
rect 2369 5064 2381 5104
rect 2434 5064 2446 5122
rect 2470 5064 2482 5124
rect 2511 5064 2523 5084
rect 2531 5064 2543 5084
rect 2551 5064 2563 5084
rect 2577 5064 2589 5084
rect 2597 5064 2609 5084
rect 2661 5064 2673 5104
rect 2681 5064 2693 5104
rect 2711 5064 2723 5104
rect 2737 5064 2749 5084
rect 2757 5064 2769 5084
rect 2777 5064 2789 5084
rect 2839 5064 2851 5104
rect 2869 5064 2881 5104
rect 2919 5064 2931 5104
rect 2949 5064 2961 5104
rect 2977 5064 2989 5084
rect 2997 5064 3009 5084
rect 3017 5064 3029 5084
rect 3037 5064 3049 5104
rect 3101 5064 3113 5104
rect 3121 5064 3133 5104
rect 3151 5064 3163 5104
rect 3179 5064 3191 5104
rect 3209 5064 3221 5104
rect 3294 5064 3306 5122
rect 3330 5064 3342 5124
rect 3371 5064 3383 5084
rect 3391 5064 3403 5084
rect 3438 5064 3450 5084
rect 3460 5064 3472 5104
rect 3488 5064 3500 5104
rect 3531 5064 3543 5084
rect 3551 5064 3563 5084
rect 3571 5064 3583 5084
rect 3597 5064 3609 5104
rect 3617 5064 3629 5092
rect 3637 5064 3649 5104
rect 3657 5064 3669 5104
rect 3711 5064 3723 5104
rect 3731 5064 3743 5104
rect 3751 5064 3763 5092
rect 3771 5064 3783 5104
rect 3797 5064 3809 5084
rect 3817 5064 3829 5084
rect 3837 5064 3849 5084
rect 3879 5064 3891 5104
rect 3909 5064 3921 5104
rect 3979 5064 3991 5104
rect 4009 5064 4021 5104
rect 4037 5064 4049 5104
rect 4057 5064 4069 5092
rect 4077 5064 4089 5104
rect 4097 5064 4109 5104
rect 4159 5064 4171 5104
rect 4189 5064 4201 5104
rect 4241 5064 4253 5104
rect 4261 5064 4273 5104
rect 4291 5064 4303 5104
rect 4339 5064 4351 5104
rect 4369 5064 4381 5104
rect 4411 5064 4423 5104
rect 4431 5064 4443 5104
rect 4451 5064 4463 5092
rect 4471 5064 4483 5104
rect 4511 5064 4523 5104
rect 4531 5064 4543 5104
rect 4551 5064 4563 5092
rect 4571 5064 4583 5104
rect 4599 5064 4611 5104
rect 4629 5064 4641 5104
rect 4679 5064 4691 5104
rect 4709 5064 4721 5104
rect 4757 5064 4769 5084
rect 4777 5064 4789 5084
rect 4854 5064 4866 5122
rect 4890 5064 4902 5124
rect 4917 5064 4929 5104
rect 4937 5064 4949 5092
rect 4957 5064 4969 5104
rect 4977 5064 4989 5104
rect 5017 5064 5029 5104
rect 5037 5064 5049 5104
rect 5079 5064 5091 5104
rect 5109 5064 5121 5104
rect 5157 5064 5169 5104
rect 5177 5064 5189 5104
rect 5197 5064 5209 5104
rect 5239 5064 5251 5104
rect 5269 5064 5281 5104
rect 5317 5064 5329 5104
rect 5337 5064 5349 5092
rect 5357 5064 5369 5104
rect 5377 5064 5389 5104
rect 5418 5064 5430 5124
rect 5454 5064 5466 5122
rect 5518 5064 5530 5124
rect 5554 5064 5566 5122
rect 5617 5064 5629 5084
rect 5637 5064 5649 5084
rect 5678 5064 5690 5124
rect 5714 5064 5726 5122
rect 5777 5064 5789 5104
rect 5797 5064 5809 5092
rect 5817 5064 5829 5104
rect 5837 5064 5849 5104
rect 5899 5064 5911 5104
rect 5929 5064 5941 5104
rect 5958 5064 5970 5124
rect 5994 5064 6006 5122
rect 6059 5064 6071 5104
rect 6089 5064 6101 5104
rect 6158 5064 6170 5084
rect 6180 5064 6192 5104
rect 6208 5064 6220 5104
rect 6251 5064 6263 5084
rect 6271 5064 6283 5084
rect 6334 5064 6346 5122
rect 6370 5064 6382 5124
rect 6434 5064 6446 5122
rect 6470 5064 6482 5124
rect 6497 5064 6509 5084
rect 6517 5064 6529 5084
rect 6594 5064 6606 5122
rect 6630 5064 6642 5124
rect 6659 5064 6671 5104
rect 6689 5064 6701 5104
rect 29 4996 41 5036
rect 49 4996 61 5036
rect 71 5016 83 5036
rect 109 4996 121 5036
rect 129 4996 141 5036
rect 151 5016 163 5036
rect 199 4996 211 5036
rect 229 4996 241 5036
rect 257 4996 269 5036
rect 279 5016 291 5036
rect 309 5016 321 5036
rect 337 5016 349 5036
rect 363 5016 375 5036
rect 385 5016 397 5036
rect 415 5016 427 5036
rect 447 5016 459 5036
rect 467 4996 479 5036
rect 518 5016 530 5036
rect 540 4996 552 5036
rect 568 4996 580 5036
rect 619 4996 631 5036
rect 649 4996 661 5036
rect 679 4996 691 5036
rect 709 4996 721 5036
rect 779 4996 791 5036
rect 809 4996 821 5036
rect 837 4996 849 5036
rect 859 5016 871 5036
rect 889 5016 901 5036
rect 917 5016 929 5036
rect 943 5016 955 5036
rect 965 5016 977 5036
rect 995 5016 1007 5036
rect 1027 5016 1039 5036
rect 1047 4996 1059 5036
rect 1089 4996 1101 5036
rect 1109 4996 1121 5036
rect 1131 5016 1143 5036
rect 1178 5016 1190 5036
rect 1200 4996 1212 5036
rect 1228 4996 1240 5036
rect 1279 4996 1291 5036
rect 1309 4996 1321 5036
rect 1349 4996 1361 5036
rect 1369 4996 1381 5036
rect 1391 5016 1403 5036
rect 1419 4996 1431 5036
rect 1449 4996 1461 5036
rect 1519 4996 1531 5036
rect 1549 4996 1561 5036
rect 1591 4996 1603 5036
rect 1611 4996 1623 5036
rect 1631 5008 1643 5036
rect 1651 4996 1663 5036
rect 1699 4996 1711 5036
rect 1729 4996 1741 5036
rect 1771 4996 1783 5036
rect 1791 4996 1803 5036
rect 1811 5008 1823 5036
rect 1831 4996 1843 5036
rect 1859 4996 1871 5036
rect 1889 4996 1901 5036
rect 1951 4996 1963 5036
rect 1971 4996 1983 5036
rect 1991 5008 2003 5036
rect 2011 4996 2023 5036
rect 2051 4996 2063 5036
rect 2071 4996 2083 5036
rect 2091 5008 2103 5036
rect 2111 4996 2123 5036
rect 2161 4996 2173 5036
rect 2181 4996 2193 5036
rect 2211 4996 2223 5036
rect 2237 5016 2249 5036
rect 2257 5016 2269 5036
rect 2311 5016 2323 5036
rect 2331 5016 2343 5036
rect 2351 5016 2363 5036
rect 2391 4996 2403 5036
rect 2411 5016 2423 5036
rect 2431 5016 2443 5036
rect 2451 5016 2463 5036
rect 2499 4996 2511 5036
rect 2529 4996 2541 5036
rect 2571 4996 2583 5036
rect 2591 4996 2603 5036
rect 2611 5008 2623 5036
rect 2631 4996 2643 5036
rect 2671 4996 2683 5036
rect 2691 4996 2703 5036
rect 2711 5008 2723 5036
rect 2731 4996 2743 5036
rect 2771 5016 2783 5036
rect 2791 5016 2803 5036
rect 2817 4996 2829 5036
rect 2837 5008 2849 5036
rect 2857 4996 2869 5036
rect 2877 4996 2889 5036
rect 2931 4996 2943 5036
rect 2951 4996 2963 5036
rect 2971 5008 2983 5036
rect 2991 4996 3003 5036
rect 3031 4996 3043 5036
rect 3051 4996 3063 5036
rect 3071 5008 3083 5036
rect 3091 4996 3103 5036
rect 3131 5016 3143 5036
rect 3151 5016 3163 5036
rect 3171 5016 3183 5036
rect 3211 4996 3223 5036
rect 3231 4996 3243 5036
rect 3279 4996 3291 5036
rect 3309 4996 3321 5036
rect 3351 4996 3363 5036
rect 3371 4996 3383 5036
rect 3391 5008 3403 5036
rect 3411 4996 3423 5036
rect 3441 4996 3453 5036
rect 3461 5016 3473 5036
rect 3493 5016 3505 5036
rect 3523 5016 3535 5036
rect 3545 5016 3557 5036
rect 3571 5016 3583 5036
rect 3599 5016 3611 5036
rect 3629 5016 3641 5036
rect 3651 4996 3663 5036
rect 3677 4996 3689 5036
rect 3697 5008 3709 5036
rect 3717 4996 3729 5036
rect 3737 4996 3749 5036
rect 3798 5016 3810 5036
rect 3820 4996 3832 5036
rect 3848 4996 3860 5036
rect 3914 4978 3926 5036
rect 3950 4976 3962 5036
rect 3998 5016 4010 5036
rect 4020 4996 4032 5036
rect 4048 4996 4060 5036
rect 4091 4996 4103 5036
rect 4111 4996 4123 5036
rect 4161 4996 4173 5036
rect 4181 4996 4193 5036
rect 4211 4996 4223 5036
rect 4259 4996 4271 5036
rect 4289 4996 4301 5036
rect 4317 4996 4329 5036
rect 4347 4996 4359 5036
rect 4367 4996 4379 5036
rect 4431 4996 4443 5036
rect 4451 4996 4463 5036
rect 4471 5008 4483 5036
rect 4491 4996 4503 5036
rect 4518 4976 4530 5036
rect 4554 4978 4566 5036
rect 4617 4996 4629 5036
rect 4637 5008 4649 5036
rect 4657 4996 4669 5036
rect 4677 4996 4689 5036
rect 4739 4996 4751 5036
rect 4769 4996 4781 5036
rect 4821 4996 4833 5036
rect 4841 4996 4853 5036
rect 4871 4996 4883 5036
rect 4919 4996 4931 5036
rect 4949 4996 4961 5036
rect 4979 4996 4991 5036
rect 5009 4996 5021 5036
rect 5057 4996 5069 5036
rect 5087 4996 5099 5036
rect 5107 4996 5119 5036
rect 5179 4996 5191 5036
rect 5209 4996 5221 5036
rect 5261 4996 5273 5036
rect 5281 4996 5293 5036
rect 5311 4996 5323 5036
rect 5337 4996 5349 5036
rect 5367 4996 5379 5036
rect 5387 4996 5399 5036
rect 5472 4996 5484 5036
rect 5500 4996 5512 5036
rect 5528 4996 5540 5036
rect 5579 4996 5591 5036
rect 5609 4996 5621 5036
rect 5638 4976 5650 5036
rect 5674 4978 5686 5036
rect 5758 5016 5770 5036
rect 5780 4996 5792 5036
rect 5808 4996 5820 5036
rect 5874 4978 5886 5036
rect 5910 4976 5922 5036
rect 5959 4996 5971 5036
rect 5989 4996 6001 5036
rect 6020 4996 6032 5036
rect 6048 4996 6060 5036
rect 6076 4996 6088 5036
rect 6174 4978 6186 5036
rect 6210 4976 6222 5036
rect 6237 4996 6249 5036
rect 6257 5008 6269 5036
rect 6277 4996 6289 5036
rect 6297 4996 6309 5036
rect 6374 4978 6386 5036
rect 6410 4976 6422 5036
rect 6474 4978 6486 5036
rect 6510 4976 6522 5036
rect 6539 4996 6551 5036
rect 6569 4996 6581 5036
rect 6631 5016 6643 5036
rect 6651 5016 6663 5036
rect 17 4584 29 4624
rect 37 4584 49 4624
rect 57 4584 69 4624
rect 77 4584 89 4624
rect 97 4584 109 4624
rect 117 4584 129 4624
rect 137 4584 149 4624
rect 157 4584 169 4624
rect 177 4584 189 4624
rect 231 4584 243 4604
rect 251 4584 263 4604
rect 271 4584 283 4604
rect 311 4584 323 4604
rect 331 4584 343 4604
rect 378 4584 390 4604
rect 400 4584 412 4624
rect 428 4584 440 4624
rect 471 4584 483 4604
rect 491 4584 503 4604
rect 531 4584 543 4604
rect 551 4584 563 4604
rect 571 4584 583 4604
rect 621 4584 633 4624
rect 641 4584 653 4624
rect 671 4584 683 4624
rect 697 4584 709 4604
rect 717 4584 729 4604
rect 737 4584 749 4604
rect 789 4584 801 4624
rect 809 4584 821 4624
rect 831 4584 843 4604
rect 879 4584 891 4624
rect 909 4584 921 4624
rect 937 4584 949 4624
rect 959 4584 971 4604
rect 989 4584 1001 4604
rect 1017 4584 1029 4604
rect 1043 4584 1055 4604
rect 1065 4584 1077 4604
rect 1095 4584 1107 4604
rect 1127 4584 1139 4604
rect 1147 4584 1159 4624
rect 1191 4584 1203 4624
rect 1211 4584 1223 4624
rect 1231 4584 1243 4612
rect 1251 4584 1263 4624
rect 1299 4584 1311 4624
rect 1329 4584 1341 4624
rect 1359 4584 1371 4624
rect 1389 4584 1401 4624
rect 1451 4584 1463 4624
rect 1471 4584 1483 4624
rect 1491 4584 1503 4612
rect 1511 4584 1523 4624
rect 1537 4584 1549 4604
rect 1557 4584 1569 4604
rect 1577 4584 1589 4604
rect 1617 4584 1629 4604
rect 1637 4584 1649 4604
rect 1657 4584 1669 4604
rect 1697 4584 1709 4604
rect 1717 4584 1729 4604
rect 1757 4584 1769 4604
rect 1777 4584 1789 4604
rect 1797 4584 1809 4604
rect 1837 4584 1849 4624
rect 1857 4584 1869 4612
rect 1877 4584 1889 4624
rect 1897 4584 1909 4624
rect 1937 4584 1949 4624
rect 1959 4584 1971 4604
rect 1989 4584 2001 4604
rect 2017 4584 2029 4604
rect 2043 4584 2055 4604
rect 2065 4584 2077 4604
rect 2095 4584 2107 4604
rect 2127 4584 2139 4604
rect 2147 4584 2159 4624
rect 2199 4584 2211 4624
rect 2229 4584 2241 4624
rect 2271 4584 2283 4624
rect 2291 4584 2303 4604
rect 2311 4584 2323 4604
rect 2331 4584 2343 4604
rect 2359 4584 2371 4624
rect 2389 4584 2401 4624
rect 2437 4584 2449 4604
rect 2457 4584 2469 4604
rect 2477 4584 2489 4604
rect 2520 4584 2532 4624
rect 2548 4584 2560 4624
rect 2570 4584 2582 4604
rect 2631 4584 2643 4604
rect 2651 4584 2663 4604
rect 2677 4584 2689 4624
rect 2699 4584 2711 4604
rect 2729 4584 2741 4604
rect 2757 4584 2769 4604
rect 2783 4584 2795 4604
rect 2805 4584 2817 4604
rect 2835 4584 2847 4604
rect 2867 4584 2879 4604
rect 2887 4584 2899 4624
rect 2917 4584 2929 4624
rect 2937 4584 2949 4612
rect 2957 4584 2969 4624
rect 2977 4584 2989 4624
rect 3017 4584 3029 4624
rect 3039 4584 3051 4604
rect 3069 4584 3081 4604
rect 3097 4584 3109 4604
rect 3123 4584 3135 4604
rect 3145 4584 3157 4604
rect 3175 4584 3187 4604
rect 3207 4584 3219 4604
rect 3227 4584 3239 4624
rect 3257 4584 3269 4624
rect 3279 4584 3291 4604
rect 3309 4584 3321 4604
rect 3337 4584 3349 4604
rect 3363 4584 3375 4604
rect 3385 4584 3397 4604
rect 3415 4584 3427 4604
rect 3447 4584 3459 4604
rect 3467 4584 3479 4624
rect 3511 4584 3523 4624
rect 3531 4584 3543 4624
rect 3551 4584 3563 4612
rect 3571 4584 3583 4624
rect 3611 4584 3623 4624
rect 3631 4584 3643 4624
rect 3679 4584 3691 4624
rect 3709 4584 3721 4624
rect 3751 4584 3763 4624
rect 3771 4584 3783 4624
rect 3791 4584 3803 4612
rect 3811 4584 3823 4624
rect 3841 4584 3853 4624
rect 3861 4584 3873 4604
rect 3893 4584 3905 4604
rect 3923 4584 3935 4604
rect 3945 4584 3957 4604
rect 3971 4584 3983 4604
rect 3999 4584 4011 4604
rect 4029 4584 4041 4604
rect 4051 4584 4063 4624
rect 4091 4584 4103 4624
rect 4111 4584 4123 4624
rect 4159 4584 4171 4624
rect 4189 4584 4201 4624
rect 4217 4584 4229 4624
rect 4239 4584 4251 4604
rect 4269 4584 4281 4604
rect 4297 4584 4309 4604
rect 4323 4584 4335 4604
rect 4345 4584 4357 4604
rect 4375 4584 4387 4604
rect 4407 4584 4419 4604
rect 4427 4584 4439 4624
rect 4494 4584 4506 4642
rect 4530 4584 4542 4644
rect 4557 4584 4569 4604
rect 4577 4584 4589 4604
rect 4617 4584 4629 4624
rect 4637 4584 4649 4624
rect 4691 4584 4703 4604
rect 4711 4584 4723 4604
rect 4737 4584 4749 4624
rect 4757 4584 4769 4612
rect 4777 4584 4789 4624
rect 4797 4584 4809 4624
rect 4837 4584 4849 4604
rect 4857 4584 4869 4604
rect 4877 4584 4889 4604
rect 4919 4584 4931 4624
rect 4949 4584 4961 4624
rect 4999 4584 5011 4624
rect 5029 4584 5041 4624
rect 5099 4584 5111 4624
rect 5129 4584 5141 4624
rect 5157 4584 5169 4624
rect 5177 4584 5189 4612
rect 5197 4584 5209 4624
rect 5217 4584 5229 4624
rect 5271 4584 5283 4624
rect 5291 4596 5303 4624
rect 5311 4584 5323 4624
rect 5331 4584 5343 4614
rect 5351 4584 5363 4624
rect 5379 4584 5391 4624
rect 5409 4584 5421 4624
rect 5479 4584 5491 4624
rect 5509 4584 5521 4624
rect 5538 4584 5550 4644
rect 5574 4584 5586 4642
rect 5659 4584 5671 4624
rect 5689 4584 5701 4624
rect 5718 4584 5730 4644
rect 5754 4584 5766 4642
rect 5831 4584 5843 4604
rect 5851 4584 5863 4604
rect 5878 4584 5890 4644
rect 5914 4584 5926 4642
rect 6001 4584 6013 4624
rect 6021 4584 6033 4624
rect 6051 4584 6063 4624
rect 6077 4584 6089 4624
rect 6097 4584 6109 4612
rect 6117 4584 6129 4624
rect 6137 4584 6149 4624
rect 6199 4584 6211 4624
rect 6229 4584 6241 4624
rect 6260 4584 6272 4624
rect 6288 4584 6300 4624
rect 6310 4584 6322 4604
rect 6358 4584 6370 4644
rect 6394 4584 6406 4642
rect 6481 4584 6493 4624
rect 6501 4584 6513 4624
rect 6531 4584 6543 4624
rect 6594 4584 6606 4642
rect 6630 4584 6642 4644
rect 31 4536 43 4556
rect 51 4536 63 4556
rect 91 4536 103 4556
rect 111 4536 123 4556
rect 131 4536 143 4556
rect 171 4536 183 4556
rect 191 4536 203 4556
rect 217 4516 229 4556
rect 237 4528 249 4556
rect 257 4516 269 4556
rect 277 4516 289 4556
rect 331 4536 343 4556
rect 351 4536 363 4556
rect 371 4536 383 4556
rect 397 4516 409 4556
rect 417 4528 429 4556
rect 437 4516 449 4556
rect 457 4516 469 4556
rect 497 4536 509 4556
rect 517 4536 529 4556
rect 537 4536 549 4556
rect 557 4516 569 4556
rect 600 4516 612 4556
rect 628 4516 640 4556
rect 650 4536 662 4556
rect 711 4536 723 4556
rect 731 4536 743 4556
rect 757 4536 769 4556
rect 777 4536 789 4556
rect 797 4536 809 4556
rect 837 4536 849 4556
rect 857 4536 869 4556
rect 897 4536 909 4556
rect 917 4536 929 4556
rect 937 4536 949 4556
rect 977 4536 989 4556
rect 997 4536 1009 4556
rect 1037 4516 1049 4556
rect 1057 4516 1069 4556
rect 1077 4516 1089 4556
rect 1097 4516 1109 4556
rect 1117 4516 1129 4556
rect 1137 4516 1149 4556
rect 1157 4516 1169 4556
rect 1177 4516 1189 4556
rect 1197 4516 1209 4556
rect 1237 4536 1249 4556
rect 1259 4516 1271 4556
rect 1279 4516 1291 4556
rect 1331 4536 1343 4556
rect 1351 4536 1363 4556
rect 1391 4536 1403 4556
rect 1411 4536 1423 4556
rect 1431 4536 1443 4556
rect 1479 4516 1491 4556
rect 1509 4516 1521 4556
rect 1539 4516 1551 4556
rect 1569 4516 1581 4556
rect 1631 4516 1643 4556
rect 1651 4516 1663 4556
rect 1671 4516 1683 4556
rect 1691 4516 1703 4556
rect 1711 4516 1723 4556
rect 1741 4516 1753 4556
rect 1761 4536 1773 4556
rect 1793 4536 1805 4556
rect 1823 4536 1835 4556
rect 1845 4536 1857 4556
rect 1871 4536 1883 4556
rect 1899 4536 1911 4556
rect 1929 4536 1941 4556
rect 1951 4516 1963 4556
rect 1979 4516 1991 4556
rect 2009 4516 2021 4556
rect 2057 4516 2069 4556
rect 2079 4536 2091 4556
rect 2109 4536 2121 4556
rect 2137 4536 2149 4556
rect 2163 4536 2175 4556
rect 2185 4536 2197 4556
rect 2215 4536 2227 4556
rect 2247 4536 2259 4556
rect 2267 4516 2279 4556
rect 2297 4536 2309 4556
rect 2317 4536 2329 4556
rect 2357 4536 2369 4556
rect 2377 4536 2389 4556
rect 2397 4536 2409 4556
rect 2437 4536 2449 4556
rect 2457 4536 2469 4556
rect 2477 4536 2489 4556
rect 2517 4536 2529 4556
rect 2537 4536 2549 4556
rect 2577 4516 2589 4556
rect 2599 4536 2611 4556
rect 2629 4536 2641 4556
rect 2657 4536 2669 4556
rect 2683 4536 2695 4556
rect 2705 4536 2717 4556
rect 2735 4536 2747 4556
rect 2767 4536 2779 4556
rect 2787 4516 2799 4556
rect 2817 4516 2829 4556
rect 2837 4528 2849 4556
rect 2857 4516 2869 4556
rect 2877 4516 2889 4556
rect 2919 4516 2931 4556
rect 2949 4516 2961 4556
rect 3011 4536 3023 4556
rect 3031 4536 3043 4556
rect 3057 4516 3069 4556
rect 3077 4528 3089 4556
rect 3097 4516 3109 4556
rect 3117 4516 3129 4556
rect 3157 4516 3169 4556
rect 3179 4536 3191 4556
rect 3209 4536 3221 4556
rect 3237 4536 3249 4556
rect 3263 4536 3275 4556
rect 3285 4536 3297 4556
rect 3315 4536 3327 4556
rect 3347 4536 3359 4556
rect 3367 4516 3379 4556
rect 3397 4516 3409 4556
rect 3417 4528 3429 4556
rect 3437 4516 3449 4556
rect 3457 4516 3469 4556
rect 3511 4516 3523 4556
rect 3531 4516 3543 4556
rect 3551 4528 3563 4556
rect 3571 4516 3583 4556
rect 3601 4516 3613 4556
rect 3621 4536 3633 4556
rect 3653 4536 3665 4556
rect 3683 4536 3695 4556
rect 3705 4536 3717 4556
rect 3731 4536 3743 4556
rect 3759 4536 3771 4556
rect 3789 4536 3801 4556
rect 3811 4516 3823 4556
rect 3837 4516 3849 4556
rect 3857 4528 3869 4556
rect 3877 4516 3889 4556
rect 3897 4516 3909 4556
rect 3941 4516 3953 4556
rect 3961 4536 3973 4556
rect 3993 4536 4005 4556
rect 4023 4536 4035 4556
rect 4045 4536 4057 4556
rect 4071 4536 4083 4556
rect 4099 4536 4111 4556
rect 4129 4536 4141 4556
rect 4151 4516 4163 4556
rect 4214 4498 4226 4556
rect 4250 4496 4262 4556
rect 4277 4516 4289 4556
rect 4297 4528 4309 4556
rect 4317 4516 4329 4556
rect 4337 4516 4349 4556
rect 4391 4536 4403 4556
rect 4411 4536 4423 4556
rect 4431 4536 4443 4556
rect 4478 4536 4490 4556
rect 4500 4516 4512 4556
rect 4528 4516 4540 4556
rect 4558 4496 4570 4556
rect 4594 4498 4606 4556
rect 4671 4536 4683 4556
rect 4691 4536 4703 4556
rect 4717 4516 4729 4556
rect 4737 4528 4749 4556
rect 4757 4516 4769 4556
rect 4777 4516 4789 4556
rect 4831 4516 4843 4556
rect 4851 4536 4863 4556
rect 4871 4536 4883 4556
rect 4891 4536 4903 4556
rect 4939 4516 4951 4556
rect 4969 4516 4981 4556
rect 5034 4498 5046 4556
rect 5070 4496 5082 4556
rect 5097 4516 5109 4556
rect 5117 4528 5129 4556
rect 5137 4516 5149 4556
rect 5157 4516 5169 4556
rect 5211 4516 5223 4556
rect 5231 4536 5243 4556
rect 5251 4536 5263 4556
rect 5271 4536 5283 4556
rect 5297 4516 5309 4556
rect 5317 4528 5329 4556
rect 5337 4516 5349 4556
rect 5357 4516 5369 4556
rect 5397 4536 5409 4556
rect 5417 4536 5429 4556
rect 5494 4498 5506 4556
rect 5530 4496 5542 4556
rect 5559 4516 5571 4556
rect 5589 4516 5601 4556
rect 5637 4516 5649 4556
rect 5657 4528 5669 4556
rect 5677 4516 5689 4556
rect 5697 4516 5709 4556
rect 5759 4516 5771 4556
rect 5789 4516 5801 4556
rect 5854 4498 5866 4556
rect 5890 4496 5902 4556
rect 5931 4516 5943 4556
rect 5951 4516 5963 4556
rect 5971 4528 5983 4556
rect 5991 4516 6003 4556
rect 6017 4536 6029 4556
rect 6037 4536 6049 4556
rect 6091 4536 6103 4556
rect 6111 4536 6123 4556
rect 6138 4496 6150 4556
rect 6174 4498 6186 4556
rect 6251 4516 6263 4556
rect 6271 4516 6283 4556
rect 6291 4528 6303 4556
rect 6311 4516 6323 4556
rect 6338 4496 6350 4556
rect 6374 4498 6386 4556
rect 6438 4496 6450 4556
rect 6474 4498 6486 4556
rect 6537 4516 6549 4556
rect 6557 4528 6569 4556
rect 6577 4516 6589 4556
rect 6597 4516 6609 4556
rect 6637 4536 6649 4556
rect 6657 4536 6669 4556
rect 29 4104 41 4144
rect 49 4104 61 4144
rect 71 4104 83 4124
rect 111 4104 123 4144
rect 131 4104 143 4144
rect 151 4104 163 4132
rect 171 4104 183 4144
rect 197 4104 209 4144
rect 217 4104 229 4132
rect 237 4104 249 4144
rect 257 4104 269 4144
rect 301 4104 313 4144
rect 321 4104 333 4124
rect 353 4104 365 4124
rect 383 4104 395 4124
rect 405 4104 417 4124
rect 431 4104 443 4124
rect 459 4104 471 4124
rect 489 4104 501 4124
rect 511 4104 523 4144
rect 539 4104 551 4144
rect 569 4104 581 4144
rect 652 4104 664 4144
rect 680 4104 692 4144
rect 708 4104 720 4144
rect 751 4104 763 4124
rect 771 4104 783 4124
rect 797 4104 809 4144
rect 819 4104 831 4124
rect 849 4104 861 4124
rect 877 4104 889 4124
rect 903 4104 915 4124
rect 925 4104 937 4124
rect 955 4104 967 4124
rect 987 4104 999 4124
rect 1007 4104 1019 4144
rect 1039 4104 1051 4144
rect 1069 4104 1081 4144
rect 1117 4104 1129 4144
rect 1139 4104 1151 4124
rect 1169 4104 1181 4124
rect 1197 4104 1209 4124
rect 1223 4104 1235 4124
rect 1245 4104 1257 4124
rect 1275 4104 1287 4124
rect 1307 4104 1319 4124
rect 1327 4104 1339 4144
rect 1359 4104 1371 4144
rect 1389 4104 1401 4144
rect 1437 4104 1449 4124
rect 1457 4104 1469 4124
rect 1511 4104 1523 4144
rect 1531 4104 1543 4144
rect 1551 4104 1563 4132
rect 1571 4104 1583 4144
rect 1618 4104 1630 4124
rect 1640 4104 1652 4144
rect 1668 4104 1680 4144
rect 1719 4104 1731 4144
rect 1749 4104 1761 4144
rect 1779 4104 1791 4144
rect 1809 4104 1821 4144
rect 1857 4104 1869 4144
rect 1879 4104 1891 4124
rect 1909 4104 1921 4124
rect 1937 4104 1949 4124
rect 1963 4104 1975 4124
rect 1985 4104 1997 4124
rect 2015 4104 2027 4124
rect 2047 4104 2059 4124
rect 2067 4104 2079 4144
rect 2099 4104 2111 4144
rect 2129 4104 2141 4144
rect 2191 4104 2203 4144
rect 2211 4104 2223 4144
rect 2231 4104 2243 4132
rect 2251 4104 2263 4144
rect 2281 4104 2293 4144
rect 2301 4104 2313 4124
rect 2333 4104 2345 4124
rect 2363 4104 2375 4124
rect 2385 4104 2397 4124
rect 2411 4104 2423 4124
rect 2439 4104 2451 4124
rect 2469 4104 2481 4124
rect 2491 4104 2503 4144
rect 2531 4104 2543 4124
rect 2551 4104 2563 4124
rect 2571 4104 2583 4124
rect 2597 4104 2609 4124
rect 2617 4104 2629 4124
rect 2657 4104 2669 4144
rect 2677 4104 2689 4132
rect 2697 4104 2709 4144
rect 2717 4104 2729 4144
rect 2759 4104 2771 4144
rect 2789 4104 2801 4144
rect 2851 4104 2863 4144
rect 2871 4104 2883 4144
rect 2891 4104 2903 4132
rect 2911 4104 2923 4144
rect 2937 4104 2949 4124
rect 2957 4104 2969 4124
rect 2997 4104 3009 4124
rect 3017 4104 3029 4124
rect 3037 4104 3049 4124
rect 3091 4104 3103 4124
rect 3111 4104 3123 4124
rect 3137 4104 3149 4144
rect 3159 4104 3171 4124
rect 3189 4104 3201 4124
rect 3217 4104 3229 4124
rect 3243 4104 3255 4124
rect 3265 4104 3277 4124
rect 3295 4104 3307 4124
rect 3327 4104 3339 4124
rect 3347 4104 3359 4144
rect 3377 4104 3389 4144
rect 3397 4104 3409 4134
rect 3417 4104 3429 4144
rect 3437 4116 3449 4144
rect 3457 4104 3469 4144
rect 3499 4104 3511 4144
rect 3529 4104 3541 4144
rect 3577 4104 3589 4144
rect 3597 4104 3609 4144
rect 3617 4104 3629 4144
rect 3637 4104 3649 4144
rect 3657 4104 3669 4144
rect 3677 4104 3689 4144
rect 3697 4104 3709 4144
rect 3717 4104 3729 4144
rect 3737 4104 3749 4144
rect 3779 4104 3791 4144
rect 3809 4104 3821 4144
rect 3859 4104 3871 4144
rect 3889 4104 3901 4144
rect 3959 4104 3971 4144
rect 3989 4104 4001 4144
rect 4017 4104 4029 4124
rect 4037 4104 4049 4124
rect 4091 4104 4103 4144
rect 4111 4104 4123 4144
rect 4131 4104 4143 4132
rect 4151 4104 4163 4144
rect 4177 4104 4189 4144
rect 4197 4104 4209 4132
rect 4217 4104 4229 4144
rect 4237 4104 4249 4144
rect 4281 4104 4293 4144
rect 4301 4104 4313 4124
rect 4333 4104 4345 4124
rect 4363 4104 4375 4124
rect 4385 4104 4397 4124
rect 4411 4104 4423 4124
rect 4439 4104 4451 4124
rect 4469 4104 4481 4124
rect 4491 4104 4503 4144
rect 4531 4104 4543 4144
rect 4551 4104 4563 4144
rect 4571 4104 4583 4132
rect 4591 4104 4603 4144
rect 4621 4104 4633 4144
rect 4641 4104 4653 4124
rect 4673 4104 4685 4124
rect 4703 4104 4715 4124
rect 4725 4104 4737 4124
rect 4751 4104 4763 4124
rect 4779 4104 4791 4124
rect 4809 4104 4821 4124
rect 4831 4104 4843 4144
rect 4871 4104 4883 4144
rect 4891 4104 4903 4144
rect 4938 4104 4950 4124
rect 4960 4104 4972 4144
rect 4988 4104 5000 4144
rect 5018 4104 5030 4164
rect 5054 4104 5066 4162
rect 5131 4104 5143 4124
rect 5151 4104 5163 4124
rect 5177 4104 5189 4144
rect 5197 4104 5209 4132
rect 5217 4104 5229 4144
rect 5237 4104 5249 4144
rect 5281 4104 5293 4144
rect 5301 4104 5313 4124
rect 5333 4104 5345 4124
rect 5363 4104 5375 4124
rect 5385 4104 5397 4124
rect 5411 4104 5423 4124
rect 5439 4104 5451 4124
rect 5469 4104 5481 4124
rect 5491 4104 5503 4144
rect 5519 4104 5531 4144
rect 5549 4104 5561 4144
rect 5597 4104 5609 4124
rect 5617 4104 5629 4124
rect 5657 4104 5669 4144
rect 5677 4104 5689 4132
rect 5697 4104 5709 4144
rect 5717 4104 5729 4144
rect 5781 4104 5793 4144
rect 5801 4104 5813 4144
rect 5831 4104 5843 4144
rect 5858 4104 5870 4164
rect 5894 4104 5906 4162
rect 5971 4104 5983 4144
rect 5991 4104 6003 4144
rect 6017 4104 6029 4144
rect 6037 4104 6049 4132
rect 6057 4104 6069 4144
rect 6077 4104 6089 4144
rect 6117 4104 6129 4124
rect 6139 4104 6151 4144
rect 6159 4104 6171 4144
rect 6199 4104 6211 4144
rect 6229 4104 6241 4144
rect 6301 4104 6313 4144
rect 6321 4104 6333 4144
rect 6351 4104 6363 4144
rect 6379 4104 6391 4144
rect 6409 4104 6421 4144
rect 6457 4104 6469 4124
rect 6477 4104 6489 4124
rect 6538 4104 6550 4124
rect 6560 4104 6572 4144
rect 6588 4104 6600 4144
rect 6618 4104 6630 4164
rect 6654 4104 6666 4162
rect 29 4036 41 4076
rect 49 4036 61 4076
rect 71 4056 83 4076
rect 97 4036 109 4076
rect 119 4056 131 4076
rect 149 4056 161 4076
rect 177 4056 189 4076
rect 203 4056 215 4076
rect 225 4056 237 4076
rect 255 4056 267 4076
rect 287 4056 299 4076
rect 307 4036 319 4076
rect 339 4036 351 4076
rect 369 4036 381 4076
rect 438 4056 450 4076
rect 460 4036 472 4076
rect 488 4036 500 4076
rect 539 4036 551 4076
rect 569 4036 581 4076
rect 619 4036 631 4076
rect 649 4036 661 4076
rect 689 4036 701 4076
rect 709 4036 721 4076
rect 731 4056 743 4076
rect 757 4036 769 4076
rect 779 4056 791 4076
rect 809 4056 821 4076
rect 837 4056 849 4076
rect 863 4056 875 4076
rect 885 4056 897 4076
rect 915 4056 927 4076
rect 947 4056 959 4076
rect 967 4036 979 4076
rect 1019 4036 1031 4076
rect 1049 4036 1061 4076
rect 1079 4036 1091 4076
rect 1109 4036 1121 4076
rect 1159 4036 1171 4076
rect 1189 4036 1201 4076
rect 1258 4056 1270 4076
rect 1280 4036 1292 4076
rect 1308 4036 1320 4076
rect 1337 4036 1349 4076
rect 1359 4056 1371 4076
rect 1389 4056 1401 4076
rect 1417 4056 1429 4076
rect 1443 4056 1455 4076
rect 1465 4056 1477 4076
rect 1495 4056 1507 4076
rect 1527 4056 1539 4076
rect 1547 4036 1559 4076
rect 1599 4036 1611 4076
rect 1629 4036 1641 4076
rect 1657 4056 1669 4076
rect 1679 4036 1691 4076
rect 1699 4036 1711 4076
rect 1739 4036 1751 4076
rect 1769 4036 1781 4076
rect 1817 4036 1829 4076
rect 1839 4056 1851 4076
rect 1869 4056 1881 4076
rect 1897 4056 1909 4076
rect 1923 4056 1935 4076
rect 1945 4056 1957 4076
rect 1975 4056 1987 4076
rect 2007 4056 2019 4076
rect 2027 4036 2039 4076
rect 2059 4036 2071 4076
rect 2089 4036 2101 4076
rect 2151 4036 2163 4076
rect 2171 4036 2183 4076
rect 2191 4048 2203 4076
rect 2211 4036 2223 4076
rect 2259 4036 2271 4076
rect 2289 4036 2301 4076
rect 2319 4036 2331 4076
rect 2349 4036 2361 4076
rect 2411 4056 2423 4076
rect 2431 4056 2443 4076
rect 2471 4036 2483 4076
rect 2491 4036 2503 4076
rect 2511 4048 2523 4076
rect 2531 4036 2543 4076
rect 2557 4056 2569 4076
rect 2577 4056 2589 4076
rect 2597 4056 2609 4076
rect 2651 4056 2663 4076
rect 2671 4056 2683 4076
rect 2691 4056 2703 4076
rect 2717 4056 2729 4076
rect 2737 4056 2749 4076
rect 2791 4056 2803 4076
rect 2811 4056 2823 4076
rect 2859 4036 2871 4076
rect 2889 4036 2901 4076
rect 2917 4056 2929 4076
rect 2937 4056 2949 4076
rect 2957 4056 2969 4076
rect 2997 4036 3009 4076
rect 3017 4048 3029 4076
rect 3037 4036 3049 4076
rect 3057 4036 3069 4076
rect 3097 4056 3109 4076
rect 3117 4056 3129 4076
rect 3157 4056 3169 4076
rect 3177 4056 3189 4076
rect 3197 4056 3209 4076
rect 3259 4036 3271 4076
rect 3289 4036 3301 4076
rect 3339 4036 3351 4076
rect 3369 4036 3381 4076
rect 3401 4036 3413 4076
rect 3421 4056 3433 4076
rect 3453 4056 3465 4076
rect 3483 4056 3495 4076
rect 3505 4056 3517 4076
rect 3531 4056 3543 4076
rect 3559 4056 3571 4076
rect 3589 4056 3601 4076
rect 3611 4036 3623 4076
rect 3651 4056 3663 4076
rect 3671 4056 3683 4076
rect 3701 4036 3713 4076
rect 3721 4056 3733 4076
rect 3753 4056 3765 4076
rect 3783 4056 3795 4076
rect 3805 4056 3817 4076
rect 3831 4056 3843 4076
rect 3859 4056 3871 4076
rect 3889 4056 3901 4076
rect 3911 4036 3923 4076
rect 3974 4018 3986 4076
rect 4010 4016 4022 4076
rect 4039 4036 4051 4076
rect 4069 4036 4081 4076
rect 4131 4036 4143 4076
rect 4151 4036 4163 4076
rect 4171 4048 4183 4076
rect 4191 4036 4203 4076
rect 4217 4056 4229 4076
rect 4237 4056 4249 4076
rect 4257 4056 4269 4076
rect 4311 4056 4323 4076
rect 4331 4056 4343 4076
rect 4379 4036 4391 4076
rect 4409 4036 4421 4076
rect 4451 4036 4463 4076
rect 4471 4036 4483 4076
rect 4491 4048 4503 4076
rect 4511 4036 4523 4076
rect 4541 4036 4553 4076
rect 4561 4056 4573 4076
rect 4593 4056 4605 4076
rect 4623 4056 4635 4076
rect 4645 4056 4657 4076
rect 4671 4056 4683 4076
rect 4699 4056 4711 4076
rect 4729 4056 4741 4076
rect 4751 4036 4763 4076
rect 4799 4036 4811 4076
rect 4829 4036 4841 4076
rect 4871 4036 4883 4076
rect 4891 4036 4903 4076
rect 4911 4048 4923 4076
rect 4931 4036 4943 4076
rect 4961 4036 4973 4076
rect 4981 4056 4993 4076
rect 5013 4056 5025 4076
rect 5043 4056 5055 4076
rect 5065 4056 5077 4076
rect 5091 4056 5103 4076
rect 5119 4056 5131 4076
rect 5149 4056 5161 4076
rect 5171 4036 5183 4076
rect 5219 4036 5231 4076
rect 5249 4036 5261 4076
rect 5291 4036 5303 4076
rect 5311 4036 5323 4076
rect 5331 4048 5343 4076
rect 5351 4036 5363 4076
rect 5399 4036 5411 4076
rect 5429 4036 5441 4076
rect 5457 4036 5469 4076
rect 5477 4048 5489 4076
rect 5497 4036 5509 4076
rect 5517 4036 5529 4076
rect 5571 4056 5583 4076
rect 5591 4056 5603 4076
rect 5621 4036 5633 4076
rect 5641 4056 5653 4076
rect 5673 4056 5685 4076
rect 5703 4056 5715 4076
rect 5725 4056 5737 4076
rect 5751 4056 5763 4076
rect 5779 4056 5791 4076
rect 5809 4056 5821 4076
rect 5831 4036 5843 4076
rect 5857 4056 5869 4076
rect 5877 4056 5889 4076
rect 5954 4018 5966 4076
rect 5990 4016 6002 4076
rect 6017 4036 6029 4076
rect 6039 4056 6051 4076
rect 6069 4056 6081 4076
rect 6097 4056 6109 4076
rect 6123 4056 6135 4076
rect 6145 4056 6157 4076
rect 6175 4056 6187 4076
rect 6207 4056 6219 4076
rect 6227 4036 6239 4076
rect 6257 4036 6269 4076
rect 6279 4056 6291 4076
rect 6309 4056 6321 4076
rect 6337 4056 6349 4076
rect 6363 4056 6375 4076
rect 6385 4056 6397 4076
rect 6415 4056 6427 4076
rect 6447 4056 6459 4076
rect 6467 4036 6479 4076
rect 6497 4036 6509 4076
rect 6519 4056 6531 4076
rect 6549 4056 6561 4076
rect 6577 4056 6589 4076
rect 6603 4056 6615 4076
rect 6625 4056 6637 4076
rect 6655 4056 6667 4076
rect 6687 4056 6699 4076
rect 6707 4036 6719 4076
rect 29 3624 41 3664
rect 49 3624 61 3664
rect 71 3624 83 3644
rect 109 3624 121 3664
rect 129 3624 141 3664
rect 151 3624 163 3644
rect 199 3624 211 3664
rect 229 3624 241 3664
rect 257 3624 269 3664
rect 279 3624 291 3644
rect 309 3624 321 3644
rect 337 3624 349 3644
rect 363 3624 375 3644
rect 385 3624 397 3644
rect 415 3624 427 3644
rect 447 3624 459 3644
rect 467 3624 479 3664
rect 518 3624 530 3644
rect 540 3624 552 3664
rect 568 3624 580 3664
rect 619 3624 631 3664
rect 649 3624 661 3664
rect 679 3624 691 3664
rect 709 3624 721 3664
rect 779 3624 791 3664
rect 809 3624 821 3664
rect 837 3624 849 3664
rect 859 3624 871 3644
rect 889 3624 901 3644
rect 917 3624 929 3644
rect 943 3624 955 3644
rect 965 3624 977 3644
rect 995 3624 1007 3644
rect 1027 3624 1039 3644
rect 1047 3624 1059 3664
rect 1080 3624 1092 3664
rect 1108 3624 1120 3664
rect 1130 3624 1142 3644
rect 1199 3624 1211 3664
rect 1229 3624 1241 3664
rect 1257 3624 1269 3644
rect 1279 3624 1291 3664
rect 1299 3624 1311 3664
rect 1358 3624 1370 3644
rect 1380 3624 1392 3664
rect 1408 3624 1420 3664
rect 1459 3624 1471 3664
rect 1489 3624 1501 3664
rect 1519 3624 1531 3664
rect 1549 3624 1561 3664
rect 1597 3624 1609 3644
rect 1617 3624 1629 3644
rect 1637 3624 1649 3644
rect 1677 3624 1689 3664
rect 1699 3624 1711 3644
rect 1729 3624 1741 3644
rect 1757 3624 1769 3644
rect 1783 3624 1795 3644
rect 1805 3624 1817 3644
rect 1835 3624 1847 3644
rect 1867 3624 1879 3644
rect 1887 3624 1899 3664
rect 1939 3624 1951 3664
rect 1969 3624 1981 3664
rect 1997 3624 2009 3644
rect 2017 3624 2029 3644
rect 2037 3624 2049 3644
rect 2077 3624 2089 3644
rect 2097 3624 2109 3644
rect 2137 3624 2149 3664
rect 2157 3624 2169 3652
rect 2177 3624 2189 3664
rect 2197 3624 2209 3664
rect 2251 3624 2263 3664
rect 2271 3624 2283 3664
rect 2291 3624 2303 3652
rect 2311 3624 2323 3664
rect 2358 3624 2370 3644
rect 2380 3624 2392 3664
rect 2408 3624 2420 3664
rect 2437 3624 2449 3644
rect 2457 3624 2469 3644
rect 2511 3624 2523 3644
rect 2531 3624 2543 3644
rect 2557 3624 2569 3664
rect 2577 3624 2589 3652
rect 2597 3624 2609 3664
rect 2617 3624 2629 3664
rect 2658 3624 2670 3684
rect 2694 3624 2706 3682
rect 2771 3624 2783 3644
rect 2791 3624 2803 3644
rect 2839 3624 2851 3664
rect 2869 3624 2881 3664
rect 2897 3624 2909 3664
rect 2917 3624 2929 3652
rect 2937 3624 2949 3664
rect 2957 3624 2969 3664
rect 2997 3624 3009 3664
rect 3017 3624 3029 3652
rect 3037 3624 3049 3664
rect 3057 3624 3069 3664
rect 3100 3624 3112 3664
rect 3128 3624 3140 3664
rect 3150 3624 3162 3644
rect 3232 3624 3244 3664
rect 3260 3624 3272 3664
rect 3288 3624 3300 3664
rect 3339 3624 3351 3664
rect 3369 3624 3381 3664
rect 3419 3624 3431 3664
rect 3449 3624 3461 3664
rect 3481 3624 3493 3664
rect 3501 3624 3513 3644
rect 3533 3624 3545 3644
rect 3563 3624 3575 3644
rect 3585 3624 3597 3644
rect 3611 3624 3623 3644
rect 3639 3624 3651 3644
rect 3669 3624 3681 3644
rect 3691 3624 3703 3664
rect 3739 3624 3751 3664
rect 3769 3624 3781 3664
rect 3832 3624 3844 3664
rect 3860 3624 3872 3664
rect 3888 3624 3900 3664
rect 3917 3624 3929 3644
rect 3937 3624 3949 3644
rect 3979 3624 3991 3664
rect 4009 3624 4021 3664
rect 4057 3624 4069 3664
rect 4077 3624 4089 3652
rect 4097 3624 4109 3664
rect 4117 3624 4129 3664
rect 4161 3624 4173 3664
rect 4181 3624 4193 3644
rect 4213 3624 4225 3644
rect 4243 3624 4255 3644
rect 4265 3624 4277 3644
rect 4291 3624 4303 3644
rect 4319 3624 4331 3644
rect 4349 3624 4361 3644
rect 4371 3624 4383 3664
rect 4399 3624 4411 3664
rect 4429 3624 4441 3664
rect 4499 3624 4511 3664
rect 4529 3624 4541 3664
rect 4571 3624 4583 3664
rect 4591 3624 4603 3664
rect 4611 3624 4623 3664
rect 4631 3624 4643 3664
rect 4651 3624 4663 3664
rect 4671 3624 4683 3664
rect 4691 3624 4703 3664
rect 4711 3624 4723 3664
rect 4731 3624 4743 3664
rect 4761 3624 4773 3664
rect 4781 3624 4793 3644
rect 4813 3624 4825 3644
rect 4843 3624 4855 3644
rect 4865 3624 4877 3644
rect 4891 3624 4903 3644
rect 4919 3624 4931 3644
rect 4949 3624 4961 3644
rect 4971 3624 4983 3664
rect 4997 3624 5009 3664
rect 5017 3624 5029 3652
rect 5037 3624 5049 3664
rect 5057 3624 5069 3664
rect 5119 3624 5131 3664
rect 5149 3624 5161 3664
rect 5199 3624 5211 3664
rect 5229 3624 5241 3664
rect 5271 3624 5283 3644
rect 5291 3624 5303 3644
rect 5317 3624 5329 3664
rect 5337 3624 5349 3664
rect 5357 3624 5369 3664
rect 5377 3624 5389 3664
rect 5397 3624 5409 3664
rect 5417 3624 5429 3664
rect 5437 3624 5449 3664
rect 5457 3624 5469 3664
rect 5477 3624 5489 3664
rect 5517 3624 5529 3664
rect 5539 3624 5551 3644
rect 5569 3624 5581 3644
rect 5597 3624 5609 3644
rect 5623 3624 5635 3644
rect 5645 3624 5657 3644
rect 5675 3624 5687 3644
rect 5707 3624 5719 3644
rect 5727 3624 5739 3664
rect 5771 3624 5783 3644
rect 5791 3624 5803 3644
rect 5819 3624 5831 3664
rect 5849 3624 5861 3664
rect 5899 3624 5911 3664
rect 5929 3624 5941 3664
rect 5991 3624 6003 3644
rect 6011 3624 6023 3644
rect 6037 3624 6049 3644
rect 6057 3624 6069 3644
rect 6077 3624 6089 3644
rect 6131 3624 6143 3644
rect 6151 3624 6163 3644
rect 6171 3624 6183 3644
rect 6200 3624 6212 3664
rect 6228 3624 6240 3664
rect 6250 3624 6262 3644
rect 6297 3624 6309 3664
rect 6319 3624 6331 3644
rect 6349 3624 6361 3644
rect 6377 3624 6389 3644
rect 6403 3624 6415 3644
rect 6425 3624 6437 3644
rect 6455 3624 6467 3644
rect 6487 3624 6499 3644
rect 6507 3624 6519 3664
rect 6537 3624 6549 3664
rect 6557 3624 6569 3652
rect 6577 3624 6589 3664
rect 6597 3624 6609 3664
rect 6639 3624 6651 3664
rect 6669 3624 6681 3664
rect 29 3556 41 3596
rect 49 3556 61 3596
rect 71 3576 83 3596
rect 97 3556 109 3596
rect 119 3576 131 3596
rect 149 3576 161 3596
rect 177 3576 189 3596
rect 203 3576 215 3596
rect 225 3576 237 3596
rect 255 3576 267 3596
rect 287 3576 299 3596
rect 307 3556 319 3596
rect 339 3556 351 3596
rect 369 3556 381 3596
rect 417 3576 429 3596
rect 439 3556 451 3596
rect 459 3556 471 3596
rect 518 3576 530 3596
rect 540 3556 552 3596
rect 568 3556 580 3596
rect 619 3556 631 3596
rect 649 3556 661 3596
rect 689 3556 701 3596
rect 709 3556 721 3596
rect 731 3576 743 3596
rect 757 3576 769 3596
rect 779 3556 791 3596
rect 799 3556 811 3596
rect 839 3556 851 3596
rect 869 3556 881 3596
rect 929 3556 941 3596
rect 949 3556 961 3596
rect 971 3576 983 3596
rect 1011 3576 1023 3596
rect 1031 3576 1043 3596
rect 1069 3556 1081 3596
rect 1089 3556 1101 3596
rect 1111 3576 1123 3596
rect 1149 3556 1161 3596
rect 1169 3556 1181 3596
rect 1191 3576 1203 3596
rect 1217 3556 1229 3596
rect 1239 3576 1251 3596
rect 1269 3576 1281 3596
rect 1297 3576 1309 3596
rect 1323 3576 1335 3596
rect 1345 3576 1357 3596
rect 1375 3576 1387 3596
rect 1407 3576 1419 3596
rect 1427 3556 1439 3596
rect 1471 3576 1483 3596
rect 1491 3576 1503 3596
rect 1511 3576 1523 3596
rect 1537 3556 1549 3596
rect 1559 3576 1571 3596
rect 1589 3576 1601 3596
rect 1617 3576 1629 3596
rect 1643 3576 1655 3596
rect 1665 3576 1677 3596
rect 1695 3576 1707 3596
rect 1727 3576 1739 3596
rect 1747 3556 1759 3596
rect 1801 3556 1813 3596
rect 1821 3556 1833 3596
rect 1851 3556 1863 3596
rect 1891 3576 1903 3596
rect 1911 3576 1923 3596
rect 1951 3556 1963 3596
rect 1971 3556 1983 3596
rect 1991 3568 2003 3596
rect 2011 3556 2023 3596
rect 2037 3576 2049 3596
rect 2057 3576 2069 3596
rect 2077 3576 2089 3596
rect 2131 3576 2143 3596
rect 2151 3576 2163 3596
rect 2201 3556 2213 3596
rect 2221 3556 2233 3596
rect 2251 3556 2263 3596
rect 2291 3576 2303 3596
rect 2311 3576 2323 3596
rect 2331 3576 2343 3596
rect 2357 3556 2369 3596
rect 2379 3576 2391 3596
rect 2409 3576 2421 3596
rect 2437 3576 2449 3596
rect 2463 3576 2475 3596
rect 2485 3576 2497 3596
rect 2515 3576 2527 3596
rect 2547 3576 2559 3596
rect 2567 3556 2579 3596
rect 2597 3576 2609 3596
rect 2617 3576 2629 3596
rect 2637 3576 2649 3596
rect 2677 3556 2689 3596
rect 2697 3568 2709 3596
rect 2717 3556 2729 3596
rect 2737 3556 2749 3596
rect 2791 3576 2803 3596
rect 2811 3576 2823 3596
rect 2859 3556 2871 3596
rect 2889 3556 2901 3596
rect 2917 3556 2929 3596
rect 2937 3568 2949 3596
rect 2957 3556 2969 3596
rect 2977 3556 2989 3596
rect 3020 3556 3032 3596
rect 3048 3556 3060 3596
rect 3070 3576 3082 3596
rect 3117 3556 3129 3596
rect 3137 3556 3149 3596
rect 3212 3556 3224 3596
rect 3240 3556 3252 3596
rect 3268 3556 3280 3596
rect 3311 3576 3323 3596
rect 3331 3576 3343 3596
rect 3357 3556 3369 3596
rect 3379 3576 3391 3596
rect 3409 3576 3421 3596
rect 3437 3576 3449 3596
rect 3463 3576 3475 3596
rect 3485 3576 3497 3596
rect 3515 3576 3527 3596
rect 3547 3576 3559 3596
rect 3567 3556 3579 3596
rect 3632 3556 3644 3596
rect 3660 3556 3672 3596
rect 3688 3556 3700 3596
rect 3717 3556 3729 3596
rect 3739 3576 3751 3596
rect 3769 3576 3781 3596
rect 3797 3576 3809 3596
rect 3823 3576 3835 3596
rect 3845 3576 3857 3596
rect 3875 3576 3887 3596
rect 3907 3576 3919 3596
rect 3927 3556 3939 3596
rect 3971 3576 3983 3596
rect 3991 3576 4003 3596
rect 4017 3556 4029 3596
rect 4039 3576 4051 3596
rect 4069 3576 4081 3596
rect 4097 3576 4109 3596
rect 4123 3576 4135 3596
rect 4145 3576 4157 3596
rect 4175 3576 4187 3596
rect 4207 3576 4219 3596
rect 4227 3556 4239 3596
rect 4271 3576 4283 3596
rect 4291 3576 4303 3596
rect 4331 3576 4343 3596
rect 4351 3576 4363 3596
rect 4379 3556 4391 3596
rect 4409 3556 4421 3596
rect 4461 3556 4473 3596
rect 4481 3576 4493 3596
rect 4513 3576 4525 3596
rect 4543 3576 4555 3596
rect 4565 3576 4577 3596
rect 4591 3576 4603 3596
rect 4619 3576 4631 3596
rect 4649 3576 4661 3596
rect 4671 3556 4683 3596
rect 4711 3576 4723 3596
rect 4731 3576 4743 3596
rect 4757 3556 4769 3596
rect 4779 3576 4791 3596
rect 4809 3576 4821 3596
rect 4837 3576 4849 3596
rect 4863 3576 4875 3596
rect 4885 3576 4897 3596
rect 4915 3576 4927 3596
rect 4947 3576 4959 3596
rect 4967 3556 4979 3596
rect 5032 3556 5044 3596
rect 5060 3556 5072 3596
rect 5088 3556 5100 3596
rect 5131 3576 5143 3596
rect 5151 3576 5163 3596
rect 5177 3556 5189 3596
rect 5199 3576 5211 3596
rect 5229 3576 5241 3596
rect 5257 3576 5269 3596
rect 5283 3576 5295 3596
rect 5305 3576 5317 3596
rect 5335 3576 5347 3596
rect 5367 3576 5379 3596
rect 5387 3556 5399 3596
rect 5417 3556 5429 3596
rect 5439 3576 5451 3596
rect 5469 3576 5481 3596
rect 5497 3576 5509 3596
rect 5523 3576 5535 3596
rect 5545 3576 5557 3596
rect 5575 3576 5587 3596
rect 5607 3576 5619 3596
rect 5627 3556 5639 3596
rect 5657 3556 5669 3596
rect 5677 3568 5689 3596
rect 5697 3556 5709 3596
rect 5717 3556 5729 3596
rect 5757 3556 5769 3596
rect 5777 3568 5789 3596
rect 5797 3556 5809 3596
rect 5817 3556 5829 3596
rect 5871 3576 5883 3596
rect 5891 3576 5903 3596
rect 5952 3556 5964 3596
rect 5980 3556 5992 3596
rect 6008 3556 6020 3596
rect 6039 3556 6051 3596
rect 6069 3556 6081 3596
rect 6131 3576 6143 3596
rect 6151 3576 6163 3596
rect 6195 3576 6209 3596
rect 6217 3576 6229 3596
rect 6237 3576 6249 3596
rect 6257 3576 6269 3596
rect 6371 3576 6383 3596
rect 6391 3576 6403 3596
rect 6417 3556 6429 3596
rect 6439 3576 6451 3596
rect 6469 3576 6481 3596
rect 6497 3576 6509 3596
rect 6523 3576 6535 3596
rect 6545 3576 6557 3596
rect 6575 3576 6587 3596
rect 6607 3576 6619 3596
rect 6627 3556 6639 3596
rect 29 3144 41 3184
rect 49 3144 61 3184
rect 71 3144 83 3164
rect 97 3144 109 3184
rect 119 3144 131 3164
rect 149 3144 161 3164
rect 177 3144 189 3164
rect 203 3144 215 3164
rect 225 3144 237 3164
rect 255 3144 267 3164
rect 287 3144 299 3164
rect 307 3144 319 3184
rect 339 3144 351 3184
rect 369 3144 381 3184
rect 438 3144 450 3164
rect 460 3144 472 3184
rect 488 3144 500 3184
rect 539 3144 551 3184
rect 569 3144 581 3184
rect 597 3144 609 3164
rect 617 3144 629 3164
rect 658 3144 670 3204
rect 694 3144 706 3202
rect 759 3144 771 3184
rect 789 3144 801 3184
rect 851 3144 863 3184
rect 871 3144 883 3184
rect 891 3144 903 3172
rect 911 3144 923 3184
rect 937 3144 949 3164
rect 957 3144 969 3164
rect 997 3144 1009 3164
rect 1017 3144 1029 3164
rect 1037 3144 1049 3164
rect 1077 3144 1089 3184
rect 1097 3144 1109 3172
rect 1117 3144 1129 3184
rect 1137 3144 1149 3184
rect 1177 3144 1189 3184
rect 1197 3144 1209 3172
rect 1217 3144 1229 3184
rect 1237 3144 1249 3184
rect 1279 3144 1291 3184
rect 1309 3144 1321 3184
rect 1357 3144 1369 3184
rect 1379 3144 1391 3164
rect 1409 3144 1421 3164
rect 1437 3144 1449 3164
rect 1463 3144 1475 3164
rect 1485 3144 1497 3164
rect 1515 3144 1527 3164
rect 1547 3144 1559 3164
rect 1567 3144 1579 3184
rect 1621 3144 1633 3184
rect 1641 3144 1653 3184
rect 1671 3144 1683 3184
rect 1718 3144 1730 3164
rect 1740 3144 1752 3184
rect 1768 3144 1780 3184
rect 1834 3144 1846 3202
rect 1870 3144 1882 3204
rect 1900 3144 1912 3184
rect 1928 3144 1940 3184
rect 1950 3144 1962 3164
rect 2001 3144 2013 3184
rect 2021 3144 2033 3164
rect 2053 3144 2065 3164
rect 2083 3144 2095 3164
rect 2105 3144 2117 3164
rect 2131 3144 2143 3164
rect 2159 3144 2171 3164
rect 2189 3144 2201 3164
rect 2211 3144 2223 3184
rect 2239 3144 2251 3184
rect 2269 3144 2281 3184
rect 2317 3144 2329 3164
rect 2337 3144 2349 3164
rect 2357 3144 2369 3164
rect 2411 3144 2423 3164
rect 2431 3144 2443 3164
rect 2451 3144 2463 3164
rect 2491 3144 2503 3184
rect 2511 3144 2523 3184
rect 2531 3144 2543 3172
rect 2551 3144 2563 3184
rect 2577 3144 2589 3164
rect 2597 3144 2609 3164
rect 2641 3144 2653 3184
rect 2661 3144 2673 3164
rect 2693 3144 2705 3164
rect 2723 3144 2735 3164
rect 2745 3144 2757 3164
rect 2771 3144 2783 3164
rect 2799 3144 2811 3164
rect 2829 3144 2841 3164
rect 2851 3144 2863 3184
rect 2879 3144 2891 3184
rect 2909 3144 2921 3184
rect 2979 3144 2991 3184
rect 3009 3144 3021 3184
rect 3051 3144 3063 3184
rect 3071 3144 3083 3184
rect 3091 3144 3103 3172
rect 3111 3144 3123 3184
rect 3159 3144 3171 3184
rect 3189 3144 3201 3184
rect 3231 3144 3243 3164
rect 3251 3144 3263 3164
rect 3291 3144 3303 3184
rect 3311 3144 3323 3184
rect 3331 3144 3343 3172
rect 3351 3144 3363 3184
rect 3377 3144 3389 3164
rect 3397 3144 3409 3164
rect 3451 3144 3463 3164
rect 3471 3144 3483 3164
rect 3491 3144 3503 3164
rect 3538 3144 3550 3164
rect 3560 3144 3572 3184
rect 3588 3144 3600 3184
rect 3631 3144 3643 3164
rect 3651 3144 3663 3164
rect 3671 3144 3683 3164
rect 3697 3144 3709 3184
rect 3719 3144 3731 3164
rect 3749 3144 3761 3164
rect 3777 3144 3789 3164
rect 3803 3144 3815 3164
rect 3825 3144 3837 3164
rect 3855 3144 3867 3164
rect 3887 3144 3899 3164
rect 3907 3144 3919 3184
rect 3940 3144 3952 3184
rect 3968 3144 3980 3184
rect 3996 3144 4008 3184
rect 4092 3144 4104 3184
rect 4120 3144 4132 3184
rect 4148 3144 4160 3184
rect 4181 3144 4193 3184
rect 4201 3144 4213 3164
rect 4233 3144 4245 3164
rect 4263 3144 4275 3164
rect 4285 3144 4297 3164
rect 4311 3144 4323 3164
rect 4339 3144 4351 3164
rect 4369 3144 4381 3164
rect 4391 3144 4403 3184
rect 4417 3144 4429 3164
rect 4437 3144 4449 3164
rect 4457 3144 4469 3164
rect 4500 3144 4512 3184
rect 4528 3144 4540 3184
rect 4556 3144 4568 3184
rect 4617 3144 4629 3164
rect 4637 3144 4649 3164
rect 4657 3144 4669 3164
rect 4697 3144 4709 3164
rect 4717 3144 4729 3164
rect 4737 3144 4749 3164
rect 4777 3144 4789 3164
rect 4797 3144 4809 3164
rect 4840 3144 4852 3184
rect 4868 3144 4880 3184
rect 4896 3144 4908 3184
rect 4960 3144 4972 3184
rect 4988 3144 5000 3184
rect 5010 3144 5022 3164
rect 5057 3144 5069 3184
rect 5079 3144 5091 3164
rect 5109 3144 5121 3164
rect 5137 3144 5149 3164
rect 5163 3144 5175 3164
rect 5185 3144 5197 3164
rect 5215 3144 5227 3164
rect 5247 3144 5259 3164
rect 5267 3144 5279 3184
rect 5311 3144 5323 3164
rect 5331 3144 5343 3164
rect 5357 3152 5369 3172
rect 5377 3152 5389 3172
rect 5407 3152 5419 3184
rect 5437 3152 5449 3192
rect 5491 3144 5503 3164
rect 5511 3144 5523 3164
rect 5541 3144 5553 3184
rect 5561 3144 5573 3164
rect 5593 3144 5605 3164
rect 5623 3144 5635 3164
rect 5645 3144 5657 3164
rect 5671 3144 5683 3164
rect 5699 3144 5711 3164
rect 5729 3144 5741 3164
rect 5751 3144 5763 3184
rect 5791 3144 5803 3184
rect 5811 3144 5823 3184
rect 5831 3144 5843 3172
rect 5851 3144 5863 3184
rect 5891 3144 5903 3164
rect 5911 3144 5923 3164
rect 5958 3144 5970 3164
rect 5980 3144 5992 3184
rect 6008 3144 6020 3184
rect 6037 3144 6049 3184
rect 6057 3144 6069 3172
rect 6077 3144 6089 3184
rect 6097 3144 6109 3184
rect 6159 3144 6171 3184
rect 6189 3144 6201 3184
rect 6238 3144 6250 3164
rect 6260 3144 6272 3184
rect 6288 3144 6300 3184
rect 6339 3144 6351 3184
rect 6369 3144 6381 3184
rect 6397 3144 6409 3184
rect 6417 3144 6429 3172
rect 6437 3144 6449 3184
rect 6457 3144 6469 3184
rect 6497 3144 6509 3184
rect 6519 3144 6531 3164
rect 6549 3144 6561 3164
rect 6577 3144 6589 3164
rect 6603 3144 6615 3164
rect 6625 3144 6637 3164
rect 6655 3144 6667 3164
rect 6687 3144 6699 3164
rect 6707 3144 6719 3184
rect 17 3076 29 3116
rect 37 3076 49 3116
rect 57 3076 69 3116
rect 77 3076 89 3116
rect 97 3076 109 3116
rect 117 3076 129 3116
rect 137 3076 149 3116
rect 157 3076 169 3116
rect 177 3076 189 3116
rect 229 3076 241 3116
rect 249 3076 261 3116
rect 271 3096 283 3116
rect 301 3076 313 3116
rect 321 3096 333 3116
rect 353 3096 365 3116
rect 383 3096 395 3116
rect 405 3096 417 3116
rect 431 3096 443 3116
rect 459 3096 471 3116
rect 489 3096 501 3116
rect 511 3076 523 3116
rect 559 3076 571 3116
rect 589 3076 601 3116
rect 619 3076 631 3116
rect 649 3076 661 3116
rect 711 3076 723 3116
rect 731 3076 743 3116
rect 751 3088 763 3116
rect 771 3076 783 3116
rect 819 3076 831 3116
rect 849 3076 861 3116
rect 899 3076 911 3116
rect 929 3076 941 3116
rect 960 3076 972 3116
rect 988 3076 1000 3116
rect 1010 3096 1022 3116
rect 1057 3076 1069 3116
rect 1079 3096 1091 3116
rect 1109 3096 1121 3116
rect 1137 3096 1149 3116
rect 1163 3096 1175 3116
rect 1185 3096 1197 3116
rect 1215 3096 1227 3116
rect 1247 3096 1259 3116
rect 1267 3076 1279 3116
rect 1319 3076 1331 3116
rect 1349 3076 1361 3116
rect 1377 3076 1389 3116
rect 1399 3096 1411 3116
rect 1429 3096 1441 3116
rect 1457 3096 1469 3116
rect 1483 3096 1495 3116
rect 1505 3096 1517 3116
rect 1535 3096 1547 3116
rect 1567 3096 1579 3116
rect 1587 3076 1599 3116
rect 1631 3096 1643 3116
rect 1651 3096 1663 3116
rect 1691 3076 1703 3116
rect 1711 3076 1723 3116
rect 1731 3088 1743 3116
rect 1751 3076 1763 3116
rect 1791 3096 1803 3116
rect 1811 3096 1823 3116
rect 1831 3096 1843 3116
rect 1881 3076 1893 3116
rect 1901 3076 1913 3116
rect 1931 3076 1943 3116
rect 1957 3076 1969 3116
rect 1977 3088 1989 3116
rect 1997 3076 2009 3116
rect 2017 3076 2029 3116
rect 2078 3096 2090 3116
rect 2100 3076 2112 3116
rect 2128 3076 2140 3116
rect 2159 3076 2171 3116
rect 2189 3076 2201 3116
rect 2251 3096 2263 3116
rect 2271 3096 2283 3116
rect 2297 3076 2309 3116
rect 2327 3076 2339 3116
rect 2347 3076 2359 3116
rect 2401 3076 2413 3116
rect 2421 3096 2433 3116
rect 2453 3096 2465 3116
rect 2483 3096 2495 3116
rect 2505 3096 2517 3116
rect 2531 3096 2543 3116
rect 2559 3096 2571 3116
rect 2589 3096 2601 3116
rect 2611 3076 2623 3116
rect 2637 3096 2649 3116
rect 2657 3096 2669 3116
rect 2697 3096 2709 3116
rect 2717 3096 2729 3116
rect 2737 3096 2749 3116
rect 2791 3096 2803 3116
rect 2811 3096 2823 3116
rect 2851 3076 2863 3116
rect 2871 3076 2883 3116
rect 2891 3088 2903 3116
rect 2911 3076 2923 3116
rect 2937 3076 2949 3116
rect 2957 3076 2969 3116
rect 3034 3058 3046 3116
rect 3070 3056 3082 3116
rect 3119 3076 3131 3116
rect 3149 3076 3161 3116
rect 3191 3076 3203 3116
rect 3211 3076 3223 3116
rect 3231 3088 3243 3116
rect 3251 3076 3263 3116
rect 3279 3076 3291 3116
rect 3309 3076 3321 3116
rect 3359 3076 3371 3116
rect 3389 3076 3401 3116
rect 3437 3076 3449 3116
rect 3457 3088 3469 3116
rect 3477 3076 3489 3116
rect 3497 3076 3509 3116
rect 3537 3076 3549 3116
rect 3567 3076 3579 3116
rect 3587 3076 3599 3116
rect 3672 3076 3684 3116
rect 3700 3076 3712 3116
rect 3728 3076 3740 3116
rect 3771 3076 3783 3116
rect 3791 3076 3803 3116
rect 3811 3076 3823 3116
rect 3841 3076 3853 3116
rect 3861 3096 3873 3116
rect 3893 3096 3905 3116
rect 3923 3096 3935 3116
rect 3945 3096 3957 3116
rect 3971 3096 3983 3116
rect 3999 3096 4011 3116
rect 4029 3096 4041 3116
rect 4051 3076 4063 3116
rect 4077 3076 4089 3116
rect 4097 3088 4109 3116
rect 4117 3076 4129 3116
rect 4137 3076 4149 3116
rect 4214 3058 4226 3116
rect 4250 3056 4262 3116
rect 4281 3076 4293 3116
rect 4301 3096 4313 3116
rect 4333 3096 4345 3116
rect 4363 3096 4375 3116
rect 4385 3096 4397 3116
rect 4411 3096 4423 3116
rect 4439 3096 4451 3116
rect 4469 3096 4481 3116
rect 4491 3076 4503 3116
rect 4531 3076 4543 3116
rect 4551 3076 4563 3104
rect 4571 3076 4583 3116
rect 4591 3086 4603 3116
rect 4611 3076 4623 3116
rect 4651 3096 4663 3116
rect 4671 3096 4683 3116
rect 4711 3068 4723 3108
rect 4741 3076 4753 3108
rect 4771 3088 4783 3108
rect 4791 3088 4803 3108
rect 4820 3076 4832 3116
rect 4848 3076 4860 3116
rect 4876 3076 4888 3116
rect 4951 3096 4963 3116
rect 4971 3096 4983 3116
rect 5000 3076 5012 3116
rect 5028 3076 5040 3116
rect 5056 3076 5068 3116
rect 5117 3096 5129 3116
rect 5137 3096 5149 3116
rect 5177 3096 5189 3116
rect 5197 3096 5209 3116
rect 5217 3096 5229 3116
rect 5261 3076 5273 3116
rect 5281 3096 5293 3116
rect 5313 3096 5325 3116
rect 5343 3096 5355 3116
rect 5365 3096 5377 3116
rect 5391 3096 5403 3116
rect 5419 3096 5431 3116
rect 5449 3096 5461 3116
rect 5471 3076 5483 3116
rect 5511 3096 5523 3116
rect 5531 3096 5543 3116
rect 5551 3096 5563 3116
rect 5577 3076 5589 3116
rect 5597 3088 5609 3116
rect 5617 3076 5629 3116
rect 5637 3076 5649 3116
rect 5714 3058 5726 3116
rect 5750 3056 5762 3116
rect 5791 3076 5803 3116
rect 5811 3076 5823 3104
rect 5831 3076 5843 3116
rect 5851 3086 5863 3116
rect 5871 3076 5883 3116
rect 5897 3096 5909 3116
rect 5917 3096 5929 3116
rect 5957 3088 5969 3108
rect 5977 3088 5989 3108
rect 6007 3076 6019 3108
rect 6037 3068 6049 3108
rect 6098 3096 6110 3116
rect 6120 3076 6132 3116
rect 6148 3076 6160 3116
rect 6191 3096 6203 3116
rect 6211 3096 6223 3116
rect 6231 3096 6243 3116
rect 6257 3096 6269 3116
rect 6277 3096 6289 3116
rect 6352 3076 6364 3116
rect 6380 3076 6392 3116
rect 6408 3076 6420 3116
rect 6451 3096 6463 3116
rect 6471 3096 6483 3116
rect 6497 3096 6509 3116
rect 6517 3096 6529 3116
rect 6557 3076 6569 3116
rect 6577 3088 6589 3116
rect 6597 3076 6609 3116
rect 6617 3076 6629 3116
rect 17 2664 29 2684
rect 37 2664 49 2684
rect 91 2664 103 2684
rect 111 2664 123 2684
rect 131 2664 143 2684
rect 161 2664 173 2704
rect 181 2664 193 2684
rect 213 2664 225 2684
rect 243 2664 255 2684
rect 265 2664 277 2684
rect 291 2664 303 2684
rect 319 2664 331 2684
rect 349 2664 361 2684
rect 371 2664 383 2704
rect 397 2664 409 2684
rect 417 2664 429 2684
rect 471 2664 483 2684
rect 491 2664 503 2684
rect 511 2664 523 2684
rect 541 2664 553 2704
rect 561 2664 573 2684
rect 593 2664 605 2684
rect 623 2664 635 2684
rect 645 2664 657 2684
rect 671 2664 683 2684
rect 699 2664 711 2684
rect 729 2664 741 2684
rect 751 2664 763 2704
rect 789 2664 801 2704
rect 809 2664 821 2704
rect 831 2664 843 2684
rect 857 2664 869 2704
rect 877 2664 889 2704
rect 897 2664 909 2704
rect 939 2664 951 2704
rect 969 2664 981 2704
rect 1019 2664 1031 2704
rect 1049 2664 1061 2704
rect 1097 2664 1109 2684
rect 1117 2664 1129 2684
rect 1160 2664 1172 2704
rect 1188 2664 1200 2704
rect 1216 2664 1228 2704
rect 1298 2664 1310 2684
rect 1320 2664 1332 2704
rect 1348 2664 1360 2704
rect 1391 2664 1403 2684
rect 1411 2664 1423 2684
rect 1451 2664 1463 2704
rect 1471 2664 1483 2704
rect 1491 2664 1503 2692
rect 1511 2664 1523 2704
rect 1537 2664 1549 2684
rect 1557 2664 1569 2684
rect 1577 2664 1589 2684
rect 1619 2664 1631 2704
rect 1649 2664 1661 2704
rect 1697 2664 1709 2684
rect 1717 2664 1729 2684
rect 1737 2664 1749 2684
rect 1791 2664 1803 2704
rect 1811 2664 1823 2704
rect 1831 2664 1843 2692
rect 1851 2664 1863 2704
rect 1877 2664 1889 2684
rect 1897 2664 1909 2684
rect 1917 2664 1929 2684
rect 1937 2664 1949 2704
rect 1977 2664 1989 2704
rect 1997 2664 2009 2692
rect 2017 2664 2029 2704
rect 2037 2664 2049 2704
rect 2098 2664 2110 2684
rect 2120 2664 2132 2704
rect 2148 2664 2160 2704
rect 2181 2664 2193 2704
rect 2201 2664 2213 2684
rect 2233 2664 2245 2684
rect 2263 2664 2275 2684
rect 2285 2664 2297 2684
rect 2311 2664 2323 2684
rect 2339 2664 2351 2684
rect 2369 2664 2381 2684
rect 2391 2664 2403 2704
rect 2419 2664 2431 2704
rect 2449 2664 2461 2704
rect 2497 2664 2509 2684
rect 2517 2664 2529 2684
rect 2571 2664 2583 2684
rect 2591 2664 2603 2684
rect 2621 2664 2633 2704
rect 2641 2664 2653 2684
rect 2673 2664 2685 2684
rect 2703 2664 2715 2684
rect 2725 2664 2737 2684
rect 2751 2664 2763 2684
rect 2779 2664 2791 2684
rect 2809 2664 2821 2684
rect 2831 2664 2843 2704
rect 2857 2664 2869 2704
rect 2877 2664 2889 2692
rect 2897 2664 2909 2704
rect 2917 2664 2929 2704
rect 2978 2664 2990 2684
rect 3000 2664 3012 2704
rect 3028 2664 3040 2704
rect 3057 2664 3069 2704
rect 3079 2664 3091 2684
rect 3109 2664 3121 2684
rect 3137 2664 3149 2684
rect 3163 2664 3175 2684
rect 3185 2664 3197 2684
rect 3215 2664 3227 2684
rect 3247 2664 3259 2684
rect 3267 2664 3279 2704
rect 3297 2664 3309 2684
rect 3317 2664 3329 2684
rect 3357 2664 3369 2704
rect 3377 2664 3389 2694
rect 3397 2664 3409 2704
rect 3417 2676 3429 2704
rect 3437 2664 3449 2704
rect 3477 2664 3489 2704
rect 3497 2664 3509 2692
rect 3517 2664 3529 2704
rect 3537 2664 3549 2704
rect 3591 2664 3603 2704
rect 3611 2676 3623 2704
rect 3631 2664 3643 2704
rect 3651 2664 3663 2694
rect 3671 2664 3683 2704
rect 3697 2664 3709 2704
rect 3717 2664 3729 2692
rect 3737 2664 3749 2704
rect 3757 2664 3769 2704
rect 3811 2664 3823 2704
rect 3831 2676 3843 2704
rect 3851 2664 3863 2704
rect 3871 2664 3883 2694
rect 3891 2664 3903 2704
rect 3931 2664 3943 2684
rect 3951 2664 3963 2684
rect 3977 2664 3989 2684
rect 3997 2664 4009 2684
rect 4017 2664 4029 2684
rect 4057 2664 4069 2684
rect 4077 2664 4089 2684
rect 4097 2664 4109 2684
rect 4158 2664 4170 2684
rect 4180 2664 4192 2704
rect 4208 2664 4220 2704
rect 4237 2664 4249 2704
rect 4257 2664 4269 2692
rect 4277 2664 4289 2704
rect 4297 2664 4309 2704
rect 4374 2664 4386 2722
rect 4410 2664 4422 2724
rect 4441 2664 4453 2704
rect 4461 2664 4473 2684
rect 4493 2664 4505 2684
rect 4523 2664 4535 2684
rect 4545 2664 4557 2684
rect 4571 2664 4583 2684
rect 4599 2664 4611 2684
rect 4629 2664 4641 2684
rect 4651 2664 4663 2704
rect 4677 2664 4689 2684
rect 4697 2664 4709 2684
rect 4737 2664 4749 2684
rect 4757 2664 4769 2684
rect 4777 2664 4789 2684
rect 4817 2664 4829 2704
rect 4837 2664 4849 2692
rect 4857 2664 4869 2704
rect 4877 2664 4889 2704
rect 4931 2664 4943 2684
rect 4951 2664 4963 2684
rect 4971 2664 4983 2684
rect 5011 2664 5023 2704
rect 5031 2676 5043 2704
rect 5051 2664 5063 2704
rect 5071 2664 5083 2694
rect 5091 2664 5103 2704
rect 5120 2664 5132 2704
rect 5148 2664 5160 2704
rect 5170 2664 5182 2684
rect 5217 2664 5229 2684
rect 5239 2664 5251 2704
rect 5259 2664 5271 2704
rect 5297 2664 5309 2704
rect 5317 2664 5329 2692
rect 5337 2664 5349 2704
rect 5357 2664 5369 2704
rect 5411 2664 5423 2704
rect 5431 2676 5443 2704
rect 5451 2664 5463 2704
rect 5471 2664 5483 2694
rect 5491 2664 5503 2704
rect 5531 2664 5543 2684
rect 5551 2664 5563 2684
rect 5581 2664 5593 2704
rect 5601 2664 5613 2684
rect 5633 2664 5645 2684
rect 5663 2664 5675 2684
rect 5685 2664 5697 2684
rect 5711 2664 5723 2684
rect 5739 2664 5751 2684
rect 5769 2664 5781 2684
rect 5791 2664 5803 2704
rect 5817 2672 5829 2692
rect 5837 2672 5849 2692
rect 5867 2672 5879 2704
rect 5897 2672 5909 2712
rect 5937 2672 5949 2692
rect 5957 2672 5969 2692
rect 5987 2672 5999 2704
rect 6017 2672 6029 2712
rect 6057 2672 6069 2692
rect 6077 2672 6089 2692
rect 6107 2672 6119 2704
rect 6137 2672 6149 2712
rect 6201 2664 6213 2704
rect 6221 2664 6233 2704
rect 6251 2664 6263 2704
rect 6291 2664 6303 2704
rect 6311 2664 6323 2704
rect 6331 2664 6343 2704
rect 6357 2664 6369 2704
rect 6387 2664 6399 2704
rect 6407 2664 6419 2704
rect 6457 2664 6469 2704
rect 6479 2664 6491 2684
rect 6509 2664 6521 2684
rect 6537 2664 6549 2684
rect 6563 2664 6575 2684
rect 6585 2664 6597 2684
rect 6615 2664 6627 2684
rect 6647 2664 6659 2684
rect 6667 2664 6679 2704
rect 17 2596 29 2636
rect 39 2616 51 2636
rect 69 2616 81 2636
rect 97 2616 109 2636
rect 123 2616 135 2636
rect 145 2616 157 2636
rect 175 2616 187 2636
rect 207 2616 219 2636
rect 227 2596 239 2636
rect 269 2596 281 2636
rect 289 2596 301 2636
rect 311 2616 323 2636
rect 337 2596 349 2636
rect 359 2616 371 2636
rect 389 2616 401 2636
rect 417 2616 429 2636
rect 443 2616 455 2636
rect 465 2616 477 2636
rect 495 2616 507 2636
rect 527 2616 539 2636
rect 547 2596 559 2636
rect 598 2616 610 2636
rect 620 2596 632 2636
rect 648 2596 660 2636
rect 679 2596 691 2636
rect 709 2596 721 2636
rect 779 2596 791 2636
rect 809 2596 821 2636
rect 851 2596 863 2636
rect 871 2596 883 2636
rect 891 2596 903 2636
rect 911 2596 923 2636
rect 931 2596 943 2636
rect 951 2596 963 2636
rect 971 2596 983 2636
rect 991 2596 1003 2636
rect 1011 2596 1023 2636
rect 1037 2596 1049 2636
rect 1059 2616 1071 2636
rect 1089 2616 1101 2636
rect 1117 2616 1129 2636
rect 1143 2616 1155 2636
rect 1165 2616 1177 2636
rect 1195 2616 1207 2636
rect 1227 2616 1239 2636
rect 1247 2596 1259 2636
rect 1299 2596 1311 2636
rect 1329 2596 1341 2636
rect 1357 2616 1369 2636
rect 1377 2616 1389 2636
rect 1397 2616 1409 2636
rect 1437 2616 1449 2636
rect 1457 2616 1469 2636
rect 1511 2596 1523 2636
rect 1531 2596 1543 2636
rect 1551 2608 1563 2636
rect 1571 2596 1583 2636
rect 1601 2596 1613 2636
rect 1621 2616 1633 2636
rect 1653 2616 1665 2636
rect 1683 2616 1695 2636
rect 1705 2616 1717 2636
rect 1731 2616 1743 2636
rect 1759 2616 1771 2636
rect 1789 2616 1801 2636
rect 1811 2596 1823 2636
rect 1837 2616 1849 2636
rect 1857 2616 1869 2636
rect 1897 2616 1909 2636
rect 1917 2616 1929 2636
rect 1957 2596 1969 2636
rect 1977 2606 1989 2636
rect 1997 2596 2009 2636
rect 2017 2596 2029 2624
rect 2037 2596 2049 2636
rect 2077 2616 2089 2636
rect 2097 2616 2109 2636
rect 2117 2616 2129 2636
rect 2157 2608 2169 2628
rect 2177 2608 2189 2628
rect 2207 2596 2219 2628
rect 2237 2588 2249 2628
rect 2277 2608 2289 2628
rect 2297 2608 2309 2628
rect 2327 2596 2339 2628
rect 2357 2588 2369 2628
rect 2401 2596 2413 2636
rect 2421 2616 2433 2636
rect 2453 2616 2465 2636
rect 2483 2616 2495 2636
rect 2505 2616 2517 2636
rect 2531 2616 2543 2636
rect 2559 2616 2571 2636
rect 2589 2616 2601 2636
rect 2611 2596 2623 2636
rect 2637 2608 2649 2628
rect 2657 2608 2669 2628
rect 2687 2596 2699 2628
rect 2717 2588 2729 2628
rect 2771 2616 2783 2636
rect 2791 2616 2803 2636
rect 2811 2616 2823 2636
rect 2851 2588 2863 2628
rect 2881 2596 2893 2628
rect 2911 2608 2923 2628
rect 2931 2608 2943 2628
rect 2971 2596 2983 2636
rect 2991 2596 3003 2624
rect 3011 2596 3023 2636
rect 3031 2606 3043 2636
rect 3051 2596 3063 2636
rect 3091 2616 3103 2636
rect 3111 2616 3123 2636
rect 3141 2596 3153 2636
rect 3161 2616 3173 2636
rect 3193 2616 3205 2636
rect 3223 2616 3235 2636
rect 3245 2616 3257 2636
rect 3271 2616 3283 2636
rect 3299 2616 3311 2636
rect 3329 2616 3341 2636
rect 3351 2596 3363 2636
rect 3377 2616 3389 2636
rect 3397 2616 3409 2636
rect 3417 2616 3429 2636
rect 3479 2596 3491 2636
rect 3509 2596 3521 2636
rect 3537 2616 3549 2636
rect 3557 2616 3569 2636
rect 3598 2576 3610 2636
rect 3634 2578 3646 2636
rect 3698 2576 3710 2636
rect 3734 2578 3746 2636
rect 3834 2578 3846 2636
rect 3870 2576 3882 2636
rect 3897 2596 3909 2636
rect 3917 2608 3929 2636
rect 3937 2596 3949 2636
rect 3957 2596 3969 2636
rect 4000 2596 4012 2636
rect 4028 2596 4040 2636
rect 4050 2616 4062 2636
rect 4111 2616 4123 2636
rect 4131 2616 4143 2636
rect 4151 2616 4163 2636
rect 4191 2596 4203 2636
rect 4211 2596 4223 2624
rect 4231 2596 4243 2636
rect 4251 2606 4263 2636
rect 4271 2596 4283 2636
rect 4301 2596 4313 2636
rect 4321 2616 4333 2636
rect 4353 2616 4365 2636
rect 4383 2616 4395 2636
rect 4405 2616 4417 2636
rect 4431 2616 4443 2636
rect 4459 2616 4471 2636
rect 4489 2616 4501 2636
rect 4511 2596 4523 2636
rect 4551 2616 4563 2636
rect 4571 2616 4583 2636
rect 4611 2596 4623 2636
rect 4631 2596 4643 2624
rect 4651 2596 4663 2636
rect 4671 2606 4683 2636
rect 4691 2596 4703 2636
rect 4717 2608 4729 2628
rect 4737 2608 4749 2628
rect 4767 2596 4779 2628
rect 4797 2588 4809 2628
rect 4837 2596 4849 2636
rect 4859 2616 4871 2636
rect 4889 2616 4901 2636
rect 4917 2616 4929 2636
rect 4943 2616 4955 2636
rect 4965 2616 4977 2636
rect 4995 2616 5007 2636
rect 5027 2616 5039 2636
rect 5047 2596 5059 2636
rect 5077 2616 5089 2636
rect 5097 2616 5109 2636
rect 5137 2596 5149 2636
rect 5157 2606 5169 2636
rect 5177 2596 5189 2636
rect 5197 2596 5209 2624
rect 5217 2596 5229 2636
rect 5257 2596 5269 2636
rect 5277 2608 5289 2636
rect 5297 2596 5309 2636
rect 5317 2596 5329 2636
rect 5357 2616 5369 2636
rect 5377 2616 5389 2636
rect 5397 2616 5409 2636
rect 5451 2616 5463 2636
rect 5471 2616 5483 2636
rect 5491 2616 5503 2636
rect 5517 2596 5529 2636
rect 5537 2596 5549 2636
rect 5557 2596 5569 2636
rect 5577 2596 5589 2636
rect 5597 2596 5609 2636
rect 5617 2596 5629 2636
rect 5637 2596 5649 2636
rect 5657 2596 5669 2636
rect 5677 2596 5689 2636
rect 5731 2616 5743 2636
rect 5751 2616 5763 2636
rect 5771 2616 5783 2636
rect 5797 2596 5809 2636
rect 5817 2608 5829 2636
rect 5837 2596 5849 2636
rect 5857 2596 5869 2636
rect 5911 2596 5923 2636
rect 5931 2596 5943 2624
rect 5951 2596 5963 2636
rect 5971 2606 5983 2636
rect 5991 2596 6003 2636
rect 6031 2616 6043 2636
rect 6051 2616 6063 2636
rect 6077 2596 6089 2636
rect 6099 2616 6111 2636
rect 6129 2616 6141 2636
rect 6157 2616 6169 2636
rect 6183 2616 6195 2636
rect 6205 2616 6217 2636
rect 6235 2616 6247 2636
rect 6267 2616 6279 2636
rect 6287 2596 6299 2636
rect 6352 2596 6364 2636
rect 6380 2596 6392 2636
rect 6408 2596 6420 2636
rect 6437 2596 6449 2636
rect 6457 2596 6469 2636
rect 6477 2596 6489 2636
rect 6517 2616 6529 2636
rect 6537 2616 6549 2636
rect 6580 2596 6592 2636
rect 6608 2596 6620 2636
rect 6636 2596 6648 2636
rect 21 2184 33 2224
rect 41 2184 53 2204
rect 73 2184 85 2204
rect 103 2184 115 2204
rect 125 2184 137 2204
rect 151 2184 163 2204
rect 179 2184 191 2204
rect 209 2184 221 2204
rect 231 2184 243 2224
rect 269 2184 281 2224
rect 289 2184 301 2224
rect 311 2184 323 2204
rect 351 2184 363 2224
rect 371 2184 383 2224
rect 411 2184 423 2204
rect 431 2184 443 2204
rect 471 2184 483 2204
rect 491 2184 503 2204
rect 511 2184 523 2204
rect 537 2184 549 2224
rect 557 2184 569 2212
rect 577 2184 589 2224
rect 597 2184 609 2224
rect 661 2184 673 2224
rect 681 2184 693 2224
rect 711 2184 723 2224
rect 738 2184 750 2244
rect 774 2184 786 2242
rect 839 2184 851 2224
rect 869 2184 881 2224
rect 917 2184 929 2224
rect 939 2184 951 2204
rect 969 2184 981 2204
rect 997 2184 1009 2204
rect 1023 2184 1035 2204
rect 1045 2184 1057 2204
rect 1075 2184 1087 2204
rect 1107 2184 1119 2204
rect 1127 2184 1139 2224
rect 1157 2184 1169 2204
rect 1177 2184 1189 2204
rect 1221 2184 1233 2224
rect 1241 2184 1253 2204
rect 1273 2184 1285 2204
rect 1303 2184 1315 2204
rect 1325 2184 1337 2204
rect 1351 2184 1363 2204
rect 1379 2184 1391 2204
rect 1409 2184 1421 2204
rect 1431 2184 1443 2224
rect 1471 2184 1483 2204
rect 1491 2184 1503 2204
rect 1517 2184 1529 2224
rect 1537 2184 1549 2214
rect 1557 2184 1569 2224
rect 1577 2196 1589 2224
rect 1597 2184 1609 2224
rect 1637 2184 1649 2224
rect 1657 2184 1669 2212
rect 1677 2184 1689 2224
rect 1697 2184 1709 2224
rect 1751 2184 1763 2204
rect 1771 2184 1783 2204
rect 1791 2184 1803 2204
rect 1831 2184 1843 2204
rect 1851 2184 1863 2204
rect 1871 2184 1883 2204
rect 1911 2184 1923 2224
rect 1931 2196 1943 2224
rect 1951 2184 1963 2224
rect 1971 2184 1983 2214
rect 1991 2184 2003 2224
rect 2031 2184 2043 2204
rect 2051 2184 2063 2204
rect 2081 2184 2093 2224
rect 2101 2184 2113 2204
rect 2133 2184 2145 2204
rect 2163 2184 2175 2204
rect 2185 2184 2197 2204
rect 2211 2184 2223 2204
rect 2239 2184 2251 2204
rect 2269 2184 2281 2204
rect 2291 2184 2303 2224
rect 2331 2184 2343 2204
rect 2351 2184 2363 2204
rect 2371 2184 2383 2204
rect 2397 2184 2409 2224
rect 2417 2184 2429 2212
rect 2437 2184 2449 2224
rect 2457 2184 2469 2224
rect 2534 2184 2546 2242
rect 2570 2184 2582 2244
rect 2618 2184 2630 2204
rect 2640 2184 2652 2224
rect 2668 2184 2680 2224
rect 2697 2184 2709 2224
rect 2717 2184 2729 2212
rect 2737 2184 2749 2224
rect 2757 2184 2769 2224
rect 2811 2184 2823 2204
rect 2831 2184 2843 2204
rect 2851 2184 2863 2204
rect 2877 2184 2889 2224
rect 2899 2184 2911 2204
rect 2929 2184 2941 2204
rect 2957 2184 2969 2204
rect 2983 2184 2995 2204
rect 3005 2184 3017 2204
rect 3035 2184 3047 2204
rect 3067 2184 3079 2204
rect 3087 2184 3099 2224
rect 3117 2184 3129 2224
rect 3137 2184 3149 2212
rect 3157 2184 3169 2224
rect 3177 2184 3189 2224
rect 3231 2184 3243 2224
rect 3251 2196 3263 2224
rect 3271 2184 3283 2224
rect 3291 2184 3303 2214
rect 3311 2184 3323 2224
rect 3351 2184 3363 2204
rect 3371 2184 3383 2204
rect 3391 2184 3403 2204
rect 3431 2184 3443 2204
rect 3451 2184 3463 2204
rect 3491 2184 3503 2204
rect 3511 2184 3523 2204
rect 3531 2184 3543 2204
rect 3561 2184 3573 2224
rect 3581 2184 3593 2204
rect 3613 2184 3625 2204
rect 3643 2184 3655 2204
rect 3665 2184 3677 2204
rect 3691 2184 3703 2204
rect 3719 2184 3731 2204
rect 3749 2184 3761 2204
rect 3771 2184 3783 2224
rect 3799 2184 3811 2224
rect 3829 2184 3841 2224
rect 3878 2184 3890 2244
rect 3914 2184 3926 2242
rect 3977 2192 3989 2212
rect 3997 2192 4009 2212
rect 4027 2192 4039 2224
rect 4057 2192 4069 2232
rect 4097 2192 4109 2212
rect 4117 2192 4129 2212
rect 4147 2192 4159 2224
rect 4177 2192 4189 2232
rect 4217 2192 4229 2212
rect 4237 2192 4249 2212
rect 4267 2192 4279 2224
rect 4297 2192 4309 2232
rect 4337 2184 4349 2204
rect 4359 2184 4371 2224
rect 4379 2184 4391 2224
rect 4431 2184 4443 2204
rect 4451 2184 4463 2204
rect 4471 2184 4483 2204
rect 4497 2192 4509 2212
rect 4517 2192 4529 2212
rect 4547 2192 4559 2224
rect 4577 2192 4589 2232
rect 4631 2192 4643 2232
rect 4661 2192 4673 2224
rect 4691 2192 4703 2212
rect 4711 2192 4723 2212
rect 4737 2192 4749 2212
rect 4757 2192 4769 2212
rect 4787 2192 4799 2224
rect 4817 2192 4829 2232
rect 4857 2184 4869 2204
rect 4877 2184 4889 2204
rect 4897 2184 4909 2204
rect 4937 2192 4949 2212
rect 4957 2192 4969 2212
rect 4987 2192 4999 2224
rect 5017 2192 5029 2232
rect 5078 2184 5090 2204
rect 5100 2184 5112 2224
rect 5128 2184 5140 2224
rect 5157 2184 5169 2204
rect 5177 2184 5189 2204
rect 5217 2184 5229 2224
rect 5237 2184 5249 2214
rect 5257 2184 5269 2224
rect 5277 2196 5289 2224
rect 5297 2184 5309 2224
rect 5351 2192 5363 2232
rect 5381 2192 5393 2224
rect 5411 2192 5423 2212
rect 5431 2192 5443 2212
rect 5457 2192 5469 2212
rect 5477 2192 5489 2212
rect 5507 2192 5519 2224
rect 5537 2192 5549 2232
rect 5577 2192 5589 2212
rect 5597 2192 5609 2212
rect 5627 2192 5639 2224
rect 5657 2192 5669 2232
rect 5734 2184 5746 2242
rect 5770 2184 5782 2244
rect 5834 2184 5846 2242
rect 5870 2184 5882 2244
rect 5911 2184 5923 2204
rect 5931 2184 5943 2204
rect 5992 2184 6004 2224
rect 6020 2184 6032 2224
rect 6048 2184 6060 2224
rect 6091 2192 6103 2232
rect 6121 2192 6133 2224
rect 6151 2192 6163 2212
rect 6171 2192 6183 2212
rect 6211 2192 6223 2232
rect 6241 2192 6253 2224
rect 6271 2192 6283 2212
rect 6291 2192 6303 2212
rect 6317 2184 6329 2204
rect 6337 2184 6349 2204
rect 6377 2184 6389 2224
rect 6397 2184 6409 2212
rect 6417 2184 6429 2224
rect 6437 2184 6449 2224
rect 6479 2184 6491 2224
rect 6509 2184 6521 2224
rect 6560 2184 6572 2224
rect 6588 2184 6600 2224
rect 6610 2184 6622 2204
rect 6657 2184 6669 2204
rect 6677 2184 6689 2204
rect 31 2136 43 2156
rect 51 2136 63 2156
rect 71 2136 83 2156
rect 119 2116 131 2156
rect 149 2116 161 2156
rect 214 2098 226 2156
rect 250 2096 262 2156
rect 314 2098 326 2156
rect 350 2096 362 2156
rect 399 2116 411 2156
rect 429 2116 441 2156
rect 458 2096 470 2156
rect 494 2098 506 2156
rect 571 2136 583 2156
rect 591 2136 603 2156
rect 611 2136 623 2156
rect 637 2116 649 2156
rect 657 2128 669 2156
rect 677 2116 689 2156
rect 697 2116 709 2156
rect 738 2096 750 2156
rect 774 2098 786 2156
rect 837 2136 849 2156
rect 857 2136 869 2156
rect 877 2136 889 2156
rect 939 2116 951 2156
rect 969 2116 981 2156
rect 997 2128 1009 2148
rect 1017 2128 1029 2148
rect 1047 2116 1059 2148
rect 1077 2108 1089 2148
rect 1121 2116 1133 2156
rect 1141 2136 1153 2156
rect 1173 2136 1185 2156
rect 1203 2136 1215 2156
rect 1225 2136 1237 2156
rect 1251 2136 1263 2156
rect 1279 2136 1291 2156
rect 1309 2136 1321 2156
rect 1331 2116 1343 2156
rect 1357 2136 1369 2156
rect 1377 2136 1389 2156
rect 1417 2116 1429 2156
rect 1437 2126 1449 2156
rect 1457 2116 1469 2156
rect 1477 2116 1489 2144
rect 1497 2116 1509 2156
rect 1551 2116 1563 2156
rect 1571 2116 1583 2156
rect 1591 2128 1603 2156
rect 1611 2116 1623 2156
rect 1651 2116 1663 2156
rect 1671 2116 1683 2156
rect 1691 2128 1703 2156
rect 1711 2116 1723 2156
rect 1751 2136 1763 2156
rect 1771 2136 1783 2156
rect 1791 2136 1803 2156
rect 1831 2116 1843 2156
rect 1851 2116 1863 2156
rect 1871 2128 1883 2156
rect 1891 2116 1903 2156
rect 1931 2108 1943 2148
rect 1961 2116 1973 2148
rect 1991 2128 2003 2148
rect 2011 2128 2023 2148
rect 2051 2108 2063 2148
rect 2081 2116 2093 2148
rect 2111 2128 2123 2148
rect 2131 2128 2143 2148
rect 2161 2116 2173 2156
rect 2181 2136 2193 2156
rect 2213 2136 2225 2156
rect 2243 2136 2255 2156
rect 2265 2136 2277 2156
rect 2291 2136 2303 2156
rect 2319 2136 2331 2156
rect 2349 2136 2361 2156
rect 2371 2116 2383 2156
rect 2411 2116 2423 2156
rect 2431 2116 2443 2156
rect 2451 2128 2463 2156
rect 2471 2116 2483 2156
rect 2497 2136 2509 2156
rect 2517 2136 2529 2156
rect 2537 2136 2549 2156
rect 2614 2098 2626 2156
rect 2650 2096 2662 2156
rect 2677 2128 2689 2148
rect 2697 2128 2709 2148
rect 2727 2116 2739 2148
rect 2757 2108 2769 2148
rect 2811 2108 2823 2148
rect 2841 2116 2853 2148
rect 2871 2128 2883 2148
rect 2891 2128 2903 2148
rect 2917 2136 2929 2156
rect 2937 2136 2949 2156
rect 2977 2116 2989 2156
rect 2997 2126 3009 2156
rect 3017 2116 3029 2156
rect 3037 2116 3049 2144
rect 3057 2116 3069 2156
rect 3118 2136 3130 2156
rect 3140 2116 3152 2156
rect 3168 2116 3180 2156
rect 3197 2136 3209 2156
rect 3217 2136 3229 2156
rect 3257 2116 3269 2156
rect 3277 2126 3289 2156
rect 3297 2116 3309 2156
rect 3317 2116 3329 2144
rect 3337 2116 3349 2156
rect 3377 2136 3389 2156
rect 3397 2136 3409 2156
rect 3417 2136 3429 2156
rect 3461 2116 3473 2156
rect 3481 2136 3493 2156
rect 3513 2136 3525 2156
rect 3543 2136 3555 2156
rect 3565 2136 3577 2156
rect 3591 2136 3603 2156
rect 3619 2136 3631 2156
rect 3649 2136 3661 2156
rect 3671 2116 3683 2156
rect 3711 2136 3723 2156
rect 3731 2136 3743 2156
rect 3751 2136 3763 2156
rect 3791 2116 3803 2156
rect 3811 2116 3823 2144
rect 3831 2116 3843 2156
rect 3851 2126 3863 2156
rect 3871 2116 3883 2156
rect 3911 2136 3923 2156
rect 3931 2136 3943 2156
rect 3957 2116 3969 2156
rect 3977 2128 3989 2156
rect 3997 2116 4009 2156
rect 4017 2116 4029 2156
rect 4059 2116 4071 2156
rect 4089 2116 4101 2156
rect 4151 2136 4163 2156
rect 4171 2136 4183 2156
rect 4191 2136 4203 2156
rect 4221 2116 4233 2156
rect 4241 2136 4253 2156
rect 4273 2136 4285 2156
rect 4303 2136 4315 2156
rect 4325 2136 4337 2156
rect 4351 2136 4363 2156
rect 4379 2136 4391 2156
rect 4409 2136 4421 2156
rect 4431 2116 4443 2156
rect 4457 2136 4469 2156
rect 4477 2136 4489 2156
rect 4517 2116 4529 2156
rect 4537 2126 4549 2156
rect 4557 2116 4569 2156
rect 4577 2116 4589 2144
rect 4597 2116 4609 2156
rect 4637 2136 4649 2156
rect 4657 2136 4669 2156
rect 4677 2136 4689 2156
rect 4731 2116 4743 2156
rect 4751 2116 4763 2156
rect 4771 2128 4783 2156
rect 4791 2116 4803 2156
rect 4831 2136 4843 2156
rect 4851 2136 4863 2156
rect 4871 2136 4883 2156
rect 4897 2116 4909 2156
rect 4917 2126 4929 2156
rect 4937 2116 4949 2156
rect 4957 2116 4969 2144
rect 4977 2116 4989 2156
rect 5039 2116 5051 2156
rect 5069 2116 5081 2156
rect 5111 2136 5123 2156
rect 5131 2136 5143 2156
rect 5151 2136 5163 2156
rect 5177 2136 5189 2156
rect 5197 2136 5209 2156
rect 5217 2136 5229 2156
rect 5237 2116 5249 2156
rect 5291 2116 5303 2156
rect 5311 2116 5323 2144
rect 5331 2116 5343 2156
rect 5351 2126 5363 2156
rect 5371 2116 5383 2156
rect 5397 2116 5409 2156
rect 5417 2126 5429 2156
rect 5437 2116 5449 2156
rect 5457 2116 5469 2144
rect 5477 2116 5489 2156
rect 5531 2136 5543 2156
rect 5551 2136 5563 2156
rect 5571 2136 5583 2156
rect 5611 2116 5623 2156
rect 5631 2116 5643 2144
rect 5651 2116 5663 2156
rect 5671 2126 5683 2156
rect 5691 2116 5703 2156
rect 5731 2136 5743 2156
rect 5751 2136 5763 2156
rect 5779 2116 5791 2156
rect 5809 2116 5821 2156
rect 5857 2116 5869 2156
rect 5879 2136 5891 2156
rect 5909 2136 5921 2156
rect 5937 2136 5949 2156
rect 5963 2136 5975 2156
rect 5985 2136 5997 2156
rect 6015 2136 6027 2156
rect 6047 2136 6059 2156
rect 6067 2116 6079 2156
rect 6101 2116 6113 2156
rect 6121 2136 6133 2156
rect 6153 2136 6165 2156
rect 6183 2136 6195 2156
rect 6205 2136 6217 2156
rect 6231 2136 6243 2156
rect 6259 2136 6271 2156
rect 6289 2136 6301 2156
rect 6311 2116 6323 2156
rect 6337 2128 6349 2148
rect 6357 2128 6369 2148
rect 6387 2116 6399 2148
rect 6417 2108 6429 2148
rect 6460 2116 6472 2156
rect 6488 2116 6500 2156
rect 6510 2136 6522 2156
rect 6557 2116 6569 2156
rect 6577 2128 6589 2156
rect 6597 2116 6609 2156
rect 6617 2116 6629 2156
rect 31 1704 43 1724
rect 51 1704 63 1724
rect 77 1704 89 1744
rect 99 1704 111 1724
rect 129 1704 141 1724
rect 157 1704 169 1724
rect 183 1704 195 1724
rect 205 1704 217 1724
rect 235 1704 247 1724
rect 267 1704 279 1724
rect 287 1704 299 1744
rect 317 1704 329 1724
rect 337 1704 349 1724
rect 357 1704 369 1724
rect 411 1704 423 1724
rect 431 1704 443 1724
rect 451 1704 463 1724
rect 491 1704 503 1724
rect 511 1704 523 1724
rect 551 1704 563 1744
rect 571 1704 583 1744
rect 591 1704 603 1732
rect 611 1704 623 1744
rect 637 1704 649 1744
rect 659 1704 671 1724
rect 689 1704 701 1724
rect 717 1704 729 1724
rect 743 1704 755 1724
rect 765 1704 777 1724
rect 795 1704 807 1724
rect 827 1704 839 1724
rect 847 1704 859 1744
rect 914 1704 926 1762
rect 950 1704 962 1764
rect 977 1704 989 1744
rect 1007 1704 1019 1744
rect 1027 1704 1039 1744
rect 1077 1704 1089 1724
rect 1097 1704 1109 1724
rect 1137 1704 1149 1744
rect 1157 1704 1169 1732
rect 1177 1704 1189 1744
rect 1197 1704 1209 1744
rect 1259 1704 1271 1744
rect 1289 1704 1301 1744
rect 1354 1704 1366 1762
rect 1390 1704 1402 1764
rect 1417 1704 1429 1724
rect 1437 1704 1449 1724
rect 1481 1704 1493 1744
rect 1501 1704 1513 1724
rect 1533 1704 1545 1724
rect 1563 1704 1575 1724
rect 1585 1704 1597 1724
rect 1611 1704 1623 1724
rect 1639 1704 1651 1724
rect 1669 1704 1681 1724
rect 1691 1704 1703 1744
rect 1717 1704 1729 1724
rect 1737 1704 1749 1724
rect 1777 1704 1789 1744
rect 1797 1704 1809 1734
rect 1817 1704 1829 1744
rect 1837 1716 1849 1744
rect 1857 1704 1869 1744
rect 1897 1704 1909 1724
rect 1917 1704 1929 1724
rect 1937 1704 1949 1724
rect 1977 1704 1989 1744
rect 1997 1704 2009 1732
rect 2017 1704 2029 1744
rect 2037 1704 2049 1744
rect 2077 1704 2089 1744
rect 2099 1704 2111 1724
rect 2129 1704 2141 1724
rect 2157 1704 2169 1724
rect 2183 1704 2195 1724
rect 2205 1704 2217 1724
rect 2235 1704 2247 1724
rect 2267 1704 2279 1724
rect 2287 1704 2299 1744
rect 2331 1704 2343 1744
rect 2351 1716 2363 1744
rect 2371 1704 2383 1744
rect 2391 1704 2403 1734
rect 2411 1704 2423 1744
rect 2437 1704 2449 1724
rect 2457 1704 2469 1724
rect 2497 1704 2509 1724
rect 2517 1704 2529 1724
rect 2537 1704 2549 1724
rect 2577 1704 2589 1744
rect 2599 1704 2611 1724
rect 2629 1704 2641 1724
rect 2657 1704 2669 1724
rect 2683 1704 2695 1724
rect 2705 1704 2717 1724
rect 2735 1704 2747 1724
rect 2767 1704 2779 1724
rect 2787 1704 2799 1744
rect 2818 1704 2830 1764
rect 2854 1704 2866 1762
rect 2931 1704 2943 1744
rect 2951 1704 2963 1744
rect 2971 1704 2983 1732
rect 2991 1704 3003 1744
rect 3017 1704 3029 1724
rect 3037 1704 3049 1724
rect 3057 1704 3069 1724
rect 3118 1704 3130 1724
rect 3140 1704 3152 1744
rect 3168 1704 3180 1744
rect 3218 1704 3230 1724
rect 3240 1704 3252 1744
rect 3268 1704 3280 1744
rect 3309 1704 3321 1744
rect 3329 1704 3341 1744
rect 3351 1704 3363 1724
rect 3399 1704 3411 1744
rect 3429 1704 3441 1744
rect 3457 1704 3469 1724
rect 3477 1704 3489 1724
rect 3497 1704 3509 1724
rect 3539 1704 3551 1744
rect 3569 1704 3581 1744
rect 3617 1704 3629 1744
rect 3637 1704 3649 1732
rect 3657 1704 3669 1744
rect 3677 1704 3689 1744
rect 3739 1704 3751 1744
rect 3769 1704 3781 1744
rect 3811 1704 3823 1724
rect 3831 1704 3843 1724
rect 3859 1704 3871 1744
rect 3889 1704 3901 1744
rect 3937 1704 3949 1724
rect 3957 1704 3969 1724
rect 3977 1704 3989 1724
rect 4017 1704 4029 1744
rect 4037 1704 4049 1734
rect 4057 1704 4069 1744
rect 4077 1716 4089 1744
rect 4097 1704 4109 1744
rect 4151 1704 4163 1724
rect 4171 1704 4183 1724
rect 4191 1704 4203 1724
rect 4217 1704 4229 1744
rect 4237 1704 4249 1732
rect 4257 1704 4269 1744
rect 4277 1704 4289 1744
rect 4317 1704 4329 1744
rect 4337 1704 4349 1744
rect 4357 1704 4369 1744
rect 4397 1704 4409 1744
rect 4417 1704 4429 1732
rect 4437 1704 4449 1744
rect 4457 1704 4469 1744
rect 4511 1704 4523 1724
rect 4531 1704 4543 1724
rect 4551 1704 4563 1724
rect 4591 1704 4603 1744
rect 4611 1716 4623 1744
rect 4631 1704 4643 1744
rect 4651 1704 4663 1734
rect 4671 1704 4683 1744
rect 4711 1704 4723 1724
rect 4731 1704 4743 1724
rect 4757 1704 4769 1744
rect 4779 1704 4791 1724
rect 4809 1704 4821 1724
rect 4837 1704 4849 1724
rect 4863 1704 4875 1724
rect 4885 1704 4897 1724
rect 4915 1704 4927 1724
rect 4947 1704 4959 1724
rect 4967 1704 4979 1744
rect 5000 1704 5012 1744
rect 5028 1704 5040 1744
rect 5050 1704 5062 1724
rect 5097 1704 5109 1724
rect 5117 1704 5129 1724
rect 5137 1704 5149 1724
rect 5177 1704 5189 1744
rect 5197 1704 5209 1732
rect 5217 1704 5229 1744
rect 5237 1704 5249 1744
rect 5278 1704 5290 1764
rect 5314 1704 5326 1762
rect 5377 1704 5389 1724
rect 5399 1704 5411 1744
rect 5419 1704 5431 1744
rect 5471 1704 5483 1724
rect 5491 1704 5503 1724
rect 5531 1704 5543 1744
rect 5551 1704 5563 1744
rect 5591 1704 5603 1744
rect 5611 1704 5623 1744
rect 5631 1704 5643 1732
rect 5651 1704 5663 1744
rect 5679 1704 5691 1744
rect 5709 1704 5721 1744
rect 5792 1704 5804 1744
rect 5820 1704 5832 1744
rect 5848 1704 5860 1744
rect 5877 1704 5889 1724
rect 5899 1704 5911 1744
rect 5919 1704 5931 1744
rect 5971 1704 5983 1744
rect 5991 1704 6003 1744
rect 6011 1704 6023 1732
rect 6031 1704 6043 1744
rect 6071 1704 6083 1744
rect 6091 1716 6103 1744
rect 6111 1704 6123 1744
rect 6131 1704 6143 1734
rect 6151 1704 6163 1744
rect 6177 1712 6189 1732
rect 6197 1712 6209 1732
rect 6227 1712 6239 1744
rect 6257 1712 6269 1752
rect 6297 1712 6309 1732
rect 6317 1712 6329 1732
rect 6347 1712 6359 1744
rect 6377 1712 6389 1752
rect 6417 1704 6429 1724
rect 6437 1704 6449 1724
rect 6477 1704 6489 1744
rect 6497 1704 6509 1732
rect 6517 1704 6529 1744
rect 6537 1704 6549 1744
rect 6599 1704 6611 1744
rect 6629 1704 6641 1744
rect 31 1656 43 1676
rect 51 1656 63 1676
rect 71 1656 83 1676
rect 111 1636 123 1676
rect 131 1636 143 1676
rect 151 1636 163 1676
rect 171 1636 183 1676
rect 191 1636 203 1676
rect 211 1636 223 1676
rect 231 1636 243 1676
rect 251 1636 263 1676
rect 271 1636 283 1676
rect 301 1636 313 1676
rect 321 1656 333 1676
rect 353 1656 365 1676
rect 383 1656 395 1676
rect 405 1656 417 1676
rect 431 1656 443 1676
rect 459 1656 471 1676
rect 489 1656 501 1676
rect 511 1636 523 1676
rect 551 1656 563 1676
rect 571 1656 583 1676
rect 598 1616 610 1676
rect 634 1618 646 1676
rect 700 1636 712 1676
rect 728 1636 740 1676
rect 750 1656 762 1676
rect 801 1636 813 1676
rect 821 1656 833 1676
rect 853 1656 865 1676
rect 883 1656 895 1676
rect 905 1656 917 1676
rect 931 1656 943 1676
rect 959 1656 971 1676
rect 989 1656 1001 1676
rect 1011 1636 1023 1676
rect 1051 1656 1063 1676
rect 1071 1656 1083 1676
rect 1097 1636 1109 1676
rect 1117 1646 1129 1676
rect 1137 1636 1149 1676
rect 1157 1636 1169 1664
rect 1177 1636 1189 1676
rect 1231 1636 1243 1676
rect 1251 1636 1263 1676
rect 1271 1648 1283 1676
rect 1291 1636 1303 1676
rect 1331 1656 1343 1676
rect 1351 1656 1363 1676
rect 1371 1656 1383 1676
rect 1411 1628 1423 1668
rect 1441 1636 1453 1668
rect 1471 1648 1483 1668
rect 1491 1648 1503 1668
rect 1531 1628 1543 1668
rect 1561 1636 1573 1668
rect 1591 1648 1603 1668
rect 1611 1648 1623 1668
rect 1651 1628 1663 1668
rect 1681 1636 1693 1668
rect 1711 1648 1723 1668
rect 1731 1648 1743 1668
rect 1757 1636 1769 1676
rect 1779 1656 1791 1676
rect 1809 1656 1821 1676
rect 1837 1656 1849 1676
rect 1863 1656 1875 1676
rect 1885 1656 1897 1676
rect 1915 1656 1927 1676
rect 1947 1656 1959 1676
rect 1967 1636 1979 1676
rect 1997 1648 2009 1668
rect 2017 1648 2029 1668
rect 2047 1636 2059 1668
rect 2077 1628 2089 1668
rect 2117 1656 2129 1676
rect 2137 1656 2149 1676
rect 2177 1636 2189 1676
rect 2197 1646 2209 1676
rect 2217 1636 2229 1676
rect 2237 1636 2249 1664
rect 2257 1636 2269 1676
rect 2297 1656 2309 1676
rect 2317 1656 2329 1676
rect 2337 1656 2349 1676
rect 2391 1636 2403 1676
rect 2411 1636 2423 1676
rect 2431 1648 2443 1676
rect 2451 1636 2463 1676
rect 2489 1636 2501 1676
rect 2509 1636 2521 1676
rect 2531 1656 2543 1676
rect 2557 1656 2569 1676
rect 2577 1656 2589 1676
rect 2597 1656 2609 1676
rect 2659 1636 2671 1676
rect 2689 1636 2701 1676
rect 2719 1636 2731 1676
rect 2749 1636 2761 1676
rect 2811 1628 2823 1668
rect 2841 1636 2853 1668
rect 2871 1648 2883 1668
rect 2891 1648 2903 1668
rect 2954 1618 2966 1676
rect 2990 1616 3002 1676
rect 3031 1636 3043 1676
rect 3051 1636 3063 1676
rect 3081 1636 3093 1676
rect 3101 1656 3113 1676
rect 3133 1656 3145 1676
rect 3163 1656 3175 1676
rect 3185 1656 3197 1676
rect 3211 1656 3223 1676
rect 3239 1656 3251 1676
rect 3269 1656 3281 1676
rect 3291 1636 3303 1676
rect 3339 1636 3351 1676
rect 3369 1636 3381 1676
rect 3411 1636 3423 1676
rect 3431 1636 3443 1676
rect 3451 1648 3463 1676
rect 3471 1636 3483 1676
rect 3500 1636 3512 1676
rect 3528 1636 3540 1676
rect 3556 1636 3568 1676
rect 3631 1636 3643 1676
rect 3651 1636 3663 1676
rect 3671 1648 3683 1676
rect 3691 1636 3703 1676
rect 3731 1656 3743 1676
rect 3751 1656 3763 1676
rect 3791 1656 3803 1676
rect 3811 1656 3823 1676
rect 3831 1656 3843 1676
rect 3871 1636 3883 1676
rect 3891 1636 3903 1664
rect 3911 1636 3923 1676
rect 3931 1646 3943 1676
rect 3951 1636 3963 1676
rect 3991 1656 4003 1676
rect 4011 1656 4023 1676
rect 4041 1636 4053 1676
rect 4061 1656 4073 1676
rect 4093 1656 4105 1676
rect 4123 1656 4135 1676
rect 4145 1656 4157 1676
rect 4171 1656 4183 1676
rect 4199 1656 4211 1676
rect 4229 1656 4241 1676
rect 4251 1636 4263 1676
rect 4291 1628 4303 1668
rect 4321 1636 4333 1668
rect 4351 1648 4363 1668
rect 4371 1648 4383 1668
rect 4411 1628 4423 1668
rect 4441 1636 4453 1668
rect 4471 1648 4483 1668
rect 4491 1648 4503 1668
rect 4517 1648 4529 1668
rect 4537 1648 4549 1668
rect 4567 1636 4579 1668
rect 4597 1628 4609 1668
rect 4637 1648 4649 1668
rect 4657 1648 4669 1668
rect 4687 1636 4699 1668
rect 4717 1628 4729 1668
rect 4757 1648 4769 1668
rect 4777 1648 4789 1668
rect 4807 1636 4819 1668
rect 4837 1628 4849 1668
rect 4877 1648 4889 1668
rect 4897 1648 4909 1668
rect 4927 1636 4939 1668
rect 4957 1628 4969 1668
rect 4997 1636 5009 1676
rect 5019 1656 5031 1676
rect 5049 1656 5061 1676
rect 5077 1656 5089 1676
rect 5103 1656 5115 1676
rect 5125 1656 5137 1676
rect 5155 1656 5167 1676
rect 5187 1656 5199 1676
rect 5207 1636 5219 1676
rect 5237 1636 5249 1676
rect 5259 1656 5271 1676
rect 5289 1656 5301 1676
rect 5317 1656 5329 1676
rect 5343 1656 5355 1676
rect 5365 1656 5377 1676
rect 5395 1656 5407 1676
rect 5427 1656 5439 1676
rect 5447 1636 5459 1676
rect 5480 1636 5492 1676
rect 5508 1636 5520 1676
rect 5536 1636 5548 1676
rect 5597 1648 5609 1668
rect 5617 1648 5629 1668
rect 5647 1636 5659 1668
rect 5677 1628 5689 1668
rect 5731 1636 5743 1676
rect 5751 1636 5763 1676
rect 5771 1648 5783 1676
rect 5791 1636 5803 1676
rect 5831 1656 5843 1676
rect 5851 1656 5863 1676
rect 5871 1656 5883 1676
rect 5919 1636 5931 1676
rect 5949 1636 5961 1676
rect 5991 1636 6003 1676
rect 6011 1636 6023 1676
rect 6031 1648 6043 1676
rect 6051 1636 6063 1676
rect 6091 1656 6103 1676
rect 6111 1656 6123 1676
rect 6131 1656 6143 1676
rect 6171 1636 6183 1676
rect 6191 1636 6203 1664
rect 6211 1636 6223 1676
rect 6231 1646 6243 1676
rect 6251 1636 6263 1676
rect 6291 1628 6303 1668
rect 6321 1636 6333 1668
rect 6351 1648 6363 1668
rect 6371 1648 6383 1668
rect 6397 1656 6409 1676
rect 6417 1656 6429 1676
rect 6457 1636 6469 1676
rect 6479 1656 6491 1676
rect 6509 1656 6521 1676
rect 6537 1656 6549 1676
rect 6563 1656 6575 1676
rect 6585 1656 6597 1676
rect 6615 1656 6627 1676
rect 6647 1656 6659 1676
rect 6667 1636 6679 1676
rect 17 1224 29 1264
rect 47 1224 59 1264
rect 67 1224 79 1264
rect 117 1224 129 1244
rect 137 1224 149 1244
rect 157 1224 169 1244
rect 211 1224 223 1264
rect 231 1224 243 1264
rect 251 1224 263 1252
rect 271 1224 283 1264
rect 311 1224 323 1244
rect 331 1224 343 1244
rect 351 1224 363 1244
rect 377 1224 389 1244
rect 397 1224 409 1244
rect 437 1224 449 1244
rect 457 1224 469 1244
rect 519 1224 531 1264
rect 549 1224 561 1264
rect 580 1224 592 1264
rect 608 1224 620 1264
rect 630 1224 642 1244
rect 681 1224 693 1264
rect 701 1224 713 1244
rect 733 1224 745 1244
rect 763 1224 775 1244
rect 785 1224 797 1244
rect 811 1224 823 1244
rect 839 1224 851 1244
rect 869 1224 881 1244
rect 891 1224 903 1264
rect 939 1224 951 1264
rect 969 1224 981 1264
rect 998 1224 1010 1284
rect 1034 1224 1046 1282
rect 1097 1224 1109 1244
rect 1117 1224 1129 1244
rect 1137 1224 1149 1244
rect 1181 1224 1193 1264
rect 1201 1224 1213 1244
rect 1233 1224 1245 1244
rect 1263 1224 1275 1244
rect 1285 1224 1297 1244
rect 1311 1224 1323 1244
rect 1339 1224 1351 1244
rect 1369 1224 1381 1244
rect 1391 1224 1403 1264
rect 1431 1224 1443 1264
rect 1451 1224 1463 1264
rect 1471 1224 1483 1264
rect 1491 1224 1503 1264
rect 1511 1224 1523 1264
rect 1531 1224 1543 1264
rect 1551 1224 1563 1264
rect 1571 1224 1583 1264
rect 1591 1224 1603 1264
rect 1631 1232 1643 1272
rect 1661 1232 1673 1264
rect 1691 1232 1703 1252
rect 1711 1232 1723 1252
rect 1751 1224 1763 1244
rect 1771 1224 1783 1244
rect 1791 1224 1803 1244
rect 1831 1224 1843 1264
rect 1851 1236 1863 1264
rect 1871 1224 1883 1264
rect 1891 1224 1903 1254
rect 1911 1224 1923 1264
rect 1951 1224 1963 1264
rect 1971 1224 1983 1264
rect 1991 1224 2003 1252
rect 2011 1224 2023 1264
rect 2037 1224 2049 1244
rect 2057 1224 2069 1244
rect 2097 1224 2109 1264
rect 2117 1224 2129 1252
rect 2137 1224 2149 1264
rect 2157 1224 2169 1264
rect 2199 1224 2211 1264
rect 2229 1224 2241 1264
rect 2277 1232 2289 1252
rect 2297 1232 2309 1252
rect 2327 1232 2339 1264
rect 2357 1232 2369 1272
rect 2411 1232 2423 1272
rect 2441 1232 2453 1264
rect 2471 1232 2483 1252
rect 2491 1232 2503 1252
rect 2552 1224 2564 1264
rect 2580 1224 2592 1264
rect 2608 1224 2620 1264
rect 2640 1224 2652 1264
rect 2668 1224 2680 1264
rect 2696 1224 2708 1264
rect 2792 1224 2804 1264
rect 2820 1224 2832 1264
rect 2848 1224 2860 1264
rect 2877 1224 2889 1244
rect 2899 1224 2911 1264
rect 2919 1224 2931 1264
rect 2992 1224 3004 1264
rect 3020 1224 3032 1264
rect 3048 1224 3060 1264
rect 3091 1224 3103 1244
rect 3111 1224 3123 1244
rect 3151 1232 3163 1272
rect 3181 1232 3193 1264
rect 3211 1232 3223 1252
rect 3231 1232 3243 1252
rect 3261 1224 3273 1264
rect 3281 1224 3293 1244
rect 3313 1224 3325 1244
rect 3343 1224 3355 1244
rect 3365 1224 3377 1244
rect 3391 1224 3403 1244
rect 3419 1224 3431 1244
rect 3449 1224 3461 1244
rect 3471 1224 3483 1264
rect 3511 1224 3523 1244
rect 3531 1224 3543 1244
rect 3551 1224 3563 1244
rect 3591 1224 3603 1264
rect 3611 1236 3623 1264
rect 3631 1224 3643 1264
rect 3651 1224 3663 1254
rect 3671 1224 3683 1264
rect 3711 1224 3723 1264
rect 3731 1224 3743 1264
rect 3751 1224 3763 1252
rect 3771 1224 3783 1264
rect 3811 1224 3823 1244
rect 3831 1224 3843 1244
rect 3857 1224 3869 1264
rect 3879 1224 3891 1244
rect 3909 1224 3921 1244
rect 3937 1224 3949 1244
rect 3963 1224 3975 1244
rect 3985 1224 3997 1244
rect 4015 1224 4027 1244
rect 4047 1224 4059 1244
rect 4067 1224 4079 1264
rect 4097 1224 4109 1264
rect 4119 1224 4131 1244
rect 4149 1224 4161 1244
rect 4177 1224 4189 1244
rect 4203 1224 4215 1244
rect 4225 1224 4237 1244
rect 4255 1224 4267 1244
rect 4287 1224 4299 1244
rect 4307 1224 4319 1264
rect 4351 1224 4363 1244
rect 4371 1224 4383 1244
rect 4400 1224 4412 1264
rect 4428 1224 4440 1264
rect 4456 1224 4468 1264
rect 4517 1232 4529 1252
rect 4537 1232 4549 1252
rect 4567 1232 4579 1264
rect 4597 1232 4609 1272
rect 4672 1224 4684 1264
rect 4700 1224 4712 1264
rect 4728 1224 4740 1264
rect 4769 1224 4781 1264
rect 4789 1224 4801 1264
rect 4811 1224 4823 1244
rect 4859 1224 4871 1264
rect 4889 1224 4901 1264
rect 4939 1224 4951 1264
rect 4969 1224 4981 1264
rect 5011 1224 5023 1264
rect 5031 1236 5043 1264
rect 5051 1224 5063 1264
rect 5071 1224 5083 1254
rect 5091 1224 5103 1264
rect 5131 1224 5143 1264
rect 5151 1236 5163 1264
rect 5171 1224 5183 1264
rect 5191 1224 5203 1254
rect 5211 1224 5223 1264
rect 5237 1224 5249 1264
rect 5257 1224 5269 1264
rect 5319 1224 5331 1264
rect 5349 1224 5361 1264
rect 5377 1224 5389 1264
rect 5397 1224 5409 1254
rect 5417 1224 5429 1264
rect 5437 1236 5449 1264
rect 5457 1224 5469 1264
rect 5518 1224 5530 1244
rect 5540 1224 5552 1264
rect 5568 1224 5580 1264
rect 5597 1224 5609 1264
rect 5617 1224 5629 1264
rect 5657 1232 5669 1252
rect 5677 1232 5689 1252
rect 5707 1232 5719 1264
rect 5737 1232 5749 1272
rect 5799 1224 5811 1264
rect 5829 1224 5841 1264
rect 5871 1224 5883 1264
rect 5891 1224 5903 1264
rect 5911 1224 5923 1252
rect 5931 1224 5943 1264
rect 5971 1224 5983 1244
rect 5991 1224 6003 1244
rect 6017 1224 6029 1264
rect 6037 1224 6049 1252
rect 6057 1224 6069 1264
rect 6077 1224 6089 1264
rect 6117 1224 6129 1264
rect 6137 1224 6149 1254
rect 6157 1224 6169 1264
rect 6177 1236 6189 1264
rect 6197 1224 6209 1264
rect 6237 1224 6249 1264
rect 6259 1224 6271 1244
rect 6289 1224 6301 1244
rect 6317 1224 6329 1244
rect 6343 1224 6355 1244
rect 6365 1224 6377 1244
rect 6395 1224 6407 1244
rect 6427 1224 6439 1244
rect 6447 1224 6459 1264
rect 6477 1224 6489 1264
rect 6499 1224 6511 1244
rect 6529 1224 6541 1244
rect 6557 1224 6569 1244
rect 6583 1224 6595 1244
rect 6605 1224 6617 1244
rect 6635 1224 6647 1244
rect 6667 1224 6679 1244
rect 6687 1224 6699 1264
rect 17 1156 29 1196
rect 39 1176 51 1196
rect 69 1176 81 1196
rect 97 1176 109 1196
rect 123 1176 135 1196
rect 145 1176 157 1196
rect 175 1176 187 1196
rect 207 1176 219 1196
rect 227 1156 239 1196
rect 271 1176 283 1196
rect 291 1176 303 1196
rect 317 1156 329 1196
rect 339 1176 351 1196
rect 369 1176 381 1196
rect 397 1176 409 1196
rect 423 1176 435 1196
rect 445 1176 457 1196
rect 475 1176 487 1196
rect 507 1176 519 1196
rect 527 1156 539 1196
rect 557 1176 569 1196
rect 577 1176 589 1196
rect 618 1136 630 1196
rect 654 1138 666 1196
rect 717 1176 729 1196
rect 737 1176 749 1196
rect 757 1176 769 1196
rect 798 1136 810 1196
rect 834 1138 846 1196
rect 899 1156 911 1196
rect 929 1156 941 1196
rect 977 1176 989 1196
rect 997 1176 1009 1196
rect 1041 1156 1053 1196
rect 1061 1176 1073 1196
rect 1093 1176 1105 1196
rect 1123 1176 1135 1196
rect 1145 1176 1157 1196
rect 1171 1176 1183 1196
rect 1199 1176 1211 1196
rect 1229 1176 1241 1196
rect 1251 1156 1263 1196
rect 1277 1156 1289 1196
rect 1297 1156 1309 1196
rect 1317 1156 1329 1196
rect 1337 1156 1349 1196
rect 1357 1156 1369 1196
rect 1377 1156 1389 1196
rect 1397 1156 1409 1196
rect 1417 1156 1429 1196
rect 1437 1156 1449 1196
rect 1481 1156 1493 1196
rect 1501 1176 1513 1196
rect 1533 1176 1545 1196
rect 1563 1176 1575 1196
rect 1585 1176 1597 1196
rect 1611 1176 1623 1196
rect 1639 1176 1651 1196
rect 1669 1176 1681 1196
rect 1691 1156 1703 1196
rect 1731 1176 1743 1196
rect 1751 1176 1763 1196
rect 1771 1176 1783 1196
rect 1811 1156 1823 1196
rect 1831 1156 1843 1184
rect 1851 1156 1863 1196
rect 1871 1166 1883 1196
rect 1891 1156 1903 1196
rect 1931 1156 1943 1196
rect 1951 1156 1963 1196
rect 1971 1168 1983 1196
rect 1991 1156 2003 1196
rect 2031 1156 2043 1196
rect 2051 1156 2063 1196
rect 2071 1168 2083 1196
rect 2091 1156 2103 1196
rect 2131 1176 2143 1196
rect 2151 1176 2163 1196
rect 2171 1176 2183 1196
rect 2211 1156 2223 1196
rect 2231 1156 2243 1184
rect 2251 1156 2263 1196
rect 2271 1166 2283 1196
rect 2291 1156 2303 1196
rect 2321 1156 2333 1196
rect 2341 1176 2353 1196
rect 2373 1176 2385 1196
rect 2403 1176 2415 1196
rect 2425 1176 2437 1196
rect 2451 1176 2463 1196
rect 2479 1176 2491 1196
rect 2509 1176 2521 1196
rect 2531 1156 2543 1196
rect 2571 1176 2583 1196
rect 2591 1176 2603 1196
rect 2617 1156 2629 1196
rect 2637 1168 2649 1196
rect 2657 1156 2669 1196
rect 2677 1156 2689 1196
rect 2729 1156 2741 1196
rect 2749 1156 2761 1196
rect 2771 1176 2783 1196
rect 2797 1176 2809 1196
rect 2817 1176 2829 1196
rect 2892 1156 2904 1196
rect 2920 1156 2932 1196
rect 2948 1156 2960 1196
rect 2981 1156 2993 1196
rect 3001 1176 3013 1196
rect 3033 1176 3045 1196
rect 3063 1176 3075 1196
rect 3085 1176 3097 1196
rect 3111 1176 3123 1196
rect 3139 1176 3151 1196
rect 3169 1176 3181 1196
rect 3191 1156 3203 1196
rect 3219 1156 3231 1196
rect 3249 1156 3261 1196
rect 3311 1148 3323 1188
rect 3341 1156 3353 1188
rect 3371 1168 3383 1188
rect 3391 1168 3403 1188
rect 3417 1168 3429 1188
rect 3437 1168 3449 1188
rect 3467 1156 3479 1188
rect 3497 1148 3509 1188
rect 3549 1156 3561 1196
rect 3569 1156 3581 1196
rect 3591 1176 3603 1196
rect 3621 1156 3633 1196
rect 3641 1176 3653 1196
rect 3673 1176 3685 1196
rect 3703 1176 3715 1196
rect 3725 1176 3737 1196
rect 3751 1176 3763 1196
rect 3779 1176 3791 1196
rect 3809 1176 3821 1196
rect 3831 1156 3843 1196
rect 3857 1168 3869 1188
rect 3877 1168 3889 1188
rect 3907 1156 3919 1188
rect 3937 1148 3949 1188
rect 3991 1148 4003 1188
rect 4021 1156 4033 1188
rect 4051 1168 4063 1188
rect 4071 1168 4083 1188
rect 4097 1176 4109 1196
rect 4117 1176 4129 1196
rect 4157 1156 4169 1196
rect 4177 1166 4189 1196
rect 4197 1156 4209 1196
rect 4217 1156 4229 1184
rect 4237 1156 4249 1196
rect 4277 1176 4289 1196
rect 4297 1176 4309 1196
rect 4317 1176 4329 1196
rect 4371 1156 4383 1196
rect 4391 1156 4403 1196
rect 4411 1168 4423 1196
rect 4431 1156 4443 1196
rect 4478 1176 4490 1196
rect 4500 1156 4512 1196
rect 4528 1156 4540 1196
rect 4561 1156 4573 1196
rect 4581 1176 4593 1196
rect 4613 1176 4625 1196
rect 4643 1176 4655 1196
rect 4665 1176 4677 1196
rect 4691 1176 4703 1196
rect 4719 1176 4731 1196
rect 4749 1176 4761 1196
rect 4771 1156 4783 1196
rect 4797 1156 4809 1196
rect 4817 1166 4829 1196
rect 4837 1156 4849 1196
rect 4857 1156 4869 1184
rect 4877 1156 4889 1196
rect 4931 1176 4943 1196
rect 4951 1176 4963 1196
rect 4971 1176 4983 1196
rect 5011 1156 5023 1196
rect 5031 1156 5043 1196
rect 5051 1168 5063 1196
rect 5071 1156 5083 1196
rect 5111 1176 5123 1196
rect 5131 1176 5143 1196
rect 5151 1176 5163 1196
rect 5177 1176 5189 1196
rect 5197 1176 5209 1196
rect 5217 1176 5229 1196
rect 5257 1176 5269 1196
rect 5277 1176 5289 1196
rect 5297 1176 5309 1196
rect 5349 1156 5361 1196
rect 5369 1156 5381 1196
rect 5391 1176 5403 1196
rect 5417 1176 5429 1196
rect 5437 1176 5449 1196
rect 5457 1176 5469 1196
rect 5497 1176 5509 1196
rect 5517 1176 5529 1196
rect 5537 1176 5549 1196
rect 5580 1156 5592 1196
rect 5608 1156 5620 1196
rect 5630 1176 5642 1196
rect 5677 1176 5689 1196
rect 5697 1176 5709 1196
rect 5717 1176 5729 1196
rect 5737 1156 5749 1196
rect 5791 1176 5803 1196
rect 5811 1176 5823 1196
rect 5831 1176 5843 1196
rect 5857 1156 5869 1196
rect 5877 1168 5889 1196
rect 5897 1156 5909 1196
rect 5917 1156 5929 1196
rect 5994 1138 6006 1196
rect 6030 1136 6042 1196
rect 6057 1156 6069 1196
rect 6077 1168 6089 1196
rect 6097 1156 6109 1196
rect 6117 1156 6129 1196
rect 6171 1176 6183 1196
rect 6191 1176 6203 1196
rect 6211 1176 6223 1196
rect 6237 1176 6249 1196
rect 6257 1176 6269 1196
rect 6277 1176 6289 1196
rect 6317 1156 6329 1196
rect 6339 1176 6351 1196
rect 6369 1176 6381 1196
rect 6397 1176 6409 1196
rect 6423 1176 6435 1196
rect 6445 1176 6457 1196
rect 6475 1176 6487 1196
rect 6507 1176 6519 1196
rect 6527 1156 6539 1196
rect 6557 1156 6569 1196
rect 6577 1166 6589 1196
rect 6597 1156 6609 1196
rect 6617 1156 6629 1184
rect 6637 1156 6649 1196
rect 17 744 29 764
rect 37 744 49 764
rect 57 744 69 764
rect 77 744 89 784
rect 139 744 151 784
rect 169 744 181 784
rect 197 744 209 784
rect 219 744 231 764
rect 249 744 261 764
rect 277 744 289 764
rect 303 744 315 764
rect 325 744 337 764
rect 355 744 367 764
rect 387 744 399 764
rect 407 744 419 784
rect 451 744 463 764
rect 471 744 483 764
rect 511 744 523 764
rect 531 744 543 764
rect 551 744 563 764
rect 577 744 589 764
rect 597 744 609 764
rect 617 744 629 764
rect 659 744 671 784
rect 689 744 701 784
rect 738 744 750 804
rect 774 744 786 802
rect 837 744 849 784
rect 857 744 869 774
rect 877 744 889 784
rect 897 756 909 784
rect 917 744 929 784
rect 957 744 969 784
rect 977 744 989 772
rect 997 744 1009 784
rect 1017 744 1029 784
rect 1057 744 1069 784
rect 1077 744 1089 772
rect 1097 744 1109 784
rect 1117 744 1129 784
rect 1231 744 1243 764
rect 1251 744 1263 764
rect 1271 744 1283 764
rect 1291 744 1305 764
rect 1337 744 1349 784
rect 1357 744 1369 772
rect 1377 744 1389 784
rect 1397 744 1409 784
rect 1451 744 1463 764
rect 1471 744 1483 764
rect 1501 744 1513 784
rect 1521 744 1533 764
rect 1553 744 1565 764
rect 1583 744 1595 764
rect 1605 744 1617 764
rect 1631 744 1643 764
rect 1659 744 1671 764
rect 1689 744 1701 764
rect 1711 744 1723 784
rect 1737 744 1749 764
rect 1757 744 1769 764
rect 1797 752 1809 772
rect 1817 752 1829 772
rect 1847 752 1859 784
rect 1877 752 1889 792
rect 1917 744 1929 784
rect 1937 744 1949 772
rect 1957 744 1969 784
rect 1977 744 1989 784
rect 2019 744 2031 784
rect 2049 744 2061 784
rect 2097 744 2109 784
rect 2119 744 2131 764
rect 2149 744 2161 764
rect 2177 744 2189 764
rect 2203 744 2215 764
rect 2225 744 2237 764
rect 2255 744 2267 764
rect 2287 744 2299 764
rect 2307 744 2319 784
rect 2337 744 2349 764
rect 2357 744 2369 764
rect 2397 744 2409 784
rect 2417 744 2429 774
rect 2437 744 2449 784
rect 2457 756 2469 784
rect 2477 744 2489 784
rect 2517 744 2529 764
rect 2537 744 2549 764
rect 2557 744 2569 764
rect 2611 744 2623 784
rect 2631 744 2643 784
rect 2651 744 2663 772
rect 2671 744 2683 784
rect 2711 744 2723 784
rect 2731 744 2743 784
rect 2751 744 2763 784
rect 2771 744 2783 784
rect 2791 744 2803 784
rect 2811 744 2823 784
rect 2831 744 2843 784
rect 2851 744 2863 784
rect 2871 744 2883 784
rect 2900 744 2912 784
rect 2928 744 2940 784
rect 2950 744 2962 764
rect 3018 744 3030 764
rect 3040 744 3052 784
rect 3068 744 3080 784
rect 3111 752 3123 792
rect 3141 752 3153 784
rect 3171 752 3183 772
rect 3191 752 3203 772
rect 3231 752 3243 792
rect 3261 752 3273 784
rect 3291 752 3303 772
rect 3311 752 3323 772
rect 3351 744 3363 784
rect 3371 744 3383 784
rect 3391 744 3403 772
rect 3411 744 3423 784
rect 3439 744 3451 784
rect 3469 744 3481 784
rect 3517 752 3529 772
rect 3537 752 3549 772
rect 3567 752 3579 784
rect 3597 752 3609 792
rect 3651 744 3663 764
rect 3671 744 3683 764
rect 3711 752 3723 792
rect 3741 752 3753 784
rect 3771 752 3783 772
rect 3791 752 3803 772
rect 3821 744 3833 784
rect 3841 744 3853 764
rect 3873 744 3885 764
rect 3903 744 3915 764
rect 3925 744 3937 764
rect 3951 744 3963 764
rect 3979 744 3991 764
rect 4009 744 4021 764
rect 4031 744 4043 784
rect 4057 752 4069 772
rect 4077 752 4089 772
rect 4107 752 4119 784
rect 4137 752 4149 792
rect 4180 744 4192 784
rect 4208 744 4220 784
rect 4230 744 4242 764
rect 4277 744 4289 784
rect 4297 744 4309 772
rect 4317 744 4329 784
rect 4337 744 4349 784
rect 4414 744 4426 802
rect 4450 744 4462 804
rect 4477 744 4489 764
rect 4497 744 4509 764
rect 4537 744 4549 784
rect 4557 744 4569 772
rect 4577 744 4589 784
rect 4597 744 4609 784
rect 4639 744 4651 784
rect 4669 744 4681 784
rect 4731 744 4743 764
rect 4751 744 4763 764
rect 4777 744 4789 784
rect 4797 744 4809 772
rect 4817 744 4829 784
rect 4837 744 4849 784
rect 4879 744 4891 784
rect 4909 744 4921 784
rect 4957 752 4969 772
rect 4977 752 4989 772
rect 5007 752 5019 784
rect 5037 752 5049 792
rect 5091 752 5103 792
rect 5121 752 5133 784
rect 5151 752 5163 772
rect 5171 752 5183 772
rect 5197 744 5209 784
rect 5217 744 5229 784
rect 5237 744 5249 784
rect 5257 744 5269 784
rect 5277 744 5289 784
rect 5297 744 5309 784
rect 5317 744 5329 784
rect 5337 744 5349 784
rect 5357 744 5369 784
rect 5400 744 5412 784
rect 5428 744 5440 784
rect 5450 744 5462 764
rect 5511 744 5523 764
rect 5531 744 5543 764
rect 5557 744 5569 784
rect 5577 744 5589 772
rect 5597 744 5609 784
rect 5617 744 5629 784
rect 5659 744 5671 784
rect 5689 744 5701 784
rect 5737 744 5749 784
rect 5757 744 5769 772
rect 5777 744 5789 784
rect 5797 744 5809 784
rect 5874 744 5886 802
rect 5910 744 5922 804
rect 5941 744 5953 784
rect 5961 744 5973 764
rect 5993 744 6005 764
rect 6023 744 6035 764
rect 6045 744 6057 764
rect 6071 744 6083 764
rect 6099 744 6111 764
rect 6129 744 6141 764
rect 6151 744 6163 784
rect 6177 744 6189 784
rect 6197 744 6209 772
rect 6217 744 6229 784
rect 6237 744 6249 784
rect 6277 744 6289 784
rect 6297 744 6309 772
rect 6317 744 6329 784
rect 6337 744 6349 784
rect 6399 744 6411 784
rect 6429 744 6441 784
rect 6461 744 6473 784
rect 6481 744 6493 764
rect 6513 744 6525 764
rect 6543 744 6555 764
rect 6565 744 6577 764
rect 6591 744 6603 764
rect 6619 744 6631 764
rect 6649 744 6661 764
rect 6671 744 6683 784
rect 17 696 29 716
rect 37 696 49 716
rect 79 676 91 716
rect 109 676 121 716
rect 160 676 172 716
rect 188 676 200 716
rect 210 696 222 716
rect 257 696 269 716
rect 277 696 289 716
rect 338 696 350 716
rect 360 676 372 716
rect 388 676 400 716
rect 418 656 430 716
rect 454 658 466 716
rect 539 676 551 716
rect 569 676 581 716
rect 634 658 646 716
rect 670 656 682 716
rect 697 696 709 716
rect 717 696 729 716
rect 757 696 769 716
rect 777 696 789 716
rect 831 696 843 716
rect 851 696 863 716
rect 871 696 883 716
rect 971 696 983 716
rect 991 696 1003 716
rect 1011 696 1023 716
rect 1031 696 1045 716
rect 1081 676 1093 716
rect 1101 696 1113 716
rect 1133 696 1145 716
rect 1163 696 1175 716
rect 1185 696 1197 716
rect 1211 696 1223 716
rect 1239 696 1251 716
rect 1269 696 1281 716
rect 1291 676 1303 716
rect 1317 696 1329 716
rect 1339 676 1351 716
rect 1359 676 1371 716
rect 1399 676 1411 716
rect 1429 676 1441 716
rect 1481 676 1493 716
rect 1501 696 1513 716
rect 1533 696 1545 716
rect 1563 696 1575 716
rect 1585 696 1597 716
rect 1611 696 1623 716
rect 1639 696 1651 716
rect 1669 696 1681 716
rect 1691 676 1703 716
rect 1721 676 1733 716
rect 1741 696 1753 716
rect 1773 696 1785 716
rect 1803 696 1815 716
rect 1825 696 1837 716
rect 1851 696 1863 716
rect 1879 696 1891 716
rect 1909 696 1921 716
rect 1931 676 1943 716
rect 1961 676 1973 716
rect 1981 696 1993 716
rect 2013 696 2025 716
rect 2043 696 2055 716
rect 2065 696 2077 716
rect 2091 696 2103 716
rect 2119 696 2131 716
rect 2149 696 2161 716
rect 2171 676 2183 716
rect 2201 676 2213 716
rect 2221 696 2233 716
rect 2253 696 2265 716
rect 2283 696 2295 716
rect 2305 696 2317 716
rect 2331 696 2343 716
rect 2359 696 2371 716
rect 2389 696 2401 716
rect 2411 676 2423 716
rect 2437 676 2449 716
rect 2459 696 2471 716
rect 2489 696 2501 716
rect 2517 696 2529 716
rect 2543 696 2555 716
rect 2565 696 2577 716
rect 2595 696 2607 716
rect 2627 696 2639 716
rect 2647 676 2659 716
rect 2712 676 2724 716
rect 2740 676 2752 716
rect 2768 676 2780 716
rect 2811 696 2823 716
rect 2831 696 2843 716
rect 2878 696 2890 716
rect 2900 676 2912 716
rect 2928 676 2940 716
rect 2957 696 2969 716
rect 2977 696 2989 716
rect 3017 676 3029 716
rect 3037 688 3049 716
rect 3057 676 3069 716
rect 3077 676 3089 716
rect 3119 676 3131 716
rect 3149 676 3161 716
rect 3198 656 3210 716
rect 3234 658 3246 716
rect 3297 696 3309 716
rect 3317 696 3329 716
rect 3357 676 3369 716
rect 3377 688 3389 716
rect 3397 676 3409 716
rect 3417 676 3429 716
rect 3459 676 3471 716
rect 3489 676 3501 716
rect 3540 676 3552 716
rect 3568 676 3580 716
rect 3590 696 3602 716
rect 3637 696 3649 716
rect 3657 696 3669 716
rect 3677 696 3689 716
rect 3717 676 3729 716
rect 3737 688 3749 716
rect 3757 676 3769 716
rect 3777 676 3789 716
rect 3854 658 3866 716
rect 3890 656 3902 716
rect 3917 676 3929 716
rect 3939 696 3951 716
rect 3969 696 3981 716
rect 3997 696 4009 716
rect 4023 696 4035 716
rect 4045 696 4057 716
rect 4075 696 4087 716
rect 4107 696 4119 716
rect 4127 676 4139 716
rect 4171 696 4183 716
rect 4191 696 4203 716
rect 4211 696 4223 716
rect 4237 676 4249 716
rect 4259 696 4271 716
rect 4289 696 4301 716
rect 4317 696 4329 716
rect 4343 696 4355 716
rect 4365 696 4377 716
rect 4395 696 4407 716
rect 4427 696 4439 716
rect 4447 676 4459 716
rect 4477 696 4489 716
rect 4497 696 4509 716
rect 4540 676 4552 716
rect 4568 676 4580 716
rect 4596 676 4608 716
rect 4678 696 4690 716
rect 4700 676 4712 716
rect 4728 676 4740 716
rect 4771 676 4783 716
rect 4791 676 4803 716
rect 4811 688 4823 716
rect 4831 676 4843 716
rect 4859 676 4871 716
rect 4889 676 4901 716
rect 4951 696 4963 716
rect 4971 696 4983 716
rect 5011 668 5023 708
rect 5041 676 5053 708
rect 5071 688 5083 708
rect 5091 688 5103 708
rect 5118 656 5130 716
rect 5154 658 5166 716
rect 5217 676 5229 716
rect 5239 696 5251 716
rect 5269 696 5281 716
rect 5297 696 5309 716
rect 5323 696 5335 716
rect 5345 696 5357 716
rect 5375 696 5387 716
rect 5407 696 5419 716
rect 5427 676 5439 716
rect 5457 676 5469 716
rect 5477 676 5489 716
rect 5517 688 5529 708
rect 5537 688 5549 708
rect 5567 676 5579 708
rect 5597 668 5609 708
rect 5651 696 5663 716
rect 5671 696 5683 716
rect 5691 696 5703 716
rect 5731 696 5743 716
rect 5751 696 5763 716
rect 5771 696 5783 716
rect 5811 696 5823 716
rect 5831 696 5843 716
rect 5851 696 5863 716
rect 5877 696 5889 716
rect 5897 696 5909 716
rect 5917 696 5929 716
rect 5971 696 5983 716
rect 5991 696 6003 716
rect 6011 696 6023 716
rect 6037 676 6049 716
rect 6057 688 6069 716
rect 6077 676 6089 716
rect 6097 676 6109 716
rect 6137 676 6149 716
rect 6157 688 6169 716
rect 6177 676 6189 716
rect 6197 676 6209 716
rect 6259 676 6271 716
rect 6289 676 6301 716
rect 6321 676 6333 716
rect 6341 696 6353 716
rect 6373 696 6385 716
rect 6403 696 6415 716
rect 6425 696 6437 716
rect 6451 696 6463 716
rect 6479 696 6491 716
rect 6509 696 6521 716
rect 6531 676 6543 716
rect 6557 696 6569 716
rect 6577 696 6589 716
rect 6617 696 6629 716
rect 6637 696 6649 716
rect 17 264 29 304
rect 39 264 51 284
rect 69 264 81 284
rect 97 264 109 284
rect 123 264 135 284
rect 145 264 157 284
rect 175 264 187 284
rect 207 264 219 284
rect 227 264 239 304
rect 261 264 273 304
rect 281 264 293 284
rect 313 264 325 284
rect 343 264 355 284
rect 365 264 377 284
rect 391 264 403 284
rect 419 264 431 284
rect 449 264 461 284
rect 471 264 483 304
rect 498 264 510 324
rect 534 264 546 322
rect 597 264 609 284
rect 617 264 629 284
rect 637 264 649 284
rect 691 264 703 284
rect 711 264 723 284
rect 731 264 743 284
rect 759 264 771 304
rect 789 264 801 304
rect 851 264 863 284
rect 871 264 883 284
rect 901 264 913 304
rect 921 264 933 284
rect 953 264 965 284
rect 983 264 995 284
rect 1005 264 1017 284
rect 1031 264 1043 284
rect 1059 264 1071 284
rect 1089 264 1101 284
rect 1111 264 1123 304
rect 1149 264 1161 304
rect 1169 264 1181 304
rect 1191 264 1203 284
rect 1217 264 1229 284
rect 1239 264 1251 304
rect 1259 264 1271 304
rect 1297 264 1309 284
rect 1319 264 1331 304
rect 1339 264 1351 304
rect 1391 264 1403 284
rect 1411 264 1423 284
rect 1437 264 1449 304
rect 1457 264 1469 292
rect 1477 264 1489 304
rect 1497 264 1509 304
rect 1551 264 1563 284
rect 1571 264 1583 284
rect 1597 264 1609 304
rect 1617 264 1629 292
rect 1637 264 1649 304
rect 1657 264 1669 304
rect 1701 264 1713 304
rect 1721 264 1733 284
rect 1753 264 1765 284
rect 1783 264 1795 284
rect 1805 264 1817 284
rect 1831 264 1843 284
rect 1859 264 1871 284
rect 1889 264 1901 284
rect 1911 264 1923 304
rect 1951 264 1963 284
rect 1971 264 1983 284
rect 2011 264 2023 284
rect 2031 264 2043 284
rect 2057 264 2069 304
rect 2077 264 2089 292
rect 2097 264 2109 304
rect 2117 264 2129 304
rect 2157 264 2169 284
rect 2177 264 2189 284
rect 2217 264 2229 304
rect 2237 264 2249 294
rect 2257 264 2269 304
rect 2277 276 2289 304
rect 2297 264 2309 304
rect 2351 264 2363 304
rect 2371 264 2383 304
rect 2391 264 2403 292
rect 2411 264 2423 304
rect 2437 264 2449 284
rect 2457 264 2469 284
rect 2477 264 2489 284
rect 2521 264 2533 304
rect 2541 264 2553 284
rect 2573 264 2585 284
rect 2603 264 2615 284
rect 2625 264 2637 284
rect 2651 264 2663 284
rect 2679 264 2691 284
rect 2709 264 2721 284
rect 2731 264 2743 304
rect 2771 264 2783 304
rect 2791 264 2803 304
rect 2811 264 2823 292
rect 2831 264 2843 304
rect 2857 264 2869 284
rect 2877 264 2889 284
rect 2897 264 2909 284
rect 2941 264 2953 304
rect 2961 264 2973 284
rect 2993 264 3005 284
rect 3023 264 3035 284
rect 3045 264 3057 284
rect 3071 264 3083 284
rect 3099 264 3111 284
rect 3129 264 3141 284
rect 3151 264 3163 304
rect 3179 264 3191 304
rect 3209 264 3221 304
rect 3271 264 3283 304
rect 3291 264 3303 304
rect 3311 264 3323 292
rect 3331 264 3343 304
rect 3357 264 3369 284
rect 3377 264 3389 284
rect 3397 264 3409 284
rect 3458 264 3470 284
rect 3480 264 3492 304
rect 3508 264 3520 304
rect 3537 264 3549 304
rect 3557 264 3569 292
rect 3577 264 3589 304
rect 3597 264 3609 304
rect 3637 264 3649 284
rect 3657 264 3669 284
rect 3677 264 3689 284
rect 3720 264 3732 304
rect 3748 264 3760 304
rect 3770 264 3782 284
rect 3831 264 3843 284
rect 3851 264 3863 284
rect 3871 264 3883 284
rect 3897 264 3909 304
rect 3917 264 3929 292
rect 3937 264 3949 304
rect 3957 264 3969 304
rect 4034 264 4046 322
rect 4070 264 4082 324
rect 4097 264 4109 284
rect 4117 264 4129 284
rect 4137 264 4149 284
rect 4177 264 4189 304
rect 4199 264 4211 284
rect 4229 264 4241 284
rect 4257 264 4269 284
rect 4283 264 4295 284
rect 4305 264 4317 284
rect 4335 264 4347 284
rect 4367 264 4379 284
rect 4387 264 4399 304
rect 4417 264 4429 284
rect 4437 264 4449 284
rect 4457 264 4469 284
rect 4511 264 4523 304
rect 4531 264 4543 304
rect 4551 264 4563 292
rect 4571 264 4583 304
rect 4597 264 4609 284
rect 4617 264 4629 284
rect 4637 264 4649 284
rect 4691 264 4703 304
rect 4711 276 4723 304
rect 4731 264 4743 304
rect 4751 264 4763 294
rect 4771 264 4783 304
rect 4811 264 4823 284
rect 4831 264 4843 284
rect 4861 264 4873 304
rect 4881 264 4893 284
rect 4913 264 4925 284
rect 4943 264 4955 284
rect 4965 264 4977 284
rect 4991 264 5003 284
rect 5019 264 5031 284
rect 5049 264 5061 284
rect 5071 264 5083 304
rect 5118 264 5130 284
rect 5140 264 5152 304
rect 5168 264 5180 304
rect 5197 264 5209 284
rect 5217 264 5229 284
rect 5237 264 5249 284
rect 5291 264 5303 304
rect 5311 264 5323 304
rect 5331 264 5343 292
rect 5351 264 5363 304
rect 5377 264 5389 284
rect 5397 264 5409 284
rect 5417 264 5429 284
rect 5460 264 5472 304
rect 5488 264 5500 304
rect 5510 264 5522 284
rect 5558 264 5570 324
rect 5594 264 5606 322
rect 5657 264 5669 304
rect 5677 264 5689 292
rect 5697 264 5709 304
rect 5717 264 5729 304
rect 5779 264 5791 304
rect 5809 264 5821 304
rect 5851 264 5863 304
rect 5871 264 5883 304
rect 5891 264 5903 292
rect 5911 264 5923 304
rect 5937 264 5949 304
rect 5957 264 5969 292
rect 5977 264 5989 304
rect 5997 264 6009 304
rect 6037 264 6049 304
rect 6057 264 6069 292
rect 6077 264 6089 304
rect 6097 264 6109 304
rect 6151 264 6163 284
rect 6171 264 6183 284
rect 6191 264 6203 284
rect 6231 264 6243 284
rect 6251 264 6263 284
rect 6271 264 6283 284
rect 6311 264 6323 304
rect 6331 276 6343 304
rect 6351 264 6363 304
rect 6371 264 6383 294
rect 6391 264 6403 304
rect 6421 264 6433 304
rect 6441 264 6453 284
rect 6473 264 6485 284
rect 6503 264 6515 284
rect 6525 264 6537 284
rect 6551 264 6563 284
rect 6579 264 6591 284
rect 6609 264 6621 284
rect 6631 264 6643 304
rect 17 196 29 236
rect 39 216 51 236
rect 69 216 81 236
rect 97 216 109 236
rect 123 216 135 236
rect 145 216 157 236
rect 175 216 187 236
rect 207 216 219 236
rect 227 196 239 236
rect 257 196 269 236
rect 279 216 291 236
rect 309 216 321 236
rect 337 216 349 236
rect 363 216 375 236
rect 385 216 397 236
rect 415 216 427 236
rect 447 216 459 236
rect 467 196 479 236
rect 509 196 521 236
rect 529 196 541 236
rect 551 216 563 236
rect 577 216 589 236
rect 599 196 611 236
rect 619 196 631 236
rect 669 196 681 236
rect 689 196 701 236
rect 711 216 723 236
rect 737 196 749 236
rect 759 216 771 236
rect 789 216 801 236
rect 817 216 829 236
rect 843 216 855 236
rect 865 216 877 236
rect 895 216 907 236
rect 927 216 939 236
rect 947 196 959 236
rect 977 216 989 236
rect 999 196 1011 236
rect 1019 196 1031 236
rect 1079 196 1091 236
rect 1109 196 1121 236
rect 1151 196 1163 236
rect 1171 196 1183 236
rect 1191 208 1203 236
rect 1211 196 1223 236
rect 1241 196 1253 236
rect 1261 216 1273 236
rect 1293 216 1305 236
rect 1323 216 1335 236
rect 1345 216 1357 236
rect 1371 216 1383 236
rect 1399 216 1411 236
rect 1429 216 1441 236
rect 1451 196 1463 236
rect 1491 216 1503 236
rect 1511 216 1523 236
rect 1539 196 1551 236
rect 1569 196 1581 236
rect 1631 196 1643 236
rect 1651 196 1663 236
rect 1671 208 1683 236
rect 1691 196 1703 236
rect 1717 216 1729 236
rect 1737 216 1749 236
rect 1779 196 1791 236
rect 1809 196 1821 236
rect 1859 196 1871 236
rect 1889 196 1901 236
rect 1939 196 1951 236
rect 1969 196 1981 236
rect 2031 196 2043 236
rect 2051 196 2063 236
rect 2071 208 2083 236
rect 2091 196 2103 236
rect 2121 196 2133 236
rect 2141 216 2153 236
rect 2173 216 2185 236
rect 2203 216 2215 236
rect 2225 216 2237 236
rect 2251 216 2263 236
rect 2279 216 2291 236
rect 2309 216 2321 236
rect 2331 196 2343 236
rect 2359 196 2371 236
rect 2389 196 2401 236
rect 2459 196 2471 236
rect 2489 196 2501 236
rect 2531 196 2543 236
rect 2551 196 2563 236
rect 2571 208 2583 236
rect 2591 196 2603 236
rect 2631 216 2643 236
rect 2651 216 2663 236
rect 2681 196 2693 236
rect 2701 216 2713 236
rect 2733 216 2745 236
rect 2763 216 2775 236
rect 2785 216 2797 236
rect 2811 216 2823 236
rect 2839 216 2851 236
rect 2869 216 2881 236
rect 2891 196 2903 236
rect 2931 196 2943 236
rect 2951 196 2963 236
rect 2971 208 2983 236
rect 2991 196 3003 236
rect 3031 216 3043 236
rect 3051 216 3063 236
rect 3071 216 3083 236
rect 3111 196 3123 236
rect 3131 196 3143 224
rect 3151 196 3163 236
rect 3171 206 3183 236
rect 3191 196 3203 236
rect 3231 216 3243 236
rect 3251 216 3263 236
rect 3277 196 3289 236
rect 3299 216 3311 236
rect 3329 216 3341 236
rect 3357 216 3369 236
rect 3383 216 3395 236
rect 3405 216 3417 236
rect 3435 216 3447 236
rect 3467 216 3479 236
rect 3487 196 3499 236
rect 3539 196 3551 236
rect 3569 196 3581 236
rect 3611 196 3623 236
rect 3631 196 3643 236
rect 3651 208 3663 236
rect 3671 196 3683 236
rect 3697 196 3709 236
rect 3717 208 3729 236
rect 3737 196 3749 236
rect 3757 196 3769 236
rect 3797 196 3809 236
rect 3819 216 3831 236
rect 3849 216 3861 236
rect 3877 216 3889 236
rect 3903 216 3915 236
rect 3925 216 3937 236
rect 3955 216 3967 236
rect 3987 216 3999 236
rect 4007 196 4019 236
rect 4037 196 4049 236
rect 4057 208 4069 236
rect 4077 196 4089 236
rect 4097 196 4109 236
rect 4137 196 4149 236
rect 4157 208 4169 236
rect 4177 196 4189 236
rect 4197 196 4209 236
rect 4239 196 4251 236
rect 4269 196 4281 236
rect 4317 196 4329 236
rect 4339 216 4351 236
rect 4369 216 4381 236
rect 4397 216 4409 236
rect 4423 216 4435 236
rect 4445 216 4457 236
rect 4475 216 4487 236
rect 4507 216 4519 236
rect 4527 196 4539 236
rect 4557 196 4569 236
rect 4577 208 4589 236
rect 4597 196 4609 236
rect 4617 196 4629 236
rect 4657 196 4669 236
rect 4677 208 4689 236
rect 4697 196 4709 236
rect 4717 196 4729 236
rect 4759 196 4771 236
rect 4789 196 4801 236
rect 4837 196 4849 236
rect 4859 216 4871 236
rect 4889 216 4901 236
rect 4917 216 4929 236
rect 4943 216 4955 236
rect 4965 216 4977 236
rect 4995 216 5007 236
rect 5027 216 5039 236
rect 5047 196 5059 236
rect 5091 196 5103 236
rect 5111 196 5123 236
rect 5131 208 5143 236
rect 5151 196 5163 236
rect 5177 196 5189 236
rect 5197 208 5209 236
rect 5217 196 5229 236
rect 5237 196 5249 236
rect 5279 196 5291 236
rect 5309 196 5321 236
rect 5357 196 5369 236
rect 5379 216 5391 236
rect 5409 216 5421 236
rect 5437 216 5449 236
rect 5463 216 5475 236
rect 5485 216 5497 236
rect 5515 216 5527 236
rect 5547 216 5559 236
rect 5567 196 5579 236
rect 5597 196 5609 236
rect 5619 216 5631 236
rect 5649 216 5661 236
rect 5677 216 5689 236
rect 5703 216 5715 236
rect 5725 216 5737 236
rect 5755 216 5767 236
rect 5787 216 5799 236
rect 5807 196 5819 236
rect 5837 196 5849 236
rect 5859 216 5871 236
rect 5889 216 5901 236
rect 5917 216 5929 236
rect 5943 216 5955 236
rect 5965 216 5977 236
rect 5995 216 6007 236
rect 6027 216 6039 236
rect 6047 196 6059 236
rect 6091 196 6103 236
rect 6111 196 6123 236
rect 6137 196 6149 236
rect 6157 208 6169 236
rect 6177 196 6189 236
rect 6197 196 6209 236
rect 6251 196 6263 236
rect 6271 196 6283 224
rect 6291 196 6303 236
rect 6311 206 6323 236
rect 6331 196 6343 236
rect 6371 216 6383 236
rect 6391 216 6403 236
rect 6417 196 6429 236
rect 6439 216 6451 236
rect 6469 216 6481 236
rect 6497 216 6509 236
rect 6523 216 6535 236
rect 6545 216 6557 236
rect 6575 216 6587 236
rect 6607 216 6619 236
rect 6627 196 6639 236
<< pdcontact >>
rect 21 6264 33 6344
rect 41 6264 53 6304
rect 75 6264 87 6304
rect 107 6264 119 6304
rect 127 6264 139 6304
rect 153 6264 165 6304
rect 181 6264 193 6284
rect 211 6264 223 6284
rect 231 6264 243 6344
rect 276 6264 288 6304
rect 298 6264 310 6344
rect 326 6264 338 6344
rect 357 6264 369 6304
rect 377 6264 389 6304
rect 397 6264 409 6304
rect 451 6264 463 6304
rect 471 6264 483 6304
rect 491 6264 503 6304
rect 517 6264 529 6304
rect 537 6264 549 6304
rect 557 6264 569 6304
rect 597 6264 609 6344
rect 617 6264 629 6284
rect 647 6264 659 6284
rect 675 6264 687 6304
rect 701 6264 713 6304
rect 721 6264 733 6304
rect 753 6264 765 6304
rect 787 6264 799 6304
rect 807 6264 819 6344
rect 837 6264 849 6304
rect 857 6264 869 6304
rect 897 6264 909 6342
rect 917 6264 929 6330
rect 937 6264 949 6342
rect 957 6276 969 6344
rect 977 6264 989 6344
rect 1031 6264 1043 6304
rect 1051 6264 1063 6304
rect 1077 6264 1089 6344
rect 1097 6264 1109 6284
rect 1127 6264 1139 6284
rect 1155 6264 1167 6304
rect 1181 6264 1193 6304
rect 1201 6264 1213 6304
rect 1233 6264 1245 6304
rect 1267 6264 1279 6304
rect 1287 6264 1299 6344
rect 1317 6264 1329 6344
rect 1347 6264 1369 6344
rect 1387 6264 1399 6344
rect 1456 6264 1468 6304
rect 1478 6264 1490 6344
rect 1506 6264 1518 6344
rect 1547 6264 1559 6344
rect 1567 6264 1579 6344
rect 1591 6264 1603 6304
rect 1611 6264 1623 6304
rect 1651 6264 1663 6304
rect 1671 6264 1683 6304
rect 1697 6264 1709 6344
rect 1717 6264 1729 6284
rect 1747 6264 1759 6284
rect 1775 6264 1787 6304
rect 1801 6264 1813 6304
rect 1821 6264 1833 6304
rect 1853 6264 1865 6304
rect 1887 6264 1899 6304
rect 1907 6264 1919 6344
rect 1942 6264 1954 6344
rect 1970 6264 1982 6344
rect 1992 6264 2004 6304
rect 2037 6264 2049 6304
rect 2057 6264 2069 6304
rect 2077 6264 2089 6304
rect 2136 6264 2148 6304
rect 2158 6264 2170 6344
rect 2186 6264 2198 6344
rect 2231 6264 2243 6344
rect 2251 6264 2263 6344
rect 2271 6264 2283 6332
rect 2291 6264 2303 6336
rect 2331 6264 2343 6304
rect 2351 6264 2363 6304
rect 2371 6264 2383 6304
rect 2423 6264 2435 6344
rect 2451 6264 2463 6344
rect 2477 6264 2489 6344
rect 2505 6264 2517 6344
rect 2557 6264 2569 6304
rect 2577 6264 2589 6304
rect 2597 6264 2609 6304
rect 2651 6264 2663 6304
rect 2671 6264 2683 6300
rect 2691 6264 2703 6304
rect 2711 6264 2723 6304
rect 2737 6264 2749 6304
rect 2757 6264 2769 6304
rect 2777 6264 2789 6304
rect 2831 6264 2843 6304
rect 2851 6264 2863 6300
rect 2871 6264 2883 6304
rect 2891 6264 2903 6304
rect 2936 6264 2948 6304
rect 2958 6264 2970 6344
rect 2986 6264 2998 6344
rect 3036 6264 3048 6304
rect 3058 6264 3070 6344
rect 3086 6264 3098 6344
rect 3131 6264 3143 6304
rect 3151 6264 3163 6304
rect 3191 6264 3203 6304
rect 3211 6264 3223 6304
rect 3237 6264 3249 6336
rect 3257 6264 3269 6332
rect 3277 6264 3289 6344
rect 3297 6264 3309 6344
rect 3342 6264 3354 6344
rect 3370 6264 3382 6344
rect 3392 6264 3404 6304
rect 3451 6264 3463 6344
rect 3471 6264 3483 6344
rect 3491 6264 3503 6332
rect 3511 6264 3523 6336
rect 3551 6264 3563 6344
rect 3571 6264 3583 6344
rect 3591 6264 3603 6332
rect 3611 6264 3623 6336
rect 3637 6264 3649 6304
rect 3657 6264 3669 6304
rect 3677 6264 3689 6300
rect 3697 6264 3709 6304
rect 3756 6264 3768 6304
rect 3778 6264 3790 6344
rect 3806 6264 3818 6344
rect 3842 6264 3854 6344
rect 3870 6264 3882 6344
rect 3892 6264 3904 6304
rect 3937 6264 3949 6304
rect 3957 6264 3969 6304
rect 3997 6264 4009 6304
rect 4017 6264 4029 6304
rect 4037 6264 4049 6304
rect 4087 6264 4099 6344
rect 4107 6264 4119 6344
rect 4131 6264 4143 6304
rect 4151 6264 4163 6304
rect 4177 6264 4189 6304
rect 4197 6264 4209 6304
rect 4217 6264 4229 6304
rect 4271 6264 4283 6304
rect 4291 6264 4303 6300
rect 4311 6264 4323 6304
rect 4331 6264 4343 6304
rect 4371 6264 4383 6304
rect 4391 6264 4403 6300
rect 4411 6264 4423 6304
rect 4431 6264 4443 6304
rect 4471 6264 4483 6304
rect 4491 6264 4503 6300
rect 4511 6264 4523 6304
rect 4531 6264 4543 6304
rect 4557 6264 4569 6304
rect 4577 6264 4589 6304
rect 4617 6264 4629 6336
rect 4637 6264 4649 6332
rect 4657 6264 4669 6344
rect 4677 6264 4689 6344
rect 4717 6264 4729 6336
rect 4737 6264 4749 6332
rect 4757 6264 4769 6344
rect 4777 6264 4789 6344
rect 4822 6264 4834 6344
rect 4850 6264 4862 6344
rect 4872 6264 4884 6304
rect 4936 6264 4948 6304
rect 4958 6264 4970 6344
rect 4986 6264 4998 6344
rect 5022 6264 5034 6344
rect 5050 6264 5062 6344
rect 5072 6264 5084 6304
rect 5131 6264 5143 6304
rect 5151 6264 5163 6300
rect 5171 6264 5183 6304
rect 5191 6264 5203 6304
rect 5231 6264 5243 6304
rect 5251 6264 5263 6300
rect 5271 6264 5283 6304
rect 5291 6264 5303 6304
rect 5331 6264 5343 6304
rect 5351 6264 5363 6300
rect 5371 6264 5383 6304
rect 5391 6264 5403 6304
rect 5417 6264 5429 6336
rect 5437 6264 5449 6332
rect 5457 6264 5469 6344
rect 5477 6264 5489 6344
rect 5531 6264 5543 6344
rect 5551 6264 5563 6344
rect 5571 6264 5583 6332
rect 5591 6264 5603 6336
rect 5631 6264 5643 6304
rect 5651 6264 5663 6304
rect 5677 6264 5689 6336
rect 5697 6264 5709 6332
rect 5717 6264 5729 6344
rect 5737 6264 5749 6344
rect 5777 6264 5789 6304
rect 5797 6264 5809 6304
rect 5817 6264 5829 6300
rect 5837 6264 5849 6304
rect 5891 6264 5903 6344
rect 5911 6264 5923 6344
rect 5931 6264 5943 6332
rect 5951 6264 5963 6336
rect 5991 6264 6003 6304
rect 6011 6264 6023 6304
rect 6051 6264 6063 6344
rect 6071 6264 6083 6344
rect 6091 6264 6103 6332
rect 6111 6264 6123 6336
rect 6156 6264 6168 6304
rect 6178 6264 6190 6344
rect 6206 6264 6218 6344
rect 6251 6264 6263 6344
rect 6271 6264 6283 6344
rect 6291 6264 6303 6332
rect 6311 6264 6323 6336
rect 6337 6264 6349 6304
rect 6357 6264 6369 6304
rect 6377 6264 6389 6300
rect 6397 6264 6409 6304
rect 6451 6264 6463 6304
rect 6471 6264 6483 6300
rect 6491 6264 6503 6304
rect 6511 6264 6523 6304
rect 6537 6264 6549 6304
rect 6557 6264 6569 6304
rect 6597 6264 6609 6342
rect 6617 6264 6629 6330
rect 6637 6264 6649 6342
rect 6657 6276 6669 6344
rect 6677 6264 6689 6344
rect 17 6156 29 6236
rect 37 6216 49 6236
rect 67 6216 79 6236
rect 95 6196 107 6236
rect 121 6196 133 6236
rect 141 6196 153 6236
rect 173 6196 185 6236
rect 207 6196 219 6236
rect 227 6156 239 6236
rect 271 6156 283 6236
rect 291 6156 303 6236
rect 311 6168 323 6236
rect 331 6164 343 6236
rect 371 6196 383 6236
rect 391 6196 403 6236
rect 411 6196 423 6236
rect 437 6156 449 6236
rect 465 6156 477 6236
rect 531 6196 543 6236
rect 551 6196 563 6236
rect 571 6196 583 6236
rect 602 6156 614 6236
rect 630 6156 642 6236
rect 652 6196 664 6236
rect 716 6196 728 6236
rect 738 6156 750 6236
rect 766 6156 778 6236
rect 797 6156 809 6236
rect 825 6156 837 6236
rect 891 6156 903 6236
rect 911 6156 923 6236
rect 931 6168 943 6236
rect 951 6164 963 6236
rect 977 6156 989 6236
rect 1007 6157 1019 6236
rect 1027 6157 1039 6236
rect 1091 6196 1103 6236
rect 1111 6196 1123 6236
rect 1137 6156 1149 6236
rect 1165 6156 1177 6236
rect 1236 6196 1248 6236
rect 1258 6156 1270 6236
rect 1286 6156 1298 6236
rect 1331 6196 1343 6236
rect 1351 6196 1363 6236
rect 1391 6196 1403 6236
rect 1411 6196 1423 6236
rect 1437 6156 1449 6236
rect 1465 6156 1477 6236
rect 1517 6156 1529 6236
rect 1545 6156 1557 6236
rect 1597 6196 1609 6236
rect 1617 6196 1629 6236
rect 1657 6156 1669 6236
rect 1685 6156 1697 6236
rect 1737 6156 1749 6236
rect 1765 6156 1777 6236
rect 1822 6156 1834 6236
rect 1850 6156 1862 6236
rect 1872 6196 1884 6236
rect 1917 6196 1929 6236
rect 1937 6196 1949 6236
rect 1991 6156 2003 6236
rect 2011 6156 2023 6236
rect 2031 6168 2043 6236
rect 2051 6164 2063 6236
rect 2077 6196 2089 6236
rect 2097 6196 2109 6236
rect 2156 6196 2168 6236
rect 2178 6156 2190 6236
rect 2206 6156 2218 6236
rect 2237 6196 2249 6236
rect 2257 6196 2269 6236
rect 2316 6196 2328 6236
rect 2338 6156 2350 6236
rect 2366 6156 2378 6236
rect 2411 6196 2423 6236
rect 2431 6200 2443 6236
rect 2451 6196 2463 6236
rect 2471 6196 2483 6236
rect 2511 6156 2523 6236
rect 2531 6156 2543 6236
rect 2551 6168 2563 6236
rect 2571 6164 2583 6236
rect 2623 6156 2635 6236
rect 2651 6156 2663 6236
rect 2691 6196 2703 6236
rect 2711 6200 2723 6236
rect 2731 6196 2743 6236
rect 2751 6196 2763 6236
rect 2791 6156 2803 6236
rect 2811 6156 2823 6224
rect 2831 6158 2843 6236
rect 2851 6170 2863 6236
rect 2871 6158 2883 6236
rect 2911 6196 2923 6236
rect 2931 6196 2943 6236
rect 2957 6196 2969 6236
rect 2977 6196 2989 6236
rect 2997 6200 3009 6236
rect 3017 6196 3029 6236
rect 3071 6156 3083 6236
rect 3091 6156 3103 6236
rect 3111 6168 3123 6236
rect 3131 6164 3143 6236
rect 3171 6196 3183 6236
rect 3191 6200 3203 6236
rect 3211 6196 3223 6236
rect 3231 6196 3243 6236
rect 3271 6156 3283 6236
rect 3291 6156 3303 6236
rect 3311 6168 3323 6236
rect 3331 6164 3343 6236
rect 3371 6196 3383 6236
rect 3391 6196 3403 6236
rect 3431 6196 3443 6236
rect 3451 6200 3463 6236
rect 3471 6196 3483 6236
rect 3491 6196 3503 6236
rect 3517 6196 3529 6236
rect 3537 6196 3549 6236
rect 3557 6200 3569 6236
rect 3577 6196 3589 6236
rect 3617 6196 3629 6236
rect 3637 6196 3649 6236
rect 3677 6164 3689 6236
rect 3697 6168 3709 6236
rect 3717 6156 3729 6236
rect 3737 6156 3749 6236
rect 3791 6196 3803 6236
rect 3811 6196 3823 6236
rect 3831 6196 3843 6236
rect 3857 6196 3869 6236
rect 3877 6196 3889 6236
rect 3897 6196 3909 6236
rect 3956 6196 3968 6236
rect 3978 6156 3990 6236
rect 4006 6156 4018 6236
rect 4042 6156 4054 6236
rect 4070 6156 4082 6236
rect 4092 6196 4104 6236
rect 4163 6156 4175 6236
rect 4191 6156 4203 6236
rect 4217 6196 4229 6236
rect 4237 6196 4249 6236
rect 4291 6196 4303 6236
rect 4311 6196 4323 6236
rect 4331 6196 4343 6236
rect 4357 6196 4369 6236
rect 4377 6196 4389 6236
rect 4401 6156 4413 6236
rect 4421 6156 4433 6236
rect 4476 6196 4488 6236
rect 4498 6156 4510 6236
rect 4526 6156 4538 6236
rect 4571 6156 4583 6236
rect 4591 6156 4603 6236
rect 4611 6168 4623 6236
rect 4631 6164 4643 6236
rect 4657 6196 4669 6236
rect 4677 6196 4689 6236
rect 4697 6200 4709 6236
rect 4717 6196 4729 6236
rect 4771 6156 4783 6236
rect 4791 6156 4803 6236
rect 4811 6168 4823 6236
rect 4831 6164 4843 6236
rect 4871 6196 4883 6236
rect 4891 6200 4903 6236
rect 4911 6196 4923 6236
rect 4931 6196 4943 6236
rect 4957 6196 4969 6236
rect 4977 6196 4989 6236
rect 4997 6200 5009 6236
rect 5017 6196 5029 6236
rect 5076 6196 5088 6236
rect 5098 6156 5110 6236
rect 5126 6156 5138 6236
rect 5171 6196 5183 6236
rect 5191 6196 5203 6236
rect 5211 6196 5223 6236
rect 5237 6196 5249 6236
rect 5257 6196 5269 6236
rect 5281 6156 5293 6236
rect 5301 6156 5313 6236
rect 5342 6156 5354 6236
rect 5370 6156 5382 6236
rect 5392 6196 5404 6236
rect 5451 6156 5463 6236
rect 5471 6156 5483 6236
rect 5491 6168 5503 6236
rect 5511 6164 5523 6236
rect 5551 6196 5563 6236
rect 5571 6200 5583 6236
rect 5591 6196 5603 6236
rect 5611 6196 5623 6236
rect 5637 6196 5649 6236
rect 5657 6196 5669 6236
rect 5677 6200 5689 6236
rect 5697 6196 5709 6236
rect 5751 6156 5763 6236
rect 5771 6156 5783 6236
rect 5791 6168 5803 6236
rect 5811 6164 5823 6236
rect 5837 6196 5849 6236
rect 5857 6196 5869 6236
rect 5877 6200 5889 6236
rect 5897 6196 5909 6236
rect 5942 6156 5954 6236
rect 5970 6156 5982 6236
rect 5992 6196 6004 6236
rect 6042 6156 6054 6236
rect 6070 6156 6082 6236
rect 6092 6196 6104 6236
rect 6137 6196 6149 6236
rect 6157 6196 6169 6236
rect 6177 6200 6189 6236
rect 6197 6196 6209 6236
rect 6237 6196 6249 6236
rect 6257 6196 6269 6236
rect 6277 6200 6289 6236
rect 6297 6196 6309 6236
rect 6351 6196 6363 6236
rect 6371 6200 6383 6236
rect 6391 6196 6403 6236
rect 6411 6196 6423 6236
rect 6451 6156 6463 6236
rect 6471 6156 6483 6236
rect 6491 6168 6503 6236
rect 6511 6164 6523 6236
rect 6537 6196 6549 6236
rect 6557 6196 6569 6236
rect 6597 6196 6609 6236
rect 6617 6196 6629 6236
rect 29 5784 41 5864
rect 49 5784 61 5864
rect 71 5784 83 5824
rect 97 5784 109 5824
rect 117 5784 129 5824
rect 137 5784 149 5824
rect 177 5784 189 5824
rect 197 5784 209 5824
rect 217 5784 229 5824
rect 271 5784 283 5864
rect 291 5784 303 5864
rect 311 5784 323 5852
rect 331 5784 343 5856
rect 371 5784 383 5824
rect 391 5784 403 5824
rect 411 5784 423 5824
rect 437 5784 449 5824
rect 457 5784 469 5824
rect 523 5784 535 5864
rect 551 5784 563 5864
rect 577 5784 589 5864
rect 605 5784 617 5864
rect 662 5784 674 5864
rect 690 5784 702 5864
rect 712 5784 724 5824
rect 771 5784 783 5824
rect 791 5784 803 5824
rect 817 5784 829 5864
rect 845 5784 857 5864
rect 911 5784 923 5824
rect 931 5784 943 5824
rect 951 5784 963 5824
rect 996 5784 1008 5824
rect 1018 5784 1030 5864
rect 1046 5784 1058 5864
rect 1077 5784 1089 5864
rect 1105 5784 1117 5864
rect 1171 5784 1183 5824
rect 1191 5784 1203 5824
rect 1217 5784 1229 5864
rect 1237 5784 1249 5804
rect 1267 5784 1279 5804
rect 1295 5784 1307 5824
rect 1321 5784 1333 5824
rect 1341 5784 1353 5824
rect 1373 5784 1385 5824
rect 1407 5784 1419 5824
rect 1427 5784 1439 5864
rect 1457 5784 1469 5824
rect 1477 5784 1489 5824
rect 1497 5784 1509 5824
rect 1551 5784 1563 5824
rect 1571 5784 1583 5820
rect 1591 5784 1603 5824
rect 1611 5784 1623 5824
rect 1656 5784 1668 5824
rect 1678 5784 1690 5864
rect 1706 5784 1718 5864
rect 1763 5784 1775 5864
rect 1791 5784 1803 5864
rect 1831 5784 1843 5824
rect 1851 5784 1863 5820
rect 1871 5784 1883 5824
rect 1891 5784 1903 5824
rect 1917 5784 1929 5824
rect 1937 5784 1949 5824
rect 1996 5784 2008 5824
rect 2018 5784 2030 5864
rect 2046 5784 2058 5864
rect 2077 5784 2089 5824
rect 2097 5784 2109 5824
rect 2117 5784 2129 5820
rect 2137 5784 2149 5824
rect 2191 5784 2203 5864
rect 2211 5784 2223 5864
rect 2231 5784 2243 5852
rect 2251 5784 2263 5856
rect 2282 5784 2294 5864
rect 2310 5784 2322 5864
rect 2332 5784 2344 5824
rect 2391 5784 2403 5824
rect 2411 5784 2423 5824
rect 2431 5784 2443 5824
rect 2471 5784 2483 5824
rect 2491 5784 2503 5820
rect 2511 5784 2523 5824
rect 2531 5784 2543 5824
rect 2571 5784 2583 5864
rect 2591 5784 2603 5864
rect 2611 5784 2623 5852
rect 2631 5784 2643 5856
rect 2657 5784 2669 5824
rect 2677 5784 2689 5824
rect 2697 5784 2709 5824
rect 2751 5784 2763 5824
rect 2771 5784 2783 5820
rect 2791 5784 2803 5824
rect 2811 5784 2823 5824
rect 2851 5784 2863 5824
rect 2871 5784 2883 5820
rect 2891 5784 2903 5824
rect 2911 5784 2923 5824
rect 2951 5784 2963 5824
rect 2971 5784 2983 5820
rect 2991 5784 3003 5824
rect 3011 5784 3023 5824
rect 3051 5784 3063 5824
rect 3071 5784 3083 5820
rect 3091 5784 3103 5824
rect 3111 5784 3123 5824
rect 3137 5784 3149 5824
rect 3157 5784 3169 5824
rect 3177 5784 3189 5820
rect 3197 5784 3209 5824
rect 3256 5784 3268 5824
rect 3278 5784 3290 5864
rect 3306 5784 3318 5864
rect 3342 5784 3354 5864
rect 3370 5784 3382 5864
rect 3392 5784 3404 5824
rect 3451 5784 3463 5864
rect 3471 5784 3483 5864
rect 3491 5784 3503 5852
rect 3511 5784 3523 5856
rect 3556 5784 3568 5824
rect 3578 5784 3590 5864
rect 3606 5784 3618 5864
rect 3651 5784 3663 5824
rect 3671 5784 3683 5820
rect 3691 5784 3703 5824
rect 3711 5784 3723 5824
rect 3737 5784 3749 5856
rect 3757 5784 3769 5852
rect 3777 5784 3789 5864
rect 3797 5784 3809 5864
rect 3851 5784 3863 5824
rect 3871 5784 3883 5820
rect 3891 5784 3903 5824
rect 3911 5784 3923 5824
rect 3951 5784 3963 5864
rect 3971 5784 3983 5864
rect 3991 5784 4003 5852
rect 4011 5784 4023 5856
rect 4051 5784 4063 5824
rect 4071 5784 4083 5820
rect 4091 5784 4103 5824
rect 4111 5784 4123 5824
rect 4151 5784 4163 5864
rect 4171 5784 4183 5864
rect 4191 5784 4203 5852
rect 4211 5784 4223 5856
rect 4237 5784 4249 5824
rect 4257 5784 4269 5824
rect 4277 5784 4289 5820
rect 4297 5784 4309 5824
rect 4337 5784 4349 5824
rect 4357 5784 4369 5824
rect 4377 5784 4389 5824
rect 4436 5784 4448 5824
rect 4458 5784 4470 5864
rect 4486 5784 4498 5864
rect 4543 5784 4555 5864
rect 4571 5784 4583 5864
rect 4597 5784 4609 5824
rect 4617 5784 4629 5824
rect 4641 5784 4653 5864
rect 4661 5784 4673 5864
rect 4711 5784 4723 5864
rect 4731 5784 4743 5864
rect 4751 5784 4763 5852
rect 4771 5784 4783 5856
rect 4797 5784 4809 5824
rect 4817 5784 4829 5824
rect 4837 5784 4849 5824
rect 4891 5784 4903 5824
rect 4911 5784 4923 5824
rect 4951 5784 4963 5824
rect 4971 5784 4983 5820
rect 4991 5784 5003 5824
rect 5011 5784 5023 5824
rect 5037 5784 5049 5856
rect 5057 5784 5069 5852
rect 5077 5784 5089 5864
rect 5097 5784 5109 5864
rect 5142 5784 5154 5864
rect 5170 5784 5182 5864
rect 5192 5784 5204 5824
rect 5242 5784 5254 5864
rect 5270 5784 5282 5864
rect 5292 5784 5304 5824
rect 5337 5784 5349 5862
rect 5357 5784 5369 5850
rect 5377 5784 5389 5862
rect 5397 5796 5409 5864
rect 5417 5784 5429 5864
rect 5471 5784 5483 5824
rect 5491 5784 5503 5824
rect 5511 5784 5523 5824
rect 5537 5784 5549 5824
rect 5557 5784 5569 5824
rect 5611 5784 5623 5824
rect 5631 5784 5643 5820
rect 5651 5784 5663 5824
rect 5671 5784 5683 5824
rect 5697 5784 5709 5856
rect 5717 5784 5729 5852
rect 5737 5784 5749 5864
rect 5757 5784 5769 5864
rect 5816 5784 5828 5824
rect 5838 5784 5850 5864
rect 5866 5784 5878 5864
rect 5902 5784 5914 5864
rect 5930 5784 5942 5864
rect 5952 5784 5964 5824
rect 6016 5784 6028 5824
rect 6038 5784 6050 5864
rect 6066 5784 6078 5864
rect 6097 5784 6109 5862
rect 6117 5784 6129 5850
rect 6137 5784 6149 5862
rect 6157 5796 6169 5864
rect 6177 5784 6189 5864
rect 6231 5784 6243 5824
rect 6251 5784 6263 5824
rect 6271 5784 6283 5824
rect 6297 5784 6309 5824
rect 6317 5784 6329 5824
rect 6341 5784 6353 5864
rect 6361 5784 6373 5864
rect 6402 5784 6414 5864
rect 6430 5784 6442 5864
rect 6452 5784 6464 5824
rect 6497 5784 6509 5824
rect 6517 5784 6529 5824
rect 6537 5784 6549 5820
rect 6557 5784 6569 5824
rect 6597 5784 6609 5824
rect 6617 5784 6629 5824
rect 6637 5784 6649 5824
rect 29 5676 41 5756
rect 49 5676 61 5756
rect 71 5716 83 5756
rect 109 5676 121 5756
rect 129 5676 141 5756
rect 151 5716 163 5756
rect 177 5676 189 5756
rect 197 5736 209 5756
rect 227 5736 239 5756
rect 255 5716 267 5756
rect 281 5716 293 5756
rect 301 5716 313 5756
rect 333 5716 345 5756
rect 367 5716 379 5756
rect 387 5676 399 5756
rect 443 5676 455 5756
rect 471 5676 483 5756
rect 497 5684 509 5756
rect 517 5688 529 5756
rect 537 5676 549 5756
rect 557 5676 569 5756
rect 597 5716 609 5756
rect 617 5716 629 5756
rect 637 5716 649 5756
rect 677 5716 689 5756
rect 697 5716 709 5756
rect 721 5676 733 5756
rect 741 5676 753 5756
rect 777 5716 789 5756
rect 797 5716 809 5756
rect 817 5716 829 5756
rect 857 5716 869 5756
rect 877 5716 889 5756
rect 897 5716 909 5756
rect 937 5676 949 5756
rect 965 5676 977 5756
rect 1017 5716 1029 5756
rect 1037 5716 1049 5756
rect 1077 5676 1089 5756
rect 1107 5677 1119 5756
rect 1127 5677 1139 5756
rect 1177 5676 1189 5756
rect 1205 5676 1217 5756
rect 1257 5716 1269 5756
rect 1277 5716 1289 5756
rect 1317 5676 1329 5756
rect 1345 5676 1357 5756
rect 1397 5716 1409 5756
rect 1417 5716 1429 5756
rect 1457 5676 1469 5756
rect 1477 5736 1489 5756
rect 1507 5736 1519 5756
rect 1535 5716 1547 5756
rect 1561 5716 1573 5756
rect 1581 5716 1593 5756
rect 1613 5716 1625 5756
rect 1647 5716 1659 5756
rect 1667 5676 1679 5756
rect 1697 5676 1709 5756
rect 1727 5676 1749 5756
rect 1767 5676 1779 5756
rect 1836 5716 1848 5756
rect 1858 5676 1870 5756
rect 1886 5676 1898 5756
rect 1931 5716 1943 5756
rect 1951 5716 1963 5756
rect 1971 5716 1983 5756
rect 1997 5716 2009 5756
rect 2017 5716 2029 5756
rect 2071 5676 2083 5756
rect 2091 5676 2103 5756
rect 2111 5688 2123 5756
rect 2131 5684 2143 5756
rect 2157 5676 2169 5756
rect 2185 5676 2197 5756
rect 2237 5716 2249 5756
rect 2257 5716 2269 5756
rect 2277 5716 2289 5756
rect 2327 5688 2339 5748
rect 2347 5692 2359 5744
rect 2367 5688 2379 5748
rect 2391 5698 2403 5756
rect 2411 5696 2423 5744
rect 2431 5696 2443 5756
rect 2451 5696 2463 5756
rect 2471 5696 2483 5756
rect 2511 5716 2523 5756
rect 2531 5716 2543 5756
rect 2551 5716 2563 5756
rect 2591 5716 2603 5756
rect 2611 5720 2623 5756
rect 2631 5716 2643 5756
rect 2651 5716 2663 5756
rect 2691 5716 2703 5756
rect 2711 5720 2723 5756
rect 2731 5716 2743 5756
rect 2751 5716 2763 5756
rect 2777 5716 2789 5756
rect 2797 5716 2809 5756
rect 2817 5716 2829 5756
rect 2862 5676 2874 5756
rect 2890 5676 2902 5756
rect 2912 5716 2924 5756
rect 2971 5716 2983 5756
rect 2991 5720 3003 5756
rect 3011 5716 3023 5756
rect 3031 5716 3043 5756
rect 3057 5684 3069 5756
rect 3077 5688 3089 5756
rect 3097 5676 3109 5756
rect 3117 5676 3129 5756
rect 3176 5716 3188 5756
rect 3198 5676 3210 5756
rect 3226 5676 3238 5756
rect 3271 5716 3283 5756
rect 3291 5716 3303 5756
rect 3317 5716 3329 5756
rect 3337 5716 3349 5756
rect 3357 5720 3369 5756
rect 3377 5716 3389 5756
rect 3431 5716 3443 5756
rect 3451 5720 3463 5756
rect 3471 5716 3483 5756
rect 3491 5716 3503 5756
rect 3531 5716 3543 5756
rect 3551 5720 3563 5756
rect 3571 5716 3583 5756
rect 3591 5716 3603 5756
rect 3631 5716 3643 5756
rect 3651 5716 3663 5756
rect 3696 5716 3708 5756
rect 3718 5676 3730 5756
rect 3746 5676 3758 5756
rect 3803 5676 3815 5756
rect 3831 5676 3843 5756
rect 3862 5676 3874 5756
rect 3890 5676 3902 5756
rect 3912 5716 3924 5756
rect 3971 5716 3983 5756
rect 3991 5716 4003 5756
rect 4031 5676 4043 5756
rect 4051 5676 4063 5744
rect 4071 5678 4083 5756
rect 4091 5690 4103 5756
rect 4111 5678 4123 5756
rect 4156 5716 4168 5756
rect 4178 5676 4190 5756
rect 4206 5676 4218 5756
rect 4251 5716 4263 5756
rect 4271 5720 4283 5756
rect 4291 5716 4303 5756
rect 4311 5716 4323 5756
rect 4337 5716 4349 5756
rect 4357 5716 4369 5756
rect 4416 5716 4428 5756
rect 4438 5676 4450 5756
rect 4466 5676 4478 5756
rect 4507 5676 4519 5756
rect 4527 5676 4539 5756
rect 4551 5716 4563 5756
rect 4571 5716 4583 5756
rect 4597 5716 4609 5756
rect 4617 5716 4629 5756
rect 4637 5716 4649 5756
rect 4696 5716 4708 5756
rect 4718 5676 4730 5756
rect 4746 5676 4758 5756
rect 4782 5676 4794 5756
rect 4810 5676 4822 5756
rect 4832 5716 4844 5756
rect 4891 5716 4903 5756
rect 4911 5720 4923 5756
rect 4931 5716 4943 5756
rect 4951 5716 4963 5756
rect 4977 5684 4989 5756
rect 4997 5688 5009 5756
rect 5017 5676 5029 5756
rect 5037 5676 5049 5756
rect 5082 5676 5094 5756
rect 5110 5676 5122 5756
rect 5132 5716 5144 5756
rect 5177 5716 5189 5756
rect 5197 5716 5209 5756
rect 5217 5720 5229 5756
rect 5237 5716 5249 5756
rect 5277 5716 5289 5756
rect 5297 5716 5309 5756
rect 5317 5716 5329 5756
rect 5357 5716 5369 5756
rect 5377 5716 5389 5756
rect 5397 5720 5409 5756
rect 5417 5716 5429 5756
rect 5457 5684 5469 5756
rect 5477 5688 5489 5756
rect 5497 5676 5509 5756
rect 5517 5676 5529 5756
rect 5557 5716 5569 5756
rect 5577 5716 5589 5756
rect 5597 5716 5609 5756
rect 5651 5716 5663 5756
rect 5671 5716 5683 5756
rect 5691 5716 5703 5756
rect 5717 5678 5729 5756
rect 5737 5690 5749 5756
rect 5757 5678 5769 5756
rect 5777 5676 5789 5744
rect 5797 5676 5809 5756
rect 5856 5716 5868 5756
rect 5878 5676 5890 5756
rect 5906 5676 5918 5756
rect 5937 5716 5949 5756
rect 5957 5716 5969 5756
rect 5997 5678 6009 5756
rect 6017 5690 6029 5756
rect 6037 5678 6049 5756
rect 6057 5676 6069 5744
rect 6077 5676 6089 5756
rect 6117 5716 6129 5756
rect 6137 5716 6149 5756
rect 6157 5720 6169 5756
rect 6177 5716 6189 5756
rect 6231 5716 6243 5756
rect 6251 5716 6263 5756
rect 6277 5684 6289 5756
rect 6297 5688 6309 5756
rect 6317 5676 6329 5756
rect 6337 5676 6349 5756
rect 6377 5716 6389 5756
rect 6397 5716 6409 5756
rect 6417 5720 6429 5756
rect 6437 5716 6449 5756
rect 6477 5716 6489 5756
rect 6497 5716 6509 5756
rect 6517 5720 6529 5756
rect 6537 5716 6549 5756
rect 6577 5716 6589 5756
rect 6597 5716 6609 5756
rect 6617 5720 6629 5756
rect 6637 5716 6649 5756
rect 17 5304 29 5384
rect 37 5304 49 5324
rect 67 5304 79 5324
rect 95 5304 107 5344
rect 121 5304 133 5344
rect 141 5304 153 5344
rect 173 5304 185 5344
rect 207 5304 219 5344
rect 227 5304 239 5384
rect 257 5304 269 5344
rect 277 5304 289 5344
rect 297 5304 309 5344
rect 351 5304 363 5384
rect 371 5304 383 5384
rect 391 5304 403 5372
rect 411 5304 423 5376
rect 451 5304 463 5344
rect 471 5304 483 5344
rect 491 5304 503 5344
rect 527 5304 539 5384
rect 547 5304 559 5384
rect 571 5304 583 5344
rect 591 5304 603 5344
rect 617 5304 629 5384
rect 645 5304 657 5384
rect 697 5304 709 5384
rect 725 5304 737 5384
rect 777 5304 789 5344
rect 797 5304 809 5344
rect 817 5304 829 5344
rect 857 5304 869 5344
rect 877 5304 889 5344
rect 897 5304 909 5344
rect 937 5304 949 5344
rect 957 5304 969 5344
rect 997 5304 1009 5376
rect 1017 5304 1029 5372
rect 1037 5304 1049 5384
rect 1057 5304 1069 5384
rect 1111 5304 1123 5384
rect 1131 5316 1143 5384
rect 1151 5304 1163 5382
rect 1171 5304 1183 5370
rect 1191 5304 1203 5382
rect 1217 5304 1229 5384
rect 1237 5304 1249 5324
rect 1267 5304 1279 5324
rect 1295 5304 1307 5344
rect 1321 5304 1333 5344
rect 1341 5304 1353 5344
rect 1373 5304 1385 5344
rect 1407 5304 1419 5344
rect 1427 5304 1439 5384
rect 1471 5304 1483 5344
rect 1491 5304 1503 5340
rect 1511 5304 1523 5344
rect 1531 5304 1543 5344
rect 1571 5304 1583 5344
rect 1591 5304 1603 5340
rect 1611 5304 1623 5344
rect 1631 5304 1643 5344
rect 1671 5304 1683 5344
rect 1691 5304 1703 5344
rect 1736 5304 1748 5344
rect 1758 5304 1770 5384
rect 1786 5304 1798 5384
rect 1827 5304 1839 5384
rect 1847 5304 1859 5384
rect 1871 5304 1883 5344
rect 1891 5304 1903 5344
rect 1931 5304 1943 5344
rect 1951 5304 1963 5344
rect 1971 5304 1983 5344
rect 2016 5304 2028 5344
rect 2038 5304 2050 5384
rect 2066 5304 2078 5384
rect 2097 5304 2109 5344
rect 2117 5304 2129 5344
rect 2137 5304 2149 5344
rect 2191 5304 2203 5344
rect 2211 5304 2223 5344
rect 2256 5304 2268 5344
rect 2278 5304 2290 5384
rect 2306 5304 2318 5384
rect 2337 5304 2349 5384
rect 2365 5304 2377 5384
rect 2431 5304 2443 5344
rect 2451 5304 2463 5344
rect 2491 5304 2503 5384
rect 2511 5304 2523 5384
rect 2531 5304 2543 5372
rect 2551 5304 2563 5376
rect 2582 5304 2594 5384
rect 2610 5304 2622 5384
rect 2632 5304 2644 5344
rect 2677 5304 2689 5344
rect 2697 5304 2709 5344
rect 2717 5304 2729 5344
rect 2771 5304 2783 5344
rect 2791 5304 2803 5340
rect 2811 5304 2823 5344
rect 2831 5304 2843 5344
rect 2871 5304 2883 5344
rect 2891 5304 2903 5344
rect 2911 5304 2923 5344
rect 2963 5304 2975 5384
rect 2991 5304 3003 5384
rect 3022 5304 3034 5384
rect 3050 5304 3062 5384
rect 3072 5304 3084 5344
rect 3131 5304 3143 5344
rect 3151 5304 3163 5344
rect 3171 5304 3183 5344
rect 3202 5304 3214 5384
rect 3230 5304 3242 5384
rect 3252 5304 3264 5344
rect 3307 5304 3319 5384
rect 3327 5304 3339 5384
rect 3351 5304 3363 5344
rect 3371 5304 3383 5344
rect 3397 5304 3409 5384
rect 3425 5304 3437 5384
rect 3477 5304 3489 5384
rect 3507 5304 3519 5383
rect 3527 5304 3539 5383
rect 3582 5304 3594 5384
rect 3610 5304 3622 5384
rect 3632 5304 3644 5344
rect 3703 5304 3715 5384
rect 3731 5304 3743 5384
rect 3757 5304 3769 5384
rect 3787 5304 3809 5384
rect 3827 5304 3839 5384
rect 3903 5304 3915 5384
rect 3931 5304 3943 5384
rect 3962 5304 3974 5384
rect 3990 5304 4002 5384
rect 4012 5304 4024 5344
rect 4071 5304 4083 5344
rect 4091 5304 4103 5340
rect 4111 5304 4123 5344
rect 4131 5304 4143 5344
rect 4171 5304 4183 5344
rect 4191 5304 4203 5344
rect 4211 5304 4223 5344
rect 4237 5304 4249 5344
rect 4257 5304 4269 5344
rect 4316 5304 4328 5344
rect 4338 5304 4350 5384
rect 4366 5304 4378 5384
rect 4411 5304 4423 5344
rect 4431 5304 4443 5344
rect 4451 5304 4463 5344
rect 4477 5304 4489 5344
rect 4497 5304 4509 5344
rect 4517 5304 4529 5344
rect 4576 5304 4588 5344
rect 4598 5304 4610 5384
rect 4626 5304 4638 5384
rect 4676 5304 4688 5344
rect 4698 5304 4710 5384
rect 4726 5304 4738 5384
rect 4767 5304 4779 5384
rect 4787 5304 4799 5384
rect 4811 5304 4823 5344
rect 4831 5304 4843 5344
rect 4876 5304 4888 5344
rect 4898 5304 4910 5384
rect 4926 5304 4938 5384
rect 4971 5304 4983 5344
rect 4991 5304 5003 5344
rect 5011 5304 5023 5344
rect 5047 5304 5059 5384
rect 5067 5304 5079 5384
rect 5091 5304 5103 5344
rect 5111 5304 5123 5344
rect 5137 5304 5149 5344
rect 5157 5304 5169 5344
rect 5177 5304 5189 5344
rect 5222 5304 5234 5384
rect 5250 5304 5262 5384
rect 5272 5304 5284 5344
rect 5327 5304 5339 5384
rect 5347 5304 5359 5384
rect 5371 5304 5383 5344
rect 5391 5304 5403 5344
rect 5422 5304 5434 5384
rect 5450 5304 5462 5384
rect 5472 5304 5484 5344
rect 5517 5304 5529 5344
rect 5537 5304 5549 5344
rect 5557 5304 5569 5344
rect 5597 5304 5609 5344
rect 5617 5304 5629 5344
rect 5637 5304 5649 5340
rect 5657 5304 5669 5344
rect 5707 5304 5719 5384
rect 5727 5304 5739 5384
rect 5751 5304 5763 5344
rect 5771 5304 5783 5344
rect 5811 5304 5823 5384
rect 5831 5316 5843 5384
rect 5851 5304 5863 5382
rect 5871 5304 5883 5370
rect 5891 5304 5903 5382
rect 5917 5304 5929 5344
rect 5937 5304 5949 5344
rect 5957 5304 5969 5344
rect 5997 5304 6009 5344
rect 6017 5304 6029 5344
rect 6037 5304 6049 5340
rect 6057 5304 6069 5344
rect 6097 5304 6109 5376
rect 6117 5304 6129 5372
rect 6137 5304 6149 5384
rect 6157 5304 6169 5384
rect 6216 5304 6228 5344
rect 6238 5304 6250 5384
rect 6266 5304 6278 5384
rect 6302 5304 6314 5384
rect 6330 5304 6342 5384
rect 6352 5304 6364 5344
rect 6416 5304 6428 5344
rect 6438 5304 6450 5384
rect 6466 5304 6478 5384
rect 6511 5304 6523 5344
rect 6531 5304 6543 5340
rect 6551 5304 6563 5344
rect 6571 5304 6583 5344
rect 6611 5304 6623 5384
rect 6631 5304 6643 5384
rect 6651 5304 6663 5372
rect 6671 5304 6683 5376
rect 29 5196 41 5276
rect 49 5196 61 5276
rect 71 5236 83 5276
rect 97 5196 109 5276
rect 117 5256 129 5276
rect 147 5256 159 5276
rect 175 5236 187 5276
rect 201 5236 213 5276
rect 221 5236 233 5276
rect 253 5236 265 5276
rect 287 5236 299 5276
rect 307 5196 319 5276
rect 337 5236 349 5276
rect 357 5236 369 5276
rect 377 5236 389 5276
rect 431 5196 443 5276
rect 451 5196 463 5276
rect 471 5208 483 5276
rect 491 5204 503 5276
rect 531 5236 543 5276
rect 551 5236 563 5276
rect 571 5236 583 5276
rect 601 5196 613 5276
rect 621 5236 633 5276
rect 655 5236 667 5276
rect 687 5236 699 5276
rect 707 5236 719 5276
rect 733 5236 745 5276
rect 761 5256 773 5276
rect 791 5256 803 5276
rect 811 5196 823 5276
rect 837 5236 849 5276
rect 857 5236 869 5276
rect 877 5236 889 5276
rect 936 5236 948 5276
rect 958 5196 970 5276
rect 986 5196 998 5276
rect 1036 5236 1048 5276
rect 1058 5196 1070 5276
rect 1086 5196 1098 5276
rect 1127 5196 1139 5276
rect 1147 5196 1159 5276
rect 1171 5236 1183 5276
rect 1191 5236 1203 5276
rect 1217 5196 1229 5276
rect 1237 5256 1249 5276
rect 1267 5256 1279 5276
rect 1295 5236 1307 5276
rect 1321 5236 1333 5276
rect 1341 5236 1353 5276
rect 1373 5236 1385 5276
rect 1407 5236 1419 5276
rect 1427 5196 1439 5276
rect 1471 5236 1483 5276
rect 1491 5236 1503 5276
rect 1511 5236 1523 5276
rect 1537 5236 1549 5276
rect 1557 5236 1569 5276
rect 1577 5236 1589 5276
rect 1617 5196 1629 5276
rect 1637 5256 1649 5276
rect 1667 5256 1679 5276
rect 1695 5236 1707 5276
rect 1721 5236 1733 5276
rect 1741 5236 1753 5276
rect 1773 5236 1785 5276
rect 1807 5236 1819 5276
rect 1827 5196 1839 5276
rect 1871 5196 1883 5276
rect 1891 5196 1903 5264
rect 1911 5198 1923 5276
rect 1931 5210 1943 5276
rect 1951 5198 1963 5276
rect 1977 5236 1989 5276
rect 1997 5236 2009 5276
rect 2047 5196 2059 5276
rect 2067 5196 2079 5276
rect 2091 5236 2103 5276
rect 2111 5236 2123 5276
rect 2137 5236 2149 5276
rect 2157 5236 2169 5276
rect 2177 5236 2189 5276
rect 2241 5197 2253 5276
rect 2261 5197 2273 5276
rect 2291 5196 2303 5276
rect 2331 5236 2343 5276
rect 2351 5236 2363 5276
rect 2371 5236 2383 5276
rect 2411 5236 2423 5276
rect 2431 5240 2443 5276
rect 2451 5236 2463 5276
rect 2471 5236 2483 5276
rect 2523 5196 2535 5276
rect 2551 5196 2563 5276
rect 2577 5236 2589 5276
rect 2597 5236 2609 5276
rect 2647 5196 2659 5276
rect 2667 5196 2679 5276
rect 2691 5236 2703 5276
rect 2711 5236 2723 5276
rect 2737 5196 2749 5276
rect 2765 5196 2777 5276
rect 2831 5236 2843 5276
rect 2851 5236 2863 5276
rect 2871 5236 2883 5276
rect 2911 5236 2923 5276
rect 2931 5236 2943 5276
rect 2951 5236 2963 5276
rect 2977 5196 2989 5276
rect 3007 5197 3019 5276
rect 3027 5197 3039 5276
rect 3087 5196 3099 5276
rect 3107 5196 3119 5276
rect 3131 5236 3143 5276
rect 3151 5236 3163 5276
rect 3177 5236 3189 5276
rect 3197 5236 3209 5276
rect 3217 5236 3229 5276
rect 3271 5236 3283 5276
rect 3291 5240 3303 5276
rect 3311 5236 3323 5276
rect 3331 5236 3343 5276
rect 3371 5236 3383 5276
rect 3391 5236 3403 5276
rect 3431 5196 3443 5276
rect 3451 5196 3463 5276
rect 3471 5208 3483 5276
rect 3491 5204 3503 5276
rect 3543 5196 3555 5276
rect 3571 5196 3583 5276
rect 3602 5196 3614 5276
rect 3630 5196 3642 5276
rect 3652 5236 3664 5276
rect 3716 5236 3728 5276
rect 3738 5196 3750 5276
rect 3766 5196 3778 5276
rect 3797 5196 3809 5276
rect 3825 5196 3837 5276
rect 3877 5236 3889 5276
rect 3897 5236 3909 5276
rect 3917 5236 3929 5276
rect 3971 5236 3983 5276
rect 3991 5236 4003 5276
rect 4011 5236 4023 5276
rect 4042 5196 4054 5276
rect 4070 5196 4082 5276
rect 4092 5236 4104 5276
rect 4151 5236 4163 5276
rect 4171 5236 4183 5276
rect 4191 5236 4203 5276
rect 4227 5196 4239 5276
rect 4247 5196 4259 5276
rect 4271 5236 4283 5276
rect 4291 5236 4303 5276
rect 4331 5236 4343 5276
rect 4351 5236 4363 5276
rect 4371 5236 4383 5276
rect 4416 5236 4428 5276
rect 4438 5196 4450 5276
rect 4466 5196 4478 5276
rect 4516 5236 4528 5276
rect 4538 5196 4550 5276
rect 4566 5196 4578 5276
rect 4597 5236 4609 5276
rect 4617 5236 4629 5276
rect 4637 5236 4649 5276
rect 4677 5236 4689 5276
rect 4697 5236 4709 5276
rect 4717 5236 4729 5276
rect 4757 5236 4769 5276
rect 4777 5236 4789 5276
rect 4831 5236 4843 5276
rect 4851 5240 4863 5276
rect 4871 5236 4883 5276
rect 4891 5236 4903 5276
rect 4922 5196 4934 5276
rect 4950 5196 4962 5276
rect 4972 5236 4984 5276
rect 5017 5196 5029 5276
rect 5037 5196 5049 5276
rect 5077 5236 5089 5276
rect 5097 5236 5109 5276
rect 5117 5236 5129 5276
rect 5157 5196 5169 5274
rect 5177 5196 5189 5276
rect 5197 5196 5209 5276
rect 5237 5236 5249 5276
rect 5257 5236 5269 5276
rect 5277 5236 5289 5276
rect 5322 5196 5334 5276
rect 5350 5196 5362 5276
rect 5372 5236 5384 5276
rect 5417 5236 5429 5276
rect 5437 5236 5449 5276
rect 5457 5240 5469 5276
rect 5477 5236 5489 5276
rect 5517 5236 5529 5276
rect 5537 5236 5549 5276
rect 5557 5240 5569 5276
rect 5577 5236 5589 5276
rect 5617 5236 5629 5276
rect 5637 5236 5649 5276
rect 5677 5236 5689 5276
rect 5697 5236 5709 5276
rect 5717 5240 5729 5276
rect 5737 5236 5749 5276
rect 5782 5196 5794 5276
rect 5810 5196 5822 5276
rect 5832 5236 5844 5276
rect 5891 5236 5903 5276
rect 5911 5236 5923 5276
rect 5931 5236 5943 5276
rect 5957 5236 5969 5276
rect 5977 5236 5989 5276
rect 5997 5240 6009 5276
rect 6017 5236 6029 5276
rect 6057 5236 6069 5276
rect 6077 5236 6089 5276
rect 6097 5236 6109 5276
rect 6151 5196 6163 5276
rect 6171 5196 6183 5276
rect 6191 5208 6203 5276
rect 6211 5204 6223 5276
rect 6251 5236 6263 5276
rect 6271 5236 6283 5276
rect 6311 5236 6323 5276
rect 6331 5240 6343 5276
rect 6351 5236 6363 5276
rect 6371 5236 6383 5276
rect 6411 5236 6423 5276
rect 6431 5240 6443 5276
rect 6451 5236 6463 5276
rect 6471 5236 6483 5276
rect 6497 5236 6509 5276
rect 6517 5236 6529 5276
rect 6571 5236 6583 5276
rect 6591 5240 6603 5276
rect 6611 5236 6623 5276
rect 6631 5236 6643 5276
rect 6657 5236 6669 5276
rect 6677 5236 6689 5276
rect 6697 5236 6709 5276
rect 29 4824 41 4904
rect 49 4824 61 4904
rect 71 4824 83 4864
rect 109 4824 121 4904
rect 129 4824 141 4904
rect 151 4824 163 4864
rect 191 4824 203 4864
rect 211 4824 223 4864
rect 231 4824 243 4864
rect 257 4824 269 4904
rect 277 4824 289 4844
rect 307 4824 319 4844
rect 335 4824 347 4864
rect 361 4824 373 4864
rect 381 4824 393 4864
rect 413 4824 425 4864
rect 447 4824 459 4864
rect 467 4824 479 4904
rect 511 4824 523 4904
rect 531 4824 543 4904
rect 551 4824 563 4892
rect 571 4824 583 4896
rect 611 4824 623 4864
rect 631 4824 643 4864
rect 651 4824 663 4864
rect 677 4824 689 4864
rect 697 4824 709 4864
rect 717 4824 729 4864
rect 771 4824 783 4864
rect 791 4824 803 4864
rect 811 4824 823 4864
rect 837 4824 849 4904
rect 857 4824 869 4844
rect 887 4824 899 4844
rect 915 4824 927 4864
rect 941 4824 953 4864
rect 961 4824 973 4864
rect 993 4824 1005 4864
rect 1027 4824 1039 4864
rect 1047 4824 1059 4904
rect 1089 4824 1101 4904
rect 1109 4824 1121 4904
rect 1131 4824 1143 4864
rect 1171 4824 1183 4904
rect 1191 4824 1203 4904
rect 1211 4824 1223 4892
rect 1231 4824 1243 4896
rect 1271 4824 1283 4864
rect 1291 4824 1303 4864
rect 1311 4824 1323 4864
rect 1349 4824 1361 4904
rect 1369 4824 1381 4904
rect 1391 4824 1403 4864
rect 1417 4824 1429 4864
rect 1437 4824 1449 4864
rect 1457 4824 1469 4864
rect 1511 4824 1523 4864
rect 1531 4824 1543 4864
rect 1551 4824 1563 4864
rect 1596 4824 1608 4864
rect 1618 4824 1630 4904
rect 1646 4824 1658 4904
rect 1691 4824 1703 4864
rect 1711 4824 1723 4864
rect 1731 4824 1743 4864
rect 1776 4824 1788 4864
rect 1798 4824 1810 4904
rect 1826 4824 1838 4904
rect 1857 4824 1869 4864
rect 1877 4824 1889 4864
rect 1897 4824 1909 4864
rect 1956 4824 1968 4864
rect 1978 4824 1990 4904
rect 2006 4824 2018 4904
rect 2056 4824 2068 4864
rect 2078 4824 2090 4904
rect 2106 4824 2118 4904
rect 2147 4824 2159 4904
rect 2167 4824 2179 4904
rect 2191 4824 2203 4864
rect 2211 4824 2223 4864
rect 2237 4824 2249 4864
rect 2257 4824 2269 4864
rect 2323 4824 2335 4904
rect 2351 4824 2363 4904
rect 2401 4824 2413 4903
rect 2421 4824 2433 4903
rect 2451 4824 2463 4904
rect 2491 4824 2503 4864
rect 2511 4824 2523 4864
rect 2531 4824 2543 4864
rect 2576 4824 2588 4864
rect 2598 4824 2610 4904
rect 2626 4824 2638 4904
rect 2676 4824 2688 4864
rect 2698 4824 2710 4904
rect 2726 4824 2738 4904
rect 2771 4824 2783 4864
rect 2791 4824 2803 4864
rect 2822 4824 2834 4904
rect 2850 4824 2862 4904
rect 2872 4824 2884 4864
rect 2936 4824 2948 4864
rect 2958 4824 2970 4904
rect 2986 4824 2998 4904
rect 3036 4824 3048 4864
rect 3058 4824 3070 4904
rect 3086 4824 3098 4904
rect 3143 4824 3155 4904
rect 3171 4824 3183 4904
rect 3211 4824 3223 4904
rect 3231 4824 3243 4904
rect 3271 4824 3283 4864
rect 3291 4824 3303 4864
rect 3311 4824 3323 4864
rect 3356 4824 3368 4864
rect 3378 4824 3390 4904
rect 3406 4824 3418 4904
rect 3441 4824 3453 4904
rect 3461 4824 3473 4864
rect 3495 4824 3507 4864
rect 3527 4824 3539 4864
rect 3547 4824 3559 4864
rect 3573 4824 3585 4864
rect 3601 4824 3613 4844
rect 3631 4824 3643 4844
rect 3651 4824 3663 4904
rect 3682 4824 3694 4904
rect 3710 4824 3722 4904
rect 3732 4824 3744 4864
rect 3791 4824 3803 4904
rect 3811 4824 3823 4904
rect 3831 4824 3843 4892
rect 3851 4824 3863 4896
rect 3891 4824 3903 4864
rect 3911 4824 3923 4860
rect 3931 4824 3943 4864
rect 3951 4824 3963 4864
rect 3991 4824 4003 4904
rect 4011 4824 4023 4904
rect 4031 4824 4043 4892
rect 4051 4824 4063 4896
rect 4091 4824 4103 4904
rect 4111 4824 4123 4904
rect 4147 4824 4159 4904
rect 4167 4824 4179 4904
rect 4191 4824 4203 4864
rect 4211 4824 4223 4864
rect 4251 4824 4263 4864
rect 4271 4824 4283 4864
rect 4291 4824 4303 4864
rect 4317 4824 4329 4864
rect 4337 4824 4349 4864
rect 4361 4824 4373 4904
rect 4381 4824 4393 4904
rect 4436 4824 4448 4864
rect 4458 4824 4470 4904
rect 4486 4824 4498 4904
rect 4517 4824 4529 4864
rect 4537 4824 4549 4864
rect 4557 4824 4569 4860
rect 4577 4824 4589 4864
rect 4622 4824 4634 4904
rect 4650 4824 4662 4904
rect 4672 4824 4684 4864
rect 4731 4824 4743 4864
rect 4751 4824 4763 4864
rect 4771 4824 4783 4864
rect 4807 4824 4819 4904
rect 4827 4824 4839 4904
rect 4851 4824 4863 4864
rect 4871 4824 4883 4864
rect 4911 4824 4923 4864
rect 4931 4824 4943 4864
rect 4951 4824 4963 4864
rect 4977 4824 4989 4864
rect 4997 4824 5009 4864
rect 5017 4824 5029 4864
rect 5057 4824 5069 4864
rect 5077 4824 5089 4864
rect 5101 4824 5113 4904
rect 5121 4824 5133 4904
rect 5171 4824 5183 4864
rect 5191 4824 5203 4864
rect 5211 4824 5223 4864
rect 5247 4824 5259 4904
rect 5267 4824 5279 4904
rect 5291 4824 5303 4864
rect 5311 4824 5323 4864
rect 5337 4824 5349 4864
rect 5357 4824 5369 4864
rect 5381 4824 5393 4904
rect 5401 4824 5413 4904
rect 5451 4824 5463 4904
rect 5471 4836 5483 4904
rect 5491 4824 5503 4902
rect 5511 4824 5523 4890
rect 5531 4824 5543 4902
rect 5571 4824 5583 4864
rect 5591 4824 5603 4864
rect 5611 4824 5623 4864
rect 5637 4824 5649 4864
rect 5657 4824 5669 4864
rect 5677 4824 5689 4860
rect 5697 4824 5709 4864
rect 5751 4824 5763 4904
rect 5771 4824 5783 4904
rect 5791 4824 5803 4892
rect 5811 4824 5823 4896
rect 5851 4824 5863 4864
rect 5871 4824 5883 4860
rect 5891 4824 5903 4864
rect 5911 4824 5923 4864
rect 5951 4824 5963 4864
rect 5971 4824 5983 4864
rect 5991 4824 6003 4864
rect 6017 4824 6029 4902
rect 6037 4824 6049 4890
rect 6057 4824 6069 4902
rect 6077 4836 6089 4904
rect 6097 4824 6109 4904
rect 6151 4824 6163 4864
rect 6171 4824 6183 4860
rect 6191 4824 6203 4864
rect 6211 4824 6223 4864
rect 6242 4824 6254 4904
rect 6270 4824 6282 4904
rect 6292 4824 6304 4864
rect 6351 4824 6363 4864
rect 6371 4824 6383 4860
rect 6391 4824 6403 4864
rect 6411 4824 6423 4864
rect 6451 4824 6463 4864
rect 6471 4824 6483 4860
rect 6491 4824 6503 4864
rect 6511 4824 6523 4864
rect 6537 4824 6549 4864
rect 6557 4824 6569 4864
rect 6577 4824 6589 4864
rect 6631 4824 6643 4864
rect 6651 4824 6663 4864
rect 17 4716 29 4796
rect 37 4716 49 4796
rect 57 4716 69 4796
rect 77 4716 89 4796
rect 97 4716 109 4796
rect 117 4716 129 4796
rect 137 4716 149 4796
rect 157 4716 169 4796
rect 177 4716 189 4796
rect 243 4716 255 4796
rect 271 4716 283 4796
rect 311 4756 323 4796
rect 331 4756 343 4796
rect 371 4716 383 4796
rect 391 4716 403 4796
rect 411 4728 423 4796
rect 431 4724 443 4796
rect 471 4756 483 4796
rect 491 4756 503 4796
rect 543 4716 555 4796
rect 571 4716 583 4796
rect 607 4716 619 4796
rect 627 4716 639 4796
rect 651 4756 663 4796
rect 671 4756 683 4796
rect 697 4716 709 4796
rect 725 4716 737 4796
rect 789 4716 801 4796
rect 809 4716 821 4796
rect 831 4756 843 4796
rect 871 4756 883 4796
rect 891 4756 903 4796
rect 911 4756 923 4796
rect 937 4716 949 4796
rect 957 4776 969 4796
rect 987 4776 999 4796
rect 1015 4756 1027 4796
rect 1041 4756 1053 4796
rect 1061 4756 1073 4796
rect 1093 4756 1105 4796
rect 1127 4756 1139 4796
rect 1147 4716 1159 4796
rect 1196 4756 1208 4796
rect 1218 4716 1230 4796
rect 1246 4716 1258 4796
rect 1291 4756 1303 4796
rect 1311 4756 1323 4796
rect 1331 4756 1343 4796
rect 1357 4756 1369 4796
rect 1377 4756 1389 4796
rect 1397 4756 1409 4796
rect 1456 4756 1468 4796
rect 1478 4716 1490 4796
rect 1506 4716 1518 4796
rect 1537 4716 1549 4796
rect 1565 4716 1577 4796
rect 1617 4716 1629 4796
rect 1645 4716 1657 4796
rect 1697 4756 1709 4796
rect 1717 4756 1729 4796
rect 1757 4716 1769 4796
rect 1785 4716 1797 4796
rect 1842 4716 1854 4796
rect 1870 4716 1882 4796
rect 1892 4756 1904 4796
rect 1937 4716 1949 4796
rect 1957 4776 1969 4796
rect 1987 4776 1999 4796
rect 2015 4756 2027 4796
rect 2041 4756 2053 4796
rect 2061 4756 2073 4796
rect 2093 4756 2105 4796
rect 2127 4756 2139 4796
rect 2147 4716 2159 4796
rect 2191 4756 2203 4796
rect 2211 4756 2223 4796
rect 2231 4756 2243 4796
rect 2281 4717 2293 4796
rect 2301 4717 2313 4796
rect 2331 4716 2343 4796
rect 2357 4756 2369 4796
rect 2377 4756 2389 4796
rect 2397 4756 2409 4796
rect 2437 4716 2449 4796
rect 2465 4716 2477 4796
rect 2517 4724 2529 4796
rect 2537 4728 2549 4796
rect 2557 4716 2569 4796
rect 2577 4716 2589 4796
rect 2631 4756 2643 4796
rect 2651 4756 2663 4796
rect 2677 4716 2689 4796
rect 2697 4776 2709 4796
rect 2727 4776 2739 4796
rect 2755 4756 2767 4796
rect 2781 4756 2793 4796
rect 2801 4756 2813 4796
rect 2833 4756 2845 4796
rect 2867 4756 2879 4796
rect 2887 4716 2899 4796
rect 2922 4716 2934 4796
rect 2950 4716 2962 4796
rect 2972 4756 2984 4796
rect 3017 4716 3029 4796
rect 3037 4776 3049 4796
rect 3067 4776 3079 4796
rect 3095 4756 3107 4796
rect 3121 4756 3133 4796
rect 3141 4756 3153 4796
rect 3173 4756 3185 4796
rect 3207 4756 3219 4796
rect 3227 4716 3239 4796
rect 3257 4716 3269 4796
rect 3277 4776 3289 4796
rect 3307 4776 3319 4796
rect 3335 4756 3347 4796
rect 3361 4756 3373 4796
rect 3381 4756 3393 4796
rect 3413 4756 3425 4796
rect 3447 4756 3459 4796
rect 3467 4716 3479 4796
rect 3516 4756 3528 4796
rect 3538 4716 3550 4796
rect 3566 4716 3578 4796
rect 3611 4716 3623 4796
rect 3631 4716 3643 4796
rect 3671 4756 3683 4796
rect 3691 4756 3703 4796
rect 3711 4756 3723 4796
rect 3756 4756 3768 4796
rect 3778 4716 3790 4796
rect 3806 4716 3818 4796
rect 3841 4716 3853 4796
rect 3861 4756 3873 4796
rect 3895 4756 3907 4796
rect 3927 4756 3939 4796
rect 3947 4756 3959 4796
rect 3973 4756 3985 4796
rect 4001 4776 4013 4796
rect 4031 4776 4043 4796
rect 4051 4716 4063 4796
rect 4091 4716 4103 4796
rect 4111 4716 4123 4796
rect 4151 4756 4163 4796
rect 4171 4756 4183 4796
rect 4191 4756 4203 4796
rect 4217 4716 4229 4796
rect 4237 4776 4249 4796
rect 4267 4776 4279 4796
rect 4295 4756 4307 4796
rect 4321 4756 4333 4796
rect 4341 4756 4353 4796
rect 4373 4756 4385 4796
rect 4407 4756 4419 4796
rect 4427 4716 4439 4796
rect 4471 4756 4483 4796
rect 4491 4760 4503 4796
rect 4511 4756 4523 4796
rect 4531 4756 4543 4796
rect 4557 4756 4569 4796
rect 4577 4756 4589 4796
rect 4617 4716 4629 4796
rect 4637 4716 4649 4796
rect 4691 4756 4703 4796
rect 4711 4756 4723 4796
rect 4742 4716 4754 4796
rect 4770 4716 4782 4796
rect 4792 4756 4804 4796
rect 4837 4716 4849 4796
rect 4865 4716 4877 4796
rect 4917 4756 4929 4796
rect 4937 4756 4949 4796
rect 4957 4756 4969 4796
rect 4997 4756 5009 4796
rect 5017 4756 5029 4796
rect 5037 4756 5049 4796
rect 5091 4756 5103 4796
rect 5111 4756 5123 4796
rect 5131 4756 5143 4796
rect 5162 4716 5174 4796
rect 5190 4716 5202 4796
rect 5212 4756 5224 4796
rect 5281 4716 5293 4796
rect 5311 4716 5333 4796
rect 5351 4716 5363 4796
rect 5377 4756 5389 4796
rect 5397 4756 5409 4796
rect 5417 4756 5429 4796
rect 5471 4756 5483 4796
rect 5491 4756 5503 4796
rect 5511 4756 5523 4796
rect 5537 4756 5549 4796
rect 5557 4756 5569 4796
rect 5577 4760 5589 4796
rect 5597 4756 5609 4796
rect 5651 4756 5663 4796
rect 5671 4756 5683 4796
rect 5691 4756 5703 4796
rect 5717 4756 5729 4796
rect 5737 4756 5749 4796
rect 5757 4760 5769 4796
rect 5777 4756 5789 4796
rect 5831 4756 5843 4796
rect 5851 4756 5863 4796
rect 5877 4756 5889 4796
rect 5897 4756 5909 4796
rect 5917 4760 5929 4796
rect 5937 4756 5949 4796
rect 5987 4716 5999 4796
rect 6007 4716 6019 4796
rect 6031 4756 6043 4796
rect 6051 4756 6063 4796
rect 6082 4716 6094 4796
rect 6110 4716 6122 4796
rect 6132 4756 6144 4796
rect 6191 4756 6203 4796
rect 6211 4756 6223 4796
rect 6231 4756 6243 4796
rect 6257 4724 6269 4796
rect 6277 4728 6289 4796
rect 6297 4716 6309 4796
rect 6317 4716 6329 4796
rect 6357 4756 6369 4796
rect 6377 4756 6389 4796
rect 6397 4760 6409 4796
rect 6417 4756 6429 4796
rect 6467 4716 6479 4796
rect 6487 4716 6499 4796
rect 6511 4756 6523 4796
rect 6531 4756 6543 4796
rect 6571 4756 6583 4796
rect 6591 4760 6603 4796
rect 6611 4756 6623 4796
rect 6631 4756 6643 4796
rect 31 4344 43 4384
rect 51 4344 63 4384
rect 103 4344 115 4424
rect 131 4344 143 4424
rect 171 4344 183 4384
rect 191 4344 203 4384
rect 222 4344 234 4424
rect 250 4344 262 4424
rect 272 4344 284 4384
rect 343 4344 355 4424
rect 371 4344 383 4424
rect 402 4344 414 4424
rect 430 4344 442 4424
rect 452 4344 464 4384
rect 497 4344 509 4424
rect 527 4344 539 4423
rect 547 4344 559 4423
rect 597 4344 609 4416
rect 617 4344 629 4412
rect 637 4344 649 4424
rect 657 4344 669 4424
rect 711 4344 723 4384
rect 731 4344 743 4384
rect 757 4344 769 4424
rect 785 4344 797 4424
rect 837 4344 849 4384
rect 857 4344 869 4384
rect 897 4344 909 4424
rect 925 4344 937 4424
rect 977 4344 989 4384
rect 997 4344 1009 4384
rect 1037 4344 1049 4424
rect 1057 4344 1069 4424
rect 1077 4344 1089 4424
rect 1097 4344 1109 4424
rect 1117 4344 1129 4424
rect 1137 4344 1149 4424
rect 1157 4344 1169 4424
rect 1177 4344 1189 4424
rect 1197 4344 1209 4424
rect 1237 4344 1249 4384
rect 1259 4344 1271 4424
rect 1279 4344 1291 4424
rect 1331 4344 1343 4384
rect 1351 4344 1363 4384
rect 1403 4344 1415 4424
rect 1431 4344 1443 4424
rect 1471 4344 1483 4384
rect 1491 4344 1503 4384
rect 1511 4344 1523 4384
rect 1537 4344 1549 4384
rect 1557 4344 1569 4384
rect 1577 4344 1589 4384
rect 1631 4344 1643 4424
rect 1651 4344 1663 4424
rect 1671 4344 1683 4424
rect 1691 4344 1703 4424
rect 1711 4344 1723 4424
rect 1741 4344 1753 4424
rect 1761 4344 1773 4384
rect 1795 4344 1807 4384
rect 1827 4344 1839 4384
rect 1847 4344 1859 4384
rect 1873 4344 1885 4384
rect 1901 4344 1913 4364
rect 1931 4344 1943 4364
rect 1951 4344 1963 4424
rect 1977 4344 1989 4384
rect 1997 4344 2009 4384
rect 2017 4344 2029 4384
rect 2057 4344 2069 4424
rect 2077 4344 2089 4364
rect 2107 4344 2119 4364
rect 2135 4344 2147 4384
rect 2161 4344 2173 4384
rect 2181 4344 2193 4384
rect 2213 4344 2225 4384
rect 2247 4344 2259 4384
rect 2267 4344 2279 4424
rect 2297 4344 2309 4384
rect 2317 4344 2329 4384
rect 2357 4344 2369 4424
rect 2385 4344 2397 4424
rect 2437 4344 2449 4424
rect 2465 4344 2477 4424
rect 2517 4344 2529 4384
rect 2537 4344 2549 4384
rect 2577 4344 2589 4424
rect 2597 4344 2609 4364
rect 2627 4344 2639 4364
rect 2655 4344 2667 4384
rect 2681 4344 2693 4384
rect 2701 4344 2713 4384
rect 2733 4344 2745 4384
rect 2767 4344 2779 4384
rect 2787 4344 2799 4424
rect 2822 4344 2834 4424
rect 2850 4344 2862 4424
rect 2872 4344 2884 4384
rect 2917 4344 2929 4384
rect 2937 4344 2949 4384
rect 2957 4344 2969 4384
rect 3011 4344 3023 4384
rect 3031 4344 3043 4384
rect 3062 4344 3074 4424
rect 3090 4344 3102 4424
rect 3112 4344 3124 4384
rect 3157 4344 3169 4424
rect 3177 4344 3189 4364
rect 3207 4344 3219 4364
rect 3235 4344 3247 4384
rect 3261 4344 3273 4384
rect 3281 4344 3293 4384
rect 3313 4344 3325 4384
rect 3347 4344 3359 4384
rect 3367 4344 3379 4424
rect 3402 4344 3414 4424
rect 3430 4344 3442 4424
rect 3452 4344 3464 4384
rect 3516 4344 3528 4384
rect 3538 4344 3550 4424
rect 3566 4344 3578 4424
rect 3601 4344 3613 4424
rect 3621 4344 3633 4384
rect 3655 4344 3667 4384
rect 3687 4344 3699 4384
rect 3707 4344 3719 4384
rect 3733 4344 3745 4384
rect 3761 4344 3773 4364
rect 3791 4344 3803 4364
rect 3811 4344 3823 4424
rect 3842 4344 3854 4424
rect 3870 4344 3882 4424
rect 3892 4344 3904 4384
rect 3941 4344 3953 4424
rect 3961 4344 3973 4384
rect 3995 4344 4007 4384
rect 4027 4344 4039 4384
rect 4047 4344 4059 4384
rect 4073 4344 4085 4384
rect 4101 4344 4113 4364
rect 4131 4344 4143 4364
rect 4151 4344 4163 4424
rect 4191 4344 4203 4384
rect 4211 4344 4223 4380
rect 4231 4344 4243 4384
rect 4251 4344 4263 4384
rect 4282 4344 4294 4424
rect 4310 4344 4322 4424
rect 4332 4344 4344 4384
rect 4403 4344 4415 4424
rect 4431 4344 4443 4424
rect 4471 4344 4483 4424
rect 4491 4344 4503 4424
rect 4511 4344 4523 4412
rect 4531 4344 4543 4416
rect 4557 4344 4569 4384
rect 4577 4344 4589 4384
rect 4597 4344 4609 4380
rect 4617 4344 4629 4384
rect 4671 4344 4683 4384
rect 4691 4344 4703 4384
rect 4722 4344 4734 4424
rect 4750 4344 4762 4424
rect 4772 4344 4784 4384
rect 4841 4344 4853 4423
rect 4861 4344 4873 4423
rect 4891 4344 4903 4424
rect 4931 4344 4943 4384
rect 4951 4344 4963 4384
rect 4971 4344 4983 4384
rect 5011 4344 5023 4384
rect 5031 4344 5043 4380
rect 5051 4344 5063 4384
rect 5071 4344 5083 4384
rect 5102 4344 5114 4424
rect 5130 4344 5142 4424
rect 5152 4344 5164 4384
rect 5221 4344 5233 4423
rect 5241 4344 5253 4423
rect 5271 4344 5283 4424
rect 5302 4344 5314 4424
rect 5330 4344 5342 4424
rect 5352 4344 5364 4384
rect 5397 4344 5409 4384
rect 5417 4344 5429 4384
rect 5471 4344 5483 4384
rect 5491 4344 5503 4380
rect 5511 4344 5523 4384
rect 5531 4344 5543 4384
rect 5557 4344 5569 4384
rect 5577 4344 5589 4384
rect 5597 4344 5609 4384
rect 5642 4344 5654 4424
rect 5670 4344 5682 4424
rect 5692 4344 5704 4384
rect 5751 4344 5763 4384
rect 5771 4344 5783 4384
rect 5791 4344 5803 4384
rect 5831 4344 5843 4384
rect 5851 4344 5863 4380
rect 5871 4344 5883 4384
rect 5891 4344 5903 4384
rect 5936 4344 5948 4384
rect 5958 4344 5970 4424
rect 5986 4344 5998 4424
rect 6017 4344 6029 4384
rect 6037 4344 6049 4384
rect 6091 4344 6103 4384
rect 6111 4344 6123 4384
rect 6137 4344 6149 4384
rect 6157 4344 6169 4384
rect 6177 4344 6189 4380
rect 6197 4344 6209 4384
rect 6256 4344 6268 4384
rect 6278 4344 6290 4424
rect 6306 4344 6318 4424
rect 6337 4344 6349 4384
rect 6357 4344 6369 4384
rect 6377 4344 6389 4380
rect 6397 4344 6409 4384
rect 6437 4344 6449 4384
rect 6457 4344 6469 4384
rect 6477 4344 6489 4380
rect 6497 4344 6509 4384
rect 6542 4344 6554 4424
rect 6570 4344 6582 4424
rect 6592 4344 6604 4384
rect 6637 4344 6649 4384
rect 6657 4344 6669 4384
rect 29 4236 41 4316
rect 49 4236 61 4316
rect 71 4276 83 4316
rect 116 4276 128 4316
rect 138 4236 150 4316
rect 166 4236 178 4316
rect 202 4236 214 4316
rect 230 4236 242 4316
rect 252 4276 264 4316
rect 301 4236 313 4316
rect 321 4276 333 4316
rect 355 4276 367 4316
rect 387 4276 399 4316
rect 407 4276 419 4316
rect 433 4276 445 4316
rect 461 4296 473 4316
rect 491 4296 503 4316
rect 511 4236 523 4316
rect 537 4276 549 4316
rect 557 4276 569 4316
rect 577 4276 589 4316
rect 631 4236 643 4316
rect 651 4236 663 4304
rect 671 4238 683 4316
rect 691 4250 703 4316
rect 711 4238 723 4316
rect 751 4276 763 4316
rect 771 4276 783 4316
rect 797 4236 809 4316
rect 817 4296 829 4316
rect 847 4296 859 4316
rect 875 4276 887 4316
rect 901 4276 913 4316
rect 921 4276 933 4316
rect 953 4276 965 4316
rect 987 4276 999 4316
rect 1007 4236 1019 4316
rect 1037 4276 1049 4316
rect 1057 4276 1069 4316
rect 1077 4276 1089 4316
rect 1117 4236 1129 4316
rect 1137 4296 1149 4316
rect 1167 4296 1179 4316
rect 1195 4276 1207 4316
rect 1221 4276 1233 4316
rect 1241 4276 1253 4316
rect 1273 4276 1285 4316
rect 1307 4276 1319 4316
rect 1327 4236 1339 4316
rect 1357 4276 1369 4316
rect 1377 4276 1389 4316
rect 1397 4276 1409 4316
rect 1437 4276 1449 4316
rect 1457 4276 1469 4316
rect 1516 4276 1528 4316
rect 1538 4236 1550 4316
rect 1566 4236 1578 4316
rect 1611 4236 1623 4316
rect 1631 4236 1643 4316
rect 1651 4248 1663 4316
rect 1671 4244 1683 4316
rect 1711 4276 1723 4316
rect 1731 4276 1743 4316
rect 1751 4276 1763 4316
rect 1777 4276 1789 4316
rect 1797 4276 1809 4316
rect 1817 4276 1829 4316
rect 1857 4236 1869 4316
rect 1877 4296 1889 4316
rect 1907 4296 1919 4316
rect 1935 4276 1947 4316
rect 1961 4276 1973 4316
rect 1981 4276 1993 4316
rect 2013 4276 2025 4316
rect 2047 4276 2059 4316
rect 2067 4236 2079 4316
rect 2097 4276 2109 4316
rect 2117 4276 2129 4316
rect 2137 4276 2149 4316
rect 2196 4276 2208 4316
rect 2218 4236 2230 4316
rect 2246 4236 2258 4316
rect 2281 4236 2293 4316
rect 2301 4276 2313 4316
rect 2335 4276 2347 4316
rect 2367 4276 2379 4316
rect 2387 4276 2399 4316
rect 2413 4276 2425 4316
rect 2441 4296 2453 4316
rect 2471 4296 2483 4316
rect 2491 4236 2503 4316
rect 2543 4236 2555 4316
rect 2571 4236 2583 4316
rect 2597 4276 2609 4316
rect 2617 4276 2629 4316
rect 2662 4236 2674 4316
rect 2690 4236 2702 4316
rect 2712 4276 2724 4316
rect 2757 4276 2769 4316
rect 2777 4276 2789 4316
rect 2797 4276 2809 4316
rect 2856 4276 2868 4316
rect 2878 4236 2890 4316
rect 2906 4236 2918 4316
rect 2937 4276 2949 4316
rect 2957 4276 2969 4316
rect 2997 4236 3009 4316
rect 3025 4236 3037 4316
rect 3091 4276 3103 4316
rect 3111 4276 3123 4316
rect 3137 4236 3149 4316
rect 3157 4296 3169 4316
rect 3187 4296 3199 4316
rect 3215 4276 3227 4316
rect 3241 4276 3253 4316
rect 3261 4276 3273 4316
rect 3293 4276 3305 4316
rect 3327 4276 3339 4316
rect 3347 4236 3359 4316
rect 3377 4236 3389 4316
rect 3407 4236 3429 4316
rect 3447 4236 3459 4316
rect 3497 4276 3509 4316
rect 3517 4276 3529 4316
rect 3537 4276 3549 4316
rect 3577 4236 3589 4316
rect 3597 4236 3609 4316
rect 3617 4236 3629 4316
rect 3637 4236 3649 4316
rect 3657 4236 3669 4316
rect 3677 4236 3689 4316
rect 3697 4236 3709 4316
rect 3717 4236 3729 4316
rect 3737 4236 3749 4316
rect 3777 4276 3789 4316
rect 3797 4276 3809 4316
rect 3817 4276 3829 4316
rect 3857 4276 3869 4316
rect 3877 4276 3889 4316
rect 3897 4276 3909 4316
rect 3951 4276 3963 4316
rect 3971 4276 3983 4316
rect 3991 4276 4003 4316
rect 4017 4276 4029 4316
rect 4037 4276 4049 4316
rect 4096 4276 4108 4316
rect 4118 4236 4130 4316
rect 4146 4236 4158 4316
rect 4182 4236 4194 4316
rect 4210 4236 4222 4316
rect 4232 4276 4244 4316
rect 4281 4236 4293 4316
rect 4301 4276 4313 4316
rect 4335 4276 4347 4316
rect 4367 4276 4379 4316
rect 4387 4276 4399 4316
rect 4413 4276 4425 4316
rect 4441 4296 4453 4316
rect 4471 4296 4483 4316
rect 4491 4236 4503 4316
rect 4536 4276 4548 4316
rect 4558 4236 4570 4316
rect 4586 4236 4598 4316
rect 4621 4236 4633 4316
rect 4641 4276 4653 4316
rect 4675 4276 4687 4316
rect 4707 4276 4719 4316
rect 4727 4276 4739 4316
rect 4753 4276 4765 4316
rect 4781 4296 4793 4316
rect 4811 4296 4823 4316
rect 4831 4236 4843 4316
rect 4871 4236 4883 4316
rect 4891 4236 4903 4316
rect 4931 4236 4943 4316
rect 4951 4236 4963 4316
rect 4971 4248 4983 4316
rect 4991 4244 5003 4316
rect 5017 4276 5029 4316
rect 5037 4276 5049 4316
rect 5057 4280 5069 4316
rect 5077 4276 5089 4316
rect 5131 4276 5143 4316
rect 5151 4276 5163 4316
rect 5182 4236 5194 4316
rect 5210 4236 5222 4316
rect 5232 4276 5244 4316
rect 5281 4236 5293 4316
rect 5301 4276 5313 4316
rect 5335 4276 5347 4316
rect 5367 4276 5379 4316
rect 5387 4276 5399 4316
rect 5413 4276 5425 4316
rect 5441 4296 5453 4316
rect 5471 4296 5483 4316
rect 5491 4236 5503 4316
rect 5517 4276 5529 4316
rect 5537 4276 5549 4316
rect 5557 4276 5569 4316
rect 5597 4276 5609 4316
rect 5617 4276 5629 4316
rect 5662 4236 5674 4316
rect 5690 4236 5702 4316
rect 5712 4276 5724 4316
rect 5767 4236 5779 4316
rect 5787 4236 5799 4316
rect 5811 4276 5823 4316
rect 5831 4276 5843 4316
rect 5857 4276 5869 4316
rect 5877 4276 5889 4316
rect 5897 4280 5909 4316
rect 5917 4276 5929 4316
rect 5971 4236 5983 4316
rect 5991 4236 6003 4316
rect 6022 4236 6034 4316
rect 6050 4236 6062 4316
rect 6072 4276 6084 4316
rect 6117 4276 6129 4316
rect 6139 4236 6151 4316
rect 6159 4236 6171 4316
rect 6197 4276 6209 4316
rect 6217 4276 6229 4316
rect 6237 4276 6249 4316
rect 6287 4236 6299 4316
rect 6307 4236 6319 4316
rect 6331 4276 6343 4316
rect 6351 4276 6363 4316
rect 6377 4276 6389 4316
rect 6397 4276 6409 4316
rect 6417 4276 6429 4316
rect 6457 4276 6469 4316
rect 6477 4276 6489 4316
rect 6531 4236 6543 4316
rect 6551 4236 6563 4316
rect 6571 4248 6583 4316
rect 6591 4244 6603 4316
rect 6617 4276 6629 4316
rect 6637 4276 6649 4316
rect 6657 4280 6669 4316
rect 6677 4276 6689 4316
rect 29 3864 41 3944
rect 49 3864 61 3944
rect 71 3864 83 3904
rect 97 3864 109 3944
rect 117 3864 129 3884
rect 147 3864 159 3884
rect 175 3864 187 3904
rect 201 3864 213 3904
rect 221 3864 233 3904
rect 253 3864 265 3904
rect 287 3864 299 3904
rect 307 3864 319 3944
rect 337 3864 349 3904
rect 357 3864 369 3904
rect 377 3864 389 3904
rect 431 3864 443 3944
rect 451 3864 463 3944
rect 471 3864 483 3932
rect 491 3864 503 3936
rect 531 3864 543 3904
rect 551 3864 563 3904
rect 571 3864 583 3904
rect 611 3864 623 3904
rect 631 3864 643 3904
rect 651 3864 663 3904
rect 689 3864 701 3944
rect 709 3864 721 3944
rect 731 3864 743 3904
rect 757 3864 769 3944
rect 777 3864 789 3884
rect 807 3864 819 3884
rect 835 3864 847 3904
rect 861 3864 873 3904
rect 881 3864 893 3904
rect 913 3864 925 3904
rect 947 3864 959 3904
rect 967 3864 979 3944
rect 1011 3864 1023 3904
rect 1031 3864 1043 3904
rect 1051 3864 1063 3904
rect 1077 3864 1089 3904
rect 1097 3864 1109 3904
rect 1117 3864 1129 3904
rect 1157 3864 1169 3904
rect 1177 3864 1189 3904
rect 1197 3864 1209 3904
rect 1251 3864 1263 3944
rect 1271 3864 1283 3944
rect 1291 3864 1303 3932
rect 1311 3864 1323 3936
rect 1337 3864 1349 3944
rect 1357 3864 1369 3884
rect 1387 3864 1399 3884
rect 1415 3864 1427 3904
rect 1441 3864 1453 3904
rect 1461 3864 1473 3904
rect 1493 3864 1505 3904
rect 1527 3864 1539 3904
rect 1547 3864 1559 3944
rect 1591 3864 1603 3904
rect 1611 3864 1623 3904
rect 1631 3864 1643 3904
rect 1657 3864 1669 3904
rect 1679 3864 1691 3944
rect 1699 3864 1711 3944
rect 1737 3864 1749 3904
rect 1757 3864 1769 3904
rect 1777 3864 1789 3904
rect 1817 3864 1829 3944
rect 1837 3864 1849 3884
rect 1867 3864 1879 3884
rect 1895 3864 1907 3904
rect 1921 3864 1933 3904
rect 1941 3864 1953 3904
rect 1973 3864 1985 3904
rect 2007 3864 2019 3904
rect 2027 3864 2039 3944
rect 2057 3864 2069 3904
rect 2077 3864 2089 3904
rect 2097 3864 2109 3904
rect 2156 3864 2168 3904
rect 2178 3864 2190 3944
rect 2206 3864 2218 3944
rect 2251 3864 2263 3904
rect 2271 3864 2283 3904
rect 2291 3864 2303 3904
rect 2317 3864 2329 3904
rect 2337 3864 2349 3904
rect 2357 3864 2369 3904
rect 2411 3864 2423 3904
rect 2431 3864 2443 3904
rect 2476 3864 2488 3904
rect 2498 3864 2510 3944
rect 2526 3864 2538 3944
rect 2557 3864 2569 3944
rect 2585 3864 2597 3944
rect 2663 3864 2675 3944
rect 2691 3864 2703 3944
rect 2717 3864 2729 3904
rect 2737 3864 2749 3904
rect 2791 3864 2803 3904
rect 2811 3864 2823 3904
rect 2851 3864 2863 3904
rect 2871 3864 2883 3904
rect 2891 3864 2903 3904
rect 2917 3864 2929 3944
rect 2945 3864 2957 3944
rect 3002 3864 3014 3944
rect 3030 3864 3042 3944
rect 3052 3864 3064 3904
rect 3097 3864 3109 3904
rect 3117 3864 3129 3904
rect 3157 3864 3169 3944
rect 3185 3864 3197 3944
rect 3251 3864 3263 3904
rect 3271 3864 3283 3904
rect 3291 3864 3303 3904
rect 3331 3864 3343 3904
rect 3351 3864 3363 3904
rect 3371 3864 3383 3904
rect 3401 3864 3413 3944
rect 3421 3864 3433 3904
rect 3455 3864 3467 3904
rect 3487 3864 3499 3904
rect 3507 3864 3519 3904
rect 3533 3864 3545 3904
rect 3561 3864 3573 3884
rect 3591 3864 3603 3884
rect 3611 3864 3623 3944
rect 3651 3864 3663 3904
rect 3671 3864 3683 3904
rect 3701 3864 3713 3944
rect 3721 3864 3733 3904
rect 3755 3864 3767 3904
rect 3787 3864 3799 3904
rect 3807 3864 3819 3904
rect 3833 3864 3845 3904
rect 3861 3864 3873 3884
rect 3891 3864 3903 3884
rect 3911 3864 3923 3944
rect 3951 3864 3963 3904
rect 3971 3864 3983 3900
rect 3991 3864 4003 3904
rect 4011 3864 4023 3904
rect 4037 3864 4049 3904
rect 4057 3864 4069 3904
rect 4077 3864 4089 3904
rect 4136 3864 4148 3904
rect 4158 3864 4170 3944
rect 4186 3864 4198 3944
rect 4217 3864 4229 3944
rect 4245 3864 4257 3944
rect 4311 3864 4323 3904
rect 4331 3864 4343 3904
rect 4371 3864 4383 3904
rect 4391 3864 4403 3904
rect 4411 3864 4423 3904
rect 4456 3864 4468 3904
rect 4478 3864 4490 3944
rect 4506 3864 4518 3944
rect 4541 3864 4553 3944
rect 4561 3864 4573 3904
rect 4595 3864 4607 3904
rect 4627 3864 4639 3904
rect 4647 3864 4659 3904
rect 4673 3864 4685 3904
rect 4701 3864 4713 3884
rect 4731 3864 4743 3884
rect 4751 3864 4763 3944
rect 4791 3864 4803 3904
rect 4811 3864 4823 3904
rect 4831 3864 4843 3904
rect 4876 3864 4888 3904
rect 4898 3864 4910 3944
rect 4926 3864 4938 3944
rect 4961 3864 4973 3944
rect 4981 3864 4993 3904
rect 5015 3864 5027 3904
rect 5047 3864 5059 3904
rect 5067 3864 5079 3904
rect 5093 3864 5105 3904
rect 5121 3864 5133 3884
rect 5151 3864 5163 3884
rect 5171 3864 5183 3944
rect 5211 3864 5223 3904
rect 5231 3864 5243 3904
rect 5251 3864 5263 3904
rect 5296 3864 5308 3904
rect 5318 3864 5330 3944
rect 5346 3864 5358 3944
rect 5391 3864 5403 3904
rect 5411 3864 5423 3904
rect 5431 3864 5443 3904
rect 5462 3864 5474 3944
rect 5490 3864 5502 3944
rect 5512 3864 5524 3904
rect 5571 3864 5583 3904
rect 5591 3864 5603 3904
rect 5621 3864 5633 3944
rect 5641 3864 5653 3904
rect 5675 3864 5687 3904
rect 5707 3864 5719 3904
rect 5727 3864 5739 3904
rect 5753 3864 5765 3904
rect 5781 3864 5793 3884
rect 5811 3864 5823 3884
rect 5831 3864 5843 3944
rect 5857 3864 5869 3904
rect 5877 3864 5889 3904
rect 5931 3864 5943 3904
rect 5951 3864 5963 3900
rect 5971 3864 5983 3904
rect 5991 3864 6003 3904
rect 6017 3864 6029 3944
rect 6037 3864 6049 3884
rect 6067 3864 6079 3884
rect 6095 3864 6107 3904
rect 6121 3864 6133 3904
rect 6141 3864 6153 3904
rect 6173 3864 6185 3904
rect 6207 3864 6219 3904
rect 6227 3864 6239 3944
rect 6257 3864 6269 3944
rect 6277 3864 6289 3884
rect 6307 3864 6319 3884
rect 6335 3864 6347 3904
rect 6361 3864 6373 3904
rect 6381 3864 6393 3904
rect 6413 3864 6425 3904
rect 6447 3864 6459 3904
rect 6467 3864 6479 3944
rect 6497 3864 6509 3944
rect 6517 3864 6529 3884
rect 6547 3864 6559 3884
rect 6575 3864 6587 3904
rect 6601 3864 6613 3904
rect 6621 3864 6633 3904
rect 6653 3864 6665 3904
rect 6687 3864 6699 3904
rect 6707 3864 6719 3944
rect 29 3756 41 3836
rect 49 3756 61 3836
rect 71 3796 83 3836
rect 109 3756 121 3836
rect 129 3756 141 3836
rect 151 3796 163 3836
rect 191 3796 203 3836
rect 211 3796 223 3836
rect 231 3796 243 3836
rect 257 3756 269 3836
rect 277 3816 289 3836
rect 307 3816 319 3836
rect 335 3796 347 3836
rect 361 3796 373 3836
rect 381 3796 393 3836
rect 413 3796 425 3836
rect 447 3796 459 3836
rect 467 3756 479 3836
rect 511 3756 523 3836
rect 531 3756 543 3836
rect 551 3768 563 3836
rect 571 3764 583 3836
rect 611 3796 623 3836
rect 631 3796 643 3836
rect 651 3796 663 3836
rect 677 3796 689 3836
rect 697 3796 709 3836
rect 717 3796 729 3836
rect 771 3796 783 3836
rect 791 3796 803 3836
rect 811 3796 823 3836
rect 837 3756 849 3836
rect 857 3816 869 3836
rect 887 3816 899 3836
rect 915 3796 927 3836
rect 941 3796 953 3836
rect 961 3796 973 3836
rect 993 3796 1005 3836
rect 1027 3796 1039 3836
rect 1047 3756 1059 3836
rect 1077 3764 1089 3836
rect 1097 3768 1109 3836
rect 1117 3756 1129 3836
rect 1137 3756 1149 3836
rect 1191 3796 1203 3836
rect 1211 3796 1223 3836
rect 1231 3796 1243 3836
rect 1257 3796 1269 3836
rect 1279 3756 1291 3836
rect 1299 3756 1311 3836
rect 1351 3756 1363 3836
rect 1371 3756 1383 3836
rect 1391 3768 1403 3836
rect 1411 3764 1423 3836
rect 1451 3796 1463 3836
rect 1471 3796 1483 3836
rect 1491 3796 1503 3836
rect 1517 3796 1529 3836
rect 1537 3796 1549 3836
rect 1557 3796 1569 3836
rect 1597 3756 1609 3836
rect 1625 3756 1637 3836
rect 1677 3756 1689 3836
rect 1697 3816 1709 3836
rect 1727 3816 1739 3836
rect 1755 3796 1767 3836
rect 1781 3796 1793 3836
rect 1801 3796 1813 3836
rect 1833 3796 1845 3836
rect 1867 3796 1879 3836
rect 1887 3756 1899 3836
rect 1931 3796 1943 3836
rect 1951 3796 1963 3836
rect 1971 3796 1983 3836
rect 1997 3756 2009 3836
rect 2025 3756 2037 3836
rect 2077 3796 2089 3836
rect 2097 3796 2109 3836
rect 2142 3756 2154 3836
rect 2170 3756 2182 3836
rect 2192 3796 2204 3836
rect 2256 3796 2268 3836
rect 2278 3756 2290 3836
rect 2306 3756 2318 3836
rect 2351 3756 2363 3836
rect 2371 3756 2383 3836
rect 2391 3768 2403 3836
rect 2411 3764 2423 3836
rect 2437 3796 2449 3836
rect 2457 3796 2469 3836
rect 2511 3796 2523 3836
rect 2531 3796 2543 3836
rect 2562 3756 2574 3836
rect 2590 3756 2602 3836
rect 2612 3796 2624 3836
rect 2657 3796 2669 3836
rect 2677 3796 2689 3836
rect 2697 3800 2709 3836
rect 2717 3796 2729 3836
rect 2771 3796 2783 3836
rect 2791 3796 2803 3836
rect 2831 3796 2843 3836
rect 2851 3796 2863 3836
rect 2871 3796 2883 3836
rect 2902 3756 2914 3836
rect 2930 3756 2942 3836
rect 2952 3796 2964 3836
rect 3002 3756 3014 3836
rect 3030 3756 3042 3836
rect 3052 3796 3064 3836
rect 3097 3764 3109 3836
rect 3117 3768 3129 3836
rect 3137 3756 3149 3836
rect 3157 3756 3169 3836
rect 3211 3756 3223 3836
rect 3231 3756 3243 3824
rect 3251 3758 3263 3836
rect 3271 3770 3283 3836
rect 3291 3758 3303 3836
rect 3331 3796 3343 3836
rect 3351 3796 3363 3836
rect 3371 3796 3383 3836
rect 3411 3796 3423 3836
rect 3431 3796 3443 3836
rect 3451 3796 3463 3836
rect 3481 3756 3493 3836
rect 3501 3796 3513 3836
rect 3535 3796 3547 3836
rect 3567 3796 3579 3836
rect 3587 3796 3599 3836
rect 3613 3796 3625 3836
rect 3641 3816 3653 3836
rect 3671 3816 3683 3836
rect 3691 3756 3703 3836
rect 3731 3796 3743 3836
rect 3751 3796 3763 3836
rect 3771 3796 3783 3836
rect 3811 3756 3823 3836
rect 3831 3756 3843 3824
rect 3851 3758 3863 3836
rect 3871 3770 3883 3836
rect 3891 3758 3903 3836
rect 3917 3796 3929 3836
rect 3937 3796 3949 3836
rect 3977 3796 3989 3836
rect 3997 3796 4009 3836
rect 4017 3796 4029 3836
rect 4062 3756 4074 3836
rect 4090 3756 4102 3836
rect 4112 3796 4124 3836
rect 4161 3756 4173 3836
rect 4181 3796 4193 3836
rect 4215 3796 4227 3836
rect 4247 3796 4259 3836
rect 4267 3796 4279 3836
rect 4293 3796 4305 3836
rect 4321 3816 4333 3836
rect 4351 3816 4363 3836
rect 4371 3756 4383 3836
rect 4397 3796 4409 3836
rect 4417 3796 4429 3836
rect 4437 3796 4449 3836
rect 4491 3796 4503 3836
rect 4511 3796 4523 3836
rect 4531 3796 4543 3836
rect 4571 3756 4583 3836
rect 4591 3756 4603 3836
rect 4611 3756 4623 3836
rect 4631 3756 4643 3836
rect 4651 3756 4663 3836
rect 4671 3756 4683 3836
rect 4691 3756 4703 3836
rect 4711 3756 4723 3836
rect 4731 3756 4743 3836
rect 4761 3756 4773 3836
rect 4781 3796 4793 3836
rect 4815 3796 4827 3836
rect 4847 3796 4859 3836
rect 4867 3796 4879 3836
rect 4893 3796 4905 3836
rect 4921 3816 4933 3836
rect 4951 3816 4963 3836
rect 4971 3756 4983 3836
rect 5002 3756 5014 3836
rect 5030 3756 5042 3836
rect 5052 3796 5064 3836
rect 5111 3796 5123 3836
rect 5131 3796 5143 3836
rect 5151 3796 5163 3836
rect 5191 3796 5203 3836
rect 5211 3796 5223 3836
rect 5231 3796 5243 3836
rect 5271 3796 5283 3836
rect 5291 3796 5303 3836
rect 5317 3756 5329 3836
rect 5337 3756 5349 3836
rect 5357 3756 5369 3836
rect 5377 3756 5389 3836
rect 5397 3756 5409 3836
rect 5417 3756 5429 3836
rect 5437 3756 5449 3836
rect 5457 3756 5469 3836
rect 5477 3756 5489 3836
rect 5517 3756 5529 3836
rect 5537 3816 5549 3836
rect 5567 3816 5579 3836
rect 5595 3796 5607 3836
rect 5621 3796 5633 3836
rect 5641 3796 5653 3836
rect 5673 3796 5685 3836
rect 5707 3796 5719 3836
rect 5727 3756 5739 3836
rect 5771 3796 5783 3836
rect 5791 3796 5803 3836
rect 5817 3796 5829 3836
rect 5837 3796 5849 3836
rect 5857 3796 5869 3836
rect 5897 3796 5909 3836
rect 5917 3796 5929 3836
rect 5937 3796 5949 3836
rect 5991 3796 6003 3836
rect 6011 3796 6023 3836
rect 6037 3756 6049 3836
rect 6065 3756 6077 3836
rect 6143 3756 6155 3836
rect 6171 3756 6183 3836
rect 6197 3764 6209 3836
rect 6217 3768 6229 3836
rect 6237 3756 6249 3836
rect 6257 3756 6269 3836
rect 6297 3756 6309 3836
rect 6317 3816 6329 3836
rect 6347 3816 6359 3836
rect 6375 3796 6387 3836
rect 6401 3796 6413 3836
rect 6421 3796 6433 3836
rect 6453 3796 6465 3836
rect 6487 3796 6499 3836
rect 6507 3756 6519 3836
rect 6542 3756 6554 3836
rect 6570 3756 6582 3836
rect 6592 3796 6604 3836
rect 6637 3796 6649 3836
rect 6657 3796 6669 3836
rect 6677 3796 6689 3836
rect 29 3384 41 3464
rect 49 3384 61 3464
rect 71 3384 83 3424
rect 97 3384 109 3464
rect 117 3384 129 3404
rect 147 3384 159 3404
rect 175 3384 187 3424
rect 201 3384 213 3424
rect 221 3384 233 3424
rect 253 3384 265 3424
rect 287 3384 299 3424
rect 307 3384 319 3464
rect 337 3384 349 3424
rect 357 3384 369 3424
rect 377 3384 389 3424
rect 417 3384 429 3424
rect 439 3384 451 3464
rect 459 3384 471 3464
rect 511 3384 523 3464
rect 531 3384 543 3464
rect 551 3384 563 3452
rect 571 3384 583 3456
rect 611 3384 623 3424
rect 631 3384 643 3424
rect 651 3384 663 3424
rect 689 3384 701 3464
rect 709 3384 721 3464
rect 731 3384 743 3424
rect 757 3384 769 3424
rect 779 3384 791 3464
rect 799 3384 811 3464
rect 837 3384 849 3424
rect 857 3384 869 3424
rect 877 3384 889 3424
rect 929 3384 941 3464
rect 949 3384 961 3464
rect 971 3384 983 3424
rect 1011 3384 1023 3424
rect 1031 3384 1043 3424
rect 1069 3384 1081 3464
rect 1089 3384 1101 3464
rect 1111 3384 1123 3424
rect 1149 3384 1161 3464
rect 1169 3384 1181 3464
rect 1191 3384 1203 3424
rect 1217 3384 1229 3464
rect 1237 3384 1249 3404
rect 1267 3384 1279 3404
rect 1295 3384 1307 3424
rect 1321 3384 1333 3424
rect 1341 3384 1353 3424
rect 1373 3384 1385 3424
rect 1407 3384 1419 3424
rect 1427 3384 1439 3464
rect 1483 3384 1495 3464
rect 1511 3384 1523 3464
rect 1537 3384 1549 3464
rect 1557 3384 1569 3404
rect 1587 3384 1599 3404
rect 1615 3384 1627 3424
rect 1641 3384 1653 3424
rect 1661 3384 1673 3424
rect 1693 3384 1705 3424
rect 1727 3384 1739 3424
rect 1747 3384 1759 3464
rect 1787 3384 1799 3464
rect 1807 3384 1819 3464
rect 1831 3384 1843 3424
rect 1851 3384 1863 3424
rect 1891 3384 1903 3424
rect 1911 3384 1923 3424
rect 1956 3384 1968 3424
rect 1978 3384 1990 3464
rect 2006 3384 2018 3464
rect 2037 3384 2049 3464
rect 2065 3384 2077 3464
rect 2131 3384 2143 3424
rect 2151 3384 2163 3424
rect 2187 3384 2199 3464
rect 2207 3384 2219 3464
rect 2231 3384 2243 3424
rect 2251 3384 2263 3424
rect 2303 3384 2315 3464
rect 2331 3384 2343 3464
rect 2357 3384 2369 3464
rect 2377 3384 2389 3404
rect 2407 3384 2419 3404
rect 2435 3384 2447 3424
rect 2461 3384 2473 3424
rect 2481 3384 2493 3424
rect 2513 3384 2525 3424
rect 2547 3384 2559 3424
rect 2567 3384 2579 3464
rect 2597 3384 2609 3464
rect 2625 3384 2637 3464
rect 2682 3384 2694 3464
rect 2710 3384 2722 3464
rect 2732 3384 2744 3424
rect 2791 3384 2803 3424
rect 2811 3384 2823 3424
rect 2851 3384 2863 3424
rect 2871 3384 2883 3424
rect 2891 3384 2903 3424
rect 2922 3384 2934 3464
rect 2950 3384 2962 3464
rect 2972 3384 2984 3424
rect 3017 3384 3029 3456
rect 3037 3384 3049 3452
rect 3057 3384 3069 3464
rect 3077 3384 3089 3464
rect 3117 3384 3129 3464
rect 3137 3384 3149 3464
rect 3191 3384 3203 3464
rect 3211 3396 3223 3464
rect 3231 3384 3243 3462
rect 3251 3384 3263 3450
rect 3271 3384 3283 3462
rect 3311 3384 3323 3424
rect 3331 3384 3343 3424
rect 3357 3384 3369 3464
rect 3377 3384 3389 3404
rect 3407 3384 3419 3404
rect 3435 3384 3447 3424
rect 3461 3384 3473 3424
rect 3481 3384 3493 3424
rect 3513 3384 3525 3424
rect 3547 3384 3559 3424
rect 3567 3384 3579 3464
rect 3611 3384 3623 3464
rect 3631 3396 3643 3464
rect 3651 3384 3663 3462
rect 3671 3384 3683 3450
rect 3691 3384 3703 3462
rect 3717 3384 3729 3464
rect 3737 3384 3749 3404
rect 3767 3384 3779 3404
rect 3795 3384 3807 3424
rect 3821 3384 3833 3424
rect 3841 3384 3853 3424
rect 3873 3384 3885 3424
rect 3907 3384 3919 3424
rect 3927 3384 3939 3464
rect 3971 3384 3983 3424
rect 3991 3384 4003 3424
rect 4017 3384 4029 3464
rect 4037 3384 4049 3404
rect 4067 3384 4079 3404
rect 4095 3384 4107 3424
rect 4121 3384 4133 3424
rect 4141 3384 4153 3424
rect 4173 3384 4185 3424
rect 4207 3384 4219 3424
rect 4227 3384 4239 3464
rect 4271 3384 4283 3424
rect 4291 3384 4303 3424
rect 4331 3384 4343 3424
rect 4351 3384 4363 3424
rect 4377 3384 4389 3424
rect 4397 3384 4409 3424
rect 4417 3384 4429 3424
rect 4461 3384 4473 3464
rect 4481 3384 4493 3424
rect 4515 3384 4527 3424
rect 4547 3384 4559 3424
rect 4567 3384 4579 3424
rect 4593 3384 4605 3424
rect 4621 3384 4633 3404
rect 4651 3384 4663 3404
rect 4671 3384 4683 3464
rect 4711 3384 4723 3424
rect 4731 3384 4743 3424
rect 4757 3384 4769 3464
rect 4777 3384 4789 3404
rect 4807 3384 4819 3404
rect 4835 3384 4847 3424
rect 4861 3384 4873 3424
rect 4881 3384 4893 3424
rect 4913 3384 4925 3424
rect 4947 3384 4959 3424
rect 4967 3384 4979 3464
rect 5011 3384 5023 3464
rect 5031 3396 5043 3464
rect 5051 3384 5063 3462
rect 5071 3384 5083 3450
rect 5091 3384 5103 3462
rect 5131 3384 5143 3424
rect 5151 3384 5163 3424
rect 5177 3384 5189 3464
rect 5197 3384 5209 3404
rect 5227 3384 5239 3404
rect 5255 3384 5267 3424
rect 5281 3384 5293 3424
rect 5301 3384 5313 3424
rect 5333 3384 5345 3424
rect 5367 3384 5379 3424
rect 5387 3384 5399 3464
rect 5417 3384 5429 3464
rect 5437 3384 5449 3404
rect 5467 3384 5479 3404
rect 5495 3384 5507 3424
rect 5521 3384 5533 3424
rect 5541 3384 5553 3424
rect 5573 3384 5585 3424
rect 5607 3384 5619 3424
rect 5627 3384 5639 3464
rect 5662 3384 5674 3464
rect 5690 3384 5702 3464
rect 5712 3384 5724 3424
rect 5762 3384 5774 3464
rect 5790 3384 5802 3464
rect 5812 3384 5824 3424
rect 5871 3384 5883 3424
rect 5891 3384 5903 3424
rect 5931 3384 5943 3464
rect 5951 3396 5963 3464
rect 5971 3384 5983 3462
rect 5991 3384 6003 3450
rect 6011 3384 6023 3462
rect 6037 3384 6049 3424
rect 6057 3384 6069 3424
rect 6077 3384 6089 3424
rect 6131 3384 6143 3424
rect 6151 3384 6163 3424
rect 6177 3384 6189 3444
rect 6197 3384 6209 3444
rect 6217 3384 6229 3444
rect 6237 3396 6249 3444
rect 6257 3384 6269 3442
rect 6281 3392 6293 3452
rect 6301 3396 6313 3448
rect 6321 3392 6333 3452
rect 6371 3384 6383 3424
rect 6391 3384 6403 3424
rect 6417 3384 6429 3464
rect 6437 3384 6449 3404
rect 6467 3384 6479 3404
rect 6495 3384 6507 3424
rect 6521 3384 6533 3424
rect 6541 3384 6553 3424
rect 6573 3384 6585 3424
rect 6607 3384 6619 3424
rect 6627 3384 6639 3464
rect 29 3276 41 3356
rect 49 3276 61 3356
rect 71 3316 83 3356
rect 97 3276 109 3356
rect 117 3336 129 3356
rect 147 3336 159 3356
rect 175 3316 187 3356
rect 201 3316 213 3356
rect 221 3316 233 3356
rect 253 3316 265 3356
rect 287 3316 299 3356
rect 307 3276 319 3356
rect 337 3316 349 3356
rect 357 3316 369 3356
rect 377 3316 389 3356
rect 431 3276 443 3356
rect 451 3276 463 3356
rect 471 3288 483 3356
rect 491 3284 503 3356
rect 531 3316 543 3356
rect 551 3316 563 3356
rect 571 3316 583 3356
rect 597 3316 609 3356
rect 617 3316 629 3356
rect 657 3316 669 3356
rect 677 3316 689 3356
rect 697 3320 709 3356
rect 717 3316 729 3356
rect 757 3316 769 3356
rect 777 3316 789 3356
rect 797 3316 809 3356
rect 856 3316 868 3356
rect 878 3276 890 3356
rect 906 3276 918 3356
rect 937 3316 949 3356
rect 957 3316 969 3356
rect 997 3276 1009 3356
rect 1025 3276 1037 3356
rect 1082 3276 1094 3356
rect 1110 3276 1122 3356
rect 1132 3316 1144 3356
rect 1182 3276 1194 3356
rect 1210 3276 1222 3356
rect 1232 3316 1244 3356
rect 1277 3316 1289 3356
rect 1297 3316 1309 3356
rect 1317 3316 1329 3356
rect 1357 3276 1369 3356
rect 1377 3336 1389 3356
rect 1407 3336 1419 3356
rect 1435 3316 1447 3356
rect 1461 3316 1473 3356
rect 1481 3316 1493 3356
rect 1513 3316 1525 3356
rect 1547 3316 1559 3356
rect 1567 3276 1579 3356
rect 1607 3276 1619 3356
rect 1627 3276 1639 3356
rect 1651 3316 1663 3356
rect 1671 3316 1683 3356
rect 1711 3276 1723 3356
rect 1731 3276 1743 3356
rect 1751 3288 1763 3356
rect 1771 3284 1783 3356
rect 1811 3316 1823 3356
rect 1831 3320 1843 3356
rect 1851 3316 1863 3356
rect 1871 3316 1883 3356
rect 1897 3284 1909 3356
rect 1917 3288 1929 3356
rect 1937 3276 1949 3356
rect 1957 3276 1969 3356
rect 2001 3276 2013 3356
rect 2021 3316 2033 3356
rect 2055 3316 2067 3356
rect 2087 3316 2099 3356
rect 2107 3316 2119 3356
rect 2133 3316 2145 3356
rect 2161 3336 2173 3356
rect 2191 3336 2203 3356
rect 2211 3276 2223 3356
rect 2237 3316 2249 3356
rect 2257 3316 2269 3356
rect 2277 3316 2289 3356
rect 2317 3276 2329 3356
rect 2345 3276 2357 3356
rect 2423 3276 2435 3356
rect 2451 3276 2463 3356
rect 2496 3316 2508 3356
rect 2518 3276 2530 3356
rect 2546 3276 2558 3356
rect 2577 3316 2589 3356
rect 2597 3316 2609 3356
rect 2641 3276 2653 3356
rect 2661 3316 2673 3356
rect 2695 3316 2707 3356
rect 2727 3316 2739 3356
rect 2747 3316 2759 3356
rect 2773 3316 2785 3356
rect 2801 3336 2813 3356
rect 2831 3336 2843 3356
rect 2851 3276 2863 3356
rect 2877 3316 2889 3356
rect 2897 3316 2909 3356
rect 2917 3316 2929 3356
rect 2971 3316 2983 3356
rect 2991 3316 3003 3356
rect 3011 3316 3023 3356
rect 3056 3316 3068 3356
rect 3078 3276 3090 3356
rect 3106 3276 3118 3356
rect 3151 3316 3163 3356
rect 3171 3316 3183 3356
rect 3191 3316 3203 3356
rect 3231 3316 3243 3356
rect 3251 3316 3263 3356
rect 3296 3316 3308 3356
rect 3318 3276 3330 3356
rect 3346 3276 3358 3356
rect 3377 3316 3389 3356
rect 3397 3316 3409 3356
rect 3463 3276 3475 3356
rect 3491 3276 3503 3356
rect 3531 3276 3543 3356
rect 3551 3276 3563 3356
rect 3571 3288 3583 3356
rect 3591 3284 3603 3356
rect 3643 3276 3655 3356
rect 3671 3276 3683 3356
rect 3697 3276 3709 3356
rect 3717 3336 3729 3356
rect 3747 3336 3759 3356
rect 3775 3316 3787 3356
rect 3801 3316 3813 3356
rect 3821 3316 3833 3356
rect 3853 3316 3865 3356
rect 3887 3316 3899 3356
rect 3907 3276 3919 3356
rect 3937 3278 3949 3356
rect 3957 3290 3969 3356
rect 3977 3278 3989 3356
rect 3997 3276 4009 3344
rect 4017 3276 4029 3356
rect 4071 3276 4083 3356
rect 4091 3276 4103 3344
rect 4111 3278 4123 3356
rect 4131 3290 4143 3356
rect 4151 3278 4163 3356
rect 4181 3276 4193 3356
rect 4201 3316 4213 3356
rect 4235 3316 4247 3356
rect 4267 3316 4279 3356
rect 4287 3316 4299 3356
rect 4313 3316 4325 3356
rect 4341 3336 4353 3356
rect 4371 3336 4383 3356
rect 4391 3276 4403 3356
rect 4417 3276 4429 3356
rect 4445 3276 4457 3356
rect 4497 3278 4509 3356
rect 4517 3290 4529 3356
rect 4537 3278 4549 3356
rect 4557 3276 4569 3344
rect 4577 3276 4589 3356
rect 4617 3276 4629 3356
rect 4645 3276 4657 3356
rect 4697 3276 4709 3356
rect 4725 3276 4737 3356
rect 4777 3316 4789 3356
rect 4797 3316 4809 3356
rect 4837 3278 4849 3356
rect 4857 3290 4869 3356
rect 4877 3278 4889 3356
rect 4897 3276 4909 3344
rect 4917 3276 4929 3356
rect 4957 3284 4969 3356
rect 4977 3288 4989 3356
rect 4997 3276 5009 3356
rect 5017 3276 5029 3356
rect 5057 3276 5069 3356
rect 5077 3336 5089 3356
rect 5107 3336 5119 3356
rect 5135 3316 5147 3356
rect 5161 3316 5173 3356
rect 5181 3316 5193 3356
rect 5213 3316 5225 3356
rect 5247 3316 5259 3356
rect 5267 3276 5279 3356
rect 5311 3316 5323 3356
rect 5331 3316 5343 3356
rect 5357 3308 5369 3348
rect 5377 3308 5389 3348
rect 5407 3284 5419 3348
rect 5437 3276 5449 3356
rect 5491 3316 5503 3356
rect 5511 3316 5523 3356
rect 5541 3276 5553 3356
rect 5561 3316 5573 3356
rect 5595 3316 5607 3356
rect 5627 3316 5639 3356
rect 5647 3316 5659 3356
rect 5673 3316 5685 3356
rect 5701 3336 5713 3356
rect 5731 3336 5743 3356
rect 5751 3276 5763 3356
rect 5796 3316 5808 3356
rect 5818 3276 5830 3356
rect 5846 3276 5858 3356
rect 5891 3316 5903 3356
rect 5911 3316 5923 3356
rect 5951 3276 5963 3356
rect 5971 3276 5983 3356
rect 5991 3288 6003 3356
rect 6011 3284 6023 3356
rect 6042 3276 6054 3356
rect 6070 3276 6082 3356
rect 6092 3316 6104 3356
rect 6151 3316 6163 3356
rect 6171 3316 6183 3356
rect 6191 3316 6203 3356
rect 6231 3276 6243 3356
rect 6251 3276 6263 3356
rect 6271 3288 6283 3356
rect 6291 3284 6303 3356
rect 6331 3316 6343 3356
rect 6351 3316 6363 3356
rect 6371 3316 6383 3356
rect 6402 3276 6414 3356
rect 6430 3276 6442 3356
rect 6452 3316 6464 3356
rect 6497 3276 6509 3356
rect 6517 3336 6529 3356
rect 6547 3336 6559 3356
rect 6575 3316 6587 3356
rect 6601 3316 6613 3356
rect 6621 3316 6633 3356
rect 6653 3316 6665 3356
rect 6687 3316 6699 3356
rect 6707 3276 6719 3356
rect 17 2904 29 2984
rect 37 2904 49 2984
rect 57 2904 69 2984
rect 77 2904 89 2984
rect 97 2904 109 2984
rect 117 2904 129 2984
rect 137 2904 149 2984
rect 157 2904 169 2984
rect 177 2904 189 2984
rect 229 2904 241 2984
rect 249 2904 261 2984
rect 271 2904 283 2944
rect 301 2904 313 2984
rect 321 2904 333 2944
rect 355 2904 367 2944
rect 387 2904 399 2944
rect 407 2904 419 2944
rect 433 2904 445 2944
rect 461 2904 473 2924
rect 491 2904 503 2924
rect 511 2904 523 2984
rect 551 2904 563 2944
rect 571 2904 583 2944
rect 591 2904 603 2944
rect 617 2904 629 2944
rect 637 2904 649 2944
rect 657 2904 669 2944
rect 716 2904 728 2944
rect 738 2904 750 2984
rect 766 2904 778 2984
rect 811 2904 823 2944
rect 831 2904 843 2944
rect 851 2904 863 2944
rect 891 2904 903 2944
rect 911 2904 923 2944
rect 931 2904 943 2944
rect 957 2904 969 2976
rect 977 2904 989 2972
rect 997 2904 1009 2984
rect 1017 2904 1029 2984
rect 1057 2904 1069 2984
rect 1077 2904 1089 2924
rect 1107 2904 1119 2924
rect 1135 2904 1147 2944
rect 1161 2904 1173 2944
rect 1181 2904 1193 2944
rect 1213 2904 1225 2944
rect 1247 2904 1259 2944
rect 1267 2904 1279 2984
rect 1311 2904 1323 2944
rect 1331 2904 1343 2944
rect 1351 2904 1363 2944
rect 1377 2904 1389 2984
rect 1397 2904 1409 2924
rect 1427 2904 1439 2924
rect 1455 2904 1467 2944
rect 1481 2904 1493 2944
rect 1501 2904 1513 2944
rect 1533 2904 1545 2944
rect 1567 2904 1579 2944
rect 1587 2904 1599 2984
rect 1631 2904 1643 2944
rect 1651 2904 1663 2944
rect 1696 2904 1708 2944
rect 1718 2904 1730 2984
rect 1746 2904 1758 2984
rect 1803 2904 1815 2984
rect 1831 2904 1843 2984
rect 1867 2904 1879 2984
rect 1887 2904 1899 2984
rect 1911 2904 1923 2944
rect 1931 2904 1943 2944
rect 1962 2904 1974 2984
rect 1990 2904 2002 2984
rect 2012 2904 2024 2944
rect 2071 2904 2083 2984
rect 2091 2904 2103 2984
rect 2111 2904 2123 2972
rect 2131 2904 2143 2976
rect 2157 2904 2169 2944
rect 2177 2904 2189 2944
rect 2197 2904 2209 2944
rect 2251 2904 2263 2944
rect 2271 2904 2283 2944
rect 2297 2904 2309 2944
rect 2317 2904 2329 2944
rect 2341 2904 2353 2984
rect 2361 2904 2373 2984
rect 2401 2904 2413 2984
rect 2421 2904 2433 2944
rect 2455 2904 2467 2944
rect 2487 2904 2499 2944
rect 2507 2904 2519 2944
rect 2533 2904 2545 2944
rect 2561 2904 2573 2924
rect 2591 2904 2603 2924
rect 2611 2904 2623 2984
rect 2637 2904 2649 2944
rect 2657 2904 2669 2944
rect 2697 2904 2709 2984
rect 2725 2904 2737 2984
rect 2791 2904 2803 2944
rect 2811 2904 2823 2944
rect 2856 2904 2868 2944
rect 2878 2904 2890 2984
rect 2906 2904 2918 2984
rect 2937 2904 2949 2984
rect 2957 2904 2969 2984
rect 3011 2904 3023 2944
rect 3031 2904 3043 2940
rect 3051 2904 3063 2944
rect 3071 2904 3083 2944
rect 3111 2904 3123 2944
rect 3131 2904 3143 2944
rect 3151 2904 3163 2944
rect 3196 2904 3208 2944
rect 3218 2904 3230 2984
rect 3246 2904 3258 2984
rect 3277 2904 3289 2944
rect 3297 2904 3309 2944
rect 3317 2904 3329 2944
rect 3357 2904 3369 2944
rect 3377 2904 3389 2944
rect 3397 2904 3409 2944
rect 3442 2904 3454 2984
rect 3470 2904 3482 2984
rect 3492 2904 3504 2944
rect 3537 2904 3549 2944
rect 3557 2904 3569 2944
rect 3581 2904 3593 2984
rect 3601 2904 3613 2984
rect 3651 2904 3663 2984
rect 3671 2916 3683 2984
rect 3691 2904 3703 2982
rect 3711 2904 3723 2970
rect 3731 2904 3743 2982
rect 3771 2904 3783 2984
rect 3791 2904 3803 2984
rect 3811 2906 3823 2984
rect 3841 2904 3853 2984
rect 3861 2904 3873 2944
rect 3895 2904 3907 2944
rect 3927 2904 3939 2944
rect 3947 2904 3959 2944
rect 3973 2904 3985 2944
rect 4001 2904 4013 2924
rect 4031 2904 4043 2924
rect 4051 2904 4063 2984
rect 4082 2904 4094 2984
rect 4110 2904 4122 2984
rect 4132 2904 4144 2944
rect 4191 2904 4203 2944
rect 4211 2904 4223 2940
rect 4231 2904 4243 2944
rect 4251 2904 4263 2944
rect 4281 2904 4293 2984
rect 4301 2904 4313 2944
rect 4335 2904 4347 2944
rect 4367 2904 4379 2944
rect 4387 2904 4399 2944
rect 4413 2904 4425 2944
rect 4441 2904 4453 2924
rect 4471 2904 4483 2924
rect 4491 2904 4503 2984
rect 4541 2904 4553 2984
rect 4571 2904 4593 2984
rect 4611 2904 4623 2984
rect 4651 2904 4663 2944
rect 4671 2904 4683 2944
rect 4711 2904 4723 2984
rect 4741 2912 4753 2976
rect 4771 2912 4783 2952
rect 4791 2912 4803 2952
rect 4817 2904 4829 2982
rect 4837 2904 4849 2970
rect 4857 2904 4869 2982
rect 4877 2916 4889 2984
rect 4897 2904 4909 2984
rect 4951 2904 4963 2944
rect 4971 2904 4983 2944
rect 4997 2904 5009 2982
rect 5017 2904 5029 2970
rect 5037 2904 5049 2982
rect 5057 2916 5069 2984
rect 5077 2904 5089 2984
rect 5117 2904 5129 2944
rect 5137 2904 5149 2944
rect 5177 2904 5189 2984
rect 5205 2904 5217 2984
rect 5261 2904 5273 2984
rect 5281 2904 5293 2944
rect 5315 2904 5327 2944
rect 5347 2904 5359 2944
rect 5367 2904 5379 2944
rect 5393 2904 5405 2944
rect 5421 2904 5433 2924
rect 5451 2904 5463 2924
rect 5471 2904 5483 2984
rect 5523 2904 5535 2984
rect 5551 2904 5563 2984
rect 5582 2904 5594 2984
rect 5610 2904 5622 2984
rect 5632 2904 5644 2944
rect 5691 2904 5703 2944
rect 5711 2904 5723 2940
rect 5731 2904 5743 2944
rect 5751 2904 5763 2944
rect 5801 2904 5813 2984
rect 5831 2904 5853 2984
rect 5871 2904 5883 2984
rect 5897 2904 5909 2944
rect 5917 2904 5929 2944
rect 5957 2912 5969 2952
rect 5977 2912 5989 2952
rect 6007 2912 6019 2976
rect 6037 2904 6049 2984
rect 6091 2904 6103 2984
rect 6111 2904 6123 2984
rect 6131 2904 6143 2972
rect 6151 2904 6163 2976
rect 6203 2904 6215 2984
rect 6231 2904 6243 2984
rect 6257 2904 6269 2944
rect 6277 2904 6289 2944
rect 6331 2904 6343 2984
rect 6351 2916 6363 2984
rect 6371 2904 6383 2982
rect 6391 2904 6403 2970
rect 6411 2904 6423 2982
rect 6451 2904 6463 2944
rect 6471 2904 6483 2944
rect 6497 2904 6509 2944
rect 6517 2904 6529 2944
rect 6562 2904 6574 2984
rect 6590 2904 6602 2984
rect 6612 2904 6624 2944
rect 17 2836 29 2876
rect 37 2836 49 2876
rect 103 2796 115 2876
rect 131 2796 143 2876
rect 161 2796 173 2876
rect 181 2836 193 2876
rect 215 2836 227 2876
rect 247 2836 259 2876
rect 267 2836 279 2876
rect 293 2836 305 2876
rect 321 2856 333 2876
rect 351 2856 363 2876
rect 371 2796 383 2876
rect 397 2836 409 2876
rect 417 2836 429 2876
rect 483 2796 495 2876
rect 511 2796 523 2876
rect 541 2796 553 2876
rect 561 2836 573 2876
rect 595 2836 607 2876
rect 627 2836 639 2876
rect 647 2836 659 2876
rect 673 2836 685 2876
rect 701 2856 713 2876
rect 731 2856 743 2876
rect 751 2796 763 2876
rect 789 2796 801 2876
rect 809 2796 821 2876
rect 831 2836 843 2876
rect 857 2796 869 2874
rect 877 2796 889 2876
rect 897 2796 909 2876
rect 937 2836 949 2876
rect 957 2836 969 2876
rect 977 2836 989 2876
rect 1017 2836 1029 2876
rect 1037 2836 1049 2876
rect 1057 2836 1069 2876
rect 1097 2836 1109 2876
rect 1117 2836 1129 2876
rect 1157 2798 1169 2876
rect 1177 2810 1189 2876
rect 1197 2798 1209 2876
rect 1217 2796 1229 2864
rect 1237 2796 1249 2876
rect 1291 2796 1303 2876
rect 1311 2796 1323 2876
rect 1331 2808 1343 2876
rect 1351 2804 1363 2876
rect 1391 2836 1403 2876
rect 1411 2836 1423 2876
rect 1456 2836 1468 2876
rect 1478 2796 1490 2876
rect 1506 2796 1518 2876
rect 1537 2796 1549 2876
rect 1565 2796 1577 2876
rect 1617 2836 1629 2876
rect 1637 2836 1649 2876
rect 1657 2836 1669 2876
rect 1697 2796 1709 2876
rect 1725 2796 1737 2876
rect 1796 2836 1808 2876
rect 1818 2796 1830 2876
rect 1846 2796 1858 2876
rect 1877 2796 1889 2876
rect 1907 2797 1919 2876
rect 1927 2797 1939 2876
rect 1982 2796 1994 2876
rect 2010 2796 2022 2876
rect 2032 2836 2044 2876
rect 2091 2796 2103 2876
rect 2111 2796 2123 2876
rect 2131 2808 2143 2876
rect 2151 2804 2163 2876
rect 2181 2796 2193 2876
rect 2201 2836 2213 2876
rect 2235 2836 2247 2876
rect 2267 2836 2279 2876
rect 2287 2836 2299 2876
rect 2313 2836 2325 2876
rect 2341 2856 2353 2876
rect 2371 2856 2383 2876
rect 2391 2796 2403 2876
rect 2417 2836 2429 2876
rect 2437 2836 2449 2876
rect 2457 2836 2469 2876
rect 2497 2836 2509 2876
rect 2517 2836 2529 2876
rect 2571 2836 2583 2876
rect 2591 2836 2603 2876
rect 2621 2796 2633 2876
rect 2641 2836 2653 2876
rect 2675 2836 2687 2876
rect 2707 2836 2719 2876
rect 2727 2836 2739 2876
rect 2753 2836 2765 2876
rect 2781 2856 2793 2876
rect 2811 2856 2823 2876
rect 2831 2796 2843 2876
rect 2862 2796 2874 2876
rect 2890 2796 2902 2876
rect 2912 2836 2924 2876
rect 2971 2796 2983 2876
rect 2991 2796 3003 2876
rect 3011 2808 3023 2876
rect 3031 2804 3043 2876
rect 3057 2796 3069 2876
rect 3077 2856 3089 2876
rect 3107 2856 3119 2876
rect 3135 2836 3147 2876
rect 3161 2836 3173 2876
rect 3181 2836 3193 2876
rect 3213 2836 3225 2876
rect 3247 2836 3259 2876
rect 3267 2796 3279 2876
rect 3297 2836 3309 2876
rect 3317 2836 3329 2876
rect 3357 2796 3369 2876
rect 3387 2796 3409 2876
rect 3427 2796 3439 2876
rect 3482 2796 3494 2876
rect 3510 2796 3522 2876
rect 3532 2836 3544 2876
rect 3601 2796 3613 2876
rect 3631 2796 3653 2876
rect 3671 2796 3683 2876
rect 3702 2796 3714 2876
rect 3730 2796 3742 2876
rect 3752 2836 3764 2876
rect 3821 2796 3833 2876
rect 3851 2796 3873 2876
rect 3891 2796 3903 2876
rect 3931 2836 3943 2876
rect 3951 2836 3963 2876
rect 3977 2796 3989 2876
rect 4005 2796 4017 2876
rect 4057 2796 4069 2876
rect 4085 2796 4097 2876
rect 4151 2796 4163 2876
rect 4171 2796 4183 2876
rect 4191 2808 4203 2876
rect 4211 2804 4223 2876
rect 4242 2796 4254 2876
rect 4270 2796 4282 2876
rect 4292 2836 4304 2876
rect 4351 2836 4363 2876
rect 4371 2840 4383 2876
rect 4391 2836 4403 2876
rect 4411 2836 4423 2876
rect 4441 2796 4453 2876
rect 4461 2836 4473 2876
rect 4495 2836 4507 2876
rect 4527 2836 4539 2876
rect 4547 2836 4559 2876
rect 4573 2836 4585 2876
rect 4601 2856 4613 2876
rect 4631 2856 4643 2876
rect 4651 2796 4663 2876
rect 4677 2836 4689 2876
rect 4697 2836 4709 2876
rect 4737 2796 4749 2876
rect 4765 2796 4777 2876
rect 4822 2796 4834 2876
rect 4850 2796 4862 2876
rect 4872 2836 4884 2876
rect 4943 2796 4955 2876
rect 4971 2796 4983 2876
rect 5021 2796 5033 2876
rect 5051 2796 5073 2876
rect 5091 2796 5103 2876
rect 5117 2804 5129 2876
rect 5137 2808 5149 2876
rect 5157 2796 5169 2876
rect 5177 2796 5189 2876
rect 5217 2836 5229 2876
rect 5239 2796 5251 2876
rect 5259 2796 5271 2876
rect 5302 2796 5314 2876
rect 5330 2796 5342 2876
rect 5352 2836 5364 2876
rect 5421 2796 5433 2876
rect 5451 2796 5473 2876
rect 5491 2796 5503 2876
rect 5531 2836 5543 2876
rect 5551 2836 5563 2876
rect 5581 2796 5593 2876
rect 5601 2836 5613 2876
rect 5635 2836 5647 2876
rect 5667 2836 5679 2876
rect 5687 2836 5699 2876
rect 5713 2836 5725 2876
rect 5741 2856 5753 2876
rect 5771 2856 5783 2876
rect 5791 2796 5803 2876
rect 5817 2828 5829 2868
rect 5837 2828 5849 2868
rect 5867 2804 5879 2868
rect 5897 2796 5909 2876
rect 5937 2828 5949 2868
rect 5957 2828 5969 2868
rect 5987 2804 5999 2868
rect 6017 2796 6029 2876
rect 6057 2828 6069 2868
rect 6077 2828 6089 2868
rect 6107 2804 6119 2868
rect 6137 2796 6149 2876
rect 6187 2796 6199 2876
rect 6207 2796 6219 2876
rect 6231 2836 6243 2876
rect 6251 2836 6263 2876
rect 6291 2796 6303 2876
rect 6311 2796 6323 2876
rect 6331 2796 6343 2874
rect 6357 2836 6369 2876
rect 6377 2836 6389 2876
rect 6401 2796 6413 2876
rect 6421 2796 6433 2876
rect 6457 2796 6469 2876
rect 6477 2856 6489 2876
rect 6507 2856 6519 2876
rect 6535 2836 6547 2876
rect 6561 2836 6573 2876
rect 6581 2836 6593 2876
rect 6613 2836 6625 2876
rect 6647 2836 6659 2876
rect 6667 2796 6679 2876
rect 17 2424 29 2504
rect 37 2424 49 2444
rect 67 2424 79 2444
rect 95 2424 107 2464
rect 121 2424 133 2464
rect 141 2424 153 2464
rect 173 2424 185 2464
rect 207 2424 219 2464
rect 227 2424 239 2504
rect 269 2424 281 2504
rect 289 2424 301 2504
rect 311 2424 323 2464
rect 337 2424 349 2504
rect 357 2424 369 2444
rect 387 2424 399 2444
rect 415 2424 427 2464
rect 441 2424 453 2464
rect 461 2424 473 2464
rect 493 2424 505 2464
rect 527 2424 539 2464
rect 547 2424 559 2504
rect 591 2424 603 2504
rect 611 2424 623 2504
rect 631 2424 643 2492
rect 651 2424 663 2496
rect 677 2424 689 2464
rect 697 2424 709 2464
rect 717 2424 729 2464
rect 771 2424 783 2464
rect 791 2424 803 2464
rect 811 2424 823 2464
rect 851 2424 863 2504
rect 871 2424 883 2504
rect 891 2424 903 2504
rect 911 2424 923 2504
rect 931 2424 943 2504
rect 951 2424 963 2504
rect 971 2424 983 2504
rect 991 2424 1003 2504
rect 1011 2424 1023 2504
rect 1037 2424 1049 2504
rect 1057 2424 1069 2444
rect 1087 2424 1099 2444
rect 1115 2424 1127 2464
rect 1141 2424 1153 2464
rect 1161 2424 1173 2464
rect 1193 2424 1205 2464
rect 1227 2424 1239 2464
rect 1247 2424 1259 2504
rect 1291 2424 1303 2464
rect 1311 2424 1323 2464
rect 1331 2424 1343 2464
rect 1357 2424 1369 2504
rect 1385 2424 1397 2504
rect 1437 2424 1449 2464
rect 1457 2424 1469 2464
rect 1516 2424 1528 2464
rect 1538 2424 1550 2504
rect 1566 2424 1578 2504
rect 1601 2424 1613 2504
rect 1621 2424 1633 2464
rect 1655 2424 1667 2464
rect 1687 2424 1699 2464
rect 1707 2424 1719 2464
rect 1733 2424 1745 2464
rect 1761 2424 1773 2444
rect 1791 2424 1803 2444
rect 1811 2424 1823 2504
rect 1837 2424 1849 2464
rect 1857 2424 1869 2464
rect 1897 2424 1909 2464
rect 1917 2424 1929 2464
rect 1957 2424 1969 2504
rect 1987 2424 2009 2504
rect 2027 2424 2039 2504
rect 2077 2424 2089 2504
rect 2105 2424 2117 2504
rect 2157 2432 2169 2472
rect 2177 2432 2189 2472
rect 2207 2432 2219 2496
rect 2237 2424 2249 2504
rect 2277 2432 2289 2472
rect 2297 2432 2309 2472
rect 2327 2432 2339 2496
rect 2357 2424 2369 2504
rect 2401 2424 2413 2504
rect 2421 2424 2433 2464
rect 2455 2424 2467 2464
rect 2487 2424 2499 2464
rect 2507 2424 2519 2464
rect 2533 2424 2545 2464
rect 2561 2424 2573 2444
rect 2591 2424 2603 2444
rect 2611 2424 2623 2504
rect 2637 2432 2649 2472
rect 2657 2432 2669 2472
rect 2687 2432 2699 2496
rect 2717 2424 2729 2504
rect 2783 2424 2795 2504
rect 2811 2424 2823 2504
rect 2851 2424 2863 2504
rect 2881 2432 2893 2496
rect 2911 2432 2923 2472
rect 2931 2432 2943 2472
rect 2981 2424 2993 2504
rect 3011 2424 3033 2504
rect 3051 2424 3063 2504
rect 3091 2424 3103 2464
rect 3111 2424 3123 2464
rect 3141 2424 3153 2504
rect 3161 2424 3173 2464
rect 3195 2424 3207 2464
rect 3227 2424 3239 2464
rect 3247 2424 3259 2464
rect 3273 2424 3285 2464
rect 3301 2424 3313 2444
rect 3331 2424 3343 2444
rect 3351 2424 3363 2504
rect 3377 2424 3389 2504
rect 3405 2424 3417 2504
rect 3471 2424 3483 2464
rect 3491 2424 3503 2464
rect 3511 2424 3523 2464
rect 3537 2424 3549 2464
rect 3557 2424 3569 2464
rect 3597 2424 3609 2464
rect 3617 2424 3629 2464
rect 3637 2424 3649 2460
rect 3657 2424 3669 2464
rect 3697 2424 3709 2464
rect 3717 2424 3729 2464
rect 3737 2424 3749 2460
rect 3757 2424 3769 2464
rect 3811 2424 3823 2464
rect 3831 2424 3843 2460
rect 3851 2424 3863 2464
rect 3871 2424 3883 2464
rect 3902 2424 3914 2504
rect 3930 2424 3942 2504
rect 3952 2424 3964 2464
rect 3997 2424 4009 2496
rect 4017 2424 4029 2492
rect 4037 2424 4049 2504
rect 4057 2424 4069 2504
rect 4123 2424 4135 2504
rect 4151 2424 4163 2504
rect 4201 2424 4213 2504
rect 4231 2424 4253 2504
rect 4271 2424 4283 2504
rect 4301 2424 4313 2504
rect 4321 2424 4333 2464
rect 4355 2424 4367 2464
rect 4387 2424 4399 2464
rect 4407 2424 4419 2464
rect 4433 2424 4445 2464
rect 4461 2424 4473 2444
rect 4491 2424 4503 2444
rect 4511 2424 4523 2504
rect 4551 2424 4563 2464
rect 4571 2424 4583 2464
rect 4621 2424 4633 2504
rect 4651 2424 4673 2504
rect 4691 2424 4703 2504
rect 4717 2432 4729 2472
rect 4737 2432 4749 2472
rect 4767 2432 4779 2496
rect 4797 2424 4809 2504
rect 4837 2424 4849 2504
rect 4857 2424 4869 2444
rect 4887 2424 4899 2444
rect 4915 2424 4927 2464
rect 4941 2424 4953 2464
rect 4961 2424 4973 2464
rect 4993 2424 5005 2464
rect 5027 2424 5039 2464
rect 5047 2424 5059 2504
rect 5077 2424 5089 2464
rect 5097 2424 5109 2464
rect 5137 2424 5149 2504
rect 5167 2424 5189 2504
rect 5207 2424 5219 2504
rect 5262 2424 5274 2504
rect 5290 2424 5302 2504
rect 5312 2424 5324 2464
rect 5357 2424 5369 2504
rect 5385 2424 5397 2504
rect 5463 2424 5475 2504
rect 5491 2424 5503 2504
rect 5517 2424 5529 2504
rect 5537 2424 5549 2504
rect 5557 2424 5569 2504
rect 5577 2424 5589 2504
rect 5597 2424 5609 2504
rect 5617 2424 5629 2504
rect 5637 2424 5649 2504
rect 5657 2424 5669 2504
rect 5677 2424 5689 2504
rect 5743 2424 5755 2504
rect 5771 2424 5783 2504
rect 5802 2424 5814 2504
rect 5830 2424 5842 2504
rect 5852 2424 5864 2464
rect 5921 2424 5933 2504
rect 5951 2424 5973 2504
rect 5991 2424 6003 2504
rect 6031 2424 6043 2464
rect 6051 2424 6063 2464
rect 6077 2424 6089 2504
rect 6097 2424 6109 2444
rect 6127 2424 6139 2444
rect 6155 2424 6167 2464
rect 6181 2424 6193 2464
rect 6201 2424 6213 2464
rect 6233 2424 6245 2464
rect 6267 2424 6279 2464
rect 6287 2424 6299 2504
rect 6331 2424 6343 2504
rect 6351 2436 6363 2504
rect 6371 2424 6383 2502
rect 6391 2424 6403 2490
rect 6411 2424 6423 2502
rect 6437 2426 6449 2504
rect 6457 2424 6469 2504
rect 6477 2424 6489 2504
rect 6517 2424 6529 2464
rect 6537 2424 6549 2464
rect 6577 2424 6589 2502
rect 6597 2424 6609 2490
rect 6617 2424 6629 2502
rect 6637 2436 6649 2504
rect 6657 2424 6669 2504
rect 21 2316 33 2396
rect 41 2356 53 2396
rect 75 2356 87 2396
rect 107 2356 119 2396
rect 127 2356 139 2396
rect 153 2356 165 2396
rect 181 2376 193 2396
rect 211 2376 223 2396
rect 231 2316 243 2396
rect 269 2316 281 2396
rect 289 2316 301 2396
rect 311 2356 323 2396
rect 351 2316 363 2396
rect 371 2316 383 2396
rect 411 2356 423 2396
rect 431 2356 443 2396
rect 483 2316 495 2396
rect 511 2316 523 2396
rect 542 2316 554 2396
rect 570 2316 582 2396
rect 592 2356 604 2396
rect 647 2316 659 2396
rect 667 2316 679 2396
rect 691 2356 703 2396
rect 711 2356 723 2396
rect 737 2356 749 2396
rect 757 2356 769 2396
rect 777 2360 789 2396
rect 797 2356 809 2396
rect 837 2356 849 2396
rect 857 2356 869 2396
rect 877 2356 889 2396
rect 917 2316 929 2396
rect 937 2376 949 2396
rect 967 2376 979 2396
rect 995 2356 1007 2396
rect 1021 2356 1033 2396
rect 1041 2356 1053 2396
rect 1073 2356 1085 2396
rect 1107 2356 1119 2396
rect 1127 2316 1139 2396
rect 1157 2356 1169 2396
rect 1177 2356 1189 2396
rect 1221 2316 1233 2396
rect 1241 2356 1253 2396
rect 1275 2356 1287 2396
rect 1307 2356 1319 2396
rect 1327 2356 1339 2396
rect 1353 2356 1365 2396
rect 1381 2376 1393 2396
rect 1411 2376 1423 2396
rect 1431 2316 1443 2396
rect 1471 2356 1483 2396
rect 1491 2356 1503 2396
rect 1517 2316 1529 2396
rect 1547 2316 1569 2396
rect 1587 2316 1599 2396
rect 1642 2316 1654 2396
rect 1670 2316 1682 2396
rect 1692 2356 1704 2396
rect 1763 2316 1775 2396
rect 1791 2316 1803 2396
rect 1843 2316 1855 2396
rect 1871 2316 1883 2396
rect 1921 2316 1933 2396
rect 1951 2316 1973 2396
rect 1991 2316 2003 2396
rect 2031 2356 2043 2396
rect 2051 2356 2063 2396
rect 2081 2316 2093 2396
rect 2101 2356 2113 2396
rect 2135 2356 2147 2396
rect 2167 2356 2179 2396
rect 2187 2356 2199 2396
rect 2213 2356 2225 2396
rect 2241 2376 2253 2396
rect 2271 2376 2283 2396
rect 2291 2316 2303 2396
rect 2343 2316 2355 2396
rect 2371 2316 2383 2396
rect 2402 2316 2414 2396
rect 2430 2316 2442 2396
rect 2452 2356 2464 2396
rect 2511 2356 2523 2396
rect 2531 2360 2543 2396
rect 2551 2356 2563 2396
rect 2571 2356 2583 2396
rect 2611 2316 2623 2396
rect 2631 2316 2643 2396
rect 2651 2328 2663 2396
rect 2671 2324 2683 2396
rect 2702 2316 2714 2396
rect 2730 2316 2742 2396
rect 2752 2356 2764 2396
rect 2823 2316 2835 2396
rect 2851 2316 2863 2396
rect 2877 2316 2889 2396
rect 2897 2376 2909 2396
rect 2927 2376 2939 2396
rect 2955 2356 2967 2396
rect 2981 2356 2993 2396
rect 3001 2356 3013 2396
rect 3033 2356 3045 2396
rect 3067 2356 3079 2396
rect 3087 2316 3099 2396
rect 3122 2316 3134 2396
rect 3150 2316 3162 2396
rect 3172 2356 3184 2396
rect 3241 2316 3253 2396
rect 3271 2316 3293 2396
rect 3311 2316 3323 2396
rect 3363 2316 3375 2396
rect 3391 2316 3403 2396
rect 3431 2356 3443 2396
rect 3451 2356 3463 2396
rect 3503 2316 3515 2396
rect 3531 2316 3543 2396
rect 3561 2316 3573 2396
rect 3581 2356 3593 2396
rect 3615 2356 3627 2396
rect 3647 2356 3659 2396
rect 3667 2356 3679 2396
rect 3693 2356 3705 2396
rect 3721 2376 3733 2396
rect 3751 2376 3763 2396
rect 3771 2316 3783 2396
rect 3797 2356 3809 2396
rect 3817 2356 3829 2396
rect 3837 2356 3849 2396
rect 3877 2356 3889 2396
rect 3897 2356 3909 2396
rect 3917 2360 3929 2396
rect 3937 2356 3949 2396
rect 3977 2348 3989 2388
rect 3997 2348 4009 2388
rect 4027 2324 4039 2388
rect 4057 2316 4069 2396
rect 4097 2348 4109 2388
rect 4117 2348 4129 2388
rect 4147 2324 4159 2388
rect 4177 2316 4189 2396
rect 4217 2348 4229 2388
rect 4237 2348 4249 2388
rect 4267 2324 4279 2388
rect 4297 2316 4309 2396
rect 4337 2356 4349 2396
rect 4359 2316 4371 2396
rect 4379 2316 4391 2396
rect 4443 2316 4455 2396
rect 4471 2316 4483 2396
rect 4497 2348 4509 2388
rect 4517 2348 4529 2388
rect 4547 2324 4559 2388
rect 4577 2316 4589 2396
rect 4631 2316 4643 2396
rect 4661 2324 4673 2388
rect 4691 2348 4703 2388
rect 4711 2348 4723 2388
rect 4737 2348 4749 2388
rect 4757 2348 4769 2388
rect 4787 2324 4799 2388
rect 4817 2316 4829 2396
rect 4857 2316 4869 2396
rect 4885 2316 4897 2396
rect 4937 2348 4949 2388
rect 4957 2348 4969 2388
rect 4987 2324 4999 2388
rect 5017 2316 5029 2396
rect 5071 2316 5083 2396
rect 5091 2316 5103 2396
rect 5111 2328 5123 2396
rect 5131 2324 5143 2396
rect 5157 2356 5169 2396
rect 5177 2356 5189 2396
rect 5217 2316 5229 2396
rect 5247 2316 5269 2396
rect 5287 2316 5299 2396
rect 5351 2316 5363 2396
rect 5381 2324 5393 2388
rect 5411 2348 5423 2388
rect 5431 2348 5443 2388
rect 5457 2348 5469 2388
rect 5477 2348 5489 2388
rect 5507 2324 5519 2388
rect 5537 2316 5549 2396
rect 5577 2348 5589 2388
rect 5597 2348 5609 2388
rect 5627 2324 5639 2388
rect 5657 2316 5669 2396
rect 5711 2356 5723 2396
rect 5731 2360 5743 2396
rect 5751 2356 5763 2396
rect 5771 2356 5783 2396
rect 5811 2356 5823 2396
rect 5831 2360 5843 2396
rect 5851 2356 5863 2396
rect 5871 2356 5883 2396
rect 5911 2356 5923 2396
rect 5931 2356 5943 2396
rect 5971 2316 5983 2396
rect 5991 2316 6003 2384
rect 6011 2318 6023 2396
rect 6031 2330 6043 2396
rect 6051 2318 6063 2396
rect 6091 2316 6103 2396
rect 6121 2324 6133 2388
rect 6151 2348 6163 2388
rect 6171 2348 6183 2388
rect 6211 2316 6223 2396
rect 6241 2324 6253 2388
rect 6271 2348 6283 2388
rect 6291 2348 6303 2388
rect 6317 2356 6329 2396
rect 6337 2356 6349 2396
rect 6382 2316 6394 2396
rect 6410 2316 6422 2396
rect 6432 2356 6444 2396
rect 6477 2356 6489 2396
rect 6497 2356 6509 2396
rect 6517 2356 6529 2396
rect 6557 2324 6569 2396
rect 6577 2328 6589 2396
rect 6597 2316 6609 2396
rect 6617 2316 6629 2396
rect 6657 2356 6669 2396
rect 6677 2356 6689 2396
rect 43 1944 55 2024
rect 71 1944 83 2024
rect 111 1944 123 1984
rect 131 1944 143 1984
rect 151 1944 163 1984
rect 191 1944 203 1984
rect 211 1944 223 1980
rect 231 1944 243 1984
rect 251 1944 263 1984
rect 291 1944 303 1984
rect 311 1944 323 1980
rect 331 1944 343 1984
rect 351 1944 363 1984
rect 391 1944 403 1984
rect 411 1944 423 1984
rect 431 1944 443 1984
rect 457 1944 469 1984
rect 477 1944 489 1984
rect 497 1944 509 1980
rect 517 1944 529 1984
rect 583 1944 595 2024
rect 611 1944 623 2024
rect 642 1944 654 2024
rect 670 1944 682 2024
rect 692 1944 704 1984
rect 737 1944 749 1984
rect 757 1944 769 1984
rect 777 1944 789 1980
rect 797 1944 809 1984
rect 837 1944 849 2024
rect 865 1944 877 2024
rect 931 1944 943 1984
rect 951 1944 963 1984
rect 971 1944 983 1984
rect 997 1952 1009 1992
rect 1017 1952 1029 1992
rect 1047 1952 1059 2016
rect 1077 1944 1089 2024
rect 1121 1944 1133 2024
rect 1141 1944 1153 1984
rect 1175 1944 1187 1984
rect 1207 1944 1219 1984
rect 1227 1944 1239 1984
rect 1253 1944 1265 1984
rect 1281 1944 1293 1964
rect 1311 1944 1323 1964
rect 1331 1944 1343 2024
rect 1357 1944 1369 1984
rect 1377 1944 1389 1984
rect 1417 1944 1429 2024
rect 1447 1944 1469 2024
rect 1487 1944 1499 2024
rect 1556 1944 1568 1984
rect 1578 1944 1590 2024
rect 1606 1944 1618 2024
rect 1656 1944 1668 1984
rect 1678 1944 1690 2024
rect 1706 1944 1718 2024
rect 1763 1944 1775 2024
rect 1791 1944 1803 2024
rect 1836 1944 1848 1984
rect 1858 1944 1870 2024
rect 1886 1944 1898 2024
rect 1931 1944 1943 2024
rect 1961 1952 1973 2016
rect 1991 1952 2003 1992
rect 2011 1952 2023 1992
rect 2051 1944 2063 2024
rect 2081 1952 2093 2016
rect 2111 1952 2123 1992
rect 2131 1952 2143 1992
rect 2161 1944 2173 2024
rect 2181 1944 2193 1984
rect 2215 1944 2227 1984
rect 2247 1944 2259 1984
rect 2267 1944 2279 1984
rect 2293 1944 2305 1984
rect 2321 1944 2333 1964
rect 2351 1944 2363 1964
rect 2371 1944 2383 2024
rect 2416 1944 2428 1984
rect 2438 1944 2450 2024
rect 2466 1944 2478 2024
rect 2497 1944 2509 2024
rect 2525 1944 2537 2024
rect 2591 1944 2603 1984
rect 2611 1944 2623 1980
rect 2631 1944 2643 1984
rect 2651 1944 2663 1984
rect 2677 1952 2689 1992
rect 2697 1952 2709 1992
rect 2727 1952 2739 2016
rect 2757 1944 2769 2024
rect 2811 1944 2823 2024
rect 2841 1952 2853 2016
rect 2871 1952 2883 1992
rect 2891 1952 2903 1992
rect 2917 1944 2929 1984
rect 2937 1944 2949 1984
rect 2977 1944 2989 2024
rect 3007 1944 3029 2024
rect 3047 1944 3059 2024
rect 3111 1944 3123 2024
rect 3131 1944 3143 2024
rect 3151 1944 3163 2012
rect 3171 1944 3183 2016
rect 3197 1944 3209 1984
rect 3217 1944 3229 1984
rect 3257 1944 3269 2024
rect 3287 1944 3309 2024
rect 3327 1944 3339 2024
rect 3377 1944 3389 2024
rect 3405 1944 3417 2024
rect 3461 1944 3473 2024
rect 3481 1944 3493 1984
rect 3515 1944 3527 1984
rect 3547 1944 3559 1984
rect 3567 1944 3579 1984
rect 3593 1944 3605 1984
rect 3621 1944 3633 1964
rect 3651 1944 3663 1964
rect 3671 1944 3683 2024
rect 3723 1944 3735 2024
rect 3751 1944 3763 2024
rect 3801 1944 3813 2024
rect 3831 1944 3853 2024
rect 3871 1944 3883 2024
rect 3911 1944 3923 1984
rect 3931 1944 3943 1984
rect 3962 1944 3974 2024
rect 3990 1944 4002 2024
rect 4012 1944 4024 1984
rect 4057 1944 4069 1984
rect 4077 1944 4089 1984
rect 4097 1944 4109 1984
rect 4163 1944 4175 2024
rect 4191 1944 4203 2024
rect 4221 1944 4233 2024
rect 4241 1944 4253 1984
rect 4275 1944 4287 1984
rect 4307 1944 4319 1984
rect 4327 1944 4339 1984
rect 4353 1944 4365 1984
rect 4381 1944 4393 1964
rect 4411 1944 4423 1964
rect 4431 1944 4443 2024
rect 4457 1944 4469 1984
rect 4477 1944 4489 1984
rect 4517 1944 4529 2024
rect 4547 1944 4569 2024
rect 4587 1944 4599 2024
rect 4637 1944 4649 2024
rect 4665 1944 4677 2024
rect 4736 1944 4748 1984
rect 4758 1944 4770 2024
rect 4786 1944 4798 2024
rect 4843 1944 4855 2024
rect 4871 1944 4883 2024
rect 4897 1944 4909 2024
rect 4927 1944 4949 2024
rect 4967 1944 4979 2024
rect 5031 1944 5043 1984
rect 5051 1944 5063 1984
rect 5071 1944 5083 1984
rect 5123 1944 5135 2024
rect 5151 1944 5163 2024
rect 5177 1944 5189 2024
rect 5207 1944 5219 2023
rect 5227 1944 5239 2023
rect 5301 1944 5313 2024
rect 5331 1944 5353 2024
rect 5371 1944 5383 2024
rect 5397 1944 5409 2024
rect 5427 1944 5449 2024
rect 5467 1944 5479 2024
rect 5543 1944 5555 2024
rect 5571 1944 5583 2024
rect 5621 1944 5633 2024
rect 5651 1944 5673 2024
rect 5691 1944 5703 2024
rect 5731 1944 5743 1984
rect 5751 1944 5763 1984
rect 5777 1944 5789 1984
rect 5797 1944 5809 1984
rect 5817 1944 5829 1984
rect 5857 1944 5869 2024
rect 5877 1944 5889 1964
rect 5907 1944 5919 1964
rect 5935 1944 5947 1984
rect 5961 1944 5973 1984
rect 5981 1944 5993 1984
rect 6013 1944 6025 1984
rect 6047 1944 6059 1984
rect 6067 1944 6079 2024
rect 6101 1944 6113 2024
rect 6121 1944 6133 1984
rect 6155 1944 6167 1984
rect 6187 1944 6199 1984
rect 6207 1944 6219 1984
rect 6233 1944 6245 1984
rect 6261 1944 6273 1964
rect 6291 1944 6303 1964
rect 6311 1944 6323 2024
rect 6337 1952 6349 1992
rect 6357 1952 6369 1992
rect 6387 1952 6399 2016
rect 6417 1944 6429 2024
rect 6457 1944 6469 2016
rect 6477 1944 6489 2012
rect 6497 1944 6509 2024
rect 6517 1944 6529 2024
rect 6562 1944 6574 2024
rect 6590 1944 6602 2024
rect 6612 1944 6624 1984
rect 31 1876 43 1916
rect 51 1876 63 1916
rect 77 1836 89 1916
rect 97 1896 109 1916
rect 127 1896 139 1916
rect 155 1876 167 1916
rect 181 1876 193 1916
rect 201 1876 213 1916
rect 233 1876 245 1916
rect 267 1876 279 1916
rect 287 1836 299 1916
rect 317 1836 329 1916
rect 345 1836 357 1916
rect 423 1836 435 1916
rect 451 1836 463 1916
rect 491 1876 503 1916
rect 511 1876 523 1916
rect 556 1876 568 1916
rect 578 1836 590 1916
rect 606 1836 618 1916
rect 637 1836 649 1916
rect 657 1896 669 1916
rect 687 1896 699 1916
rect 715 1876 727 1916
rect 741 1876 753 1916
rect 761 1876 773 1916
rect 793 1876 805 1916
rect 827 1876 839 1916
rect 847 1836 859 1916
rect 891 1876 903 1916
rect 911 1880 923 1916
rect 931 1876 943 1916
rect 951 1876 963 1916
rect 977 1876 989 1916
rect 997 1876 1009 1916
rect 1021 1836 1033 1916
rect 1041 1836 1053 1916
rect 1077 1876 1089 1916
rect 1097 1876 1109 1916
rect 1142 1836 1154 1916
rect 1170 1836 1182 1916
rect 1192 1876 1204 1916
rect 1251 1876 1263 1916
rect 1271 1876 1283 1916
rect 1291 1876 1303 1916
rect 1331 1876 1343 1916
rect 1351 1880 1363 1916
rect 1371 1876 1383 1916
rect 1391 1876 1403 1916
rect 1417 1876 1429 1916
rect 1437 1876 1449 1916
rect 1481 1836 1493 1916
rect 1501 1876 1513 1916
rect 1535 1876 1547 1916
rect 1567 1876 1579 1916
rect 1587 1876 1599 1916
rect 1613 1876 1625 1916
rect 1641 1896 1653 1916
rect 1671 1896 1683 1916
rect 1691 1836 1703 1916
rect 1717 1876 1729 1916
rect 1737 1876 1749 1916
rect 1777 1836 1789 1916
rect 1807 1836 1829 1916
rect 1847 1836 1859 1916
rect 1897 1836 1909 1916
rect 1925 1836 1937 1916
rect 1982 1836 1994 1916
rect 2010 1836 2022 1916
rect 2032 1876 2044 1916
rect 2077 1836 2089 1916
rect 2097 1896 2109 1916
rect 2127 1896 2139 1916
rect 2155 1876 2167 1916
rect 2181 1876 2193 1916
rect 2201 1876 2213 1916
rect 2233 1876 2245 1916
rect 2267 1876 2279 1916
rect 2287 1836 2299 1916
rect 2341 1836 2353 1916
rect 2371 1836 2393 1916
rect 2411 1836 2423 1916
rect 2437 1876 2449 1916
rect 2457 1876 2469 1916
rect 2497 1836 2509 1916
rect 2525 1836 2537 1916
rect 2577 1836 2589 1916
rect 2597 1896 2609 1916
rect 2627 1896 2639 1916
rect 2655 1876 2667 1916
rect 2681 1876 2693 1916
rect 2701 1876 2713 1916
rect 2733 1876 2745 1916
rect 2767 1876 2779 1916
rect 2787 1836 2799 1916
rect 2817 1876 2829 1916
rect 2837 1876 2849 1916
rect 2857 1880 2869 1916
rect 2877 1876 2889 1916
rect 2936 1876 2948 1916
rect 2958 1836 2970 1916
rect 2986 1836 2998 1916
rect 3017 1836 3029 1916
rect 3045 1836 3057 1916
rect 3111 1836 3123 1916
rect 3131 1836 3143 1916
rect 3151 1848 3163 1916
rect 3171 1844 3183 1916
rect 3211 1836 3223 1916
rect 3231 1836 3243 1916
rect 3251 1848 3263 1916
rect 3271 1844 3283 1916
rect 3309 1836 3321 1916
rect 3329 1836 3341 1916
rect 3351 1876 3363 1916
rect 3391 1876 3403 1916
rect 3411 1876 3423 1916
rect 3431 1876 3443 1916
rect 3457 1836 3469 1916
rect 3485 1836 3497 1916
rect 3537 1876 3549 1916
rect 3557 1876 3569 1916
rect 3577 1876 3589 1916
rect 3622 1836 3634 1916
rect 3650 1836 3662 1916
rect 3672 1876 3684 1916
rect 3731 1876 3743 1916
rect 3751 1876 3763 1916
rect 3771 1876 3783 1916
rect 3811 1876 3823 1916
rect 3831 1876 3843 1916
rect 3857 1876 3869 1916
rect 3877 1876 3889 1916
rect 3897 1876 3909 1916
rect 3937 1836 3949 1916
rect 3965 1836 3977 1916
rect 4017 1836 4029 1916
rect 4047 1836 4069 1916
rect 4087 1836 4099 1916
rect 4163 1836 4175 1916
rect 4191 1836 4203 1916
rect 4222 1836 4234 1916
rect 4250 1836 4262 1916
rect 4272 1876 4284 1916
rect 4317 1836 4329 1914
rect 4337 1836 4349 1916
rect 4357 1836 4369 1916
rect 4402 1836 4414 1916
rect 4430 1836 4442 1916
rect 4452 1876 4464 1916
rect 4523 1836 4535 1916
rect 4551 1836 4563 1916
rect 4601 1836 4613 1916
rect 4631 1836 4653 1916
rect 4671 1836 4683 1916
rect 4711 1876 4723 1916
rect 4731 1876 4743 1916
rect 4757 1836 4769 1916
rect 4777 1896 4789 1916
rect 4807 1896 4819 1916
rect 4835 1876 4847 1916
rect 4861 1876 4873 1916
rect 4881 1876 4893 1916
rect 4913 1876 4925 1916
rect 4947 1876 4959 1916
rect 4967 1836 4979 1916
rect 4997 1844 5009 1916
rect 5017 1848 5029 1916
rect 5037 1836 5049 1916
rect 5057 1836 5069 1916
rect 5097 1836 5109 1916
rect 5125 1836 5137 1916
rect 5182 1836 5194 1916
rect 5210 1836 5222 1916
rect 5232 1876 5244 1916
rect 5277 1876 5289 1916
rect 5297 1876 5309 1916
rect 5317 1880 5329 1916
rect 5337 1876 5349 1916
rect 5377 1876 5389 1916
rect 5399 1836 5411 1916
rect 5419 1836 5431 1916
rect 5471 1876 5483 1916
rect 5491 1876 5503 1916
rect 5531 1836 5543 1916
rect 5551 1836 5563 1916
rect 5596 1876 5608 1916
rect 5618 1836 5630 1916
rect 5646 1836 5658 1916
rect 5677 1876 5689 1916
rect 5697 1876 5709 1916
rect 5717 1876 5729 1916
rect 5771 1836 5783 1916
rect 5791 1836 5803 1904
rect 5811 1838 5823 1916
rect 5831 1850 5843 1916
rect 5851 1838 5863 1916
rect 5877 1876 5889 1916
rect 5899 1836 5911 1916
rect 5919 1836 5931 1916
rect 5976 1876 5988 1916
rect 5998 1836 6010 1916
rect 6026 1836 6038 1916
rect 6081 1836 6093 1916
rect 6111 1836 6133 1916
rect 6151 1836 6163 1916
rect 6177 1868 6189 1908
rect 6197 1868 6209 1908
rect 6227 1844 6239 1908
rect 6257 1836 6269 1916
rect 6297 1868 6309 1908
rect 6317 1868 6329 1908
rect 6347 1844 6359 1908
rect 6377 1836 6389 1916
rect 6417 1876 6429 1916
rect 6437 1876 6449 1916
rect 6482 1836 6494 1916
rect 6510 1836 6522 1916
rect 6532 1876 6544 1916
rect 6591 1876 6603 1916
rect 6611 1876 6623 1916
rect 6631 1876 6643 1916
rect 43 1464 55 1544
rect 71 1464 83 1544
rect 111 1464 123 1544
rect 131 1464 143 1544
rect 151 1464 163 1544
rect 171 1464 183 1544
rect 191 1464 203 1544
rect 211 1464 223 1544
rect 231 1464 243 1544
rect 251 1464 263 1544
rect 271 1464 283 1544
rect 301 1464 313 1544
rect 321 1464 333 1504
rect 355 1464 367 1504
rect 387 1464 399 1504
rect 407 1464 419 1504
rect 433 1464 445 1504
rect 461 1464 473 1484
rect 491 1464 503 1484
rect 511 1464 523 1544
rect 551 1464 563 1504
rect 571 1464 583 1504
rect 597 1464 609 1504
rect 617 1464 629 1504
rect 637 1464 649 1500
rect 657 1464 669 1504
rect 697 1464 709 1536
rect 717 1464 729 1532
rect 737 1464 749 1544
rect 757 1464 769 1544
rect 801 1464 813 1544
rect 821 1464 833 1504
rect 855 1464 867 1504
rect 887 1464 899 1504
rect 907 1464 919 1504
rect 933 1464 945 1504
rect 961 1464 973 1484
rect 991 1464 1003 1484
rect 1011 1464 1023 1544
rect 1051 1464 1063 1504
rect 1071 1464 1083 1504
rect 1097 1464 1109 1544
rect 1127 1464 1149 1544
rect 1167 1464 1179 1544
rect 1236 1464 1248 1504
rect 1258 1464 1270 1544
rect 1286 1464 1298 1544
rect 1343 1464 1355 1544
rect 1371 1464 1383 1544
rect 1411 1464 1423 1544
rect 1441 1472 1453 1536
rect 1471 1472 1483 1512
rect 1491 1472 1503 1512
rect 1531 1464 1543 1544
rect 1561 1472 1573 1536
rect 1591 1472 1603 1512
rect 1611 1472 1623 1512
rect 1651 1464 1663 1544
rect 1681 1472 1693 1536
rect 1711 1472 1723 1512
rect 1731 1472 1743 1512
rect 1757 1464 1769 1544
rect 1777 1464 1789 1484
rect 1807 1464 1819 1484
rect 1835 1464 1847 1504
rect 1861 1464 1873 1504
rect 1881 1464 1893 1504
rect 1913 1464 1925 1504
rect 1947 1464 1959 1504
rect 1967 1464 1979 1544
rect 1997 1472 2009 1512
rect 2017 1472 2029 1512
rect 2047 1472 2059 1536
rect 2077 1464 2089 1544
rect 2117 1464 2129 1504
rect 2137 1464 2149 1504
rect 2177 1464 2189 1544
rect 2207 1464 2229 1544
rect 2247 1464 2259 1544
rect 2297 1464 2309 1544
rect 2325 1464 2337 1544
rect 2396 1464 2408 1504
rect 2418 1464 2430 1544
rect 2446 1464 2458 1544
rect 2489 1464 2501 1544
rect 2509 1464 2521 1544
rect 2531 1464 2543 1504
rect 2557 1464 2569 1544
rect 2585 1464 2597 1544
rect 2651 1464 2663 1504
rect 2671 1464 2683 1504
rect 2691 1464 2703 1504
rect 2717 1464 2729 1504
rect 2737 1464 2749 1504
rect 2757 1464 2769 1504
rect 2811 1464 2823 1544
rect 2841 1472 2853 1536
rect 2871 1472 2883 1512
rect 2891 1472 2903 1512
rect 2931 1464 2943 1504
rect 2951 1464 2963 1500
rect 2971 1464 2983 1504
rect 2991 1464 3003 1504
rect 3031 1464 3043 1544
rect 3051 1464 3063 1544
rect 3081 1464 3093 1544
rect 3101 1464 3113 1504
rect 3135 1464 3147 1504
rect 3167 1464 3179 1504
rect 3187 1464 3199 1504
rect 3213 1464 3225 1504
rect 3241 1464 3253 1484
rect 3271 1464 3283 1484
rect 3291 1464 3303 1544
rect 3331 1464 3343 1504
rect 3351 1464 3363 1504
rect 3371 1464 3383 1504
rect 3416 1464 3428 1504
rect 3438 1464 3450 1544
rect 3466 1464 3478 1544
rect 3497 1464 3509 1542
rect 3517 1464 3529 1530
rect 3537 1464 3549 1542
rect 3557 1476 3569 1544
rect 3577 1464 3589 1544
rect 3636 1464 3648 1504
rect 3658 1464 3670 1544
rect 3686 1464 3698 1544
rect 3731 1464 3743 1504
rect 3751 1464 3763 1504
rect 3803 1464 3815 1544
rect 3831 1464 3843 1544
rect 3881 1464 3893 1544
rect 3911 1464 3933 1544
rect 3951 1464 3963 1544
rect 3991 1464 4003 1504
rect 4011 1464 4023 1504
rect 4041 1464 4053 1544
rect 4061 1464 4073 1504
rect 4095 1464 4107 1504
rect 4127 1464 4139 1504
rect 4147 1464 4159 1504
rect 4173 1464 4185 1504
rect 4201 1464 4213 1484
rect 4231 1464 4243 1484
rect 4251 1464 4263 1544
rect 4291 1464 4303 1544
rect 4321 1472 4333 1536
rect 4351 1472 4363 1512
rect 4371 1472 4383 1512
rect 4411 1464 4423 1544
rect 4441 1472 4453 1536
rect 4471 1472 4483 1512
rect 4491 1472 4503 1512
rect 4517 1472 4529 1512
rect 4537 1472 4549 1512
rect 4567 1472 4579 1536
rect 4597 1464 4609 1544
rect 4637 1472 4649 1512
rect 4657 1472 4669 1512
rect 4687 1472 4699 1536
rect 4717 1464 4729 1544
rect 4757 1472 4769 1512
rect 4777 1472 4789 1512
rect 4807 1472 4819 1536
rect 4837 1464 4849 1544
rect 4877 1472 4889 1512
rect 4897 1472 4909 1512
rect 4927 1472 4939 1536
rect 4957 1464 4969 1544
rect 4997 1464 5009 1544
rect 5017 1464 5029 1484
rect 5047 1464 5059 1484
rect 5075 1464 5087 1504
rect 5101 1464 5113 1504
rect 5121 1464 5133 1504
rect 5153 1464 5165 1504
rect 5187 1464 5199 1504
rect 5207 1464 5219 1544
rect 5237 1464 5249 1544
rect 5257 1464 5269 1484
rect 5287 1464 5299 1484
rect 5315 1464 5327 1504
rect 5341 1464 5353 1504
rect 5361 1464 5373 1504
rect 5393 1464 5405 1504
rect 5427 1464 5439 1504
rect 5447 1464 5459 1544
rect 5477 1464 5489 1542
rect 5497 1464 5509 1530
rect 5517 1464 5529 1542
rect 5537 1476 5549 1544
rect 5557 1464 5569 1544
rect 5597 1472 5609 1512
rect 5617 1472 5629 1512
rect 5647 1472 5659 1536
rect 5677 1464 5689 1544
rect 5736 1464 5748 1504
rect 5758 1464 5770 1544
rect 5786 1464 5798 1544
rect 5843 1464 5855 1544
rect 5871 1464 5883 1544
rect 5911 1464 5923 1504
rect 5931 1464 5943 1504
rect 5951 1464 5963 1504
rect 5996 1464 6008 1504
rect 6018 1464 6030 1544
rect 6046 1464 6058 1544
rect 6103 1464 6115 1544
rect 6131 1464 6143 1544
rect 6181 1464 6193 1544
rect 6211 1464 6233 1544
rect 6251 1464 6263 1544
rect 6291 1464 6303 1544
rect 6321 1472 6333 1536
rect 6351 1472 6363 1512
rect 6371 1472 6383 1512
rect 6397 1464 6409 1504
rect 6417 1464 6429 1504
rect 6457 1464 6469 1544
rect 6477 1464 6489 1484
rect 6507 1464 6519 1484
rect 6535 1464 6547 1504
rect 6561 1464 6573 1504
rect 6581 1464 6593 1504
rect 6613 1464 6625 1504
rect 6647 1464 6659 1504
rect 6667 1464 6679 1544
rect 17 1396 29 1436
rect 37 1396 49 1436
rect 61 1356 73 1436
rect 81 1356 93 1436
rect 117 1356 129 1436
rect 145 1356 157 1436
rect 216 1396 228 1436
rect 238 1356 250 1436
rect 266 1356 278 1436
rect 323 1356 335 1436
rect 351 1356 363 1436
rect 377 1396 389 1436
rect 397 1396 409 1436
rect 437 1396 449 1436
rect 457 1396 469 1436
rect 511 1396 523 1436
rect 531 1396 543 1436
rect 551 1396 563 1436
rect 577 1364 589 1436
rect 597 1368 609 1436
rect 617 1356 629 1436
rect 637 1356 649 1436
rect 681 1356 693 1436
rect 701 1396 713 1436
rect 735 1396 747 1436
rect 767 1396 779 1436
rect 787 1396 799 1436
rect 813 1396 825 1436
rect 841 1416 853 1436
rect 871 1416 883 1436
rect 891 1356 903 1436
rect 931 1396 943 1436
rect 951 1396 963 1436
rect 971 1396 983 1436
rect 997 1396 1009 1436
rect 1017 1396 1029 1436
rect 1037 1400 1049 1436
rect 1057 1396 1069 1436
rect 1097 1356 1109 1436
rect 1125 1356 1137 1436
rect 1181 1356 1193 1436
rect 1201 1396 1213 1436
rect 1235 1396 1247 1436
rect 1267 1396 1279 1436
rect 1287 1396 1299 1436
rect 1313 1396 1325 1436
rect 1341 1416 1353 1436
rect 1371 1416 1383 1436
rect 1391 1356 1403 1436
rect 1431 1356 1443 1436
rect 1451 1356 1463 1436
rect 1471 1356 1483 1436
rect 1491 1356 1503 1436
rect 1511 1356 1523 1436
rect 1531 1356 1543 1436
rect 1551 1356 1563 1436
rect 1571 1356 1583 1436
rect 1591 1356 1603 1436
rect 1631 1356 1643 1436
rect 1661 1364 1673 1428
rect 1691 1388 1703 1428
rect 1711 1388 1723 1428
rect 1763 1356 1775 1436
rect 1791 1356 1803 1436
rect 1841 1356 1853 1436
rect 1871 1356 1893 1436
rect 1911 1356 1923 1436
rect 1956 1396 1968 1436
rect 1978 1356 1990 1436
rect 2006 1356 2018 1436
rect 2037 1396 2049 1436
rect 2057 1396 2069 1436
rect 2102 1356 2114 1436
rect 2130 1356 2142 1436
rect 2152 1396 2164 1436
rect 2197 1396 2209 1436
rect 2217 1396 2229 1436
rect 2237 1396 2249 1436
rect 2277 1388 2289 1428
rect 2297 1388 2309 1428
rect 2327 1364 2339 1428
rect 2357 1356 2369 1436
rect 2411 1356 2423 1436
rect 2441 1364 2453 1428
rect 2471 1388 2483 1428
rect 2491 1388 2503 1428
rect 2531 1356 2543 1436
rect 2551 1356 2563 1424
rect 2571 1358 2583 1436
rect 2591 1370 2603 1436
rect 2611 1358 2623 1436
rect 2637 1358 2649 1436
rect 2657 1370 2669 1436
rect 2677 1358 2689 1436
rect 2697 1356 2709 1424
rect 2717 1356 2729 1436
rect 2771 1356 2783 1436
rect 2791 1356 2803 1424
rect 2811 1358 2823 1436
rect 2831 1370 2843 1436
rect 2851 1358 2863 1436
rect 2877 1396 2889 1436
rect 2899 1356 2911 1436
rect 2919 1356 2931 1436
rect 2971 1356 2983 1436
rect 2991 1356 3003 1424
rect 3011 1358 3023 1436
rect 3031 1370 3043 1436
rect 3051 1358 3063 1436
rect 3091 1396 3103 1436
rect 3111 1396 3123 1436
rect 3151 1356 3163 1436
rect 3181 1364 3193 1428
rect 3211 1388 3223 1428
rect 3231 1388 3243 1428
rect 3261 1356 3273 1436
rect 3281 1396 3293 1436
rect 3315 1396 3327 1436
rect 3347 1396 3359 1436
rect 3367 1396 3379 1436
rect 3393 1396 3405 1436
rect 3421 1416 3433 1436
rect 3451 1416 3463 1436
rect 3471 1356 3483 1436
rect 3523 1356 3535 1436
rect 3551 1356 3563 1436
rect 3601 1356 3613 1436
rect 3631 1356 3653 1436
rect 3671 1356 3683 1436
rect 3716 1396 3728 1436
rect 3738 1356 3750 1436
rect 3766 1356 3778 1436
rect 3811 1396 3823 1436
rect 3831 1396 3843 1436
rect 3857 1356 3869 1436
rect 3877 1416 3889 1436
rect 3907 1416 3919 1436
rect 3935 1396 3947 1436
rect 3961 1396 3973 1436
rect 3981 1396 3993 1436
rect 4013 1396 4025 1436
rect 4047 1396 4059 1436
rect 4067 1356 4079 1436
rect 4097 1356 4109 1436
rect 4117 1416 4129 1436
rect 4147 1416 4159 1436
rect 4175 1396 4187 1436
rect 4201 1396 4213 1436
rect 4221 1396 4233 1436
rect 4253 1396 4265 1436
rect 4287 1396 4299 1436
rect 4307 1356 4319 1436
rect 4351 1396 4363 1436
rect 4371 1396 4383 1436
rect 4397 1358 4409 1436
rect 4417 1370 4429 1436
rect 4437 1358 4449 1436
rect 4457 1356 4469 1424
rect 4477 1356 4489 1436
rect 4517 1388 4529 1428
rect 4537 1388 4549 1428
rect 4567 1364 4579 1428
rect 4597 1356 4609 1436
rect 4651 1356 4663 1436
rect 4671 1356 4683 1424
rect 4691 1358 4703 1436
rect 4711 1370 4723 1436
rect 4731 1358 4743 1436
rect 4769 1356 4781 1436
rect 4789 1356 4801 1436
rect 4811 1396 4823 1436
rect 4851 1396 4863 1436
rect 4871 1396 4883 1436
rect 4891 1396 4903 1436
rect 4931 1396 4943 1436
rect 4951 1396 4963 1436
rect 4971 1396 4983 1436
rect 5021 1356 5033 1436
rect 5051 1356 5073 1436
rect 5091 1356 5103 1436
rect 5141 1356 5153 1436
rect 5171 1356 5193 1436
rect 5211 1356 5223 1436
rect 5237 1356 5249 1436
rect 5257 1356 5269 1436
rect 5311 1396 5323 1436
rect 5331 1396 5343 1436
rect 5351 1396 5363 1436
rect 5377 1356 5389 1436
rect 5407 1356 5429 1436
rect 5447 1356 5459 1436
rect 5511 1356 5523 1436
rect 5531 1356 5543 1436
rect 5551 1368 5563 1436
rect 5571 1364 5583 1436
rect 5597 1356 5609 1436
rect 5617 1356 5629 1436
rect 5657 1388 5669 1428
rect 5677 1388 5689 1428
rect 5707 1364 5719 1428
rect 5737 1356 5749 1436
rect 5791 1396 5803 1436
rect 5811 1396 5823 1436
rect 5831 1396 5843 1436
rect 5876 1396 5888 1436
rect 5898 1356 5910 1436
rect 5926 1356 5938 1436
rect 5971 1396 5983 1436
rect 5991 1396 6003 1436
rect 6022 1356 6034 1436
rect 6050 1356 6062 1436
rect 6072 1396 6084 1436
rect 6117 1356 6129 1436
rect 6147 1356 6169 1436
rect 6187 1356 6199 1436
rect 6237 1356 6249 1436
rect 6257 1416 6269 1436
rect 6287 1416 6299 1436
rect 6315 1396 6327 1436
rect 6341 1396 6353 1436
rect 6361 1396 6373 1436
rect 6393 1396 6405 1436
rect 6427 1396 6439 1436
rect 6447 1356 6459 1436
rect 6477 1356 6489 1436
rect 6497 1416 6509 1436
rect 6527 1416 6539 1436
rect 6555 1396 6567 1436
rect 6581 1396 6593 1436
rect 6601 1396 6613 1436
rect 6633 1396 6645 1436
rect 6667 1396 6679 1436
rect 6687 1356 6699 1436
rect 17 984 29 1064
rect 37 984 49 1004
rect 67 984 79 1004
rect 95 984 107 1024
rect 121 984 133 1024
rect 141 984 153 1024
rect 173 984 185 1024
rect 207 984 219 1024
rect 227 984 239 1064
rect 271 984 283 1024
rect 291 984 303 1024
rect 317 984 329 1064
rect 337 984 349 1004
rect 367 984 379 1004
rect 395 984 407 1024
rect 421 984 433 1024
rect 441 984 453 1024
rect 473 984 485 1024
rect 507 984 519 1024
rect 527 984 539 1064
rect 557 984 569 1024
rect 577 984 589 1024
rect 617 984 629 1024
rect 637 984 649 1024
rect 657 984 669 1020
rect 677 984 689 1024
rect 717 984 729 1064
rect 745 984 757 1064
rect 797 984 809 1024
rect 817 984 829 1024
rect 837 984 849 1020
rect 857 984 869 1024
rect 897 984 909 1024
rect 917 984 929 1024
rect 937 984 949 1024
rect 977 984 989 1024
rect 997 984 1009 1024
rect 1041 984 1053 1064
rect 1061 984 1073 1024
rect 1095 984 1107 1024
rect 1127 984 1139 1024
rect 1147 984 1159 1024
rect 1173 984 1185 1024
rect 1201 984 1213 1004
rect 1231 984 1243 1004
rect 1251 984 1263 1064
rect 1277 984 1289 1064
rect 1297 984 1309 1064
rect 1317 984 1329 1064
rect 1337 984 1349 1064
rect 1357 984 1369 1064
rect 1377 984 1389 1064
rect 1397 984 1409 1064
rect 1417 984 1429 1064
rect 1437 984 1449 1064
rect 1481 984 1493 1064
rect 1501 984 1513 1024
rect 1535 984 1547 1024
rect 1567 984 1579 1024
rect 1587 984 1599 1024
rect 1613 984 1625 1024
rect 1641 984 1653 1004
rect 1671 984 1683 1004
rect 1691 984 1703 1064
rect 1743 984 1755 1064
rect 1771 984 1783 1064
rect 1821 984 1833 1064
rect 1851 984 1873 1064
rect 1891 984 1903 1064
rect 1936 984 1948 1024
rect 1958 984 1970 1064
rect 1986 984 1998 1064
rect 2036 984 2048 1024
rect 2058 984 2070 1064
rect 2086 984 2098 1064
rect 2143 984 2155 1064
rect 2171 984 2183 1064
rect 2221 984 2233 1064
rect 2251 984 2273 1064
rect 2291 984 2303 1064
rect 2321 984 2333 1064
rect 2341 984 2353 1024
rect 2375 984 2387 1024
rect 2407 984 2419 1024
rect 2427 984 2439 1024
rect 2453 984 2465 1024
rect 2481 984 2493 1004
rect 2511 984 2523 1004
rect 2531 984 2543 1064
rect 2571 984 2583 1024
rect 2591 984 2603 1024
rect 2622 984 2634 1064
rect 2650 984 2662 1064
rect 2672 984 2684 1024
rect 2729 984 2741 1064
rect 2749 984 2761 1064
rect 2771 984 2783 1024
rect 2797 984 2809 1024
rect 2817 984 2829 1024
rect 2871 984 2883 1064
rect 2891 996 2903 1064
rect 2911 984 2923 1062
rect 2931 984 2943 1050
rect 2951 984 2963 1062
rect 2981 984 2993 1064
rect 3001 984 3013 1024
rect 3035 984 3047 1024
rect 3067 984 3079 1024
rect 3087 984 3099 1024
rect 3113 984 3125 1024
rect 3141 984 3153 1004
rect 3171 984 3183 1004
rect 3191 984 3203 1064
rect 3217 984 3229 1024
rect 3237 984 3249 1024
rect 3257 984 3269 1024
rect 3311 984 3323 1064
rect 3341 992 3353 1056
rect 3371 992 3383 1032
rect 3391 992 3403 1032
rect 3417 992 3429 1032
rect 3437 992 3449 1032
rect 3467 992 3479 1056
rect 3497 984 3509 1064
rect 3549 984 3561 1064
rect 3569 984 3581 1064
rect 3591 984 3603 1024
rect 3621 984 3633 1064
rect 3641 984 3653 1024
rect 3675 984 3687 1024
rect 3707 984 3719 1024
rect 3727 984 3739 1024
rect 3753 984 3765 1024
rect 3781 984 3793 1004
rect 3811 984 3823 1004
rect 3831 984 3843 1064
rect 3857 992 3869 1032
rect 3877 992 3889 1032
rect 3907 992 3919 1056
rect 3937 984 3949 1064
rect 3991 984 4003 1064
rect 4021 992 4033 1056
rect 4051 992 4063 1032
rect 4071 992 4083 1032
rect 4097 984 4109 1024
rect 4117 984 4129 1024
rect 4157 984 4169 1064
rect 4187 984 4209 1064
rect 4227 984 4239 1064
rect 4277 984 4289 1064
rect 4305 984 4317 1064
rect 4376 984 4388 1024
rect 4398 984 4410 1064
rect 4426 984 4438 1064
rect 4471 984 4483 1064
rect 4491 984 4503 1064
rect 4511 984 4523 1052
rect 4531 984 4543 1056
rect 4561 984 4573 1064
rect 4581 984 4593 1024
rect 4615 984 4627 1024
rect 4647 984 4659 1024
rect 4667 984 4679 1024
rect 4693 984 4705 1024
rect 4721 984 4733 1004
rect 4751 984 4763 1004
rect 4771 984 4783 1064
rect 4797 984 4809 1064
rect 4827 984 4849 1064
rect 4867 984 4879 1064
rect 4943 984 4955 1064
rect 4971 984 4983 1064
rect 5016 984 5028 1024
rect 5038 984 5050 1064
rect 5066 984 5078 1064
rect 5123 984 5135 1064
rect 5151 984 5163 1064
rect 5177 984 5189 1064
rect 5205 984 5217 1064
rect 5257 984 5269 1064
rect 5285 984 5297 1064
rect 5349 984 5361 1064
rect 5369 984 5381 1064
rect 5391 984 5403 1024
rect 5417 984 5429 1064
rect 5445 984 5457 1064
rect 5497 984 5509 1064
rect 5525 984 5537 1064
rect 5577 984 5589 1056
rect 5597 984 5609 1052
rect 5617 984 5629 1064
rect 5637 984 5649 1064
rect 5677 984 5689 1064
rect 5707 984 5719 1063
rect 5727 984 5739 1063
rect 5803 984 5815 1064
rect 5831 984 5843 1064
rect 5862 984 5874 1064
rect 5890 984 5902 1064
rect 5912 984 5924 1024
rect 5971 984 5983 1024
rect 5991 984 6003 1020
rect 6011 984 6023 1024
rect 6031 984 6043 1024
rect 6062 984 6074 1064
rect 6090 984 6102 1064
rect 6112 984 6124 1024
rect 6183 984 6195 1064
rect 6211 984 6223 1064
rect 6237 984 6249 1064
rect 6265 984 6277 1064
rect 6317 984 6329 1064
rect 6337 984 6349 1004
rect 6367 984 6379 1004
rect 6395 984 6407 1024
rect 6421 984 6433 1024
rect 6441 984 6453 1024
rect 6473 984 6485 1024
rect 6507 984 6519 1024
rect 6527 984 6539 1064
rect 6557 984 6569 1064
rect 6587 984 6609 1064
rect 6627 984 6639 1064
rect 17 876 29 956
rect 47 877 59 956
rect 67 877 79 956
rect 131 916 143 956
rect 151 916 163 956
rect 171 916 183 956
rect 197 876 209 956
rect 217 936 229 956
rect 247 936 259 956
rect 275 916 287 956
rect 301 916 313 956
rect 321 916 333 956
rect 353 916 365 956
rect 387 916 399 956
rect 407 876 419 956
rect 451 916 463 956
rect 471 916 483 956
rect 523 876 535 956
rect 551 876 563 956
rect 577 876 589 956
rect 605 876 617 956
rect 657 916 669 956
rect 677 916 689 956
rect 697 916 709 956
rect 737 916 749 956
rect 757 916 769 956
rect 777 920 789 956
rect 797 916 809 956
rect 837 876 849 956
rect 867 876 889 956
rect 907 876 919 956
rect 962 876 974 956
rect 990 876 1002 956
rect 1012 916 1024 956
rect 1062 876 1074 956
rect 1090 876 1102 956
rect 1112 916 1124 956
rect 1167 888 1179 948
rect 1187 892 1199 944
rect 1207 888 1219 948
rect 1231 898 1243 956
rect 1251 896 1263 944
rect 1271 896 1283 956
rect 1291 896 1303 956
rect 1311 896 1323 956
rect 1342 876 1354 956
rect 1370 876 1382 956
rect 1392 916 1404 956
rect 1451 916 1463 956
rect 1471 916 1483 956
rect 1501 876 1513 956
rect 1521 916 1533 956
rect 1555 916 1567 956
rect 1587 916 1599 956
rect 1607 916 1619 956
rect 1633 916 1645 956
rect 1661 936 1673 956
rect 1691 936 1703 956
rect 1711 876 1723 956
rect 1737 916 1749 956
rect 1757 916 1769 956
rect 1797 908 1809 948
rect 1817 908 1829 948
rect 1847 884 1859 948
rect 1877 876 1889 956
rect 1922 876 1934 956
rect 1950 876 1962 956
rect 1972 916 1984 956
rect 2017 916 2029 956
rect 2037 916 2049 956
rect 2057 916 2069 956
rect 2097 876 2109 956
rect 2117 936 2129 956
rect 2147 936 2159 956
rect 2175 916 2187 956
rect 2201 916 2213 956
rect 2221 916 2233 956
rect 2253 916 2265 956
rect 2287 916 2299 956
rect 2307 876 2319 956
rect 2337 916 2349 956
rect 2357 916 2369 956
rect 2397 876 2409 956
rect 2427 876 2449 956
rect 2467 876 2479 956
rect 2517 876 2529 956
rect 2545 876 2557 956
rect 2616 916 2628 956
rect 2638 876 2650 956
rect 2666 876 2678 956
rect 2711 876 2723 956
rect 2731 876 2743 956
rect 2751 876 2763 956
rect 2771 876 2783 956
rect 2791 876 2803 956
rect 2811 876 2823 956
rect 2831 876 2843 956
rect 2851 876 2863 956
rect 2871 876 2883 956
rect 2897 884 2909 956
rect 2917 888 2929 956
rect 2937 876 2949 956
rect 2957 876 2969 956
rect 3011 876 3023 956
rect 3031 876 3043 956
rect 3051 888 3063 956
rect 3071 884 3083 956
rect 3111 876 3123 956
rect 3141 884 3153 948
rect 3171 908 3183 948
rect 3191 908 3203 948
rect 3231 876 3243 956
rect 3261 884 3273 948
rect 3291 908 3303 948
rect 3311 908 3323 948
rect 3356 916 3368 956
rect 3378 876 3390 956
rect 3406 876 3418 956
rect 3437 916 3449 956
rect 3457 916 3469 956
rect 3477 916 3489 956
rect 3517 908 3529 948
rect 3537 908 3549 948
rect 3567 884 3579 948
rect 3597 876 3609 956
rect 3651 916 3663 956
rect 3671 916 3683 956
rect 3711 876 3723 956
rect 3741 884 3753 948
rect 3771 908 3783 948
rect 3791 908 3803 948
rect 3821 876 3833 956
rect 3841 916 3853 956
rect 3875 916 3887 956
rect 3907 916 3919 956
rect 3927 916 3939 956
rect 3953 916 3965 956
rect 3981 936 3993 956
rect 4011 936 4023 956
rect 4031 876 4043 956
rect 4057 908 4069 948
rect 4077 908 4089 948
rect 4107 884 4119 948
rect 4137 876 4149 956
rect 4177 884 4189 956
rect 4197 888 4209 956
rect 4217 876 4229 956
rect 4237 876 4249 956
rect 4282 876 4294 956
rect 4310 876 4322 956
rect 4332 916 4344 956
rect 4391 916 4403 956
rect 4411 920 4423 956
rect 4431 916 4443 956
rect 4451 916 4463 956
rect 4477 916 4489 956
rect 4497 916 4509 956
rect 4542 876 4554 956
rect 4570 876 4582 956
rect 4592 916 4604 956
rect 4637 916 4649 956
rect 4657 916 4669 956
rect 4677 916 4689 956
rect 4731 916 4743 956
rect 4751 916 4763 956
rect 4782 876 4794 956
rect 4810 876 4822 956
rect 4832 916 4844 956
rect 4877 916 4889 956
rect 4897 916 4909 956
rect 4917 916 4929 956
rect 4957 908 4969 948
rect 4977 908 4989 948
rect 5007 884 5019 948
rect 5037 876 5049 956
rect 5091 876 5103 956
rect 5121 884 5133 948
rect 5151 908 5163 948
rect 5171 908 5183 948
rect 5197 876 5209 956
rect 5217 876 5229 956
rect 5237 876 5249 956
rect 5257 876 5269 956
rect 5277 876 5289 956
rect 5297 876 5309 956
rect 5317 876 5329 956
rect 5337 876 5349 956
rect 5357 876 5369 956
rect 5397 884 5409 956
rect 5417 888 5429 956
rect 5437 876 5449 956
rect 5457 876 5469 956
rect 5511 916 5523 956
rect 5531 916 5543 956
rect 5562 876 5574 956
rect 5590 876 5602 956
rect 5612 916 5624 956
rect 5657 916 5669 956
rect 5677 916 5689 956
rect 5697 916 5709 956
rect 5742 876 5754 956
rect 5770 876 5782 956
rect 5792 916 5804 956
rect 5851 916 5863 956
rect 5871 920 5883 956
rect 5891 916 5903 956
rect 5911 916 5923 956
rect 5941 876 5953 956
rect 5961 916 5973 956
rect 5995 916 6007 956
rect 6027 916 6039 956
rect 6047 916 6059 956
rect 6073 916 6085 956
rect 6101 936 6113 956
rect 6131 936 6143 956
rect 6151 876 6163 956
rect 6182 876 6194 956
rect 6210 876 6222 956
rect 6232 916 6244 956
rect 6282 876 6294 956
rect 6310 876 6322 956
rect 6332 916 6344 956
rect 6391 916 6403 956
rect 6411 916 6423 956
rect 6431 916 6443 956
rect 6461 876 6473 956
rect 6481 916 6493 956
rect 6515 916 6527 956
rect 6547 916 6559 956
rect 6567 916 6579 956
rect 6593 916 6605 956
rect 6621 936 6633 956
rect 6651 936 6663 956
rect 6671 876 6683 956
rect 17 504 29 544
rect 37 504 49 544
rect 77 504 89 544
rect 97 504 109 544
rect 117 504 129 544
rect 157 504 169 576
rect 177 504 189 572
rect 197 504 209 584
rect 217 504 229 584
rect 257 504 269 544
rect 277 504 289 544
rect 331 504 343 584
rect 351 504 363 584
rect 371 504 383 572
rect 391 504 403 576
rect 417 504 429 544
rect 437 504 449 544
rect 457 504 469 540
rect 477 504 489 544
rect 531 504 543 544
rect 551 504 563 544
rect 571 504 583 544
rect 611 504 623 544
rect 631 504 643 540
rect 651 504 663 544
rect 671 504 683 544
rect 697 504 709 544
rect 717 504 729 544
rect 757 504 769 544
rect 777 504 789 544
rect 843 504 855 584
rect 871 504 883 584
rect 907 512 919 572
rect 927 516 939 568
rect 947 512 959 572
rect 971 504 983 562
rect 991 516 1003 564
rect 1011 504 1023 564
rect 1031 504 1043 564
rect 1051 504 1063 564
rect 1081 504 1093 584
rect 1101 504 1113 544
rect 1135 504 1147 544
rect 1167 504 1179 544
rect 1187 504 1199 544
rect 1213 504 1225 544
rect 1241 504 1253 524
rect 1271 504 1283 524
rect 1291 504 1303 584
rect 1317 504 1329 544
rect 1339 504 1351 584
rect 1359 504 1371 584
rect 1397 504 1409 544
rect 1417 504 1429 544
rect 1437 504 1449 544
rect 1481 504 1493 584
rect 1501 504 1513 544
rect 1535 504 1547 544
rect 1567 504 1579 544
rect 1587 504 1599 544
rect 1613 504 1625 544
rect 1641 504 1653 524
rect 1671 504 1683 524
rect 1691 504 1703 584
rect 1721 504 1733 584
rect 1741 504 1753 544
rect 1775 504 1787 544
rect 1807 504 1819 544
rect 1827 504 1839 544
rect 1853 504 1865 544
rect 1881 504 1893 524
rect 1911 504 1923 524
rect 1931 504 1943 584
rect 1961 504 1973 584
rect 1981 504 1993 544
rect 2015 504 2027 544
rect 2047 504 2059 544
rect 2067 504 2079 544
rect 2093 504 2105 544
rect 2121 504 2133 524
rect 2151 504 2163 524
rect 2171 504 2183 584
rect 2201 504 2213 584
rect 2221 504 2233 544
rect 2255 504 2267 544
rect 2287 504 2299 544
rect 2307 504 2319 544
rect 2333 504 2345 544
rect 2361 504 2373 524
rect 2391 504 2403 524
rect 2411 504 2423 584
rect 2437 504 2449 584
rect 2457 504 2469 524
rect 2487 504 2499 524
rect 2515 504 2527 544
rect 2541 504 2553 544
rect 2561 504 2573 544
rect 2593 504 2605 544
rect 2627 504 2639 544
rect 2647 504 2659 584
rect 2691 504 2703 584
rect 2711 516 2723 584
rect 2731 504 2743 582
rect 2751 504 2763 570
rect 2771 504 2783 582
rect 2811 504 2823 544
rect 2831 504 2843 544
rect 2871 504 2883 584
rect 2891 504 2903 584
rect 2911 504 2923 572
rect 2931 504 2943 576
rect 2957 504 2969 544
rect 2977 504 2989 544
rect 3022 504 3034 584
rect 3050 504 3062 584
rect 3072 504 3084 544
rect 3117 504 3129 544
rect 3137 504 3149 544
rect 3157 504 3169 544
rect 3197 504 3209 544
rect 3217 504 3229 544
rect 3237 504 3249 540
rect 3257 504 3269 544
rect 3297 504 3309 544
rect 3317 504 3329 544
rect 3362 504 3374 584
rect 3390 504 3402 584
rect 3412 504 3424 544
rect 3457 504 3469 544
rect 3477 504 3489 544
rect 3497 504 3509 544
rect 3537 504 3549 576
rect 3557 504 3569 572
rect 3577 504 3589 584
rect 3597 504 3609 584
rect 3637 504 3649 584
rect 3665 504 3677 584
rect 3722 504 3734 584
rect 3750 504 3762 584
rect 3772 504 3784 544
rect 3831 504 3843 544
rect 3851 504 3863 540
rect 3871 504 3883 544
rect 3891 504 3903 544
rect 3917 504 3929 584
rect 3937 504 3949 524
rect 3967 504 3979 524
rect 3995 504 4007 544
rect 4021 504 4033 544
rect 4041 504 4053 544
rect 4073 504 4085 544
rect 4107 504 4119 544
rect 4127 504 4139 584
rect 4183 504 4195 584
rect 4211 504 4223 584
rect 4237 504 4249 584
rect 4257 504 4269 524
rect 4287 504 4299 524
rect 4315 504 4327 544
rect 4341 504 4353 544
rect 4361 504 4373 544
rect 4393 504 4405 544
rect 4427 504 4439 544
rect 4447 504 4459 584
rect 4477 504 4489 544
rect 4497 504 4509 544
rect 4537 504 4549 582
rect 4557 504 4569 570
rect 4577 504 4589 582
rect 4597 516 4609 584
rect 4617 504 4629 584
rect 4671 504 4683 584
rect 4691 504 4703 584
rect 4711 504 4723 572
rect 4731 504 4743 576
rect 4776 504 4788 544
rect 4798 504 4810 584
rect 4826 504 4838 584
rect 4857 504 4869 544
rect 4877 504 4889 544
rect 4897 504 4909 544
rect 4951 504 4963 544
rect 4971 504 4983 544
rect 5011 504 5023 584
rect 5041 512 5053 576
rect 5071 512 5083 552
rect 5091 512 5103 552
rect 5117 504 5129 544
rect 5137 504 5149 544
rect 5157 504 5169 540
rect 5177 504 5189 544
rect 5217 504 5229 584
rect 5237 504 5249 524
rect 5267 504 5279 524
rect 5295 504 5307 544
rect 5321 504 5333 544
rect 5341 504 5353 544
rect 5373 504 5385 544
rect 5407 504 5419 544
rect 5427 504 5439 584
rect 5457 504 5469 584
rect 5477 504 5489 584
rect 5517 512 5529 552
rect 5537 512 5549 552
rect 5567 512 5579 576
rect 5597 504 5609 584
rect 5663 504 5675 584
rect 5691 504 5703 584
rect 5743 504 5755 584
rect 5771 504 5783 584
rect 5823 504 5835 584
rect 5851 504 5863 584
rect 5877 504 5889 584
rect 5905 504 5917 584
rect 5983 504 5995 584
rect 6011 504 6023 584
rect 6042 504 6054 584
rect 6070 504 6082 584
rect 6092 504 6104 544
rect 6142 504 6154 584
rect 6170 504 6182 584
rect 6192 504 6204 544
rect 6251 504 6263 544
rect 6271 504 6283 544
rect 6291 504 6303 544
rect 6321 504 6333 584
rect 6341 504 6353 544
rect 6375 504 6387 544
rect 6407 504 6419 544
rect 6427 504 6439 544
rect 6453 504 6465 544
rect 6481 504 6493 524
rect 6511 504 6523 524
rect 6531 504 6543 584
rect 6557 504 6569 544
rect 6577 504 6589 544
rect 6617 504 6629 544
rect 6637 504 6649 544
rect 17 396 29 476
rect 37 456 49 476
rect 67 456 79 476
rect 95 436 107 476
rect 121 436 133 476
rect 141 436 153 476
rect 173 436 185 476
rect 207 436 219 476
rect 227 396 239 476
rect 261 396 273 476
rect 281 436 293 476
rect 315 436 327 476
rect 347 436 359 476
rect 367 436 379 476
rect 393 436 405 476
rect 421 456 433 476
rect 451 456 463 476
rect 471 396 483 476
rect 497 436 509 476
rect 517 436 529 476
rect 537 440 549 476
rect 557 436 569 476
rect 597 396 609 476
rect 625 396 637 476
rect 703 396 715 476
rect 731 396 743 476
rect 757 436 769 476
rect 777 436 789 476
rect 797 436 809 476
rect 851 436 863 476
rect 871 436 883 476
rect 901 396 913 476
rect 921 436 933 476
rect 955 436 967 476
rect 987 436 999 476
rect 1007 436 1019 476
rect 1033 436 1045 476
rect 1061 456 1073 476
rect 1091 456 1103 476
rect 1111 396 1123 476
rect 1149 396 1161 476
rect 1169 396 1181 476
rect 1191 436 1203 476
rect 1217 436 1229 476
rect 1239 396 1251 476
rect 1259 396 1271 476
rect 1297 436 1309 476
rect 1319 396 1331 476
rect 1339 396 1351 476
rect 1391 436 1403 476
rect 1411 436 1423 476
rect 1442 396 1454 476
rect 1470 396 1482 476
rect 1492 436 1504 476
rect 1551 436 1563 476
rect 1571 436 1583 476
rect 1602 396 1614 476
rect 1630 396 1642 476
rect 1652 436 1664 476
rect 1701 396 1713 476
rect 1721 436 1733 476
rect 1755 436 1767 476
rect 1787 436 1799 476
rect 1807 436 1819 476
rect 1833 436 1845 476
rect 1861 456 1873 476
rect 1891 456 1903 476
rect 1911 396 1923 476
rect 1951 436 1963 476
rect 1971 436 1983 476
rect 2011 436 2023 476
rect 2031 436 2043 476
rect 2062 396 2074 476
rect 2090 396 2102 476
rect 2112 436 2124 476
rect 2157 436 2169 476
rect 2177 436 2189 476
rect 2217 396 2229 476
rect 2247 396 2269 476
rect 2287 396 2299 476
rect 2356 436 2368 476
rect 2378 396 2390 476
rect 2406 396 2418 476
rect 2437 396 2449 476
rect 2465 396 2477 476
rect 2521 396 2533 476
rect 2541 436 2553 476
rect 2575 436 2587 476
rect 2607 436 2619 476
rect 2627 436 2639 476
rect 2653 436 2665 476
rect 2681 456 2693 476
rect 2711 456 2723 476
rect 2731 396 2743 476
rect 2776 436 2788 476
rect 2798 396 2810 476
rect 2826 396 2838 476
rect 2857 396 2869 476
rect 2885 396 2897 476
rect 2941 396 2953 476
rect 2961 436 2973 476
rect 2995 436 3007 476
rect 3027 436 3039 476
rect 3047 436 3059 476
rect 3073 436 3085 476
rect 3101 456 3113 476
rect 3131 456 3143 476
rect 3151 396 3163 476
rect 3177 436 3189 476
rect 3197 436 3209 476
rect 3217 436 3229 476
rect 3276 436 3288 476
rect 3298 396 3310 476
rect 3326 396 3338 476
rect 3357 396 3369 476
rect 3385 396 3397 476
rect 3451 396 3463 476
rect 3471 396 3483 476
rect 3491 408 3503 476
rect 3511 404 3523 476
rect 3542 396 3554 476
rect 3570 396 3582 476
rect 3592 436 3604 476
rect 3637 396 3649 476
rect 3665 396 3677 476
rect 3717 404 3729 476
rect 3737 408 3749 476
rect 3757 396 3769 476
rect 3777 396 3789 476
rect 3843 396 3855 476
rect 3871 396 3883 476
rect 3902 396 3914 476
rect 3930 396 3942 476
rect 3952 436 3964 476
rect 4011 436 4023 476
rect 4031 440 4043 476
rect 4051 436 4063 476
rect 4071 436 4083 476
rect 4097 396 4109 476
rect 4125 396 4137 476
rect 4177 396 4189 476
rect 4197 456 4209 476
rect 4227 456 4239 476
rect 4255 436 4267 476
rect 4281 436 4293 476
rect 4301 436 4313 476
rect 4333 436 4345 476
rect 4367 436 4379 476
rect 4387 396 4399 476
rect 4417 396 4429 476
rect 4445 396 4457 476
rect 4516 436 4528 476
rect 4538 396 4550 476
rect 4566 396 4578 476
rect 4597 396 4609 476
rect 4625 396 4637 476
rect 4701 396 4713 476
rect 4731 396 4753 476
rect 4771 396 4783 476
rect 4811 436 4823 476
rect 4831 436 4843 476
rect 4861 396 4873 476
rect 4881 436 4893 476
rect 4915 436 4927 476
rect 4947 436 4959 476
rect 4967 436 4979 476
rect 4993 436 5005 476
rect 5021 456 5033 476
rect 5051 456 5063 476
rect 5071 396 5083 476
rect 5111 396 5123 476
rect 5131 396 5143 476
rect 5151 408 5163 476
rect 5171 404 5183 476
rect 5197 396 5209 476
rect 5225 396 5237 476
rect 5296 436 5308 476
rect 5318 396 5330 476
rect 5346 396 5358 476
rect 5377 396 5389 476
rect 5405 396 5417 476
rect 5457 404 5469 476
rect 5477 408 5489 476
rect 5497 396 5509 476
rect 5517 396 5529 476
rect 5557 436 5569 476
rect 5577 436 5589 476
rect 5597 440 5609 476
rect 5617 436 5629 476
rect 5662 396 5674 476
rect 5690 396 5702 476
rect 5712 436 5724 476
rect 5771 436 5783 476
rect 5791 436 5803 476
rect 5811 436 5823 476
rect 5856 436 5868 476
rect 5878 396 5890 476
rect 5906 396 5918 476
rect 5942 396 5954 476
rect 5970 396 5982 476
rect 5992 436 6004 476
rect 6042 396 6054 476
rect 6070 396 6082 476
rect 6092 436 6104 476
rect 6163 396 6175 476
rect 6191 396 6203 476
rect 6243 396 6255 476
rect 6271 396 6283 476
rect 6321 396 6333 476
rect 6351 396 6373 476
rect 6391 396 6403 476
rect 6421 396 6433 476
rect 6441 436 6453 476
rect 6475 436 6487 476
rect 6507 436 6519 476
rect 6527 436 6539 476
rect 6553 436 6565 476
rect 6581 456 6593 476
rect 6611 456 6623 476
rect 6631 396 6643 476
rect 17 24 29 104
rect 37 24 49 44
rect 67 24 79 44
rect 95 24 107 64
rect 121 24 133 64
rect 141 24 153 64
rect 173 24 185 64
rect 207 24 219 64
rect 227 24 239 104
rect 257 24 269 104
rect 277 24 289 44
rect 307 24 319 44
rect 335 24 347 64
rect 361 24 373 64
rect 381 24 393 64
rect 413 24 425 64
rect 447 24 459 64
rect 467 24 479 104
rect 509 24 521 104
rect 529 24 541 104
rect 551 24 563 64
rect 577 24 589 64
rect 599 24 611 104
rect 619 24 631 104
rect 669 24 681 104
rect 689 24 701 104
rect 711 24 723 64
rect 737 24 749 104
rect 757 24 769 44
rect 787 24 799 44
rect 815 24 827 64
rect 841 24 853 64
rect 861 24 873 64
rect 893 24 905 64
rect 927 24 939 64
rect 947 24 959 104
rect 977 24 989 64
rect 999 24 1011 104
rect 1019 24 1031 104
rect 1071 24 1083 64
rect 1091 24 1103 64
rect 1111 24 1123 64
rect 1156 24 1168 64
rect 1178 24 1190 104
rect 1206 24 1218 104
rect 1241 24 1253 104
rect 1261 24 1273 64
rect 1295 24 1307 64
rect 1327 24 1339 64
rect 1347 24 1359 64
rect 1373 24 1385 64
rect 1401 24 1413 44
rect 1431 24 1443 44
rect 1451 24 1463 104
rect 1491 24 1503 64
rect 1511 24 1523 64
rect 1537 24 1549 64
rect 1557 24 1569 64
rect 1577 24 1589 64
rect 1636 24 1648 64
rect 1658 24 1670 104
rect 1686 24 1698 104
rect 1717 24 1729 64
rect 1737 24 1749 64
rect 1777 24 1789 64
rect 1797 24 1809 64
rect 1817 24 1829 64
rect 1857 24 1869 64
rect 1877 24 1889 64
rect 1897 24 1909 64
rect 1937 24 1949 64
rect 1957 24 1969 64
rect 1977 24 1989 64
rect 2036 24 2048 64
rect 2058 24 2070 104
rect 2086 24 2098 104
rect 2121 24 2133 104
rect 2141 24 2153 64
rect 2175 24 2187 64
rect 2207 24 2219 64
rect 2227 24 2239 64
rect 2253 24 2265 64
rect 2281 24 2293 44
rect 2311 24 2323 44
rect 2331 24 2343 104
rect 2357 24 2369 64
rect 2377 24 2389 64
rect 2397 24 2409 64
rect 2451 24 2463 64
rect 2471 24 2483 64
rect 2491 24 2503 64
rect 2536 24 2548 64
rect 2558 24 2570 104
rect 2586 24 2598 104
rect 2631 24 2643 64
rect 2651 24 2663 64
rect 2681 24 2693 104
rect 2701 24 2713 64
rect 2735 24 2747 64
rect 2767 24 2779 64
rect 2787 24 2799 64
rect 2813 24 2825 64
rect 2841 24 2853 44
rect 2871 24 2883 44
rect 2891 24 2903 104
rect 2936 24 2948 64
rect 2958 24 2970 104
rect 2986 24 2998 104
rect 3043 24 3055 104
rect 3071 24 3083 104
rect 3121 24 3133 104
rect 3151 24 3173 104
rect 3191 24 3203 104
rect 3231 24 3243 64
rect 3251 24 3263 64
rect 3277 24 3289 104
rect 3297 24 3309 44
rect 3327 24 3339 44
rect 3355 24 3367 64
rect 3381 24 3393 64
rect 3401 24 3413 64
rect 3433 24 3445 64
rect 3467 24 3479 64
rect 3487 24 3499 104
rect 3531 24 3543 64
rect 3551 24 3563 64
rect 3571 24 3583 64
rect 3616 24 3628 64
rect 3638 24 3650 104
rect 3666 24 3678 104
rect 3702 24 3714 104
rect 3730 24 3742 104
rect 3752 24 3764 64
rect 3797 24 3809 104
rect 3817 24 3829 44
rect 3847 24 3859 44
rect 3875 24 3887 64
rect 3901 24 3913 64
rect 3921 24 3933 64
rect 3953 24 3965 64
rect 3987 24 3999 64
rect 4007 24 4019 104
rect 4042 24 4054 104
rect 4070 24 4082 104
rect 4092 24 4104 64
rect 4142 24 4154 104
rect 4170 24 4182 104
rect 4192 24 4204 64
rect 4237 24 4249 64
rect 4257 24 4269 64
rect 4277 24 4289 64
rect 4317 24 4329 104
rect 4337 24 4349 44
rect 4367 24 4379 44
rect 4395 24 4407 64
rect 4421 24 4433 64
rect 4441 24 4453 64
rect 4473 24 4485 64
rect 4507 24 4519 64
rect 4527 24 4539 104
rect 4562 24 4574 104
rect 4590 24 4602 104
rect 4612 24 4624 64
rect 4662 24 4674 104
rect 4690 24 4702 104
rect 4712 24 4724 64
rect 4757 24 4769 64
rect 4777 24 4789 64
rect 4797 24 4809 64
rect 4837 24 4849 104
rect 4857 24 4869 44
rect 4887 24 4899 44
rect 4915 24 4927 64
rect 4941 24 4953 64
rect 4961 24 4973 64
rect 4993 24 5005 64
rect 5027 24 5039 64
rect 5047 24 5059 104
rect 5096 24 5108 64
rect 5118 24 5130 104
rect 5146 24 5158 104
rect 5182 24 5194 104
rect 5210 24 5222 104
rect 5232 24 5244 64
rect 5277 24 5289 64
rect 5297 24 5309 64
rect 5317 24 5329 64
rect 5357 24 5369 104
rect 5377 24 5389 44
rect 5407 24 5419 44
rect 5435 24 5447 64
rect 5461 24 5473 64
rect 5481 24 5493 64
rect 5513 24 5525 64
rect 5547 24 5559 64
rect 5567 24 5579 104
rect 5597 24 5609 104
rect 5617 24 5629 44
rect 5647 24 5659 44
rect 5675 24 5687 64
rect 5701 24 5713 64
rect 5721 24 5733 64
rect 5753 24 5765 64
rect 5787 24 5799 64
rect 5807 24 5819 104
rect 5837 24 5849 104
rect 5857 24 5869 44
rect 5887 24 5899 44
rect 5915 24 5927 64
rect 5941 24 5953 64
rect 5961 24 5973 64
rect 5993 24 6005 64
rect 6027 24 6039 64
rect 6047 24 6059 104
rect 6091 24 6103 104
rect 6111 24 6123 104
rect 6142 24 6154 104
rect 6170 24 6182 104
rect 6192 24 6204 64
rect 6261 24 6273 104
rect 6291 24 6313 104
rect 6331 24 6343 104
rect 6371 24 6383 64
rect 6391 24 6403 64
rect 6417 24 6429 104
rect 6437 24 6449 44
rect 6467 24 6479 44
rect 6495 24 6507 64
rect 6521 24 6533 64
rect 6541 24 6553 64
rect 6573 24 6585 64
rect 6607 24 6619 64
rect 6627 24 6639 104
<< psubstratepcontact >>
rect 4 6484 6736 6496
rect 4 6004 6736 6016
rect 4 5524 6736 5536
rect 4 5044 6736 5056
rect 4 4564 6736 4576
rect 4 4084 6736 4096
rect 4 3604 6736 3616
rect 4 3124 6736 3136
rect 4 2644 6736 2656
rect 4 2164 6736 2176
rect 4 1684 6736 1696
rect 4 1204 6736 1216
rect 4 724 6736 736
rect 4 244 6736 256
<< nsubstratencontact >>
rect 4 6244 6736 6256
rect 4 5764 6736 5776
rect 4 5284 6736 5296
rect 4 4804 6736 4816
rect 4 4324 6736 4336
rect 4 3844 6736 3856
rect 4 3364 6736 3376
rect 4 2884 6736 2896
rect 4 2404 6736 2416
rect 4 1924 6736 1936
rect 4 1444 6736 1456
rect 4 964 6736 976
rect 4 484 6736 496
rect 4 4 6736 16
<< polysilicon >>
rect 35 6476 39 6480
rect 55 6476 59 6480
rect 65 6476 69 6480
rect 87 6476 91 6480
rect 97 6476 101 6480
rect 119 6476 123 6480
rect 165 6476 169 6480
rect 173 6476 177 6480
rect 193 6476 197 6480
rect 203 6476 207 6480
rect 225 6476 229 6480
rect 285 6476 289 6480
rect 305 6476 309 6480
rect 325 6476 329 6480
rect 373 6476 377 6480
rect 383 6476 387 6480
rect 473 6476 477 6480
rect 483 6476 487 6480
rect 533 6476 537 6480
rect 543 6476 547 6480
rect 611 6476 615 6480
rect 633 6476 637 6480
rect 643 6476 647 6480
rect 663 6476 667 6480
rect 671 6476 675 6480
rect 717 6476 721 6480
rect 739 6476 743 6480
rect 749 6476 753 6480
rect 771 6476 775 6480
rect 781 6476 785 6480
rect 801 6476 805 6480
rect 851 6476 855 6480
rect 914 6476 918 6480
rect 922 6476 926 6480
rect 942 6476 946 6480
rect 950 6476 954 6480
rect 1045 6476 1049 6480
rect 1091 6476 1095 6480
rect 1113 6476 1117 6480
rect 1123 6476 1127 6480
rect 1143 6476 1147 6480
rect 1151 6476 1155 6480
rect 1197 6476 1201 6480
rect 1219 6476 1223 6480
rect 1229 6476 1233 6480
rect 1251 6476 1255 6480
rect 1261 6476 1265 6480
rect 1281 6476 1285 6480
rect 1331 6476 1335 6480
rect 1351 6476 1355 6480
rect 1371 6476 1375 6480
rect 1391 6476 1395 6480
rect 1465 6476 1469 6480
rect 1485 6476 1489 6480
rect 1505 6476 1509 6480
rect 1575 6476 1579 6480
rect 1595 6476 1599 6480
rect 1605 6476 1609 6480
rect 1665 6476 1669 6480
rect 1711 6476 1715 6480
rect 1733 6476 1737 6480
rect 1743 6476 1747 6480
rect 1763 6476 1767 6480
rect 1771 6476 1775 6480
rect 1817 6476 1821 6480
rect 1839 6476 1843 6480
rect 1849 6476 1853 6480
rect 1871 6476 1875 6480
rect 1881 6476 1885 6480
rect 1901 6476 1905 6480
rect 1951 6476 1955 6480
rect 1971 6476 1975 6480
rect 1991 6476 1995 6480
rect 2053 6476 2057 6480
rect 2063 6476 2067 6480
rect 2145 6476 2149 6480
rect 2165 6476 2169 6480
rect 2185 6476 2189 6480
rect 2252 6476 2256 6480
rect 2274 6476 2278 6480
rect 2282 6476 2286 6480
rect 2353 6476 2357 6480
rect 2363 6476 2367 6480
rect 2425 6476 2429 6480
rect 2445 6476 2449 6480
rect 2491 6476 2495 6480
rect 2511 6476 2515 6480
rect 2573 6476 2577 6480
rect 2583 6476 2587 6480
rect 2688 6476 2692 6480
rect 2696 6476 2700 6480
rect 2704 6476 2708 6480
rect 2753 6476 2757 6480
rect 2763 6476 2767 6480
rect 2868 6476 2872 6480
rect 2876 6476 2880 6480
rect 2884 6476 2888 6480
rect 2945 6476 2949 6480
rect 2965 6476 2969 6480
rect 2985 6476 2989 6480
rect 3045 6476 3049 6480
rect 3065 6476 3069 6480
rect 3085 6476 3089 6480
rect 3145 6476 3149 6480
rect 3205 6476 3209 6480
rect 3254 6476 3258 6480
rect 3262 6476 3266 6480
rect 3284 6476 3288 6480
rect 3351 6476 3355 6480
rect 3371 6476 3375 6480
rect 3391 6476 3395 6480
rect 3472 6476 3476 6480
rect 3494 6476 3498 6480
rect 3502 6476 3506 6480
rect 3572 6476 3576 6480
rect 3594 6476 3598 6480
rect 3602 6476 3606 6480
rect 3652 6476 3656 6480
rect 3660 6476 3664 6480
rect 3668 6476 3672 6480
rect 3765 6476 3769 6480
rect 3785 6476 3789 6480
rect 3805 6476 3809 6480
rect 3851 6476 3855 6480
rect 3871 6476 3875 6480
rect 3891 6476 3895 6480
rect 3951 6476 3955 6480
rect 4013 6476 4017 6480
rect 4023 6476 4027 6480
rect 4115 6476 4119 6480
rect 4135 6476 4139 6480
rect 4145 6476 4149 6480
rect 4193 6476 4197 6480
rect 4203 6476 4207 6480
rect 4308 6476 4312 6480
rect 4316 6476 4320 6480
rect 4324 6476 4328 6480
rect 4408 6476 4412 6480
rect 4416 6476 4420 6480
rect 4424 6476 4428 6480
rect 4508 6476 4512 6480
rect 4516 6476 4520 6480
rect 4524 6476 4528 6480
rect 4571 6476 4575 6480
rect 4634 6476 4638 6480
rect 4642 6476 4646 6480
rect 4664 6476 4668 6480
rect 4734 6476 4738 6480
rect 4742 6476 4746 6480
rect 4764 6476 4768 6480
rect 4831 6476 4835 6480
rect 4851 6476 4855 6480
rect 4871 6476 4875 6480
rect 4945 6476 4949 6480
rect 4965 6476 4969 6480
rect 4985 6476 4989 6480
rect 5031 6476 5035 6480
rect 5051 6476 5055 6480
rect 5071 6476 5075 6480
rect 5168 6476 5172 6480
rect 5176 6476 5180 6480
rect 5184 6476 5188 6480
rect 5268 6476 5272 6480
rect 5276 6476 5280 6480
rect 5284 6476 5288 6480
rect 5368 6476 5372 6480
rect 5376 6476 5380 6480
rect 5384 6476 5388 6480
rect 5434 6476 5438 6480
rect 5442 6476 5446 6480
rect 5464 6476 5468 6480
rect 5552 6476 5556 6480
rect 5574 6476 5578 6480
rect 5582 6476 5586 6480
rect 5645 6476 5649 6480
rect 5694 6476 5698 6480
rect 5702 6476 5706 6480
rect 5724 6476 5728 6480
rect 5792 6476 5796 6480
rect 5800 6476 5804 6480
rect 5808 6476 5812 6480
rect 5912 6476 5916 6480
rect 5934 6476 5938 6480
rect 5942 6476 5946 6480
rect 6005 6476 6009 6480
rect 6072 6476 6076 6480
rect 6094 6476 6098 6480
rect 6102 6476 6106 6480
rect 6165 6476 6169 6480
rect 6185 6476 6189 6480
rect 6205 6476 6209 6480
rect 6272 6476 6276 6480
rect 6294 6476 6298 6480
rect 6302 6476 6306 6480
rect 6352 6476 6356 6480
rect 6360 6476 6364 6480
rect 6368 6476 6372 6480
rect 6488 6476 6492 6480
rect 6496 6476 6500 6480
rect 6504 6476 6508 6480
rect 6551 6476 6555 6480
rect 6614 6476 6618 6480
rect 6622 6476 6626 6480
rect 6642 6476 6646 6480
rect 6650 6476 6654 6480
rect 35 6399 39 6436
rect 55 6398 59 6456
rect 65 6424 69 6456
rect 87 6444 91 6456
rect 89 6432 91 6444
rect 97 6444 101 6456
rect 97 6432 99 6444
rect 65 6420 98 6424
rect 35 6344 39 6387
rect 55 6304 59 6386
rect 74 6371 78 6400
rect 69 6363 78 6371
rect 69 6304 73 6363
rect 94 6356 98 6420
rect 95 6344 98 6356
rect 89 6304 93 6344
rect 103 6322 107 6432
rect 119 6342 123 6456
rect 165 6452 169 6456
rect 135 6448 169 6452
rect 101 6304 105 6310
rect 121 6304 125 6330
rect 135 6322 139 6448
rect 173 6444 177 6456
rect 147 6440 177 6444
rect 159 6439 177 6440
rect 193 6435 197 6456
rect 173 6431 197 6435
rect 173 6336 179 6431
rect 203 6407 207 6456
rect 203 6349 207 6395
rect 225 6368 229 6436
rect 227 6356 229 6368
rect 285 6359 289 6436
rect 305 6413 309 6436
rect 325 6431 329 6436
rect 325 6424 338 6431
rect 305 6401 314 6413
rect 203 6343 211 6349
rect 225 6344 229 6356
rect 287 6347 294 6359
rect 147 6310 171 6312
rect 135 6308 171 6310
rect 167 6304 171 6308
rect 175 6304 179 6336
rect 195 6284 199 6324
rect 207 6314 211 6343
rect 203 6307 211 6314
rect 203 6284 207 6307
rect 290 6304 294 6347
rect 312 6344 316 6401
rect 334 6379 338 6424
rect 373 6416 377 6436
rect 369 6409 377 6416
rect 383 6416 387 6436
rect 473 6416 477 6436
rect 383 6409 397 6416
rect 369 6393 375 6409
rect 366 6381 375 6393
rect 334 6356 338 6367
rect 320 6348 338 6356
rect 320 6344 324 6348
rect 371 6304 375 6381
rect 391 6393 397 6409
rect 463 6409 477 6416
rect 483 6416 487 6436
rect 533 6416 537 6436
rect 483 6409 491 6416
rect 463 6393 469 6409
rect 391 6381 394 6393
rect 466 6381 469 6393
rect 391 6304 395 6381
rect 465 6304 469 6381
rect 485 6393 491 6409
rect 529 6409 537 6416
rect 543 6416 547 6436
rect 543 6409 557 6416
rect 529 6393 535 6409
rect 485 6381 494 6393
rect 526 6381 535 6393
rect 485 6304 489 6381
rect 531 6304 535 6381
rect 551 6393 557 6409
rect 551 6381 554 6393
rect 551 6304 555 6381
rect 611 6368 615 6436
rect 633 6407 637 6456
rect 643 6435 647 6456
rect 663 6444 667 6456
rect 671 6452 675 6456
rect 671 6448 705 6452
rect 663 6440 693 6444
rect 663 6439 681 6440
rect 643 6431 667 6435
rect 611 6356 613 6368
rect 611 6344 615 6356
rect 633 6349 637 6395
rect 629 6343 637 6349
rect 629 6314 633 6343
rect 661 6336 667 6431
rect 629 6307 637 6314
rect 633 6284 637 6307
rect 641 6284 645 6324
rect 661 6304 665 6336
rect 701 6322 705 6448
rect 717 6342 721 6456
rect 739 6444 743 6456
rect 741 6432 743 6444
rect 749 6444 753 6456
rect 749 6432 751 6444
rect 669 6310 693 6312
rect 669 6308 705 6310
rect 669 6304 673 6308
rect 715 6304 719 6330
rect 733 6322 737 6432
rect 771 6424 775 6456
rect 742 6420 775 6424
rect 742 6356 746 6420
rect 762 6371 766 6400
rect 781 6398 785 6456
rect 801 6399 805 6436
rect 851 6399 855 6456
rect 914 6428 918 6436
rect 846 6387 855 6399
rect 762 6363 771 6371
rect 742 6344 745 6356
rect 735 6304 739 6310
rect 747 6304 751 6344
rect 767 6304 771 6363
rect 781 6304 785 6386
rect 801 6344 805 6387
rect 851 6304 855 6387
rect 901 6421 918 6428
rect 901 6379 907 6421
rect 922 6413 926 6436
rect 942 6422 946 6436
rect 950 6431 954 6436
rect 950 6427 980 6431
rect 942 6415 955 6422
rect 951 6413 955 6415
rect 951 6401 953 6413
rect 922 6372 926 6401
rect 907 6367 915 6372
rect 895 6366 915 6367
rect 922 6366 935 6372
rect 911 6344 915 6366
rect 931 6344 935 6366
rect 951 6344 955 6401
rect 974 6379 980 6427
rect 1045 6399 1049 6456
rect 1045 6387 1054 6399
rect 971 6367 974 6379
rect 971 6344 975 6367
rect 1045 6304 1049 6387
rect 1091 6368 1095 6436
rect 1113 6407 1117 6456
rect 1123 6435 1127 6456
rect 1143 6444 1147 6456
rect 1151 6452 1155 6456
rect 1151 6448 1185 6452
rect 1143 6440 1173 6444
rect 1143 6439 1161 6440
rect 1123 6431 1147 6435
rect 1091 6356 1093 6368
rect 1091 6344 1095 6356
rect 1113 6349 1117 6395
rect 1109 6343 1117 6349
rect 1109 6314 1113 6343
rect 1141 6336 1147 6431
rect 1109 6307 1117 6314
rect 1113 6284 1117 6307
rect 1121 6284 1125 6324
rect 1141 6304 1145 6336
rect 1181 6322 1185 6448
rect 1197 6342 1201 6456
rect 1219 6444 1223 6456
rect 1221 6432 1223 6444
rect 1229 6444 1233 6456
rect 1229 6432 1231 6444
rect 1149 6310 1173 6312
rect 1149 6308 1185 6310
rect 1149 6304 1153 6308
rect 1195 6304 1199 6330
rect 1213 6322 1217 6432
rect 1251 6424 1255 6456
rect 1222 6420 1255 6424
rect 1222 6356 1226 6420
rect 1242 6371 1246 6400
rect 1261 6398 1265 6456
rect 1281 6399 1285 6436
rect 1331 6429 1335 6436
rect 1320 6425 1335 6429
rect 1242 6363 1251 6371
rect 1222 6344 1225 6356
rect 1215 6304 1219 6310
rect 1227 6304 1231 6344
rect 1247 6304 1251 6363
rect 1261 6304 1265 6386
rect 1281 6344 1285 6387
rect 1320 6379 1326 6425
rect 1351 6413 1355 6436
rect 1371 6413 1375 6436
rect 1346 6401 1355 6413
rect 1321 6352 1326 6367
rect 1349 6352 1355 6401
rect 1321 6348 1335 6352
rect 1331 6344 1335 6348
rect 1341 6348 1355 6352
rect 1341 6344 1345 6348
rect 1371 6344 1375 6401
rect 1391 6379 1395 6436
rect 1391 6367 1393 6379
rect 1391 6352 1395 6367
rect 1465 6359 1469 6436
rect 1485 6413 1489 6436
rect 1505 6431 1509 6436
rect 1505 6424 1518 6431
rect 1575 6430 1579 6436
rect 1485 6401 1494 6413
rect 1381 6348 1395 6352
rect 1381 6344 1385 6348
rect 1467 6347 1474 6359
rect 1470 6304 1474 6347
rect 1492 6344 1496 6401
rect 1514 6379 1518 6424
rect 1561 6418 1573 6430
rect 1514 6356 1518 6367
rect 1500 6348 1518 6356
rect 1500 6344 1504 6348
rect 1561 6344 1565 6418
rect 1595 6393 1599 6436
rect 1586 6381 1599 6393
rect 1583 6304 1587 6381
rect 1605 6379 1609 6436
rect 1665 6399 1669 6456
rect 1665 6387 1674 6399
rect 1605 6367 1614 6379
rect 1605 6304 1609 6367
rect 1665 6304 1669 6387
rect 1711 6368 1715 6436
rect 1733 6407 1737 6456
rect 1743 6435 1747 6456
rect 1763 6444 1767 6456
rect 1771 6452 1775 6456
rect 1771 6448 1805 6452
rect 1763 6440 1793 6444
rect 1763 6439 1781 6440
rect 1743 6431 1767 6435
rect 1711 6356 1713 6368
rect 1711 6344 1715 6356
rect 1733 6349 1737 6395
rect 1729 6343 1737 6349
rect 1729 6314 1733 6343
rect 1761 6336 1767 6431
rect 1729 6307 1737 6314
rect 1733 6284 1737 6307
rect 1741 6284 1745 6324
rect 1761 6304 1765 6336
rect 1801 6322 1805 6448
rect 1817 6342 1821 6456
rect 1839 6444 1843 6456
rect 1841 6432 1843 6444
rect 1849 6444 1853 6456
rect 1849 6432 1851 6444
rect 1769 6310 1793 6312
rect 1769 6308 1805 6310
rect 1769 6304 1773 6308
rect 1815 6304 1819 6330
rect 1833 6322 1837 6432
rect 1871 6424 1875 6456
rect 1842 6420 1875 6424
rect 1842 6356 1846 6420
rect 1862 6371 1866 6400
rect 1881 6398 1885 6456
rect 1901 6399 1905 6436
rect 1951 6431 1955 6436
rect 1942 6424 1955 6431
rect 1862 6363 1871 6371
rect 1842 6344 1845 6356
rect 1835 6304 1839 6310
rect 1847 6304 1851 6344
rect 1867 6304 1871 6363
rect 1881 6304 1885 6386
rect 1901 6344 1905 6387
rect 1942 6379 1946 6424
rect 1971 6413 1975 6436
rect 1966 6401 1975 6413
rect 1942 6356 1946 6367
rect 1942 6348 1960 6356
rect 1956 6344 1960 6348
rect 1964 6344 1968 6401
rect 1991 6359 1995 6436
rect 2053 6416 2057 6436
rect 2049 6409 2057 6416
rect 2063 6416 2067 6436
rect 2063 6409 2077 6416
rect 2049 6393 2055 6409
rect 2046 6381 2055 6393
rect 1986 6347 1993 6359
rect 1986 6304 1990 6347
rect 2051 6304 2055 6381
rect 2071 6393 2077 6409
rect 2071 6381 2074 6393
rect 2071 6304 2075 6381
rect 2145 6359 2149 6436
rect 2165 6413 2169 6436
rect 2185 6431 2189 6436
rect 2185 6424 2198 6431
rect 2165 6401 2174 6413
rect 2147 6347 2154 6359
rect 2150 6304 2154 6347
rect 2172 6344 2176 6401
rect 2194 6379 2198 6424
rect 2252 6413 2256 6456
rect 2245 6401 2254 6413
rect 2194 6356 2198 6367
rect 2180 6348 2198 6356
rect 2180 6344 2184 6348
rect 2245 6344 2249 6401
rect 2274 6399 2278 6436
rect 2282 6432 2286 6436
rect 2282 6426 2301 6432
rect 2294 6413 2301 6426
rect 2353 6416 2357 6436
rect 2343 6409 2357 6416
rect 2363 6416 2367 6436
rect 2363 6409 2371 6416
rect 2274 6364 2280 6387
rect 2294 6364 2301 6401
rect 2343 6393 2349 6409
rect 2346 6381 2349 6393
rect 2265 6358 2280 6364
rect 2285 6358 2301 6364
rect 2265 6344 2269 6358
rect 2285 6344 2289 6358
rect 2345 6304 2349 6381
rect 2365 6393 2371 6409
rect 2365 6381 2374 6393
rect 2365 6304 2369 6381
rect 2425 6379 2429 6456
rect 2445 6379 2449 6456
rect 2491 6379 2495 6456
rect 2511 6379 2515 6456
rect 2573 6416 2577 6436
rect 2569 6409 2577 6416
rect 2583 6416 2587 6436
rect 2753 6416 2757 6436
rect 2583 6409 2597 6416
rect 2569 6393 2575 6409
rect 2566 6381 2575 6393
rect 2426 6367 2441 6379
rect 2437 6344 2441 6367
rect 2445 6367 2454 6379
rect 2486 6367 2495 6379
rect 2445 6344 2449 6367
rect 2491 6344 2495 6367
rect 2499 6367 2514 6379
rect 2499 6344 2503 6367
rect 2571 6304 2575 6381
rect 2591 6393 2597 6409
rect 2591 6381 2594 6393
rect 2591 6304 2595 6381
rect 2688 6359 2692 6416
rect 2665 6347 2673 6359
rect 2685 6347 2692 6359
rect 2665 6304 2669 6347
rect 2696 6339 2700 6416
rect 2704 6359 2708 6416
rect 2749 6409 2757 6416
rect 2763 6416 2767 6436
rect 2763 6409 2777 6416
rect 2749 6393 2755 6409
rect 2746 6381 2755 6393
rect 2704 6347 2714 6359
rect 2694 6320 2700 6327
rect 2685 6316 2700 6320
rect 2714 6316 2720 6347
rect 2685 6304 2689 6316
rect 2705 6312 2720 6316
rect 2705 6304 2709 6312
rect 2751 6304 2755 6381
rect 2771 6393 2777 6409
rect 2771 6381 2774 6393
rect 2771 6304 2775 6381
rect 2868 6359 2872 6416
rect 2845 6347 2853 6359
rect 2865 6347 2872 6359
rect 2845 6304 2849 6347
rect 2876 6339 2880 6416
rect 2884 6359 2888 6416
rect 2945 6359 2949 6436
rect 2965 6413 2969 6436
rect 2985 6431 2989 6436
rect 2985 6424 2998 6431
rect 2965 6401 2974 6413
rect 2884 6347 2894 6359
rect 2947 6347 2954 6359
rect 2874 6320 2880 6327
rect 2865 6316 2880 6320
rect 2894 6316 2900 6347
rect 2865 6304 2869 6316
rect 2885 6312 2900 6316
rect 2885 6304 2889 6312
rect 2950 6304 2954 6347
rect 2972 6344 2976 6401
rect 2994 6379 2998 6424
rect 2994 6356 2998 6367
rect 3045 6359 3049 6436
rect 3065 6413 3069 6436
rect 3085 6431 3089 6436
rect 3085 6424 3098 6431
rect 3065 6401 3074 6413
rect 2980 6348 2998 6356
rect 2980 6344 2984 6348
rect 3047 6347 3054 6359
rect 3050 6304 3054 6347
rect 3072 6344 3076 6401
rect 3094 6379 3098 6424
rect 3145 6399 3149 6456
rect 3205 6399 3209 6456
rect 3254 6432 3258 6436
rect 3239 6426 3258 6432
rect 3239 6413 3246 6426
rect 3145 6387 3154 6399
rect 3205 6387 3214 6399
rect 3094 6356 3098 6367
rect 3080 6348 3098 6356
rect 3080 6344 3084 6348
rect 3145 6304 3149 6387
rect 3205 6304 3209 6387
rect 3239 6364 3246 6401
rect 3262 6399 3266 6436
rect 3284 6413 3288 6456
rect 3351 6431 3355 6436
rect 3342 6424 3355 6431
rect 3286 6401 3295 6413
rect 3260 6364 3266 6387
rect 3239 6358 3255 6364
rect 3260 6358 3275 6364
rect 3251 6344 3255 6358
rect 3271 6344 3275 6358
rect 3291 6344 3295 6401
rect 3342 6379 3346 6424
rect 3371 6413 3375 6436
rect 3366 6401 3375 6413
rect 3342 6356 3346 6367
rect 3342 6348 3360 6356
rect 3356 6344 3360 6348
rect 3364 6344 3368 6401
rect 3391 6359 3395 6436
rect 3472 6413 3476 6456
rect 3465 6401 3474 6413
rect 3386 6347 3393 6359
rect 3386 6304 3390 6347
rect 3465 6344 3469 6401
rect 3494 6399 3498 6436
rect 3502 6432 3506 6436
rect 3502 6426 3521 6432
rect 3514 6413 3521 6426
rect 3572 6413 3576 6456
rect 3565 6401 3574 6413
rect 3494 6364 3500 6387
rect 3514 6364 3521 6401
rect 3485 6358 3500 6364
rect 3505 6358 3521 6364
rect 3485 6344 3489 6358
rect 3505 6344 3509 6358
rect 3565 6344 3569 6401
rect 3594 6399 3598 6436
rect 3602 6432 3606 6436
rect 3602 6426 3621 6432
rect 3614 6413 3621 6426
rect 3594 6364 3600 6387
rect 3614 6364 3621 6401
rect 3585 6358 3600 6364
rect 3605 6358 3621 6364
rect 3652 6359 3656 6416
rect 3585 6344 3589 6358
rect 3605 6344 3609 6358
rect 3646 6347 3656 6359
rect 3640 6316 3646 6347
rect 3660 6339 3664 6416
rect 3668 6359 3672 6416
rect 3765 6359 3769 6436
rect 3785 6413 3789 6436
rect 3805 6431 3809 6436
rect 3851 6431 3855 6436
rect 3805 6424 3818 6431
rect 3785 6401 3794 6413
rect 3668 6347 3675 6359
rect 3687 6347 3695 6359
rect 3767 6347 3774 6359
rect 3660 6320 3666 6327
rect 3660 6316 3675 6320
rect 3640 6312 3655 6316
rect 3651 6304 3655 6312
rect 3671 6304 3675 6316
rect 3691 6304 3695 6347
rect 3770 6304 3774 6347
rect 3792 6344 3796 6401
rect 3814 6379 3818 6424
rect 3842 6424 3855 6431
rect 3842 6379 3846 6424
rect 3871 6413 3875 6436
rect 3866 6401 3875 6413
rect 3814 6356 3818 6367
rect 3800 6348 3818 6356
rect 3842 6356 3846 6367
rect 3842 6348 3860 6356
rect 3800 6344 3804 6348
rect 3856 6344 3860 6348
rect 3864 6344 3868 6401
rect 3891 6359 3895 6436
rect 3951 6399 3955 6456
rect 4013 6416 4017 6436
rect 3946 6387 3955 6399
rect 4009 6409 4017 6416
rect 4023 6416 4027 6436
rect 4115 6430 4119 6436
rect 4101 6418 4113 6430
rect 4023 6409 4037 6416
rect 4009 6393 4015 6409
rect 3886 6347 3893 6359
rect 3886 6304 3890 6347
rect 3951 6304 3955 6387
rect 4006 6381 4015 6393
rect 4011 6304 4015 6381
rect 4031 6393 4037 6409
rect 4031 6381 4034 6393
rect 4031 6304 4035 6381
rect 4101 6344 4105 6418
rect 4135 6393 4139 6436
rect 4126 6381 4139 6393
rect 4123 6304 4127 6381
rect 4145 6379 4149 6436
rect 4193 6416 4197 6436
rect 4189 6409 4197 6416
rect 4203 6416 4207 6436
rect 4203 6409 4217 6416
rect 4189 6393 4195 6409
rect 4186 6381 4195 6393
rect 4145 6367 4154 6379
rect 4145 6304 4149 6367
rect 4191 6304 4195 6381
rect 4211 6393 4217 6409
rect 4211 6381 4214 6393
rect 4211 6304 4215 6381
rect 4308 6359 4312 6416
rect 4285 6347 4293 6359
rect 4305 6347 4312 6359
rect 4285 6304 4289 6347
rect 4316 6339 4320 6416
rect 4324 6359 4328 6416
rect 4408 6359 4412 6416
rect 4324 6347 4334 6359
rect 4385 6347 4393 6359
rect 4405 6347 4412 6359
rect 4314 6320 4320 6327
rect 4305 6316 4320 6320
rect 4334 6316 4340 6347
rect 4305 6304 4309 6316
rect 4325 6312 4340 6316
rect 4325 6304 4329 6312
rect 4385 6304 4389 6347
rect 4416 6339 4420 6416
rect 4424 6359 4428 6416
rect 4508 6359 4512 6416
rect 4424 6347 4434 6359
rect 4485 6347 4493 6359
rect 4505 6347 4512 6359
rect 4414 6320 4420 6327
rect 4405 6316 4420 6320
rect 4434 6316 4440 6347
rect 4405 6304 4409 6316
rect 4425 6312 4440 6316
rect 4425 6304 4429 6312
rect 4485 6304 4489 6347
rect 4516 6339 4520 6416
rect 4524 6359 4528 6416
rect 4571 6399 4575 6456
rect 4634 6432 4638 6436
rect 4619 6426 4638 6432
rect 4619 6413 4626 6426
rect 4566 6387 4575 6399
rect 4524 6347 4534 6359
rect 4514 6320 4520 6327
rect 4505 6316 4520 6320
rect 4534 6316 4540 6347
rect 4505 6304 4509 6316
rect 4525 6312 4540 6316
rect 4525 6304 4529 6312
rect 4571 6304 4575 6387
rect 4619 6364 4626 6401
rect 4642 6399 4646 6436
rect 4664 6413 4668 6456
rect 4734 6432 4738 6436
rect 4719 6426 4738 6432
rect 4719 6413 4726 6426
rect 4666 6401 4675 6413
rect 4640 6364 4646 6387
rect 4619 6358 4635 6364
rect 4640 6358 4655 6364
rect 4631 6344 4635 6358
rect 4651 6344 4655 6358
rect 4671 6344 4675 6401
rect 4719 6364 4726 6401
rect 4742 6399 4746 6436
rect 4764 6413 4768 6456
rect 4831 6431 4835 6436
rect 4822 6424 4835 6431
rect 4766 6401 4775 6413
rect 4740 6364 4746 6387
rect 4719 6358 4735 6364
rect 4740 6358 4755 6364
rect 4731 6344 4735 6358
rect 4751 6344 4755 6358
rect 4771 6344 4775 6401
rect 4822 6379 4826 6424
rect 4851 6413 4855 6436
rect 4846 6401 4855 6413
rect 4822 6356 4826 6367
rect 4822 6348 4840 6356
rect 4836 6344 4840 6348
rect 4844 6344 4848 6401
rect 4871 6359 4875 6436
rect 4945 6359 4949 6436
rect 4965 6413 4969 6436
rect 4985 6431 4989 6436
rect 5031 6431 5035 6436
rect 4985 6424 4998 6431
rect 4965 6401 4974 6413
rect 4866 6347 4873 6359
rect 4947 6347 4954 6359
rect 4866 6304 4870 6347
rect 4950 6304 4954 6347
rect 4972 6344 4976 6401
rect 4994 6379 4998 6424
rect 5022 6424 5035 6431
rect 5022 6379 5026 6424
rect 5051 6413 5055 6436
rect 5046 6401 5055 6413
rect 4994 6356 4998 6367
rect 4980 6348 4998 6356
rect 5022 6356 5026 6367
rect 5022 6348 5040 6356
rect 4980 6344 4984 6348
rect 5036 6344 5040 6348
rect 5044 6344 5048 6401
rect 5071 6359 5075 6436
rect 5434 6432 5438 6436
rect 5419 6426 5438 6432
rect 5168 6359 5172 6416
rect 5066 6347 5073 6359
rect 5145 6347 5153 6359
rect 5165 6347 5172 6359
rect 5066 6304 5070 6347
rect 5145 6304 5149 6347
rect 5176 6339 5180 6416
rect 5184 6359 5188 6416
rect 5268 6359 5272 6416
rect 5184 6347 5194 6359
rect 5245 6347 5253 6359
rect 5265 6347 5272 6359
rect 5174 6320 5180 6327
rect 5165 6316 5180 6320
rect 5194 6316 5200 6347
rect 5165 6304 5169 6316
rect 5185 6312 5200 6316
rect 5185 6304 5189 6312
rect 5245 6304 5249 6347
rect 5276 6339 5280 6416
rect 5284 6359 5288 6416
rect 5368 6359 5372 6416
rect 5284 6347 5294 6359
rect 5345 6347 5353 6359
rect 5365 6347 5372 6359
rect 5274 6320 5280 6327
rect 5265 6316 5280 6320
rect 5294 6316 5300 6347
rect 5265 6304 5269 6316
rect 5285 6312 5300 6316
rect 5285 6304 5289 6312
rect 5345 6304 5349 6347
rect 5376 6339 5380 6416
rect 5384 6359 5388 6416
rect 5419 6413 5426 6426
rect 5419 6364 5426 6401
rect 5442 6399 5446 6436
rect 5464 6413 5468 6456
rect 5552 6413 5556 6456
rect 5466 6401 5475 6413
rect 5440 6364 5446 6387
rect 5384 6347 5394 6359
rect 5419 6358 5435 6364
rect 5440 6358 5455 6364
rect 5374 6320 5380 6327
rect 5365 6316 5380 6320
rect 5394 6316 5400 6347
rect 5431 6344 5435 6358
rect 5451 6344 5455 6358
rect 5471 6344 5475 6401
rect 5545 6401 5554 6413
rect 5545 6344 5549 6401
rect 5574 6399 5578 6436
rect 5582 6432 5586 6436
rect 5582 6426 5601 6432
rect 5594 6413 5601 6426
rect 5574 6364 5580 6387
rect 5594 6364 5601 6401
rect 5565 6358 5580 6364
rect 5585 6358 5601 6364
rect 5645 6399 5649 6456
rect 5694 6432 5698 6436
rect 5679 6426 5698 6432
rect 5679 6413 5686 6426
rect 5645 6387 5654 6399
rect 5565 6344 5569 6358
rect 5585 6344 5589 6358
rect 5365 6304 5369 6316
rect 5385 6312 5400 6316
rect 5385 6304 5389 6312
rect 5645 6304 5649 6387
rect 5679 6364 5686 6401
rect 5702 6399 5706 6436
rect 5724 6413 5728 6456
rect 5726 6401 5735 6413
rect 5700 6364 5706 6387
rect 5679 6358 5695 6364
rect 5700 6358 5715 6364
rect 5691 6344 5695 6358
rect 5711 6344 5715 6358
rect 5731 6344 5735 6401
rect 5792 6359 5796 6416
rect 5786 6347 5796 6359
rect 5780 6316 5786 6347
rect 5800 6339 5804 6416
rect 5808 6359 5812 6416
rect 5912 6413 5916 6456
rect 5905 6401 5914 6413
rect 5808 6347 5815 6359
rect 5827 6347 5835 6359
rect 5800 6320 5806 6327
rect 5800 6316 5815 6320
rect 5780 6312 5795 6316
rect 5791 6304 5795 6312
rect 5811 6304 5815 6316
rect 5831 6304 5835 6347
rect 5905 6344 5909 6401
rect 5934 6399 5938 6436
rect 5942 6432 5946 6436
rect 5942 6426 5961 6432
rect 5954 6413 5961 6426
rect 5934 6364 5940 6387
rect 5954 6364 5961 6401
rect 5925 6358 5940 6364
rect 5945 6358 5961 6364
rect 6005 6399 6009 6456
rect 6072 6413 6076 6456
rect 6065 6401 6074 6413
rect 6005 6387 6014 6399
rect 5925 6344 5929 6358
rect 5945 6344 5949 6358
rect 6005 6304 6009 6387
rect 6065 6344 6069 6401
rect 6094 6399 6098 6436
rect 6102 6432 6106 6436
rect 6102 6426 6121 6432
rect 6114 6413 6121 6426
rect 6094 6364 6100 6387
rect 6114 6364 6121 6401
rect 6085 6358 6100 6364
rect 6105 6358 6121 6364
rect 6165 6359 6169 6436
rect 6185 6413 6189 6436
rect 6205 6431 6209 6436
rect 6205 6424 6218 6431
rect 6185 6401 6194 6413
rect 6085 6344 6089 6358
rect 6105 6344 6109 6358
rect 6167 6347 6174 6359
rect 6170 6304 6174 6347
rect 6192 6344 6196 6401
rect 6214 6379 6218 6424
rect 6272 6413 6276 6456
rect 6265 6401 6274 6413
rect 6214 6356 6218 6367
rect 6200 6348 6218 6356
rect 6200 6344 6204 6348
rect 6265 6344 6269 6401
rect 6294 6399 6298 6436
rect 6302 6432 6306 6436
rect 6302 6426 6321 6432
rect 6314 6413 6321 6426
rect 6294 6364 6300 6387
rect 6314 6364 6321 6401
rect 6285 6358 6300 6364
rect 6305 6358 6321 6364
rect 6352 6359 6356 6416
rect 6285 6344 6289 6358
rect 6305 6344 6309 6358
rect 6346 6347 6356 6359
rect 6340 6316 6346 6347
rect 6360 6339 6364 6416
rect 6368 6359 6372 6416
rect 6488 6359 6492 6416
rect 6368 6347 6375 6359
rect 6387 6347 6395 6359
rect 6360 6320 6366 6327
rect 6360 6316 6375 6320
rect 6340 6312 6355 6316
rect 6351 6304 6355 6312
rect 6371 6304 6375 6316
rect 6391 6304 6395 6347
rect 6465 6347 6473 6359
rect 6485 6347 6492 6359
rect 6465 6304 6469 6347
rect 6496 6339 6500 6416
rect 6504 6359 6508 6416
rect 6551 6399 6555 6456
rect 6614 6428 6618 6436
rect 6546 6387 6555 6399
rect 6504 6347 6514 6359
rect 6494 6320 6500 6327
rect 6485 6316 6500 6320
rect 6514 6316 6520 6347
rect 6485 6304 6489 6316
rect 6505 6312 6520 6316
rect 6505 6304 6509 6312
rect 6551 6304 6555 6387
rect 6601 6421 6618 6428
rect 6601 6379 6607 6421
rect 6622 6413 6626 6436
rect 6642 6422 6646 6436
rect 6650 6431 6654 6436
rect 6650 6427 6680 6431
rect 6642 6415 6655 6422
rect 6651 6413 6655 6415
rect 6651 6401 6653 6413
rect 6622 6372 6626 6401
rect 6607 6367 6615 6372
rect 6595 6366 6615 6367
rect 6622 6366 6635 6372
rect 6611 6344 6615 6366
rect 6631 6344 6635 6366
rect 6651 6344 6655 6401
rect 6674 6379 6680 6427
rect 6671 6367 6674 6379
rect 6671 6344 6675 6367
rect 35 6260 39 6264
rect 55 6260 59 6264
rect 69 6260 73 6264
rect 89 6260 93 6264
rect 101 6260 105 6264
rect 121 6260 125 6264
rect 167 6260 171 6264
rect 175 6260 179 6264
rect 195 6260 199 6264
rect 203 6260 207 6264
rect 225 6260 229 6264
rect 290 6260 294 6264
rect 312 6260 316 6264
rect 320 6260 324 6264
rect 371 6260 375 6264
rect 391 6260 395 6264
rect 465 6260 469 6264
rect 485 6260 489 6264
rect 531 6260 535 6264
rect 551 6260 555 6264
rect 611 6260 615 6264
rect 633 6260 637 6264
rect 641 6260 645 6264
rect 661 6260 665 6264
rect 669 6260 673 6264
rect 715 6260 719 6264
rect 735 6260 739 6264
rect 747 6260 751 6264
rect 767 6260 771 6264
rect 781 6260 785 6264
rect 801 6260 805 6264
rect 851 6260 855 6264
rect 911 6260 915 6264
rect 931 6260 935 6264
rect 951 6260 955 6264
rect 971 6260 975 6264
rect 1045 6260 1049 6264
rect 1091 6260 1095 6264
rect 1113 6260 1117 6264
rect 1121 6260 1125 6264
rect 1141 6260 1145 6264
rect 1149 6260 1153 6264
rect 1195 6260 1199 6264
rect 1215 6260 1219 6264
rect 1227 6260 1231 6264
rect 1247 6260 1251 6264
rect 1261 6260 1265 6264
rect 1281 6260 1285 6264
rect 1331 6260 1335 6264
rect 1341 6260 1345 6264
rect 1371 6260 1375 6264
rect 1381 6260 1385 6264
rect 1470 6260 1474 6264
rect 1492 6260 1496 6264
rect 1500 6260 1504 6264
rect 1561 6260 1565 6264
rect 1583 6260 1587 6264
rect 1605 6260 1609 6264
rect 1665 6260 1669 6264
rect 1711 6260 1715 6264
rect 1733 6260 1737 6264
rect 1741 6260 1745 6264
rect 1761 6260 1765 6264
rect 1769 6260 1773 6264
rect 1815 6260 1819 6264
rect 1835 6260 1839 6264
rect 1847 6260 1851 6264
rect 1867 6260 1871 6264
rect 1881 6260 1885 6264
rect 1901 6260 1905 6264
rect 1956 6260 1960 6264
rect 1964 6260 1968 6264
rect 1986 6260 1990 6264
rect 2051 6260 2055 6264
rect 2071 6260 2075 6264
rect 2150 6260 2154 6264
rect 2172 6260 2176 6264
rect 2180 6260 2184 6264
rect 2245 6260 2249 6264
rect 2265 6260 2269 6264
rect 2285 6260 2289 6264
rect 2345 6260 2349 6264
rect 2365 6260 2369 6264
rect 2437 6260 2441 6264
rect 2445 6260 2449 6264
rect 2491 6260 2495 6264
rect 2499 6260 2503 6264
rect 2571 6260 2575 6264
rect 2591 6260 2595 6264
rect 2665 6260 2669 6264
rect 2685 6260 2689 6264
rect 2705 6260 2709 6264
rect 2751 6260 2755 6264
rect 2771 6260 2775 6264
rect 2845 6260 2849 6264
rect 2865 6260 2869 6264
rect 2885 6260 2889 6264
rect 2950 6260 2954 6264
rect 2972 6260 2976 6264
rect 2980 6260 2984 6264
rect 3050 6260 3054 6264
rect 3072 6260 3076 6264
rect 3080 6260 3084 6264
rect 3145 6260 3149 6264
rect 3205 6260 3209 6264
rect 3251 6260 3255 6264
rect 3271 6260 3275 6264
rect 3291 6260 3295 6264
rect 3356 6260 3360 6264
rect 3364 6260 3368 6264
rect 3386 6260 3390 6264
rect 3465 6260 3469 6264
rect 3485 6260 3489 6264
rect 3505 6260 3509 6264
rect 3565 6260 3569 6264
rect 3585 6260 3589 6264
rect 3605 6260 3609 6264
rect 3651 6260 3655 6264
rect 3671 6260 3675 6264
rect 3691 6260 3695 6264
rect 3770 6260 3774 6264
rect 3792 6260 3796 6264
rect 3800 6260 3804 6264
rect 3856 6260 3860 6264
rect 3864 6260 3868 6264
rect 3886 6260 3890 6264
rect 3951 6260 3955 6264
rect 4011 6260 4015 6264
rect 4031 6260 4035 6264
rect 4101 6260 4105 6264
rect 4123 6260 4127 6264
rect 4145 6260 4149 6264
rect 4191 6260 4195 6264
rect 4211 6260 4215 6264
rect 4285 6260 4289 6264
rect 4305 6260 4309 6264
rect 4325 6260 4329 6264
rect 4385 6260 4389 6264
rect 4405 6260 4409 6264
rect 4425 6260 4429 6264
rect 4485 6260 4489 6264
rect 4505 6260 4509 6264
rect 4525 6260 4529 6264
rect 4571 6260 4575 6264
rect 4631 6260 4635 6264
rect 4651 6260 4655 6264
rect 4671 6260 4675 6264
rect 4731 6260 4735 6264
rect 4751 6260 4755 6264
rect 4771 6260 4775 6264
rect 4836 6260 4840 6264
rect 4844 6260 4848 6264
rect 4866 6260 4870 6264
rect 4950 6260 4954 6264
rect 4972 6260 4976 6264
rect 4980 6260 4984 6264
rect 5036 6260 5040 6264
rect 5044 6260 5048 6264
rect 5066 6260 5070 6264
rect 5145 6260 5149 6264
rect 5165 6260 5169 6264
rect 5185 6260 5189 6264
rect 5245 6260 5249 6264
rect 5265 6260 5269 6264
rect 5285 6260 5289 6264
rect 5345 6260 5349 6264
rect 5365 6260 5369 6264
rect 5385 6260 5389 6264
rect 5431 6260 5435 6264
rect 5451 6260 5455 6264
rect 5471 6260 5475 6264
rect 5545 6260 5549 6264
rect 5565 6260 5569 6264
rect 5585 6260 5589 6264
rect 5645 6260 5649 6264
rect 5691 6260 5695 6264
rect 5711 6260 5715 6264
rect 5731 6260 5735 6264
rect 5791 6260 5795 6264
rect 5811 6260 5815 6264
rect 5831 6260 5835 6264
rect 5905 6260 5909 6264
rect 5925 6260 5929 6264
rect 5945 6260 5949 6264
rect 6005 6260 6009 6264
rect 6065 6260 6069 6264
rect 6085 6260 6089 6264
rect 6105 6260 6109 6264
rect 6170 6260 6174 6264
rect 6192 6260 6196 6264
rect 6200 6260 6204 6264
rect 6265 6260 6269 6264
rect 6285 6260 6289 6264
rect 6305 6260 6309 6264
rect 6351 6260 6355 6264
rect 6371 6260 6375 6264
rect 6391 6260 6395 6264
rect 6465 6260 6469 6264
rect 6485 6260 6489 6264
rect 6505 6260 6509 6264
rect 6551 6260 6555 6264
rect 6611 6260 6615 6264
rect 6631 6260 6635 6264
rect 6651 6260 6655 6264
rect 6671 6260 6675 6264
rect 31 6236 35 6240
rect 53 6236 57 6240
rect 61 6236 65 6240
rect 81 6236 85 6240
rect 89 6236 93 6240
rect 135 6236 139 6240
rect 155 6236 159 6240
rect 167 6236 171 6240
rect 187 6236 191 6240
rect 201 6236 205 6240
rect 221 6236 225 6240
rect 285 6236 289 6240
rect 305 6236 309 6240
rect 325 6236 329 6240
rect 385 6236 389 6240
rect 405 6236 409 6240
rect 451 6236 455 6240
rect 459 6236 463 6240
rect 545 6236 549 6240
rect 565 6236 569 6240
rect 616 6236 620 6240
rect 624 6236 628 6240
rect 646 6236 650 6240
rect 730 6236 734 6240
rect 752 6236 756 6240
rect 760 6236 764 6240
rect 811 6236 815 6240
rect 819 6236 823 6240
rect 905 6236 909 6240
rect 925 6236 929 6240
rect 945 6236 949 6240
rect 991 6236 995 6240
rect 1001 6236 1005 6240
rect 1021 6236 1025 6240
rect 1105 6236 1109 6240
rect 1151 6236 1155 6240
rect 1159 6236 1163 6240
rect 1250 6236 1254 6240
rect 1272 6236 1276 6240
rect 1280 6236 1284 6240
rect 1345 6236 1349 6240
rect 1405 6236 1409 6240
rect 1451 6236 1455 6240
rect 1459 6236 1463 6240
rect 1531 6236 1535 6240
rect 1539 6236 1543 6240
rect 1611 6236 1615 6240
rect 1671 6236 1675 6240
rect 1679 6236 1683 6240
rect 1751 6236 1755 6240
rect 1759 6236 1763 6240
rect 1836 6236 1840 6240
rect 1844 6236 1848 6240
rect 1866 6236 1870 6240
rect 1931 6236 1935 6240
rect 2005 6236 2009 6240
rect 2025 6236 2029 6240
rect 2045 6236 2049 6240
rect 2091 6236 2095 6240
rect 2170 6236 2174 6240
rect 2192 6236 2196 6240
rect 2200 6236 2204 6240
rect 2251 6236 2255 6240
rect 2330 6236 2334 6240
rect 2352 6236 2356 6240
rect 2360 6236 2364 6240
rect 2425 6236 2429 6240
rect 2445 6236 2449 6240
rect 2465 6236 2469 6240
rect 2525 6236 2529 6240
rect 2545 6236 2549 6240
rect 2565 6236 2569 6240
rect 2637 6236 2641 6240
rect 2645 6236 2649 6240
rect 2705 6236 2709 6240
rect 2725 6236 2729 6240
rect 2745 6236 2749 6240
rect 2805 6236 2809 6240
rect 2825 6236 2829 6240
rect 2845 6236 2849 6240
rect 2865 6236 2869 6240
rect 2925 6236 2929 6240
rect 2971 6236 2975 6240
rect 2991 6236 2995 6240
rect 3011 6236 3015 6240
rect 3085 6236 3089 6240
rect 3105 6236 3109 6240
rect 3125 6236 3129 6240
rect 3185 6236 3189 6240
rect 3205 6236 3209 6240
rect 3225 6236 3229 6240
rect 3285 6236 3289 6240
rect 3305 6236 3309 6240
rect 3325 6236 3329 6240
rect 3385 6236 3389 6240
rect 3445 6236 3449 6240
rect 3465 6236 3469 6240
rect 3485 6236 3489 6240
rect 3531 6236 3535 6240
rect 3551 6236 3555 6240
rect 3571 6236 3575 6240
rect 3631 6236 3635 6240
rect 3691 6236 3695 6240
rect 3711 6236 3715 6240
rect 3731 6236 3735 6240
rect 3805 6236 3809 6240
rect 3825 6236 3829 6240
rect 3871 6236 3875 6240
rect 3891 6236 3895 6240
rect 3970 6236 3974 6240
rect 3992 6236 3996 6240
rect 4000 6236 4004 6240
rect 4056 6236 4060 6240
rect 4064 6236 4068 6240
rect 4086 6236 4090 6240
rect 4177 6236 4181 6240
rect 4185 6236 4189 6240
rect 4231 6236 4235 6240
rect 4305 6236 4309 6240
rect 4325 6236 4329 6240
rect 4371 6236 4375 6240
rect 4393 6236 4397 6240
rect 4415 6236 4419 6240
rect 4490 6236 4494 6240
rect 4512 6236 4516 6240
rect 4520 6236 4524 6240
rect 4585 6236 4589 6240
rect 4605 6236 4609 6240
rect 4625 6236 4629 6240
rect 4671 6236 4675 6240
rect 4691 6236 4695 6240
rect 4711 6236 4715 6240
rect 4785 6236 4789 6240
rect 4805 6236 4809 6240
rect 4825 6236 4829 6240
rect 4885 6236 4889 6240
rect 4905 6236 4909 6240
rect 4925 6236 4929 6240
rect 4971 6236 4975 6240
rect 4991 6236 4995 6240
rect 5011 6236 5015 6240
rect 5090 6236 5094 6240
rect 5112 6236 5116 6240
rect 5120 6236 5124 6240
rect 5185 6236 5189 6240
rect 5205 6236 5209 6240
rect 5251 6236 5255 6240
rect 5273 6236 5277 6240
rect 5295 6236 5299 6240
rect 5356 6236 5360 6240
rect 5364 6236 5368 6240
rect 5386 6236 5390 6240
rect 5465 6236 5469 6240
rect 5485 6236 5489 6240
rect 5505 6236 5509 6240
rect 5565 6236 5569 6240
rect 5585 6236 5589 6240
rect 5605 6236 5609 6240
rect 5651 6236 5655 6240
rect 5671 6236 5675 6240
rect 5691 6236 5695 6240
rect 5765 6236 5769 6240
rect 5785 6236 5789 6240
rect 5805 6236 5809 6240
rect 5851 6236 5855 6240
rect 5871 6236 5875 6240
rect 5891 6236 5895 6240
rect 5956 6236 5960 6240
rect 5964 6236 5968 6240
rect 5986 6236 5990 6240
rect 6056 6236 6060 6240
rect 6064 6236 6068 6240
rect 6086 6236 6090 6240
rect 6151 6236 6155 6240
rect 6171 6236 6175 6240
rect 6191 6236 6195 6240
rect 6251 6236 6255 6240
rect 6271 6236 6275 6240
rect 6291 6236 6295 6240
rect 6365 6236 6369 6240
rect 6385 6236 6389 6240
rect 6405 6236 6409 6240
rect 6465 6236 6469 6240
rect 6485 6236 6489 6240
rect 6505 6236 6509 6240
rect 6551 6236 6555 6240
rect 6611 6236 6615 6240
rect 53 6193 57 6216
rect 49 6186 57 6193
rect 49 6157 53 6186
rect 61 6176 65 6216
rect 81 6164 85 6196
rect 89 6192 93 6196
rect 89 6190 125 6192
rect 89 6188 113 6190
rect 31 6144 35 6156
rect 49 6151 57 6157
rect 31 6132 33 6144
rect 31 6064 35 6132
rect 53 6105 57 6151
rect 53 6044 57 6093
rect 81 6069 87 6164
rect 63 6065 87 6069
rect 63 6044 67 6065
rect 83 6060 101 6061
rect 83 6056 113 6060
rect 83 6044 87 6056
rect 121 6052 125 6178
rect 135 6170 139 6196
rect 155 6190 159 6196
rect 91 6048 125 6052
rect 91 6044 95 6048
rect 137 6044 141 6158
rect 153 6068 157 6178
rect 167 6156 171 6196
rect 162 6144 165 6156
rect 162 6080 166 6144
rect 187 6137 191 6196
rect 182 6129 191 6137
rect 182 6100 186 6129
rect 201 6114 205 6196
rect 221 6113 225 6156
rect 162 6076 195 6080
rect 161 6056 163 6068
rect 159 6044 163 6056
rect 169 6056 171 6068
rect 169 6044 173 6056
rect 191 6044 195 6076
rect 201 6044 205 6102
rect 221 6064 225 6101
rect 285 6099 289 6156
rect 305 6142 309 6156
rect 325 6142 329 6156
rect 305 6136 320 6142
rect 325 6136 341 6142
rect 314 6113 320 6136
rect 285 6087 294 6099
rect 292 6044 296 6087
rect 314 6064 318 6101
rect 334 6099 341 6136
rect 385 6119 389 6196
rect 386 6107 389 6119
rect 383 6091 389 6107
rect 405 6119 409 6196
rect 451 6133 455 6156
rect 446 6121 455 6133
rect 459 6133 463 6156
rect 459 6121 474 6133
rect 405 6107 414 6119
rect 405 6091 411 6107
rect 334 6074 341 6087
rect 383 6084 397 6091
rect 322 6068 341 6074
rect 322 6064 326 6068
rect 393 6064 397 6084
rect 403 6084 411 6091
rect 403 6064 407 6084
rect 451 6044 455 6121
rect 471 6044 475 6121
rect 545 6119 549 6196
rect 546 6107 549 6119
rect 543 6091 549 6107
rect 565 6119 569 6196
rect 616 6152 620 6156
rect 602 6144 620 6152
rect 602 6133 606 6144
rect 565 6107 574 6119
rect 565 6091 571 6107
rect 543 6084 557 6091
rect 553 6064 557 6084
rect 563 6084 571 6091
rect 563 6064 567 6084
rect 602 6076 606 6121
rect 624 6099 628 6156
rect 646 6153 650 6196
rect 730 6153 734 6196
rect 646 6141 653 6153
rect 727 6141 734 6153
rect 626 6087 635 6099
rect 602 6069 615 6076
rect 611 6064 615 6069
rect 631 6064 635 6087
rect 651 6064 655 6141
rect 725 6064 729 6141
rect 752 6099 756 6156
rect 760 6152 764 6156
rect 760 6144 778 6152
rect 774 6133 778 6144
rect 811 6133 815 6156
rect 806 6121 815 6133
rect 819 6133 823 6156
rect 819 6121 834 6133
rect 745 6087 754 6099
rect 745 6064 749 6087
rect 774 6076 778 6121
rect 765 6069 778 6076
rect 765 6064 769 6069
rect 811 6044 815 6121
rect 831 6044 835 6121
rect 905 6099 909 6156
rect 925 6142 929 6156
rect 945 6142 949 6156
rect 991 6152 995 6156
rect 982 6147 995 6152
rect 925 6136 940 6142
rect 945 6136 961 6142
rect 934 6113 940 6136
rect 905 6087 914 6099
rect 912 6044 916 6087
rect 934 6064 938 6101
rect 954 6099 961 6136
rect 982 6113 986 6147
rect 1001 6133 1005 6156
rect 1021 6151 1025 6156
rect 954 6074 961 6087
rect 942 6068 961 6074
rect 942 6064 946 6068
rect 982 6056 986 6101
rect 1001 6057 1005 6121
rect 1105 6113 1109 6196
rect 1151 6133 1155 6156
rect 1146 6121 1155 6133
rect 1159 6133 1163 6156
rect 1250 6153 1254 6196
rect 1247 6141 1254 6153
rect 1159 6121 1174 6133
rect 1105 6101 1114 6113
rect 1025 6072 1035 6084
rect 1031 6064 1035 6072
rect 982 6051 995 6056
rect 1001 6051 1015 6057
rect 991 6044 995 6051
rect 1011 6044 1015 6051
rect 1105 6044 1109 6101
rect 1151 6044 1155 6121
rect 1171 6044 1175 6121
rect 1245 6064 1249 6141
rect 1272 6099 1276 6156
rect 1280 6152 1284 6156
rect 1280 6144 1298 6152
rect 1294 6133 1298 6144
rect 1265 6087 1274 6099
rect 1265 6064 1269 6087
rect 1294 6076 1298 6121
rect 1285 6069 1298 6076
rect 1345 6113 1349 6196
rect 1405 6113 1409 6196
rect 1451 6133 1455 6156
rect 1446 6121 1455 6133
rect 1459 6133 1463 6156
rect 1531 6133 1535 6156
rect 1459 6121 1474 6133
rect 1526 6121 1535 6133
rect 1539 6133 1543 6156
rect 1539 6121 1554 6133
rect 1345 6101 1354 6113
rect 1405 6101 1414 6113
rect 1285 6064 1289 6069
rect 1345 6044 1349 6101
rect 1405 6044 1409 6101
rect 1451 6044 1455 6121
rect 1471 6044 1475 6121
rect 1531 6044 1535 6121
rect 1551 6044 1555 6121
rect 1611 6113 1615 6196
rect 1671 6133 1675 6156
rect 1666 6121 1675 6133
rect 1679 6133 1683 6156
rect 1751 6133 1755 6156
rect 1679 6121 1694 6133
rect 1746 6121 1755 6133
rect 1759 6133 1763 6156
rect 1836 6152 1840 6156
rect 1822 6144 1840 6152
rect 1822 6133 1826 6144
rect 1759 6121 1774 6133
rect 1606 6101 1615 6113
rect 1611 6044 1615 6101
rect 1671 6044 1675 6121
rect 1691 6044 1695 6121
rect 1751 6044 1755 6121
rect 1771 6044 1775 6121
rect 1822 6076 1826 6121
rect 1844 6099 1848 6156
rect 1866 6153 1870 6196
rect 1866 6141 1873 6153
rect 1846 6087 1855 6099
rect 1822 6069 1835 6076
rect 1831 6064 1835 6069
rect 1851 6064 1855 6087
rect 1871 6064 1875 6141
rect 1931 6113 1935 6196
rect 1926 6101 1935 6113
rect 1931 6044 1935 6101
rect 2005 6099 2009 6156
rect 2025 6142 2029 6156
rect 2045 6142 2049 6156
rect 2025 6136 2040 6142
rect 2045 6136 2061 6142
rect 2034 6113 2040 6136
rect 2005 6087 2014 6099
rect 2012 6044 2016 6087
rect 2034 6064 2038 6101
rect 2054 6099 2061 6136
rect 2091 6113 2095 6196
rect 2170 6153 2174 6196
rect 2167 6141 2174 6153
rect 2086 6101 2095 6113
rect 2054 6074 2061 6087
rect 2042 6068 2061 6074
rect 2042 6064 2046 6068
rect 2091 6044 2095 6101
rect 2165 6064 2169 6141
rect 2192 6099 2196 6156
rect 2200 6152 2204 6156
rect 2200 6144 2218 6152
rect 2214 6133 2218 6144
rect 2185 6087 2194 6099
rect 2185 6064 2189 6087
rect 2214 6076 2218 6121
rect 2251 6113 2255 6196
rect 2330 6153 2334 6196
rect 2327 6141 2334 6153
rect 2246 6101 2255 6113
rect 2205 6069 2218 6076
rect 2205 6064 2209 6069
rect 2251 6044 2255 6101
rect 2325 6064 2329 6141
rect 2352 6099 2356 6156
rect 2360 6152 2364 6156
rect 2425 6153 2429 6196
rect 2445 6184 2449 6196
rect 2465 6188 2469 6196
rect 2465 6184 2480 6188
rect 2445 6180 2460 6184
rect 2454 6173 2460 6180
rect 2360 6144 2378 6152
rect 2374 6133 2378 6144
rect 2425 6141 2433 6153
rect 2445 6141 2452 6153
rect 2345 6087 2354 6099
rect 2345 6064 2349 6087
rect 2374 6076 2378 6121
rect 2448 6084 2452 6141
rect 2456 6084 2460 6161
rect 2474 6153 2480 6184
rect 2464 6141 2474 6153
rect 2464 6084 2468 6141
rect 2525 6099 2529 6156
rect 2545 6142 2549 6156
rect 2565 6142 2569 6156
rect 2545 6136 2560 6142
rect 2565 6136 2581 6142
rect 2554 6113 2560 6136
rect 2525 6087 2534 6099
rect 2365 6069 2378 6076
rect 2365 6064 2369 6069
rect 2532 6044 2536 6087
rect 2554 6064 2558 6101
rect 2574 6099 2581 6136
rect 2637 6133 2641 6156
rect 2626 6121 2641 6133
rect 2645 6133 2649 6156
rect 2705 6153 2709 6196
rect 2725 6184 2729 6196
rect 2745 6188 2749 6196
rect 2745 6184 2760 6188
rect 2725 6180 2740 6184
rect 2734 6173 2740 6180
rect 2705 6141 2713 6153
rect 2725 6141 2732 6153
rect 2645 6121 2654 6133
rect 2574 6074 2581 6087
rect 2562 6068 2581 6074
rect 2562 6064 2566 6068
rect 2625 6044 2629 6121
rect 2645 6044 2649 6121
rect 2728 6084 2732 6141
rect 2736 6084 2740 6161
rect 2754 6153 2760 6184
rect 2744 6141 2754 6153
rect 2744 6084 2748 6141
rect 2805 6133 2809 6156
rect 2806 6121 2809 6133
rect 2800 6073 2806 6121
rect 2825 6099 2829 6156
rect 2845 6134 2849 6156
rect 2865 6134 2869 6156
rect 2845 6128 2858 6134
rect 2865 6133 2885 6134
rect 2865 6128 2873 6133
rect 2854 6099 2858 6128
rect 2827 6087 2829 6099
rect 2825 6085 2829 6087
rect 2825 6078 2838 6085
rect 2800 6069 2830 6073
rect 2826 6064 2830 6069
rect 2834 6064 2838 6078
rect 2854 6064 2858 6087
rect 2873 6079 2879 6121
rect 2862 6072 2879 6079
rect 2925 6113 2929 6196
rect 2971 6188 2975 6196
rect 2960 6184 2975 6188
rect 2991 6184 2995 6196
rect 2960 6153 2966 6184
rect 2980 6180 2995 6184
rect 2980 6173 2986 6180
rect 2966 6141 2976 6153
rect 2925 6101 2934 6113
rect 2862 6064 2866 6072
rect 2925 6044 2929 6101
rect 2972 6084 2976 6141
rect 2980 6084 2984 6161
rect 3011 6153 3015 6196
rect 2988 6141 2995 6153
rect 3007 6141 3015 6153
rect 2988 6084 2992 6141
rect 3085 6099 3089 6156
rect 3105 6142 3109 6156
rect 3125 6142 3129 6156
rect 3185 6153 3189 6196
rect 3205 6184 3209 6196
rect 3225 6188 3229 6196
rect 3225 6184 3240 6188
rect 3205 6180 3220 6184
rect 3214 6173 3220 6180
rect 3105 6136 3120 6142
rect 3125 6136 3141 6142
rect 3185 6141 3193 6153
rect 3205 6141 3212 6153
rect 3114 6113 3120 6136
rect 3085 6087 3094 6099
rect 3092 6044 3096 6087
rect 3114 6064 3118 6101
rect 3134 6099 3141 6136
rect 3134 6074 3141 6087
rect 3208 6084 3212 6141
rect 3216 6084 3220 6161
rect 3234 6153 3240 6184
rect 3224 6141 3234 6153
rect 3224 6084 3228 6141
rect 3285 6099 3289 6156
rect 3305 6142 3309 6156
rect 3325 6142 3329 6156
rect 3305 6136 3320 6142
rect 3325 6136 3341 6142
rect 3314 6113 3320 6136
rect 3285 6087 3294 6099
rect 3122 6068 3141 6074
rect 3122 6064 3126 6068
rect 3292 6044 3296 6087
rect 3314 6064 3318 6101
rect 3334 6099 3341 6136
rect 3385 6113 3389 6196
rect 3445 6153 3449 6196
rect 3465 6184 3469 6196
rect 3485 6188 3489 6196
rect 3531 6188 3535 6196
rect 3485 6184 3500 6188
rect 3465 6180 3480 6184
rect 3474 6173 3480 6180
rect 3445 6141 3453 6153
rect 3465 6141 3472 6153
rect 3385 6101 3394 6113
rect 3334 6074 3341 6087
rect 3322 6068 3341 6074
rect 3322 6064 3326 6068
rect 3385 6044 3389 6101
rect 3468 6084 3472 6141
rect 3476 6084 3480 6161
rect 3494 6153 3500 6184
rect 3520 6184 3535 6188
rect 3551 6184 3555 6196
rect 3520 6153 3526 6184
rect 3540 6180 3555 6184
rect 3540 6173 3546 6180
rect 3484 6141 3494 6153
rect 3526 6141 3536 6153
rect 3484 6084 3488 6141
rect 3532 6084 3536 6141
rect 3540 6084 3544 6161
rect 3571 6153 3575 6196
rect 3548 6141 3555 6153
rect 3567 6141 3575 6153
rect 3548 6084 3552 6141
rect 3631 6113 3635 6196
rect 3691 6142 3695 6156
rect 3711 6142 3715 6156
rect 3626 6101 3635 6113
rect 3631 6044 3635 6101
rect 3679 6136 3695 6142
rect 3700 6136 3715 6142
rect 3679 6099 3686 6136
rect 3700 6113 3706 6136
rect 3679 6074 3686 6087
rect 3679 6068 3698 6074
rect 3694 6064 3698 6068
rect 3702 6064 3706 6101
rect 3731 6099 3735 6156
rect 3805 6119 3809 6196
rect 3806 6107 3809 6119
rect 3726 6087 3735 6099
rect 3803 6091 3809 6107
rect 3825 6119 3829 6196
rect 3871 6119 3875 6196
rect 3825 6107 3834 6119
rect 3866 6107 3875 6119
rect 3825 6091 3831 6107
rect 3724 6044 3728 6087
rect 3803 6084 3817 6091
rect 3813 6064 3817 6084
rect 3823 6084 3831 6091
rect 3869 6091 3875 6107
rect 3891 6119 3895 6196
rect 3970 6153 3974 6196
rect 3967 6141 3974 6153
rect 3891 6107 3894 6119
rect 3891 6091 3897 6107
rect 3869 6084 3877 6091
rect 3823 6064 3827 6084
rect 3873 6064 3877 6084
rect 3883 6084 3897 6091
rect 3883 6064 3887 6084
rect 3965 6064 3969 6141
rect 3992 6099 3996 6156
rect 4000 6152 4004 6156
rect 4056 6152 4060 6156
rect 4000 6144 4018 6152
rect 4014 6133 4018 6144
rect 4042 6144 4060 6152
rect 4042 6133 4046 6144
rect 3985 6087 3994 6099
rect 3985 6064 3989 6087
rect 4014 6076 4018 6121
rect 4005 6069 4018 6076
rect 4042 6076 4046 6121
rect 4064 6099 4068 6156
rect 4086 6153 4090 6196
rect 4086 6141 4093 6153
rect 4066 6087 4075 6099
rect 4042 6069 4055 6076
rect 4005 6064 4009 6069
rect 4051 6064 4055 6069
rect 4071 6064 4075 6087
rect 4091 6064 4095 6141
rect 4177 6133 4181 6156
rect 4166 6121 4181 6133
rect 4185 6133 4189 6156
rect 4185 6121 4194 6133
rect 4165 6044 4169 6121
rect 4185 6044 4189 6121
rect 4231 6113 4235 6196
rect 4305 6119 4309 6196
rect 4226 6101 4235 6113
rect 4306 6107 4309 6119
rect 4231 6044 4235 6101
rect 4303 6091 4309 6107
rect 4325 6119 4329 6196
rect 4371 6133 4375 6196
rect 4366 6121 4375 6133
rect 4325 6107 4334 6119
rect 4325 6091 4331 6107
rect 4303 6084 4317 6091
rect 4313 6064 4317 6084
rect 4323 6084 4331 6091
rect 4323 6064 4327 6084
rect 4371 6064 4375 6121
rect 4393 6119 4397 6196
rect 4381 6107 4394 6119
rect 4381 6064 4385 6107
rect 4415 6082 4419 6156
rect 4490 6153 4494 6196
rect 4671 6188 4675 6196
rect 4660 6184 4675 6188
rect 4691 6184 4695 6196
rect 4487 6141 4494 6153
rect 4407 6070 4419 6082
rect 4401 6064 4405 6070
rect 4485 6064 4489 6141
rect 4512 6099 4516 6156
rect 4520 6152 4524 6156
rect 4520 6144 4538 6152
rect 4534 6133 4538 6144
rect 4505 6087 4514 6099
rect 4505 6064 4509 6087
rect 4534 6076 4538 6121
rect 4585 6099 4589 6156
rect 4605 6142 4609 6156
rect 4625 6142 4629 6156
rect 4660 6153 4666 6184
rect 4680 6180 4695 6184
rect 4680 6173 4686 6180
rect 4605 6136 4620 6142
rect 4625 6136 4641 6142
rect 4666 6141 4676 6153
rect 4614 6113 4620 6136
rect 4585 6087 4594 6099
rect 4525 6069 4538 6076
rect 4525 6064 4529 6069
rect 4592 6044 4596 6087
rect 4614 6064 4618 6101
rect 4634 6099 4641 6136
rect 4634 6074 4641 6087
rect 4672 6084 4676 6141
rect 4680 6084 4684 6161
rect 4711 6153 4715 6196
rect 4688 6141 4695 6153
rect 4707 6141 4715 6153
rect 4688 6084 4692 6141
rect 4785 6099 4789 6156
rect 4805 6142 4809 6156
rect 4825 6142 4829 6156
rect 4885 6153 4889 6196
rect 4905 6184 4909 6196
rect 4925 6188 4929 6196
rect 4971 6188 4975 6196
rect 4925 6184 4940 6188
rect 4905 6180 4920 6184
rect 4914 6173 4920 6180
rect 4805 6136 4820 6142
rect 4825 6136 4841 6142
rect 4885 6141 4893 6153
rect 4905 6141 4912 6153
rect 4814 6113 4820 6136
rect 4785 6087 4794 6099
rect 4622 6068 4641 6074
rect 4622 6064 4626 6068
rect 4792 6044 4796 6087
rect 4814 6064 4818 6101
rect 4834 6099 4841 6136
rect 4834 6074 4841 6087
rect 4908 6084 4912 6141
rect 4916 6084 4920 6161
rect 4934 6153 4940 6184
rect 4960 6184 4975 6188
rect 4991 6184 4995 6196
rect 4960 6153 4966 6184
rect 4980 6180 4995 6184
rect 4980 6173 4986 6180
rect 4924 6141 4934 6153
rect 4966 6141 4976 6153
rect 4924 6084 4928 6141
rect 4972 6084 4976 6141
rect 4980 6084 4984 6161
rect 5011 6153 5015 6196
rect 5090 6153 5094 6196
rect 4988 6141 4995 6153
rect 5007 6141 5015 6153
rect 5087 6141 5094 6153
rect 4988 6084 4992 6141
rect 4822 6068 4841 6074
rect 4822 6064 4826 6068
rect 5085 6064 5089 6141
rect 5112 6099 5116 6156
rect 5120 6152 5124 6156
rect 5120 6144 5138 6152
rect 5134 6133 5138 6144
rect 5105 6087 5114 6099
rect 5105 6064 5109 6087
rect 5134 6076 5138 6121
rect 5185 6119 5189 6196
rect 5186 6107 5189 6119
rect 5183 6091 5189 6107
rect 5205 6119 5209 6196
rect 5251 6133 5255 6196
rect 5246 6121 5255 6133
rect 5205 6107 5214 6119
rect 5205 6091 5211 6107
rect 5183 6084 5197 6091
rect 5125 6069 5138 6076
rect 5125 6064 5129 6069
rect 5193 6064 5197 6084
rect 5203 6084 5211 6091
rect 5203 6064 5207 6084
rect 5251 6064 5255 6121
rect 5273 6119 5277 6196
rect 5261 6107 5274 6119
rect 5261 6064 5265 6107
rect 5295 6082 5299 6156
rect 5356 6152 5360 6156
rect 5342 6144 5360 6152
rect 5342 6133 5346 6144
rect 5287 6070 5299 6082
rect 5342 6076 5346 6121
rect 5364 6099 5368 6156
rect 5386 6153 5390 6196
rect 5386 6141 5393 6153
rect 5366 6087 5375 6099
rect 5281 6064 5285 6070
rect 5342 6069 5355 6076
rect 5351 6064 5355 6069
rect 5371 6064 5375 6087
rect 5391 6064 5395 6141
rect 5465 6099 5469 6156
rect 5485 6142 5489 6156
rect 5505 6142 5509 6156
rect 5565 6153 5569 6196
rect 5585 6184 5589 6196
rect 5605 6188 5609 6196
rect 5651 6188 5655 6196
rect 5605 6184 5620 6188
rect 5585 6180 5600 6184
rect 5594 6173 5600 6180
rect 5485 6136 5500 6142
rect 5505 6136 5521 6142
rect 5565 6141 5573 6153
rect 5585 6141 5592 6153
rect 5494 6113 5500 6136
rect 5465 6087 5474 6099
rect 5472 6044 5476 6087
rect 5494 6064 5498 6101
rect 5514 6099 5521 6136
rect 5514 6074 5521 6087
rect 5588 6084 5592 6141
rect 5596 6084 5600 6161
rect 5614 6153 5620 6184
rect 5640 6184 5655 6188
rect 5671 6184 5675 6196
rect 5640 6153 5646 6184
rect 5660 6180 5675 6184
rect 5660 6173 5666 6180
rect 5604 6141 5614 6153
rect 5646 6141 5656 6153
rect 5604 6084 5608 6141
rect 5652 6084 5656 6141
rect 5660 6084 5664 6161
rect 5691 6153 5695 6196
rect 5851 6188 5855 6196
rect 5840 6184 5855 6188
rect 5871 6184 5875 6196
rect 5668 6141 5675 6153
rect 5687 6141 5695 6153
rect 5668 6084 5672 6141
rect 5765 6099 5769 6156
rect 5785 6142 5789 6156
rect 5805 6142 5809 6156
rect 5840 6153 5846 6184
rect 5860 6180 5875 6184
rect 5860 6173 5866 6180
rect 5785 6136 5800 6142
rect 5805 6136 5821 6142
rect 5846 6141 5856 6153
rect 5794 6113 5800 6136
rect 5765 6087 5774 6099
rect 5502 6068 5521 6074
rect 5502 6064 5506 6068
rect 5772 6044 5776 6087
rect 5794 6064 5798 6101
rect 5814 6099 5821 6136
rect 5814 6074 5821 6087
rect 5852 6084 5856 6141
rect 5860 6084 5864 6161
rect 5891 6153 5895 6196
rect 5868 6141 5875 6153
rect 5887 6141 5895 6153
rect 5956 6152 5960 6156
rect 5942 6144 5960 6152
rect 5868 6084 5872 6141
rect 5942 6133 5946 6144
rect 5802 6068 5821 6074
rect 5802 6064 5806 6068
rect 5942 6076 5946 6121
rect 5964 6099 5968 6156
rect 5986 6153 5990 6196
rect 5986 6141 5993 6153
rect 6056 6152 6060 6156
rect 6042 6144 6060 6152
rect 5966 6087 5975 6099
rect 5942 6069 5955 6076
rect 5951 6064 5955 6069
rect 5971 6064 5975 6087
rect 5991 6064 5995 6141
rect 6042 6133 6046 6144
rect 6042 6076 6046 6121
rect 6064 6099 6068 6156
rect 6086 6153 6090 6196
rect 6151 6188 6155 6196
rect 6140 6184 6155 6188
rect 6171 6184 6175 6196
rect 6140 6153 6146 6184
rect 6160 6180 6175 6184
rect 6160 6173 6166 6180
rect 6086 6141 6093 6153
rect 6146 6141 6156 6153
rect 6066 6087 6075 6099
rect 6042 6069 6055 6076
rect 6051 6064 6055 6069
rect 6071 6064 6075 6087
rect 6091 6064 6095 6141
rect 6152 6084 6156 6141
rect 6160 6084 6164 6161
rect 6191 6153 6195 6196
rect 6251 6188 6255 6196
rect 6240 6184 6255 6188
rect 6271 6184 6275 6196
rect 6240 6153 6246 6184
rect 6260 6180 6275 6184
rect 6260 6173 6266 6180
rect 6168 6141 6175 6153
rect 6187 6141 6195 6153
rect 6246 6141 6256 6153
rect 6168 6084 6172 6141
rect 6252 6084 6256 6141
rect 6260 6084 6264 6161
rect 6291 6153 6295 6196
rect 6268 6141 6275 6153
rect 6287 6141 6295 6153
rect 6365 6153 6369 6196
rect 6385 6184 6389 6196
rect 6405 6188 6409 6196
rect 6405 6184 6420 6188
rect 6385 6180 6400 6184
rect 6394 6173 6400 6180
rect 6365 6141 6373 6153
rect 6385 6141 6392 6153
rect 6268 6084 6272 6141
rect 6388 6084 6392 6141
rect 6396 6084 6400 6161
rect 6414 6153 6420 6184
rect 6404 6141 6414 6153
rect 6404 6084 6408 6141
rect 6465 6099 6469 6156
rect 6485 6142 6489 6156
rect 6505 6142 6509 6156
rect 6485 6136 6500 6142
rect 6505 6136 6521 6142
rect 6494 6113 6500 6136
rect 6465 6087 6474 6099
rect 6472 6044 6476 6087
rect 6494 6064 6498 6101
rect 6514 6099 6521 6136
rect 6551 6113 6555 6196
rect 6611 6113 6615 6196
rect 6546 6101 6555 6113
rect 6606 6101 6615 6113
rect 6514 6074 6521 6087
rect 6502 6068 6521 6074
rect 6502 6064 6506 6068
rect 6551 6044 6555 6101
rect 6611 6044 6615 6101
rect 31 6020 35 6024
rect 53 6020 57 6024
rect 63 6020 67 6024
rect 83 6020 87 6024
rect 91 6020 95 6024
rect 137 6020 141 6024
rect 159 6020 163 6024
rect 169 6020 173 6024
rect 191 6020 195 6024
rect 201 6020 205 6024
rect 221 6020 225 6024
rect 292 6020 296 6024
rect 314 6020 318 6024
rect 322 6020 326 6024
rect 393 6020 397 6024
rect 403 6020 407 6024
rect 451 6020 455 6024
rect 471 6020 475 6024
rect 553 6020 557 6024
rect 563 6020 567 6024
rect 611 6020 615 6024
rect 631 6020 635 6024
rect 651 6020 655 6024
rect 725 6020 729 6024
rect 745 6020 749 6024
rect 765 6020 769 6024
rect 811 6020 815 6024
rect 831 6020 835 6024
rect 912 6020 916 6024
rect 934 6020 938 6024
rect 942 6020 946 6024
rect 991 6020 995 6024
rect 1011 6020 1015 6024
rect 1031 6020 1035 6024
rect 1105 6020 1109 6024
rect 1151 6020 1155 6024
rect 1171 6020 1175 6024
rect 1245 6020 1249 6024
rect 1265 6020 1269 6024
rect 1285 6020 1289 6024
rect 1345 6020 1349 6024
rect 1405 6020 1409 6024
rect 1451 6020 1455 6024
rect 1471 6020 1475 6024
rect 1531 6020 1535 6024
rect 1551 6020 1555 6024
rect 1611 6020 1615 6024
rect 1671 6020 1675 6024
rect 1691 6020 1695 6024
rect 1751 6020 1755 6024
rect 1771 6020 1775 6024
rect 1831 6020 1835 6024
rect 1851 6020 1855 6024
rect 1871 6020 1875 6024
rect 1931 6020 1935 6024
rect 2012 6020 2016 6024
rect 2034 6020 2038 6024
rect 2042 6020 2046 6024
rect 2091 6020 2095 6024
rect 2165 6020 2169 6024
rect 2185 6020 2189 6024
rect 2205 6020 2209 6024
rect 2251 6020 2255 6024
rect 2325 6020 2329 6024
rect 2345 6020 2349 6024
rect 2365 6020 2369 6024
rect 2448 6020 2452 6024
rect 2456 6020 2460 6024
rect 2464 6020 2468 6024
rect 2532 6020 2536 6024
rect 2554 6020 2558 6024
rect 2562 6020 2566 6024
rect 2625 6020 2629 6024
rect 2645 6020 2649 6024
rect 2728 6020 2732 6024
rect 2736 6020 2740 6024
rect 2744 6020 2748 6024
rect 2826 6020 2830 6024
rect 2834 6020 2838 6024
rect 2854 6020 2858 6024
rect 2862 6020 2866 6024
rect 2925 6020 2929 6024
rect 2972 6020 2976 6024
rect 2980 6020 2984 6024
rect 2988 6020 2992 6024
rect 3092 6020 3096 6024
rect 3114 6020 3118 6024
rect 3122 6020 3126 6024
rect 3208 6020 3212 6024
rect 3216 6020 3220 6024
rect 3224 6020 3228 6024
rect 3292 6020 3296 6024
rect 3314 6020 3318 6024
rect 3322 6020 3326 6024
rect 3385 6020 3389 6024
rect 3468 6020 3472 6024
rect 3476 6020 3480 6024
rect 3484 6020 3488 6024
rect 3532 6020 3536 6024
rect 3540 6020 3544 6024
rect 3548 6020 3552 6024
rect 3631 6020 3635 6024
rect 3694 6020 3698 6024
rect 3702 6020 3706 6024
rect 3724 6020 3728 6024
rect 3813 6020 3817 6024
rect 3823 6020 3827 6024
rect 3873 6020 3877 6024
rect 3883 6020 3887 6024
rect 3965 6020 3969 6024
rect 3985 6020 3989 6024
rect 4005 6020 4009 6024
rect 4051 6020 4055 6024
rect 4071 6020 4075 6024
rect 4091 6020 4095 6024
rect 4165 6020 4169 6024
rect 4185 6020 4189 6024
rect 4231 6020 4235 6024
rect 4313 6020 4317 6024
rect 4323 6020 4327 6024
rect 4371 6020 4375 6024
rect 4381 6020 4385 6024
rect 4401 6020 4405 6024
rect 4485 6020 4489 6024
rect 4505 6020 4509 6024
rect 4525 6020 4529 6024
rect 4592 6020 4596 6024
rect 4614 6020 4618 6024
rect 4622 6020 4626 6024
rect 4672 6020 4676 6024
rect 4680 6020 4684 6024
rect 4688 6020 4692 6024
rect 4792 6020 4796 6024
rect 4814 6020 4818 6024
rect 4822 6020 4826 6024
rect 4908 6020 4912 6024
rect 4916 6020 4920 6024
rect 4924 6020 4928 6024
rect 4972 6020 4976 6024
rect 4980 6020 4984 6024
rect 4988 6020 4992 6024
rect 5085 6020 5089 6024
rect 5105 6020 5109 6024
rect 5125 6020 5129 6024
rect 5193 6020 5197 6024
rect 5203 6020 5207 6024
rect 5251 6020 5255 6024
rect 5261 6020 5265 6024
rect 5281 6020 5285 6024
rect 5351 6020 5355 6024
rect 5371 6020 5375 6024
rect 5391 6020 5395 6024
rect 5472 6020 5476 6024
rect 5494 6020 5498 6024
rect 5502 6020 5506 6024
rect 5588 6020 5592 6024
rect 5596 6020 5600 6024
rect 5604 6020 5608 6024
rect 5652 6020 5656 6024
rect 5660 6020 5664 6024
rect 5668 6020 5672 6024
rect 5772 6020 5776 6024
rect 5794 6020 5798 6024
rect 5802 6020 5806 6024
rect 5852 6020 5856 6024
rect 5860 6020 5864 6024
rect 5868 6020 5872 6024
rect 5951 6020 5955 6024
rect 5971 6020 5975 6024
rect 5991 6020 5995 6024
rect 6051 6020 6055 6024
rect 6071 6020 6075 6024
rect 6091 6020 6095 6024
rect 6152 6020 6156 6024
rect 6160 6020 6164 6024
rect 6168 6020 6172 6024
rect 6252 6020 6256 6024
rect 6260 6020 6264 6024
rect 6268 6020 6272 6024
rect 6388 6020 6392 6024
rect 6396 6020 6400 6024
rect 6404 6020 6408 6024
rect 6472 6020 6476 6024
rect 6494 6020 6498 6024
rect 6502 6020 6506 6024
rect 6551 6020 6555 6024
rect 6611 6020 6615 6024
rect 43 5996 47 6000
rect 65 5996 69 6000
rect 113 5996 117 6000
rect 123 5996 127 6000
rect 193 5996 197 6000
rect 203 5996 207 6000
rect 292 5996 296 6000
rect 314 5996 318 6000
rect 322 5996 326 6000
rect 393 5996 397 6000
rect 403 5996 407 6000
rect 451 5996 455 6000
rect 525 5996 529 6000
rect 545 5996 549 6000
rect 591 5996 595 6000
rect 611 5996 615 6000
rect 671 5996 675 6000
rect 691 5996 695 6000
rect 711 5996 715 6000
rect 785 5996 789 6000
rect 831 5996 835 6000
rect 851 5996 855 6000
rect 933 5996 937 6000
rect 943 5996 947 6000
rect 1005 5996 1009 6000
rect 1025 5996 1029 6000
rect 1045 5996 1049 6000
rect 1091 5996 1095 6000
rect 1111 5996 1115 6000
rect 1185 5996 1189 6000
rect 1231 5996 1235 6000
rect 1253 5996 1257 6000
rect 1263 5996 1267 6000
rect 1283 5996 1287 6000
rect 1291 5996 1295 6000
rect 1337 5996 1341 6000
rect 1359 5996 1363 6000
rect 1369 5996 1373 6000
rect 1391 5996 1395 6000
rect 1401 5996 1405 6000
rect 1421 5996 1425 6000
rect 1473 5996 1477 6000
rect 1483 5996 1487 6000
rect 1588 5996 1592 6000
rect 1596 5996 1600 6000
rect 1604 5996 1608 6000
rect 1665 5996 1669 6000
rect 1685 5996 1689 6000
rect 1705 5996 1709 6000
rect 1765 5996 1769 6000
rect 1785 5996 1789 6000
rect 1868 5996 1872 6000
rect 1876 5996 1880 6000
rect 1884 5996 1888 6000
rect 1931 5996 1935 6000
rect 2005 5996 2009 6000
rect 2025 5996 2029 6000
rect 2045 5996 2049 6000
rect 2092 5996 2096 6000
rect 2100 5996 2104 6000
rect 2108 5996 2112 6000
rect 2212 5996 2216 6000
rect 2234 5996 2238 6000
rect 2242 5996 2246 6000
rect 2291 5996 2295 6000
rect 2311 5996 2315 6000
rect 2331 5996 2335 6000
rect 2413 5996 2417 6000
rect 2423 5996 2427 6000
rect 2508 5996 2512 6000
rect 2516 5996 2520 6000
rect 2524 5996 2528 6000
rect 2592 5996 2596 6000
rect 2614 5996 2618 6000
rect 2622 5996 2626 6000
rect 2673 5996 2677 6000
rect 2683 5996 2687 6000
rect 2788 5996 2792 6000
rect 2796 5996 2800 6000
rect 2804 5996 2808 6000
rect 2888 5996 2892 6000
rect 2896 5996 2900 6000
rect 2904 5996 2908 6000
rect 2988 5996 2992 6000
rect 2996 5996 3000 6000
rect 3004 5996 3008 6000
rect 3088 5996 3092 6000
rect 3096 5996 3100 6000
rect 3104 5996 3108 6000
rect 3152 5996 3156 6000
rect 3160 5996 3164 6000
rect 3168 5996 3172 6000
rect 3265 5996 3269 6000
rect 3285 5996 3289 6000
rect 3305 5996 3309 6000
rect 3351 5996 3355 6000
rect 3371 5996 3375 6000
rect 3391 5996 3395 6000
rect 3472 5996 3476 6000
rect 3494 5996 3498 6000
rect 3502 5996 3506 6000
rect 3565 5996 3569 6000
rect 3585 5996 3589 6000
rect 3605 5996 3609 6000
rect 3688 5996 3692 6000
rect 3696 5996 3700 6000
rect 3704 5996 3708 6000
rect 3754 5996 3758 6000
rect 3762 5996 3766 6000
rect 3784 5996 3788 6000
rect 3888 5996 3892 6000
rect 3896 5996 3900 6000
rect 3904 5996 3908 6000
rect 3972 5996 3976 6000
rect 3994 5996 3998 6000
rect 4002 5996 4006 6000
rect 4088 5996 4092 6000
rect 4096 5996 4100 6000
rect 4104 5996 4108 6000
rect 4172 5996 4176 6000
rect 4194 5996 4198 6000
rect 4202 5996 4206 6000
rect 4252 5996 4256 6000
rect 4260 5996 4264 6000
rect 4268 5996 4272 6000
rect 4353 5996 4357 6000
rect 4363 5996 4367 6000
rect 4445 5996 4449 6000
rect 4465 5996 4469 6000
rect 4485 5996 4489 6000
rect 4545 5996 4549 6000
rect 4565 5996 4569 6000
rect 4611 5996 4615 6000
rect 4621 5996 4625 6000
rect 4641 5996 4645 6000
rect 4732 5996 4736 6000
rect 4754 5996 4758 6000
rect 4762 5996 4766 6000
rect 4813 5996 4817 6000
rect 4823 5996 4827 6000
rect 4905 5996 4909 6000
rect 4988 5996 4992 6000
rect 4996 5996 5000 6000
rect 5004 5996 5008 6000
rect 5054 5996 5058 6000
rect 5062 5996 5066 6000
rect 5084 5996 5088 6000
rect 5151 5996 5155 6000
rect 5171 5996 5175 6000
rect 5191 5996 5195 6000
rect 5251 5996 5255 6000
rect 5271 5996 5275 6000
rect 5291 5996 5295 6000
rect 5354 5996 5358 6000
rect 5362 5996 5366 6000
rect 5382 5996 5386 6000
rect 5390 5996 5394 6000
rect 5493 5996 5497 6000
rect 5503 5996 5507 6000
rect 5551 5996 5555 6000
rect 5648 5996 5652 6000
rect 5656 5996 5660 6000
rect 5664 5996 5668 6000
rect 5714 5996 5718 6000
rect 5722 5996 5726 6000
rect 5744 5996 5748 6000
rect 5825 5996 5829 6000
rect 5845 5996 5849 6000
rect 5865 5996 5869 6000
rect 5911 5996 5915 6000
rect 5931 5996 5935 6000
rect 5951 5996 5955 6000
rect 6025 5996 6029 6000
rect 6045 5996 6049 6000
rect 6065 5996 6069 6000
rect 6114 5996 6118 6000
rect 6122 5996 6126 6000
rect 6142 5996 6146 6000
rect 6150 5996 6154 6000
rect 6253 5996 6257 6000
rect 6263 5996 6267 6000
rect 6311 5996 6315 6000
rect 6321 5996 6325 6000
rect 6341 5996 6345 6000
rect 6411 5996 6415 6000
rect 6431 5996 6435 6000
rect 6451 5996 6455 6000
rect 6512 5996 6516 6000
rect 6520 5996 6524 6000
rect 6528 5996 6532 6000
rect 6613 5996 6617 6000
rect 6623 5996 6627 6000
rect 43 5950 47 5956
rect 43 5938 45 5950
rect 65 5899 69 5976
rect 113 5936 117 5956
rect 109 5929 117 5936
rect 123 5936 127 5956
rect 193 5936 197 5956
rect 123 5929 137 5936
rect 109 5913 115 5929
rect 106 5901 115 5913
rect 65 5887 74 5899
rect 43 5870 45 5882
rect 43 5864 47 5870
rect 65 5824 69 5887
rect 111 5824 115 5901
rect 131 5913 137 5929
rect 189 5929 197 5936
rect 203 5936 207 5956
rect 203 5929 217 5936
rect 292 5933 296 5976
rect 189 5913 195 5929
rect 131 5901 134 5913
rect 186 5901 195 5913
rect 131 5824 135 5901
rect 191 5824 195 5901
rect 211 5913 217 5929
rect 285 5921 294 5933
rect 211 5901 214 5913
rect 211 5824 215 5901
rect 285 5864 289 5921
rect 314 5919 318 5956
rect 322 5952 326 5956
rect 322 5946 341 5952
rect 334 5933 341 5946
rect 393 5936 397 5956
rect 383 5929 397 5936
rect 403 5936 407 5956
rect 403 5929 411 5936
rect 314 5884 320 5907
rect 334 5884 341 5921
rect 383 5913 389 5929
rect 386 5901 389 5913
rect 305 5878 320 5884
rect 325 5878 341 5884
rect 305 5864 309 5878
rect 325 5864 329 5878
rect 385 5824 389 5901
rect 405 5913 411 5929
rect 451 5919 455 5976
rect 405 5901 414 5913
rect 446 5907 455 5919
rect 405 5824 409 5901
rect 451 5824 455 5907
rect 525 5899 529 5976
rect 545 5899 549 5976
rect 591 5899 595 5976
rect 611 5899 615 5976
rect 671 5951 675 5956
rect 662 5944 675 5951
rect 662 5899 666 5944
rect 691 5933 695 5956
rect 686 5921 695 5933
rect 526 5887 541 5899
rect 537 5864 541 5887
rect 545 5887 554 5899
rect 586 5887 595 5899
rect 545 5864 549 5887
rect 591 5864 595 5887
rect 599 5887 614 5899
rect 599 5864 603 5887
rect 662 5876 666 5887
rect 662 5868 680 5876
rect 676 5864 680 5868
rect 684 5864 688 5921
rect 711 5879 715 5956
rect 785 5919 789 5976
rect 785 5907 794 5919
rect 706 5867 713 5879
rect 706 5824 710 5867
rect 785 5824 789 5907
rect 831 5899 835 5976
rect 851 5899 855 5976
rect 933 5936 937 5956
rect 923 5929 937 5936
rect 943 5936 947 5956
rect 943 5929 951 5936
rect 923 5913 929 5929
rect 926 5901 929 5913
rect 826 5887 835 5899
rect 831 5864 835 5887
rect 839 5887 854 5899
rect 839 5864 843 5887
rect 925 5824 929 5901
rect 945 5913 951 5929
rect 945 5901 954 5913
rect 945 5824 949 5901
rect 1005 5879 1009 5956
rect 1025 5933 1029 5956
rect 1045 5951 1049 5956
rect 1045 5944 1058 5951
rect 1025 5921 1034 5933
rect 1007 5867 1014 5879
rect 1010 5824 1014 5867
rect 1032 5864 1036 5921
rect 1054 5899 1058 5944
rect 1091 5899 1095 5976
rect 1111 5899 1115 5976
rect 1185 5919 1189 5976
rect 1185 5907 1194 5919
rect 1086 5887 1095 5899
rect 1054 5876 1058 5887
rect 1040 5868 1058 5876
rect 1040 5864 1044 5868
rect 1091 5864 1095 5887
rect 1099 5887 1114 5899
rect 1099 5864 1103 5887
rect 1185 5824 1189 5907
rect 1231 5888 1235 5956
rect 1253 5927 1257 5976
rect 1263 5955 1267 5976
rect 1283 5964 1287 5976
rect 1291 5972 1295 5976
rect 1291 5968 1325 5972
rect 1283 5960 1313 5964
rect 1283 5959 1301 5960
rect 1263 5951 1287 5955
rect 1231 5876 1233 5888
rect 1231 5864 1235 5876
rect 1253 5869 1257 5915
rect 1249 5863 1257 5869
rect 1249 5834 1253 5863
rect 1281 5856 1287 5951
rect 1249 5827 1257 5834
rect 1253 5804 1257 5827
rect 1261 5804 1265 5844
rect 1281 5824 1285 5856
rect 1321 5842 1325 5968
rect 1337 5862 1341 5976
rect 1359 5964 1363 5976
rect 1361 5952 1363 5964
rect 1369 5964 1373 5976
rect 1369 5952 1371 5964
rect 1289 5830 1313 5832
rect 1289 5828 1325 5830
rect 1289 5824 1293 5828
rect 1335 5824 1339 5850
rect 1353 5842 1357 5952
rect 1391 5944 1395 5976
rect 1362 5940 1395 5944
rect 1362 5876 1366 5940
rect 1382 5891 1386 5920
rect 1401 5918 1405 5976
rect 1421 5919 1425 5956
rect 1473 5936 1477 5956
rect 1469 5929 1477 5936
rect 1483 5936 1487 5956
rect 1483 5929 1497 5936
rect 1469 5913 1475 5929
rect 1382 5883 1391 5891
rect 1362 5864 1365 5876
rect 1355 5824 1359 5830
rect 1367 5824 1371 5864
rect 1387 5824 1391 5883
rect 1401 5824 1405 5906
rect 1421 5864 1425 5907
rect 1466 5901 1475 5913
rect 1471 5824 1475 5901
rect 1491 5913 1497 5929
rect 1491 5901 1494 5913
rect 1491 5824 1495 5901
rect 1588 5879 1592 5936
rect 1565 5867 1573 5879
rect 1585 5867 1592 5879
rect 1565 5824 1569 5867
rect 1596 5859 1600 5936
rect 1604 5879 1608 5936
rect 1665 5879 1669 5956
rect 1685 5933 1689 5956
rect 1705 5951 1709 5956
rect 1705 5944 1718 5951
rect 1685 5921 1694 5933
rect 1604 5867 1614 5879
rect 1667 5867 1674 5879
rect 1594 5840 1600 5847
rect 1585 5836 1600 5840
rect 1614 5836 1620 5867
rect 1585 5824 1589 5836
rect 1605 5832 1620 5836
rect 1605 5824 1609 5832
rect 1670 5824 1674 5867
rect 1692 5864 1696 5921
rect 1714 5899 1718 5944
rect 1765 5899 1769 5976
rect 1785 5899 1789 5976
rect 1766 5887 1781 5899
rect 1714 5876 1718 5887
rect 1700 5868 1718 5876
rect 1700 5864 1704 5868
rect 1777 5864 1781 5887
rect 1785 5887 1794 5899
rect 1785 5864 1789 5887
rect 1868 5879 1872 5936
rect 1845 5867 1853 5879
rect 1865 5867 1872 5879
rect 1845 5824 1849 5867
rect 1876 5859 1880 5936
rect 1884 5879 1888 5936
rect 1931 5919 1935 5976
rect 1926 5907 1935 5919
rect 1884 5867 1894 5879
rect 1874 5840 1880 5847
rect 1865 5836 1880 5840
rect 1894 5836 1900 5867
rect 1865 5824 1869 5836
rect 1885 5832 1900 5836
rect 1885 5824 1889 5832
rect 1931 5824 1935 5907
rect 2005 5879 2009 5956
rect 2025 5933 2029 5956
rect 2045 5951 2049 5956
rect 2045 5944 2058 5951
rect 2025 5921 2034 5933
rect 2007 5867 2014 5879
rect 2010 5824 2014 5867
rect 2032 5864 2036 5921
rect 2054 5899 2058 5944
rect 2054 5876 2058 5887
rect 2092 5879 2096 5936
rect 2040 5868 2058 5876
rect 2040 5864 2044 5868
rect 2086 5867 2096 5879
rect 2080 5836 2086 5867
rect 2100 5859 2104 5936
rect 2108 5879 2112 5936
rect 2212 5933 2216 5976
rect 2205 5921 2214 5933
rect 2108 5867 2115 5879
rect 2127 5867 2135 5879
rect 2100 5840 2106 5847
rect 2100 5836 2115 5840
rect 2080 5832 2095 5836
rect 2091 5824 2095 5832
rect 2111 5824 2115 5836
rect 2131 5824 2135 5867
rect 2205 5864 2209 5921
rect 2234 5919 2238 5956
rect 2242 5952 2246 5956
rect 2242 5946 2261 5952
rect 2291 5951 2295 5956
rect 2254 5933 2261 5946
rect 2282 5944 2295 5951
rect 2234 5884 2240 5907
rect 2254 5884 2261 5921
rect 2282 5899 2286 5944
rect 2311 5933 2315 5956
rect 2306 5921 2315 5933
rect 2225 5878 2240 5884
rect 2245 5878 2261 5884
rect 2225 5864 2229 5878
rect 2245 5864 2249 5878
rect 2282 5876 2286 5887
rect 2282 5868 2300 5876
rect 2296 5864 2300 5868
rect 2304 5864 2308 5921
rect 2331 5879 2335 5956
rect 2413 5936 2417 5956
rect 2403 5929 2417 5936
rect 2423 5936 2427 5956
rect 2423 5929 2431 5936
rect 2403 5913 2409 5929
rect 2406 5901 2409 5913
rect 2326 5867 2333 5879
rect 2326 5824 2330 5867
rect 2405 5824 2409 5901
rect 2425 5913 2431 5929
rect 2425 5901 2434 5913
rect 2425 5824 2429 5901
rect 2508 5879 2512 5936
rect 2485 5867 2493 5879
rect 2505 5867 2512 5879
rect 2485 5824 2489 5867
rect 2516 5859 2520 5936
rect 2524 5879 2528 5936
rect 2592 5933 2596 5976
rect 2585 5921 2594 5933
rect 2524 5867 2534 5879
rect 2514 5840 2520 5847
rect 2505 5836 2520 5840
rect 2534 5836 2540 5867
rect 2585 5864 2589 5921
rect 2614 5919 2618 5956
rect 2622 5952 2626 5956
rect 2622 5946 2641 5952
rect 2634 5933 2641 5946
rect 2673 5936 2677 5956
rect 2669 5929 2677 5936
rect 2683 5936 2687 5956
rect 2683 5929 2697 5936
rect 2614 5884 2620 5907
rect 2634 5884 2641 5921
rect 2669 5913 2675 5929
rect 2666 5901 2675 5913
rect 2605 5878 2620 5884
rect 2625 5878 2641 5884
rect 2605 5864 2609 5878
rect 2625 5864 2629 5878
rect 2505 5824 2509 5836
rect 2525 5832 2540 5836
rect 2525 5824 2529 5832
rect 2671 5824 2675 5901
rect 2691 5913 2697 5929
rect 2691 5901 2694 5913
rect 2691 5824 2695 5901
rect 2788 5879 2792 5936
rect 2765 5867 2773 5879
rect 2785 5867 2792 5879
rect 2765 5824 2769 5867
rect 2796 5859 2800 5936
rect 2804 5879 2808 5936
rect 2888 5879 2892 5936
rect 2804 5867 2814 5879
rect 2865 5867 2873 5879
rect 2885 5867 2892 5879
rect 2794 5840 2800 5847
rect 2785 5836 2800 5840
rect 2814 5836 2820 5867
rect 2785 5824 2789 5836
rect 2805 5832 2820 5836
rect 2805 5824 2809 5832
rect 2865 5824 2869 5867
rect 2896 5859 2900 5936
rect 2904 5879 2908 5936
rect 2988 5879 2992 5936
rect 2904 5867 2914 5879
rect 2965 5867 2973 5879
rect 2985 5867 2992 5879
rect 2894 5840 2900 5847
rect 2885 5836 2900 5840
rect 2914 5836 2920 5867
rect 2885 5824 2889 5836
rect 2905 5832 2920 5836
rect 2905 5824 2909 5832
rect 2965 5824 2969 5867
rect 2996 5859 3000 5936
rect 3004 5879 3008 5936
rect 3088 5879 3092 5936
rect 3004 5867 3014 5879
rect 3065 5867 3073 5879
rect 3085 5867 3092 5879
rect 2994 5840 3000 5847
rect 2985 5836 3000 5840
rect 3014 5836 3020 5867
rect 2985 5824 2989 5836
rect 3005 5832 3020 5836
rect 3005 5824 3009 5832
rect 3065 5824 3069 5867
rect 3096 5859 3100 5936
rect 3104 5879 3108 5936
rect 3152 5879 3156 5936
rect 3104 5867 3114 5879
rect 3146 5867 3156 5879
rect 3094 5840 3100 5847
rect 3085 5836 3100 5840
rect 3114 5836 3120 5867
rect 3085 5824 3089 5836
rect 3105 5832 3120 5836
rect 3140 5836 3146 5867
rect 3160 5859 3164 5936
rect 3168 5879 3172 5936
rect 3265 5879 3269 5956
rect 3285 5933 3289 5956
rect 3305 5951 3309 5956
rect 3351 5951 3355 5956
rect 3305 5944 3318 5951
rect 3285 5921 3294 5933
rect 3168 5867 3175 5879
rect 3187 5867 3195 5879
rect 3267 5867 3274 5879
rect 3160 5840 3166 5847
rect 3160 5836 3175 5840
rect 3140 5832 3155 5836
rect 3105 5824 3109 5832
rect 3151 5824 3155 5832
rect 3171 5824 3175 5836
rect 3191 5824 3195 5867
rect 3270 5824 3274 5867
rect 3292 5864 3296 5921
rect 3314 5899 3318 5944
rect 3342 5944 3355 5951
rect 3342 5899 3346 5944
rect 3371 5933 3375 5956
rect 3366 5921 3375 5933
rect 3314 5876 3318 5887
rect 3300 5868 3318 5876
rect 3342 5876 3346 5887
rect 3342 5868 3360 5876
rect 3300 5864 3304 5868
rect 3356 5864 3360 5868
rect 3364 5864 3368 5921
rect 3391 5879 3395 5956
rect 3472 5933 3476 5976
rect 3465 5921 3474 5933
rect 3386 5867 3393 5879
rect 3386 5824 3390 5867
rect 3465 5864 3469 5921
rect 3494 5919 3498 5956
rect 3502 5952 3506 5956
rect 3502 5946 3521 5952
rect 3514 5933 3521 5946
rect 3494 5884 3500 5907
rect 3514 5884 3521 5921
rect 3485 5878 3500 5884
rect 3505 5878 3521 5884
rect 3565 5879 3569 5956
rect 3585 5933 3589 5956
rect 3605 5951 3609 5956
rect 3605 5944 3618 5951
rect 3585 5921 3594 5933
rect 3485 5864 3489 5878
rect 3505 5864 3509 5878
rect 3567 5867 3574 5879
rect 3570 5824 3574 5867
rect 3592 5864 3596 5921
rect 3614 5899 3618 5944
rect 3754 5952 3758 5956
rect 3739 5946 3758 5952
rect 3614 5876 3618 5887
rect 3688 5879 3692 5936
rect 3600 5868 3618 5876
rect 3600 5864 3604 5868
rect 3665 5867 3673 5879
rect 3685 5867 3692 5879
rect 3665 5824 3669 5867
rect 3696 5859 3700 5936
rect 3704 5879 3708 5936
rect 3739 5933 3746 5946
rect 3739 5884 3746 5921
rect 3762 5919 3766 5956
rect 3784 5933 3788 5976
rect 3786 5921 3795 5933
rect 3760 5884 3766 5907
rect 3704 5867 3714 5879
rect 3739 5878 3755 5884
rect 3760 5878 3775 5884
rect 3694 5840 3700 5847
rect 3685 5836 3700 5840
rect 3714 5836 3720 5867
rect 3751 5864 3755 5878
rect 3771 5864 3775 5878
rect 3791 5864 3795 5921
rect 3888 5879 3892 5936
rect 3865 5867 3873 5879
rect 3885 5867 3892 5879
rect 3685 5824 3689 5836
rect 3705 5832 3720 5836
rect 3705 5824 3709 5832
rect 3865 5824 3869 5867
rect 3896 5859 3900 5936
rect 3904 5879 3908 5936
rect 3972 5933 3976 5976
rect 3965 5921 3974 5933
rect 3904 5867 3914 5879
rect 3894 5840 3900 5847
rect 3885 5836 3900 5840
rect 3914 5836 3920 5867
rect 3965 5864 3969 5921
rect 3994 5919 3998 5956
rect 4002 5952 4006 5956
rect 4002 5946 4021 5952
rect 4014 5933 4021 5946
rect 3994 5884 4000 5907
rect 4014 5884 4021 5921
rect 3985 5878 4000 5884
rect 4005 5878 4021 5884
rect 4088 5879 4092 5936
rect 3985 5864 3989 5878
rect 4005 5864 4009 5878
rect 4065 5867 4073 5879
rect 4085 5867 4092 5879
rect 3885 5824 3889 5836
rect 3905 5832 3920 5836
rect 3905 5824 3909 5832
rect 4065 5824 4069 5867
rect 4096 5859 4100 5936
rect 4104 5879 4108 5936
rect 4172 5933 4176 5976
rect 4165 5921 4174 5933
rect 4104 5867 4114 5879
rect 4094 5840 4100 5847
rect 4085 5836 4100 5840
rect 4114 5836 4120 5867
rect 4165 5864 4169 5921
rect 4194 5919 4198 5956
rect 4202 5952 4206 5956
rect 4202 5946 4221 5952
rect 4214 5933 4221 5946
rect 4353 5936 4357 5956
rect 4194 5884 4200 5907
rect 4214 5884 4221 5921
rect 4185 5878 4200 5884
rect 4205 5878 4221 5884
rect 4252 5879 4256 5936
rect 4185 5864 4189 5878
rect 4205 5864 4209 5878
rect 4246 5867 4256 5879
rect 4085 5824 4089 5836
rect 4105 5832 4120 5836
rect 4105 5824 4109 5832
rect 4240 5836 4246 5867
rect 4260 5859 4264 5936
rect 4268 5879 4272 5936
rect 4349 5929 4357 5936
rect 4363 5936 4367 5956
rect 4363 5929 4377 5936
rect 4349 5913 4355 5929
rect 4346 5901 4355 5913
rect 4268 5867 4275 5879
rect 4287 5867 4295 5879
rect 4260 5840 4266 5847
rect 4260 5836 4275 5840
rect 4240 5832 4255 5836
rect 4251 5824 4255 5832
rect 4271 5824 4275 5836
rect 4291 5824 4295 5867
rect 4351 5824 4355 5901
rect 4371 5913 4377 5929
rect 4371 5901 4374 5913
rect 4371 5824 4375 5901
rect 4445 5879 4449 5956
rect 4465 5933 4469 5956
rect 4485 5951 4489 5956
rect 4485 5944 4498 5951
rect 4465 5921 4474 5933
rect 4447 5867 4454 5879
rect 4450 5824 4454 5867
rect 4472 5864 4476 5921
rect 4494 5899 4498 5944
rect 4545 5899 4549 5976
rect 4565 5899 4569 5976
rect 4611 5899 4615 5956
rect 4621 5913 4625 5956
rect 4641 5950 4645 5956
rect 4647 5938 4659 5950
rect 4621 5901 4634 5913
rect 4546 5887 4561 5899
rect 4494 5876 4498 5887
rect 4480 5868 4498 5876
rect 4480 5864 4484 5868
rect 4557 5864 4561 5887
rect 4565 5887 4574 5899
rect 4606 5887 4615 5899
rect 4565 5864 4569 5887
rect 4611 5824 4615 5887
rect 4633 5824 4637 5901
rect 4655 5864 4659 5938
rect 4732 5933 4736 5976
rect 4725 5921 4734 5933
rect 4725 5864 4729 5921
rect 4754 5919 4758 5956
rect 4762 5952 4766 5956
rect 4762 5946 4781 5952
rect 4774 5933 4781 5946
rect 4813 5936 4817 5956
rect 4809 5929 4817 5936
rect 4823 5936 4827 5956
rect 4823 5929 4837 5936
rect 4754 5884 4760 5907
rect 4774 5884 4781 5921
rect 4809 5913 4815 5929
rect 4806 5901 4815 5913
rect 4745 5878 4760 5884
rect 4765 5878 4781 5884
rect 4745 5864 4749 5878
rect 4765 5864 4769 5878
rect 4811 5824 4815 5901
rect 4831 5913 4837 5929
rect 4905 5919 4909 5976
rect 5054 5952 5058 5956
rect 5039 5946 5058 5952
rect 4831 5901 4834 5913
rect 4905 5907 4914 5919
rect 4831 5824 4835 5901
rect 4905 5824 4909 5907
rect 4988 5879 4992 5936
rect 4965 5867 4973 5879
rect 4985 5867 4992 5879
rect 4965 5824 4969 5867
rect 4996 5859 5000 5936
rect 5004 5879 5008 5936
rect 5039 5933 5046 5946
rect 5039 5884 5046 5921
rect 5062 5919 5066 5956
rect 5084 5933 5088 5976
rect 5151 5951 5155 5956
rect 5142 5944 5155 5951
rect 5086 5921 5095 5933
rect 5060 5884 5066 5907
rect 5004 5867 5014 5879
rect 5039 5878 5055 5884
rect 5060 5878 5075 5884
rect 4994 5840 5000 5847
rect 4985 5836 5000 5840
rect 5014 5836 5020 5867
rect 5051 5864 5055 5878
rect 5071 5864 5075 5878
rect 5091 5864 5095 5921
rect 5142 5899 5146 5944
rect 5171 5933 5175 5956
rect 5166 5921 5175 5933
rect 5142 5876 5146 5887
rect 5142 5868 5160 5876
rect 5156 5864 5160 5868
rect 5164 5864 5168 5921
rect 5191 5879 5195 5956
rect 5251 5951 5255 5956
rect 5242 5944 5255 5951
rect 5242 5899 5246 5944
rect 5271 5933 5275 5956
rect 5266 5921 5275 5933
rect 5186 5867 5193 5879
rect 5242 5876 5246 5887
rect 5242 5868 5260 5876
rect 4985 5824 4989 5836
rect 5005 5832 5020 5836
rect 5005 5824 5009 5832
rect 5186 5824 5190 5867
rect 5256 5864 5260 5868
rect 5264 5864 5268 5921
rect 5291 5879 5295 5956
rect 5354 5948 5358 5956
rect 5341 5941 5358 5948
rect 5341 5899 5347 5941
rect 5362 5933 5366 5956
rect 5382 5942 5386 5956
rect 5390 5951 5394 5956
rect 5390 5947 5420 5951
rect 5382 5935 5395 5942
rect 5391 5933 5395 5935
rect 5391 5921 5393 5933
rect 5362 5892 5366 5921
rect 5347 5887 5355 5892
rect 5335 5886 5355 5887
rect 5362 5886 5375 5892
rect 5286 5867 5293 5879
rect 5286 5824 5290 5867
rect 5351 5864 5355 5886
rect 5371 5864 5375 5886
rect 5391 5864 5395 5921
rect 5414 5899 5420 5947
rect 5493 5936 5497 5956
rect 5483 5929 5497 5936
rect 5503 5936 5507 5956
rect 5503 5929 5511 5936
rect 5483 5913 5489 5929
rect 5486 5901 5489 5913
rect 5411 5887 5414 5899
rect 5411 5864 5415 5887
rect 5485 5824 5489 5901
rect 5505 5913 5511 5929
rect 5551 5919 5555 5976
rect 5714 5952 5718 5956
rect 5699 5946 5718 5952
rect 5505 5901 5514 5913
rect 5546 5907 5555 5919
rect 5505 5824 5509 5901
rect 5551 5824 5555 5907
rect 5648 5879 5652 5936
rect 5625 5867 5633 5879
rect 5645 5867 5652 5879
rect 5625 5824 5629 5867
rect 5656 5859 5660 5936
rect 5664 5879 5668 5936
rect 5699 5933 5706 5946
rect 5699 5884 5706 5921
rect 5722 5919 5726 5956
rect 5744 5933 5748 5976
rect 5746 5921 5755 5933
rect 5720 5884 5726 5907
rect 5664 5867 5674 5879
rect 5699 5878 5715 5884
rect 5720 5878 5735 5884
rect 5654 5840 5660 5847
rect 5645 5836 5660 5840
rect 5674 5836 5680 5867
rect 5711 5864 5715 5878
rect 5731 5864 5735 5878
rect 5751 5864 5755 5921
rect 5825 5879 5829 5956
rect 5845 5933 5849 5956
rect 5865 5951 5869 5956
rect 5911 5951 5915 5956
rect 5865 5944 5878 5951
rect 5845 5921 5854 5933
rect 5827 5867 5834 5879
rect 5645 5824 5649 5836
rect 5665 5832 5680 5836
rect 5665 5824 5669 5832
rect 5830 5824 5834 5867
rect 5852 5864 5856 5921
rect 5874 5899 5878 5944
rect 5902 5944 5915 5951
rect 5902 5899 5906 5944
rect 5931 5933 5935 5956
rect 5926 5921 5935 5933
rect 5874 5876 5878 5887
rect 5860 5868 5878 5876
rect 5902 5876 5906 5887
rect 5902 5868 5920 5876
rect 5860 5864 5864 5868
rect 5916 5864 5920 5868
rect 5924 5864 5928 5921
rect 5951 5879 5955 5956
rect 6025 5879 6029 5956
rect 6045 5933 6049 5956
rect 6065 5951 6069 5956
rect 6065 5944 6078 5951
rect 6114 5948 6118 5956
rect 6045 5921 6054 5933
rect 5946 5867 5953 5879
rect 6027 5867 6034 5879
rect 5946 5824 5950 5867
rect 6030 5824 6034 5867
rect 6052 5864 6056 5921
rect 6074 5899 6078 5944
rect 6101 5941 6118 5948
rect 6101 5899 6107 5941
rect 6122 5933 6126 5956
rect 6142 5942 6146 5956
rect 6150 5951 6154 5956
rect 6150 5947 6180 5951
rect 6142 5935 6155 5942
rect 6151 5933 6155 5935
rect 6151 5921 6153 5933
rect 6122 5892 6126 5921
rect 6107 5887 6115 5892
rect 6074 5876 6078 5887
rect 6095 5886 6115 5887
rect 6122 5886 6135 5892
rect 6060 5868 6078 5876
rect 6060 5864 6064 5868
rect 6111 5864 6115 5886
rect 6131 5864 6135 5886
rect 6151 5864 6155 5921
rect 6174 5899 6180 5947
rect 6253 5936 6257 5956
rect 6243 5929 6257 5936
rect 6263 5936 6267 5956
rect 6263 5929 6271 5936
rect 6243 5913 6249 5929
rect 6246 5901 6249 5913
rect 6171 5887 6174 5899
rect 6171 5864 6175 5887
rect 6245 5824 6249 5901
rect 6265 5913 6271 5929
rect 6265 5901 6274 5913
rect 6265 5824 6269 5901
rect 6311 5899 6315 5956
rect 6321 5913 6325 5956
rect 6341 5950 6345 5956
rect 6411 5951 6415 5956
rect 6347 5938 6359 5950
rect 6321 5901 6334 5913
rect 6306 5887 6315 5899
rect 6311 5824 6315 5887
rect 6333 5824 6337 5901
rect 6355 5864 6359 5938
rect 6402 5944 6415 5951
rect 6402 5899 6406 5944
rect 6431 5933 6435 5956
rect 6426 5921 6435 5933
rect 6402 5876 6406 5887
rect 6402 5868 6420 5876
rect 6416 5864 6420 5868
rect 6424 5864 6428 5921
rect 6451 5879 6455 5956
rect 6613 5936 6617 5956
rect 6512 5879 6516 5936
rect 6446 5867 6453 5879
rect 6506 5867 6516 5879
rect 6446 5824 6450 5867
rect 6500 5836 6506 5867
rect 6520 5859 6524 5936
rect 6528 5879 6532 5936
rect 6609 5929 6617 5936
rect 6623 5936 6627 5956
rect 6623 5929 6637 5936
rect 6609 5913 6615 5929
rect 6606 5901 6615 5913
rect 6528 5867 6535 5879
rect 6547 5867 6555 5879
rect 6520 5840 6526 5847
rect 6520 5836 6535 5840
rect 6500 5832 6515 5836
rect 6511 5824 6515 5832
rect 6531 5824 6535 5836
rect 6551 5824 6555 5867
rect 6611 5824 6615 5901
rect 6631 5913 6637 5929
rect 6631 5901 6634 5913
rect 6631 5824 6635 5901
rect 43 5780 47 5784
rect 65 5780 69 5784
rect 111 5780 115 5784
rect 131 5780 135 5784
rect 191 5780 195 5784
rect 211 5780 215 5784
rect 285 5780 289 5784
rect 305 5780 309 5784
rect 325 5780 329 5784
rect 385 5780 389 5784
rect 405 5780 409 5784
rect 451 5780 455 5784
rect 537 5780 541 5784
rect 545 5780 549 5784
rect 591 5780 595 5784
rect 599 5780 603 5784
rect 676 5780 680 5784
rect 684 5780 688 5784
rect 706 5780 710 5784
rect 785 5780 789 5784
rect 831 5780 835 5784
rect 839 5780 843 5784
rect 925 5780 929 5784
rect 945 5780 949 5784
rect 1010 5780 1014 5784
rect 1032 5780 1036 5784
rect 1040 5780 1044 5784
rect 1091 5780 1095 5784
rect 1099 5780 1103 5784
rect 1185 5780 1189 5784
rect 1231 5780 1235 5784
rect 1253 5780 1257 5784
rect 1261 5780 1265 5784
rect 1281 5780 1285 5784
rect 1289 5780 1293 5784
rect 1335 5780 1339 5784
rect 1355 5780 1359 5784
rect 1367 5780 1371 5784
rect 1387 5780 1391 5784
rect 1401 5780 1405 5784
rect 1421 5780 1425 5784
rect 1471 5780 1475 5784
rect 1491 5780 1495 5784
rect 1565 5780 1569 5784
rect 1585 5780 1589 5784
rect 1605 5780 1609 5784
rect 1670 5780 1674 5784
rect 1692 5780 1696 5784
rect 1700 5780 1704 5784
rect 1777 5780 1781 5784
rect 1785 5780 1789 5784
rect 1845 5780 1849 5784
rect 1865 5780 1869 5784
rect 1885 5780 1889 5784
rect 1931 5780 1935 5784
rect 2010 5780 2014 5784
rect 2032 5780 2036 5784
rect 2040 5780 2044 5784
rect 2091 5780 2095 5784
rect 2111 5780 2115 5784
rect 2131 5780 2135 5784
rect 2205 5780 2209 5784
rect 2225 5780 2229 5784
rect 2245 5780 2249 5784
rect 2296 5780 2300 5784
rect 2304 5780 2308 5784
rect 2326 5780 2330 5784
rect 2405 5780 2409 5784
rect 2425 5780 2429 5784
rect 2485 5780 2489 5784
rect 2505 5780 2509 5784
rect 2525 5780 2529 5784
rect 2585 5780 2589 5784
rect 2605 5780 2609 5784
rect 2625 5780 2629 5784
rect 2671 5780 2675 5784
rect 2691 5780 2695 5784
rect 2765 5780 2769 5784
rect 2785 5780 2789 5784
rect 2805 5780 2809 5784
rect 2865 5780 2869 5784
rect 2885 5780 2889 5784
rect 2905 5780 2909 5784
rect 2965 5780 2969 5784
rect 2985 5780 2989 5784
rect 3005 5780 3009 5784
rect 3065 5780 3069 5784
rect 3085 5780 3089 5784
rect 3105 5780 3109 5784
rect 3151 5780 3155 5784
rect 3171 5780 3175 5784
rect 3191 5780 3195 5784
rect 3270 5780 3274 5784
rect 3292 5780 3296 5784
rect 3300 5780 3304 5784
rect 3356 5780 3360 5784
rect 3364 5780 3368 5784
rect 3386 5780 3390 5784
rect 3465 5780 3469 5784
rect 3485 5780 3489 5784
rect 3505 5780 3509 5784
rect 3570 5780 3574 5784
rect 3592 5780 3596 5784
rect 3600 5780 3604 5784
rect 3665 5780 3669 5784
rect 3685 5780 3689 5784
rect 3705 5780 3709 5784
rect 3751 5780 3755 5784
rect 3771 5780 3775 5784
rect 3791 5780 3795 5784
rect 3865 5780 3869 5784
rect 3885 5780 3889 5784
rect 3905 5780 3909 5784
rect 3965 5780 3969 5784
rect 3985 5780 3989 5784
rect 4005 5780 4009 5784
rect 4065 5780 4069 5784
rect 4085 5780 4089 5784
rect 4105 5780 4109 5784
rect 4165 5780 4169 5784
rect 4185 5780 4189 5784
rect 4205 5780 4209 5784
rect 4251 5780 4255 5784
rect 4271 5780 4275 5784
rect 4291 5780 4295 5784
rect 4351 5780 4355 5784
rect 4371 5780 4375 5784
rect 4450 5780 4454 5784
rect 4472 5780 4476 5784
rect 4480 5780 4484 5784
rect 4557 5780 4561 5784
rect 4565 5780 4569 5784
rect 4611 5780 4615 5784
rect 4633 5780 4637 5784
rect 4655 5780 4659 5784
rect 4725 5780 4729 5784
rect 4745 5780 4749 5784
rect 4765 5780 4769 5784
rect 4811 5780 4815 5784
rect 4831 5780 4835 5784
rect 4905 5780 4909 5784
rect 4965 5780 4969 5784
rect 4985 5780 4989 5784
rect 5005 5780 5009 5784
rect 5051 5780 5055 5784
rect 5071 5780 5075 5784
rect 5091 5780 5095 5784
rect 5156 5780 5160 5784
rect 5164 5780 5168 5784
rect 5186 5780 5190 5784
rect 5256 5780 5260 5784
rect 5264 5780 5268 5784
rect 5286 5780 5290 5784
rect 5351 5780 5355 5784
rect 5371 5780 5375 5784
rect 5391 5780 5395 5784
rect 5411 5780 5415 5784
rect 5485 5780 5489 5784
rect 5505 5780 5509 5784
rect 5551 5780 5555 5784
rect 5625 5780 5629 5784
rect 5645 5780 5649 5784
rect 5665 5780 5669 5784
rect 5711 5780 5715 5784
rect 5731 5780 5735 5784
rect 5751 5780 5755 5784
rect 5830 5780 5834 5784
rect 5852 5780 5856 5784
rect 5860 5780 5864 5784
rect 5916 5780 5920 5784
rect 5924 5780 5928 5784
rect 5946 5780 5950 5784
rect 6030 5780 6034 5784
rect 6052 5780 6056 5784
rect 6060 5780 6064 5784
rect 6111 5780 6115 5784
rect 6131 5780 6135 5784
rect 6151 5780 6155 5784
rect 6171 5780 6175 5784
rect 6245 5780 6249 5784
rect 6265 5780 6269 5784
rect 6311 5780 6315 5784
rect 6333 5780 6337 5784
rect 6355 5780 6359 5784
rect 6416 5780 6420 5784
rect 6424 5780 6428 5784
rect 6446 5780 6450 5784
rect 6511 5780 6515 5784
rect 6531 5780 6535 5784
rect 6551 5780 6555 5784
rect 6611 5780 6615 5784
rect 6631 5780 6635 5784
rect 43 5756 47 5760
rect 65 5756 69 5760
rect 123 5756 127 5760
rect 145 5756 149 5760
rect 191 5756 195 5760
rect 213 5756 217 5760
rect 221 5756 225 5760
rect 241 5756 245 5760
rect 249 5756 253 5760
rect 295 5756 299 5760
rect 315 5756 319 5760
rect 327 5756 331 5760
rect 347 5756 351 5760
rect 361 5756 365 5760
rect 381 5756 385 5760
rect 457 5756 461 5760
rect 465 5756 469 5760
rect 511 5756 515 5760
rect 531 5756 535 5760
rect 551 5756 555 5760
rect 611 5756 615 5760
rect 631 5756 635 5760
rect 691 5756 695 5760
rect 713 5756 717 5760
rect 735 5756 739 5760
rect 791 5756 795 5760
rect 811 5756 815 5760
rect 871 5756 875 5760
rect 891 5756 895 5760
rect 951 5756 955 5760
rect 959 5756 963 5760
rect 1031 5756 1035 5760
rect 1091 5756 1095 5760
rect 1101 5756 1105 5760
rect 1121 5756 1125 5760
rect 1191 5756 1195 5760
rect 1199 5756 1203 5760
rect 1271 5756 1275 5760
rect 1331 5756 1335 5760
rect 1339 5756 1343 5760
rect 1411 5756 1415 5760
rect 1471 5756 1475 5760
rect 1493 5756 1497 5760
rect 1501 5756 1505 5760
rect 1521 5756 1525 5760
rect 1529 5756 1533 5760
rect 1575 5756 1579 5760
rect 1595 5756 1599 5760
rect 1607 5756 1611 5760
rect 1627 5756 1631 5760
rect 1641 5756 1645 5760
rect 1661 5756 1665 5760
rect 1711 5756 1715 5760
rect 1721 5756 1725 5760
rect 1751 5756 1755 5760
rect 1761 5756 1765 5760
rect 1850 5756 1854 5760
rect 1872 5756 1876 5760
rect 1880 5756 1884 5760
rect 1945 5756 1949 5760
rect 1965 5756 1969 5760
rect 2011 5756 2015 5760
rect 2085 5756 2089 5760
rect 2105 5756 2109 5760
rect 2125 5756 2129 5760
rect 2171 5756 2175 5760
rect 2179 5756 2183 5760
rect 2251 5756 2255 5760
rect 2271 5756 2275 5760
rect 2405 5756 2409 5760
rect 2425 5756 2429 5760
rect 2445 5756 2449 5760
rect 2465 5756 2469 5760
rect 2525 5756 2529 5760
rect 2545 5756 2549 5760
rect 2605 5756 2609 5760
rect 2625 5756 2629 5760
rect 2645 5756 2649 5760
rect 2705 5756 2709 5760
rect 2725 5756 2729 5760
rect 2745 5756 2749 5760
rect 2791 5756 2795 5760
rect 2811 5756 2815 5760
rect 2876 5756 2880 5760
rect 2884 5756 2888 5760
rect 2906 5756 2910 5760
rect 2985 5756 2989 5760
rect 3005 5756 3009 5760
rect 3025 5756 3029 5760
rect 3071 5756 3075 5760
rect 3091 5756 3095 5760
rect 3111 5756 3115 5760
rect 3190 5756 3194 5760
rect 3212 5756 3216 5760
rect 3220 5756 3224 5760
rect 3285 5756 3289 5760
rect 3331 5756 3335 5760
rect 3351 5756 3355 5760
rect 3371 5756 3375 5760
rect 3445 5756 3449 5760
rect 3465 5756 3469 5760
rect 3485 5756 3489 5760
rect 3545 5756 3549 5760
rect 3565 5756 3569 5760
rect 3585 5756 3589 5760
rect 3645 5756 3649 5760
rect 3710 5756 3714 5760
rect 3732 5756 3736 5760
rect 3740 5756 3744 5760
rect 3817 5756 3821 5760
rect 3825 5756 3829 5760
rect 3876 5756 3880 5760
rect 3884 5756 3888 5760
rect 3906 5756 3910 5760
rect 3985 5756 3989 5760
rect 4045 5756 4049 5760
rect 4065 5756 4069 5760
rect 4085 5756 4089 5760
rect 4105 5756 4109 5760
rect 4170 5756 4174 5760
rect 4192 5756 4196 5760
rect 4200 5756 4204 5760
rect 4265 5756 4269 5760
rect 4285 5756 4289 5760
rect 4305 5756 4309 5760
rect 4351 5756 4355 5760
rect 4430 5756 4434 5760
rect 4452 5756 4456 5760
rect 4460 5756 4464 5760
rect 4521 5756 4525 5760
rect 4543 5756 4547 5760
rect 4565 5756 4569 5760
rect 4611 5756 4615 5760
rect 4631 5756 4635 5760
rect 4710 5756 4714 5760
rect 4732 5756 4736 5760
rect 4740 5756 4744 5760
rect 4796 5756 4800 5760
rect 4804 5756 4808 5760
rect 4826 5756 4830 5760
rect 4905 5756 4909 5760
rect 4925 5756 4929 5760
rect 4945 5756 4949 5760
rect 4991 5756 4995 5760
rect 5011 5756 5015 5760
rect 5031 5756 5035 5760
rect 5096 5756 5100 5760
rect 5104 5756 5108 5760
rect 5126 5756 5130 5760
rect 5191 5756 5195 5760
rect 5211 5756 5215 5760
rect 5231 5756 5235 5760
rect 5291 5756 5295 5760
rect 5311 5756 5315 5760
rect 5371 5756 5375 5760
rect 5391 5756 5395 5760
rect 5411 5756 5415 5760
rect 5471 5756 5475 5760
rect 5491 5756 5495 5760
rect 5511 5756 5515 5760
rect 5571 5756 5575 5760
rect 5591 5756 5595 5760
rect 5665 5756 5669 5760
rect 5685 5756 5689 5760
rect 5731 5756 5735 5760
rect 5751 5756 5755 5760
rect 5771 5756 5775 5760
rect 5791 5756 5795 5760
rect 5870 5756 5874 5760
rect 5892 5756 5896 5760
rect 5900 5756 5904 5760
rect 5951 5756 5955 5760
rect 6011 5756 6015 5760
rect 6031 5756 6035 5760
rect 6051 5756 6055 5760
rect 6071 5756 6075 5760
rect 6131 5756 6135 5760
rect 6151 5756 6155 5760
rect 6171 5756 6175 5760
rect 6245 5756 6249 5760
rect 6291 5756 6295 5760
rect 6311 5756 6315 5760
rect 6331 5756 6335 5760
rect 6391 5756 6395 5760
rect 6411 5756 6415 5760
rect 6431 5756 6435 5760
rect 6491 5756 6495 5760
rect 6511 5756 6515 5760
rect 6531 5756 6535 5760
rect 6591 5756 6595 5760
rect 6611 5756 6615 5760
rect 6631 5756 6635 5760
rect 43 5670 47 5676
rect 43 5658 45 5670
rect 65 5653 69 5716
rect 123 5670 127 5676
rect 123 5658 125 5670
rect 145 5653 149 5716
rect 213 5713 217 5736
rect 209 5706 217 5713
rect 209 5677 213 5706
rect 221 5696 225 5736
rect 241 5684 245 5716
rect 249 5712 253 5716
rect 249 5710 285 5712
rect 249 5708 273 5710
rect 191 5664 195 5676
rect 209 5671 217 5677
rect 65 5641 74 5653
rect 145 5641 154 5653
rect 191 5652 193 5664
rect 43 5590 45 5602
rect 43 5584 47 5590
rect 65 5564 69 5641
rect 123 5590 125 5602
rect 123 5584 127 5590
rect 145 5564 149 5641
rect 191 5584 195 5652
rect 213 5625 217 5671
rect 213 5564 217 5613
rect 241 5589 247 5684
rect 223 5585 247 5589
rect 223 5564 227 5585
rect 243 5580 261 5581
rect 243 5576 273 5580
rect 243 5564 247 5576
rect 281 5572 285 5698
rect 295 5690 299 5716
rect 315 5710 319 5716
rect 251 5568 285 5572
rect 251 5564 255 5568
rect 297 5564 301 5678
rect 313 5588 317 5698
rect 327 5676 331 5716
rect 322 5664 325 5676
rect 322 5600 326 5664
rect 347 5657 351 5716
rect 342 5649 351 5657
rect 342 5620 346 5649
rect 361 5634 365 5716
rect 381 5633 385 5676
rect 457 5653 461 5676
rect 446 5641 461 5653
rect 465 5653 469 5676
rect 511 5662 515 5676
rect 531 5662 535 5676
rect 499 5656 515 5662
rect 520 5656 535 5662
rect 465 5641 474 5653
rect 322 5596 355 5600
rect 321 5576 323 5588
rect 319 5564 323 5576
rect 329 5576 331 5588
rect 329 5564 333 5576
rect 351 5564 355 5596
rect 361 5564 365 5622
rect 381 5584 385 5621
rect 445 5564 449 5641
rect 465 5564 469 5641
rect 499 5619 506 5656
rect 520 5633 526 5656
rect 499 5594 506 5607
rect 499 5588 518 5594
rect 514 5584 518 5588
rect 522 5584 526 5621
rect 551 5619 555 5676
rect 611 5639 615 5716
rect 606 5627 615 5639
rect 546 5607 555 5619
rect 609 5611 615 5627
rect 631 5639 635 5716
rect 691 5653 695 5716
rect 686 5641 695 5653
rect 631 5627 634 5639
rect 631 5611 637 5627
rect 544 5564 548 5607
rect 609 5604 617 5611
rect 613 5584 617 5604
rect 623 5604 637 5611
rect 623 5584 627 5604
rect 691 5584 695 5641
rect 713 5639 717 5716
rect 701 5627 714 5639
rect 701 5584 705 5627
rect 735 5602 739 5676
rect 791 5639 795 5716
rect 786 5627 795 5639
rect 789 5611 795 5627
rect 811 5639 815 5716
rect 871 5639 875 5716
rect 811 5627 814 5639
rect 866 5627 875 5639
rect 811 5611 817 5627
rect 789 5604 797 5611
rect 727 5590 739 5602
rect 721 5584 725 5590
rect 793 5584 797 5604
rect 803 5604 817 5611
rect 869 5611 875 5627
rect 891 5639 895 5716
rect 951 5653 955 5676
rect 946 5641 955 5653
rect 959 5653 963 5676
rect 959 5641 974 5653
rect 891 5627 894 5639
rect 891 5611 897 5627
rect 869 5604 877 5611
rect 803 5584 807 5604
rect 873 5584 877 5604
rect 883 5604 897 5611
rect 883 5584 887 5604
rect 951 5564 955 5641
rect 971 5564 975 5641
rect 1031 5633 1035 5716
rect 1091 5672 1095 5676
rect 1082 5667 1095 5672
rect 1082 5633 1086 5667
rect 1101 5653 1105 5676
rect 1121 5671 1125 5676
rect 1191 5653 1195 5676
rect 1186 5641 1195 5653
rect 1199 5653 1203 5676
rect 1199 5641 1214 5653
rect 1026 5621 1035 5633
rect 1031 5564 1035 5621
rect 1082 5576 1086 5621
rect 1101 5577 1105 5641
rect 1125 5592 1135 5604
rect 1131 5584 1135 5592
rect 1082 5571 1095 5576
rect 1101 5571 1115 5577
rect 1091 5564 1095 5571
rect 1111 5564 1115 5571
rect 1191 5564 1195 5641
rect 1211 5564 1215 5641
rect 1271 5633 1275 5716
rect 1331 5653 1335 5676
rect 1326 5641 1335 5653
rect 1339 5653 1343 5676
rect 1339 5641 1354 5653
rect 1266 5621 1275 5633
rect 1271 5564 1275 5621
rect 1331 5564 1335 5641
rect 1351 5564 1355 5641
rect 1411 5633 1415 5716
rect 1493 5713 1497 5736
rect 1489 5706 1497 5713
rect 1489 5677 1493 5706
rect 1501 5696 1505 5736
rect 1521 5684 1525 5716
rect 1529 5712 1533 5716
rect 1529 5710 1565 5712
rect 1529 5708 1553 5710
rect 1406 5621 1415 5633
rect 1411 5564 1415 5621
rect 1471 5664 1475 5676
rect 1489 5671 1497 5677
rect 1471 5652 1473 5664
rect 1471 5584 1475 5652
rect 1493 5625 1497 5671
rect 1493 5564 1497 5613
rect 1521 5589 1527 5684
rect 1503 5585 1527 5589
rect 1503 5564 1507 5585
rect 1523 5580 1541 5581
rect 1523 5576 1553 5580
rect 1523 5564 1527 5576
rect 1561 5572 1565 5698
rect 1575 5690 1579 5716
rect 1595 5710 1599 5716
rect 1531 5568 1565 5572
rect 1531 5564 1535 5568
rect 1577 5564 1581 5678
rect 1593 5588 1597 5698
rect 1607 5676 1611 5716
rect 1602 5664 1605 5676
rect 1602 5600 1606 5664
rect 1627 5657 1631 5716
rect 1622 5649 1631 5657
rect 1622 5620 1626 5649
rect 1641 5634 1645 5716
rect 1661 5633 1665 5676
rect 1711 5672 1715 5676
rect 1701 5668 1715 5672
rect 1721 5672 1725 5676
rect 1721 5668 1735 5672
rect 1701 5653 1706 5668
rect 1602 5596 1635 5600
rect 1601 5576 1603 5588
rect 1599 5564 1603 5576
rect 1609 5576 1611 5588
rect 1609 5564 1613 5576
rect 1631 5564 1635 5596
rect 1641 5564 1645 5622
rect 1661 5584 1665 5621
rect 1700 5595 1706 5641
rect 1729 5619 1735 5668
rect 1751 5619 1755 5676
rect 1761 5672 1765 5676
rect 1850 5673 1854 5716
rect 1761 5668 1775 5672
rect 1771 5653 1775 5668
rect 1847 5661 1854 5673
rect 1771 5641 1773 5653
rect 1726 5607 1735 5619
rect 1700 5591 1715 5595
rect 1711 5584 1715 5591
rect 1731 5584 1735 5607
rect 1751 5584 1755 5607
rect 1771 5584 1775 5641
rect 1845 5584 1849 5661
rect 1872 5619 1876 5676
rect 1880 5672 1884 5676
rect 1880 5664 1898 5672
rect 1894 5653 1898 5664
rect 1865 5607 1874 5619
rect 1865 5584 1869 5607
rect 1894 5596 1898 5641
rect 1945 5639 1949 5716
rect 1946 5627 1949 5639
rect 1943 5611 1949 5627
rect 1965 5639 1969 5716
rect 1965 5627 1974 5639
rect 2011 5633 2015 5716
rect 2341 5748 2345 5752
rect 2361 5748 2365 5752
rect 1965 5611 1971 5627
rect 2006 5621 2015 5633
rect 1943 5604 1957 5611
rect 1885 5589 1898 5596
rect 1885 5584 1889 5589
rect 1953 5584 1957 5604
rect 1963 5604 1971 5611
rect 1963 5584 1967 5604
rect 2011 5564 2015 5621
rect 2085 5619 2089 5676
rect 2105 5662 2109 5676
rect 2125 5662 2129 5676
rect 2105 5656 2120 5662
rect 2125 5656 2141 5662
rect 2114 5633 2120 5656
rect 2085 5607 2094 5619
rect 2092 5564 2096 5607
rect 2114 5584 2118 5621
rect 2134 5619 2141 5656
rect 2171 5653 2175 5676
rect 2166 5641 2175 5653
rect 2179 5653 2183 5676
rect 2179 5641 2194 5653
rect 2134 5594 2141 5607
rect 2122 5588 2141 5594
rect 2122 5584 2126 5588
rect 2171 5564 2175 5641
rect 2191 5564 2195 5641
rect 2251 5639 2255 5716
rect 2246 5627 2255 5639
rect 2249 5611 2255 5627
rect 2271 5639 2275 5716
rect 2405 5692 2409 5696
rect 2425 5692 2429 5696
rect 2405 5688 2429 5692
rect 2341 5680 2345 5688
rect 2361 5680 2365 5688
rect 2341 5676 2391 5680
rect 2385 5653 2391 5676
rect 2385 5641 2394 5653
rect 2271 5627 2274 5639
rect 2271 5611 2277 5627
rect 2249 5604 2257 5611
rect 2253 5584 2257 5604
rect 2263 5604 2277 5611
rect 2263 5584 2267 5604
rect 2385 5586 2391 5641
rect 2425 5619 2429 5688
rect 2426 5607 2429 5619
rect 2385 5580 2409 5586
rect 2405 5564 2409 5580
rect 2425 5564 2429 5607
rect 2445 5692 2449 5696
rect 2465 5692 2469 5696
rect 2445 5688 2469 5692
rect 2445 5653 2449 5688
rect 2445 5641 2454 5653
rect 2445 5564 2449 5641
rect 2525 5639 2529 5716
rect 2526 5627 2529 5639
rect 2523 5611 2529 5627
rect 2545 5639 2549 5716
rect 2605 5673 2609 5716
rect 2625 5704 2629 5716
rect 2645 5708 2649 5716
rect 2645 5704 2660 5708
rect 2625 5700 2640 5704
rect 2634 5693 2640 5700
rect 2605 5661 2613 5673
rect 2625 5661 2632 5673
rect 2545 5627 2554 5639
rect 2545 5611 2551 5627
rect 2523 5604 2537 5611
rect 2533 5584 2537 5604
rect 2543 5604 2551 5611
rect 2628 5604 2632 5661
rect 2636 5604 2640 5681
rect 2654 5673 2660 5704
rect 2705 5673 2709 5716
rect 2725 5704 2729 5716
rect 2745 5708 2749 5716
rect 2745 5704 2760 5708
rect 2725 5700 2740 5704
rect 2734 5693 2740 5700
rect 2644 5661 2654 5673
rect 2705 5661 2713 5673
rect 2725 5661 2732 5673
rect 2644 5604 2648 5661
rect 2728 5604 2732 5661
rect 2736 5604 2740 5681
rect 2754 5673 2760 5704
rect 2744 5661 2754 5673
rect 2744 5604 2748 5661
rect 2791 5639 2795 5716
rect 2786 5627 2795 5639
rect 2789 5611 2795 5627
rect 2811 5639 2815 5716
rect 2876 5672 2880 5676
rect 2862 5664 2880 5672
rect 2862 5653 2866 5664
rect 2811 5627 2814 5639
rect 2811 5611 2817 5627
rect 2789 5604 2797 5611
rect 2543 5584 2547 5604
rect 2793 5584 2797 5604
rect 2803 5604 2817 5611
rect 2803 5584 2807 5604
rect 2862 5596 2866 5641
rect 2884 5619 2888 5676
rect 2906 5673 2910 5716
rect 2985 5673 2989 5716
rect 3005 5704 3009 5716
rect 3025 5708 3029 5716
rect 3025 5704 3040 5708
rect 3005 5700 3020 5704
rect 3014 5693 3020 5700
rect 2906 5661 2913 5673
rect 2985 5661 2993 5673
rect 3005 5661 3012 5673
rect 2886 5607 2895 5619
rect 2862 5589 2875 5596
rect 2871 5584 2875 5589
rect 2891 5584 2895 5607
rect 2911 5584 2915 5661
rect 3008 5604 3012 5661
rect 3016 5604 3020 5681
rect 3034 5673 3040 5704
rect 3024 5661 3034 5673
rect 3071 5662 3075 5676
rect 3091 5662 3095 5676
rect 3024 5604 3028 5661
rect 3059 5656 3075 5662
rect 3080 5656 3095 5662
rect 3059 5619 3066 5656
rect 3080 5633 3086 5656
rect 3059 5594 3066 5607
rect 3059 5588 3078 5594
rect 3074 5584 3078 5588
rect 3082 5584 3086 5621
rect 3111 5619 3115 5676
rect 3190 5673 3194 5716
rect 3187 5661 3194 5673
rect 3106 5607 3115 5619
rect 3104 5564 3108 5607
rect 3185 5584 3189 5661
rect 3212 5619 3216 5676
rect 3220 5672 3224 5676
rect 3220 5664 3238 5672
rect 3234 5653 3238 5664
rect 3205 5607 3214 5619
rect 3205 5584 3209 5607
rect 3234 5596 3238 5641
rect 3225 5589 3238 5596
rect 3285 5633 3289 5716
rect 3331 5708 3335 5716
rect 3320 5704 3335 5708
rect 3351 5704 3355 5716
rect 3320 5673 3326 5704
rect 3340 5700 3355 5704
rect 3340 5693 3346 5700
rect 3326 5661 3336 5673
rect 3285 5621 3294 5633
rect 3225 5584 3229 5589
rect 3285 5564 3289 5621
rect 3332 5604 3336 5661
rect 3340 5604 3344 5681
rect 3371 5673 3375 5716
rect 3348 5661 3355 5673
rect 3367 5661 3375 5673
rect 3445 5673 3449 5716
rect 3465 5704 3469 5716
rect 3485 5708 3489 5716
rect 3485 5704 3500 5708
rect 3465 5700 3480 5704
rect 3474 5693 3480 5700
rect 3445 5661 3453 5673
rect 3465 5661 3472 5673
rect 3348 5604 3352 5661
rect 3468 5604 3472 5661
rect 3476 5604 3480 5681
rect 3494 5673 3500 5704
rect 3545 5673 3549 5716
rect 3565 5704 3569 5716
rect 3585 5708 3589 5716
rect 3585 5704 3600 5708
rect 3565 5700 3580 5704
rect 3574 5693 3580 5700
rect 3484 5661 3494 5673
rect 3545 5661 3553 5673
rect 3565 5661 3572 5673
rect 3484 5604 3488 5661
rect 3568 5604 3572 5661
rect 3576 5604 3580 5681
rect 3594 5673 3600 5704
rect 3584 5661 3594 5673
rect 3584 5604 3588 5661
rect 3645 5633 3649 5716
rect 3710 5673 3714 5716
rect 3707 5661 3714 5673
rect 3645 5621 3654 5633
rect 3645 5564 3649 5621
rect 3705 5584 3709 5661
rect 3732 5619 3736 5676
rect 3740 5672 3744 5676
rect 3740 5664 3758 5672
rect 3754 5653 3758 5664
rect 3817 5653 3821 5676
rect 3806 5641 3821 5653
rect 3825 5653 3829 5676
rect 3876 5672 3880 5676
rect 3862 5664 3880 5672
rect 3862 5653 3866 5664
rect 3825 5641 3834 5653
rect 3725 5607 3734 5619
rect 3725 5584 3729 5607
rect 3754 5596 3758 5641
rect 3745 5589 3758 5596
rect 3745 5584 3749 5589
rect 3805 5564 3809 5641
rect 3825 5564 3829 5641
rect 3862 5596 3866 5641
rect 3884 5619 3888 5676
rect 3906 5673 3910 5716
rect 3906 5661 3913 5673
rect 3886 5607 3895 5619
rect 3862 5589 3875 5596
rect 3871 5584 3875 5589
rect 3891 5584 3895 5607
rect 3911 5584 3915 5661
rect 3985 5633 3989 5716
rect 4045 5653 4049 5676
rect 4046 5641 4049 5653
rect 3985 5621 3994 5633
rect 3985 5564 3989 5621
rect 4040 5593 4046 5641
rect 4065 5619 4069 5676
rect 4085 5654 4089 5676
rect 4105 5654 4109 5676
rect 4170 5673 4174 5716
rect 4167 5661 4174 5673
rect 4085 5648 4098 5654
rect 4105 5653 4125 5654
rect 4105 5648 4113 5653
rect 4094 5619 4098 5648
rect 4067 5607 4069 5619
rect 4065 5605 4069 5607
rect 4065 5598 4078 5605
rect 4040 5589 4070 5593
rect 4066 5584 4070 5589
rect 4074 5584 4078 5598
rect 4094 5584 4098 5607
rect 4113 5599 4119 5641
rect 4102 5592 4119 5599
rect 4102 5584 4106 5592
rect 4165 5584 4169 5661
rect 4192 5619 4196 5676
rect 4200 5672 4204 5676
rect 4265 5673 4269 5716
rect 4285 5704 4289 5716
rect 4305 5708 4309 5716
rect 4305 5704 4320 5708
rect 4285 5700 4300 5704
rect 4294 5693 4300 5700
rect 4200 5664 4218 5672
rect 4214 5653 4218 5664
rect 4265 5661 4273 5673
rect 4285 5661 4292 5673
rect 4185 5607 4194 5619
rect 4185 5584 4189 5607
rect 4214 5596 4218 5641
rect 4288 5604 4292 5661
rect 4296 5604 4300 5681
rect 4314 5673 4320 5704
rect 4304 5661 4314 5673
rect 4304 5604 4308 5661
rect 4351 5633 4355 5716
rect 4430 5673 4434 5716
rect 4427 5661 4434 5673
rect 4346 5621 4355 5633
rect 4205 5589 4218 5596
rect 4205 5584 4209 5589
rect 4351 5564 4355 5621
rect 4425 5584 4429 5661
rect 4452 5619 4456 5676
rect 4460 5672 4464 5676
rect 4460 5664 4478 5672
rect 4474 5653 4478 5664
rect 4445 5607 4454 5619
rect 4445 5584 4449 5607
rect 4474 5596 4478 5641
rect 4465 5589 4478 5596
rect 4521 5602 4525 5676
rect 4543 5639 4547 5716
rect 4565 5653 4569 5716
rect 4565 5641 4574 5653
rect 4546 5627 4559 5639
rect 4521 5590 4533 5602
rect 4465 5584 4469 5589
rect 4535 5584 4539 5590
rect 4555 5584 4559 5627
rect 4565 5584 4569 5641
rect 4611 5639 4615 5716
rect 4606 5627 4615 5639
rect 4609 5611 4615 5627
rect 4631 5639 4635 5716
rect 4710 5673 4714 5716
rect 4707 5661 4714 5673
rect 4631 5627 4634 5639
rect 4631 5611 4637 5627
rect 4609 5604 4617 5611
rect 4613 5584 4617 5604
rect 4623 5604 4637 5611
rect 4623 5584 4627 5604
rect 4705 5584 4709 5661
rect 4732 5619 4736 5676
rect 4740 5672 4744 5676
rect 4796 5672 4800 5676
rect 4740 5664 4758 5672
rect 4754 5653 4758 5664
rect 4782 5664 4800 5672
rect 4782 5653 4786 5664
rect 4725 5607 4734 5619
rect 4725 5584 4729 5607
rect 4754 5596 4758 5641
rect 4745 5589 4758 5596
rect 4782 5596 4786 5641
rect 4804 5619 4808 5676
rect 4826 5673 4830 5716
rect 4905 5673 4909 5716
rect 4925 5704 4929 5716
rect 4945 5708 4949 5716
rect 4945 5704 4960 5708
rect 4925 5700 4940 5704
rect 4934 5693 4940 5700
rect 4826 5661 4833 5673
rect 4905 5661 4913 5673
rect 4925 5661 4932 5673
rect 4806 5607 4815 5619
rect 4782 5589 4795 5596
rect 4745 5584 4749 5589
rect 4791 5584 4795 5589
rect 4811 5584 4815 5607
rect 4831 5584 4835 5661
rect 4928 5604 4932 5661
rect 4936 5604 4940 5681
rect 4954 5673 4960 5704
rect 4944 5661 4954 5673
rect 4991 5662 4995 5676
rect 5011 5662 5015 5676
rect 4944 5604 4948 5661
rect 4979 5656 4995 5662
rect 5000 5656 5015 5662
rect 4979 5619 4986 5656
rect 5000 5633 5006 5656
rect 4979 5594 4986 5607
rect 4979 5588 4998 5594
rect 4994 5584 4998 5588
rect 5002 5584 5006 5621
rect 5031 5619 5035 5676
rect 5096 5672 5100 5676
rect 5082 5664 5100 5672
rect 5082 5653 5086 5664
rect 5026 5607 5035 5619
rect 5024 5564 5028 5607
rect 5082 5596 5086 5641
rect 5104 5619 5108 5676
rect 5126 5673 5130 5716
rect 5191 5708 5195 5716
rect 5180 5704 5195 5708
rect 5211 5704 5215 5716
rect 5180 5673 5186 5704
rect 5200 5700 5215 5704
rect 5200 5693 5206 5700
rect 5126 5661 5133 5673
rect 5186 5661 5196 5673
rect 5106 5607 5115 5619
rect 5082 5589 5095 5596
rect 5091 5584 5095 5589
rect 5111 5584 5115 5607
rect 5131 5584 5135 5661
rect 5192 5604 5196 5661
rect 5200 5604 5204 5681
rect 5231 5673 5235 5716
rect 5208 5661 5215 5673
rect 5227 5661 5235 5673
rect 5208 5604 5212 5661
rect 5291 5639 5295 5716
rect 5286 5627 5295 5639
rect 5289 5611 5295 5627
rect 5311 5639 5315 5716
rect 5371 5708 5375 5716
rect 5360 5704 5375 5708
rect 5391 5704 5395 5716
rect 5360 5673 5366 5704
rect 5380 5700 5395 5704
rect 5380 5693 5386 5700
rect 5366 5661 5376 5673
rect 5311 5627 5314 5639
rect 5311 5611 5317 5627
rect 5289 5604 5297 5611
rect 5293 5584 5297 5604
rect 5303 5604 5317 5611
rect 5372 5604 5376 5661
rect 5380 5604 5384 5681
rect 5411 5673 5415 5716
rect 5388 5661 5395 5673
rect 5407 5661 5415 5673
rect 5471 5662 5475 5676
rect 5491 5662 5495 5676
rect 5388 5604 5392 5661
rect 5459 5656 5475 5662
rect 5480 5656 5495 5662
rect 5459 5619 5466 5656
rect 5480 5633 5486 5656
rect 5303 5584 5307 5604
rect 5459 5594 5466 5607
rect 5459 5588 5478 5594
rect 5474 5584 5478 5588
rect 5482 5584 5486 5621
rect 5511 5619 5515 5676
rect 5571 5639 5575 5716
rect 5566 5627 5575 5639
rect 5506 5607 5515 5619
rect 5569 5611 5575 5627
rect 5591 5639 5595 5716
rect 5665 5639 5669 5716
rect 5591 5627 5594 5639
rect 5666 5627 5669 5639
rect 5591 5611 5597 5627
rect 5504 5564 5508 5607
rect 5569 5604 5577 5611
rect 5573 5584 5577 5604
rect 5583 5604 5597 5611
rect 5663 5611 5669 5627
rect 5685 5639 5689 5716
rect 5731 5654 5735 5676
rect 5751 5654 5755 5676
rect 5715 5653 5735 5654
rect 5727 5648 5735 5653
rect 5742 5648 5755 5654
rect 5685 5627 5694 5639
rect 5685 5611 5691 5627
rect 5663 5604 5677 5611
rect 5583 5584 5587 5604
rect 5673 5584 5677 5604
rect 5683 5604 5691 5611
rect 5683 5584 5687 5604
rect 5721 5599 5727 5641
rect 5742 5619 5746 5648
rect 5771 5619 5775 5676
rect 5791 5653 5795 5676
rect 5870 5673 5874 5716
rect 5867 5661 5874 5673
rect 5791 5641 5794 5653
rect 5771 5607 5773 5619
rect 5721 5592 5738 5599
rect 5734 5584 5738 5592
rect 5742 5584 5746 5607
rect 5771 5605 5775 5607
rect 5762 5598 5775 5605
rect 5762 5584 5766 5598
rect 5794 5593 5800 5641
rect 5770 5589 5800 5593
rect 5770 5584 5774 5589
rect 5865 5584 5869 5661
rect 5892 5619 5896 5676
rect 5900 5672 5904 5676
rect 5900 5664 5918 5672
rect 5914 5653 5918 5664
rect 5885 5607 5894 5619
rect 5885 5584 5889 5607
rect 5914 5596 5918 5641
rect 5951 5633 5955 5716
rect 6131 5708 6135 5716
rect 6120 5704 6135 5708
rect 6151 5704 6155 5716
rect 6011 5654 6015 5676
rect 6031 5654 6035 5676
rect 5995 5653 6015 5654
rect 6007 5648 6015 5653
rect 6022 5648 6035 5654
rect 5946 5621 5955 5633
rect 5905 5589 5918 5596
rect 5905 5584 5909 5589
rect 5951 5564 5955 5621
rect 6001 5599 6007 5641
rect 6022 5619 6026 5648
rect 6051 5619 6055 5676
rect 6071 5653 6075 5676
rect 6120 5673 6126 5704
rect 6140 5700 6155 5704
rect 6140 5693 6146 5700
rect 6126 5661 6136 5673
rect 6071 5641 6074 5653
rect 6051 5607 6053 5619
rect 6001 5592 6018 5599
rect 6014 5584 6018 5592
rect 6022 5584 6026 5607
rect 6051 5605 6055 5607
rect 6042 5598 6055 5605
rect 6042 5584 6046 5598
rect 6074 5593 6080 5641
rect 6132 5604 6136 5661
rect 6140 5604 6144 5681
rect 6171 5673 6175 5716
rect 6148 5661 6155 5673
rect 6167 5661 6175 5673
rect 6148 5604 6152 5661
rect 6245 5633 6249 5716
rect 6391 5708 6395 5716
rect 6380 5704 6395 5708
rect 6411 5704 6415 5716
rect 6291 5662 6295 5676
rect 6311 5662 6315 5676
rect 6279 5656 6295 5662
rect 6300 5656 6315 5662
rect 6245 5621 6254 5633
rect 6050 5589 6080 5593
rect 6050 5584 6054 5589
rect 6245 5564 6249 5621
rect 6279 5619 6286 5656
rect 6300 5633 6306 5656
rect 6279 5594 6286 5607
rect 6279 5588 6298 5594
rect 6294 5584 6298 5588
rect 6302 5584 6306 5621
rect 6331 5619 6335 5676
rect 6380 5673 6386 5704
rect 6400 5700 6415 5704
rect 6400 5693 6406 5700
rect 6386 5661 6396 5673
rect 6326 5607 6335 5619
rect 6324 5564 6328 5607
rect 6392 5604 6396 5661
rect 6400 5604 6404 5681
rect 6431 5673 6435 5716
rect 6491 5708 6495 5716
rect 6480 5704 6495 5708
rect 6511 5704 6515 5716
rect 6480 5673 6486 5704
rect 6500 5700 6515 5704
rect 6500 5693 6506 5700
rect 6408 5661 6415 5673
rect 6427 5661 6435 5673
rect 6486 5661 6496 5673
rect 6408 5604 6412 5661
rect 6492 5604 6496 5661
rect 6500 5604 6504 5681
rect 6531 5673 6535 5716
rect 6591 5708 6595 5716
rect 6580 5704 6595 5708
rect 6611 5704 6615 5716
rect 6580 5673 6586 5704
rect 6600 5700 6615 5704
rect 6600 5693 6606 5700
rect 6508 5661 6515 5673
rect 6527 5661 6535 5673
rect 6586 5661 6596 5673
rect 6508 5604 6512 5661
rect 6592 5604 6596 5661
rect 6600 5604 6604 5681
rect 6631 5673 6635 5716
rect 6608 5661 6615 5673
rect 6627 5661 6635 5673
rect 6608 5604 6612 5661
rect 43 5540 47 5544
rect 65 5540 69 5544
rect 123 5540 127 5544
rect 145 5540 149 5544
rect 191 5540 195 5544
rect 213 5540 217 5544
rect 223 5540 227 5544
rect 243 5540 247 5544
rect 251 5540 255 5544
rect 297 5540 301 5544
rect 319 5540 323 5544
rect 329 5540 333 5544
rect 351 5540 355 5544
rect 361 5540 365 5544
rect 381 5540 385 5544
rect 445 5540 449 5544
rect 465 5540 469 5544
rect 514 5540 518 5544
rect 522 5540 526 5544
rect 544 5540 548 5544
rect 613 5540 617 5544
rect 623 5540 627 5544
rect 691 5540 695 5544
rect 701 5540 705 5544
rect 721 5540 725 5544
rect 793 5540 797 5544
rect 803 5540 807 5544
rect 873 5540 877 5544
rect 883 5540 887 5544
rect 951 5540 955 5544
rect 971 5540 975 5544
rect 1031 5540 1035 5544
rect 1091 5540 1095 5544
rect 1111 5540 1115 5544
rect 1131 5540 1135 5544
rect 1191 5540 1195 5544
rect 1211 5540 1215 5544
rect 1271 5540 1275 5544
rect 1331 5540 1335 5544
rect 1351 5540 1355 5544
rect 1411 5540 1415 5544
rect 1471 5540 1475 5544
rect 1493 5540 1497 5544
rect 1503 5540 1507 5544
rect 1523 5540 1527 5544
rect 1531 5540 1535 5544
rect 1577 5540 1581 5544
rect 1599 5540 1603 5544
rect 1609 5540 1613 5544
rect 1631 5540 1635 5544
rect 1641 5540 1645 5544
rect 1661 5540 1665 5544
rect 1711 5540 1715 5544
rect 1731 5540 1735 5544
rect 1751 5540 1755 5544
rect 1771 5540 1775 5544
rect 1845 5540 1849 5544
rect 1865 5540 1869 5544
rect 1885 5540 1889 5544
rect 1953 5540 1957 5544
rect 1963 5540 1967 5544
rect 2011 5540 2015 5544
rect 2092 5540 2096 5544
rect 2114 5540 2118 5544
rect 2122 5540 2126 5544
rect 2171 5540 2175 5544
rect 2191 5540 2195 5544
rect 2253 5540 2257 5544
rect 2263 5540 2267 5544
rect 2405 5540 2409 5544
rect 2425 5540 2429 5544
rect 2445 5540 2449 5544
rect 2533 5540 2537 5544
rect 2543 5540 2547 5544
rect 2628 5540 2632 5544
rect 2636 5540 2640 5544
rect 2644 5540 2648 5544
rect 2728 5540 2732 5544
rect 2736 5540 2740 5544
rect 2744 5540 2748 5544
rect 2793 5540 2797 5544
rect 2803 5540 2807 5544
rect 2871 5540 2875 5544
rect 2891 5540 2895 5544
rect 2911 5540 2915 5544
rect 3008 5540 3012 5544
rect 3016 5540 3020 5544
rect 3024 5540 3028 5544
rect 3074 5540 3078 5544
rect 3082 5540 3086 5544
rect 3104 5540 3108 5544
rect 3185 5540 3189 5544
rect 3205 5540 3209 5544
rect 3225 5540 3229 5544
rect 3285 5540 3289 5544
rect 3332 5540 3336 5544
rect 3340 5540 3344 5544
rect 3348 5540 3352 5544
rect 3468 5540 3472 5544
rect 3476 5540 3480 5544
rect 3484 5540 3488 5544
rect 3568 5540 3572 5544
rect 3576 5540 3580 5544
rect 3584 5540 3588 5544
rect 3645 5540 3649 5544
rect 3705 5540 3709 5544
rect 3725 5540 3729 5544
rect 3745 5540 3749 5544
rect 3805 5540 3809 5544
rect 3825 5540 3829 5544
rect 3871 5540 3875 5544
rect 3891 5540 3895 5544
rect 3911 5540 3915 5544
rect 3985 5540 3989 5544
rect 4066 5540 4070 5544
rect 4074 5540 4078 5544
rect 4094 5540 4098 5544
rect 4102 5540 4106 5544
rect 4165 5540 4169 5544
rect 4185 5540 4189 5544
rect 4205 5540 4209 5544
rect 4288 5540 4292 5544
rect 4296 5540 4300 5544
rect 4304 5540 4308 5544
rect 4351 5540 4355 5544
rect 4425 5540 4429 5544
rect 4445 5540 4449 5544
rect 4465 5540 4469 5544
rect 4535 5540 4539 5544
rect 4555 5540 4559 5544
rect 4565 5540 4569 5544
rect 4613 5540 4617 5544
rect 4623 5540 4627 5544
rect 4705 5540 4709 5544
rect 4725 5540 4729 5544
rect 4745 5540 4749 5544
rect 4791 5540 4795 5544
rect 4811 5540 4815 5544
rect 4831 5540 4835 5544
rect 4928 5540 4932 5544
rect 4936 5540 4940 5544
rect 4944 5540 4948 5544
rect 4994 5540 4998 5544
rect 5002 5540 5006 5544
rect 5024 5540 5028 5544
rect 5091 5540 5095 5544
rect 5111 5540 5115 5544
rect 5131 5540 5135 5544
rect 5192 5540 5196 5544
rect 5200 5540 5204 5544
rect 5208 5540 5212 5544
rect 5293 5540 5297 5544
rect 5303 5540 5307 5544
rect 5372 5540 5376 5544
rect 5380 5540 5384 5544
rect 5388 5540 5392 5544
rect 5474 5540 5478 5544
rect 5482 5540 5486 5544
rect 5504 5540 5508 5544
rect 5573 5540 5577 5544
rect 5583 5540 5587 5544
rect 5673 5540 5677 5544
rect 5683 5540 5687 5544
rect 5734 5540 5738 5544
rect 5742 5540 5746 5544
rect 5762 5540 5766 5544
rect 5770 5540 5774 5544
rect 5865 5540 5869 5544
rect 5885 5540 5889 5544
rect 5905 5540 5909 5544
rect 5951 5540 5955 5544
rect 6014 5540 6018 5544
rect 6022 5540 6026 5544
rect 6042 5540 6046 5544
rect 6050 5540 6054 5544
rect 6132 5540 6136 5544
rect 6140 5540 6144 5544
rect 6148 5540 6152 5544
rect 6245 5540 6249 5544
rect 6294 5540 6298 5544
rect 6302 5540 6306 5544
rect 6324 5540 6328 5544
rect 6392 5540 6396 5544
rect 6400 5540 6404 5544
rect 6408 5540 6412 5544
rect 6492 5540 6496 5544
rect 6500 5540 6504 5544
rect 6508 5540 6512 5544
rect 6592 5540 6596 5544
rect 6600 5540 6604 5544
rect 6608 5540 6612 5544
rect 31 5516 35 5520
rect 53 5516 57 5520
rect 63 5516 67 5520
rect 83 5516 87 5520
rect 91 5516 95 5520
rect 137 5516 141 5520
rect 159 5516 163 5520
rect 169 5516 173 5520
rect 191 5516 195 5520
rect 201 5516 205 5520
rect 221 5516 225 5520
rect 273 5516 277 5520
rect 283 5516 287 5520
rect 372 5516 376 5520
rect 394 5516 398 5520
rect 402 5516 406 5520
rect 473 5516 477 5520
rect 483 5516 487 5520
rect 555 5516 559 5520
rect 575 5516 579 5520
rect 585 5516 589 5520
rect 631 5516 635 5520
rect 651 5516 655 5520
rect 711 5516 715 5520
rect 731 5516 735 5520
rect 793 5516 797 5520
rect 803 5516 807 5520
rect 873 5516 877 5520
rect 883 5516 887 5520
rect 951 5516 955 5520
rect 1014 5516 1018 5520
rect 1022 5516 1026 5520
rect 1044 5516 1048 5520
rect 1146 5516 1150 5520
rect 1154 5516 1158 5520
rect 1174 5516 1178 5520
rect 1182 5516 1186 5520
rect 1231 5516 1235 5520
rect 1253 5516 1257 5520
rect 1263 5516 1267 5520
rect 1283 5516 1287 5520
rect 1291 5516 1295 5520
rect 1337 5516 1341 5520
rect 1359 5516 1363 5520
rect 1369 5516 1373 5520
rect 1391 5516 1395 5520
rect 1401 5516 1405 5520
rect 1421 5516 1425 5520
rect 1508 5516 1512 5520
rect 1516 5516 1520 5520
rect 1524 5516 1528 5520
rect 1608 5516 1612 5520
rect 1616 5516 1620 5520
rect 1624 5516 1628 5520
rect 1685 5516 1689 5520
rect 1745 5516 1749 5520
rect 1765 5516 1769 5520
rect 1785 5516 1789 5520
rect 1855 5516 1859 5520
rect 1875 5516 1879 5520
rect 1885 5516 1889 5520
rect 1953 5516 1957 5520
rect 1963 5516 1967 5520
rect 2025 5516 2029 5520
rect 2045 5516 2049 5520
rect 2065 5516 2069 5520
rect 2113 5516 2117 5520
rect 2123 5516 2127 5520
rect 2205 5516 2209 5520
rect 2265 5516 2269 5520
rect 2285 5516 2289 5520
rect 2305 5516 2309 5520
rect 2351 5516 2355 5520
rect 2371 5516 2375 5520
rect 2445 5516 2449 5520
rect 2512 5516 2516 5520
rect 2534 5516 2538 5520
rect 2542 5516 2546 5520
rect 2591 5516 2595 5520
rect 2611 5516 2615 5520
rect 2631 5516 2635 5520
rect 2693 5516 2697 5520
rect 2703 5516 2707 5520
rect 2808 5516 2812 5520
rect 2816 5516 2820 5520
rect 2824 5516 2828 5520
rect 2893 5516 2897 5520
rect 2903 5516 2907 5520
rect 2965 5516 2969 5520
rect 2985 5516 2989 5520
rect 3031 5516 3035 5520
rect 3051 5516 3055 5520
rect 3071 5516 3075 5520
rect 3153 5516 3157 5520
rect 3163 5516 3167 5520
rect 3211 5516 3215 5520
rect 3231 5516 3235 5520
rect 3251 5516 3255 5520
rect 3335 5516 3339 5520
rect 3355 5516 3359 5520
rect 3365 5516 3369 5520
rect 3411 5516 3415 5520
rect 3431 5516 3435 5520
rect 3491 5516 3495 5520
rect 3511 5516 3515 5520
rect 3531 5516 3535 5520
rect 3591 5516 3595 5520
rect 3611 5516 3615 5520
rect 3631 5516 3635 5520
rect 3705 5516 3709 5520
rect 3725 5516 3729 5520
rect 3771 5516 3775 5520
rect 3791 5516 3795 5520
rect 3811 5516 3815 5520
rect 3831 5516 3835 5520
rect 3905 5516 3909 5520
rect 3925 5516 3929 5520
rect 3971 5516 3975 5520
rect 3991 5516 3995 5520
rect 4011 5516 4015 5520
rect 4108 5516 4112 5520
rect 4116 5516 4120 5520
rect 4124 5516 4128 5520
rect 4193 5516 4197 5520
rect 4203 5516 4207 5520
rect 4251 5516 4255 5520
rect 4325 5516 4329 5520
rect 4345 5516 4349 5520
rect 4365 5516 4369 5520
rect 4433 5516 4437 5520
rect 4443 5516 4447 5520
rect 4493 5516 4497 5520
rect 4503 5516 4507 5520
rect 4585 5516 4589 5520
rect 4605 5516 4609 5520
rect 4625 5516 4629 5520
rect 4685 5516 4689 5520
rect 4705 5516 4709 5520
rect 4725 5516 4729 5520
rect 4795 5516 4799 5520
rect 4815 5516 4819 5520
rect 4825 5516 4829 5520
rect 4885 5516 4889 5520
rect 4905 5516 4909 5520
rect 4925 5516 4929 5520
rect 4993 5516 4997 5520
rect 5003 5516 5007 5520
rect 5075 5516 5079 5520
rect 5095 5516 5099 5520
rect 5105 5516 5109 5520
rect 5153 5516 5157 5520
rect 5163 5516 5167 5520
rect 5231 5516 5235 5520
rect 5251 5516 5255 5520
rect 5271 5516 5275 5520
rect 5355 5516 5359 5520
rect 5375 5516 5379 5520
rect 5385 5516 5389 5520
rect 5431 5516 5435 5520
rect 5451 5516 5455 5520
rect 5471 5516 5475 5520
rect 5533 5516 5537 5520
rect 5543 5516 5547 5520
rect 5612 5516 5616 5520
rect 5620 5516 5624 5520
rect 5628 5516 5632 5520
rect 5735 5516 5739 5520
rect 5755 5516 5759 5520
rect 5765 5516 5769 5520
rect 5846 5516 5850 5520
rect 5854 5516 5858 5520
rect 5874 5516 5878 5520
rect 5882 5516 5886 5520
rect 5933 5516 5937 5520
rect 5943 5516 5947 5520
rect 6012 5516 6016 5520
rect 6020 5516 6024 5520
rect 6028 5516 6032 5520
rect 6114 5516 6118 5520
rect 6122 5516 6126 5520
rect 6144 5516 6148 5520
rect 6225 5516 6229 5520
rect 6245 5516 6249 5520
rect 6265 5516 6269 5520
rect 6311 5516 6315 5520
rect 6331 5516 6335 5520
rect 6351 5516 6355 5520
rect 6425 5516 6429 5520
rect 6445 5516 6449 5520
rect 6465 5516 6469 5520
rect 6548 5516 6552 5520
rect 6556 5516 6560 5520
rect 6564 5516 6568 5520
rect 6632 5516 6636 5520
rect 6654 5516 6658 5520
rect 6662 5516 6666 5520
rect 31 5408 35 5476
rect 53 5447 57 5496
rect 63 5475 67 5496
rect 83 5484 87 5496
rect 91 5492 95 5496
rect 91 5488 125 5492
rect 83 5480 113 5484
rect 83 5479 101 5480
rect 63 5471 87 5475
rect 31 5396 33 5408
rect 31 5384 35 5396
rect 53 5389 57 5435
rect 49 5383 57 5389
rect 49 5354 53 5383
rect 81 5376 87 5471
rect 49 5347 57 5354
rect 53 5324 57 5347
rect 61 5324 65 5364
rect 81 5344 85 5376
rect 121 5362 125 5488
rect 137 5382 141 5496
rect 159 5484 163 5496
rect 161 5472 163 5484
rect 169 5484 173 5496
rect 169 5472 171 5484
rect 89 5350 113 5352
rect 89 5348 125 5350
rect 89 5344 93 5348
rect 135 5344 139 5370
rect 153 5362 157 5472
rect 191 5464 195 5496
rect 162 5460 195 5464
rect 162 5396 166 5460
rect 182 5411 186 5440
rect 201 5438 205 5496
rect 221 5439 225 5476
rect 273 5456 277 5476
rect 269 5449 277 5456
rect 283 5456 287 5476
rect 283 5449 297 5456
rect 372 5453 376 5496
rect 269 5433 275 5449
rect 182 5403 191 5411
rect 162 5384 165 5396
rect 155 5344 159 5350
rect 167 5344 171 5384
rect 187 5344 191 5403
rect 201 5344 205 5426
rect 221 5384 225 5427
rect 266 5421 275 5433
rect 271 5344 275 5421
rect 291 5433 297 5449
rect 365 5441 374 5453
rect 291 5421 294 5433
rect 291 5344 295 5421
rect 365 5384 369 5441
rect 394 5439 398 5476
rect 402 5472 406 5476
rect 402 5466 421 5472
rect 414 5453 421 5466
rect 473 5456 477 5476
rect 463 5449 477 5456
rect 483 5456 487 5476
rect 555 5470 559 5476
rect 541 5458 553 5470
rect 483 5449 491 5456
rect 394 5404 400 5427
rect 414 5404 421 5441
rect 463 5433 469 5449
rect 466 5421 469 5433
rect 385 5398 400 5404
rect 405 5398 421 5404
rect 385 5384 389 5398
rect 405 5384 409 5398
rect 465 5344 469 5421
rect 485 5433 491 5449
rect 485 5421 494 5433
rect 485 5344 489 5421
rect 541 5384 545 5458
rect 575 5433 579 5476
rect 566 5421 579 5433
rect 563 5344 567 5421
rect 585 5419 589 5476
rect 631 5419 635 5496
rect 651 5419 655 5496
rect 711 5419 715 5496
rect 731 5419 735 5496
rect 793 5456 797 5476
rect 789 5449 797 5456
rect 803 5456 807 5476
rect 873 5456 877 5476
rect 803 5449 817 5456
rect 789 5433 795 5449
rect 786 5421 795 5433
rect 585 5407 594 5419
rect 626 5407 635 5419
rect 585 5344 589 5407
rect 631 5384 635 5407
rect 639 5407 654 5419
rect 706 5407 715 5419
rect 639 5384 643 5407
rect 711 5384 715 5407
rect 719 5407 734 5419
rect 719 5384 723 5407
rect 791 5344 795 5421
rect 811 5433 817 5449
rect 869 5449 877 5456
rect 883 5456 887 5476
rect 883 5449 897 5456
rect 869 5433 875 5449
rect 811 5421 814 5433
rect 866 5421 875 5433
rect 811 5344 815 5421
rect 871 5344 875 5421
rect 891 5433 897 5449
rect 951 5439 955 5496
rect 1014 5472 1018 5476
rect 999 5466 1018 5472
rect 999 5453 1006 5466
rect 891 5421 894 5433
rect 946 5427 955 5439
rect 891 5344 895 5421
rect 951 5344 955 5427
rect 999 5404 1006 5441
rect 1022 5439 1026 5476
rect 1044 5453 1048 5496
rect 1146 5471 1150 5476
rect 1120 5467 1150 5471
rect 1046 5441 1055 5453
rect 1020 5404 1026 5427
rect 999 5398 1015 5404
rect 1020 5398 1035 5404
rect 1011 5384 1015 5398
rect 1031 5384 1035 5398
rect 1051 5384 1055 5441
rect 1120 5419 1126 5467
rect 1154 5462 1158 5476
rect 1145 5455 1158 5462
rect 1145 5453 1149 5455
rect 1174 5453 1178 5476
rect 1182 5468 1186 5476
rect 1182 5461 1199 5468
rect 1147 5441 1149 5453
rect 1126 5407 1129 5419
rect 1125 5384 1129 5407
rect 1145 5384 1149 5441
rect 1174 5412 1178 5441
rect 1193 5419 1199 5461
rect 1165 5406 1178 5412
rect 1185 5407 1193 5412
rect 1185 5406 1205 5407
rect 1231 5408 1235 5476
rect 1253 5447 1257 5496
rect 1263 5475 1267 5496
rect 1283 5484 1287 5496
rect 1291 5492 1295 5496
rect 1291 5488 1325 5492
rect 1283 5480 1313 5484
rect 1283 5479 1301 5480
rect 1263 5471 1287 5475
rect 1165 5384 1169 5406
rect 1185 5384 1189 5406
rect 1231 5396 1233 5408
rect 1231 5384 1235 5396
rect 1253 5389 1257 5435
rect 1249 5383 1257 5389
rect 1249 5354 1253 5383
rect 1281 5376 1287 5471
rect 1249 5347 1257 5354
rect 1253 5324 1257 5347
rect 1261 5324 1265 5364
rect 1281 5344 1285 5376
rect 1321 5362 1325 5488
rect 1337 5382 1341 5496
rect 1359 5484 1363 5496
rect 1361 5472 1363 5484
rect 1369 5484 1373 5496
rect 1369 5472 1371 5484
rect 1289 5350 1313 5352
rect 1289 5348 1325 5350
rect 1289 5344 1293 5348
rect 1335 5344 1339 5370
rect 1353 5362 1357 5472
rect 1391 5464 1395 5496
rect 1362 5460 1395 5464
rect 1362 5396 1366 5460
rect 1382 5411 1386 5440
rect 1401 5438 1405 5496
rect 1421 5439 1425 5476
rect 1382 5403 1391 5411
rect 1362 5384 1365 5396
rect 1355 5344 1359 5350
rect 1367 5344 1371 5384
rect 1387 5344 1391 5403
rect 1401 5344 1405 5426
rect 1421 5384 1425 5427
rect 1508 5399 1512 5456
rect 1485 5387 1493 5399
rect 1505 5387 1512 5399
rect 1485 5344 1489 5387
rect 1516 5379 1520 5456
rect 1524 5399 1528 5456
rect 1608 5399 1612 5456
rect 1524 5387 1534 5399
rect 1585 5387 1593 5399
rect 1605 5387 1612 5399
rect 1514 5360 1520 5367
rect 1505 5356 1520 5360
rect 1534 5356 1540 5387
rect 1505 5344 1509 5356
rect 1525 5352 1540 5356
rect 1525 5344 1529 5352
rect 1585 5344 1589 5387
rect 1616 5379 1620 5456
rect 1624 5399 1628 5456
rect 1685 5439 1689 5496
rect 1685 5427 1694 5439
rect 1624 5387 1634 5399
rect 1614 5360 1620 5367
rect 1605 5356 1620 5360
rect 1634 5356 1640 5387
rect 1605 5344 1609 5356
rect 1625 5352 1640 5356
rect 1625 5344 1629 5352
rect 1685 5344 1689 5427
rect 1745 5399 1749 5476
rect 1765 5453 1769 5476
rect 1785 5471 1789 5476
rect 1785 5464 1798 5471
rect 1855 5470 1859 5476
rect 1765 5441 1774 5453
rect 1747 5387 1754 5399
rect 1750 5344 1754 5387
rect 1772 5384 1776 5441
rect 1794 5419 1798 5464
rect 1841 5458 1853 5470
rect 1794 5396 1798 5407
rect 1780 5388 1798 5396
rect 1780 5384 1784 5388
rect 1841 5384 1845 5458
rect 1875 5433 1879 5476
rect 1866 5421 1879 5433
rect 1863 5344 1867 5421
rect 1885 5419 1889 5476
rect 1953 5456 1957 5476
rect 1943 5449 1957 5456
rect 1963 5456 1967 5476
rect 1963 5449 1971 5456
rect 1943 5433 1949 5449
rect 1946 5421 1949 5433
rect 1885 5407 1894 5419
rect 1885 5344 1889 5407
rect 1945 5344 1949 5421
rect 1965 5433 1971 5449
rect 1965 5421 1974 5433
rect 1965 5344 1969 5421
rect 2025 5399 2029 5476
rect 2045 5453 2049 5476
rect 2065 5471 2069 5476
rect 2065 5464 2078 5471
rect 2045 5441 2054 5453
rect 2027 5387 2034 5399
rect 2030 5344 2034 5387
rect 2052 5384 2056 5441
rect 2074 5419 2078 5464
rect 2113 5456 2117 5476
rect 2109 5449 2117 5456
rect 2123 5456 2127 5476
rect 2123 5449 2137 5456
rect 2109 5433 2115 5449
rect 2106 5421 2115 5433
rect 2074 5396 2078 5407
rect 2060 5388 2078 5396
rect 2060 5384 2064 5388
rect 2111 5344 2115 5421
rect 2131 5433 2137 5449
rect 2205 5439 2209 5496
rect 2131 5421 2134 5433
rect 2205 5427 2214 5439
rect 2131 5344 2135 5421
rect 2205 5344 2209 5427
rect 2265 5399 2269 5476
rect 2285 5453 2289 5476
rect 2305 5471 2309 5476
rect 2305 5464 2318 5471
rect 2285 5441 2294 5453
rect 2267 5387 2274 5399
rect 2270 5344 2274 5387
rect 2292 5384 2296 5441
rect 2314 5419 2318 5464
rect 2351 5419 2355 5496
rect 2371 5419 2375 5496
rect 2445 5439 2449 5496
rect 2512 5453 2516 5496
rect 2505 5441 2514 5453
rect 2445 5427 2454 5439
rect 2346 5407 2355 5419
rect 2314 5396 2318 5407
rect 2300 5388 2318 5396
rect 2300 5384 2304 5388
rect 2351 5384 2355 5407
rect 2359 5407 2374 5419
rect 2359 5384 2363 5407
rect 2445 5344 2449 5427
rect 2505 5384 2509 5441
rect 2534 5439 2538 5476
rect 2542 5472 2546 5476
rect 2542 5466 2561 5472
rect 2591 5471 2595 5476
rect 2554 5453 2561 5466
rect 2582 5464 2595 5471
rect 2534 5404 2540 5427
rect 2554 5404 2561 5441
rect 2582 5419 2586 5464
rect 2611 5453 2615 5476
rect 2606 5441 2615 5453
rect 2525 5398 2540 5404
rect 2545 5398 2561 5404
rect 2525 5384 2529 5398
rect 2545 5384 2549 5398
rect 2582 5396 2586 5407
rect 2582 5388 2600 5396
rect 2596 5384 2600 5388
rect 2604 5384 2608 5441
rect 2631 5399 2635 5476
rect 2693 5456 2697 5476
rect 2689 5449 2697 5456
rect 2703 5456 2707 5476
rect 2893 5456 2897 5476
rect 2703 5449 2717 5456
rect 2689 5433 2695 5449
rect 2686 5421 2695 5433
rect 2626 5387 2633 5399
rect 2626 5344 2630 5387
rect 2691 5344 2695 5421
rect 2711 5433 2717 5449
rect 2711 5421 2714 5433
rect 2711 5344 2715 5421
rect 2808 5399 2812 5456
rect 2785 5387 2793 5399
rect 2805 5387 2812 5399
rect 2785 5344 2789 5387
rect 2816 5379 2820 5456
rect 2824 5399 2828 5456
rect 2883 5449 2897 5456
rect 2903 5456 2907 5476
rect 2903 5449 2911 5456
rect 2883 5433 2889 5449
rect 2886 5421 2889 5433
rect 2824 5387 2834 5399
rect 2814 5360 2820 5367
rect 2805 5356 2820 5360
rect 2834 5356 2840 5387
rect 2805 5344 2809 5356
rect 2825 5352 2840 5356
rect 2825 5344 2829 5352
rect 2885 5344 2889 5421
rect 2905 5433 2911 5449
rect 2905 5421 2914 5433
rect 2905 5344 2909 5421
rect 2965 5419 2969 5496
rect 2985 5419 2989 5496
rect 3031 5471 3035 5476
rect 3022 5464 3035 5471
rect 3022 5419 3026 5464
rect 3051 5453 3055 5476
rect 3046 5441 3055 5453
rect 2966 5407 2981 5419
rect 2977 5384 2981 5407
rect 2985 5407 2994 5419
rect 2985 5384 2989 5407
rect 3022 5396 3026 5407
rect 3022 5388 3040 5396
rect 3036 5384 3040 5388
rect 3044 5384 3048 5441
rect 3071 5399 3075 5476
rect 3153 5456 3157 5476
rect 3143 5449 3157 5456
rect 3163 5456 3167 5476
rect 3211 5471 3215 5476
rect 3202 5464 3215 5471
rect 3163 5449 3171 5456
rect 3143 5433 3149 5449
rect 3146 5421 3149 5433
rect 3066 5387 3073 5399
rect 3066 5344 3070 5387
rect 3145 5344 3149 5421
rect 3165 5433 3171 5449
rect 3165 5421 3174 5433
rect 3165 5344 3169 5421
rect 3202 5419 3206 5464
rect 3231 5453 3235 5476
rect 3226 5441 3235 5453
rect 3202 5396 3206 5407
rect 3202 5388 3220 5396
rect 3216 5384 3220 5388
rect 3224 5384 3228 5441
rect 3251 5399 3255 5476
rect 3335 5470 3339 5476
rect 3321 5458 3333 5470
rect 3246 5387 3253 5399
rect 3246 5344 3250 5387
rect 3321 5384 3325 5458
rect 3355 5433 3359 5476
rect 3346 5421 3359 5433
rect 3343 5344 3347 5421
rect 3365 5419 3369 5476
rect 3411 5419 3415 5496
rect 3431 5419 3435 5496
rect 3491 5489 3495 5496
rect 3511 5489 3515 5496
rect 3482 5484 3495 5489
rect 3482 5439 3486 5484
rect 3365 5407 3374 5419
rect 3406 5407 3415 5419
rect 3365 5344 3369 5407
rect 3411 5384 3415 5407
rect 3419 5407 3434 5419
rect 3419 5384 3423 5407
rect 3482 5393 3486 5427
rect 3501 5483 3515 5489
rect 3501 5419 3505 5483
rect 3531 5468 3535 5476
rect 3591 5471 3595 5476
rect 3525 5456 3535 5468
rect 3582 5464 3595 5471
rect 3582 5419 3586 5464
rect 3611 5453 3615 5476
rect 3606 5441 3615 5453
rect 3482 5388 3495 5393
rect 3491 5384 3495 5388
rect 3501 5384 3505 5407
rect 3521 5384 3525 5389
rect 3582 5396 3586 5407
rect 3582 5388 3600 5396
rect 3596 5384 3600 5388
rect 3604 5384 3608 5441
rect 3631 5399 3635 5476
rect 3705 5419 3709 5496
rect 3725 5419 3729 5496
rect 3771 5469 3775 5476
rect 3760 5465 3775 5469
rect 3760 5419 3766 5465
rect 3791 5453 3795 5476
rect 3811 5453 3815 5476
rect 3786 5441 3795 5453
rect 3706 5407 3721 5419
rect 3626 5387 3633 5399
rect 3626 5344 3630 5387
rect 3717 5384 3721 5407
rect 3725 5407 3734 5419
rect 3725 5384 3729 5407
rect 3761 5392 3766 5407
rect 3789 5392 3795 5441
rect 3761 5388 3775 5392
rect 3771 5384 3775 5388
rect 3781 5388 3795 5392
rect 3781 5384 3785 5388
rect 3811 5384 3815 5441
rect 3831 5419 3835 5476
rect 3905 5419 3909 5496
rect 3925 5419 3929 5496
rect 3971 5471 3975 5476
rect 3962 5464 3975 5471
rect 3962 5419 3966 5464
rect 3991 5453 3995 5476
rect 3986 5441 3995 5453
rect 3831 5407 3833 5419
rect 3906 5407 3921 5419
rect 3831 5392 3835 5407
rect 3821 5388 3835 5392
rect 3821 5384 3825 5388
rect 3917 5384 3921 5407
rect 3925 5407 3934 5419
rect 3925 5384 3929 5407
rect 3962 5396 3966 5407
rect 3962 5388 3980 5396
rect 3976 5384 3980 5388
rect 3984 5384 3988 5441
rect 4011 5399 4015 5476
rect 4193 5456 4197 5476
rect 4108 5399 4112 5456
rect 4006 5387 4013 5399
rect 4085 5387 4093 5399
rect 4105 5387 4112 5399
rect 4006 5344 4010 5387
rect 4085 5344 4089 5387
rect 4116 5379 4120 5456
rect 4124 5399 4128 5456
rect 4183 5449 4197 5456
rect 4203 5456 4207 5476
rect 4203 5449 4211 5456
rect 4183 5433 4189 5449
rect 4186 5421 4189 5433
rect 4124 5387 4134 5399
rect 4114 5360 4120 5367
rect 4105 5356 4120 5360
rect 4134 5356 4140 5387
rect 4105 5344 4109 5356
rect 4125 5352 4140 5356
rect 4125 5344 4129 5352
rect 4185 5344 4189 5421
rect 4205 5433 4211 5449
rect 4251 5439 4255 5496
rect 4205 5421 4214 5433
rect 4246 5427 4255 5439
rect 4205 5344 4209 5421
rect 4251 5344 4255 5427
rect 4325 5399 4329 5476
rect 4345 5453 4349 5476
rect 4365 5471 4369 5476
rect 4365 5464 4378 5471
rect 4345 5441 4354 5453
rect 4327 5387 4334 5399
rect 4330 5344 4334 5387
rect 4352 5384 4356 5441
rect 4374 5419 4378 5464
rect 4433 5456 4437 5476
rect 4423 5449 4437 5456
rect 4443 5456 4447 5476
rect 4493 5456 4497 5476
rect 4443 5449 4451 5456
rect 4423 5433 4429 5449
rect 4426 5421 4429 5433
rect 4374 5396 4378 5407
rect 4360 5388 4378 5396
rect 4360 5384 4364 5388
rect 4425 5344 4429 5421
rect 4445 5433 4451 5449
rect 4489 5449 4497 5456
rect 4503 5456 4507 5476
rect 4503 5449 4517 5456
rect 4489 5433 4495 5449
rect 4445 5421 4454 5433
rect 4486 5421 4495 5433
rect 4445 5344 4449 5421
rect 4491 5344 4495 5421
rect 4511 5433 4517 5449
rect 4511 5421 4514 5433
rect 4511 5344 4515 5421
rect 4585 5399 4589 5476
rect 4605 5453 4609 5476
rect 4625 5471 4629 5476
rect 4625 5464 4638 5471
rect 4605 5441 4614 5453
rect 4587 5387 4594 5399
rect 4590 5344 4594 5387
rect 4612 5384 4616 5441
rect 4634 5419 4638 5464
rect 4634 5396 4638 5407
rect 4685 5399 4689 5476
rect 4705 5453 4709 5476
rect 4725 5471 4729 5476
rect 4725 5464 4738 5471
rect 4795 5470 4799 5476
rect 4705 5441 4714 5453
rect 4620 5388 4638 5396
rect 4620 5384 4624 5388
rect 4687 5387 4694 5399
rect 4690 5344 4694 5387
rect 4712 5384 4716 5441
rect 4734 5419 4738 5464
rect 4781 5458 4793 5470
rect 4734 5396 4738 5407
rect 4720 5388 4738 5396
rect 4720 5384 4724 5388
rect 4781 5384 4785 5458
rect 4815 5433 4819 5476
rect 4806 5421 4819 5433
rect 4803 5344 4807 5421
rect 4825 5419 4829 5476
rect 4825 5407 4834 5419
rect 4825 5344 4829 5407
rect 4885 5399 4889 5476
rect 4905 5453 4909 5476
rect 4925 5471 4929 5476
rect 4925 5464 4938 5471
rect 4905 5441 4914 5453
rect 4887 5387 4894 5399
rect 4890 5344 4894 5387
rect 4912 5384 4916 5441
rect 4934 5419 4938 5464
rect 4993 5456 4997 5476
rect 4983 5449 4997 5456
rect 5003 5456 5007 5476
rect 5075 5470 5079 5476
rect 5061 5458 5073 5470
rect 5003 5449 5011 5456
rect 4983 5433 4989 5449
rect 4986 5421 4989 5433
rect 4934 5396 4938 5407
rect 4920 5388 4938 5396
rect 4920 5384 4924 5388
rect 4985 5344 4989 5421
rect 5005 5433 5011 5449
rect 5005 5421 5014 5433
rect 5005 5344 5009 5421
rect 5061 5384 5065 5458
rect 5095 5433 5099 5476
rect 5086 5421 5099 5433
rect 5083 5344 5087 5421
rect 5105 5419 5109 5476
rect 5153 5456 5157 5476
rect 5149 5449 5157 5456
rect 5163 5456 5167 5476
rect 5231 5471 5235 5476
rect 5222 5464 5235 5471
rect 5163 5449 5177 5456
rect 5149 5433 5155 5449
rect 5146 5421 5155 5433
rect 5105 5407 5114 5419
rect 5105 5344 5109 5407
rect 5151 5344 5155 5421
rect 5171 5433 5177 5449
rect 5171 5421 5174 5433
rect 5171 5344 5175 5421
rect 5222 5419 5226 5464
rect 5251 5453 5255 5476
rect 5246 5441 5255 5453
rect 5222 5396 5226 5407
rect 5222 5388 5240 5396
rect 5236 5384 5240 5388
rect 5244 5384 5248 5441
rect 5271 5399 5275 5476
rect 5355 5470 5359 5476
rect 5341 5458 5353 5470
rect 5266 5387 5273 5399
rect 5266 5344 5270 5387
rect 5341 5384 5345 5458
rect 5375 5433 5379 5476
rect 5366 5421 5379 5433
rect 5363 5344 5367 5421
rect 5385 5419 5389 5476
rect 5431 5471 5435 5476
rect 5422 5464 5435 5471
rect 5422 5419 5426 5464
rect 5451 5453 5455 5476
rect 5446 5441 5455 5453
rect 5385 5407 5394 5419
rect 5385 5344 5389 5407
rect 5422 5396 5426 5407
rect 5422 5388 5440 5396
rect 5436 5384 5440 5388
rect 5444 5384 5448 5441
rect 5471 5399 5475 5476
rect 5533 5456 5537 5476
rect 5529 5449 5537 5456
rect 5543 5456 5547 5476
rect 5735 5470 5739 5476
rect 5721 5458 5733 5470
rect 5543 5449 5557 5456
rect 5529 5433 5535 5449
rect 5526 5421 5535 5433
rect 5466 5387 5473 5399
rect 5466 5344 5470 5387
rect 5531 5344 5535 5421
rect 5551 5433 5557 5449
rect 5551 5421 5554 5433
rect 5551 5344 5555 5421
rect 5612 5399 5616 5456
rect 5606 5387 5616 5399
rect 5600 5356 5606 5387
rect 5620 5379 5624 5456
rect 5628 5399 5632 5456
rect 5628 5387 5635 5399
rect 5647 5387 5655 5399
rect 5620 5360 5626 5367
rect 5620 5356 5635 5360
rect 5600 5352 5615 5356
rect 5611 5344 5615 5352
rect 5631 5344 5635 5356
rect 5651 5344 5655 5387
rect 5721 5384 5725 5458
rect 5755 5433 5759 5476
rect 5746 5421 5759 5433
rect 5743 5344 5747 5421
rect 5765 5419 5769 5476
rect 5846 5471 5850 5476
rect 5820 5467 5850 5471
rect 5820 5419 5826 5467
rect 5854 5462 5858 5476
rect 5845 5455 5858 5462
rect 5845 5453 5849 5455
rect 5874 5453 5878 5476
rect 5882 5468 5886 5476
rect 5882 5461 5899 5468
rect 5847 5441 5849 5453
rect 5765 5407 5774 5419
rect 5826 5407 5829 5419
rect 5765 5344 5769 5407
rect 5825 5384 5829 5407
rect 5845 5384 5849 5441
rect 5874 5412 5878 5441
rect 5893 5419 5899 5461
rect 5933 5456 5937 5476
rect 5929 5449 5937 5456
rect 5943 5456 5947 5476
rect 6114 5472 6118 5476
rect 6099 5466 6118 5472
rect 5943 5449 5957 5456
rect 5929 5433 5935 5449
rect 5926 5421 5935 5433
rect 5865 5406 5878 5412
rect 5885 5407 5893 5412
rect 5885 5406 5905 5407
rect 5865 5384 5869 5406
rect 5885 5384 5889 5406
rect 5931 5344 5935 5421
rect 5951 5433 5957 5449
rect 5951 5421 5954 5433
rect 5951 5344 5955 5421
rect 6012 5399 6016 5456
rect 6006 5387 6016 5399
rect 6000 5356 6006 5387
rect 6020 5379 6024 5456
rect 6028 5399 6032 5456
rect 6099 5453 6106 5466
rect 6099 5404 6106 5441
rect 6122 5439 6126 5476
rect 6144 5453 6148 5496
rect 6146 5441 6155 5453
rect 6120 5404 6126 5427
rect 6028 5387 6035 5399
rect 6047 5387 6055 5399
rect 6099 5398 6115 5404
rect 6120 5398 6135 5404
rect 6020 5360 6026 5367
rect 6020 5356 6035 5360
rect 6000 5352 6015 5356
rect 6011 5344 6015 5352
rect 6031 5344 6035 5356
rect 6051 5344 6055 5387
rect 6111 5384 6115 5398
rect 6131 5384 6135 5398
rect 6151 5384 6155 5441
rect 6225 5399 6229 5476
rect 6245 5453 6249 5476
rect 6265 5471 6269 5476
rect 6311 5471 6315 5476
rect 6265 5464 6278 5471
rect 6245 5441 6254 5453
rect 6227 5387 6234 5399
rect 6230 5344 6234 5387
rect 6252 5384 6256 5441
rect 6274 5419 6278 5464
rect 6302 5464 6315 5471
rect 6302 5419 6306 5464
rect 6331 5453 6335 5476
rect 6326 5441 6335 5453
rect 6274 5396 6278 5407
rect 6260 5388 6278 5396
rect 6302 5396 6306 5407
rect 6302 5388 6320 5396
rect 6260 5384 6264 5388
rect 6316 5384 6320 5388
rect 6324 5384 6328 5441
rect 6351 5399 6355 5476
rect 6425 5399 6429 5476
rect 6445 5453 6449 5476
rect 6465 5471 6469 5476
rect 6465 5464 6478 5471
rect 6445 5441 6454 5453
rect 6346 5387 6353 5399
rect 6427 5387 6434 5399
rect 6346 5344 6350 5387
rect 6430 5344 6434 5387
rect 6452 5384 6456 5441
rect 6474 5419 6478 5464
rect 6474 5396 6478 5407
rect 6548 5399 6552 5456
rect 6460 5388 6478 5396
rect 6460 5384 6464 5388
rect 6525 5387 6533 5399
rect 6545 5387 6552 5399
rect 6525 5344 6529 5387
rect 6556 5379 6560 5456
rect 6564 5399 6568 5456
rect 6632 5453 6636 5496
rect 6625 5441 6634 5453
rect 6564 5387 6574 5399
rect 6554 5360 6560 5367
rect 6545 5356 6560 5360
rect 6574 5356 6580 5387
rect 6625 5384 6629 5441
rect 6654 5439 6658 5476
rect 6662 5472 6666 5476
rect 6662 5466 6681 5472
rect 6674 5453 6681 5466
rect 6654 5404 6660 5427
rect 6674 5404 6681 5441
rect 6645 5398 6660 5404
rect 6665 5398 6681 5404
rect 6645 5384 6649 5398
rect 6665 5384 6669 5398
rect 6545 5344 6549 5356
rect 6565 5352 6580 5356
rect 6565 5344 6569 5352
rect 31 5300 35 5304
rect 53 5300 57 5304
rect 61 5300 65 5304
rect 81 5300 85 5304
rect 89 5300 93 5304
rect 135 5300 139 5304
rect 155 5300 159 5304
rect 167 5300 171 5304
rect 187 5300 191 5304
rect 201 5300 205 5304
rect 221 5300 225 5304
rect 271 5300 275 5304
rect 291 5300 295 5304
rect 365 5300 369 5304
rect 385 5300 389 5304
rect 405 5300 409 5304
rect 465 5300 469 5304
rect 485 5300 489 5304
rect 541 5300 545 5304
rect 563 5300 567 5304
rect 585 5300 589 5304
rect 631 5300 635 5304
rect 639 5300 643 5304
rect 711 5300 715 5304
rect 719 5300 723 5304
rect 791 5300 795 5304
rect 811 5300 815 5304
rect 871 5300 875 5304
rect 891 5300 895 5304
rect 951 5300 955 5304
rect 1011 5300 1015 5304
rect 1031 5300 1035 5304
rect 1051 5300 1055 5304
rect 1125 5300 1129 5304
rect 1145 5300 1149 5304
rect 1165 5300 1169 5304
rect 1185 5300 1189 5304
rect 1231 5300 1235 5304
rect 1253 5300 1257 5304
rect 1261 5300 1265 5304
rect 1281 5300 1285 5304
rect 1289 5300 1293 5304
rect 1335 5300 1339 5304
rect 1355 5300 1359 5304
rect 1367 5300 1371 5304
rect 1387 5300 1391 5304
rect 1401 5300 1405 5304
rect 1421 5300 1425 5304
rect 1485 5300 1489 5304
rect 1505 5300 1509 5304
rect 1525 5300 1529 5304
rect 1585 5300 1589 5304
rect 1605 5300 1609 5304
rect 1625 5300 1629 5304
rect 1685 5300 1689 5304
rect 1750 5300 1754 5304
rect 1772 5300 1776 5304
rect 1780 5300 1784 5304
rect 1841 5300 1845 5304
rect 1863 5300 1867 5304
rect 1885 5300 1889 5304
rect 1945 5300 1949 5304
rect 1965 5300 1969 5304
rect 2030 5300 2034 5304
rect 2052 5300 2056 5304
rect 2060 5300 2064 5304
rect 2111 5300 2115 5304
rect 2131 5300 2135 5304
rect 2205 5300 2209 5304
rect 2270 5300 2274 5304
rect 2292 5300 2296 5304
rect 2300 5300 2304 5304
rect 2351 5300 2355 5304
rect 2359 5300 2363 5304
rect 2445 5300 2449 5304
rect 2505 5300 2509 5304
rect 2525 5300 2529 5304
rect 2545 5300 2549 5304
rect 2596 5300 2600 5304
rect 2604 5300 2608 5304
rect 2626 5300 2630 5304
rect 2691 5300 2695 5304
rect 2711 5300 2715 5304
rect 2785 5300 2789 5304
rect 2805 5300 2809 5304
rect 2825 5300 2829 5304
rect 2885 5300 2889 5304
rect 2905 5300 2909 5304
rect 2977 5300 2981 5304
rect 2985 5300 2989 5304
rect 3036 5300 3040 5304
rect 3044 5300 3048 5304
rect 3066 5300 3070 5304
rect 3145 5300 3149 5304
rect 3165 5300 3169 5304
rect 3216 5300 3220 5304
rect 3224 5300 3228 5304
rect 3246 5300 3250 5304
rect 3321 5300 3325 5304
rect 3343 5300 3347 5304
rect 3365 5300 3369 5304
rect 3411 5300 3415 5304
rect 3419 5300 3423 5304
rect 3491 5300 3495 5304
rect 3501 5300 3505 5304
rect 3521 5300 3525 5304
rect 3596 5300 3600 5304
rect 3604 5300 3608 5304
rect 3626 5300 3630 5304
rect 3717 5300 3721 5304
rect 3725 5300 3729 5304
rect 3771 5300 3775 5304
rect 3781 5300 3785 5304
rect 3811 5300 3815 5304
rect 3821 5300 3825 5304
rect 3917 5300 3921 5304
rect 3925 5300 3929 5304
rect 3976 5300 3980 5304
rect 3984 5300 3988 5304
rect 4006 5300 4010 5304
rect 4085 5300 4089 5304
rect 4105 5300 4109 5304
rect 4125 5300 4129 5304
rect 4185 5300 4189 5304
rect 4205 5300 4209 5304
rect 4251 5300 4255 5304
rect 4330 5300 4334 5304
rect 4352 5300 4356 5304
rect 4360 5300 4364 5304
rect 4425 5300 4429 5304
rect 4445 5300 4449 5304
rect 4491 5300 4495 5304
rect 4511 5300 4515 5304
rect 4590 5300 4594 5304
rect 4612 5300 4616 5304
rect 4620 5300 4624 5304
rect 4690 5300 4694 5304
rect 4712 5300 4716 5304
rect 4720 5300 4724 5304
rect 4781 5300 4785 5304
rect 4803 5300 4807 5304
rect 4825 5300 4829 5304
rect 4890 5300 4894 5304
rect 4912 5300 4916 5304
rect 4920 5300 4924 5304
rect 4985 5300 4989 5304
rect 5005 5300 5009 5304
rect 5061 5300 5065 5304
rect 5083 5300 5087 5304
rect 5105 5300 5109 5304
rect 5151 5300 5155 5304
rect 5171 5300 5175 5304
rect 5236 5300 5240 5304
rect 5244 5300 5248 5304
rect 5266 5300 5270 5304
rect 5341 5300 5345 5304
rect 5363 5300 5367 5304
rect 5385 5300 5389 5304
rect 5436 5300 5440 5304
rect 5444 5300 5448 5304
rect 5466 5300 5470 5304
rect 5531 5300 5535 5304
rect 5551 5300 5555 5304
rect 5611 5300 5615 5304
rect 5631 5300 5635 5304
rect 5651 5300 5655 5304
rect 5721 5300 5725 5304
rect 5743 5300 5747 5304
rect 5765 5300 5769 5304
rect 5825 5300 5829 5304
rect 5845 5300 5849 5304
rect 5865 5300 5869 5304
rect 5885 5300 5889 5304
rect 5931 5300 5935 5304
rect 5951 5300 5955 5304
rect 6011 5300 6015 5304
rect 6031 5300 6035 5304
rect 6051 5300 6055 5304
rect 6111 5300 6115 5304
rect 6131 5300 6135 5304
rect 6151 5300 6155 5304
rect 6230 5300 6234 5304
rect 6252 5300 6256 5304
rect 6260 5300 6264 5304
rect 6316 5300 6320 5304
rect 6324 5300 6328 5304
rect 6346 5300 6350 5304
rect 6430 5300 6434 5304
rect 6452 5300 6456 5304
rect 6460 5300 6464 5304
rect 6525 5300 6529 5304
rect 6545 5300 6549 5304
rect 6565 5300 6569 5304
rect 6625 5300 6629 5304
rect 6645 5300 6649 5304
rect 6665 5300 6669 5304
rect 43 5276 47 5280
rect 65 5276 69 5280
rect 111 5276 115 5280
rect 133 5276 137 5280
rect 141 5276 145 5280
rect 161 5276 165 5280
rect 169 5276 173 5280
rect 215 5276 219 5280
rect 235 5276 239 5280
rect 247 5276 251 5280
rect 267 5276 271 5280
rect 281 5276 285 5280
rect 301 5276 305 5280
rect 351 5276 355 5280
rect 371 5276 375 5280
rect 445 5276 449 5280
rect 465 5276 469 5280
rect 485 5276 489 5280
rect 545 5276 549 5280
rect 565 5276 569 5280
rect 615 5276 619 5280
rect 635 5276 639 5280
rect 649 5276 653 5280
rect 669 5276 673 5280
rect 681 5276 685 5280
rect 701 5276 705 5280
rect 747 5276 751 5280
rect 755 5276 759 5280
rect 775 5276 779 5280
rect 783 5276 787 5280
rect 805 5276 809 5280
rect 851 5276 855 5280
rect 871 5276 875 5280
rect 950 5276 954 5280
rect 972 5276 976 5280
rect 980 5276 984 5280
rect 1050 5276 1054 5280
rect 1072 5276 1076 5280
rect 1080 5276 1084 5280
rect 1141 5276 1145 5280
rect 1163 5276 1167 5280
rect 1185 5276 1189 5280
rect 1231 5276 1235 5280
rect 1253 5276 1257 5280
rect 1261 5276 1265 5280
rect 1281 5276 1285 5280
rect 1289 5276 1293 5280
rect 1335 5276 1339 5280
rect 1355 5276 1359 5280
rect 1367 5276 1371 5280
rect 1387 5276 1391 5280
rect 1401 5276 1405 5280
rect 1421 5276 1425 5280
rect 1485 5276 1489 5280
rect 1505 5276 1509 5280
rect 1551 5276 1555 5280
rect 1571 5276 1575 5280
rect 1631 5276 1635 5280
rect 1653 5276 1657 5280
rect 1661 5276 1665 5280
rect 1681 5276 1685 5280
rect 1689 5276 1693 5280
rect 1735 5276 1739 5280
rect 1755 5276 1759 5280
rect 1767 5276 1771 5280
rect 1787 5276 1791 5280
rect 1801 5276 1805 5280
rect 1821 5276 1825 5280
rect 1885 5276 1889 5280
rect 1905 5276 1909 5280
rect 1925 5276 1929 5280
rect 1945 5276 1949 5280
rect 1991 5276 1995 5280
rect 2061 5276 2065 5280
rect 2083 5276 2087 5280
rect 2105 5276 2109 5280
rect 2151 5276 2155 5280
rect 2171 5276 2175 5280
rect 2255 5276 2259 5280
rect 2275 5276 2279 5280
rect 2285 5276 2289 5280
rect 2345 5276 2349 5280
rect 2365 5276 2369 5280
rect 2425 5276 2429 5280
rect 2445 5276 2449 5280
rect 2465 5276 2469 5280
rect 2537 5276 2541 5280
rect 2545 5276 2549 5280
rect 2591 5276 2595 5280
rect 2661 5276 2665 5280
rect 2683 5276 2687 5280
rect 2705 5276 2709 5280
rect 2751 5276 2755 5280
rect 2759 5276 2763 5280
rect 2845 5276 2849 5280
rect 2865 5276 2869 5280
rect 2925 5276 2929 5280
rect 2945 5276 2949 5280
rect 2991 5276 2995 5280
rect 3001 5276 3005 5280
rect 3021 5276 3025 5280
rect 3101 5276 3105 5280
rect 3123 5276 3127 5280
rect 3145 5276 3149 5280
rect 3191 5276 3195 5280
rect 3211 5276 3215 5280
rect 3285 5276 3289 5280
rect 3305 5276 3309 5280
rect 3325 5276 3329 5280
rect 3385 5276 3389 5280
rect 3445 5276 3449 5280
rect 3465 5276 3469 5280
rect 3485 5276 3489 5280
rect 3557 5276 3561 5280
rect 3565 5276 3569 5280
rect 3616 5276 3620 5280
rect 3624 5276 3628 5280
rect 3646 5276 3650 5280
rect 3730 5276 3734 5280
rect 3752 5276 3756 5280
rect 3760 5276 3764 5280
rect 3811 5276 3815 5280
rect 3819 5276 3823 5280
rect 3891 5276 3895 5280
rect 3911 5276 3915 5280
rect 3985 5276 3989 5280
rect 4005 5276 4009 5280
rect 4056 5276 4060 5280
rect 4064 5276 4068 5280
rect 4086 5276 4090 5280
rect 4165 5276 4169 5280
rect 4185 5276 4189 5280
rect 4241 5276 4245 5280
rect 4263 5276 4267 5280
rect 4285 5276 4289 5280
rect 4345 5276 4349 5280
rect 4365 5276 4369 5280
rect 4430 5276 4434 5280
rect 4452 5276 4456 5280
rect 4460 5276 4464 5280
rect 4530 5276 4534 5280
rect 4552 5276 4556 5280
rect 4560 5276 4564 5280
rect 4611 5276 4615 5280
rect 4631 5276 4635 5280
rect 4691 5276 4695 5280
rect 4711 5276 4715 5280
rect 4771 5276 4775 5280
rect 4845 5276 4849 5280
rect 4865 5276 4869 5280
rect 4885 5276 4889 5280
rect 4936 5276 4940 5280
rect 4944 5276 4948 5280
rect 4966 5276 4970 5280
rect 5031 5276 5035 5280
rect 5091 5276 5095 5280
rect 5111 5276 5115 5280
rect 5171 5276 5175 5280
rect 5191 5276 5195 5280
rect 5251 5276 5255 5280
rect 5271 5276 5275 5280
rect 5336 5276 5340 5280
rect 5344 5276 5348 5280
rect 5366 5276 5370 5280
rect 5431 5276 5435 5280
rect 5451 5276 5455 5280
rect 5471 5276 5475 5280
rect 5531 5276 5535 5280
rect 5551 5276 5555 5280
rect 5571 5276 5575 5280
rect 5631 5276 5635 5280
rect 5691 5276 5695 5280
rect 5711 5276 5715 5280
rect 5731 5276 5735 5280
rect 5796 5276 5800 5280
rect 5804 5276 5808 5280
rect 5826 5276 5830 5280
rect 5905 5276 5909 5280
rect 5925 5276 5929 5280
rect 5971 5276 5975 5280
rect 5991 5276 5995 5280
rect 6011 5276 6015 5280
rect 6071 5276 6075 5280
rect 6091 5276 6095 5280
rect 6165 5276 6169 5280
rect 6185 5276 6189 5280
rect 6205 5276 6209 5280
rect 6265 5276 6269 5280
rect 6325 5276 6329 5280
rect 6345 5276 6349 5280
rect 6365 5276 6369 5280
rect 6425 5276 6429 5280
rect 6445 5276 6449 5280
rect 6465 5276 6469 5280
rect 6511 5276 6515 5280
rect 6585 5276 6589 5280
rect 6605 5276 6609 5280
rect 6625 5276 6629 5280
rect 6671 5276 6675 5280
rect 6691 5276 6695 5280
rect 43 5190 47 5196
rect 43 5178 45 5190
rect 65 5173 69 5236
rect 133 5233 137 5256
rect 129 5226 137 5233
rect 129 5197 133 5226
rect 141 5216 145 5256
rect 161 5204 165 5236
rect 169 5232 173 5236
rect 169 5230 205 5232
rect 169 5228 193 5230
rect 111 5184 115 5196
rect 129 5191 137 5197
rect 65 5161 74 5173
rect 111 5172 113 5184
rect 43 5110 45 5122
rect 43 5104 47 5110
rect 65 5084 69 5161
rect 111 5104 115 5172
rect 133 5145 137 5191
rect 133 5084 137 5133
rect 161 5109 167 5204
rect 143 5105 167 5109
rect 143 5084 147 5105
rect 163 5100 181 5101
rect 163 5096 193 5100
rect 163 5084 167 5096
rect 201 5092 205 5218
rect 215 5210 219 5236
rect 235 5230 239 5236
rect 171 5088 205 5092
rect 171 5084 175 5088
rect 217 5084 221 5198
rect 233 5108 237 5218
rect 247 5196 251 5236
rect 242 5184 245 5196
rect 242 5120 246 5184
rect 267 5177 271 5236
rect 262 5169 271 5177
rect 262 5140 266 5169
rect 281 5154 285 5236
rect 301 5153 305 5196
rect 351 5159 355 5236
rect 242 5116 275 5120
rect 241 5096 243 5108
rect 239 5084 243 5096
rect 249 5096 251 5108
rect 249 5084 253 5096
rect 271 5084 275 5116
rect 281 5084 285 5142
rect 346 5147 355 5159
rect 301 5104 305 5141
rect 349 5131 355 5147
rect 371 5159 375 5236
rect 371 5147 374 5159
rect 371 5131 377 5147
rect 349 5124 357 5131
rect 353 5104 357 5124
rect 363 5124 377 5131
rect 445 5139 449 5196
rect 465 5182 469 5196
rect 485 5182 489 5196
rect 465 5176 480 5182
rect 485 5176 501 5182
rect 474 5153 480 5176
rect 445 5127 454 5139
rect 363 5104 367 5124
rect 452 5084 456 5127
rect 474 5104 478 5141
rect 494 5139 501 5176
rect 545 5159 549 5236
rect 546 5147 549 5159
rect 543 5131 549 5147
rect 565 5159 569 5236
rect 565 5147 574 5159
rect 615 5153 619 5196
rect 635 5154 639 5236
rect 649 5177 653 5236
rect 669 5196 673 5236
rect 681 5230 685 5236
rect 675 5184 678 5196
rect 649 5169 658 5177
rect 565 5131 571 5147
rect 494 5114 501 5127
rect 543 5124 557 5131
rect 482 5108 501 5114
rect 482 5104 486 5108
rect 553 5104 557 5124
rect 563 5124 571 5131
rect 563 5104 567 5124
rect 615 5104 619 5141
rect 635 5084 639 5142
rect 654 5140 658 5169
rect 674 5120 678 5184
rect 645 5116 678 5120
rect 645 5084 649 5116
rect 683 5108 687 5218
rect 701 5210 705 5236
rect 747 5232 751 5236
rect 715 5230 751 5232
rect 727 5228 751 5230
rect 669 5096 671 5108
rect 667 5084 671 5096
rect 677 5096 679 5108
rect 677 5084 681 5096
rect 699 5084 703 5198
rect 715 5092 719 5218
rect 755 5204 759 5236
rect 775 5216 779 5256
rect 783 5233 787 5256
rect 783 5226 791 5233
rect 753 5109 759 5204
rect 787 5197 791 5226
rect 783 5191 791 5197
rect 783 5145 787 5191
rect 805 5184 809 5196
rect 807 5172 809 5184
rect 753 5105 777 5109
rect 739 5100 757 5101
rect 727 5096 757 5100
rect 715 5088 749 5092
rect 745 5084 749 5088
rect 753 5084 757 5096
rect 773 5084 777 5105
rect 783 5084 787 5133
rect 805 5104 809 5172
rect 851 5159 855 5236
rect 846 5147 855 5159
rect 849 5131 855 5147
rect 871 5159 875 5236
rect 950 5193 954 5236
rect 947 5181 954 5193
rect 871 5147 874 5159
rect 871 5131 877 5147
rect 849 5124 857 5131
rect 853 5104 857 5124
rect 863 5124 877 5131
rect 863 5104 867 5124
rect 945 5104 949 5181
rect 972 5139 976 5196
rect 980 5192 984 5196
rect 1050 5193 1054 5236
rect 980 5184 998 5192
rect 994 5173 998 5184
rect 1047 5181 1054 5193
rect 965 5127 974 5139
rect 965 5104 969 5127
rect 994 5116 998 5161
rect 985 5109 998 5116
rect 985 5104 989 5109
rect 1045 5104 1049 5181
rect 1072 5139 1076 5196
rect 1080 5192 1084 5196
rect 1080 5184 1098 5192
rect 1094 5173 1098 5184
rect 1065 5127 1074 5139
rect 1065 5104 1069 5127
rect 1094 5116 1098 5161
rect 1085 5109 1098 5116
rect 1141 5122 1145 5196
rect 1163 5159 1167 5236
rect 1185 5173 1189 5236
rect 1253 5233 1257 5256
rect 1249 5226 1257 5233
rect 1249 5197 1253 5226
rect 1261 5216 1265 5256
rect 1281 5204 1285 5236
rect 1289 5232 1293 5236
rect 1289 5230 1325 5232
rect 1289 5228 1313 5230
rect 1231 5184 1235 5196
rect 1249 5191 1257 5197
rect 1185 5161 1194 5173
rect 1231 5172 1233 5184
rect 1166 5147 1179 5159
rect 1141 5110 1153 5122
rect 1085 5104 1089 5109
rect 1155 5104 1159 5110
rect 1175 5104 1179 5147
rect 1185 5104 1189 5161
rect 1231 5104 1235 5172
rect 1253 5145 1257 5191
rect 1253 5084 1257 5133
rect 1281 5109 1287 5204
rect 1263 5105 1287 5109
rect 1263 5084 1267 5105
rect 1283 5100 1301 5101
rect 1283 5096 1313 5100
rect 1283 5084 1287 5096
rect 1321 5092 1325 5218
rect 1335 5210 1339 5236
rect 1355 5230 1359 5236
rect 1291 5088 1325 5092
rect 1291 5084 1295 5088
rect 1337 5084 1341 5198
rect 1353 5108 1357 5218
rect 1367 5196 1371 5236
rect 1362 5184 1365 5196
rect 1362 5120 1366 5184
rect 1387 5177 1391 5236
rect 1382 5169 1391 5177
rect 1382 5140 1386 5169
rect 1401 5154 1405 5236
rect 1421 5153 1425 5196
rect 1485 5159 1489 5236
rect 1362 5116 1395 5120
rect 1361 5096 1363 5108
rect 1359 5084 1363 5096
rect 1369 5096 1371 5108
rect 1369 5084 1373 5096
rect 1391 5084 1395 5116
rect 1401 5084 1405 5142
rect 1486 5147 1489 5159
rect 1421 5104 1425 5141
rect 1483 5131 1489 5147
rect 1505 5159 1509 5236
rect 1551 5159 1555 5236
rect 1505 5147 1514 5159
rect 1546 5147 1555 5159
rect 1505 5131 1511 5147
rect 1483 5124 1497 5131
rect 1493 5104 1497 5124
rect 1503 5124 1511 5131
rect 1549 5131 1555 5147
rect 1571 5159 1575 5236
rect 1653 5233 1657 5256
rect 1649 5226 1657 5233
rect 1649 5197 1653 5226
rect 1661 5216 1665 5256
rect 1681 5204 1685 5236
rect 1689 5232 1693 5236
rect 1689 5230 1725 5232
rect 1689 5228 1713 5230
rect 1631 5184 1635 5196
rect 1649 5191 1657 5197
rect 1631 5172 1633 5184
rect 1571 5147 1574 5159
rect 1571 5131 1577 5147
rect 1549 5124 1557 5131
rect 1503 5104 1507 5124
rect 1553 5104 1557 5124
rect 1563 5124 1577 5131
rect 1563 5104 1567 5124
rect 1631 5104 1635 5172
rect 1653 5145 1657 5191
rect 1653 5084 1657 5133
rect 1681 5109 1687 5204
rect 1663 5105 1687 5109
rect 1663 5084 1667 5105
rect 1683 5100 1701 5101
rect 1683 5096 1713 5100
rect 1683 5084 1687 5096
rect 1721 5092 1725 5218
rect 1735 5210 1739 5236
rect 1755 5230 1759 5236
rect 1691 5088 1725 5092
rect 1691 5084 1695 5088
rect 1737 5084 1741 5198
rect 1753 5108 1757 5218
rect 1767 5196 1771 5236
rect 1762 5184 1765 5196
rect 1762 5120 1766 5184
rect 1787 5177 1791 5236
rect 1782 5169 1791 5177
rect 1782 5140 1786 5169
rect 1801 5154 1805 5236
rect 1821 5153 1825 5196
rect 1885 5173 1889 5196
rect 1886 5161 1889 5173
rect 1762 5116 1795 5120
rect 1761 5096 1763 5108
rect 1759 5084 1763 5096
rect 1769 5096 1771 5108
rect 1769 5084 1773 5096
rect 1791 5084 1795 5116
rect 1801 5084 1805 5142
rect 1821 5104 1825 5141
rect 1880 5113 1886 5161
rect 1905 5139 1909 5196
rect 1925 5174 1929 5196
rect 1945 5174 1949 5196
rect 1925 5168 1938 5174
rect 1945 5173 1965 5174
rect 1945 5168 1953 5173
rect 1934 5139 1938 5168
rect 1907 5127 1909 5139
rect 1905 5125 1909 5127
rect 1905 5118 1918 5125
rect 1880 5109 1910 5113
rect 1906 5104 1910 5109
rect 1914 5104 1918 5118
rect 1934 5104 1938 5127
rect 1953 5119 1959 5161
rect 1991 5153 1995 5236
rect 1986 5141 1995 5153
rect 1942 5112 1959 5119
rect 1942 5104 1946 5112
rect 1991 5084 1995 5141
rect 2061 5122 2065 5196
rect 2083 5159 2087 5236
rect 2105 5173 2109 5236
rect 2105 5161 2114 5173
rect 2086 5147 2099 5159
rect 2061 5110 2073 5122
rect 2075 5104 2079 5110
rect 2095 5104 2099 5147
rect 2105 5104 2109 5161
rect 2151 5159 2155 5236
rect 2146 5147 2155 5159
rect 2149 5131 2155 5147
rect 2171 5159 2175 5236
rect 2255 5191 2259 5196
rect 2275 5173 2279 5196
rect 2285 5192 2289 5196
rect 2285 5187 2298 5192
rect 2171 5147 2174 5159
rect 2171 5131 2177 5147
rect 2149 5124 2157 5131
rect 2153 5104 2157 5124
rect 2163 5124 2177 5131
rect 2163 5104 2167 5124
rect 2245 5112 2255 5124
rect 2245 5104 2249 5112
rect 2275 5097 2279 5161
rect 2265 5091 2279 5097
rect 2294 5153 2298 5187
rect 2345 5159 2349 5236
rect 2346 5147 2349 5159
rect 2294 5096 2298 5141
rect 2343 5131 2349 5147
rect 2365 5159 2369 5236
rect 2425 5193 2429 5236
rect 2445 5224 2449 5236
rect 2465 5228 2469 5236
rect 2465 5224 2480 5228
rect 2445 5220 2460 5224
rect 2454 5213 2460 5220
rect 2425 5181 2433 5193
rect 2445 5181 2452 5193
rect 2365 5147 2374 5159
rect 2365 5131 2371 5147
rect 2343 5124 2357 5131
rect 2353 5104 2357 5124
rect 2363 5124 2371 5131
rect 2448 5124 2452 5181
rect 2456 5124 2460 5201
rect 2474 5193 2480 5224
rect 2464 5181 2474 5193
rect 2464 5124 2468 5181
rect 2537 5173 2541 5196
rect 2526 5161 2541 5173
rect 2545 5173 2549 5196
rect 2545 5161 2554 5173
rect 2363 5104 2367 5124
rect 2285 5091 2298 5096
rect 2265 5084 2269 5091
rect 2285 5084 2289 5091
rect 2525 5084 2529 5161
rect 2545 5084 2549 5161
rect 2591 5153 2595 5236
rect 2586 5141 2595 5153
rect 2591 5084 2595 5141
rect 2661 5122 2665 5196
rect 2683 5159 2687 5236
rect 2705 5173 2709 5236
rect 2751 5173 2755 5196
rect 2705 5161 2714 5173
rect 2746 5161 2755 5173
rect 2759 5173 2763 5196
rect 2759 5161 2774 5173
rect 2686 5147 2699 5159
rect 2661 5110 2673 5122
rect 2675 5104 2679 5110
rect 2695 5104 2699 5147
rect 2705 5104 2709 5161
rect 2751 5084 2755 5161
rect 2771 5084 2775 5161
rect 2845 5159 2849 5236
rect 2846 5147 2849 5159
rect 2843 5131 2849 5147
rect 2865 5159 2869 5236
rect 2925 5159 2929 5236
rect 2865 5147 2874 5159
rect 2926 5147 2929 5159
rect 2865 5131 2871 5147
rect 2843 5124 2857 5131
rect 2853 5104 2857 5124
rect 2863 5124 2871 5131
rect 2923 5131 2929 5147
rect 2945 5159 2949 5236
rect 2991 5192 2995 5196
rect 2982 5187 2995 5192
rect 2945 5147 2954 5159
rect 2982 5153 2986 5187
rect 3001 5173 3005 5196
rect 3021 5191 3025 5196
rect 2945 5131 2951 5147
rect 2923 5124 2937 5131
rect 2863 5104 2867 5124
rect 2933 5104 2937 5124
rect 2943 5124 2951 5131
rect 2943 5104 2947 5124
rect 2982 5096 2986 5141
rect 3001 5097 3005 5161
rect 3025 5112 3035 5124
rect 3031 5104 3035 5112
rect 3101 5122 3105 5196
rect 3123 5159 3127 5236
rect 3145 5173 3149 5236
rect 3145 5161 3154 5173
rect 3126 5147 3139 5159
rect 3101 5110 3113 5122
rect 3115 5104 3119 5110
rect 3135 5104 3139 5147
rect 3145 5104 3149 5161
rect 3191 5159 3195 5236
rect 3186 5147 3195 5159
rect 3189 5131 3195 5147
rect 3211 5159 3215 5236
rect 3285 5193 3289 5236
rect 3305 5224 3309 5236
rect 3325 5228 3329 5236
rect 3325 5224 3340 5228
rect 3305 5220 3320 5224
rect 3314 5213 3320 5220
rect 3285 5181 3293 5193
rect 3305 5181 3312 5193
rect 3211 5147 3214 5159
rect 3211 5131 3217 5147
rect 3189 5124 3197 5131
rect 3193 5104 3197 5124
rect 3203 5124 3217 5131
rect 3308 5124 3312 5181
rect 3316 5124 3320 5201
rect 3334 5193 3340 5224
rect 3324 5181 3334 5193
rect 3324 5124 3328 5181
rect 3385 5153 3389 5236
rect 3385 5141 3394 5153
rect 3203 5104 3207 5124
rect 2982 5091 2995 5096
rect 3001 5091 3015 5097
rect 2991 5084 2995 5091
rect 3011 5084 3015 5091
rect 3385 5084 3389 5141
rect 3445 5139 3449 5196
rect 3465 5182 3469 5196
rect 3485 5182 3489 5196
rect 3465 5176 3480 5182
rect 3485 5176 3501 5182
rect 3474 5153 3480 5176
rect 3445 5127 3454 5139
rect 3452 5084 3456 5127
rect 3474 5104 3478 5141
rect 3494 5139 3501 5176
rect 3557 5173 3561 5196
rect 3546 5161 3561 5173
rect 3565 5173 3569 5196
rect 3616 5192 3620 5196
rect 3602 5184 3620 5192
rect 3602 5173 3606 5184
rect 3565 5161 3574 5173
rect 3494 5114 3501 5127
rect 3482 5108 3501 5114
rect 3482 5104 3486 5108
rect 3545 5084 3549 5161
rect 3565 5084 3569 5161
rect 3602 5116 3606 5161
rect 3624 5139 3628 5196
rect 3646 5193 3650 5236
rect 3730 5193 3734 5236
rect 3646 5181 3653 5193
rect 3727 5181 3734 5193
rect 3626 5127 3635 5139
rect 3602 5109 3615 5116
rect 3611 5104 3615 5109
rect 3631 5104 3635 5127
rect 3651 5104 3655 5181
rect 3725 5104 3729 5181
rect 3752 5139 3756 5196
rect 3760 5192 3764 5196
rect 3760 5184 3778 5192
rect 3774 5173 3778 5184
rect 3811 5173 3815 5196
rect 3806 5161 3815 5173
rect 3819 5173 3823 5196
rect 3819 5161 3834 5173
rect 3745 5127 3754 5139
rect 3745 5104 3749 5127
rect 3774 5116 3778 5161
rect 3765 5109 3778 5116
rect 3765 5104 3769 5109
rect 3811 5084 3815 5161
rect 3831 5084 3835 5161
rect 3891 5159 3895 5236
rect 3886 5147 3895 5159
rect 3889 5131 3895 5147
rect 3911 5159 3915 5236
rect 3985 5159 3989 5236
rect 3911 5147 3914 5159
rect 3986 5147 3989 5159
rect 3911 5131 3917 5147
rect 3889 5124 3897 5131
rect 3893 5104 3897 5124
rect 3903 5124 3917 5131
rect 3983 5131 3989 5147
rect 4005 5159 4009 5236
rect 4056 5192 4060 5196
rect 4042 5184 4060 5192
rect 4042 5173 4046 5184
rect 4005 5147 4014 5159
rect 4005 5131 4011 5147
rect 3983 5124 3997 5131
rect 3903 5104 3907 5124
rect 3993 5104 3997 5124
rect 4003 5124 4011 5131
rect 4003 5104 4007 5124
rect 4042 5116 4046 5161
rect 4064 5139 4068 5196
rect 4086 5193 4090 5236
rect 4086 5181 4093 5193
rect 4066 5127 4075 5139
rect 4042 5109 4055 5116
rect 4051 5104 4055 5109
rect 4071 5104 4075 5127
rect 4091 5104 4095 5181
rect 4165 5159 4169 5236
rect 4166 5147 4169 5159
rect 4163 5131 4169 5147
rect 4185 5159 4189 5236
rect 4185 5147 4194 5159
rect 4185 5131 4191 5147
rect 4163 5124 4177 5131
rect 4173 5104 4177 5124
rect 4183 5124 4191 5131
rect 4183 5104 4187 5124
rect 4241 5122 4245 5196
rect 4263 5159 4267 5236
rect 4285 5173 4289 5236
rect 4285 5161 4294 5173
rect 4266 5147 4279 5159
rect 4241 5110 4253 5122
rect 4255 5104 4259 5110
rect 4275 5104 4279 5147
rect 4285 5104 4289 5161
rect 4345 5159 4349 5236
rect 4346 5147 4349 5159
rect 4343 5131 4349 5147
rect 4365 5159 4369 5236
rect 4430 5193 4434 5236
rect 4427 5181 4434 5193
rect 4365 5147 4374 5159
rect 4365 5131 4371 5147
rect 4343 5124 4357 5131
rect 4353 5104 4357 5124
rect 4363 5124 4371 5131
rect 4363 5104 4367 5124
rect 4425 5104 4429 5181
rect 4452 5139 4456 5196
rect 4460 5192 4464 5196
rect 4530 5193 4534 5236
rect 4460 5184 4478 5192
rect 4474 5173 4478 5184
rect 4527 5181 4534 5193
rect 4445 5127 4454 5139
rect 4445 5104 4449 5127
rect 4474 5116 4478 5161
rect 4465 5109 4478 5116
rect 4465 5104 4469 5109
rect 4525 5104 4529 5181
rect 4552 5139 4556 5196
rect 4560 5192 4564 5196
rect 4560 5184 4578 5192
rect 4574 5173 4578 5184
rect 4545 5127 4554 5139
rect 4545 5104 4549 5127
rect 4574 5116 4578 5161
rect 4611 5159 4615 5236
rect 4606 5147 4615 5159
rect 4609 5131 4615 5147
rect 4631 5159 4635 5236
rect 4691 5159 4695 5236
rect 4631 5147 4634 5159
rect 4686 5147 4695 5159
rect 4631 5131 4637 5147
rect 4609 5124 4617 5131
rect 4565 5109 4578 5116
rect 4565 5104 4569 5109
rect 4613 5104 4617 5124
rect 4623 5124 4637 5131
rect 4689 5131 4695 5147
rect 4711 5159 4715 5236
rect 4711 5147 4714 5159
rect 4771 5153 4775 5236
rect 4845 5193 4849 5236
rect 4865 5224 4869 5236
rect 4885 5228 4889 5236
rect 4885 5224 4900 5228
rect 4865 5220 4880 5224
rect 4874 5213 4880 5220
rect 4845 5181 4853 5193
rect 4865 5181 4872 5193
rect 4711 5131 4717 5147
rect 4766 5141 4775 5153
rect 4689 5124 4697 5131
rect 4623 5104 4627 5124
rect 4693 5104 4697 5124
rect 4703 5124 4717 5131
rect 4703 5104 4707 5124
rect 4771 5084 4775 5141
rect 4868 5124 4872 5181
rect 4876 5124 4880 5201
rect 4894 5193 4900 5224
rect 4884 5181 4894 5193
rect 4936 5192 4940 5196
rect 4922 5184 4940 5192
rect 4884 5124 4888 5181
rect 4922 5173 4926 5184
rect 4922 5116 4926 5161
rect 4944 5139 4948 5196
rect 4966 5193 4970 5236
rect 4966 5181 4973 5193
rect 4946 5127 4955 5139
rect 4922 5109 4935 5116
rect 4931 5104 4935 5109
rect 4951 5104 4955 5127
rect 4971 5104 4975 5181
rect 5031 5139 5035 5196
rect 5091 5159 5095 5236
rect 5086 5147 5095 5159
rect 5026 5127 5035 5139
rect 5031 5104 5035 5127
rect 5089 5131 5095 5147
rect 5111 5159 5115 5236
rect 5171 5192 5175 5196
rect 5191 5192 5195 5196
rect 5171 5188 5195 5192
rect 5111 5147 5114 5159
rect 5111 5131 5117 5147
rect 5171 5139 5175 5188
rect 5251 5159 5255 5236
rect 5246 5147 5255 5159
rect 5089 5124 5097 5131
rect 5093 5104 5097 5124
rect 5103 5124 5117 5131
rect 5166 5127 5175 5139
rect 5103 5104 5107 5124
rect 5171 5112 5175 5127
rect 5249 5131 5255 5147
rect 5271 5159 5275 5236
rect 5336 5192 5340 5196
rect 5322 5184 5340 5192
rect 5322 5173 5326 5184
rect 5271 5147 5274 5159
rect 5271 5131 5277 5147
rect 5249 5124 5257 5131
rect 5171 5108 5195 5112
rect 5171 5104 5175 5108
rect 5191 5104 5195 5108
rect 5253 5104 5257 5124
rect 5263 5124 5277 5131
rect 5263 5104 5267 5124
rect 5322 5116 5326 5161
rect 5344 5139 5348 5196
rect 5366 5193 5370 5236
rect 5431 5228 5435 5236
rect 5420 5224 5435 5228
rect 5451 5224 5455 5236
rect 5420 5193 5426 5224
rect 5440 5220 5455 5224
rect 5440 5213 5446 5220
rect 5366 5181 5373 5193
rect 5426 5181 5436 5193
rect 5346 5127 5355 5139
rect 5322 5109 5335 5116
rect 5331 5104 5335 5109
rect 5351 5104 5355 5127
rect 5371 5104 5375 5181
rect 5432 5124 5436 5181
rect 5440 5124 5444 5201
rect 5471 5193 5475 5236
rect 5531 5228 5535 5236
rect 5520 5224 5535 5228
rect 5551 5224 5555 5236
rect 5520 5193 5526 5224
rect 5540 5220 5555 5224
rect 5540 5213 5546 5220
rect 5448 5181 5455 5193
rect 5467 5181 5475 5193
rect 5526 5181 5536 5193
rect 5448 5124 5452 5181
rect 5532 5124 5536 5181
rect 5540 5124 5544 5201
rect 5571 5193 5575 5236
rect 5548 5181 5555 5193
rect 5567 5181 5575 5193
rect 5548 5124 5552 5181
rect 5631 5153 5635 5236
rect 5691 5228 5695 5236
rect 5680 5224 5695 5228
rect 5711 5224 5715 5236
rect 5680 5193 5686 5224
rect 5700 5220 5715 5224
rect 5700 5213 5706 5220
rect 5686 5181 5696 5193
rect 5626 5141 5635 5153
rect 5631 5084 5635 5141
rect 5692 5124 5696 5181
rect 5700 5124 5704 5201
rect 5731 5193 5735 5236
rect 5708 5181 5715 5193
rect 5727 5181 5735 5193
rect 5796 5192 5800 5196
rect 5782 5184 5800 5192
rect 5708 5124 5712 5181
rect 5782 5173 5786 5184
rect 5782 5116 5786 5161
rect 5804 5139 5808 5196
rect 5826 5193 5830 5236
rect 5826 5181 5833 5193
rect 5806 5127 5815 5139
rect 5782 5109 5795 5116
rect 5791 5104 5795 5109
rect 5811 5104 5815 5127
rect 5831 5104 5835 5181
rect 5905 5159 5909 5236
rect 5906 5147 5909 5159
rect 5903 5131 5909 5147
rect 5925 5159 5929 5236
rect 5971 5228 5975 5236
rect 5960 5224 5975 5228
rect 5991 5224 5995 5236
rect 5960 5193 5966 5224
rect 5980 5220 5995 5224
rect 5980 5213 5986 5220
rect 5966 5181 5976 5193
rect 5925 5147 5934 5159
rect 5925 5131 5931 5147
rect 5903 5124 5917 5131
rect 5913 5104 5917 5124
rect 5923 5124 5931 5131
rect 5972 5124 5976 5181
rect 5980 5124 5984 5201
rect 6011 5193 6015 5236
rect 5988 5181 5995 5193
rect 6007 5181 6015 5193
rect 5988 5124 5992 5181
rect 6071 5159 6075 5236
rect 6066 5147 6075 5159
rect 6069 5131 6075 5147
rect 6091 5159 6095 5236
rect 6091 5147 6094 5159
rect 6091 5131 6097 5147
rect 6069 5124 6077 5131
rect 5923 5104 5927 5124
rect 6073 5104 6077 5124
rect 6083 5124 6097 5131
rect 6165 5139 6169 5196
rect 6185 5182 6189 5196
rect 6205 5182 6209 5196
rect 6185 5176 6200 5182
rect 6205 5176 6221 5182
rect 6194 5153 6200 5176
rect 6165 5127 6174 5139
rect 6083 5104 6087 5124
rect 6172 5084 6176 5127
rect 6194 5104 6198 5141
rect 6214 5139 6221 5176
rect 6265 5153 6269 5236
rect 6325 5193 6329 5236
rect 6345 5224 6349 5236
rect 6365 5228 6369 5236
rect 6365 5224 6380 5228
rect 6345 5220 6360 5224
rect 6354 5213 6360 5220
rect 6325 5181 6333 5193
rect 6345 5181 6352 5193
rect 6265 5141 6274 5153
rect 6214 5114 6221 5127
rect 6202 5108 6221 5114
rect 6202 5104 6206 5108
rect 6265 5084 6269 5141
rect 6348 5124 6352 5181
rect 6356 5124 6360 5201
rect 6374 5193 6380 5224
rect 6425 5193 6429 5236
rect 6445 5224 6449 5236
rect 6465 5228 6469 5236
rect 6465 5224 6480 5228
rect 6445 5220 6460 5224
rect 6454 5213 6460 5220
rect 6364 5181 6374 5193
rect 6425 5181 6433 5193
rect 6445 5181 6452 5193
rect 6364 5124 6368 5181
rect 6448 5124 6452 5181
rect 6456 5124 6460 5201
rect 6474 5193 6480 5224
rect 6464 5181 6474 5193
rect 6464 5124 6468 5181
rect 6511 5153 6515 5236
rect 6585 5193 6589 5236
rect 6605 5224 6609 5236
rect 6625 5228 6629 5236
rect 6625 5224 6640 5228
rect 6605 5220 6620 5224
rect 6614 5213 6620 5220
rect 6585 5181 6593 5193
rect 6605 5181 6612 5193
rect 6506 5141 6515 5153
rect 6511 5084 6515 5141
rect 6608 5124 6612 5181
rect 6616 5124 6620 5201
rect 6634 5193 6640 5224
rect 6624 5181 6634 5193
rect 6624 5124 6628 5181
rect 6671 5159 6675 5236
rect 6666 5147 6675 5159
rect 6669 5131 6675 5147
rect 6691 5159 6695 5236
rect 6691 5147 6694 5159
rect 6691 5131 6697 5147
rect 6669 5124 6677 5131
rect 6673 5104 6677 5124
rect 6683 5124 6697 5131
rect 6683 5104 6687 5124
rect 43 5060 47 5064
rect 65 5060 69 5064
rect 111 5060 115 5064
rect 133 5060 137 5064
rect 143 5060 147 5064
rect 163 5060 167 5064
rect 171 5060 175 5064
rect 217 5060 221 5064
rect 239 5060 243 5064
rect 249 5060 253 5064
rect 271 5060 275 5064
rect 281 5060 285 5064
rect 301 5060 305 5064
rect 353 5060 357 5064
rect 363 5060 367 5064
rect 452 5060 456 5064
rect 474 5060 478 5064
rect 482 5060 486 5064
rect 553 5060 557 5064
rect 563 5060 567 5064
rect 615 5060 619 5064
rect 635 5060 639 5064
rect 645 5060 649 5064
rect 667 5060 671 5064
rect 677 5060 681 5064
rect 699 5060 703 5064
rect 745 5060 749 5064
rect 753 5060 757 5064
rect 773 5060 777 5064
rect 783 5060 787 5064
rect 805 5060 809 5064
rect 853 5060 857 5064
rect 863 5060 867 5064
rect 945 5060 949 5064
rect 965 5060 969 5064
rect 985 5060 989 5064
rect 1045 5060 1049 5064
rect 1065 5060 1069 5064
rect 1085 5060 1089 5064
rect 1155 5060 1159 5064
rect 1175 5060 1179 5064
rect 1185 5060 1189 5064
rect 1231 5060 1235 5064
rect 1253 5060 1257 5064
rect 1263 5060 1267 5064
rect 1283 5060 1287 5064
rect 1291 5060 1295 5064
rect 1337 5060 1341 5064
rect 1359 5060 1363 5064
rect 1369 5060 1373 5064
rect 1391 5060 1395 5064
rect 1401 5060 1405 5064
rect 1421 5060 1425 5064
rect 1493 5060 1497 5064
rect 1503 5060 1507 5064
rect 1553 5060 1557 5064
rect 1563 5060 1567 5064
rect 1631 5060 1635 5064
rect 1653 5060 1657 5064
rect 1663 5060 1667 5064
rect 1683 5060 1687 5064
rect 1691 5060 1695 5064
rect 1737 5060 1741 5064
rect 1759 5060 1763 5064
rect 1769 5060 1773 5064
rect 1791 5060 1795 5064
rect 1801 5060 1805 5064
rect 1821 5060 1825 5064
rect 1906 5060 1910 5064
rect 1914 5060 1918 5064
rect 1934 5060 1938 5064
rect 1942 5060 1946 5064
rect 1991 5060 1995 5064
rect 2075 5060 2079 5064
rect 2095 5060 2099 5064
rect 2105 5060 2109 5064
rect 2153 5060 2157 5064
rect 2163 5060 2167 5064
rect 2245 5060 2249 5064
rect 2265 5060 2269 5064
rect 2285 5060 2289 5064
rect 2353 5060 2357 5064
rect 2363 5060 2367 5064
rect 2448 5060 2452 5064
rect 2456 5060 2460 5064
rect 2464 5060 2468 5064
rect 2525 5060 2529 5064
rect 2545 5060 2549 5064
rect 2591 5060 2595 5064
rect 2675 5060 2679 5064
rect 2695 5060 2699 5064
rect 2705 5060 2709 5064
rect 2751 5060 2755 5064
rect 2771 5060 2775 5064
rect 2853 5060 2857 5064
rect 2863 5060 2867 5064
rect 2933 5060 2937 5064
rect 2943 5060 2947 5064
rect 2991 5060 2995 5064
rect 3011 5060 3015 5064
rect 3031 5060 3035 5064
rect 3115 5060 3119 5064
rect 3135 5060 3139 5064
rect 3145 5060 3149 5064
rect 3193 5060 3197 5064
rect 3203 5060 3207 5064
rect 3308 5060 3312 5064
rect 3316 5060 3320 5064
rect 3324 5060 3328 5064
rect 3385 5060 3389 5064
rect 3452 5060 3456 5064
rect 3474 5060 3478 5064
rect 3482 5060 3486 5064
rect 3545 5060 3549 5064
rect 3565 5060 3569 5064
rect 3611 5060 3615 5064
rect 3631 5060 3635 5064
rect 3651 5060 3655 5064
rect 3725 5060 3729 5064
rect 3745 5060 3749 5064
rect 3765 5060 3769 5064
rect 3811 5060 3815 5064
rect 3831 5060 3835 5064
rect 3893 5060 3897 5064
rect 3903 5060 3907 5064
rect 3993 5060 3997 5064
rect 4003 5060 4007 5064
rect 4051 5060 4055 5064
rect 4071 5060 4075 5064
rect 4091 5060 4095 5064
rect 4173 5060 4177 5064
rect 4183 5060 4187 5064
rect 4255 5060 4259 5064
rect 4275 5060 4279 5064
rect 4285 5060 4289 5064
rect 4353 5060 4357 5064
rect 4363 5060 4367 5064
rect 4425 5060 4429 5064
rect 4445 5060 4449 5064
rect 4465 5060 4469 5064
rect 4525 5060 4529 5064
rect 4545 5060 4549 5064
rect 4565 5060 4569 5064
rect 4613 5060 4617 5064
rect 4623 5060 4627 5064
rect 4693 5060 4697 5064
rect 4703 5060 4707 5064
rect 4771 5060 4775 5064
rect 4868 5060 4872 5064
rect 4876 5060 4880 5064
rect 4884 5060 4888 5064
rect 4931 5060 4935 5064
rect 4951 5060 4955 5064
rect 4971 5060 4975 5064
rect 5031 5060 5035 5064
rect 5093 5060 5097 5064
rect 5103 5060 5107 5064
rect 5171 5060 5175 5064
rect 5191 5060 5195 5064
rect 5253 5060 5257 5064
rect 5263 5060 5267 5064
rect 5331 5060 5335 5064
rect 5351 5060 5355 5064
rect 5371 5060 5375 5064
rect 5432 5060 5436 5064
rect 5440 5060 5444 5064
rect 5448 5060 5452 5064
rect 5532 5060 5536 5064
rect 5540 5060 5544 5064
rect 5548 5060 5552 5064
rect 5631 5060 5635 5064
rect 5692 5060 5696 5064
rect 5700 5060 5704 5064
rect 5708 5060 5712 5064
rect 5791 5060 5795 5064
rect 5811 5060 5815 5064
rect 5831 5060 5835 5064
rect 5913 5060 5917 5064
rect 5923 5060 5927 5064
rect 5972 5060 5976 5064
rect 5980 5060 5984 5064
rect 5988 5060 5992 5064
rect 6073 5060 6077 5064
rect 6083 5060 6087 5064
rect 6172 5060 6176 5064
rect 6194 5060 6198 5064
rect 6202 5060 6206 5064
rect 6265 5060 6269 5064
rect 6348 5060 6352 5064
rect 6356 5060 6360 5064
rect 6364 5060 6368 5064
rect 6448 5060 6452 5064
rect 6456 5060 6460 5064
rect 6464 5060 6468 5064
rect 6511 5060 6515 5064
rect 6608 5060 6612 5064
rect 6616 5060 6620 5064
rect 6624 5060 6628 5064
rect 6673 5060 6677 5064
rect 6683 5060 6687 5064
rect 43 5036 47 5040
rect 65 5036 69 5040
rect 123 5036 127 5040
rect 145 5036 149 5040
rect 213 5036 217 5040
rect 223 5036 227 5040
rect 271 5036 275 5040
rect 293 5036 297 5040
rect 303 5036 307 5040
rect 323 5036 327 5040
rect 331 5036 335 5040
rect 377 5036 381 5040
rect 399 5036 403 5040
rect 409 5036 413 5040
rect 431 5036 435 5040
rect 441 5036 445 5040
rect 461 5036 465 5040
rect 532 5036 536 5040
rect 554 5036 558 5040
rect 562 5036 566 5040
rect 633 5036 637 5040
rect 643 5036 647 5040
rect 693 5036 697 5040
rect 703 5036 707 5040
rect 793 5036 797 5040
rect 803 5036 807 5040
rect 851 5036 855 5040
rect 873 5036 877 5040
rect 883 5036 887 5040
rect 903 5036 907 5040
rect 911 5036 915 5040
rect 957 5036 961 5040
rect 979 5036 983 5040
rect 989 5036 993 5040
rect 1011 5036 1015 5040
rect 1021 5036 1025 5040
rect 1041 5036 1045 5040
rect 1103 5036 1107 5040
rect 1125 5036 1129 5040
rect 1192 5036 1196 5040
rect 1214 5036 1218 5040
rect 1222 5036 1226 5040
rect 1293 5036 1297 5040
rect 1303 5036 1307 5040
rect 1363 5036 1367 5040
rect 1385 5036 1389 5040
rect 1433 5036 1437 5040
rect 1443 5036 1447 5040
rect 1533 5036 1537 5040
rect 1543 5036 1547 5040
rect 1605 5036 1609 5040
rect 1625 5036 1629 5040
rect 1645 5036 1649 5040
rect 1713 5036 1717 5040
rect 1723 5036 1727 5040
rect 1785 5036 1789 5040
rect 1805 5036 1809 5040
rect 1825 5036 1829 5040
rect 1873 5036 1877 5040
rect 1883 5036 1887 5040
rect 1965 5036 1969 5040
rect 1985 5036 1989 5040
rect 2005 5036 2009 5040
rect 2065 5036 2069 5040
rect 2085 5036 2089 5040
rect 2105 5036 2109 5040
rect 2175 5036 2179 5040
rect 2195 5036 2199 5040
rect 2205 5036 2209 5040
rect 2251 5036 2255 5040
rect 2325 5036 2329 5040
rect 2345 5036 2349 5040
rect 2405 5036 2409 5040
rect 2425 5036 2429 5040
rect 2445 5036 2449 5040
rect 2513 5036 2517 5040
rect 2523 5036 2527 5040
rect 2585 5036 2589 5040
rect 2605 5036 2609 5040
rect 2625 5036 2629 5040
rect 2685 5036 2689 5040
rect 2705 5036 2709 5040
rect 2725 5036 2729 5040
rect 2785 5036 2789 5040
rect 2831 5036 2835 5040
rect 2851 5036 2855 5040
rect 2871 5036 2875 5040
rect 2945 5036 2949 5040
rect 2965 5036 2969 5040
rect 2985 5036 2989 5040
rect 3045 5036 3049 5040
rect 3065 5036 3069 5040
rect 3085 5036 3089 5040
rect 3145 5036 3149 5040
rect 3165 5036 3169 5040
rect 3225 5036 3229 5040
rect 3293 5036 3297 5040
rect 3303 5036 3307 5040
rect 3365 5036 3369 5040
rect 3385 5036 3389 5040
rect 3405 5036 3409 5040
rect 3455 5036 3459 5040
rect 3475 5036 3479 5040
rect 3485 5036 3489 5040
rect 3507 5036 3511 5040
rect 3517 5036 3521 5040
rect 3539 5036 3543 5040
rect 3585 5036 3589 5040
rect 3593 5036 3597 5040
rect 3613 5036 3617 5040
rect 3623 5036 3627 5040
rect 3645 5036 3649 5040
rect 3691 5036 3695 5040
rect 3711 5036 3715 5040
rect 3731 5036 3735 5040
rect 3812 5036 3816 5040
rect 3834 5036 3838 5040
rect 3842 5036 3846 5040
rect 3928 5036 3932 5040
rect 3936 5036 3940 5040
rect 3944 5036 3948 5040
rect 4012 5036 4016 5040
rect 4034 5036 4038 5040
rect 4042 5036 4046 5040
rect 4105 5036 4109 5040
rect 4175 5036 4179 5040
rect 4195 5036 4199 5040
rect 4205 5036 4209 5040
rect 4273 5036 4277 5040
rect 4283 5036 4287 5040
rect 4331 5036 4335 5040
rect 4341 5036 4345 5040
rect 4361 5036 4365 5040
rect 4445 5036 4449 5040
rect 4465 5036 4469 5040
rect 4485 5036 4489 5040
rect 4532 5036 4536 5040
rect 4540 5036 4544 5040
rect 4548 5036 4552 5040
rect 4631 5036 4635 5040
rect 4651 5036 4655 5040
rect 4671 5036 4675 5040
rect 4753 5036 4757 5040
rect 4763 5036 4767 5040
rect 4835 5036 4839 5040
rect 4855 5036 4859 5040
rect 4865 5036 4869 5040
rect 4933 5036 4937 5040
rect 4943 5036 4947 5040
rect 4993 5036 4997 5040
rect 5003 5036 5007 5040
rect 5071 5036 5075 5040
rect 5081 5036 5085 5040
rect 5101 5036 5105 5040
rect 5193 5036 5197 5040
rect 5203 5036 5207 5040
rect 5275 5036 5279 5040
rect 5295 5036 5299 5040
rect 5305 5036 5309 5040
rect 5351 5036 5355 5040
rect 5361 5036 5365 5040
rect 5381 5036 5385 5040
rect 5486 5036 5490 5040
rect 5494 5036 5498 5040
rect 5514 5036 5518 5040
rect 5522 5036 5526 5040
rect 5593 5036 5597 5040
rect 5603 5036 5607 5040
rect 5652 5036 5656 5040
rect 5660 5036 5664 5040
rect 5668 5036 5672 5040
rect 5772 5036 5776 5040
rect 5794 5036 5798 5040
rect 5802 5036 5806 5040
rect 5888 5036 5892 5040
rect 5896 5036 5900 5040
rect 5904 5036 5908 5040
rect 5973 5036 5977 5040
rect 5983 5036 5987 5040
rect 6034 5036 6038 5040
rect 6042 5036 6046 5040
rect 6062 5036 6066 5040
rect 6070 5036 6074 5040
rect 6188 5036 6192 5040
rect 6196 5036 6200 5040
rect 6204 5036 6208 5040
rect 6251 5036 6255 5040
rect 6271 5036 6275 5040
rect 6291 5036 6295 5040
rect 6388 5036 6392 5040
rect 6396 5036 6400 5040
rect 6404 5036 6408 5040
rect 6488 5036 6492 5040
rect 6496 5036 6500 5040
rect 6504 5036 6508 5040
rect 6553 5036 6557 5040
rect 6563 5036 6567 5040
rect 6645 5036 6649 5040
rect 43 4990 47 4996
rect 43 4978 45 4990
rect 65 4939 69 5016
rect 123 4990 127 4996
rect 123 4978 125 4990
rect 145 4939 149 5016
rect 213 4976 217 4996
rect 203 4969 217 4976
rect 223 4976 227 4996
rect 223 4969 231 4976
rect 203 4953 209 4969
rect 206 4941 209 4953
rect 65 4927 74 4939
rect 145 4927 154 4939
rect 43 4910 45 4922
rect 43 4904 47 4910
rect 65 4864 69 4927
rect 123 4910 125 4922
rect 123 4904 127 4910
rect 145 4864 149 4927
rect 205 4864 209 4941
rect 225 4953 231 4969
rect 225 4941 234 4953
rect 225 4864 229 4941
rect 271 4928 275 4996
rect 293 4967 297 5016
rect 303 4995 307 5016
rect 323 5004 327 5016
rect 331 5012 335 5016
rect 331 5008 365 5012
rect 323 5000 353 5004
rect 323 4999 341 5000
rect 303 4991 327 4995
rect 271 4916 273 4928
rect 271 4904 275 4916
rect 293 4909 297 4955
rect 289 4903 297 4909
rect 289 4874 293 4903
rect 321 4896 327 4991
rect 289 4867 297 4874
rect 293 4844 297 4867
rect 301 4844 305 4884
rect 321 4864 325 4896
rect 361 4882 365 5008
rect 377 4902 381 5016
rect 399 5004 403 5016
rect 401 4992 403 5004
rect 409 5004 413 5016
rect 409 4992 411 5004
rect 329 4870 353 4872
rect 329 4868 365 4870
rect 329 4864 333 4868
rect 375 4864 379 4890
rect 393 4882 397 4992
rect 431 4984 435 5016
rect 402 4980 435 4984
rect 402 4916 406 4980
rect 422 4931 426 4960
rect 441 4958 445 5016
rect 461 4959 465 4996
rect 532 4973 536 5016
rect 525 4961 534 4973
rect 422 4923 431 4931
rect 402 4904 405 4916
rect 395 4864 399 4870
rect 407 4864 411 4904
rect 427 4864 431 4923
rect 441 4864 445 4946
rect 461 4904 465 4947
rect 525 4904 529 4961
rect 554 4959 558 4996
rect 562 4992 566 4996
rect 562 4986 581 4992
rect 574 4973 581 4986
rect 633 4976 637 4996
rect 623 4969 637 4976
rect 643 4976 647 4996
rect 693 4976 697 4996
rect 643 4969 651 4976
rect 554 4924 560 4947
rect 574 4924 581 4961
rect 623 4953 629 4969
rect 626 4941 629 4953
rect 545 4918 560 4924
rect 565 4918 581 4924
rect 545 4904 549 4918
rect 565 4904 569 4918
rect 625 4864 629 4941
rect 645 4953 651 4969
rect 689 4969 697 4976
rect 703 4976 707 4996
rect 793 4976 797 4996
rect 703 4969 717 4976
rect 689 4953 695 4969
rect 645 4941 654 4953
rect 686 4941 695 4953
rect 645 4864 649 4941
rect 691 4864 695 4941
rect 711 4953 717 4969
rect 783 4969 797 4976
rect 803 4976 807 4996
rect 803 4969 811 4976
rect 783 4953 789 4969
rect 711 4941 714 4953
rect 786 4941 789 4953
rect 711 4864 715 4941
rect 785 4864 789 4941
rect 805 4953 811 4969
rect 805 4941 814 4953
rect 805 4864 809 4941
rect 851 4928 855 4996
rect 873 4967 877 5016
rect 883 4995 887 5016
rect 903 5004 907 5016
rect 911 5012 915 5016
rect 911 5008 945 5012
rect 903 5000 933 5004
rect 903 4999 921 5000
rect 883 4991 907 4995
rect 851 4916 853 4928
rect 851 4904 855 4916
rect 873 4909 877 4955
rect 869 4903 877 4909
rect 869 4874 873 4903
rect 901 4896 907 4991
rect 869 4867 877 4874
rect 873 4844 877 4867
rect 881 4844 885 4884
rect 901 4864 905 4896
rect 941 4882 945 5008
rect 957 4902 961 5016
rect 979 5004 983 5016
rect 981 4992 983 5004
rect 989 5004 993 5016
rect 989 4992 991 5004
rect 909 4870 933 4872
rect 909 4868 945 4870
rect 909 4864 913 4868
rect 955 4864 959 4890
rect 973 4882 977 4992
rect 1011 4984 1015 5016
rect 982 4980 1015 4984
rect 982 4916 986 4980
rect 1002 4931 1006 4960
rect 1021 4958 1025 5016
rect 1041 4959 1045 4996
rect 1103 4990 1107 4996
rect 1103 4978 1105 4990
rect 1002 4923 1011 4931
rect 982 4904 985 4916
rect 975 4864 979 4870
rect 987 4864 991 4904
rect 1007 4864 1011 4923
rect 1021 4864 1025 4946
rect 1041 4904 1045 4947
rect 1125 4939 1129 5016
rect 1192 4973 1196 5016
rect 1185 4961 1194 4973
rect 1125 4927 1134 4939
rect 1103 4910 1105 4922
rect 1103 4904 1107 4910
rect 1125 4864 1129 4927
rect 1185 4904 1189 4961
rect 1214 4959 1218 4996
rect 1222 4992 1226 4996
rect 1222 4986 1241 4992
rect 1234 4973 1241 4986
rect 1293 4976 1297 4996
rect 1283 4969 1297 4976
rect 1303 4976 1307 4996
rect 1363 4990 1367 4996
rect 1363 4978 1365 4990
rect 1303 4969 1311 4976
rect 1214 4924 1220 4947
rect 1234 4924 1241 4961
rect 1283 4953 1289 4969
rect 1286 4941 1289 4953
rect 1205 4918 1220 4924
rect 1225 4918 1241 4924
rect 1205 4904 1209 4918
rect 1225 4904 1229 4918
rect 1285 4864 1289 4941
rect 1305 4953 1311 4969
rect 1305 4941 1314 4953
rect 1305 4864 1309 4941
rect 1385 4939 1389 5016
rect 1433 4976 1437 4996
rect 1429 4969 1437 4976
rect 1443 4976 1447 4996
rect 1533 4976 1537 4996
rect 1443 4969 1457 4976
rect 1429 4953 1435 4969
rect 1426 4941 1435 4953
rect 1385 4927 1394 4939
rect 1363 4910 1365 4922
rect 1363 4904 1367 4910
rect 1385 4864 1389 4927
rect 1431 4864 1435 4941
rect 1451 4953 1457 4969
rect 1523 4969 1537 4976
rect 1543 4976 1547 4996
rect 1543 4969 1551 4976
rect 1523 4953 1529 4969
rect 1451 4941 1454 4953
rect 1526 4941 1529 4953
rect 1451 4864 1455 4941
rect 1525 4864 1529 4941
rect 1545 4953 1551 4969
rect 1545 4941 1554 4953
rect 1545 4864 1549 4941
rect 1605 4919 1609 4996
rect 1625 4973 1629 4996
rect 1645 4991 1649 4996
rect 1645 4984 1658 4991
rect 1625 4961 1634 4973
rect 1607 4907 1614 4919
rect 1610 4864 1614 4907
rect 1632 4904 1636 4961
rect 1654 4939 1658 4984
rect 1713 4976 1717 4996
rect 1703 4969 1717 4976
rect 1723 4976 1727 4996
rect 1723 4969 1731 4976
rect 1703 4953 1709 4969
rect 1706 4941 1709 4953
rect 1654 4916 1658 4927
rect 1640 4908 1658 4916
rect 1640 4904 1644 4908
rect 1705 4864 1709 4941
rect 1725 4953 1731 4969
rect 1725 4941 1734 4953
rect 1725 4864 1729 4941
rect 1785 4919 1789 4996
rect 1805 4973 1809 4996
rect 1825 4991 1829 4996
rect 1825 4984 1838 4991
rect 1805 4961 1814 4973
rect 1787 4907 1794 4919
rect 1790 4864 1794 4907
rect 1812 4904 1816 4961
rect 1834 4939 1838 4984
rect 1873 4976 1877 4996
rect 1869 4969 1877 4976
rect 1883 4976 1887 4996
rect 1883 4969 1897 4976
rect 1869 4953 1875 4969
rect 1866 4941 1875 4953
rect 1834 4916 1838 4927
rect 1820 4908 1838 4916
rect 1820 4904 1824 4908
rect 1871 4864 1875 4941
rect 1891 4953 1897 4969
rect 1891 4941 1894 4953
rect 1891 4864 1895 4941
rect 1965 4919 1969 4996
rect 1985 4973 1989 4996
rect 2005 4991 2009 4996
rect 2005 4984 2018 4991
rect 1985 4961 1994 4973
rect 1967 4907 1974 4919
rect 1970 4864 1974 4907
rect 1992 4904 1996 4961
rect 2014 4939 2018 4984
rect 2014 4916 2018 4927
rect 2065 4919 2069 4996
rect 2085 4973 2089 4996
rect 2105 4991 2109 4996
rect 2105 4984 2118 4991
rect 2175 4990 2179 4996
rect 2085 4961 2094 4973
rect 2000 4908 2018 4916
rect 2000 4904 2004 4908
rect 2067 4907 2074 4919
rect 2070 4864 2074 4907
rect 2092 4904 2096 4961
rect 2114 4939 2118 4984
rect 2161 4978 2173 4990
rect 2114 4916 2118 4927
rect 2100 4908 2118 4916
rect 2100 4904 2104 4908
rect 2161 4904 2165 4978
rect 2195 4953 2199 4996
rect 2186 4941 2199 4953
rect 2183 4864 2187 4941
rect 2205 4939 2209 4996
rect 2251 4959 2255 5016
rect 2246 4947 2255 4959
rect 2205 4927 2214 4939
rect 2205 4864 2209 4927
rect 2251 4864 2255 4947
rect 2325 4939 2329 5016
rect 2345 4939 2349 5016
rect 2425 5009 2429 5016
rect 2445 5009 2449 5016
rect 2425 5003 2439 5009
rect 2445 5004 2458 5009
rect 2405 4988 2409 4996
rect 2405 4976 2415 4988
rect 2435 4939 2439 5003
rect 2454 4959 2458 5004
rect 2513 4976 2517 4996
rect 2503 4969 2517 4976
rect 2523 4976 2527 4996
rect 2523 4969 2531 4976
rect 2503 4953 2509 4969
rect 2326 4927 2341 4939
rect 2337 4904 2341 4927
rect 2345 4927 2354 4939
rect 2345 4904 2349 4927
rect 2415 4904 2419 4909
rect 2435 4904 2439 4927
rect 2454 4913 2458 4947
rect 2506 4941 2509 4953
rect 2445 4908 2458 4913
rect 2445 4904 2449 4908
rect 2505 4864 2509 4941
rect 2525 4953 2531 4969
rect 2525 4941 2534 4953
rect 2525 4864 2529 4941
rect 2585 4919 2589 4996
rect 2605 4973 2609 4996
rect 2625 4991 2629 4996
rect 2625 4984 2638 4991
rect 2605 4961 2614 4973
rect 2587 4907 2594 4919
rect 2590 4864 2594 4907
rect 2612 4904 2616 4961
rect 2634 4939 2638 4984
rect 2634 4916 2638 4927
rect 2685 4919 2689 4996
rect 2705 4973 2709 4996
rect 2725 4991 2729 4996
rect 2725 4984 2738 4991
rect 2705 4961 2714 4973
rect 2620 4908 2638 4916
rect 2620 4904 2624 4908
rect 2687 4907 2694 4919
rect 2690 4864 2694 4907
rect 2712 4904 2716 4961
rect 2734 4939 2738 4984
rect 2785 4959 2789 5016
rect 2831 4991 2835 4996
rect 2822 4984 2835 4991
rect 2785 4947 2794 4959
rect 2734 4916 2738 4927
rect 2720 4908 2738 4916
rect 2720 4904 2724 4908
rect 2785 4864 2789 4947
rect 2822 4939 2826 4984
rect 2851 4973 2855 4996
rect 2846 4961 2855 4973
rect 2822 4916 2826 4927
rect 2822 4908 2840 4916
rect 2836 4904 2840 4908
rect 2844 4904 2848 4961
rect 2871 4919 2875 4996
rect 2945 4919 2949 4996
rect 2965 4973 2969 4996
rect 2985 4991 2989 4996
rect 2985 4984 2998 4991
rect 2965 4961 2974 4973
rect 2866 4907 2873 4919
rect 2947 4907 2954 4919
rect 2866 4864 2870 4907
rect 2950 4864 2954 4907
rect 2972 4904 2976 4961
rect 2994 4939 2998 4984
rect 2994 4916 2998 4927
rect 3045 4919 3049 4996
rect 3065 4973 3069 4996
rect 3085 4991 3089 4996
rect 3085 4984 3098 4991
rect 3065 4961 3074 4973
rect 2980 4908 2998 4916
rect 2980 4904 2984 4908
rect 3047 4907 3054 4919
rect 3050 4864 3054 4907
rect 3072 4904 3076 4961
rect 3094 4939 3098 4984
rect 3145 4939 3149 5016
rect 3165 4939 3169 5016
rect 3225 4973 3229 4996
rect 3293 4976 3297 4996
rect 3225 4961 3234 4973
rect 3283 4969 3297 4976
rect 3303 4976 3307 4996
rect 3303 4969 3311 4976
rect 3146 4927 3161 4939
rect 3094 4916 3098 4927
rect 3080 4908 3098 4916
rect 3080 4904 3084 4908
rect 3157 4904 3161 4927
rect 3165 4927 3174 4939
rect 3165 4904 3169 4927
rect 3225 4904 3229 4961
rect 3283 4953 3289 4969
rect 3286 4941 3289 4953
rect 3285 4864 3289 4941
rect 3305 4953 3311 4969
rect 3305 4941 3314 4953
rect 3305 4864 3309 4941
rect 3365 4919 3369 4996
rect 3385 4973 3389 4996
rect 3405 4991 3409 4996
rect 3405 4984 3418 4991
rect 3385 4961 3394 4973
rect 3367 4907 3374 4919
rect 3370 4864 3374 4907
rect 3392 4904 3396 4961
rect 3414 4939 3418 4984
rect 3455 4959 3459 4996
rect 3475 4958 3479 5016
rect 3485 4984 3489 5016
rect 3507 5004 3511 5016
rect 3509 4992 3511 5004
rect 3517 5004 3521 5016
rect 3517 4992 3519 5004
rect 3485 4980 3518 4984
rect 3414 4916 3418 4927
rect 3400 4908 3418 4916
rect 3400 4904 3404 4908
rect 3455 4904 3459 4947
rect 3475 4864 3479 4946
rect 3494 4931 3498 4960
rect 3489 4923 3498 4931
rect 3489 4864 3493 4923
rect 3514 4916 3518 4980
rect 3515 4904 3518 4916
rect 3509 4864 3513 4904
rect 3523 4882 3527 4992
rect 3539 4902 3543 5016
rect 3585 5012 3589 5016
rect 3555 5008 3589 5012
rect 3521 4864 3525 4870
rect 3541 4864 3545 4890
rect 3555 4882 3559 5008
rect 3593 5004 3597 5016
rect 3567 5000 3597 5004
rect 3579 4999 3597 5000
rect 3613 4995 3617 5016
rect 3593 4991 3617 4995
rect 3593 4896 3599 4991
rect 3623 4967 3627 5016
rect 3623 4909 3627 4955
rect 3645 4928 3649 4996
rect 3691 4991 3695 4996
rect 3682 4984 3695 4991
rect 3682 4939 3686 4984
rect 3711 4973 3715 4996
rect 3706 4961 3715 4973
rect 3647 4916 3649 4928
rect 3623 4903 3631 4909
rect 3645 4904 3649 4916
rect 3682 4916 3686 4927
rect 3682 4908 3700 4916
rect 3696 4904 3700 4908
rect 3704 4904 3708 4961
rect 3731 4919 3735 4996
rect 3812 4973 3816 5016
rect 3805 4961 3814 4973
rect 3726 4907 3733 4919
rect 3567 4870 3591 4872
rect 3555 4868 3591 4870
rect 3587 4864 3591 4868
rect 3595 4864 3599 4896
rect 3615 4844 3619 4884
rect 3627 4874 3631 4903
rect 3623 4867 3631 4874
rect 3623 4844 3627 4867
rect 3726 4864 3730 4907
rect 3805 4904 3809 4961
rect 3834 4959 3838 4996
rect 3842 4992 3846 4996
rect 3842 4986 3861 4992
rect 3854 4973 3861 4986
rect 3834 4924 3840 4947
rect 3854 4924 3861 4961
rect 3825 4918 3840 4924
rect 3845 4918 3861 4924
rect 3928 4919 3932 4976
rect 3825 4904 3829 4918
rect 3845 4904 3849 4918
rect 3905 4907 3913 4919
rect 3925 4907 3932 4919
rect 3905 4864 3909 4907
rect 3936 4899 3940 4976
rect 3944 4919 3948 4976
rect 4012 4973 4016 5016
rect 4005 4961 4014 4973
rect 3944 4907 3954 4919
rect 3934 4880 3940 4887
rect 3925 4876 3940 4880
rect 3954 4876 3960 4907
rect 4005 4904 4009 4961
rect 4034 4959 4038 4996
rect 4042 4992 4046 4996
rect 4042 4986 4061 4992
rect 4054 4973 4061 4986
rect 4105 4973 4109 4996
rect 4175 4990 4179 4996
rect 4161 4978 4173 4990
rect 4105 4961 4114 4973
rect 4034 4924 4040 4947
rect 4054 4924 4061 4961
rect 4025 4918 4040 4924
rect 4045 4918 4061 4924
rect 4025 4904 4029 4918
rect 4045 4904 4049 4918
rect 4105 4904 4109 4961
rect 4161 4904 4165 4978
rect 4195 4953 4199 4996
rect 4186 4941 4199 4953
rect 3925 4864 3929 4876
rect 3945 4872 3960 4876
rect 3945 4864 3949 4872
rect 4183 4864 4187 4941
rect 4205 4939 4209 4996
rect 4273 4976 4277 4996
rect 4263 4969 4277 4976
rect 4283 4976 4287 4996
rect 4283 4969 4291 4976
rect 4263 4953 4269 4969
rect 4266 4941 4269 4953
rect 4205 4927 4214 4939
rect 4205 4864 4209 4927
rect 4265 4864 4269 4941
rect 4285 4953 4291 4969
rect 4285 4941 4294 4953
rect 4285 4864 4289 4941
rect 4331 4939 4335 4996
rect 4341 4953 4345 4996
rect 4361 4990 4365 4996
rect 4367 4978 4379 4990
rect 4341 4941 4354 4953
rect 4326 4927 4335 4939
rect 4331 4864 4335 4927
rect 4353 4864 4357 4941
rect 4375 4904 4379 4978
rect 4445 4919 4449 4996
rect 4465 4973 4469 4996
rect 4485 4991 4489 4996
rect 4485 4984 4498 4991
rect 4465 4961 4474 4973
rect 4447 4907 4454 4919
rect 4450 4864 4454 4907
rect 4472 4904 4476 4961
rect 4494 4939 4498 4984
rect 4631 4991 4635 4996
rect 4622 4984 4635 4991
rect 4494 4916 4498 4927
rect 4532 4919 4536 4976
rect 4480 4908 4498 4916
rect 4480 4904 4484 4908
rect 4526 4907 4536 4919
rect 4520 4876 4526 4907
rect 4540 4899 4544 4976
rect 4548 4919 4552 4976
rect 4622 4939 4626 4984
rect 4651 4973 4655 4996
rect 4646 4961 4655 4973
rect 4548 4907 4555 4919
rect 4567 4907 4575 4919
rect 4622 4916 4626 4927
rect 4622 4908 4640 4916
rect 4540 4880 4546 4887
rect 4540 4876 4555 4880
rect 4520 4872 4535 4876
rect 4531 4864 4535 4872
rect 4551 4864 4555 4876
rect 4571 4864 4575 4907
rect 4636 4904 4640 4908
rect 4644 4904 4648 4961
rect 4671 4919 4675 4996
rect 4753 4976 4757 4996
rect 4743 4969 4757 4976
rect 4763 4976 4767 4996
rect 4835 4990 4839 4996
rect 4821 4978 4833 4990
rect 4763 4969 4771 4976
rect 4743 4953 4749 4969
rect 4746 4941 4749 4953
rect 4666 4907 4673 4919
rect 4666 4864 4670 4907
rect 4745 4864 4749 4941
rect 4765 4953 4771 4969
rect 4765 4941 4774 4953
rect 4765 4864 4769 4941
rect 4821 4904 4825 4978
rect 4855 4953 4859 4996
rect 4846 4941 4859 4953
rect 4843 4864 4847 4941
rect 4865 4939 4869 4996
rect 4933 4976 4937 4996
rect 4923 4969 4937 4976
rect 4943 4976 4947 4996
rect 4993 4976 4997 4996
rect 4943 4969 4951 4976
rect 4923 4953 4929 4969
rect 4926 4941 4929 4953
rect 4865 4927 4874 4939
rect 4865 4864 4869 4927
rect 4925 4864 4929 4941
rect 4945 4953 4951 4969
rect 4989 4969 4997 4976
rect 5003 4976 5007 4996
rect 5003 4969 5017 4976
rect 4989 4953 4995 4969
rect 4945 4941 4954 4953
rect 4986 4941 4995 4953
rect 4945 4864 4949 4941
rect 4991 4864 4995 4941
rect 5011 4953 5017 4969
rect 5011 4941 5014 4953
rect 5011 4864 5015 4941
rect 5071 4939 5075 4996
rect 5081 4953 5085 4996
rect 5101 4990 5105 4996
rect 5107 4978 5119 4990
rect 5081 4941 5094 4953
rect 5066 4927 5075 4939
rect 5071 4864 5075 4927
rect 5093 4864 5097 4941
rect 5115 4904 5119 4978
rect 5193 4976 5197 4996
rect 5183 4969 5197 4976
rect 5203 4976 5207 4996
rect 5275 4990 5279 4996
rect 5261 4978 5273 4990
rect 5203 4969 5211 4976
rect 5183 4953 5189 4969
rect 5186 4941 5189 4953
rect 5185 4864 5189 4941
rect 5205 4953 5211 4969
rect 5205 4941 5214 4953
rect 5205 4864 5209 4941
rect 5261 4904 5265 4978
rect 5295 4953 5299 4996
rect 5286 4941 5299 4953
rect 5283 4864 5287 4941
rect 5305 4939 5309 4996
rect 5351 4939 5355 4996
rect 5361 4953 5365 4996
rect 5381 4990 5385 4996
rect 5486 4991 5490 4996
rect 5387 4978 5399 4990
rect 5361 4941 5374 4953
rect 5305 4927 5314 4939
rect 5346 4927 5355 4939
rect 5305 4864 5309 4927
rect 5351 4864 5355 4927
rect 5373 4864 5377 4941
rect 5395 4904 5399 4978
rect 5460 4987 5490 4991
rect 5460 4939 5466 4987
rect 5494 4982 5498 4996
rect 5485 4975 5498 4982
rect 5485 4973 5489 4975
rect 5514 4973 5518 4996
rect 5522 4988 5526 4996
rect 5522 4981 5539 4988
rect 5487 4961 5489 4973
rect 5466 4927 5469 4939
rect 5465 4904 5469 4927
rect 5485 4904 5489 4961
rect 5514 4932 5518 4961
rect 5533 4939 5539 4981
rect 5593 4976 5597 4996
rect 5583 4969 5597 4976
rect 5603 4976 5607 4996
rect 5603 4969 5611 4976
rect 5583 4953 5589 4969
rect 5586 4941 5589 4953
rect 5505 4926 5518 4932
rect 5525 4927 5533 4932
rect 5525 4926 5545 4927
rect 5505 4904 5509 4926
rect 5525 4904 5529 4926
rect 5585 4864 5589 4941
rect 5605 4953 5611 4969
rect 5605 4941 5614 4953
rect 5605 4864 5609 4941
rect 5652 4919 5656 4976
rect 5646 4907 5656 4919
rect 5640 4876 5646 4907
rect 5660 4899 5664 4976
rect 5668 4919 5672 4976
rect 5772 4973 5776 5016
rect 5765 4961 5774 4973
rect 5668 4907 5675 4919
rect 5687 4907 5695 4919
rect 5660 4880 5666 4887
rect 5660 4876 5675 4880
rect 5640 4872 5655 4876
rect 5651 4864 5655 4872
rect 5671 4864 5675 4876
rect 5691 4864 5695 4907
rect 5765 4904 5769 4961
rect 5794 4959 5798 4996
rect 5802 4992 5806 4996
rect 5802 4986 5821 4992
rect 5814 4973 5821 4986
rect 5973 4976 5977 4996
rect 5794 4924 5800 4947
rect 5814 4924 5821 4961
rect 5785 4918 5800 4924
rect 5805 4918 5821 4924
rect 5888 4919 5892 4976
rect 5785 4904 5789 4918
rect 5805 4904 5809 4918
rect 5865 4907 5873 4919
rect 5885 4907 5892 4919
rect 5865 4864 5869 4907
rect 5896 4899 5900 4976
rect 5904 4919 5908 4976
rect 5963 4969 5977 4976
rect 5983 4976 5987 4996
rect 6034 4988 6038 4996
rect 6021 4981 6038 4988
rect 5983 4969 5991 4976
rect 5963 4953 5969 4969
rect 5966 4941 5969 4953
rect 5904 4907 5914 4919
rect 5894 4880 5900 4887
rect 5885 4876 5900 4880
rect 5914 4876 5920 4907
rect 5885 4864 5889 4876
rect 5905 4872 5920 4876
rect 5905 4864 5909 4872
rect 5965 4864 5969 4941
rect 5985 4953 5991 4969
rect 5985 4941 5994 4953
rect 5985 4864 5989 4941
rect 6021 4939 6027 4981
rect 6042 4973 6046 4996
rect 6062 4982 6066 4996
rect 6070 4991 6074 4996
rect 6070 4987 6100 4991
rect 6062 4975 6075 4982
rect 6071 4973 6075 4975
rect 6071 4961 6073 4973
rect 6042 4932 6046 4961
rect 6027 4927 6035 4932
rect 6015 4926 6035 4927
rect 6042 4926 6055 4932
rect 6031 4904 6035 4926
rect 6051 4904 6055 4926
rect 6071 4904 6075 4961
rect 6094 4939 6100 4987
rect 6251 4991 6255 4996
rect 6242 4984 6255 4991
rect 6091 4927 6094 4939
rect 6091 4904 6095 4927
rect 6188 4919 6192 4976
rect 6165 4907 6173 4919
rect 6185 4907 6192 4919
rect 6165 4864 6169 4907
rect 6196 4899 6200 4976
rect 6204 4919 6208 4976
rect 6242 4939 6246 4984
rect 6271 4973 6275 4996
rect 6266 4961 6275 4973
rect 6204 4907 6214 4919
rect 6242 4916 6246 4927
rect 6242 4908 6260 4916
rect 6194 4880 6200 4887
rect 6185 4876 6200 4880
rect 6214 4876 6220 4907
rect 6256 4904 6260 4908
rect 6264 4904 6268 4961
rect 6291 4919 6295 4996
rect 6553 4976 6557 4996
rect 6388 4919 6392 4976
rect 6286 4907 6293 4919
rect 6365 4907 6373 4919
rect 6385 4907 6392 4919
rect 6185 4864 6189 4876
rect 6205 4872 6220 4876
rect 6205 4864 6209 4872
rect 6286 4864 6290 4907
rect 6365 4864 6369 4907
rect 6396 4899 6400 4976
rect 6404 4919 6408 4976
rect 6488 4919 6492 4976
rect 6404 4907 6414 4919
rect 6465 4907 6473 4919
rect 6485 4907 6492 4919
rect 6394 4880 6400 4887
rect 6385 4876 6400 4880
rect 6414 4876 6420 4907
rect 6385 4864 6389 4876
rect 6405 4872 6420 4876
rect 6405 4864 6409 4872
rect 6465 4864 6469 4907
rect 6496 4899 6500 4976
rect 6504 4919 6508 4976
rect 6549 4969 6557 4976
rect 6563 4976 6567 4996
rect 6563 4969 6577 4976
rect 6549 4953 6555 4969
rect 6546 4941 6555 4953
rect 6504 4907 6514 4919
rect 6494 4880 6500 4887
rect 6485 4876 6500 4880
rect 6514 4876 6520 4907
rect 6485 4864 6489 4876
rect 6505 4872 6520 4876
rect 6505 4864 6509 4872
rect 6551 4864 6555 4941
rect 6571 4953 6577 4969
rect 6645 4959 6649 5016
rect 6571 4941 6574 4953
rect 6645 4947 6654 4959
rect 6571 4864 6575 4941
rect 6645 4864 6649 4947
rect 43 4820 47 4824
rect 65 4820 69 4824
rect 123 4820 127 4824
rect 145 4820 149 4824
rect 205 4820 209 4824
rect 225 4820 229 4824
rect 271 4820 275 4824
rect 293 4820 297 4824
rect 301 4820 305 4824
rect 321 4820 325 4824
rect 329 4820 333 4824
rect 375 4820 379 4824
rect 395 4820 399 4824
rect 407 4820 411 4824
rect 427 4820 431 4824
rect 441 4820 445 4824
rect 461 4820 465 4824
rect 525 4820 529 4824
rect 545 4820 549 4824
rect 565 4820 569 4824
rect 625 4820 629 4824
rect 645 4820 649 4824
rect 691 4820 695 4824
rect 711 4820 715 4824
rect 785 4820 789 4824
rect 805 4820 809 4824
rect 851 4820 855 4824
rect 873 4820 877 4824
rect 881 4820 885 4824
rect 901 4820 905 4824
rect 909 4820 913 4824
rect 955 4820 959 4824
rect 975 4820 979 4824
rect 987 4820 991 4824
rect 1007 4820 1011 4824
rect 1021 4820 1025 4824
rect 1041 4820 1045 4824
rect 1103 4820 1107 4824
rect 1125 4820 1129 4824
rect 1185 4820 1189 4824
rect 1205 4820 1209 4824
rect 1225 4820 1229 4824
rect 1285 4820 1289 4824
rect 1305 4820 1309 4824
rect 1363 4820 1367 4824
rect 1385 4820 1389 4824
rect 1431 4820 1435 4824
rect 1451 4820 1455 4824
rect 1525 4820 1529 4824
rect 1545 4820 1549 4824
rect 1610 4820 1614 4824
rect 1632 4820 1636 4824
rect 1640 4820 1644 4824
rect 1705 4820 1709 4824
rect 1725 4820 1729 4824
rect 1790 4820 1794 4824
rect 1812 4820 1816 4824
rect 1820 4820 1824 4824
rect 1871 4820 1875 4824
rect 1891 4820 1895 4824
rect 1970 4820 1974 4824
rect 1992 4820 1996 4824
rect 2000 4820 2004 4824
rect 2070 4820 2074 4824
rect 2092 4820 2096 4824
rect 2100 4820 2104 4824
rect 2161 4820 2165 4824
rect 2183 4820 2187 4824
rect 2205 4820 2209 4824
rect 2251 4820 2255 4824
rect 2337 4820 2341 4824
rect 2345 4820 2349 4824
rect 2415 4820 2419 4824
rect 2435 4820 2439 4824
rect 2445 4820 2449 4824
rect 2505 4820 2509 4824
rect 2525 4820 2529 4824
rect 2590 4820 2594 4824
rect 2612 4820 2616 4824
rect 2620 4820 2624 4824
rect 2690 4820 2694 4824
rect 2712 4820 2716 4824
rect 2720 4820 2724 4824
rect 2785 4820 2789 4824
rect 2836 4820 2840 4824
rect 2844 4820 2848 4824
rect 2866 4820 2870 4824
rect 2950 4820 2954 4824
rect 2972 4820 2976 4824
rect 2980 4820 2984 4824
rect 3050 4820 3054 4824
rect 3072 4820 3076 4824
rect 3080 4820 3084 4824
rect 3157 4820 3161 4824
rect 3165 4820 3169 4824
rect 3225 4820 3229 4824
rect 3285 4820 3289 4824
rect 3305 4820 3309 4824
rect 3370 4820 3374 4824
rect 3392 4820 3396 4824
rect 3400 4820 3404 4824
rect 3455 4820 3459 4824
rect 3475 4820 3479 4824
rect 3489 4820 3493 4824
rect 3509 4820 3513 4824
rect 3521 4820 3525 4824
rect 3541 4820 3545 4824
rect 3587 4820 3591 4824
rect 3595 4820 3599 4824
rect 3615 4820 3619 4824
rect 3623 4820 3627 4824
rect 3645 4820 3649 4824
rect 3696 4820 3700 4824
rect 3704 4820 3708 4824
rect 3726 4820 3730 4824
rect 3805 4820 3809 4824
rect 3825 4820 3829 4824
rect 3845 4820 3849 4824
rect 3905 4820 3909 4824
rect 3925 4820 3929 4824
rect 3945 4820 3949 4824
rect 4005 4820 4009 4824
rect 4025 4820 4029 4824
rect 4045 4820 4049 4824
rect 4105 4820 4109 4824
rect 4161 4820 4165 4824
rect 4183 4820 4187 4824
rect 4205 4820 4209 4824
rect 4265 4820 4269 4824
rect 4285 4820 4289 4824
rect 4331 4820 4335 4824
rect 4353 4820 4357 4824
rect 4375 4820 4379 4824
rect 4450 4820 4454 4824
rect 4472 4820 4476 4824
rect 4480 4820 4484 4824
rect 4531 4820 4535 4824
rect 4551 4820 4555 4824
rect 4571 4820 4575 4824
rect 4636 4820 4640 4824
rect 4644 4820 4648 4824
rect 4666 4820 4670 4824
rect 4745 4820 4749 4824
rect 4765 4820 4769 4824
rect 4821 4820 4825 4824
rect 4843 4820 4847 4824
rect 4865 4820 4869 4824
rect 4925 4820 4929 4824
rect 4945 4820 4949 4824
rect 4991 4820 4995 4824
rect 5011 4820 5015 4824
rect 5071 4820 5075 4824
rect 5093 4820 5097 4824
rect 5115 4820 5119 4824
rect 5185 4820 5189 4824
rect 5205 4820 5209 4824
rect 5261 4820 5265 4824
rect 5283 4820 5287 4824
rect 5305 4820 5309 4824
rect 5351 4820 5355 4824
rect 5373 4820 5377 4824
rect 5395 4820 5399 4824
rect 5465 4820 5469 4824
rect 5485 4820 5489 4824
rect 5505 4820 5509 4824
rect 5525 4820 5529 4824
rect 5585 4820 5589 4824
rect 5605 4820 5609 4824
rect 5651 4820 5655 4824
rect 5671 4820 5675 4824
rect 5691 4820 5695 4824
rect 5765 4820 5769 4824
rect 5785 4820 5789 4824
rect 5805 4820 5809 4824
rect 5865 4820 5869 4824
rect 5885 4820 5889 4824
rect 5905 4820 5909 4824
rect 5965 4820 5969 4824
rect 5985 4820 5989 4824
rect 6031 4820 6035 4824
rect 6051 4820 6055 4824
rect 6071 4820 6075 4824
rect 6091 4820 6095 4824
rect 6165 4820 6169 4824
rect 6185 4820 6189 4824
rect 6205 4820 6209 4824
rect 6256 4820 6260 4824
rect 6264 4820 6268 4824
rect 6286 4820 6290 4824
rect 6365 4820 6369 4824
rect 6385 4820 6389 4824
rect 6405 4820 6409 4824
rect 6465 4820 6469 4824
rect 6485 4820 6489 4824
rect 6505 4820 6509 4824
rect 6551 4820 6555 4824
rect 6571 4820 6575 4824
rect 6645 4820 6649 4824
rect 31 4796 35 4800
rect 51 4796 55 4800
rect 71 4796 75 4800
rect 91 4796 95 4800
rect 111 4796 115 4800
rect 131 4796 135 4800
rect 151 4796 155 4800
rect 171 4796 175 4800
rect 257 4796 261 4800
rect 265 4796 269 4800
rect 325 4796 329 4800
rect 385 4796 389 4800
rect 405 4796 409 4800
rect 425 4796 429 4800
rect 485 4796 489 4800
rect 557 4796 561 4800
rect 565 4796 569 4800
rect 621 4796 625 4800
rect 643 4796 647 4800
rect 665 4796 669 4800
rect 711 4796 715 4800
rect 719 4796 723 4800
rect 803 4796 807 4800
rect 825 4796 829 4800
rect 885 4796 889 4800
rect 905 4796 909 4800
rect 951 4796 955 4800
rect 973 4796 977 4800
rect 981 4796 985 4800
rect 1001 4796 1005 4800
rect 1009 4796 1013 4800
rect 1055 4796 1059 4800
rect 1075 4796 1079 4800
rect 1087 4796 1091 4800
rect 1107 4796 1111 4800
rect 1121 4796 1125 4800
rect 1141 4796 1145 4800
rect 1210 4796 1214 4800
rect 1232 4796 1236 4800
rect 1240 4796 1244 4800
rect 1305 4796 1309 4800
rect 1325 4796 1329 4800
rect 1371 4796 1375 4800
rect 1391 4796 1395 4800
rect 1470 4796 1474 4800
rect 1492 4796 1496 4800
rect 1500 4796 1504 4800
rect 1551 4796 1555 4800
rect 1559 4796 1563 4800
rect 1631 4796 1635 4800
rect 1639 4796 1643 4800
rect 1711 4796 1715 4800
rect 1771 4796 1775 4800
rect 1779 4796 1783 4800
rect 1856 4796 1860 4800
rect 1864 4796 1868 4800
rect 1886 4796 1890 4800
rect 1951 4796 1955 4800
rect 1973 4796 1977 4800
rect 1981 4796 1985 4800
rect 2001 4796 2005 4800
rect 2009 4796 2013 4800
rect 2055 4796 2059 4800
rect 2075 4796 2079 4800
rect 2087 4796 2091 4800
rect 2107 4796 2111 4800
rect 2121 4796 2125 4800
rect 2141 4796 2145 4800
rect 2205 4796 2209 4800
rect 2225 4796 2229 4800
rect 2295 4796 2299 4800
rect 2315 4796 2319 4800
rect 2325 4796 2329 4800
rect 2371 4796 2375 4800
rect 2391 4796 2395 4800
rect 2451 4796 2455 4800
rect 2459 4796 2463 4800
rect 2531 4796 2535 4800
rect 2551 4796 2555 4800
rect 2571 4796 2575 4800
rect 2645 4796 2649 4800
rect 2691 4796 2695 4800
rect 2713 4796 2717 4800
rect 2721 4796 2725 4800
rect 2741 4796 2745 4800
rect 2749 4796 2753 4800
rect 2795 4796 2799 4800
rect 2815 4796 2819 4800
rect 2827 4796 2831 4800
rect 2847 4796 2851 4800
rect 2861 4796 2865 4800
rect 2881 4796 2885 4800
rect 2936 4796 2940 4800
rect 2944 4796 2948 4800
rect 2966 4796 2970 4800
rect 3031 4796 3035 4800
rect 3053 4796 3057 4800
rect 3061 4796 3065 4800
rect 3081 4796 3085 4800
rect 3089 4796 3093 4800
rect 3135 4796 3139 4800
rect 3155 4796 3159 4800
rect 3167 4796 3171 4800
rect 3187 4796 3191 4800
rect 3201 4796 3205 4800
rect 3221 4796 3225 4800
rect 3271 4796 3275 4800
rect 3293 4796 3297 4800
rect 3301 4796 3305 4800
rect 3321 4796 3325 4800
rect 3329 4796 3333 4800
rect 3375 4796 3379 4800
rect 3395 4796 3399 4800
rect 3407 4796 3411 4800
rect 3427 4796 3431 4800
rect 3441 4796 3445 4800
rect 3461 4796 3465 4800
rect 3530 4796 3534 4800
rect 3552 4796 3556 4800
rect 3560 4796 3564 4800
rect 3625 4796 3629 4800
rect 3685 4796 3689 4800
rect 3705 4796 3709 4800
rect 3770 4796 3774 4800
rect 3792 4796 3796 4800
rect 3800 4796 3804 4800
rect 3855 4796 3859 4800
rect 3875 4796 3879 4800
rect 3889 4796 3893 4800
rect 3909 4796 3913 4800
rect 3921 4796 3925 4800
rect 3941 4796 3945 4800
rect 3987 4796 3991 4800
rect 3995 4796 3999 4800
rect 4015 4796 4019 4800
rect 4023 4796 4027 4800
rect 4045 4796 4049 4800
rect 4105 4796 4109 4800
rect 4165 4796 4169 4800
rect 4185 4796 4189 4800
rect 4231 4796 4235 4800
rect 4253 4796 4257 4800
rect 4261 4796 4265 4800
rect 4281 4796 4285 4800
rect 4289 4796 4293 4800
rect 4335 4796 4339 4800
rect 4355 4796 4359 4800
rect 4367 4796 4371 4800
rect 4387 4796 4391 4800
rect 4401 4796 4405 4800
rect 4421 4796 4425 4800
rect 4485 4796 4489 4800
rect 4505 4796 4509 4800
rect 4525 4796 4529 4800
rect 4571 4796 4575 4800
rect 4631 4796 4635 4800
rect 4705 4796 4709 4800
rect 4756 4796 4760 4800
rect 4764 4796 4768 4800
rect 4786 4796 4790 4800
rect 4851 4796 4855 4800
rect 4859 4796 4863 4800
rect 4931 4796 4935 4800
rect 4951 4796 4955 4800
rect 5011 4796 5015 4800
rect 5031 4796 5035 4800
rect 5105 4796 5109 4800
rect 5125 4796 5129 4800
rect 5176 4796 5180 4800
rect 5184 4796 5188 4800
rect 5206 4796 5210 4800
rect 5295 4796 5299 4800
rect 5305 4796 5309 4800
rect 5335 4796 5339 4800
rect 5345 4796 5349 4800
rect 5391 4796 5395 4800
rect 5411 4796 5415 4800
rect 5485 4796 5489 4800
rect 5505 4796 5509 4800
rect 5551 4796 5555 4800
rect 5571 4796 5575 4800
rect 5591 4796 5595 4800
rect 5665 4796 5669 4800
rect 5685 4796 5689 4800
rect 5731 4796 5735 4800
rect 5751 4796 5755 4800
rect 5771 4796 5775 4800
rect 5845 4796 5849 4800
rect 5891 4796 5895 4800
rect 5911 4796 5915 4800
rect 5931 4796 5935 4800
rect 6001 4796 6005 4800
rect 6023 4796 6027 4800
rect 6045 4796 6049 4800
rect 6096 4796 6100 4800
rect 6104 4796 6108 4800
rect 6126 4796 6130 4800
rect 6205 4796 6209 4800
rect 6225 4796 6229 4800
rect 6271 4796 6275 4800
rect 6291 4796 6295 4800
rect 6311 4796 6315 4800
rect 6371 4796 6375 4800
rect 6391 4796 6395 4800
rect 6411 4796 6415 4800
rect 6481 4796 6485 4800
rect 6503 4796 6507 4800
rect 6525 4796 6529 4800
rect 6585 4796 6589 4800
rect 6605 4796 6609 4800
rect 6625 4796 6629 4800
rect 31 4659 35 4716
rect 51 4659 55 4716
rect 31 4647 34 4659
rect 46 4647 55 4659
rect 71 4656 75 4716
rect 91 4656 95 4716
rect 111 4656 115 4716
rect 131 4656 135 4716
rect 151 4656 155 4716
rect 171 4656 175 4716
rect 257 4693 261 4716
rect 246 4681 261 4693
rect 265 4693 269 4716
rect 265 4681 274 4693
rect 31 4624 35 4647
rect 51 4624 55 4647
rect 82 4644 95 4656
rect 122 4644 135 4656
rect 162 4644 175 4656
rect 71 4624 75 4644
rect 91 4624 95 4644
rect 111 4624 115 4644
rect 131 4624 135 4644
rect 151 4624 155 4644
rect 171 4624 175 4644
rect 245 4604 249 4681
rect 265 4604 269 4681
rect 325 4673 329 4756
rect 325 4661 334 4673
rect 325 4604 329 4661
rect 385 4659 389 4716
rect 405 4702 409 4716
rect 425 4702 429 4716
rect 405 4696 420 4702
rect 425 4696 441 4702
rect 414 4673 420 4696
rect 385 4647 394 4659
rect 392 4604 396 4647
rect 414 4624 418 4661
rect 434 4659 441 4696
rect 485 4673 489 4756
rect 557 4693 561 4716
rect 546 4681 561 4693
rect 565 4693 569 4716
rect 565 4681 574 4693
rect 485 4661 494 4673
rect 434 4634 441 4647
rect 422 4628 441 4634
rect 422 4624 426 4628
rect 485 4604 489 4661
rect 545 4604 549 4681
rect 565 4604 569 4681
rect 621 4642 625 4716
rect 643 4679 647 4756
rect 665 4693 669 4756
rect 711 4693 715 4716
rect 665 4681 674 4693
rect 706 4681 715 4693
rect 719 4693 723 4716
rect 803 4710 807 4716
rect 803 4698 805 4710
rect 825 4693 829 4756
rect 719 4681 734 4693
rect 825 4681 834 4693
rect 646 4667 659 4679
rect 621 4630 633 4642
rect 635 4624 639 4630
rect 655 4624 659 4667
rect 665 4624 669 4681
rect 711 4604 715 4681
rect 731 4604 735 4681
rect 803 4630 805 4642
rect 803 4624 807 4630
rect 825 4604 829 4681
rect 885 4679 889 4756
rect 886 4667 889 4679
rect 883 4651 889 4667
rect 905 4679 909 4756
rect 973 4753 977 4776
rect 969 4746 977 4753
rect 969 4717 973 4746
rect 981 4736 985 4776
rect 1001 4724 1005 4756
rect 1009 4752 1013 4756
rect 1009 4750 1045 4752
rect 1009 4748 1033 4750
rect 951 4704 955 4716
rect 969 4711 977 4717
rect 951 4692 953 4704
rect 905 4667 914 4679
rect 905 4651 911 4667
rect 883 4644 897 4651
rect 893 4624 897 4644
rect 903 4644 911 4651
rect 903 4624 907 4644
rect 951 4624 955 4692
rect 973 4665 977 4711
rect 973 4604 977 4653
rect 1001 4629 1007 4724
rect 983 4625 1007 4629
rect 983 4604 987 4625
rect 1003 4620 1021 4621
rect 1003 4616 1033 4620
rect 1003 4604 1007 4616
rect 1041 4612 1045 4738
rect 1055 4730 1059 4756
rect 1075 4750 1079 4756
rect 1011 4608 1045 4612
rect 1011 4604 1015 4608
rect 1057 4604 1061 4718
rect 1073 4628 1077 4738
rect 1087 4716 1091 4756
rect 1082 4704 1085 4716
rect 1082 4640 1086 4704
rect 1107 4697 1111 4756
rect 1102 4689 1111 4697
rect 1102 4660 1106 4689
rect 1121 4674 1125 4756
rect 1141 4673 1145 4716
rect 1210 4713 1214 4756
rect 1207 4701 1214 4713
rect 1082 4636 1115 4640
rect 1081 4616 1083 4628
rect 1079 4604 1083 4616
rect 1089 4616 1091 4628
rect 1089 4604 1093 4616
rect 1111 4604 1115 4636
rect 1121 4604 1125 4662
rect 1141 4624 1145 4661
rect 1205 4624 1209 4701
rect 1232 4659 1236 4716
rect 1240 4712 1244 4716
rect 1240 4704 1258 4712
rect 1254 4693 1258 4704
rect 1225 4647 1234 4659
rect 1225 4624 1229 4647
rect 1254 4636 1258 4681
rect 1305 4679 1309 4756
rect 1306 4667 1309 4679
rect 1303 4651 1309 4667
rect 1325 4679 1329 4756
rect 1371 4679 1375 4756
rect 1325 4667 1334 4679
rect 1366 4667 1375 4679
rect 1325 4651 1331 4667
rect 1303 4644 1317 4651
rect 1245 4629 1258 4636
rect 1245 4624 1249 4629
rect 1313 4624 1317 4644
rect 1323 4644 1331 4651
rect 1369 4651 1375 4667
rect 1391 4679 1395 4756
rect 1470 4713 1474 4756
rect 1467 4701 1474 4713
rect 1391 4667 1394 4679
rect 1391 4651 1397 4667
rect 1369 4644 1377 4651
rect 1323 4624 1327 4644
rect 1373 4624 1377 4644
rect 1383 4644 1397 4651
rect 1383 4624 1387 4644
rect 1465 4624 1469 4701
rect 1492 4659 1496 4716
rect 1500 4712 1504 4716
rect 1500 4704 1518 4712
rect 1514 4693 1518 4704
rect 1551 4693 1555 4716
rect 1546 4681 1555 4693
rect 1559 4693 1563 4716
rect 1631 4693 1635 4716
rect 1559 4681 1574 4693
rect 1626 4681 1635 4693
rect 1639 4693 1643 4716
rect 1639 4681 1654 4693
rect 1485 4647 1494 4659
rect 1485 4624 1489 4647
rect 1514 4636 1518 4681
rect 1505 4629 1518 4636
rect 1505 4624 1509 4629
rect 1551 4604 1555 4681
rect 1571 4604 1575 4681
rect 1631 4604 1635 4681
rect 1651 4604 1655 4681
rect 1711 4673 1715 4756
rect 1771 4693 1775 4716
rect 1766 4681 1775 4693
rect 1779 4693 1783 4716
rect 1856 4712 1860 4716
rect 1842 4704 1860 4712
rect 1842 4693 1846 4704
rect 1779 4681 1794 4693
rect 1706 4661 1715 4673
rect 1711 4604 1715 4661
rect 1771 4604 1775 4681
rect 1791 4604 1795 4681
rect 1842 4636 1846 4681
rect 1864 4659 1868 4716
rect 1886 4713 1890 4756
rect 1973 4753 1977 4776
rect 1969 4746 1977 4753
rect 1969 4717 1973 4746
rect 1981 4736 1985 4776
rect 2001 4724 2005 4756
rect 2009 4752 2013 4756
rect 2009 4750 2045 4752
rect 2009 4748 2033 4750
rect 1886 4701 1893 4713
rect 1951 4704 1955 4716
rect 1969 4711 1977 4717
rect 1866 4647 1875 4659
rect 1842 4629 1855 4636
rect 1851 4624 1855 4629
rect 1871 4624 1875 4647
rect 1891 4624 1895 4701
rect 1951 4692 1953 4704
rect 1951 4624 1955 4692
rect 1973 4665 1977 4711
rect 1973 4604 1977 4653
rect 2001 4629 2007 4724
rect 1983 4625 2007 4629
rect 1983 4604 1987 4625
rect 2003 4620 2021 4621
rect 2003 4616 2033 4620
rect 2003 4604 2007 4616
rect 2041 4612 2045 4738
rect 2055 4730 2059 4756
rect 2075 4750 2079 4756
rect 2011 4608 2045 4612
rect 2011 4604 2015 4608
rect 2057 4604 2061 4718
rect 2073 4628 2077 4738
rect 2087 4716 2091 4756
rect 2082 4704 2085 4716
rect 2082 4640 2086 4704
rect 2107 4697 2111 4756
rect 2102 4689 2111 4697
rect 2102 4660 2106 4689
rect 2121 4674 2125 4756
rect 2141 4673 2145 4716
rect 2205 4679 2209 4756
rect 2082 4636 2115 4640
rect 2081 4616 2083 4628
rect 2079 4604 2083 4616
rect 2089 4616 2091 4628
rect 2089 4604 2093 4616
rect 2111 4604 2115 4636
rect 2121 4604 2125 4662
rect 2206 4667 2209 4679
rect 2141 4624 2145 4661
rect 2203 4651 2209 4667
rect 2225 4679 2229 4756
rect 2295 4711 2299 4716
rect 2315 4693 2319 4716
rect 2325 4712 2329 4716
rect 2325 4707 2338 4712
rect 2225 4667 2234 4679
rect 2225 4651 2231 4667
rect 2203 4644 2217 4651
rect 2213 4624 2217 4644
rect 2223 4644 2231 4651
rect 2223 4624 2227 4644
rect 2285 4632 2295 4644
rect 2285 4624 2289 4632
rect 2315 4617 2319 4681
rect 2305 4611 2319 4617
rect 2334 4673 2338 4707
rect 2371 4679 2375 4756
rect 2366 4667 2375 4679
rect 2334 4616 2338 4661
rect 2369 4651 2375 4667
rect 2391 4679 2395 4756
rect 2451 4693 2455 4716
rect 2446 4681 2455 4693
rect 2459 4693 2463 4716
rect 2531 4702 2535 4716
rect 2551 4702 2555 4716
rect 2519 4696 2535 4702
rect 2540 4696 2555 4702
rect 2459 4681 2474 4693
rect 2391 4667 2394 4679
rect 2391 4651 2397 4667
rect 2369 4644 2377 4651
rect 2373 4624 2377 4644
rect 2383 4644 2397 4651
rect 2383 4624 2387 4644
rect 2325 4611 2338 4616
rect 2305 4604 2309 4611
rect 2325 4604 2329 4611
rect 2451 4604 2455 4681
rect 2471 4604 2475 4681
rect 2519 4659 2526 4696
rect 2540 4673 2546 4696
rect 2519 4634 2526 4647
rect 2519 4628 2538 4634
rect 2534 4624 2538 4628
rect 2542 4624 2546 4661
rect 2571 4659 2575 4716
rect 2566 4647 2575 4659
rect 2645 4673 2649 4756
rect 2713 4753 2717 4776
rect 2709 4746 2717 4753
rect 2709 4717 2713 4746
rect 2721 4736 2725 4776
rect 2741 4724 2745 4756
rect 2749 4752 2753 4756
rect 2749 4750 2785 4752
rect 2749 4748 2773 4750
rect 2691 4704 2695 4716
rect 2709 4711 2717 4717
rect 2691 4692 2693 4704
rect 2645 4661 2654 4673
rect 2564 4604 2568 4647
rect 2645 4604 2649 4661
rect 2691 4624 2695 4692
rect 2713 4665 2717 4711
rect 2713 4604 2717 4653
rect 2741 4629 2747 4724
rect 2723 4625 2747 4629
rect 2723 4604 2727 4625
rect 2743 4620 2761 4621
rect 2743 4616 2773 4620
rect 2743 4604 2747 4616
rect 2781 4612 2785 4738
rect 2795 4730 2799 4756
rect 2815 4750 2819 4756
rect 2751 4608 2785 4612
rect 2751 4604 2755 4608
rect 2797 4604 2801 4718
rect 2813 4628 2817 4738
rect 2827 4716 2831 4756
rect 2822 4704 2825 4716
rect 2822 4640 2826 4704
rect 2847 4697 2851 4756
rect 2842 4689 2851 4697
rect 2842 4660 2846 4689
rect 2861 4674 2865 4756
rect 2881 4673 2885 4716
rect 2936 4712 2940 4716
rect 2922 4704 2940 4712
rect 2922 4693 2926 4704
rect 2822 4636 2855 4640
rect 2821 4616 2823 4628
rect 2819 4604 2823 4616
rect 2829 4616 2831 4628
rect 2829 4604 2833 4616
rect 2851 4604 2855 4636
rect 2861 4604 2865 4662
rect 2881 4624 2885 4661
rect 2922 4636 2926 4681
rect 2944 4659 2948 4716
rect 2966 4713 2970 4756
rect 3053 4753 3057 4776
rect 3049 4746 3057 4753
rect 3049 4717 3053 4746
rect 3061 4736 3065 4776
rect 3081 4724 3085 4756
rect 3089 4752 3093 4756
rect 3089 4750 3125 4752
rect 3089 4748 3113 4750
rect 2966 4701 2973 4713
rect 3031 4704 3035 4716
rect 3049 4711 3057 4717
rect 2946 4647 2955 4659
rect 2922 4629 2935 4636
rect 2931 4624 2935 4629
rect 2951 4624 2955 4647
rect 2971 4624 2975 4701
rect 3031 4692 3033 4704
rect 3031 4624 3035 4692
rect 3053 4665 3057 4711
rect 3053 4604 3057 4653
rect 3081 4629 3087 4724
rect 3063 4625 3087 4629
rect 3063 4604 3067 4625
rect 3083 4620 3101 4621
rect 3083 4616 3113 4620
rect 3083 4604 3087 4616
rect 3121 4612 3125 4738
rect 3135 4730 3139 4756
rect 3155 4750 3159 4756
rect 3091 4608 3125 4612
rect 3091 4604 3095 4608
rect 3137 4604 3141 4718
rect 3153 4628 3157 4738
rect 3167 4716 3171 4756
rect 3162 4704 3165 4716
rect 3162 4640 3166 4704
rect 3187 4697 3191 4756
rect 3182 4689 3191 4697
rect 3182 4660 3186 4689
rect 3201 4674 3205 4756
rect 3293 4753 3297 4776
rect 3289 4746 3297 4753
rect 3289 4717 3293 4746
rect 3301 4736 3305 4776
rect 3321 4724 3325 4756
rect 3329 4752 3333 4756
rect 3329 4750 3365 4752
rect 3329 4748 3353 4750
rect 3221 4673 3225 4716
rect 3271 4704 3275 4716
rect 3289 4711 3297 4717
rect 3271 4692 3273 4704
rect 3162 4636 3195 4640
rect 3161 4616 3163 4628
rect 3159 4604 3163 4616
rect 3169 4616 3171 4628
rect 3169 4604 3173 4616
rect 3191 4604 3195 4636
rect 3201 4604 3205 4662
rect 3221 4624 3225 4661
rect 3271 4624 3275 4692
rect 3293 4665 3297 4711
rect 3293 4604 3297 4653
rect 3321 4629 3327 4724
rect 3303 4625 3327 4629
rect 3303 4604 3307 4625
rect 3323 4620 3341 4621
rect 3323 4616 3353 4620
rect 3323 4604 3327 4616
rect 3361 4612 3365 4738
rect 3375 4730 3379 4756
rect 3395 4750 3399 4756
rect 3331 4608 3365 4612
rect 3331 4604 3335 4608
rect 3377 4604 3381 4718
rect 3393 4628 3397 4738
rect 3407 4716 3411 4756
rect 3402 4704 3405 4716
rect 3402 4640 3406 4704
rect 3427 4697 3431 4756
rect 3422 4689 3431 4697
rect 3422 4660 3426 4689
rect 3441 4674 3445 4756
rect 3461 4673 3465 4716
rect 3530 4713 3534 4756
rect 3527 4701 3534 4713
rect 3402 4636 3435 4640
rect 3401 4616 3403 4628
rect 3399 4604 3403 4616
rect 3409 4616 3411 4628
rect 3409 4604 3413 4616
rect 3431 4604 3435 4636
rect 3441 4604 3445 4662
rect 3461 4624 3465 4661
rect 3525 4624 3529 4701
rect 3552 4659 3556 4716
rect 3560 4712 3564 4716
rect 3560 4704 3578 4712
rect 3574 4693 3578 4704
rect 3545 4647 3554 4659
rect 3545 4624 3549 4647
rect 3574 4636 3578 4681
rect 3565 4629 3578 4636
rect 3625 4659 3629 4716
rect 3685 4679 3689 4756
rect 3686 4667 3689 4679
rect 3625 4647 3634 4659
rect 3683 4651 3689 4667
rect 3705 4679 3709 4756
rect 3770 4713 3774 4756
rect 3767 4701 3774 4713
rect 3705 4667 3714 4679
rect 3705 4651 3711 4667
rect 3565 4624 3569 4629
rect 3625 4624 3629 4647
rect 3683 4644 3697 4651
rect 3693 4624 3697 4644
rect 3703 4644 3711 4651
rect 3703 4624 3707 4644
rect 3765 4624 3769 4701
rect 3792 4659 3796 4716
rect 3800 4712 3804 4716
rect 3800 4704 3818 4712
rect 3814 4693 3818 4704
rect 3785 4647 3794 4659
rect 3785 4624 3789 4647
rect 3814 4636 3818 4681
rect 3855 4673 3859 4716
rect 3875 4674 3879 4756
rect 3889 4697 3893 4756
rect 3909 4716 3913 4756
rect 3921 4750 3925 4756
rect 3915 4704 3918 4716
rect 3889 4689 3898 4697
rect 3805 4629 3818 4636
rect 3805 4624 3809 4629
rect 3855 4624 3859 4661
rect 3875 4604 3879 4662
rect 3894 4660 3898 4689
rect 3914 4640 3918 4704
rect 3885 4636 3918 4640
rect 3885 4604 3889 4636
rect 3923 4628 3927 4738
rect 3941 4730 3945 4756
rect 3987 4752 3991 4756
rect 3955 4750 3991 4752
rect 3967 4748 3991 4750
rect 3909 4616 3911 4628
rect 3907 4604 3911 4616
rect 3917 4616 3919 4628
rect 3917 4604 3921 4616
rect 3939 4604 3943 4718
rect 3955 4612 3959 4738
rect 3995 4724 3999 4756
rect 4015 4736 4019 4776
rect 4023 4753 4027 4776
rect 4023 4746 4031 4753
rect 3993 4629 3999 4724
rect 4027 4717 4031 4746
rect 4023 4711 4031 4717
rect 4023 4665 4027 4711
rect 4045 4704 4049 4716
rect 4047 4692 4049 4704
rect 3993 4625 4017 4629
rect 3979 4620 3997 4621
rect 3967 4616 3997 4620
rect 3955 4608 3989 4612
rect 3985 4604 3989 4608
rect 3993 4604 3997 4616
rect 4013 4604 4017 4625
rect 4023 4604 4027 4653
rect 4045 4624 4049 4692
rect 4105 4659 4109 4716
rect 4165 4679 4169 4756
rect 4166 4667 4169 4679
rect 4105 4647 4114 4659
rect 4163 4651 4169 4667
rect 4185 4679 4189 4756
rect 4253 4753 4257 4776
rect 4249 4746 4257 4753
rect 4249 4717 4253 4746
rect 4261 4736 4265 4776
rect 4281 4724 4285 4756
rect 4289 4752 4293 4756
rect 4289 4750 4325 4752
rect 4289 4748 4313 4750
rect 4231 4704 4235 4716
rect 4249 4711 4257 4717
rect 4231 4692 4233 4704
rect 4185 4667 4194 4679
rect 4185 4651 4191 4667
rect 4105 4624 4109 4647
rect 4163 4644 4177 4651
rect 4173 4624 4177 4644
rect 4183 4644 4191 4651
rect 4183 4624 4187 4644
rect 4231 4624 4235 4692
rect 4253 4665 4257 4711
rect 4253 4604 4257 4653
rect 4281 4629 4287 4724
rect 4263 4625 4287 4629
rect 4263 4604 4267 4625
rect 4283 4620 4301 4621
rect 4283 4616 4313 4620
rect 4283 4604 4287 4616
rect 4321 4612 4325 4738
rect 4335 4730 4339 4756
rect 4355 4750 4359 4756
rect 4291 4608 4325 4612
rect 4291 4604 4295 4608
rect 4337 4604 4341 4718
rect 4353 4628 4357 4738
rect 4367 4716 4371 4756
rect 4362 4704 4365 4716
rect 4362 4640 4366 4704
rect 4387 4697 4391 4756
rect 4382 4689 4391 4697
rect 4382 4660 4386 4689
rect 4401 4674 4405 4756
rect 4421 4673 4425 4716
rect 4485 4713 4489 4756
rect 4505 4744 4509 4756
rect 4525 4748 4529 4756
rect 4525 4744 4540 4748
rect 4505 4740 4520 4744
rect 4514 4733 4520 4740
rect 4485 4701 4493 4713
rect 4505 4701 4512 4713
rect 4362 4636 4395 4640
rect 4361 4616 4363 4628
rect 4359 4604 4363 4616
rect 4369 4616 4371 4628
rect 4369 4604 4373 4616
rect 4391 4604 4395 4636
rect 4401 4604 4405 4662
rect 4421 4624 4425 4661
rect 4508 4644 4512 4701
rect 4516 4644 4520 4721
rect 4534 4713 4540 4744
rect 4524 4701 4534 4713
rect 4524 4644 4528 4701
rect 4571 4673 4575 4756
rect 4566 4661 4575 4673
rect 4571 4604 4575 4661
rect 4631 4659 4635 4716
rect 4626 4647 4635 4659
rect 4631 4624 4635 4647
rect 4705 4673 4709 4756
rect 4756 4712 4760 4716
rect 4742 4704 4760 4712
rect 4742 4693 4746 4704
rect 4705 4661 4714 4673
rect 4705 4604 4709 4661
rect 4742 4636 4746 4681
rect 4764 4659 4768 4716
rect 4786 4713 4790 4756
rect 4786 4701 4793 4713
rect 4766 4647 4775 4659
rect 4742 4629 4755 4636
rect 4751 4624 4755 4629
rect 4771 4624 4775 4647
rect 4791 4624 4795 4701
rect 4851 4693 4855 4716
rect 4846 4681 4855 4693
rect 4859 4693 4863 4716
rect 4859 4681 4874 4693
rect 4851 4604 4855 4681
rect 4871 4604 4875 4681
rect 4931 4679 4935 4756
rect 4926 4667 4935 4679
rect 4929 4651 4935 4667
rect 4951 4679 4955 4756
rect 5011 4679 5015 4756
rect 4951 4667 4954 4679
rect 5006 4667 5015 4679
rect 4951 4651 4957 4667
rect 4929 4644 4937 4651
rect 4933 4624 4937 4644
rect 4943 4644 4957 4651
rect 5009 4651 5015 4667
rect 5031 4679 5035 4756
rect 5105 4679 5109 4756
rect 5031 4667 5034 4679
rect 5106 4667 5109 4679
rect 5031 4651 5037 4667
rect 5009 4644 5017 4651
rect 4943 4624 4947 4644
rect 5013 4624 5017 4644
rect 5023 4644 5037 4651
rect 5103 4651 5109 4667
rect 5125 4679 5129 4756
rect 5176 4712 5180 4716
rect 5162 4704 5180 4712
rect 5162 4693 5166 4704
rect 5125 4667 5134 4679
rect 5125 4651 5131 4667
rect 5103 4644 5117 4651
rect 5023 4624 5027 4644
rect 5113 4624 5117 4644
rect 5123 4644 5131 4651
rect 5123 4624 5127 4644
rect 5162 4636 5166 4681
rect 5184 4659 5188 4716
rect 5206 4713 5210 4756
rect 5206 4701 5213 4713
rect 5295 4712 5299 4716
rect 5285 4708 5299 4712
rect 5186 4647 5195 4659
rect 5162 4629 5175 4636
rect 5171 4624 5175 4629
rect 5191 4624 5195 4647
rect 5211 4624 5215 4701
rect 5285 4693 5289 4708
rect 5287 4681 5289 4693
rect 5285 4624 5289 4681
rect 5305 4659 5309 4716
rect 5335 4712 5339 4716
rect 5325 4708 5339 4712
rect 5345 4712 5349 4716
rect 5345 4708 5359 4712
rect 5325 4659 5331 4708
rect 5354 4693 5359 4708
rect 5325 4647 5334 4659
rect 5305 4624 5309 4647
rect 5325 4624 5329 4647
rect 5354 4635 5360 4681
rect 5391 4679 5395 4756
rect 5386 4667 5395 4679
rect 5389 4651 5395 4667
rect 5411 4679 5415 4756
rect 5485 4679 5489 4756
rect 5411 4667 5414 4679
rect 5486 4667 5489 4679
rect 5411 4651 5417 4667
rect 5389 4644 5397 4651
rect 5345 4631 5360 4635
rect 5345 4624 5349 4631
rect 5393 4624 5397 4644
rect 5403 4644 5417 4651
rect 5483 4651 5489 4667
rect 5505 4679 5509 4756
rect 5551 4748 5555 4756
rect 5540 4744 5555 4748
rect 5571 4744 5575 4756
rect 5540 4713 5546 4744
rect 5560 4740 5575 4744
rect 5560 4733 5566 4740
rect 5546 4701 5556 4713
rect 5505 4667 5514 4679
rect 5505 4651 5511 4667
rect 5483 4644 5497 4651
rect 5403 4624 5407 4644
rect 5493 4624 5497 4644
rect 5503 4644 5511 4651
rect 5552 4644 5556 4701
rect 5560 4644 5564 4721
rect 5591 4713 5595 4756
rect 5568 4701 5575 4713
rect 5587 4701 5595 4713
rect 5568 4644 5572 4701
rect 5665 4679 5669 4756
rect 5666 4667 5669 4679
rect 5663 4651 5669 4667
rect 5685 4679 5689 4756
rect 5731 4748 5735 4756
rect 5720 4744 5735 4748
rect 5751 4744 5755 4756
rect 5720 4713 5726 4744
rect 5740 4740 5755 4744
rect 5740 4733 5746 4740
rect 5726 4701 5736 4713
rect 5685 4667 5694 4679
rect 5685 4651 5691 4667
rect 5663 4644 5677 4651
rect 5503 4624 5507 4644
rect 5673 4624 5677 4644
rect 5683 4644 5691 4651
rect 5732 4644 5736 4701
rect 5740 4644 5744 4721
rect 5771 4713 5775 4756
rect 5748 4701 5755 4713
rect 5767 4701 5775 4713
rect 5748 4644 5752 4701
rect 5845 4673 5849 4756
rect 5891 4748 5895 4756
rect 5880 4744 5895 4748
rect 5911 4744 5915 4756
rect 5880 4713 5886 4744
rect 5900 4740 5915 4744
rect 5900 4733 5906 4740
rect 5886 4701 5896 4713
rect 5845 4661 5854 4673
rect 5683 4624 5687 4644
rect 5845 4604 5849 4661
rect 5892 4644 5896 4701
rect 5900 4644 5904 4721
rect 5931 4713 5935 4756
rect 5908 4701 5915 4713
rect 5927 4701 5935 4713
rect 5908 4644 5912 4701
rect 6001 4642 6005 4716
rect 6023 4679 6027 4756
rect 6045 4693 6049 4756
rect 6096 4712 6100 4716
rect 6082 4704 6100 4712
rect 6082 4693 6086 4704
rect 6045 4681 6054 4693
rect 6026 4667 6039 4679
rect 6001 4630 6013 4642
rect 6015 4624 6019 4630
rect 6035 4624 6039 4667
rect 6045 4624 6049 4681
rect 6082 4636 6086 4681
rect 6104 4659 6108 4716
rect 6126 4713 6130 4756
rect 6126 4701 6133 4713
rect 6106 4647 6115 4659
rect 6082 4629 6095 4636
rect 6091 4624 6095 4629
rect 6111 4624 6115 4647
rect 6131 4624 6135 4701
rect 6205 4679 6209 4756
rect 6206 4667 6209 4679
rect 6203 4651 6209 4667
rect 6225 4679 6229 4756
rect 6371 4748 6375 4756
rect 6360 4744 6375 4748
rect 6391 4744 6395 4756
rect 6271 4702 6275 4716
rect 6291 4702 6295 4716
rect 6259 4696 6275 4702
rect 6280 4696 6295 4702
rect 6225 4667 6234 4679
rect 6225 4651 6231 4667
rect 6259 4659 6266 4696
rect 6280 4673 6286 4696
rect 6203 4644 6217 4651
rect 6213 4624 6217 4644
rect 6223 4644 6231 4651
rect 6223 4624 6227 4644
rect 6259 4634 6266 4647
rect 6259 4628 6278 4634
rect 6274 4624 6278 4628
rect 6282 4624 6286 4661
rect 6311 4659 6315 4716
rect 6360 4713 6366 4744
rect 6380 4740 6395 4744
rect 6380 4733 6386 4740
rect 6366 4701 6376 4713
rect 6306 4647 6315 4659
rect 6304 4604 6308 4647
rect 6372 4644 6376 4701
rect 6380 4644 6384 4721
rect 6411 4713 6415 4756
rect 6388 4701 6395 4713
rect 6407 4701 6415 4713
rect 6388 4644 6392 4701
rect 6481 4642 6485 4716
rect 6503 4679 6507 4756
rect 6525 4693 6529 4756
rect 6585 4713 6589 4756
rect 6605 4744 6609 4756
rect 6625 4748 6629 4756
rect 6625 4744 6640 4748
rect 6605 4740 6620 4744
rect 6614 4733 6620 4740
rect 6585 4701 6593 4713
rect 6605 4701 6612 4713
rect 6525 4681 6534 4693
rect 6506 4667 6519 4679
rect 6481 4630 6493 4642
rect 6495 4624 6499 4630
rect 6515 4624 6519 4667
rect 6525 4624 6529 4681
rect 6608 4644 6612 4701
rect 6616 4644 6620 4721
rect 6634 4713 6640 4744
rect 6624 4701 6634 4713
rect 6624 4644 6628 4701
rect 31 4580 35 4584
rect 51 4580 55 4584
rect 71 4580 75 4584
rect 91 4580 95 4584
rect 111 4580 115 4584
rect 131 4580 135 4584
rect 151 4580 155 4584
rect 171 4580 175 4584
rect 245 4580 249 4584
rect 265 4580 269 4584
rect 325 4580 329 4584
rect 392 4580 396 4584
rect 414 4580 418 4584
rect 422 4580 426 4584
rect 485 4580 489 4584
rect 545 4580 549 4584
rect 565 4580 569 4584
rect 635 4580 639 4584
rect 655 4580 659 4584
rect 665 4580 669 4584
rect 711 4580 715 4584
rect 731 4580 735 4584
rect 803 4580 807 4584
rect 825 4580 829 4584
rect 893 4580 897 4584
rect 903 4580 907 4584
rect 951 4580 955 4584
rect 973 4580 977 4584
rect 983 4580 987 4584
rect 1003 4580 1007 4584
rect 1011 4580 1015 4584
rect 1057 4580 1061 4584
rect 1079 4580 1083 4584
rect 1089 4580 1093 4584
rect 1111 4580 1115 4584
rect 1121 4580 1125 4584
rect 1141 4580 1145 4584
rect 1205 4580 1209 4584
rect 1225 4580 1229 4584
rect 1245 4580 1249 4584
rect 1313 4580 1317 4584
rect 1323 4580 1327 4584
rect 1373 4580 1377 4584
rect 1383 4580 1387 4584
rect 1465 4580 1469 4584
rect 1485 4580 1489 4584
rect 1505 4580 1509 4584
rect 1551 4580 1555 4584
rect 1571 4580 1575 4584
rect 1631 4580 1635 4584
rect 1651 4580 1655 4584
rect 1711 4580 1715 4584
rect 1771 4580 1775 4584
rect 1791 4580 1795 4584
rect 1851 4580 1855 4584
rect 1871 4580 1875 4584
rect 1891 4580 1895 4584
rect 1951 4580 1955 4584
rect 1973 4580 1977 4584
rect 1983 4580 1987 4584
rect 2003 4580 2007 4584
rect 2011 4580 2015 4584
rect 2057 4580 2061 4584
rect 2079 4580 2083 4584
rect 2089 4580 2093 4584
rect 2111 4580 2115 4584
rect 2121 4580 2125 4584
rect 2141 4580 2145 4584
rect 2213 4580 2217 4584
rect 2223 4580 2227 4584
rect 2285 4580 2289 4584
rect 2305 4580 2309 4584
rect 2325 4580 2329 4584
rect 2373 4580 2377 4584
rect 2383 4580 2387 4584
rect 2451 4580 2455 4584
rect 2471 4580 2475 4584
rect 2534 4580 2538 4584
rect 2542 4580 2546 4584
rect 2564 4580 2568 4584
rect 2645 4580 2649 4584
rect 2691 4580 2695 4584
rect 2713 4580 2717 4584
rect 2723 4580 2727 4584
rect 2743 4580 2747 4584
rect 2751 4580 2755 4584
rect 2797 4580 2801 4584
rect 2819 4580 2823 4584
rect 2829 4580 2833 4584
rect 2851 4580 2855 4584
rect 2861 4580 2865 4584
rect 2881 4580 2885 4584
rect 2931 4580 2935 4584
rect 2951 4580 2955 4584
rect 2971 4580 2975 4584
rect 3031 4580 3035 4584
rect 3053 4580 3057 4584
rect 3063 4580 3067 4584
rect 3083 4580 3087 4584
rect 3091 4580 3095 4584
rect 3137 4580 3141 4584
rect 3159 4580 3163 4584
rect 3169 4580 3173 4584
rect 3191 4580 3195 4584
rect 3201 4580 3205 4584
rect 3221 4580 3225 4584
rect 3271 4580 3275 4584
rect 3293 4580 3297 4584
rect 3303 4580 3307 4584
rect 3323 4580 3327 4584
rect 3331 4580 3335 4584
rect 3377 4580 3381 4584
rect 3399 4580 3403 4584
rect 3409 4580 3413 4584
rect 3431 4580 3435 4584
rect 3441 4580 3445 4584
rect 3461 4580 3465 4584
rect 3525 4580 3529 4584
rect 3545 4580 3549 4584
rect 3565 4580 3569 4584
rect 3625 4580 3629 4584
rect 3693 4580 3697 4584
rect 3703 4580 3707 4584
rect 3765 4580 3769 4584
rect 3785 4580 3789 4584
rect 3805 4580 3809 4584
rect 3855 4580 3859 4584
rect 3875 4580 3879 4584
rect 3885 4580 3889 4584
rect 3907 4580 3911 4584
rect 3917 4580 3921 4584
rect 3939 4580 3943 4584
rect 3985 4580 3989 4584
rect 3993 4580 3997 4584
rect 4013 4580 4017 4584
rect 4023 4580 4027 4584
rect 4045 4580 4049 4584
rect 4105 4580 4109 4584
rect 4173 4580 4177 4584
rect 4183 4580 4187 4584
rect 4231 4580 4235 4584
rect 4253 4580 4257 4584
rect 4263 4580 4267 4584
rect 4283 4580 4287 4584
rect 4291 4580 4295 4584
rect 4337 4580 4341 4584
rect 4359 4580 4363 4584
rect 4369 4580 4373 4584
rect 4391 4580 4395 4584
rect 4401 4580 4405 4584
rect 4421 4580 4425 4584
rect 4508 4580 4512 4584
rect 4516 4580 4520 4584
rect 4524 4580 4528 4584
rect 4571 4580 4575 4584
rect 4631 4580 4635 4584
rect 4705 4580 4709 4584
rect 4751 4580 4755 4584
rect 4771 4580 4775 4584
rect 4791 4580 4795 4584
rect 4851 4580 4855 4584
rect 4871 4580 4875 4584
rect 4933 4580 4937 4584
rect 4943 4580 4947 4584
rect 5013 4580 5017 4584
rect 5023 4580 5027 4584
rect 5113 4580 5117 4584
rect 5123 4580 5127 4584
rect 5171 4580 5175 4584
rect 5191 4580 5195 4584
rect 5211 4580 5215 4584
rect 5285 4580 5289 4584
rect 5305 4580 5309 4584
rect 5325 4580 5329 4584
rect 5345 4580 5349 4584
rect 5393 4580 5397 4584
rect 5403 4580 5407 4584
rect 5493 4580 5497 4584
rect 5503 4580 5507 4584
rect 5552 4580 5556 4584
rect 5560 4580 5564 4584
rect 5568 4580 5572 4584
rect 5673 4580 5677 4584
rect 5683 4580 5687 4584
rect 5732 4580 5736 4584
rect 5740 4580 5744 4584
rect 5748 4580 5752 4584
rect 5845 4580 5849 4584
rect 5892 4580 5896 4584
rect 5900 4580 5904 4584
rect 5908 4580 5912 4584
rect 6015 4580 6019 4584
rect 6035 4580 6039 4584
rect 6045 4580 6049 4584
rect 6091 4580 6095 4584
rect 6111 4580 6115 4584
rect 6131 4580 6135 4584
rect 6213 4580 6217 4584
rect 6223 4580 6227 4584
rect 6274 4580 6278 4584
rect 6282 4580 6286 4584
rect 6304 4580 6308 4584
rect 6372 4580 6376 4584
rect 6380 4580 6384 4584
rect 6388 4580 6392 4584
rect 6495 4580 6499 4584
rect 6515 4580 6519 4584
rect 6525 4580 6529 4584
rect 6608 4580 6612 4584
rect 6616 4580 6620 4584
rect 6624 4580 6628 4584
rect 45 4556 49 4560
rect 105 4556 109 4560
rect 125 4556 129 4560
rect 185 4556 189 4560
rect 231 4556 235 4560
rect 251 4556 255 4560
rect 271 4556 275 4560
rect 345 4556 349 4560
rect 365 4556 369 4560
rect 411 4556 415 4560
rect 431 4556 435 4560
rect 451 4556 455 4560
rect 511 4556 515 4560
rect 531 4556 535 4560
rect 551 4556 555 4560
rect 614 4556 618 4560
rect 622 4556 626 4560
rect 644 4556 648 4560
rect 725 4556 729 4560
rect 771 4556 775 4560
rect 791 4556 795 4560
rect 851 4556 855 4560
rect 911 4556 915 4560
rect 931 4556 935 4560
rect 991 4556 995 4560
rect 1051 4556 1055 4560
rect 1071 4556 1075 4560
rect 1091 4556 1095 4560
rect 1111 4556 1115 4560
rect 1131 4556 1135 4560
rect 1151 4556 1155 4560
rect 1171 4556 1175 4560
rect 1191 4556 1195 4560
rect 1251 4556 1255 4560
rect 1273 4556 1277 4560
rect 1345 4556 1349 4560
rect 1405 4556 1409 4560
rect 1425 4556 1429 4560
rect 1493 4556 1497 4560
rect 1503 4556 1507 4560
rect 1553 4556 1557 4560
rect 1563 4556 1567 4560
rect 1645 4556 1649 4560
rect 1665 4556 1669 4560
rect 1685 4556 1689 4560
rect 1705 4556 1709 4560
rect 1755 4556 1759 4560
rect 1775 4556 1779 4560
rect 1785 4556 1789 4560
rect 1807 4556 1811 4560
rect 1817 4556 1821 4560
rect 1839 4556 1843 4560
rect 1885 4556 1889 4560
rect 1893 4556 1897 4560
rect 1913 4556 1917 4560
rect 1923 4556 1927 4560
rect 1945 4556 1949 4560
rect 1993 4556 1997 4560
rect 2003 4556 2007 4560
rect 2071 4556 2075 4560
rect 2093 4556 2097 4560
rect 2103 4556 2107 4560
rect 2123 4556 2127 4560
rect 2131 4556 2135 4560
rect 2177 4556 2181 4560
rect 2199 4556 2203 4560
rect 2209 4556 2213 4560
rect 2231 4556 2235 4560
rect 2241 4556 2245 4560
rect 2261 4556 2265 4560
rect 2311 4556 2315 4560
rect 2371 4556 2375 4560
rect 2391 4556 2395 4560
rect 2451 4556 2455 4560
rect 2471 4556 2475 4560
rect 2531 4556 2535 4560
rect 2591 4556 2595 4560
rect 2613 4556 2617 4560
rect 2623 4556 2627 4560
rect 2643 4556 2647 4560
rect 2651 4556 2655 4560
rect 2697 4556 2701 4560
rect 2719 4556 2723 4560
rect 2729 4556 2733 4560
rect 2751 4556 2755 4560
rect 2761 4556 2765 4560
rect 2781 4556 2785 4560
rect 2831 4556 2835 4560
rect 2851 4556 2855 4560
rect 2871 4556 2875 4560
rect 2933 4556 2937 4560
rect 2943 4556 2947 4560
rect 3025 4556 3029 4560
rect 3071 4556 3075 4560
rect 3091 4556 3095 4560
rect 3111 4556 3115 4560
rect 3171 4556 3175 4560
rect 3193 4556 3197 4560
rect 3203 4556 3207 4560
rect 3223 4556 3227 4560
rect 3231 4556 3235 4560
rect 3277 4556 3281 4560
rect 3299 4556 3303 4560
rect 3309 4556 3313 4560
rect 3331 4556 3335 4560
rect 3341 4556 3345 4560
rect 3361 4556 3365 4560
rect 3411 4556 3415 4560
rect 3431 4556 3435 4560
rect 3451 4556 3455 4560
rect 3525 4556 3529 4560
rect 3545 4556 3549 4560
rect 3565 4556 3569 4560
rect 3615 4556 3619 4560
rect 3635 4556 3639 4560
rect 3645 4556 3649 4560
rect 3667 4556 3671 4560
rect 3677 4556 3681 4560
rect 3699 4556 3703 4560
rect 3745 4556 3749 4560
rect 3753 4556 3757 4560
rect 3773 4556 3777 4560
rect 3783 4556 3787 4560
rect 3805 4556 3809 4560
rect 3851 4556 3855 4560
rect 3871 4556 3875 4560
rect 3891 4556 3895 4560
rect 3955 4556 3959 4560
rect 3975 4556 3979 4560
rect 3985 4556 3989 4560
rect 4007 4556 4011 4560
rect 4017 4556 4021 4560
rect 4039 4556 4043 4560
rect 4085 4556 4089 4560
rect 4093 4556 4097 4560
rect 4113 4556 4117 4560
rect 4123 4556 4127 4560
rect 4145 4556 4149 4560
rect 4228 4556 4232 4560
rect 4236 4556 4240 4560
rect 4244 4556 4248 4560
rect 4291 4556 4295 4560
rect 4311 4556 4315 4560
rect 4331 4556 4335 4560
rect 4405 4556 4409 4560
rect 4425 4556 4429 4560
rect 4492 4556 4496 4560
rect 4514 4556 4518 4560
rect 4522 4556 4526 4560
rect 4572 4556 4576 4560
rect 4580 4556 4584 4560
rect 4588 4556 4592 4560
rect 4685 4556 4689 4560
rect 4731 4556 4735 4560
rect 4751 4556 4755 4560
rect 4771 4556 4775 4560
rect 4845 4556 4849 4560
rect 4865 4556 4869 4560
rect 4885 4556 4889 4560
rect 4953 4556 4957 4560
rect 4963 4556 4967 4560
rect 5048 4556 5052 4560
rect 5056 4556 5060 4560
rect 5064 4556 5068 4560
rect 5111 4556 5115 4560
rect 5131 4556 5135 4560
rect 5151 4556 5155 4560
rect 5225 4556 5229 4560
rect 5245 4556 5249 4560
rect 5265 4556 5269 4560
rect 5311 4556 5315 4560
rect 5331 4556 5335 4560
rect 5351 4556 5355 4560
rect 5411 4556 5415 4560
rect 5508 4556 5512 4560
rect 5516 4556 5520 4560
rect 5524 4556 5528 4560
rect 5573 4556 5577 4560
rect 5583 4556 5587 4560
rect 5651 4556 5655 4560
rect 5671 4556 5675 4560
rect 5691 4556 5695 4560
rect 5773 4556 5777 4560
rect 5783 4556 5787 4560
rect 5868 4556 5872 4560
rect 5876 4556 5880 4560
rect 5884 4556 5888 4560
rect 5945 4556 5949 4560
rect 5965 4556 5969 4560
rect 5985 4556 5989 4560
rect 6031 4556 6035 4560
rect 6105 4556 6109 4560
rect 6152 4556 6156 4560
rect 6160 4556 6164 4560
rect 6168 4556 6172 4560
rect 6265 4556 6269 4560
rect 6285 4556 6289 4560
rect 6305 4556 6309 4560
rect 6352 4556 6356 4560
rect 6360 4556 6364 4560
rect 6368 4556 6372 4560
rect 6452 4556 6456 4560
rect 6460 4556 6464 4560
rect 6468 4556 6472 4560
rect 6551 4556 6555 4560
rect 6571 4556 6575 4560
rect 6591 4556 6595 4560
rect 6651 4556 6655 4560
rect 45 4479 49 4536
rect 45 4467 54 4479
rect 45 4384 49 4467
rect 105 4459 109 4536
rect 125 4459 129 4536
rect 185 4479 189 4536
rect 231 4511 235 4516
rect 222 4504 235 4511
rect 185 4467 194 4479
rect 106 4447 121 4459
rect 117 4424 121 4447
rect 125 4447 134 4459
rect 125 4424 129 4447
rect 185 4384 189 4467
rect 222 4459 226 4504
rect 251 4493 255 4516
rect 246 4481 255 4493
rect 222 4436 226 4447
rect 222 4428 240 4436
rect 236 4424 240 4428
rect 244 4424 248 4481
rect 271 4439 275 4516
rect 345 4459 349 4536
rect 365 4459 369 4536
rect 511 4529 515 4536
rect 531 4529 535 4536
rect 502 4524 515 4529
rect 411 4511 415 4516
rect 402 4504 415 4511
rect 402 4459 406 4504
rect 431 4493 435 4516
rect 426 4481 435 4493
rect 346 4447 361 4459
rect 266 4427 273 4439
rect 266 4384 270 4427
rect 357 4424 361 4447
rect 365 4447 374 4459
rect 365 4424 369 4447
rect 402 4436 406 4447
rect 402 4428 420 4436
rect 416 4424 420 4428
rect 424 4424 428 4481
rect 451 4439 455 4516
rect 502 4479 506 4524
rect 446 4427 453 4439
rect 502 4433 506 4467
rect 521 4523 535 4529
rect 521 4459 525 4523
rect 551 4508 555 4516
rect 614 4512 618 4516
rect 545 4496 555 4508
rect 599 4506 618 4512
rect 599 4493 606 4506
rect 502 4428 515 4433
rect 446 4384 450 4427
rect 511 4424 515 4428
rect 521 4424 525 4447
rect 599 4444 606 4481
rect 622 4479 626 4516
rect 644 4493 648 4536
rect 646 4481 655 4493
rect 620 4444 626 4467
rect 599 4438 615 4444
rect 620 4438 635 4444
rect 541 4424 545 4429
rect 611 4424 615 4438
rect 631 4424 635 4438
rect 651 4424 655 4481
rect 725 4479 729 4536
rect 725 4467 734 4479
rect 725 4384 729 4467
rect 771 4459 775 4536
rect 791 4459 795 4536
rect 851 4479 855 4536
rect 846 4467 855 4479
rect 766 4447 775 4459
rect 771 4424 775 4447
rect 779 4447 794 4459
rect 779 4424 783 4447
rect 851 4384 855 4467
rect 911 4459 915 4536
rect 931 4459 935 4536
rect 991 4479 995 4536
rect 986 4467 995 4479
rect 906 4447 915 4459
rect 911 4424 915 4447
rect 919 4447 934 4459
rect 919 4424 923 4447
rect 991 4384 995 4467
rect 1051 4493 1055 4516
rect 1071 4493 1075 4516
rect 1091 4496 1095 4516
rect 1111 4496 1115 4516
rect 1131 4496 1135 4516
rect 1151 4496 1155 4516
rect 1171 4496 1175 4516
rect 1191 4496 1195 4516
rect 1051 4481 1054 4493
rect 1066 4481 1075 4493
rect 1102 4484 1115 4496
rect 1142 4484 1155 4496
rect 1182 4484 1195 4496
rect 1051 4424 1055 4481
rect 1071 4424 1075 4481
rect 1091 4424 1095 4484
rect 1111 4424 1115 4484
rect 1131 4424 1135 4484
rect 1151 4424 1155 4484
rect 1171 4424 1175 4484
rect 1191 4424 1195 4484
rect 1251 4459 1255 4536
rect 1273 4510 1277 4516
rect 1275 4498 1277 4510
rect 1246 4447 1255 4459
rect 1251 4384 1255 4447
rect 1345 4479 1349 4536
rect 1345 4467 1354 4479
rect 1275 4430 1277 4442
rect 1273 4424 1277 4430
rect 1345 4384 1349 4467
rect 1405 4459 1409 4536
rect 1425 4459 1429 4536
rect 1493 4496 1497 4516
rect 1483 4489 1497 4496
rect 1503 4496 1507 4516
rect 1553 4496 1557 4516
rect 1503 4489 1511 4496
rect 1483 4473 1489 4489
rect 1486 4461 1489 4473
rect 1406 4447 1421 4459
rect 1417 4424 1421 4447
rect 1425 4447 1434 4459
rect 1425 4424 1429 4447
rect 1485 4384 1489 4461
rect 1505 4473 1511 4489
rect 1549 4489 1557 4496
rect 1563 4496 1567 4516
rect 1645 4512 1649 4516
rect 1665 4512 1669 4516
rect 1685 4512 1689 4516
rect 1705 4512 1709 4516
rect 1645 4508 1709 4512
rect 1563 4489 1577 4496
rect 1549 4473 1555 4489
rect 1505 4461 1514 4473
rect 1546 4461 1555 4473
rect 1505 4384 1509 4461
rect 1551 4384 1555 4461
rect 1571 4473 1577 4489
rect 1571 4461 1574 4473
rect 1571 4384 1575 4461
rect 1703 4459 1709 4508
rect 1755 4479 1759 4516
rect 1775 4478 1779 4536
rect 1785 4504 1789 4536
rect 1807 4524 1811 4536
rect 1809 4512 1811 4524
rect 1817 4524 1821 4536
rect 1817 4512 1819 4524
rect 1785 4500 1818 4504
rect 1706 4447 1709 4459
rect 1703 4432 1709 4447
rect 1645 4428 1709 4432
rect 1645 4424 1649 4428
rect 1665 4424 1669 4428
rect 1685 4424 1689 4428
rect 1705 4424 1709 4428
rect 1755 4424 1759 4467
rect 1775 4384 1779 4466
rect 1794 4451 1798 4480
rect 1789 4443 1798 4451
rect 1789 4384 1793 4443
rect 1814 4436 1818 4500
rect 1815 4424 1818 4436
rect 1809 4384 1813 4424
rect 1823 4402 1827 4512
rect 1839 4422 1843 4536
rect 1885 4532 1889 4536
rect 1855 4528 1889 4532
rect 1821 4384 1825 4390
rect 1841 4384 1845 4410
rect 1855 4402 1859 4528
rect 1893 4524 1897 4536
rect 1867 4520 1897 4524
rect 1879 4519 1897 4520
rect 1913 4515 1917 4536
rect 1893 4511 1917 4515
rect 1893 4416 1899 4511
rect 1923 4487 1927 4536
rect 1923 4429 1927 4475
rect 1945 4448 1949 4516
rect 1993 4496 1997 4516
rect 1989 4489 1997 4496
rect 2003 4496 2007 4516
rect 2003 4489 2017 4496
rect 1989 4473 1995 4489
rect 1986 4461 1995 4473
rect 1947 4436 1949 4448
rect 1923 4423 1931 4429
rect 1945 4424 1949 4436
rect 1867 4390 1891 4392
rect 1855 4388 1891 4390
rect 1887 4384 1891 4388
rect 1895 4384 1899 4416
rect 1915 4364 1919 4404
rect 1927 4394 1931 4423
rect 1923 4387 1931 4394
rect 1923 4364 1927 4387
rect 1991 4384 1995 4461
rect 2011 4473 2017 4489
rect 2011 4461 2014 4473
rect 2011 4384 2015 4461
rect 2071 4448 2075 4516
rect 2093 4487 2097 4536
rect 2103 4515 2107 4536
rect 2123 4524 2127 4536
rect 2131 4532 2135 4536
rect 2131 4528 2165 4532
rect 2123 4520 2153 4524
rect 2123 4519 2141 4520
rect 2103 4511 2127 4515
rect 2071 4436 2073 4448
rect 2071 4424 2075 4436
rect 2093 4429 2097 4475
rect 2089 4423 2097 4429
rect 2089 4394 2093 4423
rect 2121 4416 2127 4511
rect 2089 4387 2097 4394
rect 2093 4364 2097 4387
rect 2101 4364 2105 4404
rect 2121 4384 2125 4416
rect 2161 4402 2165 4528
rect 2177 4422 2181 4536
rect 2199 4524 2203 4536
rect 2201 4512 2203 4524
rect 2209 4524 2213 4536
rect 2209 4512 2211 4524
rect 2129 4390 2153 4392
rect 2129 4388 2165 4390
rect 2129 4384 2133 4388
rect 2175 4384 2179 4410
rect 2193 4402 2197 4512
rect 2231 4504 2235 4536
rect 2202 4500 2235 4504
rect 2202 4436 2206 4500
rect 2222 4451 2226 4480
rect 2241 4478 2245 4536
rect 2261 4479 2265 4516
rect 2311 4479 2315 4536
rect 2306 4467 2315 4479
rect 2222 4443 2231 4451
rect 2202 4424 2205 4436
rect 2195 4384 2199 4390
rect 2207 4384 2211 4424
rect 2227 4384 2231 4443
rect 2241 4384 2245 4466
rect 2261 4424 2265 4467
rect 2311 4384 2315 4467
rect 2371 4459 2375 4536
rect 2391 4459 2395 4536
rect 2451 4459 2455 4536
rect 2471 4459 2475 4536
rect 2531 4479 2535 4536
rect 2526 4467 2535 4479
rect 2366 4447 2375 4459
rect 2371 4424 2375 4447
rect 2379 4447 2394 4459
rect 2446 4447 2455 4459
rect 2379 4424 2383 4447
rect 2451 4424 2455 4447
rect 2459 4447 2474 4459
rect 2459 4424 2463 4447
rect 2531 4384 2535 4467
rect 2591 4448 2595 4516
rect 2613 4487 2617 4536
rect 2623 4515 2627 4536
rect 2643 4524 2647 4536
rect 2651 4532 2655 4536
rect 2651 4528 2685 4532
rect 2643 4520 2673 4524
rect 2643 4519 2661 4520
rect 2623 4511 2647 4515
rect 2591 4436 2593 4448
rect 2591 4424 2595 4436
rect 2613 4429 2617 4475
rect 2609 4423 2617 4429
rect 2609 4394 2613 4423
rect 2641 4416 2647 4511
rect 2609 4387 2617 4394
rect 2613 4364 2617 4387
rect 2621 4364 2625 4404
rect 2641 4384 2645 4416
rect 2681 4402 2685 4528
rect 2697 4422 2701 4536
rect 2719 4524 2723 4536
rect 2721 4512 2723 4524
rect 2729 4524 2733 4536
rect 2729 4512 2731 4524
rect 2649 4390 2673 4392
rect 2649 4388 2685 4390
rect 2649 4384 2653 4388
rect 2695 4384 2699 4410
rect 2713 4402 2717 4512
rect 2751 4504 2755 4536
rect 2722 4500 2755 4504
rect 2722 4436 2726 4500
rect 2742 4451 2746 4480
rect 2761 4478 2765 4536
rect 2781 4479 2785 4516
rect 2831 4511 2835 4516
rect 2822 4504 2835 4511
rect 2742 4443 2751 4451
rect 2722 4424 2725 4436
rect 2715 4384 2719 4390
rect 2727 4384 2731 4424
rect 2747 4384 2751 4443
rect 2761 4384 2765 4466
rect 2781 4424 2785 4467
rect 2822 4459 2826 4504
rect 2851 4493 2855 4516
rect 2846 4481 2855 4493
rect 2822 4436 2826 4447
rect 2822 4428 2840 4436
rect 2836 4424 2840 4428
rect 2844 4424 2848 4481
rect 2871 4439 2875 4516
rect 2933 4496 2937 4516
rect 2929 4489 2937 4496
rect 2943 4496 2947 4516
rect 2943 4489 2957 4496
rect 2929 4473 2935 4489
rect 2926 4461 2935 4473
rect 2866 4427 2873 4439
rect 2866 4384 2870 4427
rect 2931 4384 2935 4461
rect 2951 4473 2957 4489
rect 3025 4479 3029 4536
rect 3071 4511 3075 4516
rect 3062 4504 3075 4511
rect 2951 4461 2954 4473
rect 3025 4467 3034 4479
rect 2951 4384 2955 4461
rect 3025 4384 3029 4467
rect 3062 4459 3066 4504
rect 3091 4493 3095 4516
rect 3086 4481 3095 4493
rect 3062 4436 3066 4447
rect 3062 4428 3080 4436
rect 3076 4424 3080 4428
rect 3084 4424 3088 4481
rect 3111 4439 3115 4516
rect 3171 4448 3175 4516
rect 3193 4487 3197 4536
rect 3203 4515 3207 4536
rect 3223 4524 3227 4536
rect 3231 4532 3235 4536
rect 3231 4528 3265 4532
rect 3223 4520 3253 4524
rect 3223 4519 3241 4520
rect 3203 4511 3227 4515
rect 3106 4427 3113 4439
rect 3171 4436 3173 4448
rect 3106 4384 3110 4427
rect 3171 4424 3175 4436
rect 3193 4429 3197 4475
rect 3189 4423 3197 4429
rect 3189 4394 3193 4423
rect 3221 4416 3227 4511
rect 3189 4387 3197 4394
rect 3193 4364 3197 4387
rect 3201 4364 3205 4404
rect 3221 4384 3225 4416
rect 3261 4402 3265 4528
rect 3277 4422 3281 4536
rect 3299 4524 3303 4536
rect 3301 4512 3303 4524
rect 3309 4524 3313 4536
rect 3309 4512 3311 4524
rect 3229 4390 3253 4392
rect 3229 4388 3265 4390
rect 3229 4384 3233 4388
rect 3275 4384 3279 4410
rect 3293 4402 3297 4512
rect 3331 4504 3335 4536
rect 3302 4500 3335 4504
rect 3302 4436 3306 4500
rect 3322 4451 3326 4480
rect 3341 4478 3345 4536
rect 3361 4479 3365 4516
rect 3411 4511 3415 4516
rect 3402 4504 3415 4511
rect 3322 4443 3331 4451
rect 3302 4424 3305 4436
rect 3295 4384 3299 4390
rect 3307 4384 3311 4424
rect 3327 4384 3331 4443
rect 3341 4384 3345 4466
rect 3361 4424 3365 4467
rect 3402 4459 3406 4504
rect 3431 4493 3435 4516
rect 3426 4481 3435 4493
rect 3402 4436 3406 4447
rect 3402 4428 3420 4436
rect 3416 4424 3420 4428
rect 3424 4424 3428 4481
rect 3451 4439 3455 4516
rect 3525 4439 3529 4516
rect 3545 4493 3549 4516
rect 3565 4511 3569 4516
rect 3565 4504 3578 4511
rect 3545 4481 3554 4493
rect 3446 4427 3453 4439
rect 3527 4427 3534 4439
rect 3446 4384 3450 4427
rect 3530 4384 3534 4427
rect 3552 4424 3556 4481
rect 3574 4459 3578 4504
rect 3615 4479 3619 4516
rect 3635 4478 3639 4536
rect 3645 4504 3649 4536
rect 3667 4524 3671 4536
rect 3669 4512 3671 4524
rect 3677 4524 3681 4536
rect 3677 4512 3679 4524
rect 3645 4500 3678 4504
rect 3574 4436 3578 4447
rect 3560 4428 3578 4436
rect 3560 4424 3564 4428
rect 3615 4424 3619 4467
rect 3635 4384 3639 4466
rect 3654 4451 3658 4480
rect 3649 4443 3658 4451
rect 3649 4384 3653 4443
rect 3674 4436 3678 4500
rect 3675 4424 3678 4436
rect 3669 4384 3673 4424
rect 3683 4402 3687 4512
rect 3699 4422 3703 4536
rect 3745 4532 3749 4536
rect 3715 4528 3749 4532
rect 3681 4384 3685 4390
rect 3701 4384 3705 4410
rect 3715 4402 3719 4528
rect 3753 4524 3757 4536
rect 3727 4520 3757 4524
rect 3739 4519 3757 4520
rect 3773 4515 3777 4536
rect 3753 4511 3777 4515
rect 3753 4416 3759 4511
rect 3783 4487 3787 4536
rect 3783 4429 3787 4475
rect 3805 4448 3809 4516
rect 3851 4511 3855 4516
rect 3842 4504 3855 4511
rect 3842 4459 3846 4504
rect 3871 4493 3875 4516
rect 3866 4481 3875 4493
rect 3807 4436 3809 4448
rect 3783 4423 3791 4429
rect 3805 4424 3809 4436
rect 3842 4436 3846 4447
rect 3842 4428 3860 4436
rect 3856 4424 3860 4428
rect 3864 4424 3868 4481
rect 3891 4439 3895 4516
rect 3955 4479 3959 4516
rect 3975 4478 3979 4536
rect 3985 4504 3989 4536
rect 4007 4524 4011 4536
rect 4009 4512 4011 4524
rect 4017 4524 4021 4536
rect 4017 4512 4019 4524
rect 3985 4500 4018 4504
rect 3886 4427 3893 4439
rect 3727 4390 3751 4392
rect 3715 4388 3751 4390
rect 3747 4384 3751 4388
rect 3755 4384 3759 4416
rect 3775 4364 3779 4404
rect 3787 4394 3791 4423
rect 3783 4387 3791 4394
rect 3783 4364 3787 4387
rect 3886 4384 3890 4427
rect 3955 4424 3959 4467
rect 3975 4384 3979 4466
rect 3994 4451 3998 4480
rect 3989 4443 3998 4451
rect 3989 4384 3993 4443
rect 4014 4436 4018 4500
rect 4015 4424 4018 4436
rect 4009 4384 4013 4424
rect 4023 4402 4027 4512
rect 4039 4422 4043 4536
rect 4085 4532 4089 4536
rect 4055 4528 4089 4532
rect 4021 4384 4025 4390
rect 4041 4384 4045 4410
rect 4055 4402 4059 4528
rect 4093 4524 4097 4536
rect 4067 4520 4097 4524
rect 4079 4519 4097 4520
rect 4113 4515 4117 4536
rect 4093 4511 4117 4515
rect 4093 4416 4099 4511
rect 4123 4487 4127 4536
rect 4123 4429 4127 4475
rect 4145 4448 4149 4516
rect 4291 4511 4295 4516
rect 4282 4504 4295 4511
rect 4147 4436 4149 4448
rect 4228 4439 4232 4496
rect 4123 4423 4131 4429
rect 4145 4424 4149 4436
rect 4205 4427 4213 4439
rect 4225 4427 4232 4439
rect 4067 4390 4091 4392
rect 4055 4388 4091 4390
rect 4087 4384 4091 4388
rect 4095 4384 4099 4416
rect 4115 4364 4119 4404
rect 4127 4394 4131 4423
rect 4123 4387 4131 4394
rect 4123 4364 4127 4387
rect 4205 4384 4209 4427
rect 4236 4419 4240 4496
rect 4244 4439 4248 4496
rect 4282 4459 4286 4504
rect 4311 4493 4315 4516
rect 4306 4481 4315 4493
rect 4244 4427 4254 4439
rect 4282 4436 4286 4447
rect 4282 4428 4300 4436
rect 4234 4400 4240 4407
rect 4225 4396 4240 4400
rect 4254 4396 4260 4427
rect 4296 4424 4300 4428
rect 4304 4424 4308 4481
rect 4331 4439 4335 4516
rect 4405 4459 4409 4536
rect 4425 4459 4429 4536
rect 4492 4493 4496 4536
rect 4485 4481 4494 4493
rect 4406 4447 4421 4459
rect 4326 4427 4333 4439
rect 4225 4384 4229 4396
rect 4245 4392 4260 4396
rect 4245 4384 4249 4392
rect 4326 4384 4330 4427
rect 4417 4424 4421 4447
rect 4425 4447 4434 4459
rect 4425 4424 4429 4447
rect 4485 4424 4489 4481
rect 4514 4479 4518 4516
rect 4522 4512 4526 4516
rect 4522 4506 4541 4512
rect 4534 4493 4541 4506
rect 4514 4444 4520 4467
rect 4534 4444 4541 4481
rect 4505 4438 4520 4444
rect 4525 4438 4541 4444
rect 4572 4439 4576 4496
rect 4505 4424 4509 4438
rect 4525 4424 4529 4438
rect 4566 4427 4576 4439
rect 4560 4396 4566 4427
rect 4580 4419 4584 4496
rect 4588 4439 4592 4496
rect 4685 4479 4689 4536
rect 4865 4529 4869 4536
rect 4885 4529 4889 4536
rect 4865 4523 4879 4529
rect 4885 4524 4898 4529
rect 4731 4511 4735 4516
rect 4722 4504 4735 4511
rect 4685 4467 4694 4479
rect 4588 4427 4595 4439
rect 4607 4427 4615 4439
rect 4580 4400 4586 4407
rect 4580 4396 4595 4400
rect 4560 4392 4575 4396
rect 4571 4384 4575 4392
rect 4591 4384 4595 4396
rect 4611 4384 4615 4427
rect 4685 4384 4689 4467
rect 4722 4459 4726 4504
rect 4751 4493 4755 4516
rect 4746 4481 4755 4493
rect 4722 4436 4726 4447
rect 4722 4428 4740 4436
rect 4736 4424 4740 4428
rect 4744 4424 4748 4481
rect 4771 4439 4775 4516
rect 4845 4508 4849 4516
rect 4845 4496 4855 4508
rect 4875 4459 4879 4523
rect 4894 4479 4898 4524
rect 4953 4496 4957 4516
rect 4943 4489 4957 4496
rect 4963 4496 4967 4516
rect 5245 4529 5249 4536
rect 5265 4529 5269 4536
rect 5245 4523 5259 4529
rect 5265 4524 5278 4529
rect 5111 4511 5115 4516
rect 5102 4504 5115 4511
rect 4963 4489 4971 4496
rect 4943 4473 4949 4489
rect 4766 4427 4773 4439
rect 4766 4384 4770 4427
rect 4855 4424 4859 4429
rect 4875 4424 4879 4447
rect 4894 4433 4898 4467
rect 4946 4461 4949 4473
rect 4885 4428 4898 4433
rect 4885 4424 4889 4428
rect 4945 4384 4949 4461
rect 4965 4473 4971 4489
rect 4965 4461 4974 4473
rect 4965 4384 4969 4461
rect 5048 4439 5052 4496
rect 5025 4427 5033 4439
rect 5045 4427 5052 4439
rect 5025 4384 5029 4427
rect 5056 4419 5060 4496
rect 5064 4439 5068 4496
rect 5102 4459 5106 4504
rect 5131 4493 5135 4516
rect 5126 4481 5135 4493
rect 5064 4427 5074 4439
rect 5102 4436 5106 4447
rect 5102 4428 5120 4436
rect 5054 4400 5060 4407
rect 5045 4396 5060 4400
rect 5074 4396 5080 4427
rect 5116 4424 5120 4428
rect 5124 4424 5128 4481
rect 5151 4439 5155 4516
rect 5225 4508 5229 4516
rect 5225 4496 5235 4508
rect 5255 4459 5259 4523
rect 5274 4479 5278 4524
rect 5311 4511 5315 4516
rect 5302 4504 5315 4511
rect 5146 4427 5153 4439
rect 5045 4384 5049 4396
rect 5065 4392 5080 4396
rect 5065 4384 5069 4392
rect 5146 4384 5150 4427
rect 5235 4424 5239 4429
rect 5255 4424 5259 4447
rect 5274 4433 5278 4467
rect 5302 4459 5306 4504
rect 5331 4493 5335 4516
rect 5326 4481 5335 4493
rect 5265 4428 5278 4433
rect 5302 4436 5306 4447
rect 5302 4428 5320 4436
rect 5265 4424 5269 4428
rect 5316 4424 5320 4428
rect 5324 4424 5328 4481
rect 5351 4439 5355 4516
rect 5411 4479 5415 4536
rect 5573 4496 5577 4516
rect 5406 4467 5415 4479
rect 5346 4427 5353 4439
rect 5346 4384 5350 4427
rect 5411 4384 5415 4467
rect 5508 4439 5512 4496
rect 5485 4427 5493 4439
rect 5505 4427 5512 4439
rect 5485 4384 5489 4427
rect 5516 4419 5520 4496
rect 5524 4439 5528 4496
rect 5569 4489 5577 4496
rect 5583 4496 5587 4516
rect 5651 4511 5655 4516
rect 5642 4504 5655 4511
rect 5583 4489 5597 4496
rect 5569 4473 5575 4489
rect 5566 4461 5575 4473
rect 5524 4427 5534 4439
rect 5514 4400 5520 4407
rect 5505 4396 5520 4400
rect 5534 4396 5540 4427
rect 5505 4384 5509 4396
rect 5525 4392 5540 4396
rect 5525 4384 5529 4392
rect 5571 4384 5575 4461
rect 5591 4473 5597 4489
rect 5591 4461 5594 4473
rect 5591 4384 5595 4461
rect 5642 4459 5646 4504
rect 5671 4493 5675 4516
rect 5666 4481 5675 4493
rect 5642 4436 5646 4447
rect 5642 4428 5660 4436
rect 5656 4424 5660 4428
rect 5664 4424 5668 4481
rect 5691 4439 5695 4516
rect 5773 4496 5777 4516
rect 5763 4489 5777 4496
rect 5783 4496 5787 4516
rect 5783 4489 5791 4496
rect 5763 4473 5769 4489
rect 5766 4461 5769 4473
rect 5686 4427 5693 4439
rect 5686 4384 5690 4427
rect 5765 4384 5769 4461
rect 5785 4473 5791 4489
rect 5785 4461 5794 4473
rect 5785 4384 5789 4461
rect 5868 4439 5872 4496
rect 5845 4427 5853 4439
rect 5865 4427 5872 4439
rect 5845 4384 5849 4427
rect 5876 4419 5880 4496
rect 5884 4439 5888 4496
rect 5945 4439 5949 4516
rect 5965 4493 5969 4516
rect 5985 4511 5989 4516
rect 5985 4504 5998 4511
rect 5965 4481 5974 4493
rect 5884 4427 5894 4439
rect 5947 4427 5954 4439
rect 5874 4400 5880 4407
rect 5865 4396 5880 4400
rect 5894 4396 5900 4427
rect 5865 4384 5869 4396
rect 5885 4392 5900 4396
rect 5885 4384 5889 4392
rect 5950 4384 5954 4427
rect 5972 4424 5976 4481
rect 5994 4459 5998 4504
rect 6031 4479 6035 4536
rect 6026 4467 6035 4479
rect 5994 4436 5998 4447
rect 5980 4428 5998 4436
rect 5980 4424 5984 4428
rect 6031 4384 6035 4467
rect 6105 4479 6109 4536
rect 6105 4467 6114 4479
rect 6105 4384 6109 4467
rect 6152 4439 6156 4496
rect 6146 4427 6156 4439
rect 6140 4396 6146 4427
rect 6160 4419 6164 4496
rect 6168 4439 6172 4496
rect 6265 4439 6269 4516
rect 6285 4493 6289 4516
rect 6305 4511 6309 4516
rect 6305 4504 6318 4511
rect 6285 4481 6294 4493
rect 6168 4427 6175 4439
rect 6187 4427 6195 4439
rect 6267 4427 6274 4439
rect 6160 4400 6166 4407
rect 6160 4396 6175 4400
rect 6140 4392 6155 4396
rect 6151 4384 6155 4392
rect 6171 4384 6175 4396
rect 6191 4384 6195 4427
rect 6270 4384 6274 4427
rect 6292 4424 6296 4481
rect 6314 4459 6318 4504
rect 6551 4511 6555 4516
rect 6542 4504 6555 4511
rect 6314 4436 6318 4447
rect 6352 4439 6356 4496
rect 6300 4428 6318 4436
rect 6300 4424 6304 4428
rect 6346 4427 6356 4439
rect 6340 4396 6346 4427
rect 6360 4419 6364 4496
rect 6368 4439 6372 4496
rect 6452 4439 6456 4496
rect 6368 4427 6375 4439
rect 6387 4427 6395 4439
rect 6446 4427 6456 4439
rect 6360 4400 6366 4407
rect 6360 4396 6375 4400
rect 6340 4392 6355 4396
rect 6351 4384 6355 4392
rect 6371 4384 6375 4396
rect 6391 4384 6395 4427
rect 6440 4396 6446 4427
rect 6460 4419 6464 4496
rect 6468 4439 6472 4496
rect 6542 4459 6546 4504
rect 6571 4493 6575 4516
rect 6566 4481 6575 4493
rect 6468 4427 6475 4439
rect 6487 4427 6495 4439
rect 6542 4436 6546 4447
rect 6542 4428 6560 4436
rect 6460 4400 6466 4407
rect 6460 4396 6475 4400
rect 6440 4392 6455 4396
rect 6451 4384 6455 4392
rect 6471 4384 6475 4396
rect 6491 4384 6495 4427
rect 6556 4424 6560 4428
rect 6564 4424 6568 4481
rect 6591 4439 6595 4516
rect 6651 4479 6655 4536
rect 6646 4467 6655 4479
rect 6586 4427 6593 4439
rect 6586 4384 6590 4427
rect 6651 4384 6655 4467
rect 45 4340 49 4344
rect 117 4340 121 4344
rect 125 4340 129 4344
rect 185 4340 189 4344
rect 236 4340 240 4344
rect 244 4340 248 4344
rect 266 4340 270 4344
rect 357 4340 361 4344
rect 365 4340 369 4344
rect 416 4340 420 4344
rect 424 4340 428 4344
rect 446 4340 450 4344
rect 511 4340 515 4344
rect 521 4340 525 4344
rect 541 4340 545 4344
rect 611 4340 615 4344
rect 631 4340 635 4344
rect 651 4340 655 4344
rect 725 4340 729 4344
rect 771 4340 775 4344
rect 779 4340 783 4344
rect 851 4340 855 4344
rect 911 4340 915 4344
rect 919 4340 923 4344
rect 991 4340 995 4344
rect 1051 4340 1055 4344
rect 1071 4340 1075 4344
rect 1091 4340 1095 4344
rect 1111 4340 1115 4344
rect 1131 4340 1135 4344
rect 1151 4340 1155 4344
rect 1171 4340 1175 4344
rect 1191 4340 1195 4344
rect 1251 4340 1255 4344
rect 1273 4340 1277 4344
rect 1345 4340 1349 4344
rect 1417 4340 1421 4344
rect 1425 4340 1429 4344
rect 1485 4340 1489 4344
rect 1505 4340 1509 4344
rect 1551 4340 1555 4344
rect 1571 4340 1575 4344
rect 1645 4340 1649 4344
rect 1665 4340 1669 4344
rect 1685 4340 1689 4344
rect 1705 4340 1709 4344
rect 1755 4340 1759 4344
rect 1775 4340 1779 4344
rect 1789 4340 1793 4344
rect 1809 4340 1813 4344
rect 1821 4340 1825 4344
rect 1841 4340 1845 4344
rect 1887 4340 1891 4344
rect 1895 4340 1899 4344
rect 1915 4340 1919 4344
rect 1923 4340 1927 4344
rect 1945 4340 1949 4344
rect 1991 4340 1995 4344
rect 2011 4340 2015 4344
rect 2071 4340 2075 4344
rect 2093 4340 2097 4344
rect 2101 4340 2105 4344
rect 2121 4340 2125 4344
rect 2129 4340 2133 4344
rect 2175 4340 2179 4344
rect 2195 4340 2199 4344
rect 2207 4340 2211 4344
rect 2227 4340 2231 4344
rect 2241 4340 2245 4344
rect 2261 4340 2265 4344
rect 2311 4340 2315 4344
rect 2371 4340 2375 4344
rect 2379 4340 2383 4344
rect 2451 4340 2455 4344
rect 2459 4340 2463 4344
rect 2531 4340 2535 4344
rect 2591 4340 2595 4344
rect 2613 4340 2617 4344
rect 2621 4340 2625 4344
rect 2641 4340 2645 4344
rect 2649 4340 2653 4344
rect 2695 4340 2699 4344
rect 2715 4340 2719 4344
rect 2727 4340 2731 4344
rect 2747 4340 2751 4344
rect 2761 4340 2765 4344
rect 2781 4340 2785 4344
rect 2836 4340 2840 4344
rect 2844 4340 2848 4344
rect 2866 4340 2870 4344
rect 2931 4340 2935 4344
rect 2951 4340 2955 4344
rect 3025 4340 3029 4344
rect 3076 4340 3080 4344
rect 3084 4340 3088 4344
rect 3106 4340 3110 4344
rect 3171 4340 3175 4344
rect 3193 4340 3197 4344
rect 3201 4340 3205 4344
rect 3221 4340 3225 4344
rect 3229 4340 3233 4344
rect 3275 4340 3279 4344
rect 3295 4340 3299 4344
rect 3307 4340 3311 4344
rect 3327 4340 3331 4344
rect 3341 4340 3345 4344
rect 3361 4340 3365 4344
rect 3416 4340 3420 4344
rect 3424 4340 3428 4344
rect 3446 4340 3450 4344
rect 3530 4340 3534 4344
rect 3552 4340 3556 4344
rect 3560 4340 3564 4344
rect 3615 4340 3619 4344
rect 3635 4340 3639 4344
rect 3649 4340 3653 4344
rect 3669 4340 3673 4344
rect 3681 4340 3685 4344
rect 3701 4340 3705 4344
rect 3747 4340 3751 4344
rect 3755 4340 3759 4344
rect 3775 4340 3779 4344
rect 3783 4340 3787 4344
rect 3805 4340 3809 4344
rect 3856 4340 3860 4344
rect 3864 4340 3868 4344
rect 3886 4340 3890 4344
rect 3955 4340 3959 4344
rect 3975 4340 3979 4344
rect 3989 4340 3993 4344
rect 4009 4340 4013 4344
rect 4021 4340 4025 4344
rect 4041 4340 4045 4344
rect 4087 4340 4091 4344
rect 4095 4340 4099 4344
rect 4115 4340 4119 4344
rect 4123 4340 4127 4344
rect 4145 4340 4149 4344
rect 4205 4340 4209 4344
rect 4225 4340 4229 4344
rect 4245 4340 4249 4344
rect 4296 4340 4300 4344
rect 4304 4340 4308 4344
rect 4326 4340 4330 4344
rect 4417 4340 4421 4344
rect 4425 4340 4429 4344
rect 4485 4340 4489 4344
rect 4505 4340 4509 4344
rect 4525 4340 4529 4344
rect 4571 4340 4575 4344
rect 4591 4340 4595 4344
rect 4611 4340 4615 4344
rect 4685 4340 4689 4344
rect 4736 4340 4740 4344
rect 4744 4340 4748 4344
rect 4766 4340 4770 4344
rect 4855 4340 4859 4344
rect 4875 4340 4879 4344
rect 4885 4340 4889 4344
rect 4945 4340 4949 4344
rect 4965 4340 4969 4344
rect 5025 4340 5029 4344
rect 5045 4340 5049 4344
rect 5065 4340 5069 4344
rect 5116 4340 5120 4344
rect 5124 4340 5128 4344
rect 5146 4340 5150 4344
rect 5235 4340 5239 4344
rect 5255 4340 5259 4344
rect 5265 4340 5269 4344
rect 5316 4340 5320 4344
rect 5324 4340 5328 4344
rect 5346 4340 5350 4344
rect 5411 4340 5415 4344
rect 5485 4340 5489 4344
rect 5505 4340 5509 4344
rect 5525 4340 5529 4344
rect 5571 4340 5575 4344
rect 5591 4340 5595 4344
rect 5656 4340 5660 4344
rect 5664 4340 5668 4344
rect 5686 4340 5690 4344
rect 5765 4340 5769 4344
rect 5785 4340 5789 4344
rect 5845 4340 5849 4344
rect 5865 4340 5869 4344
rect 5885 4340 5889 4344
rect 5950 4340 5954 4344
rect 5972 4340 5976 4344
rect 5980 4340 5984 4344
rect 6031 4340 6035 4344
rect 6105 4340 6109 4344
rect 6151 4340 6155 4344
rect 6171 4340 6175 4344
rect 6191 4340 6195 4344
rect 6270 4340 6274 4344
rect 6292 4340 6296 4344
rect 6300 4340 6304 4344
rect 6351 4340 6355 4344
rect 6371 4340 6375 4344
rect 6391 4340 6395 4344
rect 6451 4340 6455 4344
rect 6471 4340 6475 4344
rect 6491 4340 6495 4344
rect 6556 4340 6560 4344
rect 6564 4340 6568 4344
rect 6586 4340 6590 4344
rect 6651 4340 6655 4344
rect 43 4316 47 4320
rect 65 4316 69 4320
rect 130 4316 134 4320
rect 152 4316 156 4320
rect 160 4316 164 4320
rect 216 4316 220 4320
rect 224 4316 228 4320
rect 246 4316 250 4320
rect 315 4316 319 4320
rect 335 4316 339 4320
rect 349 4316 353 4320
rect 369 4316 373 4320
rect 381 4316 385 4320
rect 401 4316 405 4320
rect 447 4316 451 4320
rect 455 4316 459 4320
rect 475 4316 479 4320
rect 483 4316 487 4320
rect 505 4316 509 4320
rect 551 4316 555 4320
rect 571 4316 575 4320
rect 645 4316 649 4320
rect 665 4316 669 4320
rect 685 4316 689 4320
rect 705 4316 709 4320
rect 765 4316 769 4320
rect 811 4316 815 4320
rect 833 4316 837 4320
rect 841 4316 845 4320
rect 861 4316 865 4320
rect 869 4316 873 4320
rect 915 4316 919 4320
rect 935 4316 939 4320
rect 947 4316 951 4320
rect 967 4316 971 4320
rect 981 4316 985 4320
rect 1001 4316 1005 4320
rect 1051 4316 1055 4320
rect 1071 4316 1075 4320
rect 1131 4316 1135 4320
rect 1153 4316 1157 4320
rect 1161 4316 1165 4320
rect 1181 4316 1185 4320
rect 1189 4316 1193 4320
rect 1235 4316 1239 4320
rect 1255 4316 1259 4320
rect 1267 4316 1271 4320
rect 1287 4316 1291 4320
rect 1301 4316 1305 4320
rect 1321 4316 1325 4320
rect 1371 4316 1375 4320
rect 1391 4316 1395 4320
rect 1451 4316 1455 4320
rect 1530 4316 1534 4320
rect 1552 4316 1556 4320
rect 1560 4316 1564 4320
rect 1625 4316 1629 4320
rect 1645 4316 1649 4320
rect 1665 4316 1669 4320
rect 1725 4316 1729 4320
rect 1745 4316 1749 4320
rect 1791 4316 1795 4320
rect 1811 4316 1815 4320
rect 1871 4316 1875 4320
rect 1893 4316 1897 4320
rect 1901 4316 1905 4320
rect 1921 4316 1925 4320
rect 1929 4316 1933 4320
rect 1975 4316 1979 4320
rect 1995 4316 1999 4320
rect 2007 4316 2011 4320
rect 2027 4316 2031 4320
rect 2041 4316 2045 4320
rect 2061 4316 2065 4320
rect 2111 4316 2115 4320
rect 2131 4316 2135 4320
rect 2210 4316 2214 4320
rect 2232 4316 2236 4320
rect 2240 4316 2244 4320
rect 2295 4316 2299 4320
rect 2315 4316 2319 4320
rect 2329 4316 2333 4320
rect 2349 4316 2353 4320
rect 2361 4316 2365 4320
rect 2381 4316 2385 4320
rect 2427 4316 2431 4320
rect 2435 4316 2439 4320
rect 2455 4316 2459 4320
rect 2463 4316 2467 4320
rect 2485 4316 2489 4320
rect 2557 4316 2561 4320
rect 2565 4316 2569 4320
rect 2611 4316 2615 4320
rect 2676 4316 2680 4320
rect 2684 4316 2688 4320
rect 2706 4316 2710 4320
rect 2771 4316 2775 4320
rect 2791 4316 2795 4320
rect 2870 4316 2874 4320
rect 2892 4316 2896 4320
rect 2900 4316 2904 4320
rect 2951 4316 2955 4320
rect 3011 4316 3015 4320
rect 3019 4316 3023 4320
rect 3105 4316 3109 4320
rect 3151 4316 3155 4320
rect 3173 4316 3177 4320
rect 3181 4316 3185 4320
rect 3201 4316 3205 4320
rect 3209 4316 3213 4320
rect 3255 4316 3259 4320
rect 3275 4316 3279 4320
rect 3287 4316 3291 4320
rect 3307 4316 3311 4320
rect 3321 4316 3325 4320
rect 3341 4316 3345 4320
rect 3391 4316 3395 4320
rect 3401 4316 3405 4320
rect 3431 4316 3435 4320
rect 3441 4316 3445 4320
rect 3511 4316 3515 4320
rect 3531 4316 3535 4320
rect 3591 4316 3595 4320
rect 3611 4316 3615 4320
rect 3631 4316 3635 4320
rect 3651 4316 3655 4320
rect 3671 4316 3675 4320
rect 3691 4316 3695 4320
rect 3711 4316 3715 4320
rect 3731 4316 3735 4320
rect 3791 4316 3795 4320
rect 3811 4316 3815 4320
rect 3871 4316 3875 4320
rect 3891 4316 3895 4320
rect 3965 4316 3969 4320
rect 3985 4316 3989 4320
rect 4031 4316 4035 4320
rect 4110 4316 4114 4320
rect 4132 4316 4136 4320
rect 4140 4316 4144 4320
rect 4196 4316 4200 4320
rect 4204 4316 4208 4320
rect 4226 4316 4230 4320
rect 4295 4316 4299 4320
rect 4315 4316 4319 4320
rect 4329 4316 4333 4320
rect 4349 4316 4353 4320
rect 4361 4316 4365 4320
rect 4381 4316 4385 4320
rect 4427 4316 4431 4320
rect 4435 4316 4439 4320
rect 4455 4316 4459 4320
rect 4463 4316 4467 4320
rect 4485 4316 4489 4320
rect 4550 4316 4554 4320
rect 4572 4316 4576 4320
rect 4580 4316 4584 4320
rect 4635 4316 4639 4320
rect 4655 4316 4659 4320
rect 4669 4316 4673 4320
rect 4689 4316 4693 4320
rect 4701 4316 4705 4320
rect 4721 4316 4725 4320
rect 4767 4316 4771 4320
rect 4775 4316 4779 4320
rect 4795 4316 4799 4320
rect 4803 4316 4807 4320
rect 4825 4316 4829 4320
rect 4885 4316 4889 4320
rect 4945 4316 4949 4320
rect 4965 4316 4969 4320
rect 4985 4316 4989 4320
rect 5031 4316 5035 4320
rect 5051 4316 5055 4320
rect 5071 4316 5075 4320
rect 5145 4316 5149 4320
rect 5196 4316 5200 4320
rect 5204 4316 5208 4320
rect 5226 4316 5230 4320
rect 5295 4316 5299 4320
rect 5315 4316 5319 4320
rect 5329 4316 5333 4320
rect 5349 4316 5353 4320
rect 5361 4316 5365 4320
rect 5381 4316 5385 4320
rect 5427 4316 5431 4320
rect 5435 4316 5439 4320
rect 5455 4316 5459 4320
rect 5463 4316 5467 4320
rect 5485 4316 5489 4320
rect 5531 4316 5535 4320
rect 5551 4316 5555 4320
rect 5611 4316 5615 4320
rect 5676 4316 5680 4320
rect 5684 4316 5688 4320
rect 5706 4316 5710 4320
rect 5781 4316 5785 4320
rect 5803 4316 5807 4320
rect 5825 4316 5829 4320
rect 5871 4316 5875 4320
rect 5891 4316 5895 4320
rect 5911 4316 5915 4320
rect 5985 4316 5989 4320
rect 6036 4316 6040 4320
rect 6044 4316 6048 4320
rect 6066 4316 6070 4320
rect 6131 4316 6135 4320
rect 6153 4316 6157 4320
rect 6211 4316 6215 4320
rect 6231 4316 6235 4320
rect 6301 4316 6305 4320
rect 6323 4316 6327 4320
rect 6345 4316 6349 4320
rect 6391 4316 6395 4320
rect 6411 4316 6415 4320
rect 6471 4316 6475 4320
rect 6545 4316 6549 4320
rect 6565 4316 6569 4320
rect 6585 4316 6589 4320
rect 6631 4316 6635 4320
rect 6651 4316 6655 4320
rect 6671 4316 6675 4320
rect 43 4230 47 4236
rect 43 4218 45 4230
rect 65 4213 69 4276
rect 130 4233 134 4276
rect 127 4221 134 4233
rect 65 4201 74 4213
rect 43 4150 45 4162
rect 43 4144 47 4150
rect 65 4124 69 4201
rect 125 4144 129 4221
rect 152 4179 156 4236
rect 160 4232 164 4236
rect 216 4232 220 4236
rect 160 4224 178 4232
rect 174 4213 178 4224
rect 202 4224 220 4232
rect 202 4213 206 4224
rect 145 4167 154 4179
rect 145 4144 149 4167
rect 174 4156 178 4201
rect 165 4149 178 4156
rect 202 4156 206 4201
rect 224 4179 228 4236
rect 246 4233 250 4276
rect 246 4221 253 4233
rect 226 4167 235 4179
rect 202 4149 215 4156
rect 165 4144 169 4149
rect 211 4144 215 4149
rect 231 4144 235 4167
rect 251 4144 255 4221
rect 315 4193 319 4236
rect 335 4194 339 4276
rect 349 4217 353 4276
rect 369 4236 373 4276
rect 381 4270 385 4276
rect 375 4224 378 4236
rect 349 4209 358 4217
rect 315 4144 319 4181
rect 335 4124 339 4182
rect 354 4180 358 4209
rect 374 4160 378 4224
rect 345 4156 378 4160
rect 345 4124 349 4156
rect 383 4148 387 4258
rect 401 4250 405 4276
rect 447 4272 451 4276
rect 415 4270 451 4272
rect 427 4268 451 4270
rect 369 4136 371 4148
rect 367 4124 371 4136
rect 377 4136 379 4148
rect 377 4124 381 4136
rect 399 4124 403 4238
rect 415 4132 419 4258
rect 455 4244 459 4276
rect 475 4256 479 4296
rect 483 4273 487 4296
rect 483 4266 491 4273
rect 453 4149 459 4244
rect 487 4237 491 4266
rect 483 4231 491 4237
rect 483 4185 487 4231
rect 505 4224 509 4236
rect 507 4212 509 4224
rect 453 4145 477 4149
rect 439 4140 457 4141
rect 427 4136 457 4140
rect 415 4128 449 4132
rect 445 4124 449 4128
rect 453 4124 457 4136
rect 473 4124 477 4145
rect 483 4124 487 4173
rect 505 4144 509 4212
rect 551 4199 555 4276
rect 546 4187 555 4199
rect 549 4171 555 4187
rect 571 4199 575 4276
rect 645 4213 649 4236
rect 646 4201 649 4213
rect 571 4187 574 4199
rect 571 4171 577 4187
rect 549 4164 557 4171
rect 553 4144 557 4164
rect 563 4164 577 4171
rect 563 4144 567 4164
rect 640 4153 646 4201
rect 665 4179 669 4236
rect 685 4214 689 4236
rect 705 4214 709 4236
rect 685 4208 698 4214
rect 705 4213 725 4214
rect 705 4208 713 4213
rect 694 4179 698 4208
rect 667 4167 669 4179
rect 665 4165 669 4167
rect 665 4158 678 4165
rect 640 4149 670 4153
rect 666 4144 670 4149
rect 674 4144 678 4158
rect 694 4144 698 4167
rect 713 4159 719 4201
rect 702 4152 719 4159
rect 765 4193 769 4276
rect 833 4273 837 4296
rect 829 4266 837 4273
rect 829 4237 833 4266
rect 841 4256 845 4296
rect 861 4244 865 4276
rect 869 4272 873 4276
rect 869 4270 905 4272
rect 869 4268 893 4270
rect 811 4224 815 4236
rect 829 4231 837 4237
rect 811 4212 813 4224
rect 765 4181 774 4193
rect 702 4144 706 4152
rect 765 4124 769 4181
rect 811 4144 815 4212
rect 833 4185 837 4231
rect 833 4124 837 4173
rect 861 4149 867 4244
rect 843 4145 867 4149
rect 843 4124 847 4145
rect 863 4140 881 4141
rect 863 4136 893 4140
rect 863 4124 867 4136
rect 901 4132 905 4258
rect 915 4250 919 4276
rect 935 4270 939 4276
rect 871 4128 905 4132
rect 871 4124 875 4128
rect 917 4124 921 4238
rect 933 4148 937 4258
rect 947 4236 951 4276
rect 942 4224 945 4236
rect 942 4160 946 4224
rect 967 4217 971 4276
rect 962 4209 971 4217
rect 962 4180 966 4209
rect 981 4194 985 4276
rect 1001 4193 1005 4236
rect 1051 4199 1055 4276
rect 942 4156 975 4160
rect 941 4136 943 4148
rect 939 4124 943 4136
rect 949 4136 951 4148
rect 949 4124 953 4136
rect 971 4124 975 4156
rect 981 4124 985 4182
rect 1046 4187 1055 4199
rect 1001 4144 1005 4181
rect 1049 4171 1055 4187
rect 1071 4199 1075 4276
rect 1153 4273 1157 4296
rect 1149 4266 1157 4273
rect 1149 4237 1153 4266
rect 1161 4256 1165 4296
rect 1181 4244 1185 4276
rect 1189 4272 1193 4276
rect 1189 4270 1225 4272
rect 1189 4268 1213 4270
rect 1131 4224 1135 4236
rect 1149 4231 1157 4237
rect 1131 4212 1133 4224
rect 1071 4187 1074 4199
rect 1071 4171 1077 4187
rect 1049 4164 1057 4171
rect 1053 4144 1057 4164
rect 1063 4164 1077 4171
rect 1063 4144 1067 4164
rect 1131 4144 1135 4212
rect 1153 4185 1157 4231
rect 1153 4124 1157 4173
rect 1181 4149 1187 4244
rect 1163 4145 1187 4149
rect 1163 4124 1167 4145
rect 1183 4140 1201 4141
rect 1183 4136 1213 4140
rect 1183 4124 1187 4136
rect 1221 4132 1225 4258
rect 1235 4250 1239 4276
rect 1255 4270 1259 4276
rect 1191 4128 1225 4132
rect 1191 4124 1195 4128
rect 1237 4124 1241 4238
rect 1253 4148 1257 4258
rect 1267 4236 1271 4276
rect 1262 4224 1265 4236
rect 1262 4160 1266 4224
rect 1287 4217 1291 4276
rect 1282 4209 1291 4217
rect 1282 4180 1286 4209
rect 1301 4194 1305 4276
rect 1321 4193 1325 4236
rect 1371 4199 1375 4276
rect 1262 4156 1295 4160
rect 1261 4136 1263 4148
rect 1259 4124 1263 4136
rect 1269 4136 1271 4148
rect 1269 4124 1273 4136
rect 1291 4124 1295 4156
rect 1301 4124 1305 4182
rect 1366 4187 1375 4199
rect 1321 4144 1325 4181
rect 1369 4171 1375 4187
rect 1391 4199 1395 4276
rect 1391 4187 1394 4199
rect 1451 4193 1455 4276
rect 1530 4233 1534 4276
rect 1527 4221 1534 4233
rect 1391 4171 1397 4187
rect 1446 4181 1455 4193
rect 1369 4164 1377 4171
rect 1373 4144 1377 4164
rect 1383 4164 1397 4171
rect 1383 4144 1387 4164
rect 1451 4124 1455 4181
rect 1525 4144 1529 4221
rect 1552 4179 1556 4236
rect 1560 4232 1564 4236
rect 1560 4224 1578 4232
rect 1574 4213 1578 4224
rect 1545 4167 1554 4179
rect 1545 4144 1549 4167
rect 1574 4156 1578 4201
rect 1625 4179 1629 4236
rect 1645 4222 1649 4236
rect 1665 4222 1669 4236
rect 1645 4216 1660 4222
rect 1665 4216 1681 4222
rect 1654 4193 1660 4216
rect 1625 4167 1634 4179
rect 1565 4149 1578 4156
rect 1565 4144 1569 4149
rect 1632 4124 1636 4167
rect 1654 4144 1658 4181
rect 1674 4179 1681 4216
rect 1725 4199 1729 4276
rect 1726 4187 1729 4199
rect 1723 4171 1729 4187
rect 1745 4199 1749 4276
rect 1791 4199 1795 4276
rect 1745 4187 1754 4199
rect 1786 4187 1795 4199
rect 1745 4171 1751 4187
rect 1674 4154 1681 4167
rect 1723 4164 1737 4171
rect 1662 4148 1681 4154
rect 1662 4144 1666 4148
rect 1733 4144 1737 4164
rect 1743 4164 1751 4171
rect 1789 4171 1795 4187
rect 1811 4199 1815 4276
rect 1893 4273 1897 4296
rect 1889 4266 1897 4273
rect 1889 4237 1893 4266
rect 1901 4256 1905 4296
rect 1921 4244 1925 4276
rect 1929 4272 1933 4276
rect 1929 4270 1965 4272
rect 1929 4268 1953 4270
rect 1871 4224 1875 4236
rect 1889 4231 1897 4237
rect 1871 4212 1873 4224
rect 1811 4187 1814 4199
rect 1811 4171 1817 4187
rect 1789 4164 1797 4171
rect 1743 4144 1747 4164
rect 1793 4144 1797 4164
rect 1803 4164 1817 4171
rect 1803 4144 1807 4164
rect 1871 4144 1875 4212
rect 1893 4185 1897 4231
rect 1893 4124 1897 4173
rect 1921 4149 1927 4244
rect 1903 4145 1927 4149
rect 1903 4124 1907 4145
rect 1923 4140 1941 4141
rect 1923 4136 1953 4140
rect 1923 4124 1927 4136
rect 1961 4132 1965 4258
rect 1975 4250 1979 4276
rect 1995 4270 1999 4276
rect 1931 4128 1965 4132
rect 1931 4124 1935 4128
rect 1977 4124 1981 4238
rect 1993 4148 1997 4258
rect 2007 4236 2011 4276
rect 2002 4224 2005 4236
rect 2002 4160 2006 4224
rect 2027 4217 2031 4276
rect 2022 4209 2031 4217
rect 2022 4180 2026 4209
rect 2041 4194 2045 4276
rect 2061 4193 2065 4236
rect 2111 4199 2115 4276
rect 2002 4156 2035 4160
rect 2001 4136 2003 4148
rect 1999 4124 2003 4136
rect 2009 4136 2011 4148
rect 2009 4124 2013 4136
rect 2031 4124 2035 4156
rect 2041 4124 2045 4182
rect 2106 4187 2115 4199
rect 2061 4144 2065 4181
rect 2109 4171 2115 4187
rect 2131 4199 2135 4276
rect 2210 4233 2214 4276
rect 2207 4221 2214 4233
rect 2131 4187 2134 4199
rect 2131 4171 2137 4187
rect 2109 4164 2117 4171
rect 2113 4144 2117 4164
rect 2123 4164 2137 4171
rect 2123 4144 2127 4164
rect 2205 4144 2209 4221
rect 2232 4179 2236 4236
rect 2240 4232 2244 4236
rect 2240 4224 2258 4232
rect 2254 4213 2258 4224
rect 2225 4167 2234 4179
rect 2225 4144 2229 4167
rect 2254 4156 2258 4201
rect 2295 4193 2299 4236
rect 2315 4194 2319 4276
rect 2329 4217 2333 4276
rect 2349 4236 2353 4276
rect 2361 4270 2365 4276
rect 2355 4224 2358 4236
rect 2329 4209 2338 4217
rect 2245 4149 2258 4156
rect 2245 4144 2249 4149
rect 2295 4144 2299 4181
rect 2315 4124 2319 4182
rect 2334 4180 2338 4209
rect 2354 4160 2358 4224
rect 2325 4156 2358 4160
rect 2325 4124 2329 4156
rect 2363 4148 2367 4258
rect 2381 4250 2385 4276
rect 2427 4272 2431 4276
rect 2395 4270 2431 4272
rect 2407 4268 2431 4270
rect 2349 4136 2351 4148
rect 2347 4124 2351 4136
rect 2357 4136 2359 4148
rect 2357 4124 2361 4136
rect 2379 4124 2383 4238
rect 2395 4132 2399 4258
rect 2435 4244 2439 4276
rect 2455 4256 2459 4296
rect 2463 4273 2467 4296
rect 2463 4266 2471 4273
rect 2433 4149 2439 4244
rect 2467 4237 2471 4266
rect 2463 4231 2471 4237
rect 2463 4185 2467 4231
rect 2485 4224 2489 4236
rect 2487 4212 2489 4224
rect 2557 4213 2561 4236
rect 2433 4145 2457 4149
rect 2419 4140 2437 4141
rect 2407 4136 2437 4140
rect 2395 4128 2429 4132
rect 2425 4124 2429 4128
rect 2433 4124 2437 4136
rect 2453 4124 2457 4145
rect 2463 4124 2467 4173
rect 2485 4144 2489 4212
rect 2546 4201 2561 4213
rect 2565 4213 2569 4236
rect 2565 4201 2574 4213
rect 2545 4124 2549 4201
rect 2565 4124 2569 4201
rect 2611 4193 2615 4276
rect 2676 4232 2680 4236
rect 2662 4224 2680 4232
rect 2662 4213 2666 4224
rect 2606 4181 2615 4193
rect 2611 4124 2615 4181
rect 2662 4156 2666 4201
rect 2684 4179 2688 4236
rect 2706 4233 2710 4276
rect 2706 4221 2713 4233
rect 2686 4167 2695 4179
rect 2662 4149 2675 4156
rect 2671 4144 2675 4149
rect 2691 4144 2695 4167
rect 2711 4144 2715 4221
rect 2771 4199 2775 4276
rect 2766 4187 2775 4199
rect 2769 4171 2775 4187
rect 2791 4199 2795 4276
rect 2870 4233 2874 4276
rect 2867 4221 2874 4233
rect 2791 4187 2794 4199
rect 2791 4171 2797 4187
rect 2769 4164 2777 4171
rect 2773 4144 2777 4164
rect 2783 4164 2797 4171
rect 2783 4144 2787 4164
rect 2865 4144 2869 4221
rect 2892 4179 2896 4236
rect 2900 4232 2904 4236
rect 2900 4224 2918 4232
rect 2914 4213 2918 4224
rect 2885 4167 2894 4179
rect 2885 4144 2889 4167
rect 2914 4156 2918 4201
rect 2951 4193 2955 4276
rect 3011 4213 3015 4236
rect 3006 4201 3015 4213
rect 3019 4213 3023 4236
rect 3019 4201 3034 4213
rect 2946 4181 2955 4193
rect 2905 4149 2918 4156
rect 2905 4144 2909 4149
rect 2951 4124 2955 4181
rect 3011 4124 3015 4201
rect 3031 4124 3035 4201
rect 3105 4193 3109 4276
rect 3173 4273 3177 4296
rect 3169 4266 3177 4273
rect 3169 4237 3173 4266
rect 3181 4256 3185 4296
rect 3201 4244 3205 4276
rect 3209 4272 3213 4276
rect 3209 4270 3245 4272
rect 3209 4268 3233 4270
rect 3151 4224 3155 4236
rect 3169 4231 3177 4237
rect 3151 4212 3153 4224
rect 3105 4181 3114 4193
rect 3105 4124 3109 4181
rect 3151 4144 3155 4212
rect 3173 4185 3177 4231
rect 3173 4124 3177 4173
rect 3201 4149 3207 4244
rect 3183 4145 3207 4149
rect 3183 4124 3187 4145
rect 3203 4140 3221 4141
rect 3203 4136 3233 4140
rect 3203 4124 3207 4136
rect 3241 4132 3245 4258
rect 3255 4250 3259 4276
rect 3275 4270 3279 4276
rect 3211 4128 3245 4132
rect 3211 4124 3215 4128
rect 3257 4124 3261 4238
rect 3273 4148 3277 4258
rect 3287 4236 3291 4276
rect 3282 4224 3285 4236
rect 3282 4160 3286 4224
rect 3307 4217 3311 4276
rect 3302 4209 3311 4217
rect 3302 4180 3306 4209
rect 3321 4194 3325 4276
rect 3341 4193 3345 4236
rect 3391 4232 3395 4236
rect 3381 4228 3395 4232
rect 3401 4232 3405 4236
rect 3401 4228 3415 4232
rect 3381 4213 3386 4228
rect 3282 4156 3315 4160
rect 3281 4136 3283 4148
rect 3279 4124 3283 4136
rect 3289 4136 3291 4148
rect 3289 4124 3293 4136
rect 3311 4124 3315 4156
rect 3321 4124 3325 4182
rect 3341 4144 3345 4181
rect 3380 4155 3386 4201
rect 3409 4179 3415 4228
rect 3431 4179 3435 4236
rect 3441 4232 3445 4236
rect 3441 4228 3455 4232
rect 3451 4213 3455 4228
rect 3451 4201 3453 4213
rect 3406 4167 3415 4179
rect 3380 4151 3395 4155
rect 3391 4144 3395 4151
rect 3411 4144 3415 4167
rect 3431 4144 3435 4167
rect 3451 4144 3455 4201
rect 3511 4199 3515 4276
rect 3506 4187 3515 4199
rect 3509 4171 3515 4187
rect 3531 4199 3535 4276
rect 3531 4187 3534 4199
rect 3531 4171 3537 4187
rect 3509 4164 3517 4171
rect 3513 4144 3517 4164
rect 3523 4164 3537 4171
rect 3591 4179 3595 4236
rect 3611 4179 3615 4236
rect 3591 4167 3594 4179
rect 3606 4167 3615 4179
rect 3631 4176 3635 4236
rect 3651 4176 3655 4236
rect 3671 4176 3675 4236
rect 3691 4176 3695 4236
rect 3711 4176 3715 4236
rect 3731 4176 3735 4236
rect 3791 4199 3795 4276
rect 3786 4187 3795 4199
rect 3523 4144 3527 4164
rect 3591 4144 3595 4167
rect 3611 4144 3615 4167
rect 3642 4164 3655 4176
rect 3682 4164 3695 4176
rect 3722 4164 3735 4176
rect 3789 4171 3795 4187
rect 3811 4199 3815 4276
rect 3871 4199 3875 4276
rect 3811 4187 3814 4199
rect 3866 4187 3875 4199
rect 3811 4171 3817 4187
rect 3789 4164 3797 4171
rect 3631 4144 3635 4164
rect 3651 4144 3655 4164
rect 3671 4144 3675 4164
rect 3691 4144 3695 4164
rect 3711 4144 3715 4164
rect 3731 4144 3735 4164
rect 3793 4144 3797 4164
rect 3803 4164 3817 4171
rect 3869 4171 3875 4187
rect 3891 4199 3895 4276
rect 3965 4199 3969 4276
rect 3891 4187 3894 4199
rect 3966 4187 3969 4199
rect 3891 4171 3897 4187
rect 3869 4164 3877 4171
rect 3803 4144 3807 4164
rect 3873 4144 3877 4164
rect 3883 4164 3897 4171
rect 3963 4171 3969 4187
rect 3985 4199 3989 4276
rect 3985 4187 3994 4199
rect 4031 4193 4035 4276
rect 4110 4233 4114 4276
rect 4107 4221 4114 4233
rect 3985 4171 3991 4187
rect 4026 4181 4035 4193
rect 3963 4164 3977 4171
rect 3883 4144 3887 4164
rect 3973 4144 3977 4164
rect 3983 4164 3991 4171
rect 3983 4144 3987 4164
rect 4031 4124 4035 4181
rect 4105 4144 4109 4221
rect 4132 4179 4136 4236
rect 4140 4232 4144 4236
rect 4196 4232 4200 4236
rect 4140 4224 4158 4232
rect 4154 4213 4158 4224
rect 4182 4224 4200 4232
rect 4182 4213 4186 4224
rect 4125 4167 4134 4179
rect 4125 4144 4129 4167
rect 4154 4156 4158 4201
rect 4145 4149 4158 4156
rect 4182 4156 4186 4201
rect 4204 4179 4208 4236
rect 4226 4233 4230 4276
rect 4226 4221 4233 4233
rect 4206 4167 4215 4179
rect 4182 4149 4195 4156
rect 4145 4144 4149 4149
rect 4191 4144 4195 4149
rect 4211 4144 4215 4167
rect 4231 4144 4235 4221
rect 4295 4193 4299 4236
rect 4315 4194 4319 4276
rect 4329 4217 4333 4276
rect 4349 4236 4353 4276
rect 4361 4270 4365 4276
rect 4355 4224 4358 4236
rect 4329 4209 4338 4217
rect 4295 4144 4299 4181
rect 4315 4124 4319 4182
rect 4334 4180 4338 4209
rect 4354 4160 4358 4224
rect 4325 4156 4358 4160
rect 4325 4124 4329 4156
rect 4363 4148 4367 4258
rect 4381 4250 4385 4276
rect 4427 4272 4431 4276
rect 4395 4270 4431 4272
rect 4407 4268 4431 4270
rect 4349 4136 4351 4148
rect 4347 4124 4351 4136
rect 4357 4136 4359 4148
rect 4357 4124 4361 4136
rect 4379 4124 4383 4238
rect 4395 4132 4399 4258
rect 4435 4244 4439 4276
rect 4455 4256 4459 4296
rect 4463 4273 4467 4296
rect 4463 4266 4471 4273
rect 4433 4149 4439 4244
rect 4467 4237 4471 4266
rect 4463 4231 4471 4237
rect 4463 4185 4467 4231
rect 4485 4224 4489 4236
rect 4550 4233 4554 4276
rect 4487 4212 4489 4224
rect 4547 4221 4554 4233
rect 4433 4145 4457 4149
rect 4419 4140 4437 4141
rect 4407 4136 4437 4140
rect 4395 4128 4429 4132
rect 4425 4124 4429 4128
rect 4433 4124 4437 4136
rect 4453 4124 4457 4145
rect 4463 4124 4467 4173
rect 4485 4144 4489 4212
rect 4545 4144 4549 4221
rect 4572 4179 4576 4236
rect 4580 4232 4584 4236
rect 4580 4224 4598 4232
rect 4594 4213 4598 4224
rect 4565 4167 4574 4179
rect 4565 4144 4569 4167
rect 4594 4156 4598 4201
rect 4635 4193 4639 4236
rect 4655 4194 4659 4276
rect 4669 4217 4673 4276
rect 4689 4236 4693 4276
rect 4701 4270 4705 4276
rect 4695 4224 4698 4236
rect 4669 4209 4678 4217
rect 4585 4149 4598 4156
rect 4585 4144 4589 4149
rect 4635 4144 4639 4181
rect 4655 4124 4659 4182
rect 4674 4180 4678 4209
rect 4694 4160 4698 4224
rect 4665 4156 4698 4160
rect 4665 4124 4669 4156
rect 4703 4148 4707 4258
rect 4721 4250 4725 4276
rect 4767 4272 4771 4276
rect 4735 4270 4771 4272
rect 4747 4268 4771 4270
rect 4689 4136 4691 4148
rect 4687 4124 4691 4136
rect 4697 4136 4699 4148
rect 4697 4124 4701 4136
rect 4719 4124 4723 4238
rect 4735 4132 4739 4258
rect 4775 4244 4779 4276
rect 4795 4256 4799 4296
rect 4803 4273 4807 4296
rect 4803 4266 4811 4273
rect 4773 4149 4779 4244
rect 4807 4237 4811 4266
rect 4803 4231 4811 4237
rect 5031 4268 5035 4276
rect 5020 4264 5035 4268
rect 5051 4264 5055 4276
rect 4803 4185 4807 4231
rect 4825 4224 4829 4236
rect 4827 4212 4829 4224
rect 4773 4145 4797 4149
rect 4759 4140 4777 4141
rect 4747 4136 4777 4140
rect 4735 4128 4769 4132
rect 4765 4124 4769 4128
rect 4773 4124 4777 4136
rect 4793 4124 4797 4145
rect 4803 4124 4807 4173
rect 4825 4144 4829 4212
rect 4885 4179 4889 4236
rect 4945 4179 4949 4236
rect 4965 4222 4969 4236
rect 4985 4222 4989 4236
rect 5020 4233 5026 4264
rect 5040 4260 5055 4264
rect 5040 4253 5046 4260
rect 4965 4216 4980 4222
rect 4985 4216 5001 4222
rect 5026 4221 5036 4233
rect 4974 4193 4980 4216
rect 4885 4167 4894 4179
rect 4945 4167 4954 4179
rect 4885 4144 4889 4167
rect 4952 4124 4956 4167
rect 4974 4144 4978 4181
rect 4994 4179 5001 4216
rect 4994 4154 5001 4167
rect 5032 4164 5036 4221
rect 5040 4164 5044 4241
rect 5071 4233 5075 4276
rect 5048 4221 5055 4233
rect 5067 4221 5075 4233
rect 5048 4164 5052 4221
rect 5145 4193 5149 4276
rect 5196 4232 5200 4236
rect 5182 4224 5200 4232
rect 5182 4213 5186 4224
rect 5145 4181 5154 4193
rect 4982 4148 5001 4154
rect 4982 4144 4986 4148
rect 5145 4124 5149 4181
rect 5182 4156 5186 4201
rect 5204 4179 5208 4236
rect 5226 4233 5230 4276
rect 5226 4221 5233 4233
rect 5206 4167 5215 4179
rect 5182 4149 5195 4156
rect 5191 4144 5195 4149
rect 5211 4144 5215 4167
rect 5231 4144 5235 4221
rect 5295 4193 5299 4236
rect 5315 4194 5319 4276
rect 5329 4217 5333 4276
rect 5349 4236 5353 4276
rect 5361 4270 5365 4276
rect 5355 4224 5358 4236
rect 5329 4209 5338 4217
rect 5295 4144 5299 4181
rect 5315 4124 5319 4182
rect 5334 4180 5338 4209
rect 5354 4160 5358 4224
rect 5325 4156 5358 4160
rect 5325 4124 5329 4156
rect 5363 4148 5367 4258
rect 5381 4250 5385 4276
rect 5427 4272 5431 4276
rect 5395 4270 5431 4272
rect 5407 4268 5431 4270
rect 5349 4136 5351 4148
rect 5347 4124 5351 4136
rect 5357 4136 5359 4148
rect 5357 4124 5361 4136
rect 5379 4124 5383 4238
rect 5395 4132 5399 4258
rect 5435 4244 5439 4276
rect 5455 4256 5459 4296
rect 5463 4273 5467 4296
rect 5463 4266 5471 4273
rect 5433 4149 5439 4244
rect 5467 4237 5471 4266
rect 5463 4231 5471 4237
rect 5463 4185 5467 4231
rect 5485 4224 5489 4236
rect 5487 4212 5489 4224
rect 5433 4145 5457 4149
rect 5419 4140 5437 4141
rect 5407 4136 5437 4140
rect 5395 4128 5429 4132
rect 5425 4124 5429 4128
rect 5433 4124 5437 4136
rect 5453 4124 5457 4145
rect 5463 4124 5467 4173
rect 5485 4144 5489 4212
rect 5531 4199 5535 4276
rect 5526 4187 5535 4199
rect 5529 4171 5535 4187
rect 5551 4199 5555 4276
rect 5551 4187 5554 4199
rect 5611 4193 5615 4276
rect 5676 4232 5680 4236
rect 5662 4224 5680 4232
rect 5662 4213 5666 4224
rect 5551 4171 5557 4187
rect 5606 4181 5615 4193
rect 5529 4164 5537 4171
rect 5533 4144 5537 4164
rect 5543 4164 5557 4171
rect 5543 4144 5547 4164
rect 5611 4124 5615 4181
rect 5662 4156 5666 4201
rect 5684 4179 5688 4236
rect 5706 4233 5710 4276
rect 5706 4221 5713 4233
rect 5686 4167 5695 4179
rect 5662 4149 5675 4156
rect 5671 4144 5675 4149
rect 5691 4144 5695 4167
rect 5711 4144 5715 4221
rect 5781 4162 5785 4236
rect 5803 4199 5807 4276
rect 5825 4213 5829 4276
rect 5871 4268 5875 4276
rect 5860 4264 5875 4268
rect 5891 4264 5895 4276
rect 5860 4233 5866 4264
rect 5880 4260 5895 4264
rect 5880 4253 5886 4260
rect 5866 4221 5876 4233
rect 5825 4201 5834 4213
rect 5806 4187 5819 4199
rect 5781 4150 5793 4162
rect 5795 4144 5799 4150
rect 5815 4144 5819 4187
rect 5825 4144 5829 4201
rect 5872 4164 5876 4221
rect 5880 4164 5884 4241
rect 5911 4233 5915 4276
rect 5888 4221 5895 4233
rect 5907 4221 5915 4233
rect 5888 4164 5892 4221
rect 5985 4179 5989 4236
rect 6036 4232 6040 4236
rect 6022 4224 6040 4232
rect 6022 4213 6026 4224
rect 5985 4167 5994 4179
rect 5985 4144 5989 4167
rect 6022 4156 6026 4201
rect 6044 4179 6048 4236
rect 6066 4233 6070 4276
rect 6066 4221 6073 4233
rect 6046 4167 6055 4179
rect 6022 4149 6035 4156
rect 6031 4144 6035 4149
rect 6051 4144 6055 4167
rect 6071 4144 6075 4221
rect 6131 4213 6135 4276
rect 6153 4230 6157 4236
rect 6155 4218 6157 4230
rect 6126 4201 6135 4213
rect 6131 4124 6135 4201
rect 6211 4199 6215 4276
rect 6206 4187 6215 4199
rect 6209 4171 6215 4187
rect 6231 4199 6235 4276
rect 6231 4187 6234 4199
rect 6231 4171 6237 4187
rect 6209 4164 6217 4171
rect 6155 4150 6157 4162
rect 6153 4144 6157 4150
rect 6213 4144 6217 4164
rect 6223 4164 6237 4171
rect 6223 4144 6227 4164
rect 6301 4162 6305 4236
rect 6323 4199 6327 4276
rect 6345 4213 6349 4276
rect 6345 4201 6354 4213
rect 6326 4187 6339 4199
rect 6301 4150 6313 4162
rect 6315 4144 6319 4150
rect 6335 4144 6339 4187
rect 6345 4144 6349 4201
rect 6391 4199 6395 4276
rect 6386 4187 6395 4199
rect 6389 4171 6395 4187
rect 6411 4199 6415 4276
rect 6411 4187 6414 4199
rect 6471 4193 6475 4276
rect 6631 4268 6635 4276
rect 6620 4264 6635 4268
rect 6651 4264 6655 4276
rect 6411 4171 6417 4187
rect 6466 4181 6475 4193
rect 6389 4164 6397 4171
rect 6393 4144 6397 4164
rect 6403 4164 6417 4171
rect 6403 4144 6407 4164
rect 6471 4124 6475 4181
rect 6545 4179 6549 4236
rect 6565 4222 6569 4236
rect 6585 4222 6589 4236
rect 6620 4233 6626 4264
rect 6640 4260 6655 4264
rect 6640 4253 6646 4260
rect 6565 4216 6580 4222
rect 6585 4216 6601 4222
rect 6626 4221 6636 4233
rect 6574 4193 6580 4216
rect 6545 4167 6554 4179
rect 6552 4124 6556 4167
rect 6574 4144 6578 4181
rect 6594 4179 6601 4216
rect 6594 4154 6601 4167
rect 6632 4164 6636 4221
rect 6640 4164 6644 4241
rect 6671 4233 6675 4276
rect 6648 4221 6655 4233
rect 6667 4221 6675 4233
rect 6648 4164 6652 4221
rect 6582 4148 6601 4154
rect 6582 4144 6586 4148
rect 43 4100 47 4104
rect 65 4100 69 4104
rect 125 4100 129 4104
rect 145 4100 149 4104
rect 165 4100 169 4104
rect 211 4100 215 4104
rect 231 4100 235 4104
rect 251 4100 255 4104
rect 315 4100 319 4104
rect 335 4100 339 4104
rect 345 4100 349 4104
rect 367 4100 371 4104
rect 377 4100 381 4104
rect 399 4100 403 4104
rect 445 4100 449 4104
rect 453 4100 457 4104
rect 473 4100 477 4104
rect 483 4100 487 4104
rect 505 4100 509 4104
rect 553 4100 557 4104
rect 563 4100 567 4104
rect 666 4100 670 4104
rect 674 4100 678 4104
rect 694 4100 698 4104
rect 702 4100 706 4104
rect 765 4100 769 4104
rect 811 4100 815 4104
rect 833 4100 837 4104
rect 843 4100 847 4104
rect 863 4100 867 4104
rect 871 4100 875 4104
rect 917 4100 921 4104
rect 939 4100 943 4104
rect 949 4100 953 4104
rect 971 4100 975 4104
rect 981 4100 985 4104
rect 1001 4100 1005 4104
rect 1053 4100 1057 4104
rect 1063 4100 1067 4104
rect 1131 4100 1135 4104
rect 1153 4100 1157 4104
rect 1163 4100 1167 4104
rect 1183 4100 1187 4104
rect 1191 4100 1195 4104
rect 1237 4100 1241 4104
rect 1259 4100 1263 4104
rect 1269 4100 1273 4104
rect 1291 4100 1295 4104
rect 1301 4100 1305 4104
rect 1321 4100 1325 4104
rect 1373 4100 1377 4104
rect 1383 4100 1387 4104
rect 1451 4100 1455 4104
rect 1525 4100 1529 4104
rect 1545 4100 1549 4104
rect 1565 4100 1569 4104
rect 1632 4100 1636 4104
rect 1654 4100 1658 4104
rect 1662 4100 1666 4104
rect 1733 4100 1737 4104
rect 1743 4100 1747 4104
rect 1793 4100 1797 4104
rect 1803 4100 1807 4104
rect 1871 4100 1875 4104
rect 1893 4100 1897 4104
rect 1903 4100 1907 4104
rect 1923 4100 1927 4104
rect 1931 4100 1935 4104
rect 1977 4100 1981 4104
rect 1999 4100 2003 4104
rect 2009 4100 2013 4104
rect 2031 4100 2035 4104
rect 2041 4100 2045 4104
rect 2061 4100 2065 4104
rect 2113 4100 2117 4104
rect 2123 4100 2127 4104
rect 2205 4100 2209 4104
rect 2225 4100 2229 4104
rect 2245 4100 2249 4104
rect 2295 4100 2299 4104
rect 2315 4100 2319 4104
rect 2325 4100 2329 4104
rect 2347 4100 2351 4104
rect 2357 4100 2361 4104
rect 2379 4100 2383 4104
rect 2425 4100 2429 4104
rect 2433 4100 2437 4104
rect 2453 4100 2457 4104
rect 2463 4100 2467 4104
rect 2485 4100 2489 4104
rect 2545 4100 2549 4104
rect 2565 4100 2569 4104
rect 2611 4100 2615 4104
rect 2671 4100 2675 4104
rect 2691 4100 2695 4104
rect 2711 4100 2715 4104
rect 2773 4100 2777 4104
rect 2783 4100 2787 4104
rect 2865 4100 2869 4104
rect 2885 4100 2889 4104
rect 2905 4100 2909 4104
rect 2951 4100 2955 4104
rect 3011 4100 3015 4104
rect 3031 4100 3035 4104
rect 3105 4100 3109 4104
rect 3151 4100 3155 4104
rect 3173 4100 3177 4104
rect 3183 4100 3187 4104
rect 3203 4100 3207 4104
rect 3211 4100 3215 4104
rect 3257 4100 3261 4104
rect 3279 4100 3283 4104
rect 3289 4100 3293 4104
rect 3311 4100 3315 4104
rect 3321 4100 3325 4104
rect 3341 4100 3345 4104
rect 3391 4100 3395 4104
rect 3411 4100 3415 4104
rect 3431 4100 3435 4104
rect 3451 4100 3455 4104
rect 3513 4100 3517 4104
rect 3523 4100 3527 4104
rect 3591 4100 3595 4104
rect 3611 4100 3615 4104
rect 3631 4100 3635 4104
rect 3651 4100 3655 4104
rect 3671 4100 3675 4104
rect 3691 4100 3695 4104
rect 3711 4100 3715 4104
rect 3731 4100 3735 4104
rect 3793 4100 3797 4104
rect 3803 4100 3807 4104
rect 3873 4100 3877 4104
rect 3883 4100 3887 4104
rect 3973 4100 3977 4104
rect 3983 4100 3987 4104
rect 4031 4100 4035 4104
rect 4105 4100 4109 4104
rect 4125 4100 4129 4104
rect 4145 4100 4149 4104
rect 4191 4100 4195 4104
rect 4211 4100 4215 4104
rect 4231 4100 4235 4104
rect 4295 4100 4299 4104
rect 4315 4100 4319 4104
rect 4325 4100 4329 4104
rect 4347 4100 4351 4104
rect 4357 4100 4361 4104
rect 4379 4100 4383 4104
rect 4425 4100 4429 4104
rect 4433 4100 4437 4104
rect 4453 4100 4457 4104
rect 4463 4100 4467 4104
rect 4485 4100 4489 4104
rect 4545 4100 4549 4104
rect 4565 4100 4569 4104
rect 4585 4100 4589 4104
rect 4635 4100 4639 4104
rect 4655 4100 4659 4104
rect 4665 4100 4669 4104
rect 4687 4100 4691 4104
rect 4697 4100 4701 4104
rect 4719 4100 4723 4104
rect 4765 4100 4769 4104
rect 4773 4100 4777 4104
rect 4793 4100 4797 4104
rect 4803 4100 4807 4104
rect 4825 4100 4829 4104
rect 4885 4100 4889 4104
rect 4952 4100 4956 4104
rect 4974 4100 4978 4104
rect 4982 4100 4986 4104
rect 5032 4100 5036 4104
rect 5040 4100 5044 4104
rect 5048 4100 5052 4104
rect 5145 4100 5149 4104
rect 5191 4100 5195 4104
rect 5211 4100 5215 4104
rect 5231 4100 5235 4104
rect 5295 4100 5299 4104
rect 5315 4100 5319 4104
rect 5325 4100 5329 4104
rect 5347 4100 5351 4104
rect 5357 4100 5361 4104
rect 5379 4100 5383 4104
rect 5425 4100 5429 4104
rect 5433 4100 5437 4104
rect 5453 4100 5457 4104
rect 5463 4100 5467 4104
rect 5485 4100 5489 4104
rect 5533 4100 5537 4104
rect 5543 4100 5547 4104
rect 5611 4100 5615 4104
rect 5671 4100 5675 4104
rect 5691 4100 5695 4104
rect 5711 4100 5715 4104
rect 5795 4100 5799 4104
rect 5815 4100 5819 4104
rect 5825 4100 5829 4104
rect 5872 4100 5876 4104
rect 5880 4100 5884 4104
rect 5888 4100 5892 4104
rect 5985 4100 5989 4104
rect 6031 4100 6035 4104
rect 6051 4100 6055 4104
rect 6071 4100 6075 4104
rect 6131 4100 6135 4104
rect 6153 4100 6157 4104
rect 6213 4100 6217 4104
rect 6223 4100 6227 4104
rect 6315 4100 6319 4104
rect 6335 4100 6339 4104
rect 6345 4100 6349 4104
rect 6393 4100 6397 4104
rect 6403 4100 6407 4104
rect 6471 4100 6475 4104
rect 6552 4100 6556 4104
rect 6574 4100 6578 4104
rect 6582 4100 6586 4104
rect 6632 4100 6636 4104
rect 6640 4100 6644 4104
rect 6648 4100 6652 4104
rect 43 4076 47 4080
rect 65 4076 69 4080
rect 111 4076 115 4080
rect 133 4076 137 4080
rect 143 4076 147 4080
rect 163 4076 167 4080
rect 171 4076 175 4080
rect 217 4076 221 4080
rect 239 4076 243 4080
rect 249 4076 253 4080
rect 271 4076 275 4080
rect 281 4076 285 4080
rect 301 4076 305 4080
rect 353 4076 357 4080
rect 363 4076 367 4080
rect 452 4076 456 4080
rect 474 4076 478 4080
rect 482 4076 486 4080
rect 553 4076 557 4080
rect 563 4076 567 4080
rect 633 4076 637 4080
rect 643 4076 647 4080
rect 703 4076 707 4080
rect 725 4076 729 4080
rect 771 4076 775 4080
rect 793 4076 797 4080
rect 803 4076 807 4080
rect 823 4076 827 4080
rect 831 4076 835 4080
rect 877 4076 881 4080
rect 899 4076 903 4080
rect 909 4076 913 4080
rect 931 4076 935 4080
rect 941 4076 945 4080
rect 961 4076 965 4080
rect 1033 4076 1037 4080
rect 1043 4076 1047 4080
rect 1093 4076 1097 4080
rect 1103 4076 1107 4080
rect 1173 4076 1177 4080
rect 1183 4076 1187 4080
rect 1272 4076 1276 4080
rect 1294 4076 1298 4080
rect 1302 4076 1306 4080
rect 1351 4076 1355 4080
rect 1373 4076 1377 4080
rect 1383 4076 1387 4080
rect 1403 4076 1407 4080
rect 1411 4076 1415 4080
rect 1457 4076 1461 4080
rect 1479 4076 1483 4080
rect 1489 4076 1493 4080
rect 1511 4076 1515 4080
rect 1521 4076 1525 4080
rect 1541 4076 1545 4080
rect 1613 4076 1617 4080
rect 1623 4076 1627 4080
rect 1671 4076 1675 4080
rect 1693 4076 1697 4080
rect 1753 4076 1757 4080
rect 1763 4076 1767 4080
rect 1831 4076 1835 4080
rect 1853 4076 1857 4080
rect 1863 4076 1867 4080
rect 1883 4076 1887 4080
rect 1891 4076 1895 4080
rect 1937 4076 1941 4080
rect 1959 4076 1963 4080
rect 1969 4076 1973 4080
rect 1991 4076 1995 4080
rect 2001 4076 2005 4080
rect 2021 4076 2025 4080
rect 2073 4076 2077 4080
rect 2083 4076 2087 4080
rect 2165 4076 2169 4080
rect 2185 4076 2189 4080
rect 2205 4076 2209 4080
rect 2273 4076 2277 4080
rect 2283 4076 2287 4080
rect 2333 4076 2337 4080
rect 2343 4076 2347 4080
rect 2425 4076 2429 4080
rect 2485 4076 2489 4080
rect 2505 4076 2509 4080
rect 2525 4076 2529 4080
rect 2571 4076 2575 4080
rect 2591 4076 2595 4080
rect 2665 4076 2669 4080
rect 2685 4076 2689 4080
rect 2731 4076 2735 4080
rect 2805 4076 2809 4080
rect 2873 4076 2877 4080
rect 2883 4076 2887 4080
rect 2931 4076 2935 4080
rect 2951 4076 2955 4080
rect 3011 4076 3015 4080
rect 3031 4076 3035 4080
rect 3051 4076 3055 4080
rect 3111 4076 3115 4080
rect 3171 4076 3175 4080
rect 3191 4076 3195 4080
rect 3273 4076 3277 4080
rect 3283 4076 3287 4080
rect 3353 4076 3357 4080
rect 3363 4076 3367 4080
rect 3415 4076 3419 4080
rect 3435 4076 3439 4080
rect 3445 4076 3449 4080
rect 3467 4076 3471 4080
rect 3477 4076 3481 4080
rect 3499 4076 3503 4080
rect 3545 4076 3549 4080
rect 3553 4076 3557 4080
rect 3573 4076 3577 4080
rect 3583 4076 3587 4080
rect 3605 4076 3609 4080
rect 3665 4076 3669 4080
rect 3715 4076 3719 4080
rect 3735 4076 3739 4080
rect 3745 4076 3749 4080
rect 3767 4076 3771 4080
rect 3777 4076 3781 4080
rect 3799 4076 3803 4080
rect 3845 4076 3849 4080
rect 3853 4076 3857 4080
rect 3873 4076 3877 4080
rect 3883 4076 3887 4080
rect 3905 4076 3909 4080
rect 3988 4076 3992 4080
rect 3996 4076 4000 4080
rect 4004 4076 4008 4080
rect 4053 4076 4057 4080
rect 4063 4076 4067 4080
rect 4145 4076 4149 4080
rect 4165 4076 4169 4080
rect 4185 4076 4189 4080
rect 4231 4076 4235 4080
rect 4251 4076 4255 4080
rect 4325 4076 4329 4080
rect 4393 4076 4397 4080
rect 4403 4076 4407 4080
rect 4465 4076 4469 4080
rect 4485 4076 4489 4080
rect 4505 4076 4509 4080
rect 4555 4076 4559 4080
rect 4575 4076 4579 4080
rect 4585 4076 4589 4080
rect 4607 4076 4611 4080
rect 4617 4076 4621 4080
rect 4639 4076 4643 4080
rect 4685 4076 4689 4080
rect 4693 4076 4697 4080
rect 4713 4076 4717 4080
rect 4723 4076 4727 4080
rect 4745 4076 4749 4080
rect 4813 4076 4817 4080
rect 4823 4076 4827 4080
rect 4885 4076 4889 4080
rect 4905 4076 4909 4080
rect 4925 4076 4929 4080
rect 4975 4076 4979 4080
rect 4995 4076 4999 4080
rect 5005 4076 5009 4080
rect 5027 4076 5031 4080
rect 5037 4076 5041 4080
rect 5059 4076 5063 4080
rect 5105 4076 5109 4080
rect 5113 4076 5117 4080
rect 5133 4076 5137 4080
rect 5143 4076 5147 4080
rect 5165 4076 5169 4080
rect 5233 4076 5237 4080
rect 5243 4076 5247 4080
rect 5305 4076 5309 4080
rect 5325 4076 5329 4080
rect 5345 4076 5349 4080
rect 5413 4076 5417 4080
rect 5423 4076 5427 4080
rect 5471 4076 5475 4080
rect 5491 4076 5495 4080
rect 5511 4076 5515 4080
rect 5585 4076 5589 4080
rect 5635 4076 5639 4080
rect 5655 4076 5659 4080
rect 5665 4076 5669 4080
rect 5687 4076 5691 4080
rect 5697 4076 5701 4080
rect 5719 4076 5723 4080
rect 5765 4076 5769 4080
rect 5773 4076 5777 4080
rect 5793 4076 5797 4080
rect 5803 4076 5807 4080
rect 5825 4076 5829 4080
rect 5871 4076 5875 4080
rect 5968 4076 5972 4080
rect 5976 4076 5980 4080
rect 5984 4076 5988 4080
rect 6031 4076 6035 4080
rect 6053 4076 6057 4080
rect 6063 4076 6067 4080
rect 6083 4076 6087 4080
rect 6091 4076 6095 4080
rect 6137 4076 6141 4080
rect 6159 4076 6163 4080
rect 6169 4076 6173 4080
rect 6191 4076 6195 4080
rect 6201 4076 6205 4080
rect 6221 4076 6225 4080
rect 6271 4076 6275 4080
rect 6293 4076 6297 4080
rect 6303 4076 6307 4080
rect 6323 4076 6327 4080
rect 6331 4076 6335 4080
rect 6377 4076 6381 4080
rect 6399 4076 6403 4080
rect 6409 4076 6413 4080
rect 6431 4076 6435 4080
rect 6441 4076 6445 4080
rect 6461 4076 6465 4080
rect 6511 4076 6515 4080
rect 6533 4076 6537 4080
rect 6543 4076 6547 4080
rect 6563 4076 6567 4080
rect 6571 4076 6575 4080
rect 6617 4076 6621 4080
rect 6639 4076 6643 4080
rect 6649 4076 6653 4080
rect 6671 4076 6675 4080
rect 6681 4076 6685 4080
rect 6701 4076 6705 4080
rect 43 4030 47 4036
rect 43 4018 45 4030
rect 65 3979 69 4056
rect 65 3967 74 3979
rect 111 3968 115 4036
rect 133 4007 137 4056
rect 143 4035 147 4056
rect 163 4044 167 4056
rect 171 4052 175 4056
rect 171 4048 205 4052
rect 163 4040 193 4044
rect 163 4039 181 4040
rect 143 4031 167 4035
rect 43 3950 45 3962
rect 43 3944 47 3950
rect 65 3904 69 3967
rect 111 3956 113 3968
rect 111 3944 115 3956
rect 133 3949 137 3995
rect 129 3943 137 3949
rect 129 3914 133 3943
rect 161 3936 167 4031
rect 129 3907 137 3914
rect 133 3884 137 3907
rect 141 3884 145 3924
rect 161 3904 165 3936
rect 201 3922 205 4048
rect 217 3942 221 4056
rect 239 4044 243 4056
rect 241 4032 243 4044
rect 249 4044 253 4056
rect 249 4032 251 4044
rect 169 3910 193 3912
rect 169 3908 205 3910
rect 169 3904 173 3908
rect 215 3904 219 3930
rect 233 3922 237 4032
rect 271 4024 275 4056
rect 242 4020 275 4024
rect 242 3956 246 4020
rect 262 3971 266 4000
rect 281 3998 285 4056
rect 301 3999 305 4036
rect 353 4016 357 4036
rect 349 4009 357 4016
rect 363 4016 367 4036
rect 363 4009 377 4016
rect 452 4013 456 4056
rect 349 3993 355 4009
rect 262 3963 271 3971
rect 242 3944 245 3956
rect 235 3904 239 3910
rect 247 3904 251 3944
rect 267 3904 271 3963
rect 281 3904 285 3986
rect 301 3944 305 3987
rect 346 3981 355 3993
rect 351 3904 355 3981
rect 371 3993 377 4009
rect 445 4001 454 4013
rect 371 3981 374 3993
rect 371 3904 375 3981
rect 445 3944 449 4001
rect 474 3999 478 4036
rect 482 4032 486 4036
rect 482 4026 501 4032
rect 494 4013 501 4026
rect 553 4016 557 4036
rect 543 4009 557 4016
rect 563 4016 567 4036
rect 633 4016 637 4036
rect 563 4009 571 4016
rect 474 3964 480 3987
rect 494 3964 501 4001
rect 543 3993 549 4009
rect 546 3981 549 3993
rect 465 3958 480 3964
rect 485 3958 501 3964
rect 465 3944 469 3958
rect 485 3944 489 3958
rect 545 3904 549 3981
rect 565 3993 571 4009
rect 623 4009 637 4016
rect 643 4016 647 4036
rect 703 4030 707 4036
rect 703 4018 705 4030
rect 643 4009 651 4016
rect 623 3993 629 4009
rect 565 3981 574 3993
rect 626 3981 629 3993
rect 565 3904 569 3981
rect 625 3904 629 3981
rect 645 3993 651 4009
rect 645 3981 654 3993
rect 645 3904 649 3981
rect 725 3979 729 4056
rect 725 3967 734 3979
rect 771 3968 775 4036
rect 793 4007 797 4056
rect 803 4035 807 4056
rect 823 4044 827 4056
rect 831 4052 835 4056
rect 831 4048 865 4052
rect 823 4040 853 4044
rect 823 4039 841 4040
rect 803 4031 827 4035
rect 703 3950 705 3962
rect 703 3944 707 3950
rect 725 3904 729 3967
rect 771 3956 773 3968
rect 771 3944 775 3956
rect 793 3949 797 3995
rect 789 3943 797 3949
rect 789 3914 793 3943
rect 821 3936 827 4031
rect 789 3907 797 3914
rect 793 3884 797 3907
rect 801 3884 805 3924
rect 821 3904 825 3936
rect 861 3922 865 4048
rect 877 3942 881 4056
rect 899 4044 903 4056
rect 901 4032 903 4044
rect 909 4044 913 4056
rect 909 4032 911 4044
rect 829 3910 853 3912
rect 829 3908 865 3910
rect 829 3904 833 3908
rect 875 3904 879 3930
rect 893 3922 897 4032
rect 931 4024 935 4056
rect 902 4020 935 4024
rect 902 3956 906 4020
rect 922 3971 926 4000
rect 941 3998 945 4056
rect 961 3999 965 4036
rect 1033 4016 1037 4036
rect 1023 4009 1037 4016
rect 1043 4016 1047 4036
rect 1093 4016 1097 4036
rect 1043 4009 1051 4016
rect 1023 3993 1029 4009
rect 922 3963 931 3971
rect 902 3944 905 3956
rect 895 3904 899 3910
rect 907 3904 911 3944
rect 927 3904 931 3963
rect 941 3904 945 3986
rect 961 3944 965 3987
rect 1026 3981 1029 3993
rect 1025 3904 1029 3981
rect 1045 3993 1051 4009
rect 1089 4009 1097 4016
rect 1103 4016 1107 4036
rect 1173 4016 1177 4036
rect 1103 4009 1117 4016
rect 1089 3993 1095 4009
rect 1045 3981 1054 3993
rect 1086 3981 1095 3993
rect 1045 3904 1049 3981
rect 1091 3904 1095 3981
rect 1111 3993 1117 4009
rect 1169 4009 1177 4016
rect 1183 4016 1187 4036
rect 1183 4009 1197 4016
rect 1272 4013 1276 4056
rect 1169 3993 1175 4009
rect 1111 3981 1114 3993
rect 1166 3981 1175 3993
rect 1111 3904 1115 3981
rect 1171 3904 1175 3981
rect 1191 3993 1197 4009
rect 1265 4001 1274 4013
rect 1191 3981 1194 3993
rect 1191 3904 1195 3981
rect 1265 3944 1269 4001
rect 1294 3999 1298 4036
rect 1302 4032 1306 4036
rect 1302 4026 1321 4032
rect 1314 4013 1321 4026
rect 1294 3964 1300 3987
rect 1314 3964 1321 4001
rect 1285 3958 1300 3964
rect 1305 3958 1321 3964
rect 1351 3968 1355 4036
rect 1373 4007 1377 4056
rect 1383 4035 1387 4056
rect 1403 4044 1407 4056
rect 1411 4052 1415 4056
rect 1411 4048 1445 4052
rect 1403 4040 1433 4044
rect 1403 4039 1421 4040
rect 1383 4031 1407 4035
rect 1285 3944 1289 3958
rect 1305 3944 1309 3958
rect 1351 3956 1353 3968
rect 1351 3944 1355 3956
rect 1373 3949 1377 3995
rect 1369 3943 1377 3949
rect 1369 3914 1373 3943
rect 1401 3936 1407 4031
rect 1369 3907 1377 3914
rect 1373 3884 1377 3907
rect 1381 3884 1385 3924
rect 1401 3904 1405 3936
rect 1441 3922 1445 4048
rect 1457 3942 1461 4056
rect 1479 4044 1483 4056
rect 1481 4032 1483 4044
rect 1489 4044 1493 4056
rect 1489 4032 1491 4044
rect 1409 3910 1433 3912
rect 1409 3908 1445 3910
rect 1409 3904 1413 3908
rect 1455 3904 1459 3930
rect 1473 3922 1477 4032
rect 1511 4024 1515 4056
rect 1482 4020 1515 4024
rect 1482 3956 1486 4020
rect 1502 3971 1506 4000
rect 1521 3998 1525 4056
rect 1541 3999 1545 4036
rect 1613 4016 1617 4036
rect 1603 4009 1617 4016
rect 1623 4016 1627 4036
rect 1623 4009 1631 4016
rect 1603 3993 1609 4009
rect 1502 3963 1511 3971
rect 1482 3944 1485 3956
rect 1475 3904 1479 3910
rect 1487 3904 1491 3944
rect 1507 3904 1511 3963
rect 1521 3904 1525 3986
rect 1541 3944 1545 3987
rect 1606 3981 1609 3993
rect 1605 3904 1609 3981
rect 1625 3993 1631 4009
rect 1625 3981 1634 3993
rect 1625 3904 1629 3981
rect 1671 3979 1675 4056
rect 1693 4030 1697 4036
rect 1695 4018 1697 4030
rect 1753 4016 1757 4036
rect 1749 4009 1757 4016
rect 1763 4016 1767 4036
rect 1763 4009 1777 4016
rect 1749 3993 1755 4009
rect 1746 3981 1755 3993
rect 1666 3967 1675 3979
rect 1671 3904 1675 3967
rect 1695 3950 1697 3962
rect 1693 3944 1697 3950
rect 1751 3904 1755 3981
rect 1771 3993 1777 4009
rect 1771 3981 1774 3993
rect 1771 3904 1775 3981
rect 1831 3968 1835 4036
rect 1853 4007 1857 4056
rect 1863 4035 1867 4056
rect 1883 4044 1887 4056
rect 1891 4052 1895 4056
rect 1891 4048 1925 4052
rect 1883 4040 1913 4044
rect 1883 4039 1901 4040
rect 1863 4031 1887 4035
rect 1831 3956 1833 3968
rect 1831 3944 1835 3956
rect 1853 3949 1857 3995
rect 1849 3943 1857 3949
rect 1849 3914 1853 3943
rect 1881 3936 1887 4031
rect 1849 3907 1857 3914
rect 1853 3884 1857 3907
rect 1861 3884 1865 3924
rect 1881 3904 1885 3936
rect 1921 3922 1925 4048
rect 1937 3942 1941 4056
rect 1959 4044 1963 4056
rect 1961 4032 1963 4044
rect 1969 4044 1973 4056
rect 1969 4032 1971 4044
rect 1889 3910 1913 3912
rect 1889 3908 1925 3910
rect 1889 3904 1893 3908
rect 1935 3904 1939 3930
rect 1953 3922 1957 4032
rect 1991 4024 1995 4056
rect 1962 4020 1995 4024
rect 1962 3956 1966 4020
rect 1982 3971 1986 4000
rect 2001 3998 2005 4056
rect 2021 3999 2025 4036
rect 2073 4016 2077 4036
rect 2069 4009 2077 4016
rect 2083 4016 2087 4036
rect 2083 4009 2097 4016
rect 2069 3993 2075 4009
rect 1982 3963 1991 3971
rect 1962 3944 1965 3956
rect 1955 3904 1959 3910
rect 1967 3904 1971 3944
rect 1987 3904 1991 3963
rect 2001 3904 2005 3986
rect 2021 3944 2025 3987
rect 2066 3981 2075 3993
rect 2071 3904 2075 3981
rect 2091 3993 2097 4009
rect 2091 3981 2094 3993
rect 2091 3904 2095 3981
rect 2165 3959 2169 4036
rect 2185 4013 2189 4036
rect 2205 4031 2209 4036
rect 2205 4024 2218 4031
rect 2185 4001 2194 4013
rect 2167 3947 2174 3959
rect 2170 3904 2174 3947
rect 2192 3944 2196 4001
rect 2214 3979 2218 4024
rect 2273 4016 2277 4036
rect 2263 4009 2277 4016
rect 2283 4016 2287 4036
rect 2333 4016 2337 4036
rect 2283 4009 2291 4016
rect 2263 3993 2269 4009
rect 2266 3981 2269 3993
rect 2214 3956 2218 3967
rect 2200 3948 2218 3956
rect 2200 3944 2204 3948
rect 2265 3904 2269 3981
rect 2285 3993 2291 4009
rect 2329 4009 2337 4016
rect 2343 4016 2347 4036
rect 2343 4009 2357 4016
rect 2329 3993 2335 4009
rect 2285 3981 2294 3993
rect 2326 3981 2335 3993
rect 2285 3904 2289 3981
rect 2331 3904 2335 3981
rect 2351 3993 2357 4009
rect 2425 3999 2429 4056
rect 2351 3981 2354 3993
rect 2425 3987 2434 3999
rect 2351 3904 2355 3981
rect 2425 3904 2429 3987
rect 2485 3959 2489 4036
rect 2505 4013 2509 4036
rect 2525 4031 2529 4036
rect 2525 4024 2538 4031
rect 2505 4001 2514 4013
rect 2487 3947 2494 3959
rect 2490 3904 2494 3947
rect 2512 3944 2516 4001
rect 2534 3979 2538 4024
rect 2571 3979 2575 4056
rect 2591 3979 2595 4056
rect 2665 3979 2669 4056
rect 2685 3979 2689 4056
rect 2731 3999 2735 4056
rect 2726 3987 2735 3999
rect 2566 3967 2575 3979
rect 2534 3956 2538 3967
rect 2520 3948 2538 3956
rect 2520 3944 2524 3948
rect 2571 3944 2575 3967
rect 2579 3967 2594 3979
rect 2666 3967 2681 3979
rect 2579 3944 2583 3967
rect 2677 3944 2681 3967
rect 2685 3967 2694 3979
rect 2685 3944 2689 3967
rect 2731 3904 2735 3987
rect 2805 3999 2809 4056
rect 2873 4016 2877 4036
rect 2863 4009 2877 4016
rect 2883 4016 2887 4036
rect 2883 4009 2891 4016
rect 2805 3987 2814 3999
rect 2863 3993 2869 4009
rect 2805 3904 2809 3987
rect 2866 3981 2869 3993
rect 2865 3904 2869 3981
rect 2885 3993 2891 4009
rect 2885 3981 2894 3993
rect 2885 3904 2889 3981
rect 2931 3979 2935 4056
rect 2951 3979 2955 4056
rect 3011 4031 3015 4036
rect 3002 4024 3015 4031
rect 3002 3979 3006 4024
rect 3031 4013 3035 4036
rect 3026 4001 3035 4013
rect 2926 3967 2935 3979
rect 2931 3944 2935 3967
rect 2939 3967 2954 3979
rect 2939 3944 2943 3967
rect 3002 3956 3006 3967
rect 3002 3948 3020 3956
rect 3016 3944 3020 3948
rect 3024 3944 3028 4001
rect 3051 3959 3055 4036
rect 3111 3999 3115 4056
rect 3106 3987 3115 3999
rect 3046 3947 3053 3959
rect 3046 3904 3050 3947
rect 3111 3904 3115 3987
rect 3171 3979 3175 4056
rect 3191 3979 3195 4056
rect 3273 4016 3277 4036
rect 3263 4009 3277 4016
rect 3283 4016 3287 4036
rect 3353 4016 3357 4036
rect 3283 4009 3291 4016
rect 3263 3993 3269 4009
rect 3266 3981 3269 3993
rect 3166 3967 3175 3979
rect 3171 3944 3175 3967
rect 3179 3967 3194 3979
rect 3179 3944 3183 3967
rect 3265 3904 3269 3981
rect 3285 3993 3291 4009
rect 3343 4009 3357 4016
rect 3363 4016 3367 4036
rect 3363 4009 3371 4016
rect 3343 3993 3349 4009
rect 3285 3981 3294 3993
rect 3346 3981 3349 3993
rect 3285 3904 3289 3981
rect 3345 3904 3349 3981
rect 3365 3993 3371 4009
rect 3415 3999 3419 4036
rect 3365 3981 3374 3993
rect 3435 3998 3439 4056
rect 3445 4024 3449 4056
rect 3467 4044 3471 4056
rect 3469 4032 3471 4044
rect 3477 4044 3481 4056
rect 3477 4032 3479 4044
rect 3445 4020 3478 4024
rect 3365 3904 3369 3981
rect 3415 3944 3419 3987
rect 3435 3904 3439 3986
rect 3454 3971 3458 4000
rect 3449 3963 3458 3971
rect 3449 3904 3453 3963
rect 3474 3956 3478 4020
rect 3475 3944 3478 3956
rect 3469 3904 3473 3944
rect 3483 3922 3487 4032
rect 3499 3942 3503 4056
rect 3545 4052 3549 4056
rect 3515 4048 3549 4052
rect 3481 3904 3485 3910
rect 3501 3904 3505 3930
rect 3515 3922 3519 4048
rect 3553 4044 3557 4056
rect 3527 4040 3557 4044
rect 3539 4039 3557 4040
rect 3573 4035 3577 4056
rect 3553 4031 3577 4035
rect 3553 3936 3559 4031
rect 3583 4007 3587 4056
rect 3583 3949 3587 3995
rect 3605 3968 3609 4036
rect 3607 3956 3609 3968
rect 3583 3943 3591 3949
rect 3605 3944 3609 3956
rect 3665 3999 3669 4056
rect 3715 3999 3719 4036
rect 3665 3987 3674 3999
rect 3735 3998 3739 4056
rect 3745 4024 3749 4056
rect 3767 4044 3771 4056
rect 3769 4032 3771 4044
rect 3777 4044 3781 4056
rect 3777 4032 3779 4044
rect 3745 4020 3778 4024
rect 3527 3910 3551 3912
rect 3515 3908 3551 3910
rect 3547 3904 3551 3908
rect 3555 3904 3559 3936
rect 3575 3884 3579 3924
rect 3587 3914 3591 3943
rect 3583 3907 3591 3914
rect 3583 3884 3587 3907
rect 3665 3904 3669 3987
rect 3715 3944 3719 3987
rect 3735 3904 3739 3986
rect 3754 3971 3758 4000
rect 3749 3963 3758 3971
rect 3749 3904 3753 3963
rect 3774 3956 3778 4020
rect 3775 3944 3778 3956
rect 3769 3904 3773 3944
rect 3783 3922 3787 4032
rect 3799 3942 3803 4056
rect 3845 4052 3849 4056
rect 3815 4048 3849 4052
rect 3781 3904 3785 3910
rect 3801 3904 3805 3930
rect 3815 3922 3819 4048
rect 3853 4044 3857 4056
rect 3827 4040 3857 4044
rect 3839 4039 3857 4040
rect 3873 4035 3877 4056
rect 3853 4031 3877 4035
rect 3853 3936 3859 4031
rect 3883 4007 3887 4056
rect 3883 3949 3887 3995
rect 3905 3968 3909 4036
rect 4053 4016 4057 4036
rect 3907 3956 3909 3968
rect 3988 3959 3992 4016
rect 3883 3943 3891 3949
rect 3905 3944 3909 3956
rect 3965 3947 3973 3959
rect 3985 3947 3992 3959
rect 3827 3910 3851 3912
rect 3815 3908 3851 3910
rect 3847 3904 3851 3908
rect 3855 3904 3859 3936
rect 3875 3884 3879 3924
rect 3887 3914 3891 3943
rect 3883 3907 3891 3914
rect 3883 3884 3887 3907
rect 3965 3904 3969 3947
rect 3996 3939 4000 4016
rect 4004 3959 4008 4016
rect 4049 4009 4057 4016
rect 4063 4016 4067 4036
rect 4063 4009 4077 4016
rect 4049 3993 4055 4009
rect 4046 3981 4055 3993
rect 4004 3947 4014 3959
rect 3994 3920 4000 3927
rect 3985 3916 4000 3920
rect 4014 3916 4020 3947
rect 3985 3904 3989 3916
rect 4005 3912 4020 3916
rect 4005 3904 4009 3912
rect 4051 3904 4055 3981
rect 4071 3993 4077 4009
rect 4071 3981 4074 3993
rect 4071 3904 4075 3981
rect 4145 3959 4149 4036
rect 4165 4013 4169 4036
rect 4185 4031 4189 4036
rect 4185 4024 4198 4031
rect 4165 4001 4174 4013
rect 4147 3947 4154 3959
rect 4150 3904 4154 3947
rect 4172 3944 4176 4001
rect 4194 3979 4198 4024
rect 4231 3979 4235 4056
rect 4251 3979 4255 4056
rect 4325 3999 4329 4056
rect 4393 4016 4397 4036
rect 4383 4009 4397 4016
rect 4403 4016 4407 4036
rect 4403 4009 4411 4016
rect 4325 3987 4334 3999
rect 4383 3993 4389 4009
rect 4226 3967 4235 3979
rect 4194 3956 4198 3967
rect 4180 3948 4198 3956
rect 4180 3944 4184 3948
rect 4231 3944 4235 3967
rect 4239 3967 4254 3979
rect 4239 3944 4243 3967
rect 4325 3904 4329 3987
rect 4386 3981 4389 3993
rect 4385 3904 4389 3981
rect 4405 3993 4411 4009
rect 4405 3981 4414 3993
rect 4405 3904 4409 3981
rect 4465 3959 4469 4036
rect 4485 4013 4489 4036
rect 4505 4031 4509 4036
rect 4505 4024 4518 4031
rect 4485 4001 4494 4013
rect 4467 3947 4474 3959
rect 4470 3904 4474 3947
rect 4492 3944 4496 4001
rect 4514 3979 4518 4024
rect 4555 3999 4559 4036
rect 4575 3998 4579 4056
rect 4585 4024 4589 4056
rect 4607 4044 4611 4056
rect 4609 4032 4611 4044
rect 4617 4044 4621 4056
rect 4617 4032 4619 4044
rect 4585 4020 4618 4024
rect 4514 3956 4518 3967
rect 4500 3948 4518 3956
rect 4500 3944 4504 3948
rect 4555 3944 4559 3987
rect 4575 3904 4579 3986
rect 4594 3971 4598 4000
rect 4589 3963 4598 3971
rect 4589 3904 4593 3963
rect 4614 3956 4618 4020
rect 4615 3944 4618 3956
rect 4609 3904 4613 3944
rect 4623 3922 4627 4032
rect 4639 3942 4643 4056
rect 4685 4052 4689 4056
rect 4655 4048 4689 4052
rect 4621 3904 4625 3910
rect 4641 3904 4645 3930
rect 4655 3922 4659 4048
rect 4693 4044 4697 4056
rect 4667 4040 4697 4044
rect 4679 4039 4697 4040
rect 4713 4035 4717 4056
rect 4693 4031 4717 4035
rect 4693 3936 4699 4031
rect 4723 4007 4727 4056
rect 4723 3949 4727 3995
rect 4745 3968 4749 4036
rect 4813 4016 4817 4036
rect 4803 4009 4817 4016
rect 4823 4016 4827 4036
rect 4823 4009 4831 4016
rect 4803 3993 4809 4009
rect 4806 3981 4809 3993
rect 4747 3956 4749 3968
rect 4723 3943 4731 3949
rect 4745 3944 4749 3956
rect 4667 3910 4691 3912
rect 4655 3908 4691 3910
rect 4687 3904 4691 3908
rect 4695 3904 4699 3936
rect 4715 3884 4719 3924
rect 4727 3914 4731 3943
rect 4723 3907 4731 3914
rect 4723 3884 4727 3907
rect 4805 3904 4809 3981
rect 4825 3993 4831 4009
rect 4825 3981 4834 3993
rect 4825 3904 4829 3981
rect 4885 3959 4889 4036
rect 4905 4013 4909 4036
rect 4925 4031 4929 4036
rect 4925 4024 4938 4031
rect 4905 4001 4914 4013
rect 4887 3947 4894 3959
rect 4890 3904 4894 3947
rect 4912 3944 4916 4001
rect 4934 3979 4938 4024
rect 4975 3999 4979 4036
rect 4995 3998 4999 4056
rect 5005 4024 5009 4056
rect 5027 4044 5031 4056
rect 5029 4032 5031 4044
rect 5037 4044 5041 4056
rect 5037 4032 5039 4044
rect 5005 4020 5038 4024
rect 4934 3956 4938 3967
rect 4920 3948 4938 3956
rect 4920 3944 4924 3948
rect 4975 3944 4979 3987
rect 4995 3904 4999 3986
rect 5014 3971 5018 4000
rect 5009 3963 5018 3971
rect 5009 3904 5013 3963
rect 5034 3956 5038 4020
rect 5035 3944 5038 3956
rect 5029 3904 5033 3944
rect 5043 3922 5047 4032
rect 5059 3942 5063 4056
rect 5105 4052 5109 4056
rect 5075 4048 5109 4052
rect 5041 3904 5045 3910
rect 5061 3904 5065 3930
rect 5075 3922 5079 4048
rect 5113 4044 5117 4056
rect 5087 4040 5117 4044
rect 5099 4039 5117 4040
rect 5133 4035 5137 4056
rect 5113 4031 5137 4035
rect 5113 3936 5119 4031
rect 5143 4007 5147 4056
rect 5143 3949 5147 3995
rect 5165 3968 5169 4036
rect 5233 4016 5237 4036
rect 5223 4009 5237 4016
rect 5243 4016 5247 4036
rect 5243 4009 5251 4016
rect 5223 3993 5229 4009
rect 5226 3981 5229 3993
rect 5167 3956 5169 3968
rect 5143 3943 5151 3949
rect 5165 3944 5169 3956
rect 5087 3910 5111 3912
rect 5075 3908 5111 3910
rect 5107 3904 5111 3908
rect 5115 3904 5119 3936
rect 5135 3884 5139 3924
rect 5147 3914 5151 3943
rect 5143 3907 5151 3914
rect 5143 3884 5147 3907
rect 5225 3904 5229 3981
rect 5245 3993 5251 4009
rect 5245 3981 5254 3993
rect 5245 3904 5249 3981
rect 5305 3959 5309 4036
rect 5325 4013 5329 4036
rect 5345 4031 5349 4036
rect 5345 4024 5358 4031
rect 5325 4001 5334 4013
rect 5307 3947 5314 3959
rect 5310 3904 5314 3947
rect 5332 3944 5336 4001
rect 5354 3979 5358 4024
rect 5413 4016 5417 4036
rect 5403 4009 5417 4016
rect 5423 4016 5427 4036
rect 5471 4031 5475 4036
rect 5462 4024 5475 4031
rect 5423 4009 5431 4016
rect 5403 3993 5409 4009
rect 5406 3981 5409 3993
rect 5354 3956 5358 3967
rect 5340 3948 5358 3956
rect 5340 3944 5344 3948
rect 5405 3904 5409 3981
rect 5425 3993 5431 4009
rect 5425 3981 5434 3993
rect 5425 3904 5429 3981
rect 5462 3979 5466 4024
rect 5491 4013 5495 4036
rect 5486 4001 5495 4013
rect 5462 3956 5466 3967
rect 5462 3948 5480 3956
rect 5476 3944 5480 3948
rect 5484 3944 5488 4001
rect 5511 3959 5515 4036
rect 5585 3999 5589 4056
rect 5635 3999 5639 4036
rect 5585 3987 5594 3999
rect 5655 3998 5659 4056
rect 5665 4024 5669 4056
rect 5687 4044 5691 4056
rect 5689 4032 5691 4044
rect 5697 4044 5701 4056
rect 5697 4032 5699 4044
rect 5665 4020 5698 4024
rect 5506 3947 5513 3959
rect 5506 3904 5510 3947
rect 5585 3904 5589 3987
rect 5635 3944 5639 3987
rect 5655 3904 5659 3986
rect 5674 3971 5678 4000
rect 5669 3963 5678 3971
rect 5669 3904 5673 3963
rect 5694 3956 5698 4020
rect 5695 3944 5698 3956
rect 5689 3904 5693 3944
rect 5703 3922 5707 4032
rect 5719 3942 5723 4056
rect 5765 4052 5769 4056
rect 5735 4048 5769 4052
rect 5701 3904 5705 3910
rect 5721 3904 5725 3930
rect 5735 3922 5739 4048
rect 5773 4044 5777 4056
rect 5747 4040 5777 4044
rect 5759 4039 5777 4040
rect 5793 4035 5797 4056
rect 5773 4031 5797 4035
rect 5773 3936 5779 4031
rect 5803 4007 5807 4056
rect 5803 3949 5807 3995
rect 5825 3968 5829 4036
rect 5871 3999 5875 4056
rect 5866 3987 5875 3999
rect 5827 3956 5829 3968
rect 5803 3943 5811 3949
rect 5825 3944 5829 3956
rect 5747 3910 5771 3912
rect 5735 3908 5771 3910
rect 5767 3904 5771 3908
rect 5775 3904 5779 3936
rect 5795 3884 5799 3924
rect 5807 3914 5811 3943
rect 5803 3907 5811 3914
rect 5803 3884 5807 3907
rect 5871 3904 5875 3987
rect 5968 3959 5972 4016
rect 5945 3947 5953 3959
rect 5965 3947 5972 3959
rect 5945 3904 5949 3947
rect 5976 3939 5980 4016
rect 5984 3959 5988 4016
rect 6031 3968 6035 4036
rect 6053 4007 6057 4056
rect 6063 4035 6067 4056
rect 6083 4044 6087 4056
rect 6091 4052 6095 4056
rect 6091 4048 6125 4052
rect 6083 4040 6113 4044
rect 6083 4039 6101 4040
rect 6063 4031 6087 4035
rect 5984 3947 5994 3959
rect 6031 3956 6033 3968
rect 5974 3920 5980 3927
rect 5965 3916 5980 3920
rect 5994 3916 6000 3947
rect 6031 3944 6035 3956
rect 6053 3949 6057 3995
rect 5965 3904 5969 3916
rect 5985 3912 6000 3916
rect 5985 3904 5989 3912
rect 6049 3943 6057 3949
rect 6049 3914 6053 3943
rect 6081 3936 6087 4031
rect 6049 3907 6057 3914
rect 6053 3884 6057 3907
rect 6061 3884 6065 3924
rect 6081 3904 6085 3936
rect 6121 3922 6125 4048
rect 6137 3942 6141 4056
rect 6159 4044 6163 4056
rect 6161 4032 6163 4044
rect 6169 4044 6173 4056
rect 6169 4032 6171 4044
rect 6089 3910 6113 3912
rect 6089 3908 6125 3910
rect 6089 3904 6093 3908
rect 6135 3904 6139 3930
rect 6153 3922 6157 4032
rect 6191 4024 6195 4056
rect 6162 4020 6195 4024
rect 6162 3956 6166 4020
rect 6182 3971 6186 4000
rect 6201 3998 6205 4056
rect 6221 3999 6225 4036
rect 6182 3963 6191 3971
rect 6162 3944 6165 3956
rect 6155 3904 6159 3910
rect 6167 3904 6171 3944
rect 6187 3904 6191 3963
rect 6201 3904 6205 3986
rect 6221 3944 6225 3987
rect 6271 3968 6275 4036
rect 6293 4007 6297 4056
rect 6303 4035 6307 4056
rect 6323 4044 6327 4056
rect 6331 4052 6335 4056
rect 6331 4048 6365 4052
rect 6323 4040 6353 4044
rect 6323 4039 6341 4040
rect 6303 4031 6327 4035
rect 6271 3956 6273 3968
rect 6271 3944 6275 3956
rect 6293 3949 6297 3995
rect 6289 3943 6297 3949
rect 6289 3914 6293 3943
rect 6321 3936 6327 4031
rect 6289 3907 6297 3914
rect 6293 3884 6297 3907
rect 6301 3884 6305 3924
rect 6321 3904 6325 3936
rect 6361 3922 6365 4048
rect 6377 3942 6381 4056
rect 6399 4044 6403 4056
rect 6401 4032 6403 4044
rect 6409 4044 6413 4056
rect 6409 4032 6411 4044
rect 6329 3910 6353 3912
rect 6329 3908 6365 3910
rect 6329 3904 6333 3908
rect 6375 3904 6379 3930
rect 6393 3922 6397 4032
rect 6431 4024 6435 4056
rect 6402 4020 6435 4024
rect 6402 3956 6406 4020
rect 6422 3971 6426 4000
rect 6441 3998 6445 4056
rect 6461 3999 6465 4036
rect 6422 3963 6431 3971
rect 6402 3944 6405 3956
rect 6395 3904 6399 3910
rect 6407 3904 6411 3944
rect 6427 3904 6431 3963
rect 6441 3904 6445 3986
rect 6461 3944 6465 3987
rect 6511 3968 6515 4036
rect 6533 4007 6537 4056
rect 6543 4035 6547 4056
rect 6563 4044 6567 4056
rect 6571 4052 6575 4056
rect 6571 4048 6605 4052
rect 6563 4040 6593 4044
rect 6563 4039 6581 4040
rect 6543 4031 6567 4035
rect 6511 3956 6513 3968
rect 6511 3944 6515 3956
rect 6533 3949 6537 3995
rect 6529 3943 6537 3949
rect 6529 3914 6533 3943
rect 6561 3936 6567 4031
rect 6529 3907 6537 3914
rect 6533 3884 6537 3907
rect 6541 3884 6545 3924
rect 6561 3904 6565 3936
rect 6601 3922 6605 4048
rect 6617 3942 6621 4056
rect 6639 4044 6643 4056
rect 6641 4032 6643 4044
rect 6649 4044 6653 4056
rect 6649 4032 6651 4044
rect 6569 3910 6593 3912
rect 6569 3908 6605 3910
rect 6569 3904 6573 3908
rect 6615 3904 6619 3930
rect 6633 3922 6637 4032
rect 6671 4024 6675 4056
rect 6642 4020 6675 4024
rect 6642 3956 6646 4020
rect 6662 3971 6666 4000
rect 6681 3998 6685 4056
rect 6701 3999 6705 4036
rect 6662 3963 6671 3971
rect 6642 3944 6645 3956
rect 6635 3904 6639 3910
rect 6647 3904 6651 3944
rect 6667 3904 6671 3963
rect 6681 3904 6685 3986
rect 6701 3944 6705 3987
rect 43 3860 47 3864
rect 65 3860 69 3864
rect 111 3860 115 3864
rect 133 3860 137 3864
rect 141 3860 145 3864
rect 161 3860 165 3864
rect 169 3860 173 3864
rect 215 3860 219 3864
rect 235 3860 239 3864
rect 247 3860 251 3864
rect 267 3860 271 3864
rect 281 3860 285 3864
rect 301 3860 305 3864
rect 351 3860 355 3864
rect 371 3860 375 3864
rect 445 3860 449 3864
rect 465 3860 469 3864
rect 485 3860 489 3864
rect 545 3860 549 3864
rect 565 3860 569 3864
rect 625 3860 629 3864
rect 645 3860 649 3864
rect 703 3860 707 3864
rect 725 3860 729 3864
rect 771 3860 775 3864
rect 793 3860 797 3864
rect 801 3860 805 3864
rect 821 3860 825 3864
rect 829 3860 833 3864
rect 875 3860 879 3864
rect 895 3860 899 3864
rect 907 3860 911 3864
rect 927 3860 931 3864
rect 941 3860 945 3864
rect 961 3860 965 3864
rect 1025 3860 1029 3864
rect 1045 3860 1049 3864
rect 1091 3860 1095 3864
rect 1111 3860 1115 3864
rect 1171 3860 1175 3864
rect 1191 3860 1195 3864
rect 1265 3860 1269 3864
rect 1285 3860 1289 3864
rect 1305 3860 1309 3864
rect 1351 3860 1355 3864
rect 1373 3860 1377 3864
rect 1381 3860 1385 3864
rect 1401 3860 1405 3864
rect 1409 3860 1413 3864
rect 1455 3860 1459 3864
rect 1475 3860 1479 3864
rect 1487 3860 1491 3864
rect 1507 3860 1511 3864
rect 1521 3860 1525 3864
rect 1541 3860 1545 3864
rect 1605 3860 1609 3864
rect 1625 3860 1629 3864
rect 1671 3860 1675 3864
rect 1693 3860 1697 3864
rect 1751 3860 1755 3864
rect 1771 3860 1775 3864
rect 1831 3860 1835 3864
rect 1853 3860 1857 3864
rect 1861 3860 1865 3864
rect 1881 3860 1885 3864
rect 1889 3860 1893 3864
rect 1935 3860 1939 3864
rect 1955 3860 1959 3864
rect 1967 3860 1971 3864
rect 1987 3860 1991 3864
rect 2001 3860 2005 3864
rect 2021 3860 2025 3864
rect 2071 3860 2075 3864
rect 2091 3860 2095 3864
rect 2170 3860 2174 3864
rect 2192 3860 2196 3864
rect 2200 3860 2204 3864
rect 2265 3860 2269 3864
rect 2285 3860 2289 3864
rect 2331 3860 2335 3864
rect 2351 3860 2355 3864
rect 2425 3860 2429 3864
rect 2490 3860 2494 3864
rect 2512 3860 2516 3864
rect 2520 3860 2524 3864
rect 2571 3860 2575 3864
rect 2579 3860 2583 3864
rect 2677 3860 2681 3864
rect 2685 3860 2689 3864
rect 2731 3860 2735 3864
rect 2805 3860 2809 3864
rect 2865 3860 2869 3864
rect 2885 3860 2889 3864
rect 2931 3860 2935 3864
rect 2939 3860 2943 3864
rect 3016 3860 3020 3864
rect 3024 3860 3028 3864
rect 3046 3860 3050 3864
rect 3111 3860 3115 3864
rect 3171 3860 3175 3864
rect 3179 3860 3183 3864
rect 3265 3860 3269 3864
rect 3285 3860 3289 3864
rect 3345 3860 3349 3864
rect 3365 3860 3369 3864
rect 3415 3860 3419 3864
rect 3435 3860 3439 3864
rect 3449 3860 3453 3864
rect 3469 3860 3473 3864
rect 3481 3860 3485 3864
rect 3501 3860 3505 3864
rect 3547 3860 3551 3864
rect 3555 3860 3559 3864
rect 3575 3860 3579 3864
rect 3583 3860 3587 3864
rect 3605 3860 3609 3864
rect 3665 3860 3669 3864
rect 3715 3860 3719 3864
rect 3735 3860 3739 3864
rect 3749 3860 3753 3864
rect 3769 3860 3773 3864
rect 3781 3860 3785 3864
rect 3801 3860 3805 3864
rect 3847 3860 3851 3864
rect 3855 3860 3859 3864
rect 3875 3860 3879 3864
rect 3883 3860 3887 3864
rect 3905 3860 3909 3864
rect 3965 3860 3969 3864
rect 3985 3860 3989 3864
rect 4005 3860 4009 3864
rect 4051 3860 4055 3864
rect 4071 3860 4075 3864
rect 4150 3860 4154 3864
rect 4172 3860 4176 3864
rect 4180 3860 4184 3864
rect 4231 3860 4235 3864
rect 4239 3860 4243 3864
rect 4325 3860 4329 3864
rect 4385 3860 4389 3864
rect 4405 3860 4409 3864
rect 4470 3860 4474 3864
rect 4492 3860 4496 3864
rect 4500 3860 4504 3864
rect 4555 3860 4559 3864
rect 4575 3860 4579 3864
rect 4589 3860 4593 3864
rect 4609 3860 4613 3864
rect 4621 3860 4625 3864
rect 4641 3860 4645 3864
rect 4687 3860 4691 3864
rect 4695 3860 4699 3864
rect 4715 3860 4719 3864
rect 4723 3860 4727 3864
rect 4745 3860 4749 3864
rect 4805 3860 4809 3864
rect 4825 3860 4829 3864
rect 4890 3860 4894 3864
rect 4912 3860 4916 3864
rect 4920 3860 4924 3864
rect 4975 3860 4979 3864
rect 4995 3860 4999 3864
rect 5009 3860 5013 3864
rect 5029 3860 5033 3864
rect 5041 3860 5045 3864
rect 5061 3860 5065 3864
rect 5107 3860 5111 3864
rect 5115 3860 5119 3864
rect 5135 3860 5139 3864
rect 5143 3860 5147 3864
rect 5165 3860 5169 3864
rect 5225 3860 5229 3864
rect 5245 3860 5249 3864
rect 5310 3860 5314 3864
rect 5332 3860 5336 3864
rect 5340 3860 5344 3864
rect 5405 3860 5409 3864
rect 5425 3860 5429 3864
rect 5476 3860 5480 3864
rect 5484 3860 5488 3864
rect 5506 3860 5510 3864
rect 5585 3860 5589 3864
rect 5635 3860 5639 3864
rect 5655 3860 5659 3864
rect 5669 3860 5673 3864
rect 5689 3860 5693 3864
rect 5701 3860 5705 3864
rect 5721 3860 5725 3864
rect 5767 3860 5771 3864
rect 5775 3860 5779 3864
rect 5795 3860 5799 3864
rect 5803 3860 5807 3864
rect 5825 3860 5829 3864
rect 5871 3860 5875 3864
rect 5945 3860 5949 3864
rect 5965 3860 5969 3864
rect 5985 3860 5989 3864
rect 6031 3860 6035 3864
rect 6053 3860 6057 3864
rect 6061 3860 6065 3864
rect 6081 3860 6085 3864
rect 6089 3860 6093 3864
rect 6135 3860 6139 3864
rect 6155 3860 6159 3864
rect 6167 3860 6171 3864
rect 6187 3860 6191 3864
rect 6201 3860 6205 3864
rect 6221 3860 6225 3864
rect 6271 3860 6275 3864
rect 6293 3860 6297 3864
rect 6301 3860 6305 3864
rect 6321 3860 6325 3864
rect 6329 3860 6333 3864
rect 6375 3860 6379 3864
rect 6395 3860 6399 3864
rect 6407 3860 6411 3864
rect 6427 3860 6431 3864
rect 6441 3860 6445 3864
rect 6461 3860 6465 3864
rect 6511 3860 6515 3864
rect 6533 3860 6537 3864
rect 6541 3860 6545 3864
rect 6561 3860 6565 3864
rect 6569 3860 6573 3864
rect 6615 3860 6619 3864
rect 6635 3860 6639 3864
rect 6647 3860 6651 3864
rect 6667 3860 6671 3864
rect 6681 3860 6685 3864
rect 6701 3860 6705 3864
rect 43 3836 47 3840
rect 65 3836 69 3840
rect 123 3836 127 3840
rect 145 3836 149 3840
rect 205 3836 209 3840
rect 225 3836 229 3840
rect 271 3836 275 3840
rect 293 3836 297 3840
rect 301 3836 305 3840
rect 321 3836 325 3840
rect 329 3836 333 3840
rect 375 3836 379 3840
rect 395 3836 399 3840
rect 407 3836 411 3840
rect 427 3836 431 3840
rect 441 3836 445 3840
rect 461 3836 465 3840
rect 525 3836 529 3840
rect 545 3836 549 3840
rect 565 3836 569 3840
rect 625 3836 629 3840
rect 645 3836 649 3840
rect 691 3836 695 3840
rect 711 3836 715 3840
rect 785 3836 789 3840
rect 805 3836 809 3840
rect 851 3836 855 3840
rect 873 3836 877 3840
rect 881 3836 885 3840
rect 901 3836 905 3840
rect 909 3836 913 3840
rect 955 3836 959 3840
rect 975 3836 979 3840
rect 987 3836 991 3840
rect 1007 3836 1011 3840
rect 1021 3836 1025 3840
rect 1041 3836 1045 3840
rect 1091 3836 1095 3840
rect 1111 3836 1115 3840
rect 1131 3836 1135 3840
rect 1205 3836 1209 3840
rect 1225 3836 1229 3840
rect 1271 3836 1275 3840
rect 1293 3836 1297 3840
rect 1365 3836 1369 3840
rect 1385 3836 1389 3840
rect 1405 3836 1409 3840
rect 1465 3836 1469 3840
rect 1485 3836 1489 3840
rect 1531 3836 1535 3840
rect 1551 3836 1555 3840
rect 1611 3836 1615 3840
rect 1619 3836 1623 3840
rect 1691 3836 1695 3840
rect 1713 3836 1717 3840
rect 1721 3836 1725 3840
rect 1741 3836 1745 3840
rect 1749 3836 1753 3840
rect 1795 3836 1799 3840
rect 1815 3836 1819 3840
rect 1827 3836 1831 3840
rect 1847 3836 1851 3840
rect 1861 3836 1865 3840
rect 1881 3836 1885 3840
rect 1945 3836 1949 3840
rect 1965 3836 1969 3840
rect 2011 3836 2015 3840
rect 2019 3836 2023 3840
rect 2091 3836 2095 3840
rect 2156 3836 2160 3840
rect 2164 3836 2168 3840
rect 2186 3836 2190 3840
rect 2270 3836 2274 3840
rect 2292 3836 2296 3840
rect 2300 3836 2304 3840
rect 2365 3836 2369 3840
rect 2385 3836 2389 3840
rect 2405 3836 2409 3840
rect 2451 3836 2455 3840
rect 2525 3836 2529 3840
rect 2576 3836 2580 3840
rect 2584 3836 2588 3840
rect 2606 3836 2610 3840
rect 2671 3836 2675 3840
rect 2691 3836 2695 3840
rect 2711 3836 2715 3840
rect 2785 3836 2789 3840
rect 2845 3836 2849 3840
rect 2865 3836 2869 3840
rect 2916 3836 2920 3840
rect 2924 3836 2928 3840
rect 2946 3836 2950 3840
rect 3016 3836 3020 3840
rect 3024 3836 3028 3840
rect 3046 3836 3050 3840
rect 3111 3836 3115 3840
rect 3131 3836 3135 3840
rect 3151 3836 3155 3840
rect 3225 3836 3229 3840
rect 3245 3836 3249 3840
rect 3265 3836 3269 3840
rect 3285 3836 3289 3840
rect 3345 3836 3349 3840
rect 3365 3836 3369 3840
rect 3425 3836 3429 3840
rect 3445 3836 3449 3840
rect 3495 3836 3499 3840
rect 3515 3836 3519 3840
rect 3529 3836 3533 3840
rect 3549 3836 3553 3840
rect 3561 3836 3565 3840
rect 3581 3836 3585 3840
rect 3627 3836 3631 3840
rect 3635 3836 3639 3840
rect 3655 3836 3659 3840
rect 3663 3836 3667 3840
rect 3685 3836 3689 3840
rect 3745 3836 3749 3840
rect 3765 3836 3769 3840
rect 3825 3836 3829 3840
rect 3845 3836 3849 3840
rect 3865 3836 3869 3840
rect 3885 3836 3889 3840
rect 3931 3836 3935 3840
rect 3991 3836 3995 3840
rect 4011 3836 4015 3840
rect 4076 3836 4080 3840
rect 4084 3836 4088 3840
rect 4106 3836 4110 3840
rect 4175 3836 4179 3840
rect 4195 3836 4199 3840
rect 4209 3836 4213 3840
rect 4229 3836 4233 3840
rect 4241 3836 4245 3840
rect 4261 3836 4265 3840
rect 4307 3836 4311 3840
rect 4315 3836 4319 3840
rect 4335 3836 4339 3840
rect 4343 3836 4347 3840
rect 4365 3836 4369 3840
rect 4411 3836 4415 3840
rect 4431 3836 4435 3840
rect 4505 3836 4509 3840
rect 4525 3836 4529 3840
rect 4585 3836 4589 3840
rect 4605 3836 4609 3840
rect 4625 3836 4629 3840
rect 4645 3836 4649 3840
rect 4665 3836 4669 3840
rect 4685 3836 4689 3840
rect 4705 3836 4709 3840
rect 4725 3836 4729 3840
rect 4775 3836 4779 3840
rect 4795 3836 4799 3840
rect 4809 3836 4813 3840
rect 4829 3836 4833 3840
rect 4841 3836 4845 3840
rect 4861 3836 4865 3840
rect 4907 3836 4911 3840
rect 4915 3836 4919 3840
rect 4935 3836 4939 3840
rect 4943 3836 4947 3840
rect 4965 3836 4969 3840
rect 5016 3836 5020 3840
rect 5024 3836 5028 3840
rect 5046 3836 5050 3840
rect 5125 3836 5129 3840
rect 5145 3836 5149 3840
rect 5205 3836 5209 3840
rect 5225 3836 5229 3840
rect 5285 3836 5289 3840
rect 5331 3836 5335 3840
rect 5351 3836 5355 3840
rect 5371 3836 5375 3840
rect 5391 3836 5395 3840
rect 5411 3836 5415 3840
rect 5431 3836 5435 3840
rect 5451 3836 5455 3840
rect 5471 3836 5475 3840
rect 5531 3836 5535 3840
rect 5553 3836 5557 3840
rect 5561 3836 5565 3840
rect 5581 3836 5585 3840
rect 5589 3836 5593 3840
rect 5635 3836 5639 3840
rect 5655 3836 5659 3840
rect 5667 3836 5671 3840
rect 5687 3836 5691 3840
rect 5701 3836 5705 3840
rect 5721 3836 5725 3840
rect 5785 3836 5789 3840
rect 5831 3836 5835 3840
rect 5851 3836 5855 3840
rect 5911 3836 5915 3840
rect 5931 3836 5935 3840
rect 6005 3836 6009 3840
rect 6051 3836 6055 3840
rect 6059 3836 6063 3840
rect 6157 3836 6161 3840
rect 6165 3836 6169 3840
rect 6211 3836 6215 3840
rect 6231 3836 6235 3840
rect 6251 3836 6255 3840
rect 6311 3836 6315 3840
rect 6333 3836 6337 3840
rect 6341 3836 6345 3840
rect 6361 3836 6365 3840
rect 6369 3836 6373 3840
rect 6415 3836 6419 3840
rect 6435 3836 6439 3840
rect 6447 3836 6451 3840
rect 6467 3836 6471 3840
rect 6481 3836 6485 3840
rect 6501 3836 6505 3840
rect 6556 3836 6560 3840
rect 6564 3836 6568 3840
rect 6586 3836 6590 3840
rect 6651 3836 6655 3840
rect 6671 3836 6675 3840
rect 43 3750 47 3756
rect 43 3738 45 3750
rect 65 3733 69 3796
rect 123 3750 127 3756
rect 123 3738 125 3750
rect 145 3733 149 3796
rect 65 3721 74 3733
rect 145 3721 154 3733
rect 43 3670 45 3682
rect 43 3664 47 3670
rect 65 3644 69 3721
rect 123 3670 125 3682
rect 123 3664 127 3670
rect 145 3644 149 3721
rect 205 3719 209 3796
rect 206 3707 209 3719
rect 203 3691 209 3707
rect 225 3719 229 3796
rect 293 3793 297 3816
rect 289 3786 297 3793
rect 289 3757 293 3786
rect 301 3776 305 3816
rect 321 3764 325 3796
rect 329 3792 333 3796
rect 329 3790 365 3792
rect 329 3788 353 3790
rect 271 3744 275 3756
rect 289 3751 297 3757
rect 271 3732 273 3744
rect 225 3707 234 3719
rect 225 3691 231 3707
rect 203 3684 217 3691
rect 213 3664 217 3684
rect 223 3684 231 3691
rect 223 3664 227 3684
rect 271 3664 275 3732
rect 293 3705 297 3751
rect 293 3644 297 3693
rect 321 3669 327 3764
rect 303 3665 327 3669
rect 303 3644 307 3665
rect 323 3660 341 3661
rect 323 3656 353 3660
rect 323 3644 327 3656
rect 361 3652 365 3778
rect 375 3770 379 3796
rect 395 3790 399 3796
rect 331 3648 365 3652
rect 331 3644 335 3648
rect 377 3644 381 3758
rect 393 3668 397 3778
rect 407 3756 411 3796
rect 402 3744 405 3756
rect 402 3680 406 3744
rect 427 3737 431 3796
rect 422 3729 431 3737
rect 422 3700 426 3729
rect 441 3714 445 3796
rect 461 3713 465 3756
rect 402 3676 435 3680
rect 401 3656 403 3668
rect 399 3644 403 3656
rect 409 3656 411 3668
rect 409 3644 413 3656
rect 431 3644 435 3676
rect 441 3644 445 3702
rect 461 3664 465 3701
rect 525 3699 529 3756
rect 545 3742 549 3756
rect 565 3742 569 3756
rect 545 3736 560 3742
rect 565 3736 581 3742
rect 554 3713 560 3736
rect 525 3687 534 3699
rect 532 3644 536 3687
rect 554 3664 558 3701
rect 574 3699 581 3736
rect 625 3719 629 3796
rect 626 3707 629 3719
rect 623 3691 629 3707
rect 645 3719 649 3796
rect 691 3719 695 3796
rect 645 3707 654 3719
rect 686 3707 695 3719
rect 645 3691 651 3707
rect 574 3674 581 3687
rect 623 3684 637 3691
rect 562 3668 581 3674
rect 562 3664 566 3668
rect 633 3664 637 3684
rect 643 3684 651 3691
rect 689 3691 695 3707
rect 711 3719 715 3796
rect 785 3719 789 3796
rect 711 3707 714 3719
rect 786 3707 789 3719
rect 711 3691 717 3707
rect 689 3684 697 3691
rect 643 3664 647 3684
rect 693 3664 697 3684
rect 703 3684 717 3691
rect 783 3691 789 3707
rect 805 3719 809 3796
rect 873 3793 877 3816
rect 869 3786 877 3793
rect 869 3757 873 3786
rect 881 3776 885 3816
rect 901 3764 905 3796
rect 909 3792 913 3796
rect 909 3790 945 3792
rect 909 3788 933 3790
rect 851 3744 855 3756
rect 869 3751 877 3757
rect 851 3732 853 3744
rect 805 3707 814 3719
rect 805 3691 811 3707
rect 783 3684 797 3691
rect 703 3664 707 3684
rect 793 3664 797 3684
rect 803 3684 811 3691
rect 803 3664 807 3684
rect 851 3664 855 3732
rect 873 3705 877 3751
rect 873 3644 877 3693
rect 901 3669 907 3764
rect 883 3665 907 3669
rect 883 3644 887 3665
rect 903 3660 921 3661
rect 903 3656 933 3660
rect 903 3644 907 3656
rect 941 3652 945 3778
rect 955 3770 959 3796
rect 975 3790 979 3796
rect 911 3648 945 3652
rect 911 3644 915 3648
rect 957 3644 961 3758
rect 973 3668 977 3778
rect 987 3756 991 3796
rect 982 3744 985 3756
rect 982 3680 986 3744
rect 1007 3737 1011 3796
rect 1002 3729 1011 3737
rect 1002 3700 1006 3729
rect 1021 3714 1025 3796
rect 1041 3713 1045 3756
rect 1091 3742 1095 3756
rect 1111 3742 1115 3756
rect 1079 3736 1095 3742
rect 1100 3736 1115 3742
rect 982 3676 1015 3680
rect 981 3656 983 3668
rect 979 3644 983 3656
rect 989 3656 991 3668
rect 989 3644 993 3656
rect 1011 3644 1015 3676
rect 1021 3644 1025 3702
rect 1041 3664 1045 3701
rect 1079 3699 1086 3736
rect 1100 3713 1106 3736
rect 1079 3674 1086 3687
rect 1079 3668 1098 3674
rect 1094 3664 1098 3668
rect 1102 3664 1106 3701
rect 1131 3699 1135 3756
rect 1205 3719 1209 3796
rect 1206 3707 1209 3719
rect 1126 3687 1135 3699
rect 1203 3691 1209 3707
rect 1225 3719 1229 3796
rect 1271 3733 1275 3796
rect 1293 3750 1297 3756
rect 1295 3738 1297 3750
rect 1266 3721 1275 3733
rect 1225 3707 1234 3719
rect 1225 3691 1231 3707
rect 1124 3644 1128 3687
rect 1203 3684 1217 3691
rect 1213 3664 1217 3684
rect 1223 3684 1231 3691
rect 1223 3664 1227 3684
rect 1271 3644 1275 3721
rect 1365 3699 1369 3756
rect 1385 3742 1389 3756
rect 1405 3742 1409 3756
rect 1385 3736 1400 3742
rect 1405 3736 1421 3742
rect 1394 3713 1400 3736
rect 1365 3687 1374 3699
rect 1295 3670 1297 3682
rect 1293 3664 1297 3670
rect 1372 3644 1376 3687
rect 1394 3664 1398 3701
rect 1414 3699 1421 3736
rect 1465 3719 1469 3796
rect 1466 3707 1469 3719
rect 1463 3691 1469 3707
rect 1485 3719 1489 3796
rect 1531 3719 1535 3796
rect 1485 3707 1494 3719
rect 1526 3707 1535 3719
rect 1485 3691 1491 3707
rect 1414 3674 1421 3687
rect 1463 3684 1477 3691
rect 1402 3668 1421 3674
rect 1402 3664 1406 3668
rect 1473 3664 1477 3684
rect 1483 3684 1491 3691
rect 1529 3691 1535 3707
rect 1551 3719 1555 3796
rect 1713 3793 1717 3816
rect 1709 3786 1717 3793
rect 1709 3757 1713 3786
rect 1721 3776 1725 3816
rect 1741 3764 1745 3796
rect 1749 3792 1753 3796
rect 1749 3790 1785 3792
rect 1749 3788 1773 3790
rect 1611 3733 1615 3756
rect 1606 3721 1615 3733
rect 1619 3733 1623 3756
rect 1691 3744 1695 3756
rect 1709 3751 1717 3757
rect 1619 3721 1634 3733
rect 1691 3732 1693 3744
rect 1551 3707 1554 3719
rect 1551 3691 1557 3707
rect 1529 3684 1537 3691
rect 1483 3664 1487 3684
rect 1533 3664 1537 3684
rect 1543 3684 1557 3691
rect 1543 3664 1547 3684
rect 1611 3644 1615 3721
rect 1631 3644 1635 3721
rect 1691 3664 1695 3732
rect 1713 3705 1717 3751
rect 1713 3644 1717 3693
rect 1741 3669 1747 3764
rect 1723 3665 1747 3669
rect 1723 3644 1727 3665
rect 1743 3660 1761 3661
rect 1743 3656 1773 3660
rect 1743 3644 1747 3656
rect 1781 3652 1785 3778
rect 1795 3770 1799 3796
rect 1815 3790 1819 3796
rect 1751 3648 1785 3652
rect 1751 3644 1755 3648
rect 1797 3644 1801 3758
rect 1813 3668 1817 3778
rect 1827 3756 1831 3796
rect 1822 3744 1825 3756
rect 1822 3680 1826 3744
rect 1847 3737 1851 3796
rect 1842 3729 1851 3737
rect 1842 3700 1846 3729
rect 1861 3714 1865 3796
rect 1881 3713 1885 3756
rect 1945 3719 1949 3796
rect 1822 3676 1855 3680
rect 1821 3656 1823 3668
rect 1819 3644 1823 3656
rect 1829 3656 1831 3668
rect 1829 3644 1833 3656
rect 1851 3644 1855 3676
rect 1861 3644 1865 3702
rect 1946 3707 1949 3719
rect 1881 3664 1885 3701
rect 1943 3691 1949 3707
rect 1965 3719 1969 3796
rect 2011 3733 2015 3756
rect 2006 3721 2015 3733
rect 2019 3733 2023 3756
rect 2019 3721 2034 3733
rect 1965 3707 1974 3719
rect 1965 3691 1971 3707
rect 1943 3684 1957 3691
rect 1953 3664 1957 3684
rect 1963 3684 1971 3691
rect 1963 3664 1967 3684
rect 2011 3644 2015 3721
rect 2031 3644 2035 3721
rect 2091 3713 2095 3796
rect 2156 3752 2160 3756
rect 2142 3744 2160 3752
rect 2142 3733 2146 3744
rect 2086 3701 2095 3713
rect 2091 3644 2095 3701
rect 2142 3676 2146 3721
rect 2164 3699 2168 3756
rect 2186 3753 2190 3796
rect 2270 3753 2274 3796
rect 2186 3741 2193 3753
rect 2267 3741 2274 3753
rect 2166 3687 2175 3699
rect 2142 3669 2155 3676
rect 2151 3664 2155 3669
rect 2171 3664 2175 3687
rect 2191 3664 2195 3741
rect 2265 3664 2269 3741
rect 2292 3699 2296 3756
rect 2300 3752 2304 3756
rect 2300 3744 2318 3752
rect 2314 3733 2318 3744
rect 2285 3687 2294 3699
rect 2285 3664 2289 3687
rect 2314 3676 2318 3721
rect 2365 3699 2369 3756
rect 2385 3742 2389 3756
rect 2405 3742 2409 3756
rect 2385 3736 2400 3742
rect 2405 3736 2421 3742
rect 2394 3713 2400 3736
rect 2365 3687 2374 3699
rect 2305 3669 2318 3676
rect 2305 3664 2309 3669
rect 2372 3644 2376 3687
rect 2394 3664 2398 3701
rect 2414 3699 2421 3736
rect 2451 3713 2455 3796
rect 2446 3701 2455 3713
rect 2414 3674 2421 3687
rect 2402 3668 2421 3674
rect 2402 3664 2406 3668
rect 2451 3644 2455 3701
rect 2525 3713 2529 3796
rect 2576 3752 2580 3756
rect 2562 3744 2580 3752
rect 2562 3733 2566 3744
rect 2525 3701 2534 3713
rect 2525 3644 2529 3701
rect 2562 3676 2566 3721
rect 2584 3699 2588 3756
rect 2606 3753 2610 3796
rect 2671 3788 2675 3796
rect 2660 3784 2675 3788
rect 2691 3784 2695 3796
rect 2660 3753 2666 3784
rect 2680 3780 2695 3784
rect 2680 3773 2686 3780
rect 2606 3741 2613 3753
rect 2666 3741 2676 3753
rect 2586 3687 2595 3699
rect 2562 3669 2575 3676
rect 2571 3664 2575 3669
rect 2591 3664 2595 3687
rect 2611 3664 2615 3741
rect 2672 3684 2676 3741
rect 2680 3684 2684 3761
rect 2711 3753 2715 3796
rect 2688 3741 2695 3753
rect 2707 3741 2715 3753
rect 2688 3684 2692 3741
rect 2785 3713 2789 3796
rect 2845 3719 2849 3796
rect 2785 3701 2794 3713
rect 2846 3707 2849 3719
rect 2785 3644 2789 3701
rect 2843 3691 2849 3707
rect 2865 3719 2869 3796
rect 2916 3752 2920 3756
rect 2902 3744 2920 3752
rect 2902 3733 2906 3744
rect 2865 3707 2874 3719
rect 2865 3691 2871 3707
rect 2843 3684 2857 3691
rect 2853 3664 2857 3684
rect 2863 3684 2871 3691
rect 2863 3664 2867 3684
rect 2902 3676 2906 3721
rect 2924 3699 2928 3756
rect 2946 3753 2950 3796
rect 2946 3741 2953 3753
rect 3016 3752 3020 3756
rect 3002 3744 3020 3752
rect 2926 3687 2935 3699
rect 2902 3669 2915 3676
rect 2911 3664 2915 3669
rect 2931 3664 2935 3687
rect 2951 3664 2955 3741
rect 3002 3733 3006 3744
rect 3002 3676 3006 3721
rect 3024 3699 3028 3756
rect 3046 3753 3050 3796
rect 3046 3741 3053 3753
rect 3111 3742 3115 3756
rect 3131 3742 3135 3756
rect 3026 3687 3035 3699
rect 3002 3669 3015 3676
rect 3011 3664 3015 3669
rect 3031 3664 3035 3687
rect 3051 3664 3055 3741
rect 3099 3736 3115 3742
rect 3120 3736 3135 3742
rect 3099 3699 3106 3736
rect 3120 3713 3126 3736
rect 3099 3674 3106 3687
rect 3099 3668 3118 3674
rect 3114 3664 3118 3668
rect 3122 3664 3126 3701
rect 3151 3699 3155 3756
rect 3225 3733 3229 3756
rect 3226 3721 3229 3733
rect 3146 3687 3155 3699
rect 3144 3644 3148 3687
rect 3220 3673 3226 3721
rect 3245 3699 3249 3756
rect 3265 3734 3269 3756
rect 3285 3734 3289 3756
rect 3265 3728 3278 3734
rect 3285 3733 3305 3734
rect 3285 3728 3293 3733
rect 3274 3699 3278 3728
rect 3247 3687 3249 3699
rect 3245 3685 3249 3687
rect 3245 3678 3258 3685
rect 3220 3669 3250 3673
rect 3246 3664 3250 3669
rect 3254 3664 3258 3678
rect 3274 3664 3278 3687
rect 3293 3679 3299 3721
rect 3345 3719 3349 3796
rect 3346 3707 3349 3719
rect 3343 3691 3349 3707
rect 3365 3719 3369 3796
rect 3425 3719 3429 3796
rect 3365 3707 3374 3719
rect 3426 3707 3429 3719
rect 3365 3691 3371 3707
rect 3343 3684 3357 3691
rect 3282 3672 3299 3679
rect 3282 3664 3286 3672
rect 3353 3664 3357 3684
rect 3363 3684 3371 3691
rect 3423 3691 3429 3707
rect 3445 3719 3449 3796
rect 3445 3707 3454 3719
rect 3495 3713 3499 3756
rect 3515 3714 3519 3796
rect 3529 3737 3533 3796
rect 3549 3756 3553 3796
rect 3561 3790 3565 3796
rect 3555 3744 3558 3756
rect 3529 3729 3538 3737
rect 3445 3691 3451 3707
rect 3423 3684 3437 3691
rect 3363 3664 3367 3684
rect 3433 3664 3437 3684
rect 3443 3684 3451 3691
rect 3443 3664 3447 3684
rect 3495 3664 3499 3701
rect 3515 3644 3519 3702
rect 3534 3700 3538 3729
rect 3554 3680 3558 3744
rect 3525 3676 3558 3680
rect 3525 3644 3529 3676
rect 3563 3668 3567 3778
rect 3581 3770 3585 3796
rect 3627 3792 3631 3796
rect 3595 3790 3631 3792
rect 3607 3788 3631 3790
rect 3549 3656 3551 3668
rect 3547 3644 3551 3656
rect 3557 3656 3559 3668
rect 3557 3644 3561 3656
rect 3579 3644 3583 3758
rect 3595 3652 3599 3778
rect 3635 3764 3639 3796
rect 3655 3776 3659 3816
rect 3663 3793 3667 3816
rect 3663 3786 3671 3793
rect 3633 3669 3639 3764
rect 3667 3757 3671 3786
rect 3663 3751 3671 3757
rect 3663 3705 3667 3751
rect 3685 3744 3689 3756
rect 3687 3732 3689 3744
rect 3633 3665 3657 3669
rect 3619 3660 3637 3661
rect 3607 3656 3637 3660
rect 3595 3648 3629 3652
rect 3625 3644 3629 3648
rect 3633 3644 3637 3656
rect 3653 3644 3657 3665
rect 3663 3644 3667 3693
rect 3685 3664 3689 3732
rect 3745 3719 3749 3796
rect 3746 3707 3749 3719
rect 3743 3691 3749 3707
rect 3765 3719 3769 3796
rect 3825 3733 3829 3756
rect 3826 3721 3829 3733
rect 3765 3707 3774 3719
rect 3765 3691 3771 3707
rect 3743 3684 3757 3691
rect 3753 3664 3757 3684
rect 3763 3684 3771 3691
rect 3763 3664 3767 3684
rect 3820 3673 3826 3721
rect 3845 3699 3849 3756
rect 3865 3734 3869 3756
rect 3885 3734 3889 3756
rect 3865 3728 3878 3734
rect 3885 3733 3905 3734
rect 3885 3728 3893 3733
rect 3874 3699 3878 3728
rect 3847 3687 3849 3699
rect 3845 3685 3849 3687
rect 3845 3678 3858 3685
rect 3820 3669 3850 3673
rect 3846 3664 3850 3669
rect 3854 3664 3858 3678
rect 3874 3664 3878 3687
rect 3893 3679 3899 3721
rect 3931 3713 3935 3796
rect 3991 3719 3995 3796
rect 3926 3701 3935 3713
rect 3986 3707 3995 3719
rect 3882 3672 3899 3679
rect 3882 3664 3886 3672
rect 3931 3644 3935 3701
rect 3989 3691 3995 3707
rect 4011 3719 4015 3796
rect 4076 3752 4080 3756
rect 4062 3744 4080 3752
rect 4062 3733 4066 3744
rect 4011 3707 4014 3719
rect 4011 3691 4017 3707
rect 3989 3684 3997 3691
rect 3993 3664 3997 3684
rect 4003 3684 4017 3691
rect 4003 3664 4007 3684
rect 4062 3676 4066 3721
rect 4084 3699 4088 3756
rect 4106 3753 4110 3796
rect 4106 3741 4113 3753
rect 4086 3687 4095 3699
rect 4062 3669 4075 3676
rect 4071 3664 4075 3669
rect 4091 3664 4095 3687
rect 4111 3664 4115 3741
rect 4175 3713 4179 3756
rect 4195 3714 4199 3796
rect 4209 3737 4213 3796
rect 4229 3756 4233 3796
rect 4241 3790 4245 3796
rect 4235 3744 4238 3756
rect 4209 3729 4218 3737
rect 4175 3664 4179 3701
rect 4195 3644 4199 3702
rect 4214 3700 4218 3729
rect 4234 3680 4238 3744
rect 4205 3676 4238 3680
rect 4205 3644 4209 3676
rect 4243 3668 4247 3778
rect 4261 3770 4265 3796
rect 4307 3792 4311 3796
rect 4275 3790 4311 3792
rect 4287 3788 4311 3790
rect 4229 3656 4231 3668
rect 4227 3644 4231 3656
rect 4237 3656 4239 3668
rect 4237 3644 4241 3656
rect 4259 3644 4263 3758
rect 4275 3652 4279 3778
rect 4315 3764 4319 3796
rect 4335 3776 4339 3816
rect 4343 3793 4347 3816
rect 4343 3786 4351 3793
rect 4313 3669 4319 3764
rect 4347 3757 4351 3786
rect 4343 3751 4351 3757
rect 4343 3705 4347 3751
rect 4365 3744 4369 3756
rect 4367 3732 4369 3744
rect 4313 3665 4337 3669
rect 4299 3660 4317 3661
rect 4287 3656 4317 3660
rect 4275 3648 4309 3652
rect 4305 3644 4309 3648
rect 4313 3644 4317 3656
rect 4333 3644 4337 3665
rect 4343 3644 4347 3693
rect 4365 3664 4369 3732
rect 4411 3719 4415 3796
rect 4406 3707 4415 3719
rect 4409 3691 4415 3707
rect 4431 3719 4435 3796
rect 4505 3719 4509 3796
rect 4431 3707 4434 3719
rect 4506 3707 4509 3719
rect 4431 3691 4437 3707
rect 4409 3684 4417 3691
rect 4413 3664 4417 3684
rect 4423 3684 4437 3691
rect 4503 3691 4509 3707
rect 4525 3719 4529 3796
rect 4525 3707 4534 3719
rect 4525 3691 4531 3707
rect 4503 3684 4517 3691
rect 4423 3664 4427 3684
rect 4513 3664 4517 3684
rect 4523 3684 4531 3691
rect 4585 3696 4589 3756
rect 4605 3696 4609 3756
rect 4625 3696 4629 3756
rect 4645 3696 4649 3756
rect 4665 3696 4669 3756
rect 4685 3696 4689 3756
rect 4705 3699 4709 3756
rect 4725 3699 4729 3756
rect 4775 3713 4779 3756
rect 4795 3714 4799 3796
rect 4809 3737 4813 3796
rect 4829 3756 4833 3796
rect 4841 3790 4845 3796
rect 4835 3744 4838 3756
rect 4809 3729 4818 3737
rect 4585 3684 4598 3696
rect 4625 3684 4638 3696
rect 4665 3684 4678 3696
rect 4705 3687 4714 3699
rect 4726 3687 4729 3699
rect 4523 3664 4527 3684
rect 4585 3664 4589 3684
rect 4605 3664 4609 3684
rect 4625 3664 4629 3684
rect 4645 3664 4649 3684
rect 4665 3664 4669 3684
rect 4685 3664 4689 3684
rect 4705 3664 4709 3687
rect 4725 3664 4729 3687
rect 4775 3664 4779 3701
rect 4795 3644 4799 3702
rect 4814 3700 4818 3729
rect 4834 3680 4838 3744
rect 4805 3676 4838 3680
rect 4805 3644 4809 3676
rect 4843 3668 4847 3778
rect 4861 3770 4865 3796
rect 4907 3792 4911 3796
rect 4875 3790 4911 3792
rect 4887 3788 4911 3790
rect 4829 3656 4831 3668
rect 4827 3644 4831 3656
rect 4837 3656 4839 3668
rect 4837 3644 4841 3656
rect 4859 3644 4863 3758
rect 4875 3652 4879 3778
rect 4915 3764 4919 3796
rect 4935 3776 4939 3816
rect 4943 3793 4947 3816
rect 4943 3786 4951 3793
rect 4913 3669 4919 3764
rect 4947 3757 4951 3786
rect 4943 3751 4951 3757
rect 4943 3705 4947 3751
rect 4965 3744 4969 3756
rect 5016 3752 5020 3756
rect 4967 3732 4969 3744
rect 5002 3744 5020 3752
rect 5002 3733 5006 3744
rect 4913 3665 4937 3669
rect 4899 3660 4917 3661
rect 4887 3656 4917 3660
rect 4875 3648 4909 3652
rect 4905 3644 4909 3648
rect 4913 3644 4917 3656
rect 4933 3644 4937 3665
rect 4943 3644 4947 3693
rect 4965 3664 4969 3732
rect 5002 3676 5006 3721
rect 5024 3699 5028 3756
rect 5046 3753 5050 3796
rect 5046 3741 5053 3753
rect 5026 3687 5035 3699
rect 5002 3669 5015 3676
rect 5011 3664 5015 3669
rect 5031 3664 5035 3687
rect 5051 3664 5055 3741
rect 5125 3719 5129 3796
rect 5126 3707 5129 3719
rect 5123 3691 5129 3707
rect 5145 3719 5149 3796
rect 5205 3719 5209 3796
rect 5145 3707 5154 3719
rect 5206 3707 5209 3719
rect 5145 3691 5151 3707
rect 5123 3684 5137 3691
rect 5133 3664 5137 3684
rect 5143 3684 5151 3691
rect 5203 3691 5209 3707
rect 5225 3719 5229 3796
rect 5225 3707 5234 3719
rect 5285 3713 5289 3796
rect 5553 3793 5557 3816
rect 5549 3786 5557 3793
rect 5549 3757 5553 3786
rect 5561 3776 5565 3816
rect 5581 3764 5585 3796
rect 5589 3792 5593 3796
rect 5589 3790 5625 3792
rect 5589 3788 5613 3790
rect 5225 3691 5231 3707
rect 5203 3684 5217 3691
rect 5143 3664 5147 3684
rect 5213 3664 5217 3684
rect 5223 3684 5231 3691
rect 5285 3701 5294 3713
rect 5223 3664 5227 3684
rect 5285 3644 5289 3701
rect 5331 3699 5335 3756
rect 5351 3699 5355 3756
rect 5331 3687 5334 3699
rect 5346 3687 5355 3699
rect 5371 3696 5375 3756
rect 5391 3696 5395 3756
rect 5411 3696 5415 3756
rect 5431 3696 5435 3756
rect 5451 3696 5455 3756
rect 5471 3696 5475 3756
rect 5331 3664 5335 3687
rect 5351 3664 5355 3687
rect 5382 3684 5395 3696
rect 5422 3684 5435 3696
rect 5462 3684 5475 3696
rect 5371 3664 5375 3684
rect 5391 3664 5395 3684
rect 5411 3664 5415 3684
rect 5431 3664 5435 3684
rect 5451 3664 5455 3684
rect 5471 3664 5475 3684
rect 5531 3744 5535 3756
rect 5549 3751 5557 3757
rect 5531 3732 5533 3744
rect 5531 3664 5535 3732
rect 5553 3705 5557 3751
rect 5553 3644 5557 3693
rect 5581 3669 5587 3764
rect 5563 3665 5587 3669
rect 5563 3644 5567 3665
rect 5583 3660 5601 3661
rect 5583 3656 5613 3660
rect 5583 3644 5587 3656
rect 5621 3652 5625 3778
rect 5635 3770 5639 3796
rect 5655 3790 5659 3796
rect 5591 3648 5625 3652
rect 5591 3644 5595 3648
rect 5637 3644 5641 3758
rect 5653 3668 5657 3778
rect 5667 3756 5671 3796
rect 5662 3744 5665 3756
rect 5662 3680 5666 3744
rect 5687 3737 5691 3796
rect 5682 3729 5691 3737
rect 5682 3700 5686 3729
rect 5701 3714 5705 3796
rect 5721 3713 5725 3756
rect 5785 3713 5789 3796
rect 5831 3719 5835 3796
rect 5662 3676 5695 3680
rect 5661 3656 5663 3668
rect 5659 3644 5663 3656
rect 5669 3656 5671 3668
rect 5669 3644 5673 3656
rect 5691 3644 5695 3676
rect 5701 3644 5705 3702
rect 5785 3701 5794 3713
rect 5826 3707 5835 3719
rect 5721 3664 5725 3701
rect 5785 3644 5789 3701
rect 5829 3691 5835 3707
rect 5851 3719 5855 3796
rect 5911 3719 5915 3796
rect 5851 3707 5854 3719
rect 5906 3707 5915 3719
rect 5851 3691 5857 3707
rect 5829 3684 5837 3691
rect 5833 3664 5837 3684
rect 5843 3684 5857 3691
rect 5909 3691 5915 3707
rect 5931 3719 5935 3796
rect 5931 3707 5934 3719
rect 6005 3713 6009 3796
rect 6333 3793 6337 3816
rect 6329 3786 6337 3793
rect 6329 3757 6333 3786
rect 6341 3776 6345 3816
rect 6361 3764 6365 3796
rect 6369 3792 6373 3796
rect 6369 3790 6405 3792
rect 6369 3788 6393 3790
rect 6051 3733 6055 3756
rect 6046 3721 6055 3733
rect 6059 3733 6063 3756
rect 6157 3733 6161 3756
rect 6059 3721 6074 3733
rect 6146 3721 6161 3733
rect 6165 3733 6169 3756
rect 6211 3742 6215 3756
rect 6231 3742 6235 3756
rect 6199 3736 6215 3742
rect 6220 3736 6235 3742
rect 6165 3721 6174 3733
rect 5931 3691 5937 3707
rect 5909 3684 5917 3691
rect 5843 3664 5847 3684
rect 5913 3664 5917 3684
rect 5923 3684 5937 3691
rect 6005 3701 6014 3713
rect 5923 3664 5927 3684
rect 6005 3644 6009 3701
rect 6051 3644 6055 3721
rect 6071 3644 6075 3721
rect 6145 3644 6149 3721
rect 6165 3644 6169 3721
rect 6199 3699 6206 3736
rect 6220 3713 6226 3736
rect 6199 3674 6206 3687
rect 6199 3668 6218 3674
rect 6214 3664 6218 3668
rect 6222 3664 6226 3701
rect 6251 3699 6255 3756
rect 6246 3687 6255 3699
rect 6311 3744 6315 3756
rect 6329 3751 6337 3757
rect 6311 3732 6313 3744
rect 6244 3644 6248 3687
rect 6311 3664 6315 3732
rect 6333 3705 6337 3751
rect 6333 3644 6337 3693
rect 6361 3669 6367 3764
rect 6343 3665 6367 3669
rect 6343 3644 6347 3665
rect 6363 3660 6381 3661
rect 6363 3656 6393 3660
rect 6363 3644 6367 3656
rect 6401 3652 6405 3778
rect 6415 3770 6419 3796
rect 6435 3790 6439 3796
rect 6371 3648 6405 3652
rect 6371 3644 6375 3648
rect 6417 3644 6421 3758
rect 6433 3668 6437 3778
rect 6447 3756 6451 3796
rect 6442 3744 6445 3756
rect 6442 3680 6446 3744
rect 6467 3737 6471 3796
rect 6462 3729 6471 3737
rect 6462 3700 6466 3729
rect 6481 3714 6485 3796
rect 6501 3713 6505 3756
rect 6556 3752 6560 3756
rect 6542 3744 6560 3752
rect 6542 3733 6546 3744
rect 6442 3676 6475 3680
rect 6441 3656 6443 3668
rect 6439 3644 6443 3656
rect 6449 3656 6451 3668
rect 6449 3644 6453 3656
rect 6471 3644 6475 3676
rect 6481 3644 6485 3702
rect 6501 3664 6505 3701
rect 6542 3676 6546 3721
rect 6564 3699 6568 3756
rect 6586 3753 6590 3796
rect 6586 3741 6593 3753
rect 6566 3687 6575 3699
rect 6542 3669 6555 3676
rect 6551 3664 6555 3669
rect 6571 3664 6575 3687
rect 6591 3664 6595 3741
rect 6651 3719 6655 3796
rect 6646 3707 6655 3719
rect 6649 3691 6655 3707
rect 6671 3719 6675 3796
rect 6671 3707 6674 3719
rect 6671 3691 6677 3707
rect 6649 3684 6657 3691
rect 6653 3664 6657 3684
rect 6663 3684 6677 3691
rect 6663 3664 6667 3684
rect 43 3620 47 3624
rect 65 3620 69 3624
rect 123 3620 127 3624
rect 145 3620 149 3624
rect 213 3620 217 3624
rect 223 3620 227 3624
rect 271 3620 275 3624
rect 293 3620 297 3624
rect 303 3620 307 3624
rect 323 3620 327 3624
rect 331 3620 335 3624
rect 377 3620 381 3624
rect 399 3620 403 3624
rect 409 3620 413 3624
rect 431 3620 435 3624
rect 441 3620 445 3624
rect 461 3620 465 3624
rect 532 3620 536 3624
rect 554 3620 558 3624
rect 562 3620 566 3624
rect 633 3620 637 3624
rect 643 3620 647 3624
rect 693 3620 697 3624
rect 703 3620 707 3624
rect 793 3620 797 3624
rect 803 3620 807 3624
rect 851 3620 855 3624
rect 873 3620 877 3624
rect 883 3620 887 3624
rect 903 3620 907 3624
rect 911 3620 915 3624
rect 957 3620 961 3624
rect 979 3620 983 3624
rect 989 3620 993 3624
rect 1011 3620 1015 3624
rect 1021 3620 1025 3624
rect 1041 3620 1045 3624
rect 1094 3620 1098 3624
rect 1102 3620 1106 3624
rect 1124 3620 1128 3624
rect 1213 3620 1217 3624
rect 1223 3620 1227 3624
rect 1271 3620 1275 3624
rect 1293 3620 1297 3624
rect 1372 3620 1376 3624
rect 1394 3620 1398 3624
rect 1402 3620 1406 3624
rect 1473 3620 1477 3624
rect 1483 3620 1487 3624
rect 1533 3620 1537 3624
rect 1543 3620 1547 3624
rect 1611 3620 1615 3624
rect 1631 3620 1635 3624
rect 1691 3620 1695 3624
rect 1713 3620 1717 3624
rect 1723 3620 1727 3624
rect 1743 3620 1747 3624
rect 1751 3620 1755 3624
rect 1797 3620 1801 3624
rect 1819 3620 1823 3624
rect 1829 3620 1833 3624
rect 1851 3620 1855 3624
rect 1861 3620 1865 3624
rect 1881 3620 1885 3624
rect 1953 3620 1957 3624
rect 1963 3620 1967 3624
rect 2011 3620 2015 3624
rect 2031 3620 2035 3624
rect 2091 3620 2095 3624
rect 2151 3620 2155 3624
rect 2171 3620 2175 3624
rect 2191 3620 2195 3624
rect 2265 3620 2269 3624
rect 2285 3620 2289 3624
rect 2305 3620 2309 3624
rect 2372 3620 2376 3624
rect 2394 3620 2398 3624
rect 2402 3620 2406 3624
rect 2451 3620 2455 3624
rect 2525 3620 2529 3624
rect 2571 3620 2575 3624
rect 2591 3620 2595 3624
rect 2611 3620 2615 3624
rect 2672 3620 2676 3624
rect 2680 3620 2684 3624
rect 2688 3620 2692 3624
rect 2785 3620 2789 3624
rect 2853 3620 2857 3624
rect 2863 3620 2867 3624
rect 2911 3620 2915 3624
rect 2931 3620 2935 3624
rect 2951 3620 2955 3624
rect 3011 3620 3015 3624
rect 3031 3620 3035 3624
rect 3051 3620 3055 3624
rect 3114 3620 3118 3624
rect 3122 3620 3126 3624
rect 3144 3620 3148 3624
rect 3246 3620 3250 3624
rect 3254 3620 3258 3624
rect 3274 3620 3278 3624
rect 3282 3620 3286 3624
rect 3353 3620 3357 3624
rect 3363 3620 3367 3624
rect 3433 3620 3437 3624
rect 3443 3620 3447 3624
rect 3495 3620 3499 3624
rect 3515 3620 3519 3624
rect 3525 3620 3529 3624
rect 3547 3620 3551 3624
rect 3557 3620 3561 3624
rect 3579 3620 3583 3624
rect 3625 3620 3629 3624
rect 3633 3620 3637 3624
rect 3653 3620 3657 3624
rect 3663 3620 3667 3624
rect 3685 3620 3689 3624
rect 3753 3620 3757 3624
rect 3763 3620 3767 3624
rect 3846 3620 3850 3624
rect 3854 3620 3858 3624
rect 3874 3620 3878 3624
rect 3882 3620 3886 3624
rect 3931 3620 3935 3624
rect 3993 3620 3997 3624
rect 4003 3620 4007 3624
rect 4071 3620 4075 3624
rect 4091 3620 4095 3624
rect 4111 3620 4115 3624
rect 4175 3620 4179 3624
rect 4195 3620 4199 3624
rect 4205 3620 4209 3624
rect 4227 3620 4231 3624
rect 4237 3620 4241 3624
rect 4259 3620 4263 3624
rect 4305 3620 4309 3624
rect 4313 3620 4317 3624
rect 4333 3620 4337 3624
rect 4343 3620 4347 3624
rect 4365 3620 4369 3624
rect 4413 3620 4417 3624
rect 4423 3620 4427 3624
rect 4513 3620 4517 3624
rect 4523 3620 4527 3624
rect 4585 3620 4589 3624
rect 4605 3620 4609 3624
rect 4625 3620 4629 3624
rect 4645 3620 4649 3624
rect 4665 3620 4669 3624
rect 4685 3620 4689 3624
rect 4705 3620 4709 3624
rect 4725 3620 4729 3624
rect 4775 3620 4779 3624
rect 4795 3620 4799 3624
rect 4805 3620 4809 3624
rect 4827 3620 4831 3624
rect 4837 3620 4841 3624
rect 4859 3620 4863 3624
rect 4905 3620 4909 3624
rect 4913 3620 4917 3624
rect 4933 3620 4937 3624
rect 4943 3620 4947 3624
rect 4965 3620 4969 3624
rect 5011 3620 5015 3624
rect 5031 3620 5035 3624
rect 5051 3620 5055 3624
rect 5133 3620 5137 3624
rect 5143 3620 5147 3624
rect 5213 3620 5217 3624
rect 5223 3620 5227 3624
rect 5285 3620 5289 3624
rect 5331 3620 5335 3624
rect 5351 3620 5355 3624
rect 5371 3620 5375 3624
rect 5391 3620 5395 3624
rect 5411 3620 5415 3624
rect 5431 3620 5435 3624
rect 5451 3620 5455 3624
rect 5471 3620 5475 3624
rect 5531 3620 5535 3624
rect 5553 3620 5557 3624
rect 5563 3620 5567 3624
rect 5583 3620 5587 3624
rect 5591 3620 5595 3624
rect 5637 3620 5641 3624
rect 5659 3620 5663 3624
rect 5669 3620 5673 3624
rect 5691 3620 5695 3624
rect 5701 3620 5705 3624
rect 5721 3620 5725 3624
rect 5785 3620 5789 3624
rect 5833 3620 5837 3624
rect 5843 3620 5847 3624
rect 5913 3620 5917 3624
rect 5923 3620 5927 3624
rect 6005 3620 6009 3624
rect 6051 3620 6055 3624
rect 6071 3620 6075 3624
rect 6145 3620 6149 3624
rect 6165 3620 6169 3624
rect 6214 3620 6218 3624
rect 6222 3620 6226 3624
rect 6244 3620 6248 3624
rect 6311 3620 6315 3624
rect 6333 3620 6337 3624
rect 6343 3620 6347 3624
rect 6363 3620 6367 3624
rect 6371 3620 6375 3624
rect 6417 3620 6421 3624
rect 6439 3620 6443 3624
rect 6449 3620 6453 3624
rect 6471 3620 6475 3624
rect 6481 3620 6485 3624
rect 6501 3620 6505 3624
rect 6551 3620 6555 3624
rect 6571 3620 6575 3624
rect 6591 3620 6595 3624
rect 6653 3620 6657 3624
rect 6663 3620 6667 3624
rect 43 3596 47 3600
rect 65 3596 69 3600
rect 111 3596 115 3600
rect 133 3596 137 3600
rect 143 3596 147 3600
rect 163 3596 167 3600
rect 171 3596 175 3600
rect 217 3596 221 3600
rect 239 3596 243 3600
rect 249 3596 253 3600
rect 271 3596 275 3600
rect 281 3596 285 3600
rect 301 3596 305 3600
rect 353 3596 357 3600
rect 363 3596 367 3600
rect 431 3596 435 3600
rect 453 3596 457 3600
rect 532 3596 536 3600
rect 554 3596 558 3600
rect 562 3596 566 3600
rect 633 3596 637 3600
rect 643 3596 647 3600
rect 703 3596 707 3600
rect 725 3596 729 3600
rect 771 3596 775 3600
rect 793 3596 797 3600
rect 853 3596 857 3600
rect 863 3596 867 3600
rect 943 3596 947 3600
rect 965 3596 969 3600
rect 1025 3596 1029 3600
rect 1083 3596 1087 3600
rect 1105 3596 1109 3600
rect 1163 3596 1167 3600
rect 1185 3596 1189 3600
rect 1231 3596 1235 3600
rect 1253 3596 1257 3600
rect 1263 3596 1267 3600
rect 1283 3596 1287 3600
rect 1291 3596 1295 3600
rect 1337 3596 1341 3600
rect 1359 3596 1363 3600
rect 1369 3596 1373 3600
rect 1391 3596 1395 3600
rect 1401 3596 1405 3600
rect 1421 3596 1425 3600
rect 1485 3596 1489 3600
rect 1505 3596 1509 3600
rect 1551 3596 1555 3600
rect 1573 3596 1577 3600
rect 1583 3596 1587 3600
rect 1603 3596 1607 3600
rect 1611 3596 1615 3600
rect 1657 3596 1661 3600
rect 1679 3596 1683 3600
rect 1689 3596 1693 3600
rect 1711 3596 1715 3600
rect 1721 3596 1725 3600
rect 1741 3596 1745 3600
rect 1815 3596 1819 3600
rect 1835 3596 1839 3600
rect 1845 3596 1849 3600
rect 1905 3596 1909 3600
rect 1965 3596 1969 3600
rect 1985 3596 1989 3600
rect 2005 3596 2009 3600
rect 2051 3596 2055 3600
rect 2071 3596 2075 3600
rect 2145 3596 2149 3600
rect 2215 3596 2219 3600
rect 2235 3596 2239 3600
rect 2245 3596 2249 3600
rect 2305 3596 2309 3600
rect 2325 3596 2329 3600
rect 2371 3596 2375 3600
rect 2393 3596 2397 3600
rect 2403 3596 2407 3600
rect 2423 3596 2427 3600
rect 2431 3596 2435 3600
rect 2477 3596 2481 3600
rect 2499 3596 2503 3600
rect 2509 3596 2513 3600
rect 2531 3596 2535 3600
rect 2541 3596 2545 3600
rect 2561 3596 2565 3600
rect 2611 3596 2615 3600
rect 2631 3596 2635 3600
rect 2691 3596 2695 3600
rect 2711 3596 2715 3600
rect 2731 3596 2735 3600
rect 2805 3596 2809 3600
rect 2873 3596 2877 3600
rect 2883 3596 2887 3600
rect 2931 3596 2935 3600
rect 2951 3596 2955 3600
rect 2971 3596 2975 3600
rect 3034 3596 3038 3600
rect 3042 3596 3046 3600
rect 3064 3596 3068 3600
rect 3131 3596 3135 3600
rect 3226 3596 3230 3600
rect 3234 3596 3238 3600
rect 3254 3596 3258 3600
rect 3262 3596 3266 3600
rect 3325 3596 3329 3600
rect 3371 3596 3375 3600
rect 3393 3596 3397 3600
rect 3403 3596 3407 3600
rect 3423 3596 3427 3600
rect 3431 3596 3435 3600
rect 3477 3596 3481 3600
rect 3499 3596 3503 3600
rect 3509 3596 3513 3600
rect 3531 3596 3535 3600
rect 3541 3596 3545 3600
rect 3561 3596 3565 3600
rect 3646 3596 3650 3600
rect 3654 3596 3658 3600
rect 3674 3596 3678 3600
rect 3682 3596 3686 3600
rect 3731 3596 3735 3600
rect 3753 3596 3757 3600
rect 3763 3596 3767 3600
rect 3783 3596 3787 3600
rect 3791 3596 3795 3600
rect 3837 3596 3841 3600
rect 3859 3596 3863 3600
rect 3869 3596 3873 3600
rect 3891 3596 3895 3600
rect 3901 3596 3905 3600
rect 3921 3596 3925 3600
rect 3985 3596 3989 3600
rect 4031 3596 4035 3600
rect 4053 3596 4057 3600
rect 4063 3596 4067 3600
rect 4083 3596 4087 3600
rect 4091 3596 4095 3600
rect 4137 3596 4141 3600
rect 4159 3596 4163 3600
rect 4169 3596 4173 3600
rect 4191 3596 4195 3600
rect 4201 3596 4205 3600
rect 4221 3596 4225 3600
rect 4285 3596 4289 3600
rect 4345 3596 4349 3600
rect 4393 3596 4397 3600
rect 4403 3596 4407 3600
rect 4475 3596 4479 3600
rect 4495 3596 4499 3600
rect 4505 3596 4509 3600
rect 4527 3596 4531 3600
rect 4537 3596 4541 3600
rect 4559 3596 4563 3600
rect 4605 3596 4609 3600
rect 4613 3596 4617 3600
rect 4633 3596 4637 3600
rect 4643 3596 4647 3600
rect 4665 3596 4669 3600
rect 4725 3596 4729 3600
rect 4771 3596 4775 3600
rect 4793 3596 4797 3600
rect 4803 3596 4807 3600
rect 4823 3596 4827 3600
rect 4831 3596 4835 3600
rect 4877 3596 4881 3600
rect 4899 3596 4903 3600
rect 4909 3596 4913 3600
rect 4931 3596 4935 3600
rect 4941 3596 4945 3600
rect 4961 3596 4965 3600
rect 5046 3596 5050 3600
rect 5054 3596 5058 3600
rect 5074 3596 5078 3600
rect 5082 3596 5086 3600
rect 5145 3596 5149 3600
rect 5191 3596 5195 3600
rect 5213 3596 5217 3600
rect 5223 3596 5227 3600
rect 5243 3596 5247 3600
rect 5251 3596 5255 3600
rect 5297 3596 5301 3600
rect 5319 3596 5323 3600
rect 5329 3596 5333 3600
rect 5351 3596 5355 3600
rect 5361 3596 5365 3600
rect 5381 3596 5385 3600
rect 5431 3596 5435 3600
rect 5453 3596 5457 3600
rect 5463 3596 5467 3600
rect 5483 3596 5487 3600
rect 5491 3596 5495 3600
rect 5537 3596 5541 3600
rect 5559 3596 5563 3600
rect 5569 3596 5573 3600
rect 5591 3596 5595 3600
rect 5601 3596 5605 3600
rect 5621 3596 5625 3600
rect 5671 3596 5675 3600
rect 5691 3596 5695 3600
rect 5711 3596 5715 3600
rect 5771 3596 5775 3600
rect 5791 3596 5795 3600
rect 5811 3596 5815 3600
rect 5885 3596 5889 3600
rect 5966 3596 5970 3600
rect 5974 3596 5978 3600
rect 5994 3596 5998 3600
rect 6002 3596 6006 3600
rect 6053 3596 6057 3600
rect 6063 3596 6067 3600
rect 6145 3596 6149 3600
rect 6211 3596 6215 3600
rect 6231 3596 6235 3600
rect 6251 3596 6255 3600
rect 6385 3596 6389 3600
rect 6431 3596 6435 3600
rect 6453 3596 6457 3600
rect 6463 3596 6467 3600
rect 6483 3596 6487 3600
rect 6491 3596 6495 3600
rect 6537 3596 6541 3600
rect 6559 3596 6563 3600
rect 6569 3596 6573 3600
rect 6591 3596 6595 3600
rect 6601 3596 6605 3600
rect 6621 3596 6625 3600
rect 43 3550 47 3556
rect 43 3538 45 3550
rect 65 3499 69 3576
rect 65 3487 74 3499
rect 111 3488 115 3556
rect 133 3527 137 3576
rect 143 3555 147 3576
rect 163 3564 167 3576
rect 171 3572 175 3576
rect 171 3568 205 3572
rect 163 3560 193 3564
rect 163 3559 181 3560
rect 143 3551 167 3555
rect 43 3470 45 3482
rect 43 3464 47 3470
rect 65 3424 69 3487
rect 111 3476 113 3488
rect 111 3464 115 3476
rect 133 3469 137 3515
rect 129 3463 137 3469
rect 129 3434 133 3463
rect 161 3456 167 3551
rect 129 3427 137 3434
rect 133 3404 137 3427
rect 141 3404 145 3444
rect 161 3424 165 3456
rect 201 3442 205 3568
rect 217 3462 221 3576
rect 239 3564 243 3576
rect 241 3552 243 3564
rect 249 3564 253 3576
rect 249 3552 251 3564
rect 169 3430 193 3432
rect 169 3428 205 3430
rect 169 3424 173 3428
rect 215 3424 219 3450
rect 233 3442 237 3552
rect 271 3544 275 3576
rect 242 3540 275 3544
rect 242 3476 246 3540
rect 262 3491 266 3520
rect 281 3518 285 3576
rect 301 3519 305 3556
rect 353 3536 357 3556
rect 349 3529 357 3536
rect 363 3536 367 3556
rect 363 3529 377 3536
rect 349 3513 355 3529
rect 262 3483 271 3491
rect 242 3464 245 3476
rect 235 3424 239 3430
rect 247 3424 251 3464
rect 267 3424 271 3483
rect 281 3424 285 3506
rect 301 3464 305 3507
rect 346 3501 355 3513
rect 351 3424 355 3501
rect 371 3513 377 3529
rect 371 3501 374 3513
rect 371 3424 375 3501
rect 431 3499 435 3576
rect 453 3550 457 3556
rect 455 3538 457 3550
rect 532 3533 536 3576
rect 426 3487 435 3499
rect 431 3424 435 3487
rect 525 3521 534 3533
rect 455 3470 457 3482
rect 453 3464 457 3470
rect 525 3464 529 3521
rect 554 3519 558 3556
rect 562 3552 566 3556
rect 562 3546 581 3552
rect 574 3533 581 3546
rect 633 3536 637 3556
rect 623 3529 637 3536
rect 643 3536 647 3556
rect 703 3550 707 3556
rect 703 3538 705 3550
rect 643 3529 651 3536
rect 554 3484 560 3507
rect 574 3484 581 3521
rect 623 3513 629 3529
rect 626 3501 629 3513
rect 545 3478 560 3484
rect 565 3478 581 3484
rect 545 3464 549 3478
rect 565 3464 569 3478
rect 625 3424 629 3501
rect 645 3513 651 3529
rect 645 3501 654 3513
rect 645 3424 649 3501
rect 725 3499 729 3576
rect 771 3499 775 3576
rect 793 3550 797 3556
rect 795 3538 797 3550
rect 853 3536 857 3556
rect 849 3529 857 3536
rect 863 3536 867 3556
rect 943 3550 947 3556
rect 943 3538 945 3550
rect 863 3529 877 3536
rect 849 3513 855 3529
rect 846 3501 855 3513
rect 725 3487 734 3499
rect 766 3487 775 3499
rect 703 3470 705 3482
rect 703 3464 707 3470
rect 725 3424 729 3487
rect 771 3424 775 3487
rect 795 3470 797 3482
rect 793 3464 797 3470
rect 851 3424 855 3501
rect 871 3513 877 3529
rect 871 3501 874 3513
rect 871 3424 875 3501
rect 965 3499 969 3576
rect 1025 3519 1029 3576
rect 1083 3550 1087 3556
rect 1083 3538 1085 3550
rect 1025 3507 1034 3519
rect 965 3487 974 3499
rect 943 3470 945 3482
rect 943 3464 947 3470
rect 965 3424 969 3487
rect 1025 3424 1029 3507
rect 1105 3499 1109 3576
rect 1163 3550 1167 3556
rect 1163 3538 1165 3550
rect 1185 3499 1189 3576
rect 1105 3487 1114 3499
rect 1185 3487 1194 3499
rect 1231 3488 1235 3556
rect 1253 3527 1257 3576
rect 1263 3555 1267 3576
rect 1283 3564 1287 3576
rect 1291 3572 1295 3576
rect 1291 3568 1325 3572
rect 1283 3560 1313 3564
rect 1283 3559 1301 3560
rect 1263 3551 1287 3555
rect 1083 3470 1085 3482
rect 1083 3464 1087 3470
rect 1105 3424 1109 3487
rect 1163 3470 1165 3482
rect 1163 3464 1167 3470
rect 1185 3424 1189 3487
rect 1231 3476 1233 3488
rect 1231 3464 1235 3476
rect 1253 3469 1257 3515
rect 1249 3463 1257 3469
rect 1249 3434 1253 3463
rect 1281 3456 1287 3551
rect 1249 3427 1257 3434
rect 1253 3404 1257 3427
rect 1261 3404 1265 3444
rect 1281 3424 1285 3456
rect 1321 3442 1325 3568
rect 1337 3462 1341 3576
rect 1359 3564 1363 3576
rect 1361 3552 1363 3564
rect 1369 3564 1373 3576
rect 1369 3552 1371 3564
rect 1289 3430 1313 3432
rect 1289 3428 1325 3430
rect 1289 3424 1293 3428
rect 1335 3424 1339 3450
rect 1353 3442 1357 3552
rect 1391 3544 1395 3576
rect 1362 3540 1395 3544
rect 1362 3476 1366 3540
rect 1382 3491 1386 3520
rect 1401 3518 1405 3576
rect 1421 3519 1425 3556
rect 1382 3483 1391 3491
rect 1362 3464 1365 3476
rect 1355 3424 1359 3430
rect 1367 3424 1371 3464
rect 1387 3424 1391 3483
rect 1401 3424 1405 3506
rect 1421 3464 1425 3507
rect 1485 3499 1489 3576
rect 1505 3499 1509 3576
rect 1486 3487 1501 3499
rect 1497 3464 1501 3487
rect 1505 3487 1514 3499
rect 1551 3488 1555 3556
rect 1573 3527 1577 3576
rect 1583 3555 1587 3576
rect 1603 3564 1607 3576
rect 1611 3572 1615 3576
rect 1611 3568 1645 3572
rect 1603 3560 1633 3564
rect 1603 3559 1621 3560
rect 1583 3551 1607 3555
rect 1505 3464 1509 3487
rect 1551 3476 1553 3488
rect 1551 3464 1555 3476
rect 1573 3469 1577 3515
rect 1569 3463 1577 3469
rect 1569 3434 1573 3463
rect 1601 3456 1607 3551
rect 1569 3427 1577 3434
rect 1573 3404 1577 3427
rect 1581 3404 1585 3444
rect 1601 3424 1605 3456
rect 1641 3442 1645 3568
rect 1657 3462 1661 3576
rect 1679 3564 1683 3576
rect 1681 3552 1683 3564
rect 1689 3564 1693 3576
rect 1689 3552 1691 3564
rect 1609 3430 1633 3432
rect 1609 3428 1645 3430
rect 1609 3424 1613 3428
rect 1655 3424 1659 3450
rect 1673 3442 1677 3552
rect 1711 3544 1715 3576
rect 1682 3540 1715 3544
rect 1682 3476 1686 3540
rect 1702 3491 1706 3520
rect 1721 3518 1725 3576
rect 1741 3519 1745 3556
rect 1815 3550 1819 3556
rect 1801 3538 1813 3550
rect 1702 3483 1711 3491
rect 1682 3464 1685 3476
rect 1675 3424 1679 3430
rect 1687 3424 1691 3464
rect 1707 3424 1711 3483
rect 1721 3424 1725 3506
rect 1741 3464 1745 3507
rect 1801 3464 1805 3538
rect 1835 3513 1839 3556
rect 1826 3501 1839 3513
rect 1823 3424 1827 3501
rect 1845 3499 1849 3556
rect 1905 3519 1909 3576
rect 1905 3507 1914 3519
rect 1845 3487 1854 3499
rect 1845 3424 1849 3487
rect 1905 3424 1909 3507
rect 1965 3479 1969 3556
rect 1985 3533 1989 3556
rect 2005 3551 2009 3556
rect 2005 3544 2018 3551
rect 1985 3521 1994 3533
rect 1967 3467 1974 3479
rect 1970 3424 1974 3467
rect 1992 3464 1996 3521
rect 2014 3499 2018 3544
rect 2051 3499 2055 3576
rect 2071 3499 2075 3576
rect 2145 3519 2149 3576
rect 2215 3550 2219 3556
rect 2201 3538 2213 3550
rect 2145 3507 2154 3519
rect 2046 3487 2055 3499
rect 2014 3476 2018 3487
rect 2000 3468 2018 3476
rect 2000 3464 2004 3468
rect 2051 3464 2055 3487
rect 2059 3487 2074 3499
rect 2059 3464 2063 3487
rect 2145 3424 2149 3507
rect 2201 3464 2205 3538
rect 2235 3513 2239 3556
rect 2226 3501 2239 3513
rect 2223 3424 2227 3501
rect 2245 3499 2249 3556
rect 2305 3499 2309 3576
rect 2325 3499 2329 3576
rect 2245 3487 2254 3499
rect 2306 3487 2321 3499
rect 2245 3424 2249 3487
rect 2317 3464 2321 3487
rect 2325 3487 2334 3499
rect 2371 3488 2375 3556
rect 2393 3527 2397 3576
rect 2403 3555 2407 3576
rect 2423 3564 2427 3576
rect 2431 3572 2435 3576
rect 2431 3568 2465 3572
rect 2423 3560 2453 3564
rect 2423 3559 2441 3560
rect 2403 3551 2427 3555
rect 2325 3464 2329 3487
rect 2371 3476 2373 3488
rect 2371 3464 2375 3476
rect 2393 3469 2397 3515
rect 2389 3463 2397 3469
rect 2389 3434 2393 3463
rect 2421 3456 2427 3551
rect 2389 3427 2397 3434
rect 2393 3404 2397 3427
rect 2401 3404 2405 3444
rect 2421 3424 2425 3456
rect 2461 3442 2465 3568
rect 2477 3462 2481 3576
rect 2499 3564 2503 3576
rect 2501 3552 2503 3564
rect 2509 3564 2513 3576
rect 2509 3552 2511 3564
rect 2429 3430 2453 3432
rect 2429 3428 2465 3430
rect 2429 3424 2433 3428
rect 2475 3424 2479 3450
rect 2493 3442 2497 3552
rect 2531 3544 2535 3576
rect 2502 3540 2535 3544
rect 2502 3476 2506 3540
rect 2522 3491 2526 3520
rect 2541 3518 2545 3576
rect 2561 3519 2565 3556
rect 2522 3483 2531 3491
rect 2502 3464 2505 3476
rect 2495 3424 2499 3430
rect 2507 3424 2511 3464
rect 2527 3424 2531 3483
rect 2541 3424 2545 3506
rect 2561 3464 2565 3507
rect 2611 3499 2615 3576
rect 2631 3499 2635 3576
rect 2691 3551 2695 3556
rect 2682 3544 2695 3551
rect 2682 3499 2686 3544
rect 2711 3533 2715 3556
rect 2706 3521 2715 3533
rect 2606 3487 2615 3499
rect 2611 3464 2615 3487
rect 2619 3487 2634 3499
rect 2619 3464 2623 3487
rect 2682 3476 2686 3487
rect 2682 3468 2700 3476
rect 2696 3464 2700 3468
rect 2704 3464 2708 3521
rect 2731 3479 2735 3556
rect 2805 3519 2809 3576
rect 2873 3536 2877 3556
rect 2863 3529 2877 3536
rect 2883 3536 2887 3556
rect 2931 3551 2935 3556
rect 2922 3544 2935 3551
rect 2883 3529 2891 3536
rect 2805 3507 2814 3519
rect 2863 3513 2869 3529
rect 2726 3467 2733 3479
rect 2726 3424 2730 3467
rect 2805 3424 2809 3507
rect 2866 3501 2869 3513
rect 2865 3424 2869 3501
rect 2885 3513 2891 3529
rect 2885 3501 2894 3513
rect 2885 3424 2889 3501
rect 2922 3499 2926 3544
rect 2951 3533 2955 3556
rect 2946 3521 2955 3533
rect 2922 3476 2926 3487
rect 2922 3468 2940 3476
rect 2936 3464 2940 3468
rect 2944 3464 2948 3521
rect 2971 3479 2975 3556
rect 3034 3552 3038 3556
rect 3019 3546 3038 3552
rect 3019 3533 3026 3546
rect 3019 3484 3026 3521
rect 3042 3519 3046 3556
rect 3064 3533 3068 3576
rect 3131 3533 3135 3556
rect 3226 3551 3230 3556
rect 3066 3521 3075 3533
rect 3126 3521 3135 3533
rect 3040 3484 3046 3507
rect 2966 3467 2973 3479
rect 3019 3478 3035 3484
rect 3040 3478 3055 3484
rect 2966 3424 2970 3467
rect 3031 3464 3035 3478
rect 3051 3464 3055 3478
rect 3071 3464 3075 3521
rect 3131 3464 3135 3521
rect 3200 3547 3230 3551
rect 3200 3499 3206 3547
rect 3234 3542 3238 3556
rect 3225 3535 3238 3542
rect 3225 3533 3229 3535
rect 3254 3533 3258 3556
rect 3262 3548 3266 3556
rect 3262 3541 3279 3548
rect 3227 3521 3229 3533
rect 3206 3487 3209 3499
rect 3205 3464 3209 3487
rect 3225 3464 3229 3521
rect 3254 3492 3258 3521
rect 3273 3499 3279 3541
rect 3325 3519 3329 3576
rect 3325 3507 3334 3519
rect 3245 3486 3258 3492
rect 3265 3487 3273 3492
rect 3265 3486 3285 3487
rect 3245 3464 3249 3486
rect 3265 3464 3269 3486
rect 3325 3424 3329 3507
rect 3371 3488 3375 3556
rect 3393 3527 3397 3576
rect 3403 3555 3407 3576
rect 3423 3564 3427 3576
rect 3431 3572 3435 3576
rect 3431 3568 3465 3572
rect 3423 3560 3453 3564
rect 3423 3559 3441 3560
rect 3403 3551 3427 3555
rect 3371 3476 3373 3488
rect 3371 3464 3375 3476
rect 3393 3469 3397 3515
rect 3389 3463 3397 3469
rect 3389 3434 3393 3463
rect 3421 3456 3427 3551
rect 3389 3427 3397 3434
rect 3393 3404 3397 3427
rect 3401 3404 3405 3444
rect 3421 3424 3425 3456
rect 3461 3442 3465 3568
rect 3477 3462 3481 3576
rect 3499 3564 3503 3576
rect 3501 3552 3503 3564
rect 3509 3564 3513 3576
rect 3509 3552 3511 3564
rect 3429 3430 3453 3432
rect 3429 3428 3465 3430
rect 3429 3424 3433 3428
rect 3475 3424 3479 3450
rect 3493 3442 3497 3552
rect 3531 3544 3535 3576
rect 3502 3540 3535 3544
rect 3502 3476 3506 3540
rect 3522 3491 3526 3520
rect 3541 3518 3545 3576
rect 3561 3519 3565 3556
rect 3646 3551 3650 3556
rect 3620 3547 3650 3551
rect 3522 3483 3531 3491
rect 3502 3464 3505 3476
rect 3495 3424 3499 3430
rect 3507 3424 3511 3464
rect 3527 3424 3531 3483
rect 3541 3424 3545 3506
rect 3561 3464 3565 3507
rect 3620 3499 3626 3547
rect 3654 3542 3658 3556
rect 3645 3535 3658 3542
rect 3645 3533 3649 3535
rect 3674 3533 3678 3556
rect 3682 3548 3686 3556
rect 3682 3541 3699 3548
rect 3647 3521 3649 3533
rect 3626 3487 3629 3499
rect 3625 3464 3629 3487
rect 3645 3464 3649 3521
rect 3674 3492 3678 3521
rect 3693 3499 3699 3541
rect 3665 3486 3678 3492
rect 3685 3487 3693 3492
rect 3685 3486 3705 3487
rect 3731 3488 3735 3556
rect 3753 3527 3757 3576
rect 3763 3555 3767 3576
rect 3783 3564 3787 3576
rect 3791 3572 3795 3576
rect 3791 3568 3825 3572
rect 3783 3560 3813 3564
rect 3783 3559 3801 3560
rect 3763 3551 3787 3555
rect 3665 3464 3669 3486
rect 3685 3464 3689 3486
rect 3731 3476 3733 3488
rect 3731 3464 3735 3476
rect 3753 3469 3757 3515
rect 3749 3463 3757 3469
rect 3749 3434 3753 3463
rect 3781 3456 3787 3551
rect 3749 3427 3757 3434
rect 3753 3404 3757 3427
rect 3761 3404 3765 3444
rect 3781 3424 3785 3456
rect 3821 3442 3825 3568
rect 3837 3462 3841 3576
rect 3859 3564 3863 3576
rect 3861 3552 3863 3564
rect 3869 3564 3873 3576
rect 3869 3552 3871 3564
rect 3789 3430 3813 3432
rect 3789 3428 3825 3430
rect 3789 3424 3793 3428
rect 3835 3424 3839 3450
rect 3853 3442 3857 3552
rect 3891 3544 3895 3576
rect 3862 3540 3895 3544
rect 3862 3476 3866 3540
rect 3882 3491 3886 3520
rect 3901 3518 3905 3576
rect 3921 3519 3925 3556
rect 3985 3519 3989 3576
rect 3985 3507 3994 3519
rect 3882 3483 3891 3491
rect 3862 3464 3865 3476
rect 3855 3424 3859 3430
rect 3867 3424 3871 3464
rect 3887 3424 3891 3483
rect 3901 3424 3905 3506
rect 3921 3464 3925 3507
rect 3985 3424 3989 3507
rect 4031 3488 4035 3556
rect 4053 3527 4057 3576
rect 4063 3555 4067 3576
rect 4083 3564 4087 3576
rect 4091 3572 4095 3576
rect 4091 3568 4125 3572
rect 4083 3560 4113 3564
rect 4083 3559 4101 3560
rect 4063 3551 4087 3555
rect 4031 3476 4033 3488
rect 4031 3464 4035 3476
rect 4053 3469 4057 3515
rect 4049 3463 4057 3469
rect 4049 3434 4053 3463
rect 4081 3456 4087 3551
rect 4049 3427 4057 3434
rect 4053 3404 4057 3427
rect 4061 3404 4065 3444
rect 4081 3424 4085 3456
rect 4121 3442 4125 3568
rect 4137 3462 4141 3576
rect 4159 3564 4163 3576
rect 4161 3552 4163 3564
rect 4169 3564 4173 3576
rect 4169 3552 4171 3564
rect 4089 3430 4113 3432
rect 4089 3428 4125 3430
rect 4089 3424 4093 3428
rect 4135 3424 4139 3450
rect 4153 3442 4157 3552
rect 4191 3544 4195 3576
rect 4162 3540 4195 3544
rect 4162 3476 4166 3540
rect 4182 3491 4186 3520
rect 4201 3518 4205 3576
rect 4221 3519 4225 3556
rect 4285 3519 4289 3576
rect 4345 3519 4349 3576
rect 4393 3536 4397 3556
rect 4389 3529 4397 3536
rect 4403 3536 4407 3556
rect 4403 3529 4417 3536
rect 4285 3507 4294 3519
rect 4345 3507 4354 3519
rect 4389 3513 4395 3529
rect 4182 3483 4191 3491
rect 4162 3464 4165 3476
rect 4155 3424 4159 3430
rect 4167 3424 4171 3464
rect 4187 3424 4191 3483
rect 4201 3424 4205 3506
rect 4221 3464 4225 3507
rect 4285 3424 4289 3507
rect 4345 3424 4349 3507
rect 4386 3501 4395 3513
rect 4391 3424 4395 3501
rect 4411 3513 4417 3529
rect 4475 3519 4479 3556
rect 4411 3501 4414 3513
rect 4495 3518 4499 3576
rect 4505 3544 4509 3576
rect 4527 3564 4531 3576
rect 4529 3552 4531 3564
rect 4537 3564 4541 3576
rect 4537 3552 4539 3564
rect 4505 3540 4538 3544
rect 4411 3424 4415 3501
rect 4475 3464 4479 3507
rect 4495 3424 4499 3506
rect 4514 3491 4518 3520
rect 4509 3483 4518 3491
rect 4509 3424 4513 3483
rect 4534 3476 4538 3540
rect 4535 3464 4538 3476
rect 4529 3424 4533 3464
rect 4543 3442 4547 3552
rect 4559 3462 4563 3576
rect 4605 3572 4609 3576
rect 4575 3568 4609 3572
rect 4541 3424 4545 3430
rect 4561 3424 4565 3450
rect 4575 3442 4579 3568
rect 4613 3564 4617 3576
rect 4587 3560 4617 3564
rect 4599 3559 4617 3560
rect 4633 3555 4637 3576
rect 4613 3551 4637 3555
rect 4613 3456 4619 3551
rect 4643 3527 4647 3576
rect 4643 3469 4647 3515
rect 4665 3488 4669 3556
rect 4667 3476 4669 3488
rect 4643 3463 4651 3469
rect 4665 3464 4669 3476
rect 4725 3519 4729 3576
rect 4725 3507 4734 3519
rect 4587 3430 4611 3432
rect 4575 3428 4611 3430
rect 4607 3424 4611 3428
rect 4615 3424 4619 3456
rect 4635 3404 4639 3444
rect 4647 3434 4651 3463
rect 4643 3427 4651 3434
rect 4643 3404 4647 3427
rect 4725 3424 4729 3507
rect 4771 3488 4775 3556
rect 4793 3527 4797 3576
rect 4803 3555 4807 3576
rect 4823 3564 4827 3576
rect 4831 3572 4835 3576
rect 4831 3568 4865 3572
rect 4823 3560 4853 3564
rect 4823 3559 4841 3560
rect 4803 3551 4827 3555
rect 4771 3476 4773 3488
rect 4771 3464 4775 3476
rect 4793 3469 4797 3515
rect 4789 3463 4797 3469
rect 4789 3434 4793 3463
rect 4821 3456 4827 3551
rect 4789 3427 4797 3434
rect 4793 3404 4797 3427
rect 4801 3404 4805 3444
rect 4821 3424 4825 3456
rect 4861 3442 4865 3568
rect 4877 3462 4881 3576
rect 4899 3564 4903 3576
rect 4901 3552 4903 3564
rect 4909 3564 4913 3576
rect 4909 3552 4911 3564
rect 4829 3430 4853 3432
rect 4829 3428 4865 3430
rect 4829 3424 4833 3428
rect 4875 3424 4879 3450
rect 4893 3442 4897 3552
rect 4931 3544 4935 3576
rect 4902 3540 4935 3544
rect 4902 3476 4906 3540
rect 4922 3491 4926 3520
rect 4941 3518 4945 3576
rect 4961 3519 4965 3556
rect 5046 3551 5050 3556
rect 5020 3547 5050 3551
rect 4922 3483 4931 3491
rect 4902 3464 4905 3476
rect 4895 3424 4899 3430
rect 4907 3424 4911 3464
rect 4927 3424 4931 3483
rect 4941 3424 4945 3506
rect 4961 3464 4965 3507
rect 5020 3499 5026 3547
rect 5054 3542 5058 3556
rect 5045 3535 5058 3542
rect 5045 3533 5049 3535
rect 5074 3533 5078 3556
rect 5082 3548 5086 3556
rect 5082 3541 5099 3548
rect 5047 3521 5049 3533
rect 5026 3487 5029 3499
rect 5025 3464 5029 3487
rect 5045 3464 5049 3521
rect 5074 3492 5078 3521
rect 5093 3499 5099 3541
rect 5145 3519 5149 3576
rect 5145 3507 5154 3519
rect 5065 3486 5078 3492
rect 5085 3487 5093 3492
rect 5085 3486 5105 3487
rect 5065 3464 5069 3486
rect 5085 3464 5089 3486
rect 5145 3424 5149 3507
rect 5191 3488 5195 3556
rect 5213 3527 5217 3576
rect 5223 3555 5227 3576
rect 5243 3564 5247 3576
rect 5251 3572 5255 3576
rect 5251 3568 5285 3572
rect 5243 3560 5273 3564
rect 5243 3559 5261 3560
rect 5223 3551 5247 3555
rect 5191 3476 5193 3488
rect 5191 3464 5195 3476
rect 5213 3469 5217 3515
rect 5209 3463 5217 3469
rect 5209 3434 5213 3463
rect 5241 3456 5247 3551
rect 5209 3427 5217 3434
rect 5213 3404 5217 3427
rect 5221 3404 5225 3444
rect 5241 3424 5245 3456
rect 5281 3442 5285 3568
rect 5297 3462 5301 3576
rect 5319 3564 5323 3576
rect 5321 3552 5323 3564
rect 5329 3564 5333 3576
rect 5329 3552 5331 3564
rect 5249 3430 5273 3432
rect 5249 3428 5285 3430
rect 5249 3424 5253 3428
rect 5295 3424 5299 3450
rect 5313 3442 5317 3552
rect 5351 3544 5355 3576
rect 5322 3540 5355 3544
rect 5322 3476 5326 3540
rect 5342 3491 5346 3520
rect 5361 3518 5365 3576
rect 5381 3519 5385 3556
rect 5342 3483 5351 3491
rect 5322 3464 5325 3476
rect 5315 3424 5319 3430
rect 5327 3424 5331 3464
rect 5347 3424 5351 3483
rect 5361 3424 5365 3506
rect 5381 3464 5385 3507
rect 5431 3488 5435 3556
rect 5453 3527 5457 3576
rect 5463 3555 5467 3576
rect 5483 3564 5487 3576
rect 5491 3572 5495 3576
rect 5491 3568 5525 3572
rect 5483 3560 5513 3564
rect 5483 3559 5501 3560
rect 5463 3551 5487 3555
rect 5431 3476 5433 3488
rect 5431 3464 5435 3476
rect 5453 3469 5457 3515
rect 5449 3463 5457 3469
rect 5449 3434 5453 3463
rect 5481 3456 5487 3551
rect 5449 3427 5457 3434
rect 5453 3404 5457 3427
rect 5461 3404 5465 3444
rect 5481 3424 5485 3456
rect 5521 3442 5525 3568
rect 5537 3462 5541 3576
rect 5559 3564 5563 3576
rect 5561 3552 5563 3564
rect 5569 3564 5573 3576
rect 5569 3552 5571 3564
rect 5489 3430 5513 3432
rect 5489 3428 5525 3430
rect 5489 3424 5493 3428
rect 5535 3424 5539 3450
rect 5553 3442 5557 3552
rect 5591 3544 5595 3576
rect 5562 3540 5595 3544
rect 5562 3476 5566 3540
rect 5582 3491 5586 3520
rect 5601 3518 5605 3576
rect 5621 3519 5625 3556
rect 5671 3551 5675 3556
rect 5662 3544 5675 3551
rect 5582 3483 5591 3491
rect 5562 3464 5565 3476
rect 5555 3424 5559 3430
rect 5567 3424 5571 3464
rect 5587 3424 5591 3483
rect 5601 3424 5605 3506
rect 5621 3464 5625 3507
rect 5662 3499 5666 3544
rect 5691 3533 5695 3556
rect 5686 3521 5695 3533
rect 5662 3476 5666 3487
rect 5662 3468 5680 3476
rect 5676 3464 5680 3468
rect 5684 3464 5688 3521
rect 5711 3479 5715 3556
rect 5771 3551 5775 3556
rect 5762 3544 5775 3551
rect 5762 3499 5766 3544
rect 5791 3533 5795 3556
rect 5786 3521 5795 3533
rect 5706 3467 5713 3479
rect 5762 3476 5766 3487
rect 5762 3468 5780 3476
rect 5706 3424 5710 3467
rect 5776 3464 5780 3468
rect 5784 3464 5788 3521
rect 5811 3479 5815 3556
rect 5885 3519 5889 3576
rect 5966 3551 5970 3556
rect 5940 3547 5970 3551
rect 5885 3507 5894 3519
rect 5806 3467 5813 3479
rect 5806 3424 5810 3467
rect 5885 3424 5889 3507
rect 5940 3499 5946 3547
rect 5974 3542 5978 3556
rect 5965 3535 5978 3542
rect 5965 3533 5969 3535
rect 5994 3533 5998 3556
rect 6002 3548 6006 3556
rect 6002 3541 6019 3548
rect 5967 3521 5969 3533
rect 5946 3487 5949 3499
rect 5945 3464 5949 3487
rect 5965 3464 5969 3521
rect 5994 3492 5998 3521
rect 6013 3499 6019 3541
rect 6053 3536 6057 3556
rect 6049 3529 6057 3536
rect 6063 3536 6067 3556
rect 6063 3529 6077 3536
rect 6049 3513 6055 3529
rect 6046 3501 6055 3513
rect 5985 3486 5998 3492
rect 6005 3487 6013 3492
rect 6005 3486 6025 3487
rect 5985 3464 5989 3486
rect 6005 3464 6009 3486
rect 6051 3424 6055 3501
rect 6071 3513 6077 3529
rect 6145 3519 6149 3576
rect 6071 3501 6074 3513
rect 6145 3507 6154 3519
rect 6071 3424 6075 3501
rect 6145 3424 6149 3507
rect 6211 3499 6215 3576
rect 6206 3487 6215 3499
rect 6211 3452 6215 3487
rect 6191 3448 6215 3452
rect 6191 3444 6195 3448
rect 6211 3444 6215 3448
rect 6231 3533 6235 3576
rect 6251 3560 6255 3576
rect 6251 3554 6275 3560
rect 6231 3521 6234 3533
rect 6231 3452 6235 3521
rect 6269 3499 6275 3554
rect 6266 3487 6275 3499
rect 6269 3464 6275 3487
rect 6385 3519 6389 3576
rect 6385 3507 6394 3519
rect 6269 3460 6319 3464
rect 6295 3452 6299 3460
rect 6315 3452 6319 3460
rect 6231 3448 6255 3452
rect 6231 3444 6235 3448
rect 6251 3444 6255 3448
rect 6385 3424 6389 3507
rect 6431 3488 6435 3556
rect 6453 3527 6457 3576
rect 6463 3555 6467 3576
rect 6483 3564 6487 3576
rect 6491 3572 6495 3576
rect 6491 3568 6525 3572
rect 6483 3560 6513 3564
rect 6483 3559 6501 3560
rect 6463 3551 6487 3555
rect 6431 3476 6433 3488
rect 6431 3464 6435 3476
rect 6453 3469 6457 3515
rect 6295 3388 6299 3392
rect 6315 3388 6319 3392
rect 6449 3463 6457 3469
rect 6449 3434 6453 3463
rect 6481 3456 6487 3551
rect 6449 3427 6457 3434
rect 6453 3404 6457 3427
rect 6461 3404 6465 3444
rect 6481 3424 6485 3456
rect 6521 3442 6525 3568
rect 6537 3462 6541 3576
rect 6559 3564 6563 3576
rect 6561 3552 6563 3564
rect 6569 3564 6573 3576
rect 6569 3552 6571 3564
rect 6489 3430 6513 3432
rect 6489 3428 6525 3430
rect 6489 3424 6493 3428
rect 6535 3424 6539 3450
rect 6553 3442 6557 3552
rect 6591 3544 6595 3576
rect 6562 3540 6595 3544
rect 6562 3476 6566 3540
rect 6582 3491 6586 3520
rect 6601 3518 6605 3576
rect 6621 3519 6625 3556
rect 6582 3483 6591 3491
rect 6562 3464 6565 3476
rect 6555 3424 6559 3430
rect 6567 3424 6571 3464
rect 6587 3424 6591 3483
rect 6601 3424 6605 3506
rect 6621 3464 6625 3507
rect 43 3380 47 3384
rect 65 3380 69 3384
rect 111 3380 115 3384
rect 133 3380 137 3384
rect 141 3380 145 3384
rect 161 3380 165 3384
rect 169 3380 173 3384
rect 215 3380 219 3384
rect 235 3380 239 3384
rect 247 3380 251 3384
rect 267 3380 271 3384
rect 281 3380 285 3384
rect 301 3380 305 3384
rect 351 3380 355 3384
rect 371 3380 375 3384
rect 431 3380 435 3384
rect 453 3380 457 3384
rect 525 3380 529 3384
rect 545 3380 549 3384
rect 565 3380 569 3384
rect 625 3380 629 3384
rect 645 3380 649 3384
rect 703 3380 707 3384
rect 725 3380 729 3384
rect 771 3380 775 3384
rect 793 3380 797 3384
rect 851 3380 855 3384
rect 871 3380 875 3384
rect 943 3380 947 3384
rect 965 3380 969 3384
rect 1025 3380 1029 3384
rect 1083 3380 1087 3384
rect 1105 3380 1109 3384
rect 1163 3380 1167 3384
rect 1185 3380 1189 3384
rect 1231 3380 1235 3384
rect 1253 3380 1257 3384
rect 1261 3380 1265 3384
rect 1281 3380 1285 3384
rect 1289 3380 1293 3384
rect 1335 3380 1339 3384
rect 1355 3380 1359 3384
rect 1367 3380 1371 3384
rect 1387 3380 1391 3384
rect 1401 3380 1405 3384
rect 1421 3380 1425 3384
rect 1497 3380 1501 3384
rect 1505 3380 1509 3384
rect 1551 3380 1555 3384
rect 1573 3380 1577 3384
rect 1581 3380 1585 3384
rect 1601 3380 1605 3384
rect 1609 3380 1613 3384
rect 1655 3380 1659 3384
rect 1675 3380 1679 3384
rect 1687 3380 1691 3384
rect 1707 3380 1711 3384
rect 1721 3380 1725 3384
rect 1741 3380 1745 3384
rect 1801 3380 1805 3384
rect 1823 3380 1827 3384
rect 1845 3380 1849 3384
rect 1905 3380 1909 3384
rect 1970 3380 1974 3384
rect 1992 3380 1996 3384
rect 2000 3380 2004 3384
rect 2051 3380 2055 3384
rect 2059 3380 2063 3384
rect 2145 3380 2149 3384
rect 2201 3380 2205 3384
rect 2223 3380 2227 3384
rect 2245 3380 2249 3384
rect 2317 3380 2321 3384
rect 2325 3380 2329 3384
rect 2371 3380 2375 3384
rect 2393 3380 2397 3384
rect 2401 3380 2405 3384
rect 2421 3380 2425 3384
rect 2429 3380 2433 3384
rect 2475 3380 2479 3384
rect 2495 3380 2499 3384
rect 2507 3380 2511 3384
rect 2527 3380 2531 3384
rect 2541 3380 2545 3384
rect 2561 3380 2565 3384
rect 2611 3380 2615 3384
rect 2619 3380 2623 3384
rect 2696 3380 2700 3384
rect 2704 3380 2708 3384
rect 2726 3380 2730 3384
rect 2805 3380 2809 3384
rect 2865 3380 2869 3384
rect 2885 3380 2889 3384
rect 2936 3380 2940 3384
rect 2944 3380 2948 3384
rect 2966 3380 2970 3384
rect 3031 3380 3035 3384
rect 3051 3380 3055 3384
rect 3071 3380 3075 3384
rect 3131 3380 3135 3384
rect 3205 3380 3209 3384
rect 3225 3380 3229 3384
rect 3245 3380 3249 3384
rect 3265 3380 3269 3384
rect 3325 3380 3329 3384
rect 3371 3380 3375 3384
rect 3393 3380 3397 3384
rect 3401 3380 3405 3384
rect 3421 3380 3425 3384
rect 3429 3380 3433 3384
rect 3475 3380 3479 3384
rect 3495 3380 3499 3384
rect 3507 3380 3511 3384
rect 3527 3380 3531 3384
rect 3541 3380 3545 3384
rect 3561 3380 3565 3384
rect 3625 3380 3629 3384
rect 3645 3380 3649 3384
rect 3665 3380 3669 3384
rect 3685 3380 3689 3384
rect 3731 3380 3735 3384
rect 3753 3380 3757 3384
rect 3761 3380 3765 3384
rect 3781 3380 3785 3384
rect 3789 3380 3793 3384
rect 3835 3380 3839 3384
rect 3855 3380 3859 3384
rect 3867 3380 3871 3384
rect 3887 3380 3891 3384
rect 3901 3380 3905 3384
rect 3921 3380 3925 3384
rect 3985 3380 3989 3384
rect 4031 3380 4035 3384
rect 4053 3380 4057 3384
rect 4061 3380 4065 3384
rect 4081 3380 4085 3384
rect 4089 3380 4093 3384
rect 4135 3380 4139 3384
rect 4155 3380 4159 3384
rect 4167 3380 4171 3384
rect 4187 3380 4191 3384
rect 4201 3380 4205 3384
rect 4221 3380 4225 3384
rect 4285 3380 4289 3384
rect 4345 3380 4349 3384
rect 4391 3380 4395 3384
rect 4411 3380 4415 3384
rect 4475 3380 4479 3384
rect 4495 3380 4499 3384
rect 4509 3380 4513 3384
rect 4529 3380 4533 3384
rect 4541 3380 4545 3384
rect 4561 3380 4565 3384
rect 4607 3380 4611 3384
rect 4615 3380 4619 3384
rect 4635 3380 4639 3384
rect 4643 3380 4647 3384
rect 4665 3380 4669 3384
rect 4725 3380 4729 3384
rect 4771 3380 4775 3384
rect 4793 3380 4797 3384
rect 4801 3380 4805 3384
rect 4821 3380 4825 3384
rect 4829 3380 4833 3384
rect 4875 3380 4879 3384
rect 4895 3380 4899 3384
rect 4907 3380 4911 3384
rect 4927 3380 4931 3384
rect 4941 3380 4945 3384
rect 4961 3380 4965 3384
rect 5025 3380 5029 3384
rect 5045 3380 5049 3384
rect 5065 3380 5069 3384
rect 5085 3380 5089 3384
rect 5145 3380 5149 3384
rect 5191 3380 5195 3384
rect 5213 3380 5217 3384
rect 5221 3380 5225 3384
rect 5241 3380 5245 3384
rect 5249 3380 5253 3384
rect 5295 3380 5299 3384
rect 5315 3380 5319 3384
rect 5327 3380 5331 3384
rect 5347 3380 5351 3384
rect 5361 3380 5365 3384
rect 5381 3380 5385 3384
rect 5431 3380 5435 3384
rect 5453 3380 5457 3384
rect 5461 3380 5465 3384
rect 5481 3380 5485 3384
rect 5489 3380 5493 3384
rect 5535 3380 5539 3384
rect 5555 3380 5559 3384
rect 5567 3380 5571 3384
rect 5587 3380 5591 3384
rect 5601 3380 5605 3384
rect 5621 3380 5625 3384
rect 5676 3380 5680 3384
rect 5684 3380 5688 3384
rect 5706 3380 5710 3384
rect 5776 3380 5780 3384
rect 5784 3380 5788 3384
rect 5806 3380 5810 3384
rect 5885 3380 5889 3384
rect 5945 3380 5949 3384
rect 5965 3380 5969 3384
rect 5985 3380 5989 3384
rect 6005 3380 6009 3384
rect 6051 3380 6055 3384
rect 6071 3380 6075 3384
rect 6145 3380 6149 3384
rect 6191 3380 6195 3384
rect 6211 3380 6215 3384
rect 6231 3380 6235 3384
rect 6251 3380 6255 3384
rect 6385 3380 6389 3384
rect 6431 3380 6435 3384
rect 6453 3380 6457 3384
rect 6461 3380 6465 3384
rect 6481 3380 6485 3384
rect 6489 3380 6493 3384
rect 6535 3380 6539 3384
rect 6555 3380 6559 3384
rect 6567 3380 6571 3384
rect 6587 3380 6591 3384
rect 6601 3380 6605 3384
rect 6621 3380 6625 3384
rect 43 3356 47 3360
rect 65 3356 69 3360
rect 111 3356 115 3360
rect 133 3356 137 3360
rect 141 3356 145 3360
rect 161 3356 165 3360
rect 169 3356 173 3360
rect 215 3356 219 3360
rect 235 3356 239 3360
rect 247 3356 251 3360
rect 267 3356 271 3360
rect 281 3356 285 3360
rect 301 3356 305 3360
rect 351 3356 355 3360
rect 371 3356 375 3360
rect 445 3356 449 3360
rect 465 3356 469 3360
rect 485 3356 489 3360
rect 545 3356 549 3360
rect 565 3356 569 3360
rect 611 3356 615 3360
rect 671 3356 675 3360
rect 691 3356 695 3360
rect 711 3356 715 3360
rect 771 3356 775 3360
rect 791 3356 795 3360
rect 870 3356 874 3360
rect 892 3356 896 3360
rect 900 3356 904 3360
rect 951 3356 955 3360
rect 1011 3356 1015 3360
rect 1019 3356 1023 3360
rect 1096 3356 1100 3360
rect 1104 3356 1108 3360
rect 1126 3356 1130 3360
rect 1196 3356 1200 3360
rect 1204 3356 1208 3360
rect 1226 3356 1230 3360
rect 1291 3356 1295 3360
rect 1311 3356 1315 3360
rect 1371 3356 1375 3360
rect 1393 3356 1397 3360
rect 1401 3356 1405 3360
rect 1421 3356 1425 3360
rect 1429 3356 1433 3360
rect 1475 3356 1479 3360
rect 1495 3356 1499 3360
rect 1507 3356 1511 3360
rect 1527 3356 1531 3360
rect 1541 3356 1545 3360
rect 1561 3356 1565 3360
rect 1621 3356 1625 3360
rect 1643 3356 1647 3360
rect 1665 3356 1669 3360
rect 1725 3356 1729 3360
rect 1745 3356 1749 3360
rect 1765 3356 1769 3360
rect 1825 3356 1829 3360
rect 1845 3356 1849 3360
rect 1865 3356 1869 3360
rect 1911 3356 1915 3360
rect 1931 3356 1935 3360
rect 1951 3356 1955 3360
rect 2015 3356 2019 3360
rect 2035 3356 2039 3360
rect 2049 3356 2053 3360
rect 2069 3356 2073 3360
rect 2081 3356 2085 3360
rect 2101 3356 2105 3360
rect 2147 3356 2151 3360
rect 2155 3356 2159 3360
rect 2175 3356 2179 3360
rect 2183 3356 2187 3360
rect 2205 3356 2209 3360
rect 2251 3356 2255 3360
rect 2271 3356 2275 3360
rect 2331 3356 2335 3360
rect 2339 3356 2343 3360
rect 2437 3356 2441 3360
rect 2445 3356 2449 3360
rect 2510 3356 2514 3360
rect 2532 3356 2536 3360
rect 2540 3356 2544 3360
rect 2591 3356 2595 3360
rect 2655 3356 2659 3360
rect 2675 3356 2679 3360
rect 2689 3356 2693 3360
rect 2709 3356 2713 3360
rect 2721 3356 2725 3360
rect 2741 3356 2745 3360
rect 2787 3356 2791 3360
rect 2795 3356 2799 3360
rect 2815 3356 2819 3360
rect 2823 3356 2827 3360
rect 2845 3356 2849 3360
rect 2891 3356 2895 3360
rect 2911 3356 2915 3360
rect 2985 3356 2989 3360
rect 3005 3356 3009 3360
rect 3070 3356 3074 3360
rect 3092 3356 3096 3360
rect 3100 3356 3104 3360
rect 3165 3356 3169 3360
rect 3185 3356 3189 3360
rect 3245 3356 3249 3360
rect 3310 3356 3314 3360
rect 3332 3356 3336 3360
rect 3340 3356 3344 3360
rect 3391 3356 3395 3360
rect 3477 3356 3481 3360
rect 3485 3356 3489 3360
rect 3545 3356 3549 3360
rect 3565 3356 3569 3360
rect 3585 3356 3589 3360
rect 3657 3356 3661 3360
rect 3665 3356 3669 3360
rect 3711 3356 3715 3360
rect 3733 3356 3737 3360
rect 3741 3356 3745 3360
rect 3761 3356 3765 3360
rect 3769 3356 3773 3360
rect 3815 3356 3819 3360
rect 3835 3356 3839 3360
rect 3847 3356 3851 3360
rect 3867 3356 3871 3360
rect 3881 3356 3885 3360
rect 3901 3356 3905 3360
rect 3951 3356 3955 3360
rect 3971 3356 3975 3360
rect 3991 3356 3995 3360
rect 4011 3356 4015 3360
rect 4085 3356 4089 3360
rect 4105 3356 4109 3360
rect 4125 3356 4129 3360
rect 4145 3356 4149 3360
rect 4195 3356 4199 3360
rect 4215 3356 4219 3360
rect 4229 3356 4233 3360
rect 4249 3356 4253 3360
rect 4261 3356 4265 3360
rect 4281 3356 4285 3360
rect 4327 3356 4331 3360
rect 4335 3356 4339 3360
rect 4355 3356 4359 3360
rect 4363 3356 4367 3360
rect 4385 3356 4389 3360
rect 4431 3356 4435 3360
rect 4439 3356 4443 3360
rect 4511 3356 4515 3360
rect 4531 3356 4535 3360
rect 4551 3356 4555 3360
rect 4571 3356 4575 3360
rect 4631 3356 4635 3360
rect 4639 3356 4643 3360
rect 4711 3356 4715 3360
rect 4719 3356 4723 3360
rect 4791 3356 4795 3360
rect 4851 3356 4855 3360
rect 4871 3356 4875 3360
rect 4891 3356 4895 3360
rect 4911 3356 4915 3360
rect 4971 3356 4975 3360
rect 4991 3356 4995 3360
rect 5011 3356 5015 3360
rect 5071 3356 5075 3360
rect 5093 3356 5097 3360
rect 5101 3356 5105 3360
rect 5121 3356 5125 3360
rect 5129 3356 5133 3360
rect 5175 3356 5179 3360
rect 5195 3356 5199 3360
rect 5207 3356 5211 3360
rect 5227 3356 5231 3360
rect 5241 3356 5245 3360
rect 5261 3356 5265 3360
rect 5325 3356 5329 3360
rect 5371 3356 5405 3360
rect 5421 3356 5425 3360
rect 5431 3356 5435 3360
rect 5505 3356 5509 3360
rect 5555 3356 5559 3360
rect 5575 3356 5579 3360
rect 5589 3356 5593 3360
rect 5609 3356 5613 3360
rect 5621 3356 5625 3360
rect 5641 3356 5645 3360
rect 5687 3356 5691 3360
rect 5695 3356 5699 3360
rect 5715 3356 5719 3360
rect 5723 3356 5727 3360
rect 5745 3356 5749 3360
rect 5810 3356 5814 3360
rect 5832 3356 5836 3360
rect 5840 3356 5844 3360
rect 5905 3356 5909 3360
rect 5965 3356 5969 3360
rect 5985 3356 5989 3360
rect 6005 3356 6009 3360
rect 6056 3356 6060 3360
rect 6064 3356 6068 3360
rect 6086 3356 6090 3360
rect 6165 3356 6169 3360
rect 6185 3356 6189 3360
rect 6245 3356 6249 3360
rect 6265 3356 6269 3360
rect 6285 3356 6289 3360
rect 6345 3356 6349 3360
rect 6365 3356 6369 3360
rect 6416 3356 6420 3360
rect 6424 3356 6428 3360
rect 6446 3356 6450 3360
rect 6511 3356 6515 3360
rect 6533 3356 6537 3360
rect 6541 3356 6545 3360
rect 6561 3356 6565 3360
rect 6569 3356 6573 3360
rect 6615 3356 6619 3360
rect 6635 3356 6639 3360
rect 6647 3356 6651 3360
rect 6667 3356 6671 3360
rect 6681 3356 6685 3360
rect 6701 3356 6705 3360
rect 43 3270 47 3276
rect 43 3258 45 3270
rect 65 3253 69 3316
rect 133 3313 137 3336
rect 129 3306 137 3313
rect 129 3277 133 3306
rect 141 3296 145 3336
rect 161 3284 165 3316
rect 169 3312 173 3316
rect 169 3310 205 3312
rect 169 3308 193 3310
rect 111 3264 115 3276
rect 129 3271 137 3277
rect 65 3241 74 3253
rect 111 3252 113 3264
rect 43 3190 45 3202
rect 43 3184 47 3190
rect 65 3164 69 3241
rect 111 3184 115 3252
rect 133 3225 137 3271
rect 133 3164 137 3213
rect 161 3189 167 3284
rect 143 3185 167 3189
rect 143 3164 147 3185
rect 163 3180 181 3181
rect 163 3176 193 3180
rect 163 3164 167 3176
rect 201 3172 205 3298
rect 215 3290 219 3316
rect 235 3310 239 3316
rect 171 3168 205 3172
rect 171 3164 175 3168
rect 217 3164 221 3278
rect 233 3188 237 3298
rect 247 3276 251 3316
rect 242 3264 245 3276
rect 242 3200 246 3264
rect 267 3257 271 3316
rect 262 3249 271 3257
rect 262 3220 266 3249
rect 281 3234 285 3316
rect 301 3233 305 3276
rect 351 3239 355 3316
rect 242 3196 275 3200
rect 241 3176 243 3188
rect 239 3164 243 3176
rect 249 3176 251 3188
rect 249 3164 253 3176
rect 271 3164 275 3196
rect 281 3164 285 3222
rect 346 3227 355 3239
rect 301 3184 305 3221
rect 349 3211 355 3227
rect 371 3239 375 3316
rect 371 3227 374 3239
rect 371 3211 377 3227
rect 349 3204 357 3211
rect 353 3184 357 3204
rect 363 3204 377 3211
rect 445 3219 449 3276
rect 465 3262 469 3276
rect 485 3262 489 3276
rect 465 3256 480 3262
rect 485 3256 501 3262
rect 474 3233 480 3256
rect 445 3207 454 3219
rect 363 3184 367 3204
rect 452 3164 456 3207
rect 474 3184 478 3221
rect 494 3219 501 3256
rect 545 3239 549 3316
rect 546 3227 549 3239
rect 543 3211 549 3227
rect 565 3239 569 3316
rect 565 3227 574 3239
rect 611 3233 615 3316
rect 671 3308 675 3316
rect 660 3304 675 3308
rect 691 3304 695 3316
rect 660 3273 666 3304
rect 680 3300 695 3304
rect 680 3293 686 3300
rect 666 3261 676 3273
rect 565 3211 571 3227
rect 606 3221 615 3233
rect 494 3194 501 3207
rect 543 3204 557 3211
rect 482 3188 501 3194
rect 482 3184 486 3188
rect 553 3184 557 3204
rect 563 3204 571 3211
rect 563 3184 567 3204
rect 611 3164 615 3221
rect 672 3204 676 3261
rect 680 3204 684 3281
rect 711 3273 715 3316
rect 688 3261 695 3273
rect 707 3261 715 3273
rect 688 3204 692 3261
rect 771 3239 775 3316
rect 766 3227 775 3239
rect 769 3211 775 3227
rect 791 3239 795 3316
rect 870 3273 874 3316
rect 867 3261 874 3273
rect 791 3227 794 3239
rect 791 3211 797 3227
rect 769 3204 777 3211
rect 773 3184 777 3204
rect 783 3204 797 3211
rect 783 3184 787 3204
rect 865 3184 869 3261
rect 892 3219 896 3276
rect 900 3272 904 3276
rect 900 3264 918 3272
rect 914 3253 918 3264
rect 885 3207 894 3219
rect 885 3184 889 3207
rect 914 3196 918 3241
rect 951 3233 955 3316
rect 1011 3253 1015 3276
rect 1006 3241 1015 3253
rect 1019 3253 1023 3276
rect 1096 3272 1100 3276
rect 1082 3264 1100 3272
rect 1082 3253 1086 3264
rect 1019 3241 1034 3253
rect 946 3221 955 3233
rect 905 3189 918 3196
rect 905 3184 909 3189
rect 951 3164 955 3221
rect 1011 3164 1015 3241
rect 1031 3164 1035 3241
rect 1082 3196 1086 3241
rect 1104 3219 1108 3276
rect 1126 3273 1130 3316
rect 1126 3261 1133 3273
rect 1196 3272 1200 3276
rect 1182 3264 1200 3272
rect 1106 3207 1115 3219
rect 1082 3189 1095 3196
rect 1091 3184 1095 3189
rect 1111 3184 1115 3207
rect 1131 3184 1135 3261
rect 1182 3253 1186 3264
rect 1182 3196 1186 3241
rect 1204 3219 1208 3276
rect 1226 3273 1230 3316
rect 1226 3261 1233 3273
rect 1206 3207 1215 3219
rect 1182 3189 1195 3196
rect 1191 3184 1195 3189
rect 1211 3184 1215 3207
rect 1231 3184 1235 3261
rect 1291 3239 1295 3316
rect 1286 3227 1295 3239
rect 1289 3211 1295 3227
rect 1311 3239 1315 3316
rect 1393 3313 1397 3336
rect 1389 3306 1397 3313
rect 1389 3277 1393 3306
rect 1401 3296 1405 3336
rect 1421 3284 1425 3316
rect 1429 3312 1433 3316
rect 1429 3310 1465 3312
rect 1429 3308 1453 3310
rect 1371 3264 1375 3276
rect 1389 3271 1397 3277
rect 1371 3252 1373 3264
rect 1311 3227 1314 3239
rect 1311 3211 1317 3227
rect 1289 3204 1297 3211
rect 1293 3184 1297 3204
rect 1303 3204 1317 3211
rect 1303 3184 1307 3204
rect 1371 3184 1375 3252
rect 1393 3225 1397 3271
rect 1393 3164 1397 3213
rect 1421 3189 1427 3284
rect 1403 3185 1427 3189
rect 1403 3164 1407 3185
rect 1423 3180 1441 3181
rect 1423 3176 1453 3180
rect 1423 3164 1427 3176
rect 1461 3172 1465 3298
rect 1475 3290 1479 3316
rect 1495 3310 1499 3316
rect 1431 3168 1465 3172
rect 1431 3164 1435 3168
rect 1477 3164 1481 3278
rect 1493 3188 1497 3298
rect 1507 3276 1511 3316
rect 1502 3264 1505 3276
rect 1502 3200 1506 3264
rect 1527 3257 1531 3316
rect 1522 3249 1531 3257
rect 1522 3220 1526 3249
rect 1541 3234 1545 3316
rect 1561 3233 1565 3276
rect 1502 3196 1535 3200
rect 1501 3176 1503 3188
rect 1499 3164 1503 3176
rect 1509 3176 1511 3188
rect 1509 3164 1513 3176
rect 1531 3164 1535 3196
rect 1541 3164 1545 3222
rect 1561 3184 1565 3221
rect 1621 3202 1625 3276
rect 1643 3239 1647 3316
rect 1665 3253 1669 3316
rect 1665 3241 1674 3253
rect 1646 3227 1659 3239
rect 1621 3190 1633 3202
rect 1635 3184 1639 3190
rect 1655 3184 1659 3227
rect 1665 3184 1669 3241
rect 1725 3219 1729 3276
rect 1745 3262 1749 3276
rect 1765 3262 1769 3276
rect 1825 3273 1829 3316
rect 1845 3304 1849 3316
rect 1865 3308 1869 3316
rect 1865 3304 1880 3308
rect 1845 3300 1860 3304
rect 1854 3293 1860 3300
rect 1745 3256 1760 3262
rect 1765 3256 1781 3262
rect 1825 3261 1833 3273
rect 1845 3261 1852 3273
rect 1754 3233 1760 3256
rect 1725 3207 1734 3219
rect 1732 3164 1736 3207
rect 1754 3184 1758 3221
rect 1774 3219 1781 3256
rect 1774 3194 1781 3207
rect 1848 3204 1852 3261
rect 1856 3204 1860 3281
rect 1874 3273 1880 3304
rect 1864 3261 1874 3273
rect 1911 3262 1915 3276
rect 1931 3262 1935 3276
rect 1864 3204 1868 3261
rect 1899 3256 1915 3262
rect 1920 3256 1935 3262
rect 1899 3219 1906 3256
rect 1920 3233 1926 3256
rect 1762 3188 1781 3194
rect 1762 3184 1766 3188
rect 1899 3194 1906 3207
rect 1899 3188 1918 3194
rect 1914 3184 1918 3188
rect 1922 3184 1926 3221
rect 1951 3219 1955 3276
rect 2015 3233 2019 3276
rect 2035 3234 2039 3316
rect 2049 3257 2053 3316
rect 2069 3276 2073 3316
rect 2081 3310 2085 3316
rect 2075 3264 2078 3276
rect 2049 3249 2058 3257
rect 1946 3207 1955 3219
rect 1944 3164 1948 3207
rect 2015 3184 2019 3221
rect 2035 3164 2039 3222
rect 2054 3220 2058 3249
rect 2074 3200 2078 3264
rect 2045 3196 2078 3200
rect 2045 3164 2049 3196
rect 2083 3188 2087 3298
rect 2101 3290 2105 3316
rect 2147 3312 2151 3316
rect 2115 3310 2151 3312
rect 2127 3308 2151 3310
rect 2069 3176 2071 3188
rect 2067 3164 2071 3176
rect 2077 3176 2079 3188
rect 2077 3164 2081 3176
rect 2099 3164 2103 3278
rect 2115 3172 2119 3298
rect 2155 3284 2159 3316
rect 2175 3296 2179 3336
rect 2183 3313 2187 3336
rect 2183 3306 2191 3313
rect 2153 3189 2159 3284
rect 2187 3277 2191 3306
rect 2183 3271 2191 3277
rect 2183 3225 2187 3271
rect 2205 3264 2209 3276
rect 2207 3252 2209 3264
rect 2153 3185 2177 3189
rect 2139 3180 2157 3181
rect 2127 3176 2157 3180
rect 2115 3168 2149 3172
rect 2145 3164 2149 3168
rect 2153 3164 2157 3176
rect 2173 3164 2177 3185
rect 2183 3164 2187 3213
rect 2205 3184 2209 3252
rect 2251 3239 2255 3316
rect 2246 3227 2255 3239
rect 2249 3211 2255 3227
rect 2271 3239 2275 3316
rect 2331 3253 2335 3276
rect 2326 3241 2335 3253
rect 2339 3253 2343 3276
rect 2437 3253 2441 3276
rect 2339 3241 2354 3253
rect 2426 3241 2441 3253
rect 2445 3253 2449 3276
rect 2510 3273 2514 3316
rect 2507 3261 2514 3273
rect 2445 3241 2454 3253
rect 2271 3227 2274 3239
rect 2271 3211 2277 3227
rect 2249 3204 2257 3211
rect 2253 3184 2257 3204
rect 2263 3204 2277 3211
rect 2263 3184 2267 3204
rect 2331 3164 2335 3241
rect 2351 3164 2355 3241
rect 2425 3164 2429 3241
rect 2445 3164 2449 3241
rect 2505 3184 2509 3261
rect 2532 3219 2536 3276
rect 2540 3272 2544 3276
rect 2540 3264 2558 3272
rect 2554 3253 2558 3264
rect 2525 3207 2534 3219
rect 2525 3184 2529 3207
rect 2554 3196 2558 3241
rect 2591 3233 2595 3316
rect 2655 3233 2659 3276
rect 2675 3234 2679 3316
rect 2689 3257 2693 3316
rect 2709 3276 2713 3316
rect 2721 3310 2725 3316
rect 2715 3264 2718 3276
rect 2689 3249 2698 3257
rect 2586 3221 2595 3233
rect 2545 3189 2558 3196
rect 2545 3184 2549 3189
rect 2591 3164 2595 3221
rect 2655 3184 2659 3221
rect 2675 3164 2679 3222
rect 2694 3220 2698 3249
rect 2714 3200 2718 3264
rect 2685 3196 2718 3200
rect 2685 3164 2689 3196
rect 2723 3188 2727 3298
rect 2741 3290 2745 3316
rect 2787 3312 2791 3316
rect 2755 3310 2791 3312
rect 2767 3308 2791 3310
rect 2709 3176 2711 3188
rect 2707 3164 2711 3176
rect 2717 3176 2719 3188
rect 2717 3164 2721 3176
rect 2739 3164 2743 3278
rect 2755 3172 2759 3298
rect 2795 3284 2799 3316
rect 2815 3296 2819 3336
rect 2823 3313 2827 3336
rect 2823 3306 2831 3313
rect 2793 3189 2799 3284
rect 2827 3277 2831 3306
rect 2823 3271 2831 3277
rect 2823 3225 2827 3271
rect 2845 3264 2849 3276
rect 2847 3252 2849 3264
rect 2793 3185 2817 3189
rect 2779 3180 2797 3181
rect 2767 3176 2797 3180
rect 2755 3168 2789 3172
rect 2785 3164 2789 3168
rect 2793 3164 2797 3176
rect 2813 3164 2817 3185
rect 2823 3164 2827 3213
rect 2845 3184 2849 3252
rect 2891 3239 2895 3316
rect 2886 3227 2895 3239
rect 2889 3211 2895 3227
rect 2911 3239 2915 3316
rect 2985 3239 2989 3316
rect 2911 3227 2914 3239
rect 2986 3227 2989 3239
rect 2911 3211 2917 3227
rect 2889 3204 2897 3211
rect 2893 3184 2897 3204
rect 2903 3204 2917 3211
rect 2983 3211 2989 3227
rect 3005 3239 3009 3316
rect 3070 3273 3074 3316
rect 3067 3261 3074 3273
rect 3005 3227 3014 3239
rect 3005 3211 3011 3227
rect 2983 3204 2997 3211
rect 2903 3184 2907 3204
rect 2993 3184 2997 3204
rect 3003 3204 3011 3211
rect 3003 3184 3007 3204
rect 3065 3184 3069 3261
rect 3092 3219 3096 3276
rect 3100 3272 3104 3276
rect 3100 3264 3118 3272
rect 3114 3253 3118 3264
rect 3085 3207 3094 3219
rect 3085 3184 3089 3207
rect 3114 3196 3118 3241
rect 3165 3239 3169 3316
rect 3166 3227 3169 3239
rect 3163 3211 3169 3227
rect 3185 3239 3189 3316
rect 3185 3227 3194 3239
rect 3245 3233 3249 3316
rect 3310 3273 3314 3316
rect 3307 3261 3314 3273
rect 3185 3211 3191 3227
rect 3163 3204 3177 3211
rect 3105 3189 3118 3196
rect 3105 3184 3109 3189
rect 3173 3184 3177 3204
rect 3183 3204 3191 3211
rect 3245 3221 3254 3233
rect 3183 3184 3187 3204
rect 3245 3164 3249 3221
rect 3305 3184 3309 3261
rect 3332 3219 3336 3276
rect 3340 3272 3344 3276
rect 3340 3264 3358 3272
rect 3354 3253 3358 3264
rect 3325 3207 3334 3219
rect 3325 3184 3329 3207
rect 3354 3196 3358 3241
rect 3391 3233 3395 3316
rect 3733 3313 3737 3336
rect 3729 3306 3737 3313
rect 3729 3277 3733 3306
rect 3741 3296 3745 3336
rect 3761 3284 3765 3316
rect 3769 3312 3773 3316
rect 3769 3310 3805 3312
rect 3769 3308 3793 3310
rect 3477 3253 3481 3276
rect 3466 3241 3481 3253
rect 3485 3253 3489 3276
rect 3485 3241 3494 3253
rect 3386 3221 3395 3233
rect 3345 3189 3358 3196
rect 3345 3184 3349 3189
rect 3391 3164 3395 3221
rect 3465 3164 3469 3241
rect 3485 3164 3489 3241
rect 3545 3219 3549 3276
rect 3565 3262 3569 3276
rect 3585 3262 3589 3276
rect 3565 3256 3580 3262
rect 3585 3256 3601 3262
rect 3574 3233 3580 3256
rect 3545 3207 3554 3219
rect 3552 3164 3556 3207
rect 3574 3184 3578 3221
rect 3594 3219 3601 3256
rect 3657 3253 3661 3276
rect 3646 3241 3661 3253
rect 3665 3253 3669 3276
rect 3711 3264 3715 3276
rect 3729 3271 3737 3277
rect 3665 3241 3674 3253
rect 3711 3252 3713 3264
rect 3594 3194 3601 3207
rect 3582 3188 3601 3194
rect 3582 3184 3586 3188
rect 3645 3164 3649 3241
rect 3665 3164 3669 3241
rect 3711 3184 3715 3252
rect 3733 3225 3737 3271
rect 3733 3164 3737 3213
rect 3761 3189 3767 3284
rect 3743 3185 3767 3189
rect 3743 3164 3747 3185
rect 3763 3180 3781 3181
rect 3763 3176 3793 3180
rect 3763 3164 3767 3176
rect 3801 3172 3805 3298
rect 3815 3290 3819 3316
rect 3835 3310 3839 3316
rect 3771 3168 3805 3172
rect 3771 3164 3775 3168
rect 3817 3164 3821 3278
rect 3833 3188 3837 3298
rect 3847 3276 3851 3316
rect 3842 3264 3845 3276
rect 3842 3200 3846 3264
rect 3867 3257 3871 3316
rect 3862 3249 3871 3257
rect 3862 3220 3866 3249
rect 3881 3234 3885 3316
rect 3901 3233 3905 3276
rect 3951 3254 3955 3276
rect 3971 3254 3975 3276
rect 3935 3253 3955 3254
rect 3947 3248 3955 3253
rect 3962 3248 3975 3254
rect 3842 3196 3875 3200
rect 3841 3176 3843 3188
rect 3839 3164 3843 3176
rect 3849 3176 3851 3188
rect 3849 3164 3853 3176
rect 3871 3164 3875 3196
rect 3881 3164 3885 3222
rect 3901 3184 3905 3221
rect 3941 3199 3947 3241
rect 3962 3219 3966 3248
rect 3991 3219 3995 3276
rect 4011 3253 4015 3276
rect 4085 3253 4089 3276
rect 4011 3241 4014 3253
rect 4086 3241 4089 3253
rect 3991 3207 3993 3219
rect 3941 3192 3958 3199
rect 3954 3184 3958 3192
rect 3962 3184 3966 3207
rect 3991 3205 3995 3207
rect 3982 3198 3995 3205
rect 3982 3184 3986 3198
rect 4014 3193 4020 3241
rect 3990 3189 4020 3193
rect 4080 3193 4086 3241
rect 4105 3219 4109 3276
rect 4125 3254 4129 3276
rect 4145 3254 4149 3276
rect 4125 3248 4138 3254
rect 4145 3253 4165 3254
rect 4145 3248 4153 3253
rect 4134 3219 4138 3248
rect 4107 3207 4109 3219
rect 4105 3205 4109 3207
rect 4105 3198 4118 3205
rect 4080 3189 4110 3193
rect 3990 3184 3994 3189
rect 4106 3184 4110 3189
rect 4114 3184 4118 3198
rect 4134 3184 4138 3207
rect 4153 3199 4159 3241
rect 4195 3233 4199 3276
rect 4215 3234 4219 3316
rect 4229 3257 4233 3316
rect 4249 3276 4253 3316
rect 4261 3310 4265 3316
rect 4255 3264 4258 3276
rect 4229 3249 4238 3257
rect 4142 3192 4159 3199
rect 4142 3184 4146 3192
rect 4195 3184 4199 3221
rect 4215 3164 4219 3222
rect 4234 3220 4238 3249
rect 4254 3200 4258 3264
rect 4225 3196 4258 3200
rect 4225 3164 4229 3196
rect 4263 3188 4267 3298
rect 4281 3290 4285 3316
rect 4327 3312 4331 3316
rect 4295 3310 4331 3312
rect 4307 3308 4331 3310
rect 4249 3176 4251 3188
rect 4247 3164 4251 3176
rect 4257 3176 4259 3188
rect 4257 3164 4261 3176
rect 4279 3164 4283 3278
rect 4295 3172 4299 3298
rect 4335 3284 4339 3316
rect 4355 3296 4359 3336
rect 4363 3313 4367 3336
rect 4363 3306 4371 3313
rect 4333 3189 4339 3284
rect 4367 3277 4371 3306
rect 4363 3271 4371 3277
rect 4363 3225 4367 3271
rect 4385 3264 4389 3276
rect 4387 3252 4389 3264
rect 4431 3253 4435 3276
rect 4333 3185 4357 3189
rect 4319 3180 4337 3181
rect 4307 3176 4337 3180
rect 4295 3168 4329 3172
rect 4325 3164 4329 3168
rect 4333 3164 4337 3176
rect 4353 3164 4357 3185
rect 4363 3164 4367 3213
rect 4385 3184 4389 3252
rect 4426 3241 4435 3253
rect 4439 3253 4443 3276
rect 4511 3254 4515 3276
rect 4531 3254 4535 3276
rect 4495 3253 4515 3254
rect 4439 3241 4454 3253
rect 4507 3248 4515 3253
rect 4522 3248 4535 3254
rect 4431 3164 4435 3241
rect 4451 3164 4455 3241
rect 4501 3199 4507 3241
rect 4522 3219 4526 3248
rect 4551 3219 4555 3276
rect 4571 3253 4575 3276
rect 4631 3253 4635 3276
rect 4571 3241 4574 3253
rect 4626 3241 4635 3253
rect 4639 3253 4643 3276
rect 4711 3253 4715 3276
rect 4639 3241 4654 3253
rect 4706 3241 4715 3253
rect 4719 3253 4723 3276
rect 4719 3241 4734 3253
rect 4551 3207 4553 3219
rect 4501 3192 4518 3199
rect 4514 3184 4518 3192
rect 4522 3184 4526 3207
rect 4551 3205 4555 3207
rect 4542 3198 4555 3205
rect 4542 3184 4546 3198
rect 4574 3193 4580 3241
rect 4550 3189 4580 3193
rect 4550 3184 4554 3189
rect 4631 3164 4635 3241
rect 4651 3164 4655 3241
rect 4711 3164 4715 3241
rect 4731 3164 4735 3241
rect 4791 3233 4795 3316
rect 5093 3313 5097 3336
rect 5089 3306 5097 3313
rect 5089 3277 5093 3306
rect 5101 3296 5105 3336
rect 5121 3284 5125 3316
rect 5129 3312 5133 3316
rect 5129 3310 5165 3312
rect 5129 3308 5153 3310
rect 4851 3254 4855 3276
rect 4871 3254 4875 3276
rect 4835 3253 4855 3254
rect 4847 3248 4855 3253
rect 4862 3248 4875 3254
rect 4786 3221 4795 3233
rect 4791 3164 4795 3221
rect 4841 3199 4847 3241
rect 4862 3219 4866 3248
rect 4891 3219 4895 3276
rect 4911 3253 4915 3276
rect 4971 3262 4975 3276
rect 4991 3262 4995 3276
rect 4959 3256 4975 3262
rect 4980 3256 4995 3262
rect 4911 3241 4914 3253
rect 4891 3207 4893 3219
rect 4841 3192 4858 3199
rect 4854 3184 4858 3192
rect 4862 3184 4866 3207
rect 4891 3205 4895 3207
rect 4882 3198 4895 3205
rect 4882 3184 4886 3198
rect 4914 3193 4920 3241
rect 4959 3219 4966 3256
rect 4980 3233 4986 3256
rect 4890 3189 4920 3193
rect 4959 3194 4966 3207
rect 4890 3184 4894 3189
rect 4959 3188 4978 3194
rect 4974 3184 4978 3188
rect 4982 3184 4986 3221
rect 5011 3219 5015 3276
rect 5006 3207 5015 3219
rect 5071 3264 5075 3276
rect 5089 3271 5097 3277
rect 5071 3252 5073 3264
rect 5004 3164 5008 3207
rect 5071 3184 5075 3252
rect 5093 3225 5097 3271
rect 5093 3164 5097 3213
rect 5121 3189 5127 3284
rect 5103 3185 5127 3189
rect 5103 3164 5107 3185
rect 5123 3180 5141 3181
rect 5123 3176 5153 3180
rect 5123 3164 5127 3176
rect 5161 3172 5165 3298
rect 5175 3290 5179 3316
rect 5195 3310 5199 3316
rect 5131 3168 5165 3172
rect 5131 3164 5135 3168
rect 5177 3164 5181 3278
rect 5193 3188 5197 3298
rect 5207 3276 5211 3316
rect 5202 3264 5205 3276
rect 5202 3200 5206 3264
rect 5227 3257 5231 3316
rect 5222 3249 5231 3257
rect 5222 3220 5226 3249
rect 5241 3234 5245 3316
rect 5371 3348 5375 3356
rect 5391 3348 5395 3352
rect 5401 3348 5405 3356
rect 5261 3233 5265 3276
rect 5325 3233 5329 3316
rect 5371 3304 5375 3308
rect 5363 3300 5375 3304
rect 5202 3196 5235 3200
rect 5201 3176 5203 3188
rect 5199 3164 5203 3176
rect 5209 3176 5211 3188
rect 5209 3164 5213 3176
rect 5231 3164 5235 3196
rect 5241 3164 5245 3222
rect 5325 3221 5334 3233
rect 5261 3184 5265 3221
rect 5325 3164 5329 3221
rect 5363 3219 5367 3300
rect 5391 3263 5395 3268
rect 5401 3264 5405 3268
rect 5382 3259 5395 3263
rect 5382 3253 5387 3259
rect 5421 3254 5425 3276
rect 5395 3250 5425 3254
rect 5431 3253 5435 3276
rect 5363 3181 5367 3207
rect 5381 3210 5386 3241
rect 5431 3241 5434 3253
rect 5381 3204 5395 3210
rect 5391 3192 5395 3204
rect 5401 3192 5405 3238
rect 5421 3192 5425 3196
rect 5431 3192 5435 3241
rect 5505 3233 5509 3316
rect 5555 3233 5559 3276
rect 5575 3234 5579 3316
rect 5589 3257 5593 3316
rect 5609 3276 5613 3316
rect 5621 3310 5625 3316
rect 5615 3264 5618 3276
rect 5589 3249 5598 3257
rect 5505 3221 5514 3233
rect 5363 3176 5375 3181
rect 5371 3172 5375 3176
rect 5505 3164 5509 3221
rect 5555 3184 5559 3221
rect 5371 3144 5375 3152
rect 5391 3148 5395 3152
rect 5401 3148 5405 3152
rect 5421 3144 5425 3152
rect 5431 3148 5435 3152
rect 5575 3164 5579 3222
rect 5594 3220 5598 3249
rect 5614 3200 5618 3264
rect 5585 3196 5618 3200
rect 5585 3164 5589 3196
rect 5623 3188 5627 3298
rect 5641 3290 5645 3316
rect 5687 3312 5691 3316
rect 5655 3310 5691 3312
rect 5667 3308 5691 3310
rect 5609 3176 5611 3188
rect 5607 3164 5611 3176
rect 5617 3176 5619 3188
rect 5617 3164 5621 3176
rect 5639 3164 5643 3278
rect 5655 3172 5659 3298
rect 5695 3284 5699 3316
rect 5715 3296 5719 3336
rect 5723 3313 5727 3336
rect 5723 3306 5731 3313
rect 5693 3189 5699 3284
rect 5727 3277 5731 3306
rect 5723 3271 5731 3277
rect 5723 3225 5727 3271
rect 5745 3264 5749 3276
rect 5810 3273 5814 3316
rect 5747 3252 5749 3264
rect 5807 3261 5814 3273
rect 5693 3185 5717 3189
rect 5679 3180 5697 3181
rect 5667 3176 5697 3180
rect 5655 3168 5689 3172
rect 5685 3164 5689 3168
rect 5693 3164 5697 3176
rect 5713 3164 5717 3185
rect 5723 3164 5727 3213
rect 5745 3184 5749 3252
rect 5805 3184 5809 3261
rect 5832 3219 5836 3276
rect 5840 3272 5844 3276
rect 5840 3264 5858 3272
rect 5854 3253 5858 3264
rect 5825 3207 5834 3219
rect 5825 3184 5829 3207
rect 5854 3196 5858 3241
rect 5845 3189 5858 3196
rect 5905 3233 5909 3316
rect 5905 3221 5914 3233
rect 5845 3184 5849 3189
rect 5905 3164 5909 3221
rect 5965 3219 5969 3276
rect 5985 3262 5989 3276
rect 6005 3262 6009 3276
rect 6056 3272 6060 3276
rect 6042 3264 6060 3272
rect 5985 3256 6000 3262
rect 6005 3256 6021 3262
rect 5994 3233 6000 3256
rect 5965 3207 5974 3219
rect 5972 3164 5976 3207
rect 5994 3184 5998 3221
rect 6014 3219 6021 3256
rect 6042 3253 6046 3264
rect 6014 3194 6021 3207
rect 6002 3188 6021 3194
rect 6042 3196 6046 3241
rect 6064 3219 6068 3276
rect 6086 3273 6090 3316
rect 6086 3261 6093 3273
rect 6066 3207 6075 3219
rect 6042 3189 6055 3196
rect 6002 3184 6006 3188
rect 6051 3184 6055 3189
rect 6071 3184 6075 3207
rect 6091 3184 6095 3261
rect 6165 3239 6169 3316
rect 6166 3227 6169 3239
rect 6163 3211 6169 3227
rect 6185 3239 6189 3316
rect 6185 3227 6194 3239
rect 6185 3211 6191 3227
rect 6163 3204 6177 3211
rect 6173 3184 6177 3204
rect 6183 3204 6191 3211
rect 6245 3219 6249 3276
rect 6265 3262 6269 3276
rect 6285 3262 6289 3276
rect 6265 3256 6280 3262
rect 6285 3256 6301 3262
rect 6274 3233 6280 3256
rect 6245 3207 6254 3219
rect 6183 3184 6187 3204
rect 6252 3164 6256 3207
rect 6274 3184 6278 3221
rect 6294 3219 6301 3256
rect 6345 3239 6349 3316
rect 6346 3227 6349 3239
rect 6343 3211 6349 3227
rect 6365 3239 6369 3316
rect 6416 3272 6420 3276
rect 6402 3264 6420 3272
rect 6402 3253 6406 3264
rect 6365 3227 6374 3239
rect 6365 3211 6371 3227
rect 6294 3194 6301 3207
rect 6343 3204 6357 3211
rect 6282 3188 6301 3194
rect 6282 3184 6286 3188
rect 6353 3184 6357 3204
rect 6363 3204 6371 3211
rect 6363 3184 6367 3204
rect 6402 3196 6406 3241
rect 6424 3219 6428 3276
rect 6446 3273 6450 3316
rect 6533 3313 6537 3336
rect 6529 3306 6537 3313
rect 6529 3277 6533 3306
rect 6541 3296 6545 3336
rect 6561 3284 6565 3316
rect 6569 3312 6573 3316
rect 6569 3310 6605 3312
rect 6569 3308 6593 3310
rect 6446 3261 6453 3273
rect 6511 3264 6515 3276
rect 6529 3271 6537 3277
rect 6426 3207 6435 3219
rect 6402 3189 6415 3196
rect 6411 3184 6415 3189
rect 6431 3184 6435 3207
rect 6451 3184 6455 3261
rect 6511 3252 6513 3264
rect 6511 3184 6515 3252
rect 6533 3225 6537 3271
rect 6533 3164 6537 3213
rect 6561 3189 6567 3284
rect 6543 3185 6567 3189
rect 6543 3164 6547 3185
rect 6563 3180 6581 3181
rect 6563 3176 6593 3180
rect 6563 3164 6567 3176
rect 6601 3172 6605 3298
rect 6615 3290 6619 3316
rect 6635 3310 6639 3316
rect 6571 3168 6605 3172
rect 6571 3164 6575 3168
rect 6617 3164 6621 3278
rect 6633 3188 6637 3298
rect 6647 3276 6651 3316
rect 6642 3264 6645 3276
rect 6642 3200 6646 3264
rect 6667 3257 6671 3316
rect 6662 3249 6671 3257
rect 6662 3220 6666 3249
rect 6681 3234 6685 3316
rect 6701 3233 6705 3276
rect 6642 3196 6675 3200
rect 6641 3176 6643 3188
rect 6639 3164 6643 3176
rect 6649 3176 6651 3188
rect 6649 3164 6653 3176
rect 6671 3164 6675 3196
rect 6681 3164 6685 3222
rect 6701 3184 6705 3221
rect 43 3140 47 3144
rect 65 3140 69 3144
rect 111 3140 115 3144
rect 133 3140 137 3144
rect 143 3140 147 3144
rect 163 3140 167 3144
rect 171 3140 175 3144
rect 217 3140 221 3144
rect 239 3140 243 3144
rect 249 3140 253 3144
rect 271 3140 275 3144
rect 281 3140 285 3144
rect 301 3140 305 3144
rect 353 3140 357 3144
rect 363 3140 367 3144
rect 452 3140 456 3144
rect 474 3140 478 3144
rect 482 3140 486 3144
rect 553 3140 557 3144
rect 563 3140 567 3144
rect 611 3140 615 3144
rect 672 3140 676 3144
rect 680 3140 684 3144
rect 688 3140 692 3144
rect 773 3140 777 3144
rect 783 3140 787 3144
rect 865 3140 869 3144
rect 885 3140 889 3144
rect 905 3140 909 3144
rect 951 3140 955 3144
rect 1011 3140 1015 3144
rect 1031 3140 1035 3144
rect 1091 3140 1095 3144
rect 1111 3140 1115 3144
rect 1131 3140 1135 3144
rect 1191 3140 1195 3144
rect 1211 3140 1215 3144
rect 1231 3140 1235 3144
rect 1293 3140 1297 3144
rect 1303 3140 1307 3144
rect 1371 3140 1375 3144
rect 1393 3140 1397 3144
rect 1403 3140 1407 3144
rect 1423 3140 1427 3144
rect 1431 3140 1435 3144
rect 1477 3140 1481 3144
rect 1499 3140 1503 3144
rect 1509 3140 1513 3144
rect 1531 3140 1535 3144
rect 1541 3140 1545 3144
rect 1561 3140 1565 3144
rect 1635 3140 1639 3144
rect 1655 3140 1659 3144
rect 1665 3140 1669 3144
rect 1732 3140 1736 3144
rect 1754 3140 1758 3144
rect 1762 3140 1766 3144
rect 1848 3140 1852 3144
rect 1856 3140 1860 3144
rect 1864 3140 1868 3144
rect 1914 3140 1918 3144
rect 1922 3140 1926 3144
rect 1944 3140 1948 3144
rect 2015 3140 2019 3144
rect 2035 3140 2039 3144
rect 2045 3140 2049 3144
rect 2067 3140 2071 3144
rect 2077 3140 2081 3144
rect 2099 3140 2103 3144
rect 2145 3140 2149 3144
rect 2153 3140 2157 3144
rect 2173 3140 2177 3144
rect 2183 3140 2187 3144
rect 2205 3140 2209 3144
rect 2253 3140 2257 3144
rect 2263 3140 2267 3144
rect 2331 3140 2335 3144
rect 2351 3140 2355 3144
rect 2425 3140 2429 3144
rect 2445 3140 2449 3144
rect 2505 3140 2509 3144
rect 2525 3140 2529 3144
rect 2545 3140 2549 3144
rect 2591 3140 2595 3144
rect 2655 3140 2659 3144
rect 2675 3140 2679 3144
rect 2685 3140 2689 3144
rect 2707 3140 2711 3144
rect 2717 3140 2721 3144
rect 2739 3140 2743 3144
rect 2785 3140 2789 3144
rect 2793 3140 2797 3144
rect 2813 3140 2817 3144
rect 2823 3140 2827 3144
rect 2845 3140 2849 3144
rect 2893 3140 2897 3144
rect 2903 3140 2907 3144
rect 2993 3140 2997 3144
rect 3003 3140 3007 3144
rect 3065 3140 3069 3144
rect 3085 3140 3089 3144
rect 3105 3140 3109 3144
rect 3173 3140 3177 3144
rect 3183 3140 3187 3144
rect 3245 3140 3249 3144
rect 3305 3140 3309 3144
rect 3325 3140 3329 3144
rect 3345 3140 3349 3144
rect 3391 3140 3395 3144
rect 3465 3140 3469 3144
rect 3485 3140 3489 3144
rect 3552 3140 3556 3144
rect 3574 3140 3578 3144
rect 3582 3140 3586 3144
rect 3645 3140 3649 3144
rect 3665 3140 3669 3144
rect 3711 3140 3715 3144
rect 3733 3140 3737 3144
rect 3743 3140 3747 3144
rect 3763 3140 3767 3144
rect 3771 3140 3775 3144
rect 3817 3140 3821 3144
rect 3839 3140 3843 3144
rect 3849 3140 3853 3144
rect 3871 3140 3875 3144
rect 3881 3140 3885 3144
rect 3901 3140 3905 3144
rect 3954 3140 3958 3144
rect 3962 3140 3966 3144
rect 3982 3140 3986 3144
rect 3990 3140 3994 3144
rect 4106 3140 4110 3144
rect 4114 3140 4118 3144
rect 4134 3140 4138 3144
rect 4142 3140 4146 3144
rect 4195 3140 4199 3144
rect 4215 3140 4219 3144
rect 4225 3140 4229 3144
rect 4247 3140 4251 3144
rect 4257 3140 4261 3144
rect 4279 3140 4283 3144
rect 4325 3140 4329 3144
rect 4333 3140 4337 3144
rect 4353 3140 4357 3144
rect 4363 3140 4367 3144
rect 4385 3140 4389 3144
rect 4431 3140 4435 3144
rect 4451 3140 4455 3144
rect 4514 3140 4518 3144
rect 4522 3140 4526 3144
rect 4542 3140 4546 3144
rect 4550 3140 4554 3144
rect 4631 3140 4635 3144
rect 4651 3140 4655 3144
rect 4711 3140 4715 3144
rect 4731 3140 4735 3144
rect 4791 3140 4795 3144
rect 4854 3140 4858 3144
rect 4862 3140 4866 3144
rect 4882 3140 4886 3144
rect 4890 3140 4894 3144
rect 4974 3140 4978 3144
rect 4982 3140 4986 3144
rect 5004 3140 5008 3144
rect 5071 3140 5075 3144
rect 5093 3140 5097 3144
rect 5103 3140 5107 3144
rect 5123 3140 5127 3144
rect 5131 3140 5135 3144
rect 5177 3140 5181 3144
rect 5199 3140 5203 3144
rect 5209 3140 5213 3144
rect 5231 3140 5235 3144
rect 5241 3140 5245 3144
rect 5261 3140 5265 3144
rect 5325 3140 5329 3144
rect 5371 3140 5425 3144
rect 5505 3140 5509 3144
rect 5555 3140 5559 3144
rect 5575 3140 5579 3144
rect 5585 3140 5589 3144
rect 5607 3140 5611 3144
rect 5617 3140 5621 3144
rect 5639 3140 5643 3144
rect 5685 3140 5689 3144
rect 5693 3140 5697 3144
rect 5713 3140 5717 3144
rect 5723 3140 5727 3144
rect 5745 3140 5749 3144
rect 5805 3140 5809 3144
rect 5825 3140 5829 3144
rect 5845 3140 5849 3144
rect 5905 3140 5909 3144
rect 5972 3140 5976 3144
rect 5994 3140 5998 3144
rect 6002 3140 6006 3144
rect 6051 3140 6055 3144
rect 6071 3140 6075 3144
rect 6091 3140 6095 3144
rect 6173 3140 6177 3144
rect 6183 3140 6187 3144
rect 6252 3140 6256 3144
rect 6274 3140 6278 3144
rect 6282 3140 6286 3144
rect 6353 3140 6357 3144
rect 6363 3140 6367 3144
rect 6411 3140 6415 3144
rect 6431 3140 6435 3144
rect 6451 3140 6455 3144
rect 6511 3140 6515 3144
rect 6533 3140 6537 3144
rect 6543 3140 6547 3144
rect 6563 3140 6567 3144
rect 6571 3140 6575 3144
rect 6617 3140 6621 3144
rect 6639 3140 6643 3144
rect 6649 3140 6653 3144
rect 6671 3140 6675 3144
rect 6681 3140 6685 3144
rect 6701 3140 6705 3144
rect 31 3116 35 3120
rect 51 3116 55 3120
rect 71 3116 75 3120
rect 91 3116 95 3120
rect 111 3116 115 3120
rect 131 3116 135 3120
rect 151 3116 155 3120
rect 171 3116 175 3120
rect 243 3116 247 3120
rect 265 3116 269 3120
rect 315 3116 319 3120
rect 335 3116 339 3120
rect 345 3116 349 3120
rect 367 3116 371 3120
rect 377 3116 381 3120
rect 399 3116 403 3120
rect 445 3116 449 3120
rect 453 3116 457 3120
rect 473 3116 477 3120
rect 483 3116 487 3120
rect 505 3116 509 3120
rect 573 3116 577 3120
rect 583 3116 587 3120
rect 633 3116 637 3120
rect 643 3116 647 3120
rect 725 3116 729 3120
rect 745 3116 749 3120
rect 765 3116 769 3120
rect 833 3116 837 3120
rect 843 3116 847 3120
rect 913 3116 917 3120
rect 923 3116 927 3120
rect 974 3116 978 3120
rect 982 3116 986 3120
rect 1004 3116 1008 3120
rect 1071 3116 1075 3120
rect 1093 3116 1097 3120
rect 1103 3116 1107 3120
rect 1123 3116 1127 3120
rect 1131 3116 1135 3120
rect 1177 3116 1181 3120
rect 1199 3116 1203 3120
rect 1209 3116 1213 3120
rect 1231 3116 1235 3120
rect 1241 3116 1245 3120
rect 1261 3116 1265 3120
rect 1333 3116 1337 3120
rect 1343 3116 1347 3120
rect 1391 3116 1395 3120
rect 1413 3116 1417 3120
rect 1423 3116 1427 3120
rect 1443 3116 1447 3120
rect 1451 3116 1455 3120
rect 1497 3116 1501 3120
rect 1519 3116 1523 3120
rect 1529 3116 1533 3120
rect 1551 3116 1555 3120
rect 1561 3116 1565 3120
rect 1581 3116 1585 3120
rect 1645 3116 1649 3120
rect 1705 3116 1709 3120
rect 1725 3116 1729 3120
rect 1745 3116 1749 3120
rect 1805 3116 1809 3120
rect 1825 3116 1829 3120
rect 1895 3116 1899 3120
rect 1915 3116 1919 3120
rect 1925 3116 1929 3120
rect 1971 3116 1975 3120
rect 1991 3116 1995 3120
rect 2011 3116 2015 3120
rect 2092 3116 2096 3120
rect 2114 3116 2118 3120
rect 2122 3116 2126 3120
rect 2173 3116 2177 3120
rect 2183 3116 2187 3120
rect 2265 3116 2269 3120
rect 2311 3116 2315 3120
rect 2321 3116 2325 3120
rect 2341 3116 2345 3120
rect 2415 3116 2419 3120
rect 2435 3116 2439 3120
rect 2445 3116 2449 3120
rect 2467 3116 2471 3120
rect 2477 3116 2481 3120
rect 2499 3116 2503 3120
rect 2545 3116 2549 3120
rect 2553 3116 2557 3120
rect 2573 3116 2577 3120
rect 2583 3116 2587 3120
rect 2605 3116 2609 3120
rect 2651 3116 2655 3120
rect 2711 3116 2715 3120
rect 2731 3116 2735 3120
rect 2805 3116 2809 3120
rect 2865 3116 2869 3120
rect 2885 3116 2889 3120
rect 2905 3116 2909 3120
rect 2951 3116 2955 3120
rect 3048 3116 3052 3120
rect 3056 3116 3060 3120
rect 3064 3116 3068 3120
rect 3133 3116 3137 3120
rect 3143 3116 3147 3120
rect 3205 3116 3209 3120
rect 3225 3116 3229 3120
rect 3245 3116 3249 3120
rect 3293 3116 3297 3120
rect 3303 3116 3307 3120
rect 3373 3116 3377 3120
rect 3383 3116 3387 3120
rect 3451 3116 3455 3120
rect 3471 3116 3475 3120
rect 3491 3116 3495 3120
rect 3551 3116 3555 3120
rect 3561 3116 3565 3120
rect 3581 3116 3585 3120
rect 3686 3116 3690 3120
rect 3694 3116 3698 3120
rect 3714 3116 3718 3120
rect 3722 3116 3726 3120
rect 3785 3116 3789 3120
rect 3805 3116 3809 3120
rect 3855 3116 3859 3120
rect 3875 3116 3879 3120
rect 3885 3116 3889 3120
rect 3907 3116 3911 3120
rect 3917 3116 3921 3120
rect 3939 3116 3943 3120
rect 3985 3116 3989 3120
rect 3993 3116 3997 3120
rect 4013 3116 4017 3120
rect 4023 3116 4027 3120
rect 4045 3116 4049 3120
rect 4091 3116 4095 3120
rect 4111 3116 4115 3120
rect 4131 3116 4135 3120
rect 4228 3116 4232 3120
rect 4236 3116 4240 3120
rect 4244 3116 4248 3120
rect 4295 3116 4299 3120
rect 4315 3116 4319 3120
rect 4325 3116 4329 3120
rect 4347 3116 4351 3120
rect 4357 3116 4361 3120
rect 4379 3116 4383 3120
rect 4425 3116 4429 3120
rect 4433 3116 4437 3120
rect 4453 3116 4457 3120
rect 4463 3116 4467 3120
rect 4485 3116 4489 3120
rect 4545 3116 4549 3120
rect 4565 3116 4569 3120
rect 4585 3116 4589 3120
rect 4605 3116 4609 3120
rect 4665 3116 4669 3120
rect 4735 3116 4789 3120
rect 4834 3116 4838 3120
rect 4842 3116 4846 3120
rect 4862 3116 4866 3120
rect 4870 3116 4874 3120
rect 4965 3116 4969 3120
rect 5014 3116 5018 3120
rect 5022 3116 5026 3120
rect 5042 3116 5046 3120
rect 5050 3116 5054 3120
rect 5131 3116 5135 3120
rect 5191 3116 5195 3120
rect 5211 3116 5215 3120
rect 5275 3116 5279 3120
rect 5295 3116 5299 3120
rect 5305 3116 5309 3120
rect 5327 3116 5331 3120
rect 5337 3116 5341 3120
rect 5359 3116 5363 3120
rect 5405 3116 5409 3120
rect 5413 3116 5417 3120
rect 5433 3116 5437 3120
rect 5443 3116 5447 3120
rect 5465 3116 5469 3120
rect 5525 3116 5529 3120
rect 5545 3116 5549 3120
rect 5591 3116 5595 3120
rect 5611 3116 5615 3120
rect 5631 3116 5635 3120
rect 5728 3116 5732 3120
rect 5736 3116 5740 3120
rect 5744 3116 5748 3120
rect 5805 3116 5809 3120
rect 5825 3116 5829 3120
rect 5845 3116 5849 3120
rect 5865 3116 5869 3120
rect 5911 3116 5915 3120
rect 5971 3116 6025 3120
rect 6112 3116 6116 3120
rect 6134 3116 6138 3120
rect 6142 3116 6146 3120
rect 6205 3116 6209 3120
rect 6225 3116 6229 3120
rect 6271 3116 6275 3120
rect 6366 3116 6370 3120
rect 6374 3116 6378 3120
rect 6394 3116 6398 3120
rect 6402 3116 6406 3120
rect 6465 3116 6469 3120
rect 6511 3116 6515 3120
rect 6571 3116 6575 3120
rect 6591 3116 6595 3120
rect 6611 3116 6615 3120
rect 31 3053 35 3076
rect 51 3053 55 3076
rect 71 3056 75 3076
rect 91 3056 95 3076
rect 111 3056 115 3076
rect 131 3056 135 3076
rect 151 3056 155 3076
rect 171 3056 175 3076
rect 243 3070 247 3076
rect 243 3058 245 3070
rect 31 3041 34 3053
rect 46 3041 55 3053
rect 82 3044 95 3056
rect 122 3044 135 3056
rect 162 3044 175 3056
rect 31 2984 35 3041
rect 51 2984 55 3041
rect 71 2984 75 3044
rect 91 2984 95 3044
rect 111 2984 115 3044
rect 131 2984 135 3044
rect 151 2984 155 3044
rect 171 2984 175 3044
rect 265 3019 269 3096
rect 315 3039 319 3076
rect 335 3038 339 3096
rect 345 3064 349 3096
rect 367 3084 371 3096
rect 369 3072 371 3084
rect 377 3084 381 3096
rect 377 3072 379 3084
rect 345 3060 378 3064
rect 265 3007 274 3019
rect 243 2990 245 3002
rect 243 2984 247 2990
rect 265 2944 269 3007
rect 315 2984 319 3027
rect 335 2944 339 3026
rect 354 3011 358 3040
rect 349 3003 358 3011
rect 349 2944 353 3003
rect 374 2996 378 3060
rect 375 2984 378 2996
rect 369 2944 373 2984
rect 383 2962 387 3072
rect 399 2982 403 3096
rect 445 3092 449 3096
rect 415 3088 449 3092
rect 381 2944 385 2950
rect 401 2944 405 2970
rect 415 2962 419 3088
rect 453 3084 457 3096
rect 427 3080 457 3084
rect 439 3079 457 3080
rect 473 3075 477 3096
rect 453 3071 477 3075
rect 453 2976 459 3071
rect 483 3047 487 3096
rect 483 2989 487 3035
rect 505 3008 509 3076
rect 573 3056 577 3076
rect 563 3049 577 3056
rect 583 3056 587 3076
rect 633 3056 637 3076
rect 583 3049 591 3056
rect 563 3033 569 3049
rect 566 3021 569 3033
rect 507 2996 509 3008
rect 483 2983 491 2989
rect 505 2984 509 2996
rect 427 2950 451 2952
rect 415 2948 451 2950
rect 447 2944 451 2948
rect 455 2944 459 2976
rect 475 2924 479 2964
rect 487 2954 491 2983
rect 483 2947 491 2954
rect 483 2924 487 2947
rect 565 2944 569 3021
rect 585 3033 591 3049
rect 629 3049 637 3056
rect 643 3056 647 3076
rect 643 3049 657 3056
rect 629 3033 635 3049
rect 585 3021 594 3033
rect 626 3021 635 3033
rect 585 2944 589 3021
rect 631 2944 635 3021
rect 651 3033 657 3049
rect 651 3021 654 3033
rect 651 2944 655 3021
rect 725 2999 729 3076
rect 745 3053 749 3076
rect 765 3071 769 3076
rect 765 3064 778 3071
rect 745 3041 754 3053
rect 727 2987 734 2999
rect 730 2944 734 2987
rect 752 2984 756 3041
rect 774 3019 778 3064
rect 833 3056 837 3076
rect 823 3049 837 3056
rect 843 3056 847 3076
rect 913 3056 917 3076
rect 843 3049 851 3056
rect 823 3033 829 3049
rect 826 3021 829 3033
rect 774 2996 778 3007
rect 760 2988 778 2996
rect 760 2984 764 2988
rect 825 2944 829 3021
rect 845 3033 851 3049
rect 903 3049 917 3056
rect 923 3056 927 3076
rect 974 3072 978 3076
rect 959 3066 978 3072
rect 923 3049 931 3056
rect 959 3053 966 3066
rect 903 3033 909 3049
rect 845 3021 854 3033
rect 906 3021 909 3033
rect 845 2944 849 3021
rect 905 2944 909 3021
rect 925 3033 931 3049
rect 925 3021 934 3033
rect 925 2944 929 3021
rect 959 3004 966 3041
rect 982 3039 986 3076
rect 1004 3053 1008 3096
rect 1006 3041 1015 3053
rect 980 3004 986 3027
rect 959 2998 975 3004
rect 980 2998 995 3004
rect 971 2984 975 2998
rect 991 2984 995 2998
rect 1011 2984 1015 3041
rect 1071 3008 1075 3076
rect 1093 3047 1097 3096
rect 1103 3075 1107 3096
rect 1123 3084 1127 3096
rect 1131 3092 1135 3096
rect 1131 3088 1165 3092
rect 1123 3080 1153 3084
rect 1123 3079 1141 3080
rect 1103 3071 1127 3075
rect 1071 2996 1073 3008
rect 1071 2984 1075 2996
rect 1093 2989 1097 3035
rect 1089 2983 1097 2989
rect 1089 2954 1093 2983
rect 1121 2976 1127 3071
rect 1089 2947 1097 2954
rect 1093 2924 1097 2947
rect 1101 2924 1105 2964
rect 1121 2944 1125 2976
rect 1161 2962 1165 3088
rect 1177 2982 1181 3096
rect 1199 3084 1203 3096
rect 1201 3072 1203 3084
rect 1209 3084 1213 3096
rect 1209 3072 1211 3084
rect 1129 2950 1153 2952
rect 1129 2948 1165 2950
rect 1129 2944 1133 2948
rect 1175 2944 1179 2970
rect 1193 2962 1197 3072
rect 1231 3064 1235 3096
rect 1202 3060 1235 3064
rect 1202 2996 1206 3060
rect 1222 3011 1226 3040
rect 1241 3038 1245 3096
rect 1261 3039 1265 3076
rect 1333 3056 1337 3076
rect 1323 3049 1337 3056
rect 1343 3056 1347 3076
rect 1343 3049 1351 3056
rect 1323 3033 1329 3049
rect 1222 3003 1231 3011
rect 1202 2984 1205 2996
rect 1195 2944 1199 2950
rect 1207 2944 1211 2984
rect 1227 2944 1231 3003
rect 1241 2944 1245 3026
rect 1261 2984 1265 3027
rect 1326 3021 1329 3033
rect 1325 2944 1329 3021
rect 1345 3033 1351 3049
rect 1345 3021 1354 3033
rect 1345 2944 1349 3021
rect 1391 3008 1395 3076
rect 1413 3047 1417 3096
rect 1423 3075 1427 3096
rect 1443 3084 1447 3096
rect 1451 3092 1455 3096
rect 1451 3088 1485 3092
rect 1443 3080 1473 3084
rect 1443 3079 1461 3080
rect 1423 3071 1447 3075
rect 1391 2996 1393 3008
rect 1391 2984 1395 2996
rect 1413 2989 1417 3035
rect 1409 2983 1417 2989
rect 1409 2954 1413 2983
rect 1441 2976 1447 3071
rect 1409 2947 1417 2954
rect 1413 2924 1417 2947
rect 1421 2924 1425 2964
rect 1441 2944 1445 2976
rect 1481 2962 1485 3088
rect 1497 2982 1501 3096
rect 1519 3084 1523 3096
rect 1521 3072 1523 3084
rect 1529 3084 1533 3096
rect 1529 3072 1531 3084
rect 1449 2950 1473 2952
rect 1449 2948 1485 2950
rect 1449 2944 1453 2948
rect 1495 2944 1499 2970
rect 1513 2962 1517 3072
rect 1551 3064 1555 3096
rect 1522 3060 1555 3064
rect 1522 2996 1526 3060
rect 1542 3011 1546 3040
rect 1561 3038 1565 3096
rect 1581 3039 1585 3076
rect 1645 3039 1649 3096
rect 1645 3027 1654 3039
rect 1542 3003 1551 3011
rect 1522 2984 1525 2996
rect 1515 2944 1519 2950
rect 1527 2944 1531 2984
rect 1547 2944 1551 3003
rect 1561 2944 1565 3026
rect 1581 2984 1585 3027
rect 1645 2944 1649 3027
rect 1705 2999 1709 3076
rect 1725 3053 1729 3076
rect 1745 3071 1749 3076
rect 1745 3064 1758 3071
rect 1725 3041 1734 3053
rect 1707 2987 1714 2999
rect 1710 2944 1714 2987
rect 1732 2984 1736 3041
rect 1754 3019 1758 3064
rect 1805 3019 1809 3096
rect 1825 3019 1829 3096
rect 1895 3070 1899 3076
rect 1881 3058 1893 3070
rect 1806 3007 1821 3019
rect 1754 2996 1758 3007
rect 1740 2988 1758 2996
rect 1740 2984 1744 2988
rect 1817 2984 1821 3007
rect 1825 3007 1834 3019
rect 1825 2984 1829 3007
rect 1881 2984 1885 3058
rect 1915 3033 1919 3076
rect 1906 3021 1919 3033
rect 1903 2944 1907 3021
rect 1925 3019 1929 3076
rect 1971 3071 1975 3076
rect 1962 3064 1975 3071
rect 1962 3019 1966 3064
rect 1991 3053 1995 3076
rect 1986 3041 1995 3053
rect 1925 3007 1934 3019
rect 1925 2944 1929 3007
rect 1962 2996 1966 3007
rect 1962 2988 1980 2996
rect 1976 2984 1980 2988
rect 1984 2984 1988 3041
rect 2011 2999 2015 3076
rect 2092 3053 2096 3096
rect 2085 3041 2094 3053
rect 2006 2987 2013 2999
rect 2006 2944 2010 2987
rect 2085 2984 2089 3041
rect 2114 3039 2118 3076
rect 2122 3072 2126 3076
rect 2122 3066 2141 3072
rect 2134 3053 2141 3066
rect 2173 3056 2177 3076
rect 2169 3049 2177 3056
rect 2183 3056 2187 3076
rect 2183 3049 2197 3056
rect 2114 3004 2120 3027
rect 2134 3004 2141 3041
rect 2169 3033 2175 3049
rect 2166 3021 2175 3033
rect 2105 2998 2120 3004
rect 2125 2998 2141 3004
rect 2105 2984 2109 2998
rect 2125 2984 2129 2998
rect 2171 2944 2175 3021
rect 2191 3033 2197 3049
rect 2265 3039 2269 3096
rect 2191 3021 2194 3033
rect 2265 3027 2274 3039
rect 2191 2944 2195 3021
rect 2265 2944 2269 3027
rect 2311 3019 2315 3076
rect 2321 3033 2325 3076
rect 2341 3070 2345 3076
rect 2347 3058 2359 3070
rect 2321 3021 2334 3033
rect 2306 3007 2315 3019
rect 2311 2944 2315 3007
rect 2333 2944 2337 3021
rect 2355 2984 2359 3058
rect 2415 3039 2419 3076
rect 2435 3038 2439 3096
rect 2445 3064 2449 3096
rect 2467 3084 2471 3096
rect 2469 3072 2471 3084
rect 2477 3084 2481 3096
rect 2477 3072 2479 3084
rect 2445 3060 2478 3064
rect 2415 2984 2419 3027
rect 2435 2944 2439 3026
rect 2454 3011 2458 3040
rect 2449 3003 2458 3011
rect 2449 2944 2453 3003
rect 2474 2996 2478 3060
rect 2475 2984 2478 2996
rect 2469 2944 2473 2984
rect 2483 2962 2487 3072
rect 2499 2982 2503 3096
rect 2545 3092 2549 3096
rect 2515 3088 2549 3092
rect 2481 2944 2485 2950
rect 2501 2944 2505 2970
rect 2515 2962 2519 3088
rect 2553 3084 2557 3096
rect 2527 3080 2557 3084
rect 2539 3079 2557 3080
rect 2573 3075 2577 3096
rect 2553 3071 2577 3075
rect 2553 2976 2559 3071
rect 2583 3047 2587 3096
rect 2583 2989 2587 3035
rect 2605 3008 2609 3076
rect 2651 3039 2655 3096
rect 2646 3027 2655 3039
rect 2607 2996 2609 3008
rect 2583 2983 2591 2989
rect 2605 2984 2609 2996
rect 2527 2950 2551 2952
rect 2515 2948 2551 2950
rect 2547 2944 2551 2948
rect 2555 2944 2559 2976
rect 2575 2924 2579 2964
rect 2587 2954 2591 2983
rect 2583 2947 2591 2954
rect 2583 2924 2587 2947
rect 2651 2944 2655 3027
rect 2711 3019 2715 3096
rect 2731 3019 2735 3096
rect 2805 3039 2809 3096
rect 2805 3027 2814 3039
rect 2706 3007 2715 3019
rect 2711 2984 2715 3007
rect 2719 3007 2734 3019
rect 2719 2984 2723 3007
rect 2805 2944 2809 3027
rect 2865 2999 2869 3076
rect 2885 3053 2889 3076
rect 2905 3071 2909 3076
rect 2905 3064 2918 3071
rect 2885 3041 2894 3053
rect 2867 2987 2874 2999
rect 2870 2944 2874 2987
rect 2892 2984 2896 3041
rect 2914 3019 2918 3064
rect 2951 3053 2955 3076
rect 3133 3056 3137 3076
rect 2946 3041 2955 3053
rect 2914 2996 2918 3007
rect 2900 2988 2918 2996
rect 2900 2984 2904 2988
rect 2951 2984 2955 3041
rect 3048 2999 3052 3056
rect 3025 2987 3033 2999
rect 3045 2987 3052 2999
rect 3025 2944 3029 2987
rect 3056 2979 3060 3056
rect 3064 2999 3068 3056
rect 3123 3049 3137 3056
rect 3143 3056 3147 3076
rect 3143 3049 3151 3056
rect 3123 3033 3129 3049
rect 3126 3021 3129 3033
rect 3064 2987 3074 2999
rect 3054 2960 3060 2967
rect 3045 2956 3060 2960
rect 3074 2956 3080 2987
rect 3045 2944 3049 2956
rect 3065 2952 3080 2956
rect 3065 2944 3069 2952
rect 3125 2944 3129 3021
rect 3145 3033 3151 3049
rect 3145 3021 3154 3033
rect 3145 2944 3149 3021
rect 3205 2999 3209 3076
rect 3225 3053 3229 3076
rect 3245 3071 3249 3076
rect 3245 3064 3258 3071
rect 3225 3041 3234 3053
rect 3207 2987 3214 2999
rect 3210 2944 3214 2987
rect 3232 2984 3236 3041
rect 3254 3019 3258 3064
rect 3293 3056 3297 3076
rect 3289 3049 3297 3056
rect 3303 3056 3307 3076
rect 3373 3056 3377 3076
rect 3303 3049 3317 3056
rect 3289 3033 3295 3049
rect 3286 3021 3295 3033
rect 3254 2996 3258 3007
rect 3240 2988 3258 2996
rect 3240 2984 3244 2988
rect 3291 2944 3295 3021
rect 3311 3033 3317 3049
rect 3369 3049 3377 3056
rect 3383 3056 3387 3076
rect 3451 3071 3455 3076
rect 3442 3064 3455 3071
rect 3383 3049 3397 3056
rect 3369 3033 3375 3049
rect 3311 3021 3314 3033
rect 3366 3021 3375 3033
rect 3311 2944 3315 3021
rect 3371 2944 3375 3021
rect 3391 3033 3397 3049
rect 3391 3021 3394 3033
rect 3391 2944 3395 3021
rect 3442 3019 3446 3064
rect 3471 3053 3475 3076
rect 3466 3041 3475 3053
rect 3442 2996 3446 3007
rect 3442 2988 3460 2996
rect 3456 2984 3460 2988
rect 3464 2984 3468 3041
rect 3491 2999 3495 3076
rect 3551 3019 3555 3076
rect 3561 3033 3565 3076
rect 3581 3070 3585 3076
rect 3686 3071 3690 3076
rect 3587 3058 3599 3070
rect 3561 3021 3574 3033
rect 3546 3007 3555 3019
rect 3486 2987 3493 2999
rect 3486 2944 3490 2987
rect 3551 2944 3555 3007
rect 3573 2944 3577 3021
rect 3595 2984 3599 3058
rect 3660 3067 3690 3071
rect 3660 3019 3666 3067
rect 3694 3062 3698 3076
rect 3685 3055 3698 3062
rect 3685 3053 3689 3055
rect 3714 3053 3718 3076
rect 3722 3068 3726 3076
rect 3785 3072 3789 3076
rect 3805 3072 3809 3076
rect 3785 3068 3809 3072
rect 3722 3061 3739 3068
rect 3687 3041 3689 3053
rect 3666 3007 3669 3019
rect 3665 2984 3669 3007
rect 3685 2984 3689 3041
rect 3714 3012 3718 3041
rect 3733 3019 3739 3061
rect 3805 3053 3809 3068
rect 3805 3041 3814 3053
rect 3705 3006 3718 3012
rect 3725 3007 3733 3012
rect 3725 3006 3745 3007
rect 3705 2984 3709 3006
rect 3725 2984 3729 3006
rect 3805 2992 3809 3041
rect 3855 3039 3859 3076
rect 3875 3038 3879 3096
rect 3885 3064 3889 3096
rect 3907 3084 3911 3096
rect 3909 3072 3911 3084
rect 3917 3084 3921 3096
rect 3917 3072 3919 3084
rect 3885 3060 3918 3064
rect 3785 2988 3809 2992
rect 3785 2984 3789 2988
rect 3805 2984 3809 2988
rect 3855 2984 3859 3027
rect 3875 2944 3879 3026
rect 3894 3011 3898 3040
rect 3889 3003 3898 3011
rect 3889 2944 3893 3003
rect 3914 2996 3918 3060
rect 3915 2984 3918 2996
rect 3909 2944 3913 2984
rect 3923 2962 3927 3072
rect 3939 2982 3943 3096
rect 3985 3092 3989 3096
rect 3955 3088 3989 3092
rect 3921 2944 3925 2950
rect 3941 2944 3945 2970
rect 3955 2962 3959 3088
rect 3993 3084 3997 3096
rect 3967 3080 3997 3084
rect 3979 3079 3997 3080
rect 4013 3075 4017 3096
rect 3993 3071 4017 3075
rect 3993 2976 3999 3071
rect 4023 3047 4027 3096
rect 4023 2989 4027 3035
rect 4045 3008 4049 3076
rect 4091 3071 4095 3076
rect 4082 3064 4095 3071
rect 4082 3019 4086 3064
rect 4111 3053 4115 3076
rect 4106 3041 4115 3053
rect 4047 2996 4049 3008
rect 4023 2983 4031 2989
rect 4045 2984 4049 2996
rect 4082 2996 4086 3007
rect 4082 2988 4100 2996
rect 4096 2984 4100 2988
rect 4104 2984 4108 3041
rect 4131 2999 4135 3076
rect 4228 2999 4232 3056
rect 4126 2987 4133 2999
rect 4205 2987 4213 2999
rect 4225 2987 4232 2999
rect 3967 2950 3991 2952
rect 3955 2948 3991 2950
rect 3987 2944 3991 2948
rect 3995 2944 3999 2976
rect 4015 2924 4019 2964
rect 4027 2954 4031 2983
rect 4023 2947 4031 2954
rect 4023 2924 4027 2947
rect 4126 2944 4130 2987
rect 4205 2944 4209 2987
rect 4236 2979 4240 3056
rect 4244 2999 4248 3056
rect 4295 3039 4299 3076
rect 4315 3038 4319 3096
rect 4325 3064 4329 3096
rect 4347 3084 4351 3096
rect 4349 3072 4351 3084
rect 4357 3084 4361 3096
rect 4357 3072 4359 3084
rect 4325 3060 4358 3064
rect 4244 2987 4254 2999
rect 4234 2960 4240 2967
rect 4225 2956 4240 2960
rect 4254 2956 4260 2987
rect 4295 2984 4299 3027
rect 4225 2944 4229 2956
rect 4245 2952 4260 2956
rect 4245 2944 4249 2952
rect 4315 2944 4319 3026
rect 4334 3011 4338 3040
rect 4329 3003 4338 3011
rect 4329 2944 4333 3003
rect 4354 2996 4358 3060
rect 4355 2984 4358 2996
rect 4349 2944 4353 2984
rect 4363 2962 4367 3072
rect 4379 2982 4383 3096
rect 4425 3092 4429 3096
rect 4395 3088 4429 3092
rect 4361 2944 4365 2950
rect 4381 2944 4385 2970
rect 4395 2962 4399 3088
rect 4433 3084 4437 3096
rect 4407 3080 4437 3084
rect 4419 3079 4437 3080
rect 4453 3075 4457 3096
rect 4433 3071 4457 3075
rect 4433 2976 4439 3071
rect 4463 3047 4467 3096
rect 4725 3108 4729 3112
rect 4735 3108 4739 3116
rect 4755 3108 4759 3112
rect 4765 3108 4769 3112
rect 4785 3108 4789 3116
rect 4463 2989 4467 3035
rect 4485 3008 4489 3076
rect 4545 3019 4549 3076
rect 4565 3053 4569 3076
rect 4585 3053 4589 3076
rect 4605 3069 4609 3076
rect 4605 3065 4620 3069
rect 4585 3041 4594 3053
rect 4487 2996 4489 3008
rect 4547 3007 4549 3019
rect 4463 2983 4471 2989
rect 4485 2984 4489 2996
rect 4545 2992 4549 3007
rect 4545 2988 4559 2992
rect 4555 2984 4559 2988
rect 4565 2984 4569 3041
rect 4585 2992 4591 3041
rect 4614 3019 4620 3065
rect 4665 3039 4669 3096
rect 4785 3084 4789 3088
rect 4785 3079 4797 3084
rect 4665 3027 4674 3039
rect 4614 2992 4619 3007
rect 4585 2988 4599 2992
rect 4595 2984 4599 2988
rect 4605 2988 4619 2992
rect 4605 2984 4609 2988
rect 4407 2950 4431 2952
rect 4395 2948 4431 2950
rect 4427 2944 4431 2948
rect 4435 2944 4439 2976
rect 4455 2924 4459 2964
rect 4467 2954 4471 2983
rect 4463 2947 4471 2954
rect 4463 2924 4467 2947
rect 4665 2944 4669 3027
rect 4725 3019 4729 3068
rect 4735 3064 4739 3068
rect 4755 3022 4759 3068
rect 4765 3056 4769 3068
rect 4765 3050 4779 3056
rect 4726 3007 4729 3019
rect 4774 3019 4779 3050
rect 4793 3053 4797 3079
rect 4834 3068 4838 3076
rect 4821 3061 4838 3068
rect 4725 2984 4729 3007
rect 4735 3006 4765 3010
rect 4735 2984 4739 3006
rect 4773 3001 4778 3007
rect 4765 2997 4778 3001
rect 4755 2992 4759 2996
rect 4765 2992 4769 2997
rect 4793 2960 4797 3041
rect 4821 3019 4827 3061
rect 4842 3053 4846 3076
rect 4862 3062 4866 3076
rect 4870 3071 4874 3076
rect 4870 3067 4900 3071
rect 4862 3055 4875 3062
rect 4871 3053 4875 3055
rect 4871 3041 4873 3053
rect 4842 3012 4846 3041
rect 4827 3007 4835 3012
rect 4815 3006 4835 3007
rect 4842 3006 4855 3012
rect 4831 2984 4835 3006
rect 4851 2984 4855 3006
rect 4871 2984 4875 3041
rect 4894 3019 4900 3067
rect 4965 3039 4969 3096
rect 5014 3068 5018 3076
rect 5001 3061 5018 3068
rect 4965 3027 4974 3039
rect 4891 3007 4894 3019
rect 4891 2984 4895 3007
rect 4785 2956 4797 2960
rect 4785 2952 4789 2956
rect 4755 2904 4759 2912
rect 4765 2908 4769 2912
rect 4785 2904 4789 2912
rect 4965 2944 4969 3027
rect 5001 3019 5007 3061
rect 5022 3053 5026 3076
rect 5042 3062 5046 3076
rect 5050 3071 5054 3076
rect 5050 3067 5080 3071
rect 5042 3055 5055 3062
rect 5051 3053 5055 3055
rect 5051 3041 5053 3053
rect 5022 3012 5026 3041
rect 5007 3007 5015 3012
rect 4995 3006 5015 3007
rect 5022 3006 5035 3012
rect 5011 2984 5015 3006
rect 5031 2984 5035 3006
rect 5051 2984 5055 3041
rect 5074 3019 5080 3067
rect 5131 3039 5135 3096
rect 5126 3027 5135 3039
rect 5071 3007 5074 3019
rect 5071 2984 5075 3007
rect 5131 2944 5135 3027
rect 5191 3019 5195 3096
rect 5211 3019 5215 3096
rect 5275 3039 5279 3076
rect 5295 3038 5299 3096
rect 5305 3064 5309 3096
rect 5327 3084 5331 3096
rect 5329 3072 5331 3084
rect 5337 3084 5341 3096
rect 5337 3072 5339 3084
rect 5305 3060 5338 3064
rect 5186 3007 5195 3019
rect 5191 2984 5195 3007
rect 5199 3007 5214 3019
rect 5199 2984 5203 3007
rect 5275 2984 5279 3027
rect 5295 2944 5299 3026
rect 5314 3011 5318 3040
rect 5309 3003 5318 3011
rect 5309 2944 5313 3003
rect 5334 2996 5338 3060
rect 5335 2984 5338 2996
rect 5329 2944 5333 2984
rect 5343 2962 5347 3072
rect 5359 2982 5363 3096
rect 5405 3092 5409 3096
rect 5375 3088 5409 3092
rect 5341 2944 5345 2950
rect 5361 2944 5365 2970
rect 5375 2962 5379 3088
rect 5413 3084 5417 3096
rect 5387 3080 5417 3084
rect 5399 3079 5417 3080
rect 5433 3075 5437 3096
rect 5413 3071 5437 3075
rect 5413 2976 5419 3071
rect 5443 3047 5447 3096
rect 5443 2989 5447 3035
rect 5465 3008 5469 3076
rect 5525 3019 5529 3096
rect 5545 3019 5549 3096
rect 5591 3071 5595 3076
rect 5582 3064 5595 3071
rect 5582 3019 5586 3064
rect 5611 3053 5615 3076
rect 5606 3041 5615 3053
rect 5467 2996 5469 3008
rect 5526 3007 5541 3019
rect 5443 2983 5451 2989
rect 5465 2984 5469 2996
rect 5537 2984 5541 3007
rect 5545 3007 5554 3019
rect 5545 2984 5549 3007
rect 5582 2996 5586 3007
rect 5582 2988 5600 2996
rect 5596 2984 5600 2988
rect 5604 2984 5608 3041
rect 5631 2999 5635 3076
rect 5971 3108 5975 3116
rect 5991 3108 5995 3112
rect 6001 3108 6005 3112
rect 6021 3108 6025 3116
rect 6031 3108 6035 3112
rect 5728 2999 5732 3056
rect 5626 2987 5633 2999
rect 5705 2987 5713 2999
rect 5725 2987 5732 2999
rect 5387 2950 5411 2952
rect 5375 2948 5411 2950
rect 5407 2944 5411 2948
rect 5415 2944 5419 2976
rect 5435 2924 5439 2964
rect 5447 2954 5451 2983
rect 5443 2947 5451 2954
rect 5443 2924 5447 2947
rect 5626 2944 5630 2987
rect 5705 2944 5709 2987
rect 5736 2979 5740 3056
rect 5744 2999 5748 3056
rect 5805 3019 5809 3076
rect 5825 3053 5829 3076
rect 5845 3053 5849 3076
rect 5865 3069 5869 3076
rect 5865 3065 5880 3069
rect 5845 3041 5854 3053
rect 5807 3007 5809 3019
rect 5744 2987 5754 2999
rect 5805 2992 5809 3007
rect 5805 2988 5819 2992
rect 5734 2960 5740 2967
rect 5725 2956 5740 2960
rect 5754 2956 5760 2987
rect 5815 2984 5819 2988
rect 5825 2984 5829 3041
rect 5845 2992 5851 3041
rect 5874 3019 5880 3065
rect 5911 3039 5915 3096
rect 5971 3084 5975 3088
rect 5963 3079 5975 3084
rect 5963 3053 5967 3079
rect 5991 3056 5995 3068
rect 5906 3027 5915 3039
rect 5874 2992 5879 3007
rect 5845 2988 5859 2992
rect 5855 2984 5859 2988
rect 5865 2988 5879 2992
rect 5865 2984 5869 2988
rect 5725 2944 5729 2956
rect 5745 2952 5760 2956
rect 5745 2944 5749 2952
rect 5911 2944 5915 3027
rect 5963 2960 5967 3041
rect 5981 3050 5995 3056
rect 5981 3019 5986 3050
rect 6001 3022 6005 3068
rect 6021 3064 6025 3068
rect 5982 3001 5987 3007
rect 6031 3019 6035 3068
rect 6112 3053 6116 3096
rect 6105 3041 6114 3053
rect 5995 3006 6025 3010
rect 5982 2997 5995 3001
rect 5991 2992 5995 2997
rect 6001 2992 6005 2996
rect 5963 2956 5975 2960
rect 5971 2952 5975 2956
rect 6021 2984 6025 3006
rect 6031 3007 6034 3019
rect 6031 2984 6035 3007
rect 6105 2984 6109 3041
rect 6134 3039 6138 3076
rect 6142 3072 6146 3076
rect 6142 3066 6161 3072
rect 6154 3053 6161 3066
rect 6134 3004 6140 3027
rect 6154 3004 6161 3041
rect 6205 3019 6209 3096
rect 6225 3019 6229 3096
rect 6271 3039 6275 3096
rect 6366 3071 6370 3076
rect 6266 3027 6275 3039
rect 6206 3007 6221 3019
rect 6125 2998 6140 3004
rect 6145 2998 6161 3004
rect 6125 2984 6129 2998
rect 6145 2984 6149 2998
rect 6217 2984 6221 3007
rect 6225 3007 6234 3019
rect 6225 2984 6229 3007
rect 5971 2904 5975 2912
rect 5991 2908 5995 2912
rect 6001 2904 6005 2912
rect 6271 2944 6275 3027
rect 6340 3067 6370 3071
rect 6340 3019 6346 3067
rect 6374 3062 6378 3076
rect 6365 3055 6378 3062
rect 6365 3053 6369 3055
rect 6394 3053 6398 3076
rect 6402 3068 6406 3076
rect 6402 3061 6419 3068
rect 6367 3041 6369 3053
rect 6346 3007 6349 3019
rect 6345 2984 6349 3007
rect 6365 2984 6369 3041
rect 6394 3012 6398 3041
rect 6413 3019 6419 3061
rect 6465 3039 6469 3096
rect 6511 3039 6515 3096
rect 6571 3071 6575 3076
rect 6465 3027 6474 3039
rect 6506 3027 6515 3039
rect 6385 3006 6398 3012
rect 6405 3007 6413 3012
rect 6405 3006 6425 3007
rect 6385 2984 6389 3006
rect 6405 2984 6409 3006
rect 6465 2944 6469 3027
rect 6511 2944 6515 3027
rect 6562 3064 6575 3071
rect 6562 3019 6566 3064
rect 6591 3053 6595 3076
rect 6586 3041 6595 3053
rect 6562 2996 6566 3007
rect 6562 2988 6580 2996
rect 6576 2984 6580 2988
rect 6584 2984 6588 3041
rect 6611 2999 6615 3076
rect 6606 2987 6613 2999
rect 6606 2944 6610 2987
rect 31 2900 35 2904
rect 51 2900 55 2904
rect 71 2900 75 2904
rect 91 2900 95 2904
rect 111 2900 115 2904
rect 131 2900 135 2904
rect 151 2900 155 2904
rect 171 2900 175 2904
rect 243 2900 247 2904
rect 265 2900 269 2904
rect 315 2900 319 2904
rect 335 2900 339 2904
rect 349 2900 353 2904
rect 369 2900 373 2904
rect 381 2900 385 2904
rect 401 2900 405 2904
rect 447 2900 451 2904
rect 455 2900 459 2904
rect 475 2900 479 2904
rect 483 2900 487 2904
rect 505 2900 509 2904
rect 565 2900 569 2904
rect 585 2900 589 2904
rect 631 2900 635 2904
rect 651 2900 655 2904
rect 730 2900 734 2904
rect 752 2900 756 2904
rect 760 2900 764 2904
rect 825 2900 829 2904
rect 845 2900 849 2904
rect 905 2900 909 2904
rect 925 2900 929 2904
rect 971 2900 975 2904
rect 991 2900 995 2904
rect 1011 2900 1015 2904
rect 1071 2900 1075 2904
rect 1093 2900 1097 2904
rect 1101 2900 1105 2904
rect 1121 2900 1125 2904
rect 1129 2900 1133 2904
rect 1175 2900 1179 2904
rect 1195 2900 1199 2904
rect 1207 2900 1211 2904
rect 1227 2900 1231 2904
rect 1241 2900 1245 2904
rect 1261 2900 1265 2904
rect 1325 2900 1329 2904
rect 1345 2900 1349 2904
rect 1391 2900 1395 2904
rect 1413 2900 1417 2904
rect 1421 2900 1425 2904
rect 1441 2900 1445 2904
rect 1449 2900 1453 2904
rect 1495 2900 1499 2904
rect 1515 2900 1519 2904
rect 1527 2900 1531 2904
rect 1547 2900 1551 2904
rect 1561 2900 1565 2904
rect 1581 2900 1585 2904
rect 1645 2900 1649 2904
rect 1710 2900 1714 2904
rect 1732 2900 1736 2904
rect 1740 2900 1744 2904
rect 1817 2900 1821 2904
rect 1825 2900 1829 2904
rect 1881 2900 1885 2904
rect 1903 2900 1907 2904
rect 1925 2900 1929 2904
rect 1976 2900 1980 2904
rect 1984 2900 1988 2904
rect 2006 2900 2010 2904
rect 2085 2900 2089 2904
rect 2105 2900 2109 2904
rect 2125 2900 2129 2904
rect 2171 2900 2175 2904
rect 2191 2900 2195 2904
rect 2265 2900 2269 2904
rect 2311 2900 2315 2904
rect 2333 2900 2337 2904
rect 2355 2900 2359 2904
rect 2415 2900 2419 2904
rect 2435 2900 2439 2904
rect 2449 2900 2453 2904
rect 2469 2900 2473 2904
rect 2481 2900 2485 2904
rect 2501 2900 2505 2904
rect 2547 2900 2551 2904
rect 2555 2900 2559 2904
rect 2575 2900 2579 2904
rect 2583 2900 2587 2904
rect 2605 2900 2609 2904
rect 2651 2900 2655 2904
rect 2711 2900 2715 2904
rect 2719 2900 2723 2904
rect 2805 2900 2809 2904
rect 2870 2900 2874 2904
rect 2892 2900 2896 2904
rect 2900 2900 2904 2904
rect 2951 2900 2955 2904
rect 3025 2900 3029 2904
rect 3045 2900 3049 2904
rect 3065 2900 3069 2904
rect 3125 2900 3129 2904
rect 3145 2900 3149 2904
rect 3210 2900 3214 2904
rect 3232 2900 3236 2904
rect 3240 2900 3244 2904
rect 3291 2900 3295 2904
rect 3311 2900 3315 2904
rect 3371 2900 3375 2904
rect 3391 2900 3395 2904
rect 3456 2900 3460 2904
rect 3464 2900 3468 2904
rect 3486 2900 3490 2904
rect 3551 2900 3555 2904
rect 3573 2900 3577 2904
rect 3595 2900 3599 2904
rect 3665 2900 3669 2904
rect 3685 2900 3689 2904
rect 3705 2900 3709 2904
rect 3725 2900 3729 2904
rect 3785 2900 3789 2904
rect 3805 2900 3809 2904
rect 3855 2900 3859 2904
rect 3875 2900 3879 2904
rect 3889 2900 3893 2904
rect 3909 2900 3913 2904
rect 3921 2900 3925 2904
rect 3941 2900 3945 2904
rect 3987 2900 3991 2904
rect 3995 2900 3999 2904
rect 4015 2900 4019 2904
rect 4023 2900 4027 2904
rect 4045 2900 4049 2904
rect 4096 2900 4100 2904
rect 4104 2900 4108 2904
rect 4126 2900 4130 2904
rect 4205 2900 4209 2904
rect 4225 2900 4229 2904
rect 4245 2900 4249 2904
rect 4295 2900 4299 2904
rect 4315 2900 4319 2904
rect 4329 2900 4333 2904
rect 4349 2900 4353 2904
rect 4361 2900 4365 2904
rect 4381 2900 4385 2904
rect 4427 2900 4431 2904
rect 4435 2900 4439 2904
rect 4455 2900 4459 2904
rect 4463 2900 4467 2904
rect 4485 2900 4489 2904
rect 4555 2900 4559 2904
rect 4565 2900 4569 2904
rect 4595 2900 4599 2904
rect 4605 2900 4609 2904
rect 4665 2900 4669 2904
rect 4725 2900 4729 2904
rect 4735 2900 4739 2904
rect 4755 2900 4789 2904
rect 4831 2900 4835 2904
rect 4851 2900 4855 2904
rect 4871 2900 4875 2904
rect 4891 2900 4895 2904
rect 4965 2900 4969 2904
rect 5011 2900 5015 2904
rect 5031 2900 5035 2904
rect 5051 2900 5055 2904
rect 5071 2900 5075 2904
rect 5131 2900 5135 2904
rect 5191 2900 5195 2904
rect 5199 2900 5203 2904
rect 5275 2900 5279 2904
rect 5295 2900 5299 2904
rect 5309 2900 5313 2904
rect 5329 2900 5333 2904
rect 5341 2900 5345 2904
rect 5361 2900 5365 2904
rect 5407 2900 5411 2904
rect 5415 2900 5419 2904
rect 5435 2900 5439 2904
rect 5443 2900 5447 2904
rect 5465 2900 5469 2904
rect 5537 2900 5541 2904
rect 5545 2900 5549 2904
rect 5596 2900 5600 2904
rect 5604 2900 5608 2904
rect 5626 2900 5630 2904
rect 5705 2900 5709 2904
rect 5725 2900 5729 2904
rect 5745 2900 5749 2904
rect 5815 2900 5819 2904
rect 5825 2900 5829 2904
rect 5855 2900 5859 2904
rect 5865 2900 5869 2904
rect 5911 2900 5915 2904
rect 5971 2900 6005 2904
rect 6021 2900 6025 2904
rect 6031 2900 6035 2904
rect 6105 2900 6109 2904
rect 6125 2900 6129 2904
rect 6145 2900 6149 2904
rect 6217 2900 6221 2904
rect 6225 2900 6229 2904
rect 6271 2900 6275 2904
rect 6345 2900 6349 2904
rect 6365 2900 6369 2904
rect 6385 2900 6389 2904
rect 6405 2900 6409 2904
rect 6465 2900 6469 2904
rect 6511 2900 6515 2904
rect 6576 2900 6580 2904
rect 6584 2900 6588 2904
rect 6606 2900 6610 2904
rect 31 2876 35 2880
rect 117 2876 121 2880
rect 125 2876 129 2880
rect 175 2876 179 2880
rect 195 2876 199 2880
rect 209 2876 213 2880
rect 229 2876 233 2880
rect 241 2876 245 2880
rect 261 2876 265 2880
rect 307 2876 311 2880
rect 315 2876 319 2880
rect 335 2876 339 2880
rect 343 2876 347 2880
rect 365 2876 369 2880
rect 411 2876 415 2880
rect 497 2876 501 2880
rect 505 2876 509 2880
rect 555 2876 559 2880
rect 575 2876 579 2880
rect 589 2876 593 2880
rect 609 2876 613 2880
rect 621 2876 625 2880
rect 641 2876 645 2880
rect 687 2876 691 2880
rect 695 2876 699 2880
rect 715 2876 719 2880
rect 723 2876 727 2880
rect 745 2876 749 2880
rect 803 2876 807 2880
rect 825 2876 829 2880
rect 871 2876 875 2880
rect 891 2876 895 2880
rect 951 2876 955 2880
rect 971 2876 975 2880
rect 1031 2876 1035 2880
rect 1051 2876 1055 2880
rect 1111 2876 1115 2880
rect 1171 2876 1175 2880
rect 1191 2876 1195 2880
rect 1211 2876 1215 2880
rect 1231 2876 1235 2880
rect 1305 2876 1309 2880
rect 1325 2876 1329 2880
rect 1345 2876 1349 2880
rect 1405 2876 1409 2880
rect 1470 2876 1474 2880
rect 1492 2876 1496 2880
rect 1500 2876 1504 2880
rect 1551 2876 1555 2880
rect 1559 2876 1563 2880
rect 1631 2876 1635 2880
rect 1651 2876 1655 2880
rect 1711 2876 1715 2880
rect 1719 2876 1723 2880
rect 1810 2876 1814 2880
rect 1832 2876 1836 2880
rect 1840 2876 1844 2880
rect 1891 2876 1895 2880
rect 1901 2876 1905 2880
rect 1921 2876 1925 2880
rect 1996 2876 2000 2880
rect 2004 2876 2008 2880
rect 2026 2876 2030 2880
rect 2105 2876 2109 2880
rect 2125 2876 2129 2880
rect 2145 2876 2149 2880
rect 2195 2876 2199 2880
rect 2215 2876 2219 2880
rect 2229 2876 2233 2880
rect 2249 2876 2253 2880
rect 2261 2876 2265 2880
rect 2281 2876 2285 2880
rect 2327 2876 2331 2880
rect 2335 2876 2339 2880
rect 2355 2876 2359 2880
rect 2363 2876 2367 2880
rect 2385 2876 2389 2880
rect 2431 2876 2435 2880
rect 2451 2876 2455 2880
rect 2511 2876 2515 2880
rect 2585 2876 2589 2880
rect 2635 2876 2639 2880
rect 2655 2876 2659 2880
rect 2669 2876 2673 2880
rect 2689 2876 2693 2880
rect 2701 2876 2705 2880
rect 2721 2876 2725 2880
rect 2767 2876 2771 2880
rect 2775 2876 2779 2880
rect 2795 2876 2799 2880
rect 2803 2876 2807 2880
rect 2825 2876 2829 2880
rect 2876 2876 2880 2880
rect 2884 2876 2888 2880
rect 2906 2876 2910 2880
rect 2985 2876 2989 2880
rect 3005 2876 3009 2880
rect 3025 2876 3029 2880
rect 3071 2876 3075 2880
rect 3093 2876 3097 2880
rect 3101 2876 3105 2880
rect 3121 2876 3125 2880
rect 3129 2876 3133 2880
rect 3175 2876 3179 2880
rect 3195 2876 3199 2880
rect 3207 2876 3211 2880
rect 3227 2876 3231 2880
rect 3241 2876 3245 2880
rect 3261 2876 3265 2880
rect 3311 2876 3315 2880
rect 3371 2876 3375 2880
rect 3381 2876 3385 2880
rect 3411 2876 3415 2880
rect 3421 2876 3425 2880
rect 3496 2876 3500 2880
rect 3504 2876 3508 2880
rect 3526 2876 3530 2880
rect 3615 2876 3619 2880
rect 3625 2876 3629 2880
rect 3655 2876 3659 2880
rect 3665 2876 3669 2880
rect 3716 2876 3720 2880
rect 3724 2876 3728 2880
rect 3746 2876 3750 2880
rect 3835 2876 3839 2880
rect 3845 2876 3849 2880
rect 3875 2876 3879 2880
rect 3885 2876 3889 2880
rect 3945 2876 3949 2880
rect 3991 2876 3995 2880
rect 3999 2876 4003 2880
rect 4071 2876 4075 2880
rect 4079 2876 4083 2880
rect 4165 2876 4169 2880
rect 4185 2876 4189 2880
rect 4205 2876 4209 2880
rect 4256 2876 4260 2880
rect 4264 2876 4268 2880
rect 4286 2876 4290 2880
rect 4365 2876 4369 2880
rect 4385 2876 4389 2880
rect 4405 2876 4409 2880
rect 4455 2876 4459 2880
rect 4475 2876 4479 2880
rect 4489 2876 4493 2880
rect 4509 2876 4513 2880
rect 4521 2876 4525 2880
rect 4541 2876 4545 2880
rect 4587 2876 4591 2880
rect 4595 2876 4599 2880
rect 4615 2876 4619 2880
rect 4623 2876 4627 2880
rect 4645 2876 4649 2880
rect 4691 2876 4695 2880
rect 4751 2876 4755 2880
rect 4759 2876 4763 2880
rect 4836 2876 4840 2880
rect 4844 2876 4848 2880
rect 4866 2876 4870 2880
rect 4957 2876 4961 2880
rect 4965 2876 4969 2880
rect 5035 2876 5039 2880
rect 5045 2876 5049 2880
rect 5075 2876 5079 2880
rect 5085 2876 5089 2880
rect 5131 2876 5135 2880
rect 5151 2876 5155 2880
rect 5171 2876 5175 2880
rect 5231 2876 5235 2880
rect 5253 2876 5257 2880
rect 5316 2876 5320 2880
rect 5324 2876 5328 2880
rect 5346 2876 5350 2880
rect 5435 2876 5439 2880
rect 5445 2876 5449 2880
rect 5475 2876 5479 2880
rect 5485 2876 5489 2880
rect 5545 2876 5549 2880
rect 5595 2876 5599 2880
rect 5615 2876 5619 2880
rect 5629 2876 5633 2880
rect 5649 2876 5653 2880
rect 5661 2876 5665 2880
rect 5681 2876 5685 2880
rect 5727 2876 5731 2880
rect 5735 2876 5739 2880
rect 5755 2876 5759 2880
rect 5763 2876 5767 2880
rect 5785 2876 5789 2880
rect 5831 2876 5865 2880
rect 5881 2876 5885 2880
rect 5891 2876 5895 2880
rect 5951 2876 5985 2880
rect 6001 2876 6005 2880
rect 6011 2876 6015 2880
rect 6071 2876 6105 2880
rect 6121 2876 6125 2880
rect 6131 2876 6135 2880
rect 6201 2876 6205 2880
rect 6223 2876 6227 2880
rect 6245 2876 6249 2880
rect 6305 2876 6309 2880
rect 6325 2876 6329 2880
rect 6371 2876 6375 2880
rect 6393 2876 6397 2880
rect 6415 2876 6419 2880
rect 6471 2876 6475 2880
rect 6493 2876 6497 2880
rect 6501 2876 6505 2880
rect 6521 2876 6525 2880
rect 6529 2876 6533 2880
rect 6575 2876 6579 2880
rect 6595 2876 6599 2880
rect 6607 2876 6611 2880
rect 6627 2876 6631 2880
rect 6641 2876 6645 2880
rect 6661 2876 6665 2880
rect 31 2753 35 2836
rect 117 2773 121 2796
rect 106 2761 121 2773
rect 125 2773 129 2796
rect 125 2761 134 2773
rect 26 2741 35 2753
rect 31 2684 35 2741
rect 105 2684 109 2761
rect 125 2684 129 2761
rect 175 2753 179 2796
rect 195 2754 199 2836
rect 209 2777 213 2836
rect 229 2796 233 2836
rect 241 2830 245 2836
rect 235 2784 238 2796
rect 209 2769 218 2777
rect 175 2704 179 2741
rect 195 2684 199 2742
rect 214 2740 218 2769
rect 234 2720 238 2784
rect 205 2716 238 2720
rect 205 2684 209 2716
rect 243 2708 247 2818
rect 261 2810 265 2836
rect 307 2832 311 2836
rect 275 2830 311 2832
rect 287 2828 311 2830
rect 229 2696 231 2708
rect 227 2684 231 2696
rect 237 2696 239 2708
rect 237 2684 241 2696
rect 259 2684 263 2798
rect 275 2692 279 2818
rect 315 2804 319 2836
rect 335 2816 339 2856
rect 343 2833 347 2856
rect 343 2826 351 2833
rect 313 2709 319 2804
rect 347 2797 351 2826
rect 343 2791 351 2797
rect 343 2745 347 2791
rect 365 2784 369 2796
rect 367 2772 369 2784
rect 313 2705 337 2709
rect 299 2700 317 2701
rect 287 2696 317 2700
rect 275 2688 309 2692
rect 305 2684 309 2688
rect 313 2684 317 2696
rect 333 2684 337 2705
rect 343 2684 347 2733
rect 365 2704 369 2772
rect 411 2753 415 2836
rect 497 2773 501 2796
rect 486 2761 501 2773
rect 505 2773 509 2796
rect 505 2761 514 2773
rect 406 2741 415 2753
rect 411 2684 415 2741
rect 485 2684 489 2761
rect 505 2684 509 2761
rect 555 2753 559 2796
rect 575 2754 579 2836
rect 589 2777 593 2836
rect 609 2796 613 2836
rect 621 2830 625 2836
rect 615 2784 618 2796
rect 589 2769 598 2777
rect 555 2704 559 2741
rect 575 2684 579 2742
rect 594 2740 598 2769
rect 614 2720 618 2784
rect 585 2716 618 2720
rect 585 2684 589 2716
rect 623 2708 627 2818
rect 641 2810 645 2836
rect 687 2832 691 2836
rect 655 2830 691 2832
rect 667 2828 691 2830
rect 609 2696 611 2708
rect 607 2684 611 2696
rect 617 2696 619 2708
rect 617 2684 621 2696
rect 639 2684 643 2798
rect 655 2692 659 2818
rect 695 2804 699 2836
rect 715 2816 719 2856
rect 723 2833 727 2856
rect 723 2826 731 2833
rect 693 2709 699 2804
rect 727 2797 731 2826
rect 723 2791 731 2797
rect 723 2745 727 2791
rect 745 2784 749 2796
rect 747 2772 749 2784
rect 803 2790 807 2796
rect 803 2778 805 2790
rect 693 2705 717 2709
rect 679 2700 697 2701
rect 667 2696 697 2700
rect 655 2688 689 2692
rect 685 2684 689 2688
rect 693 2684 697 2696
rect 713 2684 717 2705
rect 723 2684 727 2733
rect 745 2704 749 2772
rect 825 2773 829 2836
rect 871 2792 875 2796
rect 891 2792 895 2796
rect 871 2788 895 2792
rect 825 2761 834 2773
rect 803 2710 805 2722
rect 803 2704 807 2710
rect 825 2684 829 2761
rect 871 2739 875 2788
rect 951 2759 955 2836
rect 946 2747 955 2759
rect 866 2727 875 2739
rect 871 2712 875 2727
rect 949 2731 955 2747
rect 971 2759 975 2836
rect 1031 2759 1035 2836
rect 971 2747 974 2759
rect 1026 2747 1035 2759
rect 971 2731 977 2747
rect 949 2724 957 2731
rect 871 2708 895 2712
rect 871 2704 875 2708
rect 891 2704 895 2708
rect 953 2704 957 2724
rect 963 2724 977 2731
rect 1029 2731 1035 2747
rect 1051 2759 1055 2836
rect 1051 2747 1054 2759
rect 1111 2753 1115 2836
rect 1171 2774 1175 2796
rect 1191 2774 1195 2796
rect 1155 2773 1175 2774
rect 1167 2768 1175 2773
rect 1182 2768 1195 2774
rect 1051 2731 1057 2747
rect 1106 2741 1115 2753
rect 1029 2724 1037 2731
rect 963 2704 967 2724
rect 1033 2704 1037 2724
rect 1043 2724 1057 2731
rect 1043 2704 1047 2724
rect 1111 2684 1115 2741
rect 1161 2719 1167 2761
rect 1182 2739 1186 2768
rect 1211 2739 1215 2796
rect 1231 2773 1235 2796
rect 1231 2761 1234 2773
rect 1211 2727 1213 2739
rect 1161 2712 1178 2719
rect 1174 2704 1178 2712
rect 1182 2704 1186 2727
rect 1211 2725 1215 2727
rect 1202 2718 1215 2725
rect 1202 2704 1206 2718
rect 1234 2713 1240 2761
rect 1305 2739 1309 2796
rect 1325 2782 1329 2796
rect 1345 2782 1349 2796
rect 1325 2776 1340 2782
rect 1345 2776 1361 2782
rect 1334 2753 1340 2776
rect 1305 2727 1314 2739
rect 1210 2709 1240 2713
rect 1210 2704 1214 2709
rect 1312 2684 1316 2727
rect 1334 2704 1338 2741
rect 1354 2739 1361 2776
rect 1405 2753 1409 2836
rect 1470 2793 1474 2836
rect 1467 2781 1474 2793
rect 1405 2741 1414 2753
rect 1354 2714 1361 2727
rect 1342 2708 1361 2714
rect 1342 2704 1346 2708
rect 1405 2684 1409 2741
rect 1465 2704 1469 2781
rect 1492 2739 1496 2796
rect 1500 2792 1504 2796
rect 1500 2784 1518 2792
rect 1514 2773 1518 2784
rect 1551 2773 1555 2796
rect 1546 2761 1555 2773
rect 1559 2773 1563 2796
rect 1559 2761 1574 2773
rect 1485 2727 1494 2739
rect 1485 2704 1489 2727
rect 1514 2716 1518 2761
rect 1505 2709 1518 2716
rect 1505 2704 1509 2709
rect 1551 2684 1555 2761
rect 1571 2684 1575 2761
rect 1631 2759 1635 2836
rect 1626 2747 1635 2759
rect 1629 2731 1635 2747
rect 1651 2759 1655 2836
rect 1711 2773 1715 2796
rect 1706 2761 1715 2773
rect 1719 2773 1723 2796
rect 1810 2793 1814 2836
rect 1807 2781 1814 2793
rect 1719 2761 1734 2773
rect 1651 2747 1654 2759
rect 1651 2731 1657 2747
rect 1629 2724 1637 2731
rect 1633 2704 1637 2724
rect 1643 2724 1657 2731
rect 1643 2704 1647 2724
rect 1711 2684 1715 2761
rect 1731 2684 1735 2761
rect 1805 2704 1809 2781
rect 1832 2739 1836 2796
rect 1840 2792 1844 2796
rect 1891 2792 1895 2796
rect 1840 2784 1858 2792
rect 1854 2773 1858 2784
rect 1882 2787 1895 2792
rect 1825 2727 1834 2739
rect 1825 2704 1829 2727
rect 1854 2716 1858 2761
rect 1882 2753 1886 2787
rect 1901 2773 1905 2796
rect 1921 2791 1925 2796
rect 1996 2792 2000 2796
rect 1982 2784 2000 2792
rect 1982 2773 1986 2784
rect 1845 2709 1858 2716
rect 1845 2704 1849 2709
rect 1882 2696 1886 2741
rect 1901 2697 1905 2761
rect 1925 2712 1935 2724
rect 1931 2704 1935 2712
rect 1982 2716 1986 2761
rect 2004 2739 2008 2796
rect 2026 2793 2030 2836
rect 2026 2781 2033 2793
rect 2006 2727 2015 2739
rect 1982 2709 1995 2716
rect 1991 2704 1995 2709
rect 2011 2704 2015 2727
rect 2031 2704 2035 2781
rect 2105 2739 2109 2796
rect 2125 2782 2129 2796
rect 2145 2782 2149 2796
rect 2125 2776 2140 2782
rect 2145 2776 2161 2782
rect 2134 2753 2140 2776
rect 2105 2727 2114 2739
rect 1882 2691 1895 2696
rect 1901 2691 1915 2697
rect 1891 2684 1895 2691
rect 1911 2684 1915 2691
rect 2112 2684 2116 2727
rect 2134 2704 2138 2741
rect 2154 2739 2161 2776
rect 2195 2753 2199 2796
rect 2215 2754 2219 2836
rect 2229 2777 2233 2836
rect 2249 2796 2253 2836
rect 2261 2830 2265 2836
rect 2255 2784 2258 2796
rect 2229 2769 2238 2777
rect 2154 2714 2161 2727
rect 2142 2708 2161 2714
rect 2142 2704 2146 2708
rect 2195 2704 2199 2741
rect 2215 2684 2219 2742
rect 2234 2740 2238 2769
rect 2254 2720 2258 2784
rect 2225 2716 2258 2720
rect 2225 2684 2229 2716
rect 2263 2708 2267 2818
rect 2281 2810 2285 2836
rect 2327 2832 2331 2836
rect 2295 2830 2331 2832
rect 2307 2828 2331 2830
rect 2249 2696 2251 2708
rect 2247 2684 2251 2696
rect 2257 2696 2259 2708
rect 2257 2684 2261 2696
rect 2279 2684 2283 2798
rect 2295 2692 2299 2818
rect 2335 2804 2339 2836
rect 2355 2816 2359 2856
rect 2363 2833 2367 2856
rect 2363 2826 2371 2833
rect 2333 2709 2339 2804
rect 2367 2797 2371 2826
rect 2363 2791 2371 2797
rect 2363 2745 2367 2791
rect 2385 2784 2389 2796
rect 2387 2772 2389 2784
rect 2333 2705 2357 2709
rect 2319 2700 2337 2701
rect 2307 2696 2337 2700
rect 2295 2688 2329 2692
rect 2325 2684 2329 2688
rect 2333 2684 2337 2696
rect 2353 2684 2357 2705
rect 2363 2684 2367 2733
rect 2385 2704 2389 2772
rect 2431 2759 2435 2836
rect 2426 2747 2435 2759
rect 2429 2731 2435 2747
rect 2451 2759 2455 2836
rect 2451 2747 2454 2759
rect 2511 2753 2515 2836
rect 2451 2731 2457 2747
rect 2506 2741 2515 2753
rect 2429 2724 2437 2731
rect 2433 2704 2437 2724
rect 2443 2724 2457 2731
rect 2443 2704 2447 2724
rect 2511 2684 2515 2741
rect 2585 2753 2589 2836
rect 2635 2753 2639 2796
rect 2655 2754 2659 2836
rect 2669 2777 2673 2836
rect 2689 2796 2693 2836
rect 2701 2830 2705 2836
rect 2695 2784 2698 2796
rect 2669 2769 2678 2777
rect 2585 2741 2594 2753
rect 2585 2684 2589 2741
rect 2635 2704 2639 2741
rect 2655 2684 2659 2742
rect 2674 2740 2678 2769
rect 2694 2720 2698 2784
rect 2665 2716 2698 2720
rect 2665 2684 2669 2716
rect 2703 2708 2707 2818
rect 2721 2810 2725 2836
rect 2767 2832 2771 2836
rect 2735 2830 2771 2832
rect 2747 2828 2771 2830
rect 2689 2696 2691 2708
rect 2687 2684 2691 2696
rect 2697 2696 2699 2708
rect 2697 2684 2701 2696
rect 2719 2684 2723 2798
rect 2735 2692 2739 2818
rect 2775 2804 2779 2836
rect 2795 2816 2799 2856
rect 2803 2833 2807 2856
rect 2803 2826 2811 2833
rect 2773 2709 2779 2804
rect 2807 2797 2811 2826
rect 2803 2791 2811 2797
rect 2803 2745 2807 2791
rect 2825 2784 2829 2796
rect 2876 2792 2880 2796
rect 2827 2772 2829 2784
rect 2862 2784 2880 2792
rect 2862 2773 2866 2784
rect 2773 2705 2797 2709
rect 2759 2700 2777 2701
rect 2747 2696 2777 2700
rect 2735 2688 2769 2692
rect 2765 2684 2769 2688
rect 2773 2684 2777 2696
rect 2793 2684 2797 2705
rect 2803 2684 2807 2733
rect 2825 2704 2829 2772
rect 2862 2716 2866 2761
rect 2884 2739 2888 2796
rect 2906 2793 2910 2836
rect 3093 2833 3097 2856
rect 3089 2826 3097 2833
rect 3089 2797 3093 2826
rect 3101 2816 3105 2856
rect 3121 2804 3125 2836
rect 3129 2832 3133 2836
rect 3129 2830 3165 2832
rect 3129 2828 3153 2830
rect 2906 2781 2913 2793
rect 2886 2727 2895 2739
rect 2862 2709 2875 2716
rect 2871 2704 2875 2709
rect 2891 2704 2895 2727
rect 2911 2704 2915 2781
rect 2985 2739 2989 2796
rect 3005 2782 3009 2796
rect 3025 2782 3029 2796
rect 3071 2784 3075 2796
rect 3089 2791 3097 2797
rect 3005 2776 3020 2782
rect 3025 2776 3041 2782
rect 3014 2753 3020 2776
rect 2985 2727 2994 2739
rect 2992 2684 2996 2727
rect 3014 2704 3018 2741
rect 3034 2739 3041 2776
rect 3071 2772 3073 2784
rect 3034 2714 3041 2727
rect 3022 2708 3041 2714
rect 3022 2704 3026 2708
rect 3071 2704 3075 2772
rect 3093 2745 3097 2791
rect 3093 2684 3097 2733
rect 3121 2709 3127 2804
rect 3103 2705 3127 2709
rect 3103 2684 3107 2705
rect 3123 2700 3141 2701
rect 3123 2696 3153 2700
rect 3123 2684 3127 2696
rect 3161 2692 3165 2818
rect 3175 2810 3179 2836
rect 3195 2830 3199 2836
rect 3131 2688 3165 2692
rect 3131 2684 3135 2688
rect 3177 2684 3181 2798
rect 3193 2708 3197 2818
rect 3207 2796 3211 2836
rect 3202 2784 3205 2796
rect 3202 2720 3206 2784
rect 3227 2777 3231 2836
rect 3222 2769 3231 2777
rect 3222 2740 3226 2769
rect 3241 2754 3245 2836
rect 3261 2753 3265 2796
rect 3311 2753 3315 2836
rect 3371 2792 3375 2796
rect 3361 2788 3375 2792
rect 3381 2792 3385 2796
rect 3381 2788 3395 2792
rect 3361 2773 3366 2788
rect 3202 2716 3235 2720
rect 3201 2696 3203 2708
rect 3199 2684 3203 2696
rect 3209 2696 3211 2708
rect 3209 2684 3213 2696
rect 3231 2684 3235 2716
rect 3241 2684 3245 2742
rect 3306 2741 3315 2753
rect 3261 2704 3265 2741
rect 3311 2684 3315 2741
rect 3360 2715 3366 2761
rect 3389 2739 3395 2788
rect 3411 2739 3415 2796
rect 3421 2792 3425 2796
rect 3496 2792 3500 2796
rect 3421 2788 3435 2792
rect 3431 2773 3435 2788
rect 3482 2784 3500 2792
rect 3482 2773 3486 2784
rect 3431 2761 3433 2773
rect 3386 2727 3395 2739
rect 3360 2711 3375 2715
rect 3371 2704 3375 2711
rect 3391 2704 3395 2727
rect 3411 2704 3415 2727
rect 3431 2704 3435 2761
rect 3482 2716 3486 2761
rect 3504 2739 3508 2796
rect 3526 2793 3530 2836
rect 3526 2781 3533 2793
rect 3615 2792 3619 2796
rect 3605 2788 3619 2792
rect 3506 2727 3515 2739
rect 3482 2709 3495 2716
rect 3491 2704 3495 2709
rect 3511 2704 3515 2727
rect 3531 2704 3535 2781
rect 3605 2773 3609 2788
rect 3607 2761 3609 2773
rect 3605 2704 3609 2761
rect 3625 2739 3629 2796
rect 3655 2792 3659 2796
rect 3645 2788 3659 2792
rect 3665 2792 3669 2796
rect 3716 2792 3720 2796
rect 3665 2788 3679 2792
rect 3645 2739 3651 2788
rect 3674 2773 3679 2788
rect 3702 2784 3720 2792
rect 3702 2773 3706 2784
rect 3645 2727 3654 2739
rect 3625 2704 3629 2727
rect 3645 2704 3649 2727
rect 3674 2715 3680 2761
rect 3665 2711 3680 2715
rect 3702 2716 3706 2761
rect 3724 2739 3728 2796
rect 3746 2793 3750 2836
rect 3746 2781 3753 2793
rect 3835 2792 3839 2796
rect 3825 2788 3839 2792
rect 3726 2727 3735 2739
rect 3665 2704 3669 2711
rect 3702 2709 3715 2716
rect 3711 2704 3715 2709
rect 3731 2704 3735 2727
rect 3751 2704 3755 2781
rect 3825 2773 3829 2788
rect 3827 2761 3829 2773
rect 3825 2704 3829 2761
rect 3845 2739 3849 2796
rect 3875 2792 3879 2796
rect 3865 2788 3879 2792
rect 3885 2792 3889 2796
rect 3885 2788 3899 2792
rect 3865 2739 3871 2788
rect 3894 2773 3899 2788
rect 3865 2727 3874 2739
rect 3845 2704 3849 2727
rect 3865 2704 3869 2727
rect 3894 2715 3900 2761
rect 3885 2711 3900 2715
rect 3945 2753 3949 2836
rect 3991 2773 3995 2796
rect 3986 2761 3995 2773
rect 3999 2773 4003 2796
rect 4071 2773 4075 2796
rect 3999 2761 4014 2773
rect 4066 2761 4075 2773
rect 4079 2773 4083 2796
rect 4079 2761 4094 2773
rect 3945 2741 3954 2753
rect 3885 2704 3889 2711
rect 3945 2684 3949 2741
rect 3991 2684 3995 2761
rect 4011 2684 4015 2761
rect 4071 2684 4075 2761
rect 4091 2684 4095 2761
rect 4165 2739 4169 2796
rect 4185 2782 4189 2796
rect 4205 2782 4209 2796
rect 4256 2792 4260 2796
rect 4242 2784 4260 2792
rect 4185 2776 4200 2782
rect 4205 2776 4221 2782
rect 4194 2753 4200 2776
rect 4165 2727 4174 2739
rect 4172 2684 4176 2727
rect 4194 2704 4198 2741
rect 4214 2739 4221 2776
rect 4242 2773 4246 2784
rect 4214 2714 4221 2727
rect 4202 2708 4221 2714
rect 4242 2716 4246 2761
rect 4264 2739 4268 2796
rect 4286 2793 4290 2836
rect 4365 2793 4369 2836
rect 4385 2824 4389 2836
rect 4405 2828 4409 2836
rect 4405 2824 4420 2828
rect 4385 2820 4400 2824
rect 4394 2813 4400 2820
rect 4286 2781 4293 2793
rect 4365 2781 4373 2793
rect 4385 2781 4392 2793
rect 4266 2727 4275 2739
rect 4242 2709 4255 2716
rect 4202 2704 4206 2708
rect 4251 2704 4255 2709
rect 4271 2704 4275 2727
rect 4291 2704 4295 2781
rect 4388 2724 4392 2781
rect 4396 2724 4400 2801
rect 4414 2793 4420 2824
rect 4404 2781 4414 2793
rect 4404 2724 4408 2781
rect 4455 2753 4459 2796
rect 4475 2754 4479 2836
rect 4489 2777 4493 2836
rect 4509 2796 4513 2836
rect 4521 2830 4525 2836
rect 4515 2784 4518 2796
rect 4489 2769 4498 2777
rect 4455 2704 4459 2741
rect 4475 2684 4479 2742
rect 4494 2740 4498 2769
rect 4514 2720 4518 2784
rect 4485 2716 4518 2720
rect 4485 2684 4489 2716
rect 4523 2708 4527 2818
rect 4541 2810 4545 2836
rect 4587 2832 4591 2836
rect 4555 2830 4591 2832
rect 4567 2828 4591 2830
rect 4509 2696 4511 2708
rect 4507 2684 4511 2696
rect 4517 2696 4519 2708
rect 4517 2684 4521 2696
rect 4539 2684 4543 2798
rect 4555 2692 4559 2818
rect 4595 2804 4599 2836
rect 4615 2816 4619 2856
rect 4623 2833 4627 2856
rect 4623 2826 4631 2833
rect 4593 2709 4599 2804
rect 4627 2797 4631 2826
rect 4623 2791 4631 2797
rect 4623 2745 4627 2791
rect 4645 2784 4649 2796
rect 4647 2772 4649 2784
rect 4593 2705 4617 2709
rect 4579 2700 4597 2701
rect 4567 2696 4597 2700
rect 4555 2688 4589 2692
rect 4585 2684 4589 2688
rect 4593 2684 4597 2696
rect 4613 2684 4617 2705
rect 4623 2684 4627 2733
rect 4645 2704 4649 2772
rect 4691 2753 4695 2836
rect 4751 2773 4755 2796
rect 4746 2761 4755 2773
rect 4759 2773 4763 2796
rect 4836 2792 4840 2796
rect 4822 2784 4840 2792
rect 4822 2773 4826 2784
rect 4759 2761 4774 2773
rect 4686 2741 4695 2753
rect 4691 2684 4695 2741
rect 4751 2684 4755 2761
rect 4771 2684 4775 2761
rect 4822 2716 4826 2761
rect 4844 2739 4848 2796
rect 4866 2793 4870 2836
rect 4866 2781 4873 2793
rect 4846 2727 4855 2739
rect 4822 2709 4835 2716
rect 4831 2704 4835 2709
rect 4851 2704 4855 2727
rect 4871 2704 4875 2781
rect 4957 2773 4961 2796
rect 4946 2761 4961 2773
rect 4965 2773 4969 2796
rect 5035 2792 5039 2796
rect 5025 2788 5039 2792
rect 5025 2773 5029 2788
rect 4965 2761 4974 2773
rect 5027 2761 5029 2773
rect 4945 2684 4949 2761
rect 4965 2684 4969 2761
rect 5025 2704 5029 2761
rect 5045 2739 5049 2796
rect 5075 2792 5079 2796
rect 5065 2788 5079 2792
rect 5085 2792 5089 2796
rect 5085 2788 5099 2792
rect 5065 2739 5071 2788
rect 5094 2773 5099 2788
rect 5131 2782 5135 2796
rect 5151 2782 5155 2796
rect 5119 2776 5135 2782
rect 5140 2776 5155 2782
rect 5065 2727 5074 2739
rect 5045 2704 5049 2727
rect 5065 2704 5069 2727
rect 5094 2715 5100 2761
rect 5119 2739 5126 2776
rect 5140 2753 5146 2776
rect 5085 2711 5100 2715
rect 5119 2714 5126 2727
rect 5085 2704 5089 2711
rect 5119 2708 5138 2714
rect 5134 2704 5138 2708
rect 5142 2704 5146 2741
rect 5171 2739 5175 2796
rect 5231 2773 5235 2836
rect 5253 2790 5257 2796
rect 5316 2792 5320 2796
rect 5255 2778 5257 2790
rect 5302 2784 5320 2792
rect 5302 2773 5306 2784
rect 5226 2761 5235 2773
rect 5166 2727 5175 2739
rect 5164 2684 5168 2727
rect 5231 2684 5235 2761
rect 5255 2710 5257 2722
rect 5253 2704 5257 2710
rect 5302 2716 5306 2761
rect 5324 2739 5328 2796
rect 5346 2793 5350 2836
rect 5346 2781 5353 2793
rect 5435 2792 5439 2796
rect 5425 2788 5439 2792
rect 5326 2727 5335 2739
rect 5302 2709 5315 2716
rect 5311 2704 5315 2709
rect 5331 2704 5335 2727
rect 5351 2704 5355 2781
rect 5425 2773 5429 2788
rect 5427 2761 5429 2773
rect 5425 2704 5429 2761
rect 5445 2739 5449 2796
rect 5475 2792 5479 2796
rect 5465 2788 5479 2792
rect 5485 2792 5489 2796
rect 5485 2788 5499 2792
rect 5465 2739 5471 2788
rect 5494 2773 5499 2788
rect 5465 2727 5474 2739
rect 5445 2704 5449 2727
rect 5465 2704 5469 2727
rect 5494 2715 5500 2761
rect 5485 2711 5500 2715
rect 5545 2753 5549 2836
rect 5595 2753 5599 2796
rect 5615 2754 5619 2836
rect 5629 2777 5633 2836
rect 5649 2796 5653 2836
rect 5661 2830 5665 2836
rect 5655 2784 5658 2796
rect 5629 2769 5638 2777
rect 5545 2741 5554 2753
rect 5485 2704 5489 2711
rect 5545 2684 5549 2741
rect 5595 2704 5599 2741
rect 5615 2684 5619 2742
rect 5634 2740 5638 2769
rect 5654 2720 5658 2784
rect 5625 2716 5658 2720
rect 5625 2684 5629 2716
rect 5663 2708 5667 2818
rect 5681 2810 5685 2836
rect 5727 2832 5731 2836
rect 5695 2830 5731 2832
rect 5707 2828 5731 2830
rect 5649 2696 5651 2708
rect 5647 2684 5651 2696
rect 5657 2696 5659 2708
rect 5657 2684 5661 2696
rect 5679 2684 5683 2798
rect 5695 2692 5699 2818
rect 5735 2804 5739 2836
rect 5755 2816 5759 2856
rect 5763 2833 5767 2856
rect 5763 2826 5771 2833
rect 5733 2709 5739 2804
rect 5767 2797 5771 2826
rect 5763 2791 5771 2797
rect 5831 2868 5835 2876
rect 5851 2868 5855 2872
rect 5861 2868 5865 2876
rect 5831 2824 5835 2828
rect 5823 2820 5835 2824
rect 5763 2745 5767 2791
rect 5785 2784 5789 2796
rect 5787 2772 5789 2784
rect 5733 2705 5757 2709
rect 5719 2700 5737 2701
rect 5707 2696 5737 2700
rect 5695 2688 5729 2692
rect 5725 2684 5729 2688
rect 5733 2684 5737 2696
rect 5753 2684 5757 2705
rect 5763 2684 5767 2733
rect 5785 2704 5789 2772
rect 5823 2739 5827 2820
rect 5951 2868 5955 2876
rect 5971 2868 5975 2872
rect 5981 2868 5985 2876
rect 5951 2824 5955 2828
rect 5943 2820 5955 2824
rect 5851 2783 5855 2788
rect 5861 2784 5865 2788
rect 5842 2779 5855 2783
rect 5842 2773 5847 2779
rect 5881 2774 5885 2796
rect 5855 2770 5885 2774
rect 5891 2773 5895 2796
rect 5823 2701 5827 2727
rect 5841 2730 5846 2761
rect 5891 2761 5894 2773
rect 5841 2724 5855 2730
rect 5851 2712 5855 2724
rect 5861 2712 5865 2758
rect 5881 2712 5885 2716
rect 5891 2712 5895 2761
rect 5943 2739 5947 2820
rect 6071 2868 6075 2876
rect 6091 2868 6095 2872
rect 6101 2868 6105 2876
rect 6071 2824 6075 2828
rect 6063 2820 6075 2824
rect 5971 2783 5975 2788
rect 5981 2784 5985 2788
rect 5962 2779 5975 2783
rect 5962 2773 5967 2779
rect 6001 2774 6005 2796
rect 5975 2770 6005 2774
rect 6011 2773 6015 2796
rect 5823 2696 5835 2701
rect 5831 2692 5835 2696
rect 5943 2701 5947 2727
rect 5961 2730 5966 2761
rect 6011 2761 6014 2773
rect 5961 2724 5975 2730
rect 5971 2712 5975 2724
rect 5981 2712 5985 2758
rect 6001 2712 6005 2716
rect 6011 2712 6015 2761
rect 6063 2739 6067 2820
rect 6091 2783 6095 2788
rect 6101 2784 6105 2788
rect 6082 2779 6095 2783
rect 6082 2773 6087 2779
rect 6121 2774 6125 2796
rect 6095 2770 6125 2774
rect 6131 2773 6135 2796
rect 5943 2696 5955 2701
rect 5951 2692 5955 2696
rect 6063 2701 6067 2727
rect 6081 2730 6086 2761
rect 6131 2761 6134 2773
rect 6081 2724 6095 2730
rect 6091 2712 6095 2724
rect 6101 2712 6105 2758
rect 6121 2712 6125 2716
rect 6131 2712 6135 2761
rect 6201 2722 6205 2796
rect 6223 2759 6227 2836
rect 6245 2773 6249 2836
rect 6305 2792 6309 2796
rect 6325 2792 6329 2796
rect 6305 2788 6329 2792
rect 6245 2761 6254 2773
rect 6226 2747 6239 2759
rect 6063 2696 6075 2701
rect 6071 2692 6075 2696
rect 6201 2710 6213 2722
rect 6215 2704 6219 2710
rect 6235 2704 6239 2747
rect 6245 2704 6249 2761
rect 6325 2739 6329 2788
rect 6371 2773 6375 2836
rect 6366 2761 6375 2773
rect 6325 2727 6334 2739
rect 6325 2712 6329 2727
rect 6305 2708 6329 2712
rect 6305 2704 6309 2708
rect 6325 2704 6329 2708
rect 6371 2704 6375 2761
rect 6393 2759 6397 2836
rect 6493 2833 6497 2856
rect 6489 2826 6497 2833
rect 6489 2797 6493 2826
rect 6501 2816 6505 2856
rect 6521 2804 6525 2836
rect 6529 2832 6533 2836
rect 6529 2830 6565 2832
rect 6529 2828 6553 2830
rect 6381 2747 6394 2759
rect 6381 2704 6385 2747
rect 6415 2722 6419 2796
rect 6407 2710 6419 2722
rect 6471 2784 6475 2796
rect 6489 2791 6497 2797
rect 6471 2772 6473 2784
rect 6401 2704 6405 2710
rect 6471 2704 6475 2772
rect 6493 2745 6497 2791
rect 5831 2664 5835 2672
rect 5851 2668 5855 2672
rect 5861 2668 5865 2672
rect 5881 2664 5885 2672
rect 5891 2668 5895 2672
rect 31 2660 35 2664
rect 105 2660 109 2664
rect 125 2660 129 2664
rect 175 2660 179 2664
rect 195 2660 199 2664
rect 205 2660 209 2664
rect 227 2660 231 2664
rect 237 2660 241 2664
rect 259 2660 263 2664
rect 305 2660 309 2664
rect 313 2660 317 2664
rect 333 2660 337 2664
rect 343 2660 347 2664
rect 365 2660 369 2664
rect 411 2660 415 2664
rect 485 2660 489 2664
rect 505 2660 509 2664
rect 555 2660 559 2664
rect 575 2660 579 2664
rect 585 2660 589 2664
rect 607 2660 611 2664
rect 617 2660 621 2664
rect 639 2660 643 2664
rect 685 2660 689 2664
rect 693 2660 697 2664
rect 713 2660 717 2664
rect 723 2660 727 2664
rect 745 2660 749 2664
rect 803 2660 807 2664
rect 825 2660 829 2664
rect 871 2660 875 2664
rect 891 2660 895 2664
rect 953 2660 957 2664
rect 963 2660 967 2664
rect 1033 2660 1037 2664
rect 1043 2660 1047 2664
rect 1111 2660 1115 2664
rect 1174 2660 1178 2664
rect 1182 2660 1186 2664
rect 1202 2660 1206 2664
rect 1210 2660 1214 2664
rect 1312 2660 1316 2664
rect 1334 2660 1338 2664
rect 1342 2660 1346 2664
rect 1405 2660 1409 2664
rect 1465 2660 1469 2664
rect 1485 2660 1489 2664
rect 1505 2660 1509 2664
rect 1551 2660 1555 2664
rect 1571 2660 1575 2664
rect 1633 2660 1637 2664
rect 1643 2660 1647 2664
rect 1711 2660 1715 2664
rect 1731 2660 1735 2664
rect 1805 2660 1809 2664
rect 1825 2660 1829 2664
rect 1845 2660 1849 2664
rect 1891 2660 1895 2664
rect 1911 2660 1915 2664
rect 1931 2660 1935 2664
rect 1991 2660 1995 2664
rect 2011 2660 2015 2664
rect 2031 2660 2035 2664
rect 2112 2660 2116 2664
rect 2134 2660 2138 2664
rect 2142 2660 2146 2664
rect 2195 2660 2199 2664
rect 2215 2660 2219 2664
rect 2225 2660 2229 2664
rect 2247 2660 2251 2664
rect 2257 2660 2261 2664
rect 2279 2660 2283 2664
rect 2325 2660 2329 2664
rect 2333 2660 2337 2664
rect 2353 2660 2357 2664
rect 2363 2660 2367 2664
rect 2385 2660 2389 2664
rect 2433 2660 2437 2664
rect 2443 2660 2447 2664
rect 2511 2660 2515 2664
rect 2585 2660 2589 2664
rect 2635 2660 2639 2664
rect 2655 2660 2659 2664
rect 2665 2660 2669 2664
rect 2687 2660 2691 2664
rect 2697 2660 2701 2664
rect 2719 2660 2723 2664
rect 2765 2660 2769 2664
rect 2773 2660 2777 2664
rect 2793 2660 2797 2664
rect 2803 2660 2807 2664
rect 2825 2660 2829 2664
rect 2871 2660 2875 2664
rect 2891 2660 2895 2664
rect 2911 2660 2915 2664
rect 2992 2660 2996 2664
rect 3014 2660 3018 2664
rect 3022 2660 3026 2664
rect 3071 2660 3075 2664
rect 3093 2660 3097 2664
rect 3103 2660 3107 2664
rect 3123 2660 3127 2664
rect 3131 2660 3135 2664
rect 3177 2660 3181 2664
rect 3199 2660 3203 2664
rect 3209 2660 3213 2664
rect 3231 2660 3235 2664
rect 3241 2660 3245 2664
rect 3261 2660 3265 2664
rect 3311 2660 3315 2664
rect 3371 2660 3375 2664
rect 3391 2660 3395 2664
rect 3411 2660 3415 2664
rect 3431 2660 3435 2664
rect 3491 2660 3495 2664
rect 3511 2660 3515 2664
rect 3531 2660 3535 2664
rect 3605 2660 3609 2664
rect 3625 2660 3629 2664
rect 3645 2660 3649 2664
rect 3665 2660 3669 2664
rect 3711 2660 3715 2664
rect 3731 2660 3735 2664
rect 3751 2660 3755 2664
rect 3825 2660 3829 2664
rect 3845 2660 3849 2664
rect 3865 2660 3869 2664
rect 3885 2660 3889 2664
rect 3945 2660 3949 2664
rect 3991 2660 3995 2664
rect 4011 2660 4015 2664
rect 4071 2660 4075 2664
rect 4091 2660 4095 2664
rect 4172 2660 4176 2664
rect 4194 2660 4198 2664
rect 4202 2660 4206 2664
rect 4251 2660 4255 2664
rect 4271 2660 4275 2664
rect 4291 2660 4295 2664
rect 4388 2660 4392 2664
rect 4396 2660 4400 2664
rect 4404 2660 4408 2664
rect 4455 2660 4459 2664
rect 4475 2660 4479 2664
rect 4485 2660 4489 2664
rect 4507 2660 4511 2664
rect 4517 2660 4521 2664
rect 4539 2660 4543 2664
rect 4585 2660 4589 2664
rect 4593 2660 4597 2664
rect 4613 2660 4617 2664
rect 4623 2660 4627 2664
rect 4645 2660 4649 2664
rect 4691 2660 4695 2664
rect 4751 2660 4755 2664
rect 4771 2660 4775 2664
rect 4831 2660 4835 2664
rect 4851 2660 4855 2664
rect 4871 2660 4875 2664
rect 4945 2660 4949 2664
rect 4965 2660 4969 2664
rect 5025 2660 5029 2664
rect 5045 2660 5049 2664
rect 5065 2660 5069 2664
rect 5085 2660 5089 2664
rect 5134 2660 5138 2664
rect 5142 2660 5146 2664
rect 5164 2660 5168 2664
rect 5231 2660 5235 2664
rect 5253 2660 5257 2664
rect 5311 2660 5315 2664
rect 5331 2660 5335 2664
rect 5351 2660 5355 2664
rect 5425 2660 5429 2664
rect 5445 2660 5449 2664
rect 5465 2660 5469 2664
rect 5485 2660 5489 2664
rect 5545 2660 5549 2664
rect 5595 2660 5599 2664
rect 5615 2660 5619 2664
rect 5625 2660 5629 2664
rect 5647 2660 5651 2664
rect 5657 2660 5661 2664
rect 5679 2660 5683 2664
rect 5725 2660 5729 2664
rect 5733 2660 5737 2664
rect 5753 2660 5757 2664
rect 5763 2660 5767 2664
rect 5785 2660 5789 2664
rect 5831 2660 5885 2664
rect 5951 2664 5955 2672
rect 5971 2668 5975 2672
rect 5981 2668 5985 2672
rect 6001 2664 6005 2672
rect 6011 2668 6015 2672
rect 5951 2660 6005 2664
rect 6071 2664 6075 2672
rect 6091 2668 6095 2672
rect 6101 2668 6105 2672
rect 6121 2664 6125 2672
rect 6131 2668 6135 2672
rect 6493 2684 6497 2733
rect 6521 2709 6527 2804
rect 6503 2705 6527 2709
rect 6503 2684 6507 2705
rect 6523 2700 6541 2701
rect 6523 2696 6553 2700
rect 6523 2684 6527 2696
rect 6561 2692 6565 2818
rect 6575 2810 6579 2836
rect 6595 2830 6599 2836
rect 6531 2688 6565 2692
rect 6531 2684 6535 2688
rect 6577 2684 6581 2798
rect 6593 2708 6597 2818
rect 6607 2796 6611 2836
rect 6602 2784 6605 2796
rect 6602 2720 6606 2784
rect 6627 2777 6631 2836
rect 6622 2769 6631 2777
rect 6622 2740 6626 2769
rect 6641 2754 6645 2836
rect 6661 2753 6665 2796
rect 6602 2716 6635 2720
rect 6601 2696 6603 2708
rect 6599 2684 6603 2696
rect 6609 2696 6611 2708
rect 6609 2684 6613 2696
rect 6631 2684 6635 2716
rect 6641 2684 6645 2742
rect 6661 2704 6665 2741
rect 6071 2660 6125 2664
rect 6215 2660 6219 2664
rect 6235 2660 6239 2664
rect 6245 2660 6249 2664
rect 6305 2660 6309 2664
rect 6325 2660 6329 2664
rect 6371 2660 6375 2664
rect 6381 2660 6385 2664
rect 6401 2660 6405 2664
rect 6471 2660 6475 2664
rect 6493 2660 6497 2664
rect 6503 2660 6507 2664
rect 6523 2660 6527 2664
rect 6531 2660 6535 2664
rect 6577 2660 6581 2664
rect 6599 2660 6603 2664
rect 6609 2660 6613 2664
rect 6631 2660 6635 2664
rect 6641 2660 6645 2664
rect 6661 2660 6665 2664
rect 31 2636 35 2640
rect 53 2636 57 2640
rect 63 2636 67 2640
rect 83 2636 87 2640
rect 91 2636 95 2640
rect 137 2636 141 2640
rect 159 2636 163 2640
rect 169 2636 173 2640
rect 191 2636 195 2640
rect 201 2636 205 2640
rect 221 2636 225 2640
rect 283 2636 287 2640
rect 305 2636 309 2640
rect 351 2636 355 2640
rect 373 2636 377 2640
rect 383 2636 387 2640
rect 403 2636 407 2640
rect 411 2636 415 2640
rect 457 2636 461 2640
rect 479 2636 483 2640
rect 489 2636 493 2640
rect 511 2636 515 2640
rect 521 2636 525 2640
rect 541 2636 545 2640
rect 612 2636 616 2640
rect 634 2636 638 2640
rect 642 2636 646 2640
rect 693 2636 697 2640
rect 703 2636 707 2640
rect 793 2636 797 2640
rect 803 2636 807 2640
rect 865 2636 869 2640
rect 885 2636 889 2640
rect 905 2636 909 2640
rect 925 2636 929 2640
rect 945 2636 949 2640
rect 965 2636 969 2640
rect 985 2636 989 2640
rect 1005 2636 1009 2640
rect 1051 2636 1055 2640
rect 1073 2636 1077 2640
rect 1083 2636 1087 2640
rect 1103 2636 1107 2640
rect 1111 2636 1115 2640
rect 1157 2636 1161 2640
rect 1179 2636 1183 2640
rect 1189 2636 1193 2640
rect 1211 2636 1215 2640
rect 1221 2636 1225 2640
rect 1241 2636 1245 2640
rect 1313 2636 1317 2640
rect 1323 2636 1327 2640
rect 1371 2636 1375 2640
rect 1391 2636 1395 2640
rect 1451 2636 1455 2640
rect 1525 2636 1529 2640
rect 1545 2636 1549 2640
rect 1565 2636 1569 2640
rect 1615 2636 1619 2640
rect 1635 2636 1639 2640
rect 1645 2636 1649 2640
rect 1667 2636 1671 2640
rect 1677 2636 1681 2640
rect 1699 2636 1703 2640
rect 1745 2636 1749 2640
rect 1753 2636 1757 2640
rect 1773 2636 1777 2640
rect 1783 2636 1787 2640
rect 1805 2636 1809 2640
rect 1851 2636 1855 2640
rect 1911 2636 1915 2640
rect 1971 2636 1975 2640
rect 1991 2636 1995 2640
rect 2011 2636 2015 2640
rect 2031 2636 2035 2640
rect 2091 2636 2095 2640
rect 2111 2636 2115 2640
rect 2171 2636 2225 2640
rect 31 2528 35 2596
rect 53 2567 57 2616
rect 63 2595 67 2616
rect 83 2604 87 2616
rect 91 2612 95 2616
rect 91 2608 125 2612
rect 83 2600 113 2604
rect 83 2599 101 2600
rect 63 2591 87 2595
rect 31 2516 33 2528
rect 31 2504 35 2516
rect 53 2509 57 2555
rect 49 2503 57 2509
rect 49 2474 53 2503
rect 81 2496 87 2591
rect 49 2467 57 2474
rect 53 2444 57 2467
rect 61 2444 65 2484
rect 81 2464 85 2496
rect 121 2482 125 2608
rect 137 2502 141 2616
rect 159 2604 163 2616
rect 161 2592 163 2604
rect 169 2604 173 2616
rect 169 2592 171 2604
rect 89 2470 113 2472
rect 89 2468 125 2470
rect 89 2464 93 2468
rect 135 2464 139 2490
rect 153 2482 157 2592
rect 191 2584 195 2616
rect 162 2580 195 2584
rect 162 2516 166 2580
rect 182 2531 186 2560
rect 201 2558 205 2616
rect 221 2559 225 2596
rect 283 2590 287 2596
rect 283 2578 285 2590
rect 182 2523 191 2531
rect 162 2504 165 2516
rect 155 2464 159 2470
rect 167 2464 171 2504
rect 187 2464 191 2523
rect 201 2464 205 2546
rect 221 2504 225 2547
rect 305 2539 309 2616
rect 305 2527 314 2539
rect 351 2528 355 2596
rect 373 2567 377 2616
rect 383 2595 387 2616
rect 403 2604 407 2616
rect 411 2612 415 2616
rect 411 2608 445 2612
rect 403 2600 433 2604
rect 403 2599 421 2600
rect 383 2591 407 2595
rect 283 2510 285 2522
rect 283 2504 287 2510
rect 305 2464 309 2527
rect 351 2516 353 2528
rect 351 2504 355 2516
rect 373 2509 377 2555
rect 369 2503 377 2509
rect 369 2474 373 2503
rect 401 2496 407 2591
rect 369 2467 377 2474
rect 373 2444 377 2467
rect 381 2444 385 2484
rect 401 2464 405 2496
rect 441 2482 445 2608
rect 457 2502 461 2616
rect 479 2604 483 2616
rect 481 2592 483 2604
rect 489 2604 493 2616
rect 489 2592 491 2604
rect 409 2470 433 2472
rect 409 2468 445 2470
rect 409 2464 413 2468
rect 455 2464 459 2490
rect 473 2482 477 2592
rect 511 2584 515 2616
rect 482 2580 515 2584
rect 482 2516 486 2580
rect 502 2531 506 2560
rect 521 2558 525 2616
rect 541 2559 545 2596
rect 612 2573 616 2616
rect 605 2561 614 2573
rect 502 2523 511 2531
rect 482 2504 485 2516
rect 475 2464 479 2470
rect 487 2464 491 2504
rect 507 2464 511 2523
rect 521 2464 525 2546
rect 541 2504 545 2547
rect 605 2504 609 2561
rect 634 2559 638 2596
rect 642 2592 646 2596
rect 642 2586 661 2592
rect 654 2573 661 2586
rect 693 2576 697 2596
rect 689 2569 697 2576
rect 703 2576 707 2596
rect 793 2576 797 2596
rect 703 2569 717 2576
rect 634 2524 640 2547
rect 654 2524 661 2561
rect 689 2553 695 2569
rect 686 2541 695 2553
rect 625 2518 640 2524
rect 645 2518 661 2524
rect 625 2504 629 2518
rect 645 2504 649 2518
rect 691 2464 695 2541
rect 711 2553 717 2569
rect 783 2569 797 2576
rect 803 2576 807 2596
rect 865 2576 869 2596
rect 885 2576 889 2596
rect 905 2576 909 2596
rect 925 2576 929 2596
rect 945 2576 949 2596
rect 965 2576 969 2596
rect 803 2569 811 2576
rect 783 2553 789 2569
rect 711 2541 714 2553
rect 786 2541 789 2553
rect 711 2464 715 2541
rect 785 2464 789 2541
rect 805 2553 811 2569
rect 865 2564 878 2576
rect 905 2564 918 2576
rect 945 2564 958 2576
rect 985 2573 989 2596
rect 1005 2573 1009 2596
rect 805 2541 814 2553
rect 805 2464 809 2541
rect 865 2504 869 2564
rect 885 2504 889 2564
rect 905 2504 909 2564
rect 925 2504 929 2564
rect 945 2504 949 2564
rect 965 2504 969 2564
rect 985 2561 994 2573
rect 1006 2561 1009 2573
rect 985 2504 989 2561
rect 1005 2504 1009 2561
rect 1051 2528 1055 2596
rect 1073 2567 1077 2616
rect 1083 2595 1087 2616
rect 1103 2604 1107 2616
rect 1111 2612 1115 2616
rect 1111 2608 1145 2612
rect 1103 2600 1133 2604
rect 1103 2599 1121 2600
rect 1083 2591 1107 2595
rect 1051 2516 1053 2528
rect 1051 2504 1055 2516
rect 1073 2509 1077 2555
rect 1069 2503 1077 2509
rect 1069 2474 1073 2503
rect 1101 2496 1107 2591
rect 1069 2467 1077 2474
rect 1073 2444 1077 2467
rect 1081 2444 1085 2484
rect 1101 2464 1105 2496
rect 1141 2482 1145 2608
rect 1157 2502 1161 2616
rect 1179 2604 1183 2616
rect 1181 2592 1183 2604
rect 1189 2604 1193 2616
rect 1189 2592 1191 2604
rect 1109 2470 1133 2472
rect 1109 2468 1145 2470
rect 1109 2464 1113 2468
rect 1155 2464 1159 2490
rect 1173 2482 1177 2592
rect 1211 2584 1215 2616
rect 1182 2580 1215 2584
rect 1182 2516 1186 2580
rect 1202 2531 1206 2560
rect 1221 2558 1225 2616
rect 1241 2559 1245 2596
rect 1313 2576 1317 2596
rect 1303 2569 1317 2576
rect 1323 2576 1327 2596
rect 1323 2569 1331 2576
rect 1303 2553 1309 2569
rect 1202 2523 1211 2531
rect 1182 2504 1185 2516
rect 1175 2464 1179 2470
rect 1187 2464 1191 2504
rect 1207 2464 1211 2523
rect 1221 2464 1225 2546
rect 1241 2504 1245 2547
rect 1306 2541 1309 2553
rect 1305 2464 1309 2541
rect 1325 2553 1331 2569
rect 1325 2541 1334 2553
rect 1325 2464 1329 2541
rect 1371 2539 1375 2616
rect 1391 2539 1395 2616
rect 1451 2559 1455 2616
rect 1446 2547 1455 2559
rect 1366 2527 1375 2539
rect 1371 2504 1375 2527
rect 1379 2527 1394 2539
rect 1379 2504 1383 2527
rect 1451 2464 1455 2547
rect 1525 2519 1529 2596
rect 1545 2573 1549 2596
rect 1565 2591 1569 2596
rect 1565 2584 1578 2591
rect 1545 2561 1554 2573
rect 1527 2507 1534 2519
rect 1530 2464 1534 2507
rect 1552 2504 1556 2561
rect 1574 2539 1578 2584
rect 1615 2559 1619 2596
rect 1635 2558 1639 2616
rect 1645 2584 1649 2616
rect 1667 2604 1671 2616
rect 1669 2592 1671 2604
rect 1677 2604 1681 2616
rect 1677 2592 1679 2604
rect 1645 2580 1678 2584
rect 1574 2516 1578 2527
rect 1560 2508 1578 2516
rect 1560 2504 1564 2508
rect 1615 2504 1619 2547
rect 1635 2464 1639 2546
rect 1654 2531 1658 2560
rect 1649 2523 1658 2531
rect 1649 2464 1653 2523
rect 1674 2516 1678 2580
rect 1675 2504 1678 2516
rect 1669 2464 1673 2504
rect 1683 2482 1687 2592
rect 1699 2502 1703 2616
rect 1745 2612 1749 2616
rect 1715 2608 1749 2612
rect 1681 2464 1685 2470
rect 1701 2464 1705 2490
rect 1715 2482 1719 2608
rect 1753 2604 1757 2616
rect 1727 2600 1757 2604
rect 1739 2599 1757 2600
rect 1773 2595 1777 2616
rect 1753 2591 1777 2595
rect 1753 2496 1759 2591
rect 1783 2567 1787 2616
rect 1783 2509 1787 2555
rect 1805 2528 1809 2596
rect 1851 2559 1855 2616
rect 1911 2559 1915 2616
rect 2171 2628 2175 2636
rect 2191 2628 2195 2632
rect 2201 2628 2205 2632
rect 2221 2628 2225 2636
rect 2291 2636 2345 2640
rect 2415 2636 2419 2640
rect 2435 2636 2439 2640
rect 2445 2636 2449 2640
rect 2467 2636 2471 2640
rect 2477 2636 2481 2640
rect 2499 2636 2503 2640
rect 2545 2636 2549 2640
rect 2553 2636 2557 2640
rect 2573 2636 2577 2640
rect 2583 2636 2587 2640
rect 2605 2636 2609 2640
rect 2651 2636 2705 2640
rect 2785 2636 2789 2640
rect 2805 2636 2809 2640
rect 2875 2636 2929 2640
rect 2985 2636 2989 2640
rect 3005 2636 3009 2640
rect 3025 2636 3029 2640
rect 3045 2636 3049 2640
rect 3105 2636 3109 2640
rect 3155 2636 3159 2640
rect 3175 2636 3179 2640
rect 3185 2636 3189 2640
rect 3207 2636 3211 2640
rect 3217 2636 3221 2640
rect 3239 2636 3243 2640
rect 3285 2636 3289 2640
rect 3293 2636 3297 2640
rect 3313 2636 3317 2640
rect 3323 2636 3327 2640
rect 3345 2636 3349 2640
rect 3391 2636 3395 2640
rect 3411 2636 3415 2640
rect 3493 2636 3497 2640
rect 3503 2636 3507 2640
rect 3551 2636 3555 2640
rect 3612 2636 3616 2640
rect 3620 2636 3624 2640
rect 3628 2636 3632 2640
rect 3712 2636 3716 2640
rect 3720 2636 3724 2640
rect 3728 2636 3732 2640
rect 3848 2636 3852 2640
rect 3856 2636 3860 2640
rect 3864 2636 3868 2640
rect 3911 2636 3915 2640
rect 3931 2636 3935 2640
rect 3951 2636 3955 2640
rect 4014 2636 4018 2640
rect 4022 2636 4026 2640
rect 4044 2636 4048 2640
rect 4125 2636 4129 2640
rect 4145 2636 4149 2640
rect 4205 2636 4209 2640
rect 4225 2636 4229 2640
rect 4245 2636 4249 2640
rect 4265 2636 4269 2640
rect 4315 2636 4319 2640
rect 4335 2636 4339 2640
rect 4345 2636 4349 2640
rect 4367 2636 4371 2640
rect 4377 2636 4381 2640
rect 4399 2636 4403 2640
rect 4445 2636 4449 2640
rect 4453 2636 4457 2640
rect 4473 2636 4477 2640
rect 4483 2636 4487 2640
rect 4505 2636 4509 2640
rect 4565 2636 4569 2640
rect 4625 2636 4629 2640
rect 4645 2636 4649 2640
rect 4665 2636 4669 2640
rect 4685 2636 4689 2640
rect 4731 2636 4785 2640
rect 4851 2636 4855 2640
rect 4873 2636 4877 2640
rect 4883 2636 4887 2640
rect 4903 2636 4907 2640
rect 4911 2636 4915 2640
rect 4957 2636 4961 2640
rect 4979 2636 4983 2640
rect 4989 2636 4993 2640
rect 5011 2636 5015 2640
rect 5021 2636 5025 2640
rect 5041 2636 5045 2640
rect 5091 2636 5095 2640
rect 5151 2636 5155 2640
rect 5171 2636 5175 2640
rect 5191 2636 5195 2640
rect 5211 2636 5215 2640
rect 5271 2636 5275 2640
rect 5291 2636 5295 2640
rect 5311 2636 5315 2640
rect 5371 2636 5375 2640
rect 5391 2636 5395 2640
rect 5465 2636 5469 2640
rect 5485 2636 5489 2640
rect 5531 2636 5535 2640
rect 5551 2636 5555 2640
rect 5571 2636 5575 2640
rect 5591 2636 5595 2640
rect 5611 2636 5615 2640
rect 5631 2636 5635 2640
rect 5651 2636 5655 2640
rect 5671 2636 5675 2640
rect 5745 2636 5749 2640
rect 5765 2636 5769 2640
rect 5811 2636 5815 2640
rect 5831 2636 5835 2640
rect 5851 2636 5855 2640
rect 5925 2636 5929 2640
rect 5945 2636 5949 2640
rect 5965 2636 5969 2640
rect 5985 2636 5989 2640
rect 6045 2636 6049 2640
rect 6091 2636 6095 2640
rect 6113 2636 6117 2640
rect 6123 2636 6127 2640
rect 6143 2636 6147 2640
rect 6151 2636 6155 2640
rect 6197 2636 6201 2640
rect 6219 2636 6223 2640
rect 6229 2636 6233 2640
rect 6251 2636 6255 2640
rect 6261 2636 6265 2640
rect 6281 2636 6285 2640
rect 6366 2636 6370 2640
rect 6374 2636 6378 2640
rect 6394 2636 6398 2640
rect 6402 2636 6406 2640
rect 6451 2636 6455 2640
rect 6471 2636 6475 2640
rect 6531 2636 6535 2640
rect 6594 2636 6598 2640
rect 6602 2636 6606 2640
rect 6622 2636 6626 2640
rect 6630 2636 6634 2640
rect 2231 2628 2235 2632
rect 2291 2628 2295 2636
rect 2311 2628 2315 2632
rect 2321 2628 2325 2632
rect 2341 2628 2345 2636
rect 2351 2628 2355 2632
rect 1971 2589 1975 2596
rect 1846 2547 1855 2559
rect 1906 2547 1915 2559
rect 1807 2516 1809 2528
rect 1783 2503 1791 2509
rect 1805 2504 1809 2516
rect 1727 2470 1751 2472
rect 1715 2468 1751 2470
rect 1747 2464 1751 2468
rect 1755 2464 1759 2496
rect 1775 2444 1779 2484
rect 1787 2474 1791 2503
rect 1783 2467 1791 2474
rect 1783 2444 1787 2467
rect 1851 2464 1855 2547
rect 1911 2464 1915 2547
rect 1960 2585 1975 2589
rect 1960 2539 1966 2585
rect 1991 2573 1995 2596
rect 2011 2573 2015 2596
rect 1986 2561 1995 2573
rect 1961 2512 1966 2527
rect 1989 2512 1995 2561
rect 1961 2508 1975 2512
rect 1971 2504 1975 2508
rect 1981 2508 1995 2512
rect 1981 2504 1985 2508
rect 2011 2504 2015 2561
rect 2031 2539 2035 2596
rect 2091 2539 2095 2616
rect 2111 2539 2115 2616
rect 2171 2604 2175 2608
rect 2163 2599 2175 2604
rect 2163 2573 2167 2599
rect 2291 2604 2295 2608
rect 2283 2599 2295 2604
rect 2191 2576 2195 2588
rect 2031 2527 2033 2539
rect 2086 2527 2095 2539
rect 2031 2512 2035 2527
rect 2021 2508 2035 2512
rect 2021 2504 2025 2508
rect 2091 2504 2095 2527
rect 2099 2527 2114 2539
rect 2099 2504 2103 2527
rect 2163 2480 2167 2561
rect 2181 2570 2195 2576
rect 2181 2539 2186 2570
rect 2201 2542 2205 2588
rect 2221 2584 2225 2588
rect 2182 2521 2187 2527
rect 2231 2539 2235 2588
rect 2283 2573 2287 2599
rect 2311 2576 2315 2588
rect 2195 2526 2225 2530
rect 2182 2517 2195 2521
rect 2191 2512 2195 2517
rect 2201 2512 2205 2516
rect 2163 2476 2175 2480
rect 2171 2472 2175 2476
rect 2221 2504 2225 2526
rect 2231 2527 2234 2539
rect 2231 2504 2235 2527
rect 2171 2424 2175 2432
rect 2191 2428 2195 2432
rect 2201 2424 2205 2432
rect 2283 2480 2287 2561
rect 2301 2570 2315 2576
rect 2301 2539 2306 2570
rect 2321 2542 2325 2588
rect 2341 2584 2345 2588
rect 2302 2521 2307 2527
rect 2351 2539 2355 2588
rect 2415 2559 2419 2596
rect 2435 2558 2439 2616
rect 2445 2584 2449 2616
rect 2467 2604 2471 2616
rect 2469 2592 2471 2604
rect 2477 2604 2481 2616
rect 2477 2592 2479 2604
rect 2445 2580 2478 2584
rect 2315 2526 2345 2530
rect 2302 2517 2315 2521
rect 2311 2512 2315 2517
rect 2321 2512 2325 2516
rect 2283 2476 2295 2480
rect 2291 2472 2295 2476
rect 2341 2504 2345 2526
rect 2351 2527 2354 2539
rect 2351 2504 2355 2527
rect 2415 2504 2419 2547
rect 2291 2424 2295 2432
rect 2311 2428 2315 2432
rect 2321 2424 2325 2432
rect 2435 2464 2439 2546
rect 2454 2531 2458 2560
rect 2449 2523 2458 2531
rect 2449 2464 2453 2523
rect 2474 2516 2478 2580
rect 2475 2504 2478 2516
rect 2469 2464 2473 2504
rect 2483 2482 2487 2592
rect 2499 2502 2503 2616
rect 2545 2612 2549 2616
rect 2515 2608 2549 2612
rect 2481 2464 2485 2470
rect 2501 2464 2505 2490
rect 2515 2482 2519 2608
rect 2553 2604 2557 2616
rect 2527 2600 2557 2604
rect 2539 2599 2557 2600
rect 2573 2595 2577 2616
rect 2553 2591 2577 2595
rect 2553 2496 2559 2591
rect 2583 2567 2587 2616
rect 2651 2628 2655 2636
rect 2671 2628 2675 2632
rect 2681 2628 2685 2632
rect 2701 2628 2705 2636
rect 2711 2628 2715 2632
rect 2651 2604 2655 2608
rect 2643 2599 2655 2604
rect 2583 2509 2587 2555
rect 2605 2528 2609 2596
rect 2643 2573 2647 2599
rect 2865 2628 2869 2632
rect 2875 2628 2879 2636
rect 2895 2628 2899 2632
rect 2905 2628 2909 2632
rect 2925 2628 2929 2636
rect 2671 2576 2675 2588
rect 2607 2516 2609 2528
rect 2583 2503 2591 2509
rect 2605 2504 2609 2516
rect 2527 2470 2551 2472
rect 2515 2468 2551 2470
rect 2547 2464 2551 2468
rect 2555 2464 2559 2496
rect 2575 2444 2579 2484
rect 2587 2474 2591 2503
rect 2583 2467 2591 2474
rect 2583 2444 2587 2467
rect 2643 2480 2647 2561
rect 2661 2570 2675 2576
rect 2661 2539 2666 2570
rect 2681 2542 2685 2588
rect 2701 2584 2705 2588
rect 2662 2521 2667 2527
rect 2711 2539 2715 2588
rect 2785 2539 2789 2616
rect 2805 2539 2809 2616
rect 2925 2604 2929 2608
rect 2925 2599 2937 2604
rect 2865 2539 2869 2588
rect 2875 2584 2879 2588
rect 2895 2542 2899 2588
rect 2905 2576 2909 2588
rect 2905 2570 2919 2576
rect 2675 2526 2705 2530
rect 2662 2517 2675 2521
rect 2671 2512 2675 2517
rect 2681 2512 2685 2516
rect 2643 2476 2655 2480
rect 2651 2472 2655 2476
rect 2701 2504 2705 2526
rect 2711 2527 2714 2539
rect 2786 2527 2801 2539
rect 2711 2504 2715 2527
rect 2797 2504 2801 2527
rect 2805 2527 2814 2539
rect 2866 2527 2869 2539
rect 2914 2539 2919 2570
rect 2933 2573 2937 2599
rect 2805 2504 2809 2527
rect 2865 2504 2869 2527
rect 2875 2526 2905 2530
rect 2875 2504 2879 2526
rect 2913 2521 2918 2527
rect 2905 2517 2918 2521
rect 2895 2512 2899 2516
rect 2905 2512 2909 2517
rect 2651 2424 2655 2432
rect 2671 2428 2675 2432
rect 2681 2424 2685 2432
rect 2933 2480 2937 2561
rect 2985 2539 2989 2596
rect 3005 2573 3009 2596
rect 3025 2573 3029 2596
rect 3045 2589 3049 2596
rect 3045 2585 3060 2589
rect 3025 2561 3034 2573
rect 2987 2527 2989 2539
rect 2985 2512 2989 2527
rect 2985 2508 2999 2512
rect 2995 2504 2999 2508
rect 3005 2504 3009 2561
rect 3025 2512 3031 2561
rect 3054 2539 3060 2585
rect 3105 2559 3109 2616
rect 3155 2559 3159 2596
rect 3105 2547 3114 2559
rect 3175 2558 3179 2616
rect 3185 2584 3189 2616
rect 3207 2604 3211 2616
rect 3209 2592 3211 2604
rect 3217 2604 3221 2616
rect 3217 2592 3219 2604
rect 3185 2580 3218 2584
rect 3054 2512 3059 2527
rect 3025 2508 3039 2512
rect 3035 2504 3039 2508
rect 3045 2508 3059 2512
rect 3045 2504 3049 2508
rect 2925 2476 2937 2480
rect 2925 2472 2929 2476
rect 2895 2424 2899 2432
rect 2905 2428 2909 2432
rect 2925 2424 2929 2432
rect 3105 2464 3109 2547
rect 3155 2504 3159 2547
rect 3175 2464 3179 2546
rect 3194 2531 3198 2560
rect 3189 2523 3198 2531
rect 3189 2464 3193 2523
rect 3214 2516 3218 2580
rect 3215 2504 3218 2516
rect 3209 2464 3213 2504
rect 3223 2482 3227 2592
rect 3239 2502 3243 2616
rect 3285 2612 3289 2616
rect 3255 2608 3289 2612
rect 3221 2464 3225 2470
rect 3241 2464 3245 2490
rect 3255 2482 3259 2608
rect 3293 2604 3297 2616
rect 3267 2600 3297 2604
rect 3279 2599 3297 2600
rect 3313 2595 3317 2616
rect 3293 2591 3317 2595
rect 3293 2496 3299 2591
rect 3323 2567 3327 2616
rect 3323 2509 3327 2555
rect 3345 2528 3349 2596
rect 3391 2539 3395 2616
rect 3411 2539 3415 2616
rect 3493 2576 3497 2596
rect 3483 2569 3497 2576
rect 3503 2576 3507 2596
rect 3503 2569 3511 2576
rect 3483 2553 3489 2569
rect 3486 2541 3489 2553
rect 3347 2516 3349 2528
rect 3386 2527 3395 2539
rect 3323 2503 3331 2509
rect 3345 2504 3349 2516
rect 3391 2504 3395 2527
rect 3399 2527 3414 2539
rect 3399 2504 3403 2527
rect 3267 2470 3291 2472
rect 3255 2468 3291 2470
rect 3287 2464 3291 2468
rect 3295 2464 3299 2496
rect 3315 2444 3319 2484
rect 3327 2474 3331 2503
rect 3323 2467 3331 2474
rect 3323 2444 3327 2467
rect 3485 2464 3489 2541
rect 3505 2553 3511 2569
rect 3551 2559 3555 2616
rect 3911 2591 3915 2596
rect 3902 2584 3915 2591
rect 3505 2541 3514 2553
rect 3546 2547 3555 2559
rect 3505 2464 3509 2541
rect 3551 2464 3555 2547
rect 3612 2519 3616 2576
rect 3606 2507 3616 2519
rect 3600 2476 3606 2507
rect 3620 2499 3624 2576
rect 3628 2519 3632 2576
rect 3712 2519 3716 2576
rect 3628 2507 3635 2519
rect 3647 2507 3655 2519
rect 3706 2507 3716 2519
rect 3620 2480 3626 2487
rect 3620 2476 3635 2480
rect 3600 2472 3615 2476
rect 3611 2464 3615 2472
rect 3631 2464 3635 2476
rect 3651 2464 3655 2507
rect 3700 2476 3706 2507
rect 3720 2499 3724 2576
rect 3728 2519 3732 2576
rect 3848 2519 3852 2576
rect 3728 2507 3735 2519
rect 3747 2507 3755 2519
rect 3720 2480 3726 2487
rect 3720 2476 3735 2480
rect 3700 2472 3715 2476
rect 3711 2464 3715 2472
rect 3731 2464 3735 2476
rect 3751 2464 3755 2507
rect 3825 2507 3833 2519
rect 3845 2507 3852 2519
rect 3825 2464 3829 2507
rect 3856 2499 3860 2576
rect 3864 2519 3868 2576
rect 3902 2539 3906 2584
rect 3931 2573 3935 2596
rect 3926 2561 3935 2573
rect 3864 2507 3874 2519
rect 3902 2516 3906 2527
rect 3902 2508 3920 2516
rect 3854 2480 3860 2487
rect 3845 2476 3860 2480
rect 3874 2476 3880 2507
rect 3916 2504 3920 2508
rect 3924 2504 3928 2561
rect 3951 2519 3955 2596
rect 4014 2592 4018 2596
rect 3999 2586 4018 2592
rect 3999 2573 4006 2586
rect 3999 2524 4006 2561
rect 4022 2559 4026 2596
rect 4044 2573 4048 2616
rect 4046 2561 4055 2573
rect 4020 2524 4026 2547
rect 3946 2507 3953 2519
rect 3999 2518 4015 2524
rect 4020 2518 4035 2524
rect 3845 2464 3849 2476
rect 3865 2472 3880 2476
rect 3865 2464 3869 2472
rect 3946 2464 3950 2507
rect 4011 2504 4015 2518
rect 4031 2504 4035 2518
rect 4051 2504 4055 2561
rect 4125 2539 4129 2616
rect 4145 2539 4149 2616
rect 4205 2539 4209 2596
rect 4225 2573 4229 2596
rect 4245 2573 4249 2596
rect 4265 2589 4269 2596
rect 4265 2585 4280 2589
rect 4245 2561 4254 2573
rect 4126 2527 4141 2539
rect 4137 2504 4141 2527
rect 4145 2527 4154 2539
rect 4207 2527 4209 2539
rect 4145 2504 4149 2527
rect 4205 2512 4209 2527
rect 4205 2508 4219 2512
rect 4215 2504 4219 2508
rect 4225 2504 4229 2561
rect 4245 2512 4251 2561
rect 4274 2539 4280 2585
rect 4315 2559 4319 2596
rect 4335 2558 4339 2616
rect 4345 2584 4349 2616
rect 4367 2604 4371 2616
rect 4369 2592 4371 2604
rect 4377 2604 4381 2616
rect 4377 2592 4379 2604
rect 4345 2580 4378 2584
rect 4274 2512 4279 2527
rect 4245 2508 4259 2512
rect 4255 2504 4259 2508
rect 4265 2508 4279 2512
rect 4265 2504 4269 2508
rect 4315 2504 4319 2547
rect 4335 2464 4339 2546
rect 4354 2531 4358 2560
rect 4349 2523 4358 2531
rect 4349 2464 4353 2523
rect 4374 2516 4378 2580
rect 4375 2504 4378 2516
rect 4369 2464 4373 2504
rect 4383 2482 4387 2592
rect 4399 2502 4403 2616
rect 4445 2612 4449 2616
rect 4415 2608 4449 2612
rect 4381 2464 4385 2470
rect 4401 2464 4405 2490
rect 4415 2482 4419 2608
rect 4453 2604 4457 2616
rect 4427 2600 4457 2604
rect 4439 2599 4457 2600
rect 4473 2595 4477 2616
rect 4453 2591 4477 2595
rect 4453 2496 4459 2591
rect 4483 2567 4487 2616
rect 4483 2509 4487 2555
rect 4505 2528 4509 2596
rect 4507 2516 4509 2528
rect 4483 2503 4491 2509
rect 4505 2504 4509 2516
rect 4565 2559 4569 2616
rect 4731 2628 4735 2636
rect 4751 2628 4755 2632
rect 4761 2628 4765 2632
rect 4781 2628 4785 2636
rect 4791 2628 4795 2632
rect 4731 2604 4735 2608
rect 4723 2599 4735 2604
rect 4565 2547 4574 2559
rect 4427 2470 4451 2472
rect 4415 2468 4451 2470
rect 4447 2464 4451 2468
rect 4455 2464 4459 2496
rect 4475 2444 4479 2484
rect 4487 2474 4491 2503
rect 4483 2467 4491 2474
rect 4483 2444 4487 2467
rect 4565 2464 4569 2547
rect 4625 2539 4629 2596
rect 4645 2573 4649 2596
rect 4665 2573 4669 2596
rect 4685 2589 4689 2596
rect 4685 2585 4700 2589
rect 4665 2561 4674 2573
rect 4627 2527 4629 2539
rect 4625 2512 4629 2527
rect 4625 2508 4639 2512
rect 4635 2504 4639 2508
rect 4645 2504 4649 2561
rect 4665 2512 4671 2561
rect 4694 2539 4700 2585
rect 4723 2573 4727 2599
rect 4751 2576 4755 2588
rect 4694 2512 4699 2527
rect 4665 2508 4679 2512
rect 4675 2504 4679 2508
rect 4685 2508 4699 2512
rect 4685 2504 4689 2508
rect 4723 2480 4727 2561
rect 4741 2570 4755 2576
rect 4741 2539 4746 2570
rect 4761 2542 4765 2588
rect 4781 2584 4785 2588
rect 4742 2521 4747 2527
rect 4791 2539 4795 2588
rect 4755 2526 4785 2530
rect 4742 2517 4755 2521
rect 4751 2512 4755 2517
rect 4761 2512 4765 2516
rect 4723 2476 4735 2480
rect 4731 2472 4735 2476
rect 4781 2504 4785 2526
rect 4791 2527 4794 2539
rect 4851 2528 4855 2596
rect 4873 2567 4877 2616
rect 4883 2595 4887 2616
rect 4903 2604 4907 2616
rect 4911 2612 4915 2616
rect 4911 2608 4945 2612
rect 4903 2600 4933 2604
rect 4903 2599 4921 2600
rect 4883 2591 4907 2595
rect 4791 2504 4795 2527
rect 4851 2516 4853 2528
rect 4851 2504 4855 2516
rect 4873 2509 4877 2555
rect 4731 2424 4735 2432
rect 4751 2428 4755 2432
rect 4761 2424 4765 2432
rect 4869 2503 4877 2509
rect 4869 2474 4873 2503
rect 4901 2496 4907 2591
rect 4869 2467 4877 2474
rect 4873 2444 4877 2467
rect 4881 2444 4885 2484
rect 4901 2464 4905 2496
rect 4941 2482 4945 2608
rect 4957 2502 4961 2616
rect 4979 2604 4983 2616
rect 4981 2592 4983 2604
rect 4989 2604 4993 2616
rect 4989 2592 4991 2604
rect 4909 2470 4933 2472
rect 4909 2468 4945 2470
rect 4909 2464 4913 2468
rect 4955 2464 4959 2490
rect 4973 2482 4977 2592
rect 5011 2584 5015 2616
rect 4982 2580 5015 2584
rect 4982 2516 4986 2580
rect 5002 2531 5006 2560
rect 5021 2558 5025 2616
rect 5041 2559 5045 2596
rect 5091 2559 5095 2616
rect 5151 2589 5155 2596
rect 5086 2547 5095 2559
rect 5002 2523 5011 2531
rect 4982 2504 4985 2516
rect 4975 2464 4979 2470
rect 4987 2464 4991 2504
rect 5007 2464 5011 2523
rect 5021 2464 5025 2546
rect 5041 2504 5045 2547
rect 5091 2464 5095 2547
rect 5140 2585 5155 2589
rect 5140 2539 5146 2585
rect 5171 2573 5175 2596
rect 5191 2573 5195 2596
rect 5166 2561 5175 2573
rect 5141 2512 5146 2527
rect 5169 2512 5175 2561
rect 5141 2508 5155 2512
rect 5151 2504 5155 2508
rect 5161 2508 5175 2512
rect 5161 2504 5165 2508
rect 5191 2504 5195 2561
rect 5211 2539 5215 2596
rect 5271 2591 5275 2596
rect 5262 2584 5275 2591
rect 5262 2539 5266 2584
rect 5291 2573 5295 2596
rect 5286 2561 5295 2573
rect 5211 2527 5213 2539
rect 5211 2512 5215 2527
rect 5201 2508 5215 2512
rect 5262 2516 5266 2527
rect 5262 2508 5280 2516
rect 5201 2504 5205 2508
rect 5276 2504 5280 2508
rect 5284 2504 5288 2561
rect 5311 2519 5315 2596
rect 5371 2539 5375 2616
rect 5391 2539 5395 2616
rect 5465 2539 5469 2616
rect 5485 2539 5489 2616
rect 5531 2573 5535 2596
rect 5551 2573 5555 2596
rect 5571 2576 5575 2596
rect 5591 2576 5595 2596
rect 5611 2576 5615 2596
rect 5631 2576 5635 2596
rect 5651 2576 5655 2596
rect 5671 2576 5675 2596
rect 5531 2561 5534 2573
rect 5546 2561 5555 2573
rect 5582 2564 5595 2576
rect 5622 2564 5635 2576
rect 5662 2564 5675 2576
rect 5366 2527 5375 2539
rect 5306 2507 5313 2519
rect 5306 2464 5310 2507
rect 5371 2504 5375 2527
rect 5379 2527 5394 2539
rect 5466 2527 5481 2539
rect 5379 2504 5383 2527
rect 5477 2504 5481 2527
rect 5485 2527 5494 2539
rect 5485 2504 5489 2527
rect 5531 2504 5535 2561
rect 5551 2504 5555 2561
rect 5571 2504 5575 2564
rect 5591 2504 5595 2564
rect 5611 2504 5615 2564
rect 5631 2504 5635 2564
rect 5651 2504 5655 2564
rect 5671 2504 5675 2564
rect 5745 2539 5749 2616
rect 5765 2539 5769 2616
rect 5811 2591 5815 2596
rect 5802 2584 5815 2591
rect 5802 2539 5806 2584
rect 5831 2573 5835 2596
rect 5826 2561 5835 2573
rect 5746 2527 5761 2539
rect 5757 2504 5761 2527
rect 5765 2527 5774 2539
rect 5765 2504 5769 2527
rect 5802 2516 5806 2527
rect 5802 2508 5820 2516
rect 5816 2504 5820 2508
rect 5824 2504 5828 2561
rect 5851 2519 5855 2596
rect 5925 2539 5929 2596
rect 5945 2573 5949 2596
rect 5965 2573 5969 2596
rect 5985 2589 5989 2596
rect 5985 2585 6000 2589
rect 5965 2561 5974 2573
rect 5927 2527 5929 2539
rect 5846 2507 5853 2519
rect 5925 2512 5929 2527
rect 5925 2508 5939 2512
rect 5846 2464 5850 2507
rect 5935 2504 5939 2508
rect 5945 2504 5949 2561
rect 5965 2512 5971 2561
rect 5994 2539 6000 2585
rect 6045 2559 6049 2616
rect 6045 2547 6054 2559
rect 5994 2512 5999 2527
rect 5965 2508 5979 2512
rect 5975 2504 5979 2508
rect 5985 2508 5999 2512
rect 5985 2504 5989 2508
rect 6045 2464 6049 2547
rect 6091 2528 6095 2596
rect 6113 2567 6117 2616
rect 6123 2595 6127 2616
rect 6143 2604 6147 2616
rect 6151 2612 6155 2616
rect 6151 2608 6185 2612
rect 6143 2600 6173 2604
rect 6143 2599 6161 2600
rect 6123 2591 6147 2595
rect 6091 2516 6093 2528
rect 6091 2504 6095 2516
rect 6113 2509 6117 2555
rect 6109 2503 6117 2509
rect 6109 2474 6113 2503
rect 6141 2496 6147 2591
rect 6109 2467 6117 2474
rect 6113 2444 6117 2467
rect 6121 2444 6125 2484
rect 6141 2464 6145 2496
rect 6181 2482 6185 2608
rect 6197 2502 6201 2616
rect 6219 2604 6223 2616
rect 6221 2592 6223 2604
rect 6229 2604 6233 2616
rect 6229 2592 6231 2604
rect 6149 2470 6173 2472
rect 6149 2468 6185 2470
rect 6149 2464 6153 2468
rect 6195 2464 6199 2490
rect 6213 2482 6217 2592
rect 6251 2584 6255 2616
rect 6222 2580 6255 2584
rect 6222 2516 6226 2580
rect 6242 2531 6246 2560
rect 6261 2558 6265 2616
rect 6281 2559 6285 2596
rect 6366 2591 6370 2596
rect 6340 2587 6370 2591
rect 6242 2523 6251 2531
rect 6222 2504 6225 2516
rect 6215 2464 6219 2470
rect 6227 2464 6231 2504
rect 6247 2464 6251 2523
rect 6261 2464 6265 2546
rect 6281 2504 6285 2547
rect 6340 2539 6346 2587
rect 6374 2582 6378 2596
rect 6365 2575 6378 2582
rect 6365 2573 6369 2575
rect 6394 2573 6398 2596
rect 6402 2588 6406 2596
rect 6451 2592 6455 2596
rect 6471 2592 6475 2596
rect 6451 2588 6475 2592
rect 6402 2581 6419 2588
rect 6367 2561 6369 2573
rect 6346 2527 6349 2539
rect 6345 2504 6349 2527
rect 6365 2504 6369 2561
rect 6394 2532 6398 2561
rect 6413 2539 6419 2581
rect 6451 2573 6455 2588
rect 6446 2561 6455 2573
rect 6385 2526 6398 2532
rect 6405 2527 6413 2532
rect 6405 2526 6425 2527
rect 6385 2504 6389 2526
rect 6405 2504 6409 2526
rect 6451 2512 6455 2561
rect 6531 2559 6535 2616
rect 6594 2588 6598 2596
rect 6526 2547 6535 2559
rect 6451 2508 6475 2512
rect 6451 2504 6455 2508
rect 6471 2504 6475 2508
rect 6531 2464 6535 2547
rect 6581 2581 6598 2588
rect 6581 2539 6587 2581
rect 6602 2573 6606 2596
rect 6622 2582 6626 2596
rect 6630 2591 6634 2596
rect 6630 2587 6660 2591
rect 6622 2575 6635 2582
rect 6631 2573 6635 2575
rect 6631 2561 6633 2573
rect 6602 2532 6606 2561
rect 6587 2527 6595 2532
rect 6575 2526 6595 2527
rect 6602 2526 6615 2532
rect 6591 2504 6595 2526
rect 6611 2504 6615 2526
rect 6631 2504 6635 2561
rect 6654 2539 6660 2587
rect 6651 2527 6654 2539
rect 6651 2504 6655 2527
rect 31 2420 35 2424
rect 53 2420 57 2424
rect 61 2420 65 2424
rect 81 2420 85 2424
rect 89 2420 93 2424
rect 135 2420 139 2424
rect 155 2420 159 2424
rect 167 2420 171 2424
rect 187 2420 191 2424
rect 201 2420 205 2424
rect 221 2420 225 2424
rect 283 2420 287 2424
rect 305 2420 309 2424
rect 351 2420 355 2424
rect 373 2420 377 2424
rect 381 2420 385 2424
rect 401 2420 405 2424
rect 409 2420 413 2424
rect 455 2420 459 2424
rect 475 2420 479 2424
rect 487 2420 491 2424
rect 507 2420 511 2424
rect 521 2420 525 2424
rect 541 2420 545 2424
rect 605 2420 609 2424
rect 625 2420 629 2424
rect 645 2420 649 2424
rect 691 2420 695 2424
rect 711 2420 715 2424
rect 785 2420 789 2424
rect 805 2420 809 2424
rect 865 2420 869 2424
rect 885 2420 889 2424
rect 905 2420 909 2424
rect 925 2420 929 2424
rect 945 2420 949 2424
rect 965 2420 969 2424
rect 985 2420 989 2424
rect 1005 2420 1009 2424
rect 1051 2420 1055 2424
rect 1073 2420 1077 2424
rect 1081 2420 1085 2424
rect 1101 2420 1105 2424
rect 1109 2420 1113 2424
rect 1155 2420 1159 2424
rect 1175 2420 1179 2424
rect 1187 2420 1191 2424
rect 1207 2420 1211 2424
rect 1221 2420 1225 2424
rect 1241 2420 1245 2424
rect 1305 2420 1309 2424
rect 1325 2420 1329 2424
rect 1371 2420 1375 2424
rect 1379 2420 1383 2424
rect 1451 2420 1455 2424
rect 1530 2420 1534 2424
rect 1552 2420 1556 2424
rect 1560 2420 1564 2424
rect 1615 2420 1619 2424
rect 1635 2420 1639 2424
rect 1649 2420 1653 2424
rect 1669 2420 1673 2424
rect 1681 2420 1685 2424
rect 1701 2420 1705 2424
rect 1747 2420 1751 2424
rect 1755 2420 1759 2424
rect 1775 2420 1779 2424
rect 1783 2420 1787 2424
rect 1805 2420 1809 2424
rect 1851 2420 1855 2424
rect 1911 2420 1915 2424
rect 1971 2420 1975 2424
rect 1981 2420 1985 2424
rect 2011 2420 2015 2424
rect 2021 2420 2025 2424
rect 2091 2420 2095 2424
rect 2099 2420 2103 2424
rect 2171 2420 2205 2424
rect 2221 2420 2225 2424
rect 2231 2420 2235 2424
rect 2291 2420 2325 2424
rect 2341 2420 2345 2424
rect 2351 2420 2355 2424
rect 2415 2420 2419 2424
rect 2435 2420 2439 2424
rect 2449 2420 2453 2424
rect 2469 2420 2473 2424
rect 2481 2420 2485 2424
rect 2501 2420 2505 2424
rect 2547 2420 2551 2424
rect 2555 2420 2559 2424
rect 2575 2420 2579 2424
rect 2583 2420 2587 2424
rect 2605 2420 2609 2424
rect 2651 2420 2685 2424
rect 2701 2420 2705 2424
rect 2711 2420 2715 2424
rect 2797 2420 2801 2424
rect 2805 2420 2809 2424
rect 2865 2420 2869 2424
rect 2875 2420 2879 2424
rect 2895 2420 2929 2424
rect 2995 2420 2999 2424
rect 3005 2420 3009 2424
rect 3035 2420 3039 2424
rect 3045 2420 3049 2424
rect 3105 2420 3109 2424
rect 3155 2420 3159 2424
rect 3175 2420 3179 2424
rect 3189 2420 3193 2424
rect 3209 2420 3213 2424
rect 3221 2420 3225 2424
rect 3241 2420 3245 2424
rect 3287 2420 3291 2424
rect 3295 2420 3299 2424
rect 3315 2420 3319 2424
rect 3323 2420 3327 2424
rect 3345 2420 3349 2424
rect 3391 2420 3395 2424
rect 3399 2420 3403 2424
rect 3485 2420 3489 2424
rect 3505 2420 3509 2424
rect 3551 2420 3555 2424
rect 3611 2420 3615 2424
rect 3631 2420 3635 2424
rect 3651 2420 3655 2424
rect 3711 2420 3715 2424
rect 3731 2420 3735 2424
rect 3751 2420 3755 2424
rect 3825 2420 3829 2424
rect 3845 2420 3849 2424
rect 3865 2420 3869 2424
rect 3916 2420 3920 2424
rect 3924 2420 3928 2424
rect 3946 2420 3950 2424
rect 4011 2420 4015 2424
rect 4031 2420 4035 2424
rect 4051 2420 4055 2424
rect 4137 2420 4141 2424
rect 4145 2420 4149 2424
rect 4215 2420 4219 2424
rect 4225 2420 4229 2424
rect 4255 2420 4259 2424
rect 4265 2420 4269 2424
rect 4315 2420 4319 2424
rect 4335 2420 4339 2424
rect 4349 2420 4353 2424
rect 4369 2420 4373 2424
rect 4381 2420 4385 2424
rect 4401 2420 4405 2424
rect 4447 2420 4451 2424
rect 4455 2420 4459 2424
rect 4475 2420 4479 2424
rect 4483 2420 4487 2424
rect 4505 2420 4509 2424
rect 4565 2420 4569 2424
rect 4635 2420 4639 2424
rect 4645 2420 4649 2424
rect 4675 2420 4679 2424
rect 4685 2420 4689 2424
rect 4731 2420 4765 2424
rect 4781 2420 4785 2424
rect 4791 2420 4795 2424
rect 4851 2420 4855 2424
rect 4873 2420 4877 2424
rect 4881 2420 4885 2424
rect 4901 2420 4905 2424
rect 4909 2420 4913 2424
rect 4955 2420 4959 2424
rect 4975 2420 4979 2424
rect 4987 2420 4991 2424
rect 5007 2420 5011 2424
rect 5021 2420 5025 2424
rect 5041 2420 5045 2424
rect 5091 2420 5095 2424
rect 5151 2420 5155 2424
rect 5161 2420 5165 2424
rect 5191 2420 5195 2424
rect 5201 2420 5205 2424
rect 5276 2420 5280 2424
rect 5284 2420 5288 2424
rect 5306 2420 5310 2424
rect 5371 2420 5375 2424
rect 5379 2420 5383 2424
rect 5477 2420 5481 2424
rect 5485 2420 5489 2424
rect 5531 2420 5535 2424
rect 5551 2420 5555 2424
rect 5571 2420 5575 2424
rect 5591 2420 5595 2424
rect 5611 2420 5615 2424
rect 5631 2420 5635 2424
rect 5651 2420 5655 2424
rect 5671 2420 5675 2424
rect 5757 2420 5761 2424
rect 5765 2420 5769 2424
rect 5816 2420 5820 2424
rect 5824 2420 5828 2424
rect 5846 2420 5850 2424
rect 5935 2420 5939 2424
rect 5945 2420 5949 2424
rect 5975 2420 5979 2424
rect 5985 2420 5989 2424
rect 6045 2420 6049 2424
rect 6091 2420 6095 2424
rect 6113 2420 6117 2424
rect 6121 2420 6125 2424
rect 6141 2420 6145 2424
rect 6149 2420 6153 2424
rect 6195 2420 6199 2424
rect 6215 2420 6219 2424
rect 6227 2420 6231 2424
rect 6247 2420 6251 2424
rect 6261 2420 6265 2424
rect 6281 2420 6285 2424
rect 6345 2420 6349 2424
rect 6365 2420 6369 2424
rect 6385 2420 6389 2424
rect 6405 2420 6409 2424
rect 6451 2420 6455 2424
rect 6471 2420 6475 2424
rect 6531 2420 6535 2424
rect 6591 2420 6595 2424
rect 6611 2420 6615 2424
rect 6631 2420 6635 2424
rect 6651 2420 6655 2424
rect 35 2396 39 2400
rect 55 2396 59 2400
rect 69 2396 73 2400
rect 89 2396 93 2400
rect 101 2396 105 2400
rect 121 2396 125 2400
rect 167 2396 171 2400
rect 175 2396 179 2400
rect 195 2396 199 2400
rect 203 2396 207 2400
rect 225 2396 229 2400
rect 283 2396 287 2400
rect 305 2396 309 2400
rect 365 2396 369 2400
rect 425 2396 429 2400
rect 497 2396 501 2400
rect 505 2396 509 2400
rect 556 2396 560 2400
rect 564 2396 568 2400
rect 586 2396 590 2400
rect 661 2396 665 2400
rect 683 2396 687 2400
rect 705 2396 709 2400
rect 751 2396 755 2400
rect 771 2396 775 2400
rect 791 2396 795 2400
rect 851 2396 855 2400
rect 871 2396 875 2400
rect 931 2396 935 2400
rect 953 2396 957 2400
rect 961 2396 965 2400
rect 981 2396 985 2400
rect 989 2396 993 2400
rect 1035 2396 1039 2400
rect 1055 2396 1059 2400
rect 1067 2396 1071 2400
rect 1087 2396 1091 2400
rect 1101 2396 1105 2400
rect 1121 2396 1125 2400
rect 1171 2396 1175 2400
rect 1235 2396 1239 2400
rect 1255 2396 1259 2400
rect 1269 2396 1273 2400
rect 1289 2396 1293 2400
rect 1301 2396 1305 2400
rect 1321 2396 1325 2400
rect 1367 2396 1371 2400
rect 1375 2396 1379 2400
rect 1395 2396 1399 2400
rect 1403 2396 1407 2400
rect 1425 2396 1429 2400
rect 1485 2396 1489 2400
rect 1531 2396 1535 2400
rect 1541 2396 1545 2400
rect 1571 2396 1575 2400
rect 1581 2396 1585 2400
rect 1656 2396 1660 2400
rect 1664 2396 1668 2400
rect 1686 2396 1690 2400
rect 1777 2396 1781 2400
rect 1785 2396 1789 2400
rect 1857 2396 1861 2400
rect 1865 2396 1869 2400
rect 1935 2396 1939 2400
rect 1945 2396 1949 2400
rect 1975 2396 1979 2400
rect 1985 2396 1989 2400
rect 2045 2396 2049 2400
rect 2095 2396 2099 2400
rect 2115 2396 2119 2400
rect 2129 2396 2133 2400
rect 2149 2396 2153 2400
rect 2161 2396 2165 2400
rect 2181 2396 2185 2400
rect 2227 2396 2231 2400
rect 2235 2396 2239 2400
rect 2255 2396 2259 2400
rect 2263 2396 2267 2400
rect 2285 2396 2289 2400
rect 2357 2396 2361 2400
rect 2365 2396 2369 2400
rect 2416 2396 2420 2400
rect 2424 2396 2428 2400
rect 2446 2396 2450 2400
rect 2525 2396 2529 2400
rect 2545 2396 2549 2400
rect 2565 2396 2569 2400
rect 2625 2396 2629 2400
rect 2645 2396 2649 2400
rect 2665 2396 2669 2400
rect 2716 2396 2720 2400
rect 2724 2396 2728 2400
rect 2746 2396 2750 2400
rect 2837 2396 2841 2400
rect 2845 2396 2849 2400
rect 2891 2396 2895 2400
rect 2913 2396 2917 2400
rect 2921 2396 2925 2400
rect 2941 2396 2945 2400
rect 2949 2396 2953 2400
rect 2995 2396 2999 2400
rect 3015 2396 3019 2400
rect 3027 2396 3031 2400
rect 3047 2396 3051 2400
rect 3061 2396 3065 2400
rect 3081 2396 3085 2400
rect 3136 2396 3140 2400
rect 3144 2396 3148 2400
rect 3166 2396 3170 2400
rect 3255 2396 3259 2400
rect 3265 2396 3269 2400
rect 3295 2396 3299 2400
rect 3305 2396 3309 2400
rect 3377 2396 3381 2400
rect 3385 2396 3389 2400
rect 3445 2396 3449 2400
rect 3517 2396 3521 2400
rect 3525 2396 3529 2400
rect 3575 2396 3579 2400
rect 3595 2396 3599 2400
rect 3609 2396 3613 2400
rect 3629 2396 3633 2400
rect 3641 2396 3645 2400
rect 3661 2396 3665 2400
rect 3707 2396 3711 2400
rect 3715 2396 3719 2400
rect 3735 2396 3739 2400
rect 3743 2396 3747 2400
rect 3765 2396 3769 2400
rect 3811 2396 3815 2400
rect 3831 2396 3835 2400
rect 3891 2396 3895 2400
rect 3911 2396 3915 2400
rect 3931 2396 3935 2400
rect 3991 2396 4025 2400
rect 4041 2396 4045 2400
rect 4051 2396 4055 2400
rect 4111 2396 4145 2400
rect 4161 2396 4165 2400
rect 4171 2396 4175 2400
rect 4231 2396 4265 2400
rect 4281 2396 4285 2400
rect 4291 2396 4295 2400
rect 4351 2396 4355 2400
rect 4373 2396 4377 2400
rect 4457 2396 4461 2400
rect 4465 2396 4469 2400
rect 4511 2396 4545 2400
rect 4561 2396 4565 2400
rect 4571 2396 4575 2400
rect 4645 2396 4649 2400
rect 4655 2396 4659 2400
rect 4675 2396 4709 2400
rect 35 2273 39 2316
rect 55 2274 59 2356
rect 69 2297 73 2356
rect 89 2316 93 2356
rect 101 2350 105 2356
rect 95 2304 98 2316
rect 69 2289 78 2297
rect 35 2224 39 2261
rect 55 2204 59 2262
rect 74 2260 78 2289
rect 94 2240 98 2304
rect 65 2236 98 2240
rect 65 2204 69 2236
rect 103 2228 107 2338
rect 121 2330 125 2356
rect 167 2352 171 2356
rect 135 2350 171 2352
rect 147 2348 171 2350
rect 89 2216 91 2228
rect 87 2204 91 2216
rect 97 2216 99 2228
rect 97 2204 101 2216
rect 119 2204 123 2318
rect 135 2212 139 2338
rect 175 2324 179 2356
rect 195 2336 199 2376
rect 203 2353 207 2376
rect 203 2346 211 2353
rect 173 2229 179 2324
rect 207 2317 211 2346
rect 203 2311 211 2317
rect 203 2265 207 2311
rect 225 2304 229 2316
rect 227 2292 229 2304
rect 283 2310 287 2316
rect 283 2298 285 2310
rect 173 2225 197 2229
rect 159 2220 177 2221
rect 147 2216 177 2220
rect 135 2208 169 2212
rect 165 2204 169 2208
rect 173 2204 177 2216
rect 193 2204 197 2225
rect 203 2204 207 2253
rect 225 2224 229 2292
rect 305 2293 309 2356
rect 305 2281 314 2293
rect 283 2230 285 2242
rect 283 2224 287 2230
rect 305 2204 309 2281
rect 365 2259 369 2316
rect 425 2273 429 2356
rect 497 2293 501 2316
rect 486 2281 501 2293
rect 505 2293 509 2316
rect 556 2312 560 2316
rect 542 2304 560 2312
rect 542 2293 546 2304
rect 505 2281 514 2293
rect 425 2261 434 2273
rect 365 2247 374 2259
rect 365 2224 369 2247
rect 425 2204 429 2261
rect 485 2204 489 2281
rect 505 2204 509 2281
rect 542 2236 546 2281
rect 564 2259 568 2316
rect 586 2313 590 2356
rect 586 2301 593 2313
rect 566 2247 575 2259
rect 542 2229 555 2236
rect 551 2224 555 2229
rect 571 2224 575 2247
rect 591 2224 595 2301
rect 661 2242 665 2316
rect 683 2279 687 2356
rect 705 2293 709 2356
rect 751 2348 755 2356
rect 740 2344 755 2348
rect 771 2344 775 2356
rect 740 2313 746 2344
rect 760 2340 775 2344
rect 760 2333 766 2340
rect 746 2301 756 2313
rect 705 2281 714 2293
rect 686 2267 699 2279
rect 661 2230 673 2242
rect 675 2224 679 2230
rect 695 2224 699 2267
rect 705 2224 709 2281
rect 752 2244 756 2301
rect 760 2244 764 2321
rect 791 2313 795 2356
rect 768 2301 775 2313
rect 787 2301 795 2313
rect 768 2244 772 2301
rect 851 2279 855 2356
rect 846 2267 855 2279
rect 849 2251 855 2267
rect 871 2279 875 2356
rect 953 2353 957 2376
rect 949 2346 957 2353
rect 949 2317 953 2346
rect 961 2336 965 2376
rect 981 2324 985 2356
rect 989 2352 993 2356
rect 989 2350 1025 2352
rect 989 2348 1013 2350
rect 931 2304 935 2316
rect 949 2311 957 2317
rect 931 2292 933 2304
rect 871 2267 874 2279
rect 871 2251 877 2267
rect 849 2244 857 2251
rect 853 2224 857 2244
rect 863 2244 877 2251
rect 863 2224 867 2244
rect 931 2224 935 2292
rect 953 2265 957 2311
rect 953 2204 957 2253
rect 981 2229 987 2324
rect 963 2225 987 2229
rect 963 2204 967 2225
rect 983 2220 1001 2221
rect 983 2216 1013 2220
rect 983 2204 987 2216
rect 1021 2212 1025 2338
rect 1035 2330 1039 2356
rect 1055 2350 1059 2356
rect 991 2208 1025 2212
rect 991 2204 995 2208
rect 1037 2204 1041 2318
rect 1053 2228 1057 2338
rect 1067 2316 1071 2356
rect 1062 2304 1065 2316
rect 1062 2240 1066 2304
rect 1087 2297 1091 2356
rect 1082 2289 1091 2297
rect 1082 2260 1086 2289
rect 1101 2274 1105 2356
rect 1121 2273 1125 2316
rect 1171 2273 1175 2356
rect 1235 2273 1239 2316
rect 1255 2274 1259 2356
rect 1269 2297 1273 2356
rect 1289 2316 1293 2356
rect 1301 2350 1305 2356
rect 1295 2304 1298 2316
rect 1269 2289 1278 2297
rect 1062 2236 1095 2240
rect 1061 2216 1063 2228
rect 1059 2204 1063 2216
rect 1069 2216 1071 2228
rect 1069 2204 1073 2216
rect 1091 2204 1095 2236
rect 1101 2204 1105 2262
rect 1166 2261 1175 2273
rect 1121 2224 1125 2261
rect 1171 2204 1175 2261
rect 1235 2224 1239 2261
rect 1255 2204 1259 2262
rect 1274 2260 1278 2289
rect 1294 2240 1298 2304
rect 1265 2236 1298 2240
rect 1265 2204 1269 2236
rect 1303 2228 1307 2338
rect 1321 2330 1325 2356
rect 1367 2352 1371 2356
rect 1335 2350 1371 2352
rect 1347 2348 1371 2350
rect 1289 2216 1291 2228
rect 1287 2204 1291 2216
rect 1297 2216 1299 2228
rect 1297 2204 1301 2216
rect 1319 2204 1323 2318
rect 1335 2212 1339 2338
rect 1375 2324 1379 2356
rect 1395 2336 1399 2376
rect 1403 2353 1407 2376
rect 1403 2346 1411 2353
rect 1373 2229 1379 2324
rect 1407 2317 1411 2346
rect 1403 2311 1411 2317
rect 1403 2265 1407 2311
rect 1425 2304 1429 2316
rect 1427 2292 1429 2304
rect 1373 2225 1397 2229
rect 1359 2220 1377 2221
rect 1347 2216 1377 2220
rect 1335 2208 1369 2212
rect 1365 2204 1369 2208
rect 1373 2204 1377 2216
rect 1393 2204 1397 2225
rect 1403 2204 1407 2253
rect 1425 2224 1429 2292
rect 1485 2273 1489 2356
rect 1531 2312 1535 2316
rect 1521 2308 1535 2312
rect 1541 2312 1545 2316
rect 1541 2308 1555 2312
rect 1521 2293 1526 2308
rect 1485 2261 1494 2273
rect 1485 2204 1489 2261
rect 1520 2235 1526 2281
rect 1549 2259 1555 2308
rect 1571 2259 1575 2316
rect 1581 2312 1585 2316
rect 1656 2312 1660 2316
rect 1581 2308 1595 2312
rect 1591 2293 1595 2308
rect 1642 2304 1660 2312
rect 1642 2293 1646 2304
rect 1591 2281 1593 2293
rect 1546 2247 1555 2259
rect 1520 2231 1535 2235
rect 1531 2224 1535 2231
rect 1551 2224 1555 2247
rect 1571 2224 1575 2247
rect 1591 2224 1595 2281
rect 1642 2236 1646 2281
rect 1664 2259 1668 2316
rect 1686 2313 1690 2356
rect 1686 2301 1693 2313
rect 1666 2247 1675 2259
rect 1642 2229 1655 2236
rect 1651 2224 1655 2229
rect 1671 2224 1675 2247
rect 1691 2224 1695 2301
rect 1777 2293 1781 2316
rect 1766 2281 1781 2293
rect 1785 2293 1789 2316
rect 1857 2293 1861 2316
rect 1785 2281 1794 2293
rect 1846 2281 1861 2293
rect 1865 2293 1869 2316
rect 1935 2312 1939 2316
rect 1925 2308 1939 2312
rect 1925 2293 1929 2308
rect 1865 2281 1874 2293
rect 1927 2281 1929 2293
rect 1765 2204 1769 2281
rect 1785 2204 1789 2281
rect 1845 2204 1849 2281
rect 1865 2204 1869 2281
rect 1925 2224 1929 2281
rect 1945 2259 1949 2316
rect 1975 2312 1979 2316
rect 1965 2308 1979 2312
rect 1985 2312 1989 2316
rect 1985 2308 1999 2312
rect 1965 2259 1971 2308
rect 1994 2293 1999 2308
rect 1965 2247 1974 2259
rect 1945 2224 1949 2247
rect 1965 2224 1969 2247
rect 1994 2235 2000 2281
rect 1985 2231 2000 2235
rect 2045 2273 2049 2356
rect 2095 2273 2099 2316
rect 2115 2274 2119 2356
rect 2129 2297 2133 2356
rect 2149 2316 2153 2356
rect 2161 2350 2165 2356
rect 2155 2304 2158 2316
rect 2129 2289 2138 2297
rect 2045 2261 2054 2273
rect 1985 2224 1989 2231
rect 2045 2204 2049 2261
rect 2095 2224 2099 2261
rect 2115 2204 2119 2262
rect 2134 2260 2138 2289
rect 2154 2240 2158 2304
rect 2125 2236 2158 2240
rect 2125 2204 2129 2236
rect 2163 2228 2167 2338
rect 2181 2330 2185 2356
rect 2227 2352 2231 2356
rect 2195 2350 2231 2352
rect 2207 2348 2231 2350
rect 2149 2216 2151 2228
rect 2147 2204 2151 2216
rect 2157 2216 2159 2228
rect 2157 2204 2161 2216
rect 2179 2204 2183 2318
rect 2195 2212 2199 2338
rect 2235 2324 2239 2356
rect 2255 2336 2259 2376
rect 2263 2353 2267 2376
rect 2263 2346 2271 2353
rect 2233 2229 2239 2324
rect 2267 2317 2271 2346
rect 2263 2311 2271 2317
rect 2263 2265 2267 2311
rect 2285 2304 2289 2316
rect 2287 2292 2289 2304
rect 2357 2293 2361 2316
rect 2233 2225 2257 2229
rect 2219 2220 2237 2221
rect 2207 2216 2237 2220
rect 2195 2208 2229 2212
rect 2225 2204 2229 2208
rect 2233 2204 2237 2216
rect 2253 2204 2257 2225
rect 2263 2204 2267 2253
rect 2285 2224 2289 2292
rect 2346 2281 2361 2293
rect 2365 2293 2369 2316
rect 2416 2312 2420 2316
rect 2402 2304 2420 2312
rect 2402 2293 2406 2304
rect 2365 2281 2374 2293
rect 2345 2204 2349 2281
rect 2365 2204 2369 2281
rect 2402 2236 2406 2281
rect 2424 2259 2428 2316
rect 2446 2313 2450 2356
rect 2525 2313 2529 2356
rect 2545 2344 2549 2356
rect 2565 2348 2569 2356
rect 2565 2344 2580 2348
rect 2545 2340 2560 2344
rect 2554 2333 2560 2340
rect 2446 2301 2453 2313
rect 2525 2301 2533 2313
rect 2545 2301 2552 2313
rect 2426 2247 2435 2259
rect 2402 2229 2415 2236
rect 2411 2224 2415 2229
rect 2431 2224 2435 2247
rect 2451 2224 2455 2301
rect 2548 2244 2552 2301
rect 2556 2244 2560 2321
rect 2574 2313 2580 2344
rect 2564 2301 2574 2313
rect 2564 2244 2568 2301
rect 2625 2259 2629 2316
rect 2645 2302 2649 2316
rect 2665 2302 2669 2316
rect 2716 2312 2720 2316
rect 2702 2304 2720 2312
rect 2645 2296 2660 2302
rect 2665 2296 2681 2302
rect 2654 2273 2660 2296
rect 2625 2247 2634 2259
rect 2632 2204 2636 2247
rect 2654 2224 2658 2261
rect 2674 2259 2681 2296
rect 2702 2293 2706 2304
rect 2674 2234 2681 2247
rect 2662 2228 2681 2234
rect 2702 2236 2706 2281
rect 2724 2259 2728 2316
rect 2746 2313 2750 2356
rect 2913 2353 2917 2376
rect 2909 2346 2917 2353
rect 2909 2317 2913 2346
rect 2921 2336 2925 2376
rect 2941 2324 2945 2356
rect 2949 2352 2953 2356
rect 2949 2350 2985 2352
rect 2949 2348 2973 2350
rect 2746 2301 2753 2313
rect 2726 2247 2735 2259
rect 2702 2229 2715 2236
rect 2662 2224 2666 2228
rect 2711 2224 2715 2229
rect 2731 2224 2735 2247
rect 2751 2224 2755 2301
rect 2837 2293 2841 2316
rect 2826 2281 2841 2293
rect 2845 2293 2849 2316
rect 2891 2304 2895 2316
rect 2909 2311 2917 2317
rect 2845 2281 2854 2293
rect 2891 2292 2893 2304
rect 2825 2204 2829 2281
rect 2845 2204 2849 2281
rect 2891 2224 2895 2292
rect 2913 2265 2917 2311
rect 2913 2204 2917 2253
rect 2941 2229 2947 2324
rect 2923 2225 2947 2229
rect 2923 2204 2927 2225
rect 2943 2220 2961 2221
rect 2943 2216 2973 2220
rect 2943 2204 2947 2216
rect 2981 2212 2985 2338
rect 2995 2330 2999 2356
rect 3015 2350 3019 2356
rect 2951 2208 2985 2212
rect 2951 2204 2955 2208
rect 2997 2204 3001 2318
rect 3013 2228 3017 2338
rect 3027 2316 3031 2356
rect 3022 2304 3025 2316
rect 3022 2240 3026 2304
rect 3047 2297 3051 2356
rect 3042 2289 3051 2297
rect 3042 2260 3046 2289
rect 3061 2274 3065 2356
rect 3081 2273 3085 2316
rect 3136 2312 3140 2316
rect 3122 2304 3140 2312
rect 3122 2293 3126 2304
rect 3022 2236 3055 2240
rect 3021 2216 3023 2228
rect 3019 2204 3023 2216
rect 3029 2216 3031 2228
rect 3029 2204 3033 2216
rect 3051 2204 3055 2236
rect 3061 2204 3065 2262
rect 3081 2224 3085 2261
rect 3122 2236 3126 2281
rect 3144 2259 3148 2316
rect 3166 2313 3170 2356
rect 3166 2301 3173 2313
rect 3255 2312 3259 2316
rect 3245 2308 3259 2312
rect 3146 2247 3155 2259
rect 3122 2229 3135 2236
rect 3131 2224 3135 2229
rect 3151 2224 3155 2247
rect 3171 2224 3175 2301
rect 3245 2293 3249 2308
rect 3247 2281 3249 2293
rect 3245 2224 3249 2281
rect 3265 2259 3269 2316
rect 3295 2312 3299 2316
rect 3285 2308 3299 2312
rect 3305 2312 3309 2316
rect 3305 2308 3319 2312
rect 3285 2259 3291 2308
rect 3314 2293 3319 2308
rect 3377 2293 3381 2316
rect 3366 2281 3381 2293
rect 3385 2293 3389 2316
rect 3385 2281 3394 2293
rect 3285 2247 3294 2259
rect 3265 2224 3269 2247
rect 3285 2224 3289 2247
rect 3314 2235 3320 2281
rect 3305 2231 3320 2235
rect 3305 2224 3309 2231
rect 3365 2204 3369 2281
rect 3385 2204 3389 2281
rect 3445 2273 3449 2356
rect 3517 2293 3521 2316
rect 3506 2281 3521 2293
rect 3525 2293 3529 2316
rect 3525 2281 3534 2293
rect 3445 2261 3454 2273
rect 3445 2204 3449 2261
rect 3505 2204 3509 2281
rect 3525 2204 3529 2281
rect 3575 2273 3579 2316
rect 3595 2274 3599 2356
rect 3609 2297 3613 2356
rect 3629 2316 3633 2356
rect 3641 2350 3645 2356
rect 3635 2304 3638 2316
rect 3609 2289 3618 2297
rect 3575 2224 3579 2261
rect 3595 2204 3599 2262
rect 3614 2260 3618 2289
rect 3634 2240 3638 2304
rect 3605 2236 3638 2240
rect 3605 2204 3609 2236
rect 3643 2228 3647 2338
rect 3661 2330 3665 2356
rect 3707 2352 3711 2356
rect 3675 2350 3711 2352
rect 3687 2348 3711 2350
rect 3629 2216 3631 2228
rect 3627 2204 3631 2216
rect 3637 2216 3639 2228
rect 3637 2204 3641 2216
rect 3659 2204 3663 2318
rect 3675 2212 3679 2338
rect 3715 2324 3719 2356
rect 3735 2336 3739 2376
rect 3743 2353 3747 2376
rect 3743 2346 3751 2353
rect 3713 2229 3719 2324
rect 3747 2317 3751 2346
rect 3743 2311 3751 2317
rect 3991 2388 3995 2396
rect 4011 2388 4015 2392
rect 4021 2388 4025 2396
rect 3743 2265 3747 2311
rect 3765 2304 3769 2316
rect 3767 2292 3769 2304
rect 3713 2225 3737 2229
rect 3699 2220 3717 2221
rect 3687 2216 3717 2220
rect 3675 2208 3709 2212
rect 3705 2204 3709 2208
rect 3713 2204 3717 2216
rect 3733 2204 3737 2225
rect 3743 2204 3747 2253
rect 3765 2224 3769 2292
rect 3811 2279 3815 2356
rect 3806 2267 3815 2279
rect 3809 2251 3815 2267
rect 3831 2279 3835 2356
rect 3891 2348 3895 2356
rect 3880 2344 3895 2348
rect 3911 2344 3915 2356
rect 3880 2313 3886 2344
rect 3900 2340 3915 2344
rect 3900 2333 3906 2340
rect 3886 2301 3896 2313
rect 3831 2267 3834 2279
rect 3831 2251 3837 2267
rect 3809 2244 3817 2251
rect 3813 2224 3817 2244
rect 3823 2244 3837 2251
rect 3892 2244 3896 2301
rect 3900 2244 3904 2321
rect 3931 2313 3935 2356
rect 3991 2344 3995 2348
rect 3908 2301 3915 2313
rect 3927 2301 3935 2313
rect 3983 2340 3995 2344
rect 3908 2244 3912 2301
rect 3983 2259 3987 2340
rect 4111 2388 4115 2396
rect 4131 2388 4135 2392
rect 4141 2388 4145 2396
rect 4111 2344 4115 2348
rect 4103 2340 4115 2344
rect 4011 2303 4015 2308
rect 4021 2304 4025 2308
rect 4002 2299 4015 2303
rect 4002 2293 4007 2299
rect 4041 2294 4045 2316
rect 4015 2290 4045 2294
rect 4051 2293 4055 2316
rect 3823 2224 3827 2244
rect 3983 2221 3987 2247
rect 4001 2250 4006 2281
rect 4051 2281 4054 2293
rect 4001 2244 4015 2250
rect 4011 2232 4015 2244
rect 4021 2232 4025 2278
rect 4041 2232 4045 2236
rect 4051 2232 4055 2281
rect 4103 2259 4107 2340
rect 4231 2388 4235 2396
rect 4251 2388 4255 2392
rect 4261 2388 4265 2396
rect 4231 2344 4235 2348
rect 4223 2340 4235 2344
rect 4131 2303 4135 2308
rect 4141 2304 4145 2308
rect 4122 2299 4135 2303
rect 4122 2293 4127 2299
rect 4161 2294 4165 2316
rect 4135 2290 4165 2294
rect 4171 2293 4175 2316
rect 3983 2216 3995 2221
rect 3991 2212 3995 2216
rect 4103 2221 4107 2247
rect 4121 2250 4126 2281
rect 4171 2281 4174 2293
rect 4121 2244 4135 2250
rect 4131 2232 4135 2244
rect 4141 2232 4145 2278
rect 4161 2232 4165 2236
rect 4171 2232 4175 2281
rect 4223 2259 4227 2340
rect 4251 2303 4255 2308
rect 4261 2304 4265 2308
rect 4242 2299 4255 2303
rect 4242 2293 4247 2299
rect 4281 2294 4285 2316
rect 4255 2290 4285 2294
rect 4291 2293 4295 2316
rect 4351 2293 4355 2356
rect 4511 2388 4515 2396
rect 4531 2388 4535 2392
rect 4541 2388 4545 2396
rect 4511 2344 4515 2348
rect 4503 2340 4515 2344
rect 4373 2310 4377 2316
rect 4375 2298 4377 2310
rect 4457 2293 4461 2316
rect 4103 2216 4115 2221
rect 4111 2212 4115 2216
rect 4223 2221 4227 2247
rect 4241 2250 4246 2281
rect 4291 2281 4294 2293
rect 4346 2281 4355 2293
rect 4446 2281 4461 2293
rect 4465 2293 4469 2316
rect 4465 2281 4474 2293
rect 4241 2244 4255 2250
rect 4251 2232 4255 2244
rect 4261 2232 4265 2278
rect 4281 2232 4285 2236
rect 4291 2232 4295 2281
rect 4223 2216 4235 2221
rect 4231 2212 4235 2216
rect 4351 2204 4355 2281
rect 4375 2230 4377 2242
rect 4373 2224 4377 2230
rect 3991 2184 3995 2192
rect 4011 2188 4015 2192
rect 4021 2188 4025 2192
rect 4041 2184 4045 2192
rect 4051 2188 4055 2192
rect 35 2180 39 2184
rect 55 2180 59 2184
rect 65 2180 69 2184
rect 87 2180 91 2184
rect 97 2180 101 2184
rect 119 2180 123 2184
rect 165 2180 169 2184
rect 173 2180 177 2184
rect 193 2180 197 2184
rect 203 2180 207 2184
rect 225 2180 229 2184
rect 283 2180 287 2184
rect 305 2180 309 2184
rect 365 2180 369 2184
rect 425 2180 429 2184
rect 485 2180 489 2184
rect 505 2180 509 2184
rect 551 2180 555 2184
rect 571 2180 575 2184
rect 591 2180 595 2184
rect 675 2180 679 2184
rect 695 2180 699 2184
rect 705 2180 709 2184
rect 752 2180 756 2184
rect 760 2180 764 2184
rect 768 2180 772 2184
rect 853 2180 857 2184
rect 863 2180 867 2184
rect 931 2180 935 2184
rect 953 2180 957 2184
rect 963 2180 967 2184
rect 983 2180 987 2184
rect 991 2180 995 2184
rect 1037 2180 1041 2184
rect 1059 2180 1063 2184
rect 1069 2180 1073 2184
rect 1091 2180 1095 2184
rect 1101 2180 1105 2184
rect 1121 2180 1125 2184
rect 1171 2180 1175 2184
rect 1235 2180 1239 2184
rect 1255 2180 1259 2184
rect 1265 2180 1269 2184
rect 1287 2180 1291 2184
rect 1297 2180 1301 2184
rect 1319 2180 1323 2184
rect 1365 2180 1369 2184
rect 1373 2180 1377 2184
rect 1393 2180 1397 2184
rect 1403 2180 1407 2184
rect 1425 2180 1429 2184
rect 1485 2180 1489 2184
rect 1531 2180 1535 2184
rect 1551 2180 1555 2184
rect 1571 2180 1575 2184
rect 1591 2180 1595 2184
rect 1651 2180 1655 2184
rect 1671 2180 1675 2184
rect 1691 2180 1695 2184
rect 1765 2180 1769 2184
rect 1785 2180 1789 2184
rect 1845 2180 1849 2184
rect 1865 2180 1869 2184
rect 1925 2180 1929 2184
rect 1945 2180 1949 2184
rect 1965 2180 1969 2184
rect 1985 2180 1989 2184
rect 2045 2180 2049 2184
rect 2095 2180 2099 2184
rect 2115 2180 2119 2184
rect 2125 2180 2129 2184
rect 2147 2180 2151 2184
rect 2157 2180 2161 2184
rect 2179 2180 2183 2184
rect 2225 2180 2229 2184
rect 2233 2180 2237 2184
rect 2253 2180 2257 2184
rect 2263 2180 2267 2184
rect 2285 2180 2289 2184
rect 2345 2180 2349 2184
rect 2365 2180 2369 2184
rect 2411 2180 2415 2184
rect 2431 2180 2435 2184
rect 2451 2180 2455 2184
rect 2548 2180 2552 2184
rect 2556 2180 2560 2184
rect 2564 2180 2568 2184
rect 2632 2180 2636 2184
rect 2654 2180 2658 2184
rect 2662 2180 2666 2184
rect 2711 2180 2715 2184
rect 2731 2180 2735 2184
rect 2751 2180 2755 2184
rect 2825 2180 2829 2184
rect 2845 2180 2849 2184
rect 2891 2180 2895 2184
rect 2913 2180 2917 2184
rect 2923 2180 2927 2184
rect 2943 2180 2947 2184
rect 2951 2180 2955 2184
rect 2997 2180 3001 2184
rect 3019 2180 3023 2184
rect 3029 2180 3033 2184
rect 3051 2180 3055 2184
rect 3061 2180 3065 2184
rect 3081 2180 3085 2184
rect 3131 2180 3135 2184
rect 3151 2180 3155 2184
rect 3171 2180 3175 2184
rect 3245 2180 3249 2184
rect 3265 2180 3269 2184
rect 3285 2180 3289 2184
rect 3305 2180 3309 2184
rect 3365 2180 3369 2184
rect 3385 2180 3389 2184
rect 3445 2180 3449 2184
rect 3505 2180 3509 2184
rect 3525 2180 3529 2184
rect 3575 2180 3579 2184
rect 3595 2180 3599 2184
rect 3605 2180 3609 2184
rect 3627 2180 3631 2184
rect 3637 2180 3641 2184
rect 3659 2180 3663 2184
rect 3705 2180 3709 2184
rect 3713 2180 3717 2184
rect 3733 2180 3737 2184
rect 3743 2180 3747 2184
rect 3765 2180 3769 2184
rect 3813 2180 3817 2184
rect 3823 2180 3827 2184
rect 3892 2180 3896 2184
rect 3900 2180 3904 2184
rect 3908 2180 3912 2184
rect 3991 2180 4045 2184
rect 4111 2184 4115 2192
rect 4131 2188 4135 2192
rect 4141 2188 4145 2192
rect 4161 2184 4165 2192
rect 4171 2188 4175 2192
rect 4111 2180 4165 2184
rect 4231 2184 4235 2192
rect 4251 2188 4255 2192
rect 4261 2188 4265 2192
rect 4281 2184 4285 2192
rect 4291 2188 4295 2192
rect 4445 2204 4449 2281
rect 4465 2204 4469 2281
rect 4503 2259 4507 2340
rect 4675 2388 4679 2396
rect 4685 2388 4689 2392
rect 4705 2388 4709 2396
rect 4751 2396 4785 2400
rect 4801 2396 4805 2400
rect 4811 2396 4815 2400
rect 4871 2396 4875 2400
rect 4879 2396 4883 2400
rect 4951 2396 4985 2400
rect 5001 2396 5005 2400
rect 5011 2396 5015 2400
rect 5085 2396 5089 2400
rect 5105 2396 5109 2400
rect 5125 2396 5129 2400
rect 5171 2396 5175 2400
rect 5231 2396 5235 2400
rect 5241 2396 5245 2400
rect 5271 2396 5275 2400
rect 5281 2396 5285 2400
rect 5365 2396 5369 2400
rect 5375 2396 5379 2400
rect 5395 2396 5429 2400
rect 4751 2388 4755 2396
rect 4771 2388 4775 2392
rect 4781 2388 4785 2396
rect 4531 2303 4535 2308
rect 4541 2304 4545 2308
rect 4522 2299 4535 2303
rect 4522 2293 4527 2299
rect 4561 2294 4565 2316
rect 4535 2290 4565 2294
rect 4571 2293 4575 2316
rect 4645 2293 4649 2316
rect 4503 2221 4507 2247
rect 4521 2250 4526 2281
rect 4571 2281 4574 2293
rect 4646 2281 4649 2293
rect 4655 2294 4659 2316
rect 4705 2344 4709 2348
rect 4751 2344 4755 2348
rect 4705 2340 4717 2344
rect 4675 2304 4679 2308
rect 4685 2303 4689 2308
rect 4685 2299 4698 2303
rect 4655 2290 4685 2294
rect 4521 2244 4535 2250
rect 4531 2232 4535 2244
rect 4541 2232 4545 2278
rect 4561 2232 4565 2236
rect 4571 2232 4575 2281
rect 4645 2232 4649 2281
rect 4693 2293 4698 2299
rect 4655 2232 4659 2236
rect 4675 2232 4679 2278
rect 4694 2250 4699 2281
rect 4685 2244 4699 2250
rect 4713 2259 4717 2340
rect 4743 2340 4755 2344
rect 4743 2259 4747 2340
rect 4951 2388 4955 2396
rect 4971 2388 4975 2392
rect 4981 2388 4985 2396
rect 4951 2344 4955 2348
rect 4943 2340 4955 2344
rect 4771 2303 4775 2308
rect 4781 2304 4785 2308
rect 4762 2299 4775 2303
rect 4762 2293 4767 2299
rect 4801 2294 4805 2316
rect 4775 2290 4805 2294
rect 4811 2293 4815 2316
rect 4871 2293 4875 2316
rect 4685 2232 4689 2244
rect 4503 2216 4515 2221
rect 4511 2212 4515 2216
rect 4713 2221 4717 2247
rect 4705 2216 4717 2221
rect 4743 2221 4747 2247
rect 4761 2250 4766 2281
rect 4811 2281 4814 2293
rect 4866 2281 4875 2293
rect 4879 2293 4883 2316
rect 4879 2281 4894 2293
rect 4761 2244 4775 2250
rect 4771 2232 4775 2244
rect 4781 2232 4785 2278
rect 4801 2232 4805 2236
rect 4811 2232 4815 2281
rect 4743 2216 4755 2221
rect 4705 2212 4709 2216
rect 4751 2212 4755 2216
rect 4871 2204 4875 2281
rect 4891 2204 4895 2281
rect 4943 2259 4947 2340
rect 4971 2303 4975 2308
rect 4981 2304 4985 2308
rect 4962 2299 4975 2303
rect 4962 2293 4967 2299
rect 5001 2294 5005 2316
rect 4975 2290 5005 2294
rect 5011 2293 5015 2316
rect 4943 2221 4947 2247
rect 4961 2250 4966 2281
rect 5011 2281 5014 2293
rect 4961 2244 4975 2250
rect 4971 2232 4975 2244
rect 4981 2232 4985 2278
rect 5001 2232 5005 2236
rect 5011 2232 5015 2281
rect 5085 2259 5089 2316
rect 5105 2302 5109 2316
rect 5125 2302 5129 2316
rect 5105 2296 5120 2302
rect 5125 2296 5141 2302
rect 5114 2273 5120 2296
rect 5085 2247 5094 2259
rect 4943 2216 4955 2221
rect 4951 2212 4955 2216
rect 4511 2184 4515 2192
rect 4531 2188 4535 2192
rect 4541 2188 4545 2192
rect 4561 2184 4565 2192
rect 4571 2188 4575 2192
rect 4645 2188 4649 2192
rect 4231 2180 4285 2184
rect 4351 2180 4355 2184
rect 4373 2180 4377 2184
rect 4445 2180 4449 2184
rect 4465 2180 4469 2184
rect 4511 2180 4565 2184
rect 4655 2184 4659 2192
rect 4675 2188 4679 2192
rect 4685 2188 4689 2192
rect 4705 2184 4709 2192
rect 4655 2180 4709 2184
rect 4751 2184 4755 2192
rect 4771 2188 4775 2192
rect 4781 2188 4785 2192
rect 4801 2184 4805 2192
rect 4811 2188 4815 2192
rect 5092 2204 5096 2247
rect 5114 2224 5118 2261
rect 5134 2259 5141 2296
rect 5171 2273 5175 2356
rect 5395 2388 5399 2396
rect 5405 2388 5409 2392
rect 5425 2388 5429 2396
rect 5471 2396 5505 2400
rect 5521 2396 5525 2400
rect 5531 2396 5535 2400
rect 5591 2396 5625 2400
rect 5641 2396 5645 2400
rect 5651 2396 5655 2400
rect 5725 2396 5729 2400
rect 5745 2396 5749 2400
rect 5765 2396 5769 2400
rect 5825 2396 5829 2400
rect 5845 2396 5849 2400
rect 5865 2396 5869 2400
rect 5925 2396 5929 2400
rect 5985 2396 5989 2400
rect 6005 2396 6009 2400
rect 6025 2396 6029 2400
rect 6045 2396 6049 2400
rect 6105 2396 6109 2400
rect 6115 2396 6119 2400
rect 6135 2396 6169 2400
rect 6225 2396 6229 2400
rect 6235 2396 6239 2400
rect 6255 2396 6289 2400
rect 6331 2396 6335 2400
rect 6396 2396 6400 2400
rect 6404 2396 6408 2400
rect 6426 2396 6430 2400
rect 6491 2396 6495 2400
rect 6511 2396 6515 2400
rect 6571 2396 6575 2400
rect 6591 2396 6595 2400
rect 6611 2396 6615 2400
rect 6671 2396 6675 2400
rect 5471 2388 5475 2396
rect 5491 2388 5495 2392
rect 5501 2388 5505 2396
rect 5231 2312 5235 2316
rect 5221 2308 5235 2312
rect 5241 2312 5245 2316
rect 5241 2308 5255 2312
rect 5221 2293 5226 2308
rect 5166 2261 5175 2273
rect 5134 2234 5141 2247
rect 5122 2228 5141 2234
rect 5122 2224 5126 2228
rect 4951 2184 4955 2192
rect 4971 2188 4975 2192
rect 4981 2188 4985 2192
rect 5001 2184 5005 2192
rect 5011 2188 5015 2192
rect 5171 2204 5175 2261
rect 5220 2235 5226 2281
rect 5249 2259 5255 2308
rect 5271 2259 5275 2316
rect 5281 2312 5285 2316
rect 5281 2308 5295 2312
rect 5291 2293 5295 2308
rect 5365 2293 5369 2316
rect 5291 2281 5293 2293
rect 5366 2281 5369 2293
rect 5375 2294 5379 2316
rect 5425 2344 5429 2348
rect 5471 2344 5475 2348
rect 5425 2340 5437 2344
rect 5395 2304 5399 2308
rect 5405 2303 5409 2308
rect 5405 2299 5418 2303
rect 5375 2290 5405 2294
rect 5246 2247 5255 2259
rect 5220 2231 5235 2235
rect 5231 2224 5235 2231
rect 5251 2224 5255 2247
rect 5271 2224 5275 2247
rect 5291 2224 5295 2281
rect 5365 2232 5369 2281
rect 5413 2293 5418 2299
rect 5375 2232 5379 2236
rect 5395 2232 5399 2278
rect 5414 2250 5419 2281
rect 5405 2244 5419 2250
rect 5433 2259 5437 2340
rect 5463 2340 5475 2344
rect 5463 2259 5467 2340
rect 5591 2388 5595 2396
rect 5611 2388 5615 2392
rect 5621 2388 5625 2396
rect 5591 2344 5595 2348
rect 5583 2340 5595 2344
rect 5491 2303 5495 2308
rect 5501 2304 5505 2308
rect 5482 2299 5495 2303
rect 5482 2293 5487 2299
rect 5521 2294 5525 2316
rect 5495 2290 5525 2294
rect 5531 2293 5535 2316
rect 5405 2232 5409 2244
rect 5433 2221 5437 2247
rect 5425 2216 5437 2221
rect 5463 2221 5467 2247
rect 5481 2250 5486 2281
rect 5531 2281 5534 2293
rect 5481 2244 5495 2250
rect 5491 2232 5495 2244
rect 5501 2232 5505 2278
rect 5521 2232 5525 2236
rect 5531 2232 5535 2281
rect 5583 2259 5587 2340
rect 5611 2303 5615 2308
rect 5621 2304 5625 2308
rect 5602 2299 5615 2303
rect 5602 2293 5607 2299
rect 5641 2294 5645 2316
rect 5615 2290 5645 2294
rect 5651 2293 5655 2316
rect 5725 2313 5729 2356
rect 5745 2344 5749 2356
rect 5765 2348 5769 2356
rect 5765 2344 5780 2348
rect 5745 2340 5760 2344
rect 5754 2333 5760 2340
rect 5725 2301 5733 2313
rect 5745 2301 5752 2313
rect 5463 2216 5475 2221
rect 5425 2212 5429 2216
rect 5471 2212 5475 2216
rect 5583 2221 5587 2247
rect 5601 2250 5606 2281
rect 5651 2281 5654 2293
rect 5601 2244 5615 2250
rect 5611 2232 5615 2244
rect 5621 2232 5625 2278
rect 5641 2232 5645 2236
rect 5651 2232 5655 2281
rect 5748 2244 5752 2301
rect 5756 2244 5760 2321
rect 5774 2313 5780 2344
rect 5825 2313 5829 2356
rect 5845 2344 5849 2356
rect 5865 2348 5869 2356
rect 5865 2344 5880 2348
rect 5845 2340 5860 2344
rect 5854 2333 5860 2340
rect 5764 2301 5774 2313
rect 5825 2301 5833 2313
rect 5845 2301 5852 2313
rect 5764 2244 5768 2301
rect 5848 2244 5852 2301
rect 5856 2244 5860 2321
rect 5874 2313 5880 2344
rect 5864 2301 5874 2313
rect 5864 2244 5868 2301
rect 5925 2273 5929 2356
rect 6135 2388 6139 2396
rect 6145 2388 6149 2392
rect 6165 2388 6169 2396
rect 5985 2293 5989 2316
rect 5986 2281 5989 2293
rect 5925 2261 5934 2273
rect 5583 2216 5595 2221
rect 5591 2212 5595 2216
rect 5365 2188 5369 2192
rect 5375 2184 5379 2192
rect 5395 2188 5399 2192
rect 5405 2188 5409 2192
rect 5425 2184 5429 2192
rect 4751 2180 4805 2184
rect 4871 2180 4875 2184
rect 4891 2180 4895 2184
rect 4951 2180 5005 2184
rect 5092 2180 5096 2184
rect 5114 2180 5118 2184
rect 5122 2180 5126 2184
rect 5171 2180 5175 2184
rect 5231 2180 5235 2184
rect 5251 2180 5255 2184
rect 5271 2180 5275 2184
rect 5291 2180 5295 2184
rect 5375 2180 5429 2184
rect 5471 2184 5475 2192
rect 5491 2188 5495 2192
rect 5501 2188 5505 2192
rect 5521 2184 5525 2192
rect 5531 2188 5535 2192
rect 5471 2180 5525 2184
rect 5591 2184 5595 2192
rect 5611 2188 5615 2192
rect 5621 2188 5625 2192
rect 5641 2184 5645 2192
rect 5651 2188 5655 2192
rect 5925 2204 5929 2261
rect 5980 2233 5986 2281
rect 6005 2259 6009 2316
rect 6025 2294 6029 2316
rect 6045 2294 6049 2316
rect 6025 2288 6038 2294
rect 6045 2293 6065 2294
rect 6105 2293 6109 2316
rect 6045 2288 6053 2293
rect 6034 2259 6038 2288
rect 6106 2281 6109 2293
rect 6115 2294 6119 2316
rect 6165 2344 6169 2348
rect 6165 2340 6177 2344
rect 6135 2304 6139 2308
rect 6145 2303 6149 2308
rect 6145 2299 6158 2303
rect 6115 2290 6145 2294
rect 6007 2247 6009 2259
rect 6005 2245 6009 2247
rect 6005 2238 6018 2245
rect 5980 2229 6010 2233
rect 6006 2224 6010 2229
rect 6014 2224 6018 2238
rect 6034 2224 6038 2247
rect 6053 2239 6059 2281
rect 6042 2232 6059 2239
rect 6105 2232 6109 2281
rect 6153 2293 6158 2299
rect 6115 2232 6119 2236
rect 6135 2232 6139 2278
rect 6154 2250 6159 2281
rect 6145 2244 6159 2250
rect 6173 2259 6177 2340
rect 6255 2388 6259 2396
rect 6265 2388 6269 2392
rect 6285 2388 6289 2396
rect 6225 2293 6229 2316
rect 6226 2281 6229 2293
rect 6235 2294 6239 2316
rect 6285 2344 6289 2348
rect 6285 2340 6297 2344
rect 6255 2304 6259 2308
rect 6265 2303 6269 2308
rect 6265 2299 6278 2303
rect 6235 2290 6265 2294
rect 6145 2232 6149 2244
rect 6042 2224 6046 2232
rect 6173 2221 6177 2247
rect 6225 2232 6229 2281
rect 6273 2293 6278 2299
rect 6235 2232 6239 2236
rect 6255 2232 6259 2278
rect 6274 2250 6279 2281
rect 6265 2244 6279 2250
rect 6293 2259 6297 2340
rect 6331 2273 6335 2356
rect 6396 2312 6400 2316
rect 6382 2304 6400 2312
rect 6382 2293 6386 2304
rect 6326 2261 6335 2273
rect 6265 2232 6269 2244
rect 6165 2216 6177 2221
rect 6165 2212 6169 2216
rect 6293 2221 6297 2247
rect 6285 2216 6297 2221
rect 6285 2212 6289 2216
rect 6331 2204 6335 2261
rect 6382 2236 6386 2281
rect 6404 2259 6408 2316
rect 6426 2313 6430 2356
rect 6426 2301 6433 2313
rect 6406 2247 6415 2259
rect 6382 2229 6395 2236
rect 6391 2224 6395 2229
rect 6411 2224 6415 2247
rect 6431 2224 6435 2301
rect 6491 2279 6495 2356
rect 6486 2267 6495 2279
rect 6489 2251 6495 2267
rect 6511 2279 6515 2356
rect 6571 2302 6575 2316
rect 6591 2302 6595 2316
rect 6559 2296 6575 2302
rect 6580 2296 6595 2302
rect 6511 2267 6514 2279
rect 6511 2251 6517 2267
rect 6559 2259 6566 2296
rect 6580 2273 6586 2296
rect 6489 2244 6497 2251
rect 6493 2224 6497 2244
rect 6503 2244 6517 2251
rect 6503 2224 6507 2244
rect 6559 2234 6566 2247
rect 6559 2228 6578 2234
rect 6574 2224 6578 2228
rect 6582 2224 6586 2261
rect 6611 2259 6615 2316
rect 6671 2273 6675 2356
rect 6666 2261 6675 2273
rect 6606 2247 6615 2259
rect 6105 2188 6109 2192
rect 6115 2184 6119 2192
rect 6135 2188 6139 2192
rect 6145 2188 6149 2192
rect 6165 2184 6169 2192
rect 6225 2188 6229 2192
rect 5591 2180 5645 2184
rect 5748 2180 5752 2184
rect 5756 2180 5760 2184
rect 5764 2180 5768 2184
rect 5848 2180 5852 2184
rect 5856 2180 5860 2184
rect 5864 2180 5868 2184
rect 5925 2180 5929 2184
rect 6006 2180 6010 2184
rect 6014 2180 6018 2184
rect 6034 2180 6038 2184
rect 6042 2180 6046 2184
rect 6115 2180 6169 2184
rect 6235 2184 6239 2192
rect 6255 2188 6259 2192
rect 6265 2188 6269 2192
rect 6285 2184 6289 2192
rect 6604 2204 6608 2247
rect 6671 2204 6675 2261
rect 6235 2180 6289 2184
rect 6331 2180 6335 2184
rect 6391 2180 6395 2184
rect 6411 2180 6415 2184
rect 6431 2180 6435 2184
rect 6493 2180 6497 2184
rect 6503 2180 6507 2184
rect 6574 2180 6578 2184
rect 6582 2180 6586 2184
rect 6604 2180 6608 2184
rect 6671 2180 6675 2184
rect 45 2156 49 2160
rect 65 2156 69 2160
rect 133 2156 137 2160
rect 143 2156 147 2160
rect 228 2156 232 2160
rect 236 2156 240 2160
rect 244 2156 248 2160
rect 328 2156 332 2160
rect 336 2156 340 2160
rect 344 2156 348 2160
rect 413 2156 417 2160
rect 423 2156 427 2160
rect 472 2156 476 2160
rect 480 2156 484 2160
rect 488 2156 492 2160
rect 585 2156 589 2160
rect 605 2156 609 2160
rect 651 2156 655 2160
rect 671 2156 675 2160
rect 691 2156 695 2160
rect 752 2156 756 2160
rect 760 2156 764 2160
rect 768 2156 772 2160
rect 851 2156 855 2160
rect 871 2156 875 2160
rect 953 2156 957 2160
rect 963 2156 967 2160
rect 1011 2156 1065 2160
rect 1135 2156 1139 2160
rect 1155 2156 1159 2160
rect 1165 2156 1169 2160
rect 1187 2156 1191 2160
rect 1197 2156 1201 2160
rect 1219 2156 1223 2160
rect 1265 2156 1269 2160
rect 1273 2156 1277 2160
rect 1293 2156 1297 2160
rect 1303 2156 1307 2160
rect 1325 2156 1329 2160
rect 1371 2156 1375 2160
rect 1431 2156 1435 2160
rect 1451 2156 1455 2160
rect 1471 2156 1475 2160
rect 1491 2156 1495 2160
rect 1565 2156 1569 2160
rect 1585 2156 1589 2160
rect 1605 2156 1609 2160
rect 1665 2156 1669 2160
rect 1685 2156 1689 2160
rect 1705 2156 1709 2160
rect 1765 2156 1769 2160
rect 1785 2156 1789 2160
rect 1845 2156 1849 2160
rect 1865 2156 1869 2160
rect 1885 2156 1889 2160
rect 1955 2156 2009 2160
rect 45 2059 49 2136
rect 65 2059 69 2136
rect 133 2096 137 2116
rect 123 2089 137 2096
rect 143 2096 147 2116
rect 413 2096 417 2116
rect 143 2089 151 2096
rect 123 2073 129 2089
rect 126 2061 129 2073
rect 46 2047 61 2059
rect 57 2024 61 2047
rect 65 2047 74 2059
rect 65 2024 69 2047
rect 125 1984 129 2061
rect 145 2073 151 2089
rect 145 2061 154 2073
rect 145 1984 149 2061
rect 228 2039 232 2096
rect 205 2027 213 2039
rect 225 2027 232 2039
rect 205 1984 209 2027
rect 236 2019 240 2096
rect 244 2039 248 2096
rect 328 2039 332 2096
rect 244 2027 254 2039
rect 305 2027 313 2039
rect 325 2027 332 2039
rect 234 2000 240 2007
rect 225 1996 240 2000
rect 254 1996 260 2027
rect 225 1984 229 1996
rect 245 1992 260 1996
rect 245 1984 249 1992
rect 305 1984 309 2027
rect 336 2019 340 2096
rect 344 2039 348 2096
rect 403 2089 417 2096
rect 423 2096 427 2116
rect 423 2089 431 2096
rect 403 2073 409 2089
rect 406 2061 409 2073
rect 344 2027 354 2039
rect 334 2000 340 2007
rect 325 1996 340 2000
rect 354 1996 360 2027
rect 325 1984 329 1996
rect 345 1992 360 1996
rect 345 1984 349 1992
rect 405 1984 409 2061
rect 425 2073 431 2089
rect 425 2061 434 2073
rect 425 1984 429 2061
rect 472 2039 476 2096
rect 466 2027 476 2039
rect 460 1996 466 2027
rect 480 2019 484 2096
rect 488 2039 492 2096
rect 585 2059 589 2136
rect 605 2059 609 2136
rect 651 2111 655 2116
rect 642 2104 655 2111
rect 642 2059 646 2104
rect 671 2093 675 2116
rect 666 2081 675 2093
rect 586 2047 601 2059
rect 488 2027 495 2039
rect 507 2027 515 2039
rect 480 2000 486 2007
rect 480 1996 495 2000
rect 460 1992 475 1996
rect 471 1984 475 1992
rect 491 1984 495 1996
rect 511 1984 515 2027
rect 597 2024 601 2047
rect 605 2047 614 2059
rect 605 2024 609 2047
rect 642 2036 646 2047
rect 642 2028 660 2036
rect 656 2024 660 2028
rect 664 2024 668 2081
rect 691 2039 695 2116
rect 752 2039 756 2096
rect 686 2027 693 2039
rect 746 2027 756 2039
rect 686 1984 690 2027
rect 740 1996 746 2027
rect 760 2019 764 2096
rect 768 2039 772 2096
rect 851 2059 855 2136
rect 871 2059 875 2136
rect 1011 2148 1015 2156
rect 1031 2148 1035 2152
rect 1041 2148 1045 2152
rect 1061 2148 1065 2156
rect 1071 2148 1075 2152
rect 1011 2124 1015 2128
rect 1003 2119 1015 2124
rect 953 2096 957 2116
rect 943 2089 957 2096
rect 963 2096 967 2116
rect 963 2089 971 2096
rect 1003 2093 1007 2119
rect 1031 2096 1035 2108
rect 943 2073 949 2089
rect 946 2061 949 2073
rect 846 2047 855 2059
rect 768 2027 775 2039
rect 787 2027 795 2039
rect 760 2000 766 2007
rect 760 1996 775 2000
rect 740 1992 755 1996
rect 751 1984 755 1992
rect 771 1984 775 1996
rect 791 1984 795 2027
rect 851 2024 855 2047
rect 859 2047 874 2059
rect 859 2024 863 2047
rect 945 1984 949 2061
rect 965 2073 971 2089
rect 965 2061 974 2073
rect 965 1984 969 2061
rect 1003 2000 1007 2081
rect 1021 2090 1035 2096
rect 1021 2059 1026 2090
rect 1041 2062 1045 2108
rect 1061 2104 1065 2108
rect 1022 2041 1027 2047
rect 1071 2059 1075 2108
rect 1135 2079 1139 2116
rect 1155 2078 1159 2136
rect 1165 2104 1169 2136
rect 1187 2124 1191 2136
rect 1189 2112 1191 2124
rect 1197 2124 1201 2136
rect 1197 2112 1199 2124
rect 1165 2100 1198 2104
rect 1035 2046 1065 2050
rect 1022 2037 1035 2041
rect 1031 2032 1035 2037
rect 1041 2032 1045 2036
rect 1003 1996 1015 2000
rect 1011 1992 1015 1996
rect 1061 2024 1065 2046
rect 1071 2047 1074 2059
rect 1071 2024 1075 2047
rect 1135 2024 1139 2067
rect 1011 1944 1015 1952
rect 1031 1948 1035 1952
rect 1041 1944 1045 1952
rect 1155 1984 1159 2066
rect 1174 2051 1178 2080
rect 1169 2043 1178 2051
rect 1169 1984 1173 2043
rect 1194 2036 1198 2100
rect 1195 2024 1198 2036
rect 1189 1984 1193 2024
rect 1203 2002 1207 2112
rect 1219 2022 1223 2136
rect 1265 2132 1269 2136
rect 1235 2128 1269 2132
rect 1201 1984 1205 1990
rect 1221 1984 1225 2010
rect 1235 2002 1239 2128
rect 1273 2124 1277 2136
rect 1247 2120 1277 2124
rect 1259 2119 1277 2120
rect 1293 2115 1297 2136
rect 1273 2111 1297 2115
rect 1273 2016 1279 2111
rect 1303 2087 1307 2136
rect 1303 2029 1307 2075
rect 1325 2048 1329 2116
rect 1371 2079 1375 2136
rect 1431 2109 1435 2116
rect 1366 2067 1375 2079
rect 1327 2036 1329 2048
rect 1303 2023 1311 2029
rect 1325 2024 1329 2036
rect 1247 1990 1271 1992
rect 1235 1988 1271 1990
rect 1267 1984 1271 1988
rect 1275 1984 1279 2016
rect 1295 1964 1299 2004
rect 1307 1994 1311 2023
rect 1303 1987 1311 1994
rect 1303 1964 1307 1987
rect 1371 1984 1375 2067
rect 1420 2105 1435 2109
rect 1420 2059 1426 2105
rect 1451 2093 1455 2116
rect 1471 2093 1475 2116
rect 1446 2081 1455 2093
rect 1421 2032 1426 2047
rect 1449 2032 1455 2081
rect 1421 2028 1435 2032
rect 1431 2024 1435 2028
rect 1441 2028 1455 2032
rect 1441 2024 1445 2028
rect 1471 2024 1475 2081
rect 1491 2059 1495 2116
rect 1491 2047 1493 2059
rect 1491 2032 1495 2047
rect 1565 2039 1569 2116
rect 1585 2093 1589 2116
rect 1605 2111 1609 2116
rect 1605 2104 1618 2111
rect 1585 2081 1594 2093
rect 1481 2028 1495 2032
rect 1481 2024 1485 2028
rect 1567 2027 1574 2039
rect 1570 1984 1574 2027
rect 1592 2024 1596 2081
rect 1614 2059 1618 2104
rect 1614 2036 1618 2047
rect 1665 2039 1669 2116
rect 1685 2093 1689 2116
rect 1705 2111 1709 2116
rect 1705 2104 1718 2111
rect 1685 2081 1694 2093
rect 1600 2028 1618 2036
rect 1600 2024 1604 2028
rect 1667 2027 1674 2039
rect 1670 1984 1674 2027
rect 1692 2024 1696 2081
rect 1714 2059 1718 2104
rect 1765 2059 1769 2136
rect 1785 2059 1789 2136
rect 1945 2148 1949 2152
rect 1955 2148 1959 2156
rect 1975 2148 1979 2152
rect 1985 2148 1989 2152
rect 2005 2148 2009 2156
rect 2075 2156 2129 2160
rect 2175 2156 2179 2160
rect 2195 2156 2199 2160
rect 2205 2156 2209 2160
rect 2227 2156 2231 2160
rect 2237 2156 2241 2160
rect 2259 2156 2263 2160
rect 2305 2156 2309 2160
rect 2313 2156 2317 2160
rect 2333 2156 2337 2160
rect 2343 2156 2347 2160
rect 2365 2156 2369 2160
rect 2425 2156 2429 2160
rect 2445 2156 2449 2160
rect 2465 2156 2469 2160
rect 2511 2156 2515 2160
rect 2531 2156 2535 2160
rect 2628 2156 2632 2160
rect 2636 2156 2640 2160
rect 2644 2156 2648 2160
rect 2691 2156 2745 2160
rect 2065 2148 2069 2152
rect 2075 2148 2079 2156
rect 2095 2148 2099 2152
rect 2105 2148 2109 2152
rect 2125 2148 2129 2156
rect 1766 2047 1781 2059
rect 1714 2036 1718 2047
rect 1700 2028 1718 2036
rect 1700 2024 1704 2028
rect 1777 2024 1781 2047
rect 1785 2047 1794 2059
rect 1785 2024 1789 2047
rect 1845 2039 1849 2116
rect 1865 2093 1869 2116
rect 1885 2111 1889 2116
rect 1885 2104 1898 2111
rect 2005 2124 2009 2128
rect 2005 2119 2017 2124
rect 1865 2081 1874 2093
rect 1847 2027 1854 2039
rect 1850 1984 1854 2027
rect 1872 2024 1876 2081
rect 1894 2059 1898 2104
rect 1945 2059 1949 2108
rect 1955 2104 1959 2108
rect 1975 2062 1979 2108
rect 1985 2096 1989 2108
rect 1985 2090 1999 2096
rect 1946 2047 1949 2059
rect 1994 2059 1999 2090
rect 2013 2093 2017 2119
rect 2125 2124 2129 2128
rect 2125 2119 2137 2124
rect 1894 2036 1898 2047
rect 1880 2028 1898 2036
rect 1880 2024 1884 2028
rect 1945 2024 1949 2047
rect 1955 2046 1985 2050
rect 1955 2024 1959 2046
rect 1993 2041 1998 2047
rect 1985 2037 1998 2041
rect 1975 2032 1979 2036
rect 1985 2032 1989 2037
rect 2013 2000 2017 2081
rect 2065 2059 2069 2108
rect 2075 2104 2079 2108
rect 2095 2062 2099 2108
rect 2105 2096 2109 2108
rect 2105 2090 2119 2096
rect 2066 2047 2069 2059
rect 2114 2059 2119 2090
rect 2133 2093 2137 2119
rect 2065 2024 2069 2047
rect 2075 2046 2105 2050
rect 2075 2024 2079 2046
rect 2113 2041 2118 2047
rect 2105 2037 2118 2041
rect 2095 2032 2099 2036
rect 2105 2032 2109 2037
rect 2005 1996 2017 2000
rect 2005 1992 2009 1996
rect 1975 1944 1979 1952
rect 1985 1948 1989 1952
rect 2005 1944 2009 1952
rect 2133 2000 2137 2081
rect 2175 2079 2179 2116
rect 2195 2078 2199 2136
rect 2205 2104 2209 2136
rect 2227 2124 2231 2136
rect 2229 2112 2231 2124
rect 2237 2124 2241 2136
rect 2237 2112 2239 2124
rect 2205 2100 2238 2104
rect 2175 2024 2179 2067
rect 2125 1996 2137 2000
rect 2125 1992 2129 1996
rect 2095 1944 2099 1952
rect 2105 1948 2109 1952
rect 2125 1944 2129 1952
rect 2195 1984 2199 2066
rect 2214 2051 2218 2080
rect 2209 2043 2218 2051
rect 2209 1984 2213 2043
rect 2234 2036 2238 2100
rect 2235 2024 2238 2036
rect 2229 1984 2233 2024
rect 2243 2002 2247 2112
rect 2259 2022 2263 2136
rect 2305 2132 2309 2136
rect 2275 2128 2309 2132
rect 2241 1984 2245 1990
rect 2261 1984 2265 2010
rect 2275 2002 2279 2128
rect 2313 2124 2317 2136
rect 2287 2120 2317 2124
rect 2299 2119 2317 2120
rect 2333 2115 2337 2136
rect 2313 2111 2337 2115
rect 2313 2016 2319 2111
rect 2343 2087 2347 2136
rect 2343 2029 2347 2075
rect 2365 2048 2369 2116
rect 2367 2036 2369 2048
rect 2425 2039 2429 2116
rect 2445 2093 2449 2116
rect 2465 2111 2469 2116
rect 2465 2104 2478 2111
rect 2445 2081 2454 2093
rect 2343 2023 2351 2029
rect 2365 2024 2369 2036
rect 2427 2027 2434 2039
rect 2287 1990 2311 1992
rect 2275 1988 2311 1990
rect 2307 1984 2311 1988
rect 2315 1984 2319 2016
rect 2335 1964 2339 2004
rect 2347 1994 2351 2023
rect 2343 1987 2351 1994
rect 2343 1964 2347 1987
rect 2430 1984 2434 2027
rect 2452 2024 2456 2081
rect 2474 2059 2478 2104
rect 2511 2059 2515 2136
rect 2531 2059 2535 2136
rect 2691 2148 2695 2156
rect 2711 2148 2715 2152
rect 2721 2148 2725 2152
rect 2741 2148 2745 2156
rect 2835 2156 2889 2160
rect 2931 2156 2935 2160
rect 2991 2156 2995 2160
rect 3011 2156 3015 2160
rect 3031 2156 3035 2160
rect 3051 2156 3055 2160
rect 3132 2156 3136 2160
rect 3154 2156 3158 2160
rect 3162 2156 3166 2160
rect 3211 2156 3215 2160
rect 3271 2156 3275 2160
rect 3291 2156 3295 2160
rect 3311 2156 3315 2160
rect 3331 2156 3335 2160
rect 3391 2156 3395 2160
rect 3411 2156 3415 2160
rect 3475 2156 3479 2160
rect 3495 2156 3499 2160
rect 3505 2156 3509 2160
rect 3527 2156 3531 2160
rect 3537 2156 3541 2160
rect 3559 2156 3563 2160
rect 3605 2156 3609 2160
rect 3613 2156 3617 2160
rect 3633 2156 3637 2160
rect 3643 2156 3647 2160
rect 3665 2156 3669 2160
rect 3725 2156 3729 2160
rect 3745 2156 3749 2160
rect 3805 2156 3809 2160
rect 3825 2156 3829 2160
rect 3845 2156 3849 2160
rect 3865 2156 3869 2160
rect 3925 2156 3929 2160
rect 3971 2156 3975 2160
rect 3991 2156 3995 2160
rect 4011 2156 4015 2160
rect 4073 2156 4077 2160
rect 4083 2156 4087 2160
rect 4165 2156 4169 2160
rect 4185 2156 4189 2160
rect 4235 2156 4239 2160
rect 4255 2156 4259 2160
rect 4265 2156 4269 2160
rect 4287 2156 4291 2160
rect 4297 2156 4301 2160
rect 4319 2156 4323 2160
rect 4365 2156 4369 2160
rect 4373 2156 4377 2160
rect 4393 2156 4397 2160
rect 4403 2156 4407 2160
rect 4425 2156 4429 2160
rect 4471 2156 4475 2160
rect 4531 2156 4535 2160
rect 4551 2156 4555 2160
rect 4571 2156 4575 2160
rect 4591 2156 4595 2160
rect 4651 2156 4655 2160
rect 4671 2156 4675 2160
rect 4745 2156 4749 2160
rect 4765 2156 4769 2160
rect 4785 2156 4789 2160
rect 4845 2156 4849 2160
rect 4865 2156 4869 2160
rect 4911 2156 4915 2160
rect 4931 2156 4935 2160
rect 4951 2156 4955 2160
rect 4971 2156 4975 2160
rect 5053 2156 5057 2160
rect 5063 2156 5067 2160
rect 5125 2156 5129 2160
rect 5145 2156 5149 2160
rect 5191 2156 5195 2160
rect 5211 2156 5215 2160
rect 5231 2156 5235 2160
rect 5305 2156 5309 2160
rect 5325 2156 5329 2160
rect 5345 2156 5349 2160
rect 5365 2156 5369 2160
rect 5411 2156 5415 2160
rect 5431 2156 5435 2160
rect 5451 2156 5455 2160
rect 5471 2156 5475 2160
rect 5545 2156 5549 2160
rect 5565 2156 5569 2160
rect 5625 2156 5629 2160
rect 5645 2156 5649 2160
rect 5665 2156 5669 2160
rect 5685 2156 5689 2160
rect 5745 2156 5749 2160
rect 5793 2156 5797 2160
rect 5803 2156 5807 2160
rect 5871 2156 5875 2160
rect 5893 2156 5897 2160
rect 5903 2156 5907 2160
rect 5923 2156 5927 2160
rect 5931 2156 5935 2160
rect 5977 2156 5981 2160
rect 5999 2156 6003 2160
rect 6009 2156 6013 2160
rect 6031 2156 6035 2160
rect 6041 2156 6045 2160
rect 6061 2156 6065 2160
rect 6115 2156 6119 2160
rect 6135 2156 6139 2160
rect 6145 2156 6149 2160
rect 6167 2156 6171 2160
rect 6177 2156 6181 2160
rect 6199 2156 6203 2160
rect 6245 2156 6249 2160
rect 6253 2156 6257 2160
rect 6273 2156 6277 2160
rect 6283 2156 6287 2160
rect 6305 2156 6309 2160
rect 6351 2156 6405 2160
rect 6474 2156 6478 2160
rect 6482 2156 6486 2160
rect 6504 2156 6508 2160
rect 6571 2156 6575 2160
rect 6591 2156 6595 2160
rect 6611 2156 6615 2160
rect 2751 2148 2755 2152
rect 2825 2148 2829 2152
rect 2835 2148 2839 2156
rect 2855 2148 2859 2152
rect 2865 2148 2869 2152
rect 2885 2148 2889 2156
rect 2691 2124 2695 2128
rect 2683 2119 2695 2124
rect 2506 2047 2515 2059
rect 2474 2036 2478 2047
rect 2460 2028 2478 2036
rect 2460 2024 2464 2028
rect 2511 2024 2515 2047
rect 2519 2047 2534 2059
rect 2519 2024 2523 2047
rect 2628 2039 2632 2096
rect 2605 2027 2613 2039
rect 2625 2027 2632 2039
rect 2605 1984 2609 2027
rect 2636 2019 2640 2096
rect 2644 2039 2648 2096
rect 2683 2093 2687 2119
rect 2885 2124 2889 2128
rect 2885 2119 2897 2124
rect 2711 2096 2715 2108
rect 2644 2027 2654 2039
rect 2634 2000 2640 2007
rect 2625 1996 2640 2000
rect 2654 1996 2660 2027
rect 2683 2000 2687 2081
rect 2701 2090 2715 2096
rect 2701 2059 2706 2090
rect 2721 2062 2725 2108
rect 2741 2104 2745 2108
rect 2702 2041 2707 2047
rect 2751 2059 2755 2108
rect 2825 2059 2829 2108
rect 2835 2104 2839 2108
rect 2855 2062 2859 2108
rect 2865 2096 2869 2108
rect 2865 2090 2879 2096
rect 2715 2046 2745 2050
rect 2702 2037 2715 2041
rect 2711 2032 2715 2037
rect 2721 2032 2725 2036
rect 2683 1996 2695 2000
rect 2625 1984 2629 1996
rect 2645 1992 2660 1996
rect 2691 1992 2695 1996
rect 2645 1984 2649 1992
rect 2741 2024 2745 2046
rect 2751 2047 2754 2059
rect 2826 2047 2829 2059
rect 2874 2059 2879 2090
rect 2893 2093 2897 2119
rect 2751 2024 2755 2047
rect 2825 2024 2829 2047
rect 2835 2046 2865 2050
rect 2835 2024 2839 2046
rect 2873 2041 2878 2047
rect 2865 2037 2878 2041
rect 2855 2032 2859 2036
rect 2865 2032 2869 2037
rect 2691 1944 2695 1952
rect 2711 1948 2715 1952
rect 2721 1944 2725 1952
rect 2893 2000 2897 2081
rect 2931 2079 2935 2136
rect 2991 2109 2995 2116
rect 2926 2067 2935 2079
rect 2885 1996 2897 2000
rect 2885 1992 2889 1996
rect 2931 1984 2935 2067
rect 2980 2105 2995 2109
rect 2980 2059 2986 2105
rect 3011 2093 3015 2116
rect 3031 2093 3035 2116
rect 3006 2081 3015 2093
rect 2981 2032 2986 2047
rect 3009 2032 3015 2081
rect 2981 2028 2995 2032
rect 2991 2024 2995 2028
rect 3001 2028 3015 2032
rect 3001 2024 3005 2028
rect 3031 2024 3035 2081
rect 3051 2059 3055 2116
rect 3132 2093 3136 2136
rect 3125 2081 3134 2093
rect 3051 2047 3053 2059
rect 3051 2032 3055 2047
rect 3041 2028 3055 2032
rect 3041 2024 3045 2028
rect 3125 2024 3129 2081
rect 3154 2079 3158 2116
rect 3162 2112 3166 2116
rect 3162 2106 3181 2112
rect 3174 2093 3181 2106
rect 3154 2044 3160 2067
rect 3174 2044 3181 2081
rect 3211 2079 3215 2136
rect 3271 2109 3275 2116
rect 3206 2067 3215 2079
rect 3145 2038 3160 2044
rect 3165 2038 3181 2044
rect 3145 2024 3149 2038
rect 3165 2024 3169 2038
rect 2855 1944 2859 1952
rect 2865 1948 2869 1952
rect 2885 1944 2889 1952
rect 3211 1984 3215 2067
rect 3260 2105 3275 2109
rect 3260 2059 3266 2105
rect 3291 2093 3295 2116
rect 3311 2093 3315 2116
rect 3286 2081 3295 2093
rect 3261 2032 3266 2047
rect 3289 2032 3295 2081
rect 3261 2028 3275 2032
rect 3271 2024 3275 2028
rect 3281 2028 3295 2032
rect 3281 2024 3285 2028
rect 3311 2024 3315 2081
rect 3331 2059 3335 2116
rect 3391 2059 3395 2136
rect 3411 2059 3415 2136
rect 3475 2079 3479 2116
rect 3495 2078 3499 2136
rect 3505 2104 3509 2136
rect 3527 2124 3531 2136
rect 3529 2112 3531 2124
rect 3537 2124 3541 2136
rect 3537 2112 3539 2124
rect 3505 2100 3538 2104
rect 3331 2047 3333 2059
rect 3386 2047 3395 2059
rect 3331 2032 3335 2047
rect 3321 2028 3335 2032
rect 3321 2024 3325 2028
rect 3391 2024 3395 2047
rect 3399 2047 3414 2059
rect 3399 2024 3403 2047
rect 3475 2024 3479 2067
rect 3495 1984 3499 2066
rect 3514 2051 3518 2080
rect 3509 2043 3518 2051
rect 3509 1984 3513 2043
rect 3534 2036 3538 2100
rect 3535 2024 3538 2036
rect 3529 1984 3533 2024
rect 3543 2002 3547 2112
rect 3559 2022 3563 2136
rect 3605 2132 3609 2136
rect 3575 2128 3609 2132
rect 3541 1984 3545 1990
rect 3561 1984 3565 2010
rect 3575 2002 3579 2128
rect 3613 2124 3617 2136
rect 3587 2120 3617 2124
rect 3599 2119 3617 2120
rect 3633 2115 3637 2136
rect 3613 2111 3637 2115
rect 3613 2016 3619 2111
rect 3643 2087 3647 2136
rect 3643 2029 3647 2075
rect 3665 2048 3669 2116
rect 3725 2059 3729 2136
rect 3745 2059 3749 2136
rect 3805 2059 3809 2116
rect 3825 2093 3829 2116
rect 3845 2093 3849 2116
rect 3865 2109 3869 2116
rect 3865 2105 3880 2109
rect 3845 2081 3854 2093
rect 3667 2036 3669 2048
rect 3726 2047 3741 2059
rect 3643 2023 3651 2029
rect 3665 2024 3669 2036
rect 3737 2024 3741 2047
rect 3745 2047 3754 2059
rect 3807 2047 3809 2059
rect 3745 2024 3749 2047
rect 3805 2032 3809 2047
rect 3805 2028 3819 2032
rect 3815 2024 3819 2028
rect 3825 2024 3829 2081
rect 3845 2032 3851 2081
rect 3874 2059 3880 2105
rect 3925 2079 3929 2136
rect 3971 2111 3975 2116
rect 3962 2104 3975 2111
rect 3925 2067 3934 2079
rect 3874 2032 3879 2047
rect 3845 2028 3859 2032
rect 3855 2024 3859 2028
rect 3865 2028 3879 2032
rect 3865 2024 3869 2028
rect 3587 1990 3611 1992
rect 3575 1988 3611 1990
rect 3607 1984 3611 1988
rect 3615 1984 3619 2016
rect 3635 1964 3639 2004
rect 3647 1994 3651 2023
rect 3643 1987 3651 1994
rect 3643 1964 3647 1987
rect 3925 1984 3929 2067
rect 3962 2059 3966 2104
rect 3991 2093 3995 2116
rect 3986 2081 3995 2093
rect 3962 2036 3966 2047
rect 3962 2028 3980 2036
rect 3976 2024 3980 2028
rect 3984 2024 3988 2081
rect 4011 2039 4015 2116
rect 4073 2096 4077 2116
rect 4069 2089 4077 2096
rect 4083 2096 4087 2116
rect 4083 2089 4097 2096
rect 4069 2073 4075 2089
rect 4066 2061 4075 2073
rect 4006 2027 4013 2039
rect 4006 1984 4010 2027
rect 4071 1984 4075 2061
rect 4091 2073 4097 2089
rect 4091 2061 4094 2073
rect 4091 1984 4095 2061
rect 4165 2059 4169 2136
rect 4185 2059 4189 2136
rect 4235 2079 4239 2116
rect 4255 2078 4259 2136
rect 4265 2104 4269 2136
rect 4287 2124 4291 2136
rect 4289 2112 4291 2124
rect 4297 2124 4301 2136
rect 4297 2112 4299 2124
rect 4265 2100 4298 2104
rect 4166 2047 4181 2059
rect 4177 2024 4181 2047
rect 4185 2047 4194 2059
rect 4185 2024 4189 2047
rect 4235 2024 4239 2067
rect 4255 1984 4259 2066
rect 4274 2051 4278 2080
rect 4269 2043 4278 2051
rect 4269 1984 4273 2043
rect 4294 2036 4298 2100
rect 4295 2024 4298 2036
rect 4289 1984 4293 2024
rect 4303 2002 4307 2112
rect 4319 2022 4323 2136
rect 4365 2132 4369 2136
rect 4335 2128 4369 2132
rect 4301 1984 4305 1990
rect 4321 1984 4325 2010
rect 4335 2002 4339 2128
rect 4373 2124 4377 2136
rect 4347 2120 4377 2124
rect 4359 2119 4377 2120
rect 4393 2115 4397 2136
rect 4373 2111 4397 2115
rect 4373 2016 4379 2111
rect 4403 2087 4407 2136
rect 4403 2029 4407 2075
rect 4425 2048 4429 2116
rect 4471 2079 4475 2136
rect 4531 2109 4535 2116
rect 4466 2067 4475 2079
rect 4427 2036 4429 2048
rect 4403 2023 4411 2029
rect 4425 2024 4429 2036
rect 4347 1990 4371 1992
rect 4335 1988 4371 1990
rect 4367 1984 4371 1988
rect 4375 1984 4379 2016
rect 4395 1964 4399 2004
rect 4407 1994 4411 2023
rect 4403 1987 4411 1994
rect 4403 1964 4407 1987
rect 4471 1984 4475 2067
rect 4520 2105 4535 2109
rect 4520 2059 4526 2105
rect 4551 2093 4555 2116
rect 4571 2093 4575 2116
rect 4546 2081 4555 2093
rect 4521 2032 4526 2047
rect 4549 2032 4555 2081
rect 4521 2028 4535 2032
rect 4531 2024 4535 2028
rect 4541 2028 4555 2032
rect 4541 2024 4545 2028
rect 4571 2024 4575 2081
rect 4591 2059 4595 2116
rect 4651 2059 4655 2136
rect 4671 2059 4675 2136
rect 4591 2047 4593 2059
rect 4646 2047 4655 2059
rect 4591 2032 4595 2047
rect 4581 2028 4595 2032
rect 4581 2024 4585 2028
rect 4651 2024 4655 2047
rect 4659 2047 4674 2059
rect 4659 2024 4663 2047
rect 4745 2039 4749 2116
rect 4765 2093 4769 2116
rect 4785 2111 4789 2116
rect 4785 2104 4798 2111
rect 4765 2081 4774 2093
rect 4747 2027 4754 2039
rect 4750 1984 4754 2027
rect 4772 2024 4776 2081
rect 4794 2059 4798 2104
rect 4845 2059 4849 2136
rect 4865 2059 4869 2136
rect 4911 2109 4915 2116
rect 4900 2105 4915 2109
rect 4900 2059 4906 2105
rect 4931 2093 4935 2116
rect 4951 2093 4955 2116
rect 4926 2081 4935 2093
rect 4846 2047 4861 2059
rect 4794 2036 4798 2047
rect 4780 2028 4798 2036
rect 4780 2024 4784 2028
rect 4857 2024 4861 2047
rect 4865 2047 4874 2059
rect 4865 2024 4869 2047
rect 4901 2032 4906 2047
rect 4929 2032 4935 2081
rect 4901 2028 4915 2032
rect 4911 2024 4915 2028
rect 4921 2028 4935 2032
rect 4921 2024 4925 2028
rect 4951 2024 4955 2081
rect 4971 2059 4975 2116
rect 5053 2096 5057 2116
rect 5043 2089 5057 2096
rect 5063 2096 5067 2116
rect 5063 2089 5071 2096
rect 5043 2073 5049 2089
rect 5046 2061 5049 2073
rect 4971 2047 4973 2059
rect 4971 2032 4975 2047
rect 4961 2028 4975 2032
rect 4961 2024 4965 2028
rect 5045 1984 5049 2061
rect 5065 2073 5071 2089
rect 5065 2061 5074 2073
rect 5065 1984 5069 2061
rect 5125 2059 5129 2136
rect 5145 2059 5149 2136
rect 5191 2129 5195 2136
rect 5211 2129 5215 2136
rect 5182 2124 5195 2129
rect 5182 2079 5186 2124
rect 5126 2047 5141 2059
rect 5137 2024 5141 2047
rect 5145 2047 5154 2059
rect 5145 2024 5149 2047
rect 5182 2033 5186 2067
rect 5201 2123 5215 2129
rect 5201 2059 5205 2123
rect 5231 2108 5235 2116
rect 5225 2096 5235 2108
rect 5305 2059 5309 2116
rect 5325 2093 5329 2116
rect 5345 2093 5349 2116
rect 5365 2109 5369 2116
rect 5411 2109 5415 2116
rect 5365 2105 5380 2109
rect 5345 2081 5354 2093
rect 5307 2047 5309 2059
rect 5182 2028 5195 2033
rect 5191 2024 5195 2028
rect 5201 2024 5205 2047
rect 5221 2024 5225 2029
rect 5305 2032 5309 2047
rect 5305 2028 5319 2032
rect 5315 2024 5319 2028
rect 5325 2024 5329 2081
rect 5345 2032 5351 2081
rect 5374 2059 5380 2105
rect 5400 2105 5415 2109
rect 5400 2059 5406 2105
rect 5431 2093 5435 2116
rect 5451 2093 5455 2116
rect 5426 2081 5435 2093
rect 5374 2032 5379 2047
rect 5345 2028 5359 2032
rect 5355 2024 5359 2028
rect 5365 2028 5379 2032
rect 5401 2032 5406 2047
rect 5429 2032 5435 2081
rect 5401 2028 5415 2032
rect 5365 2024 5369 2028
rect 5411 2024 5415 2028
rect 5421 2028 5435 2032
rect 5421 2024 5425 2028
rect 5451 2024 5455 2081
rect 5471 2059 5475 2116
rect 5545 2059 5549 2136
rect 5565 2059 5569 2136
rect 5625 2059 5629 2116
rect 5645 2093 5649 2116
rect 5665 2093 5669 2116
rect 5685 2109 5689 2116
rect 5685 2105 5700 2109
rect 5665 2081 5674 2093
rect 5471 2047 5473 2059
rect 5546 2047 5561 2059
rect 5471 2032 5475 2047
rect 5461 2028 5475 2032
rect 5461 2024 5465 2028
rect 5557 2024 5561 2047
rect 5565 2047 5574 2059
rect 5627 2047 5629 2059
rect 5565 2024 5569 2047
rect 5625 2032 5629 2047
rect 5625 2028 5639 2032
rect 5635 2024 5639 2028
rect 5645 2024 5649 2081
rect 5665 2032 5671 2081
rect 5694 2059 5700 2105
rect 5745 2079 5749 2136
rect 5793 2096 5797 2116
rect 5789 2089 5797 2096
rect 5803 2096 5807 2116
rect 5803 2089 5817 2096
rect 5745 2067 5754 2079
rect 5789 2073 5795 2089
rect 5694 2032 5699 2047
rect 5665 2028 5679 2032
rect 5675 2024 5679 2028
rect 5685 2028 5699 2032
rect 5685 2024 5689 2028
rect 5745 1984 5749 2067
rect 5786 2061 5795 2073
rect 5791 1984 5795 2061
rect 5811 2073 5817 2089
rect 5811 2061 5814 2073
rect 5811 1984 5815 2061
rect 5871 2048 5875 2116
rect 5893 2087 5897 2136
rect 5903 2115 5907 2136
rect 5923 2124 5927 2136
rect 5931 2132 5935 2136
rect 5931 2128 5965 2132
rect 5923 2120 5953 2124
rect 5923 2119 5941 2120
rect 5903 2111 5927 2115
rect 5871 2036 5873 2048
rect 5871 2024 5875 2036
rect 5893 2029 5897 2075
rect 5889 2023 5897 2029
rect 5889 1994 5893 2023
rect 5921 2016 5927 2111
rect 5889 1987 5897 1994
rect 5893 1964 5897 1987
rect 5901 1964 5905 2004
rect 5921 1984 5925 2016
rect 5961 2002 5965 2128
rect 5977 2022 5981 2136
rect 5999 2124 6003 2136
rect 6001 2112 6003 2124
rect 6009 2124 6013 2136
rect 6009 2112 6011 2124
rect 5929 1990 5953 1992
rect 5929 1988 5965 1990
rect 5929 1984 5933 1988
rect 5975 1984 5979 2010
rect 5993 2002 5997 2112
rect 6031 2104 6035 2136
rect 6002 2100 6035 2104
rect 6002 2036 6006 2100
rect 6022 2051 6026 2080
rect 6041 2078 6045 2136
rect 6061 2079 6065 2116
rect 6115 2079 6119 2116
rect 6135 2078 6139 2136
rect 6145 2104 6149 2136
rect 6167 2124 6171 2136
rect 6169 2112 6171 2124
rect 6177 2124 6181 2136
rect 6177 2112 6179 2124
rect 6145 2100 6178 2104
rect 6022 2043 6031 2051
rect 6002 2024 6005 2036
rect 5995 1984 5999 1990
rect 6007 1984 6011 2024
rect 6027 1984 6031 2043
rect 6041 1984 6045 2066
rect 6061 2024 6065 2067
rect 6115 2024 6119 2067
rect 6135 1984 6139 2066
rect 6154 2051 6158 2080
rect 6149 2043 6158 2051
rect 6149 1984 6153 2043
rect 6174 2036 6178 2100
rect 6175 2024 6178 2036
rect 6169 1984 6173 2024
rect 6183 2002 6187 2112
rect 6199 2022 6203 2136
rect 6245 2132 6249 2136
rect 6215 2128 6249 2132
rect 6181 1984 6185 1990
rect 6201 1984 6205 2010
rect 6215 2002 6219 2128
rect 6253 2124 6257 2136
rect 6227 2120 6257 2124
rect 6239 2119 6257 2120
rect 6273 2115 6277 2136
rect 6253 2111 6277 2115
rect 6253 2016 6259 2111
rect 6283 2087 6287 2136
rect 6351 2148 6355 2156
rect 6371 2148 6375 2152
rect 6381 2148 6385 2152
rect 6401 2148 6405 2156
rect 6411 2148 6415 2152
rect 6351 2124 6355 2128
rect 6343 2119 6355 2124
rect 6283 2029 6287 2075
rect 6305 2048 6309 2116
rect 6343 2093 6347 2119
rect 6474 2112 6478 2116
rect 6371 2096 6375 2108
rect 6307 2036 6309 2048
rect 6283 2023 6291 2029
rect 6305 2024 6309 2036
rect 6227 1990 6251 1992
rect 6215 1988 6251 1990
rect 6247 1984 6251 1988
rect 6255 1984 6259 2016
rect 6275 1964 6279 2004
rect 6287 1994 6291 2023
rect 6283 1987 6291 1994
rect 6283 1964 6287 1987
rect 6343 2000 6347 2081
rect 6361 2090 6375 2096
rect 6361 2059 6366 2090
rect 6381 2062 6385 2108
rect 6401 2104 6405 2108
rect 6362 2041 6367 2047
rect 6411 2059 6415 2108
rect 6459 2106 6478 2112
rect 6459 2093 6466 2106
rect 6375 2046 6405 2050
rect 6362 2037 6375 2041
rect 6371 2032 6375 2037
rect 6381 2032 6385 2036
rect 6343 1996 6355 2000
rect 6351 1992 6355 1996
rect 6401 2024 6405 2046
rect 6411 2047 6414 2059
rect 6411 2024 6415 2047
rect 6459 2044 6466 2081
rect 6482 2079 6486 2116
rect 6504 2093 6508 2136
rect 6571 2111 6575 2116
rect 6562 2104 6575 2111
rect 6506 2081 6515 2093
rect 6480 2044 6486 2067
rect 6459 2038 6475 2044
rect 6480 2038 6495 2044
rect 6471 2024 6475 2038
rect 6491 2024 6495 2038
rect 6511 2024 6515 2081
rect 6562 2059 6566 2104
rect 6591 2093 6595 2116
rect 6586 2081 6595 2093
rect 6562 2036 6566 2047
rect 6562 2028 6580 2036
rect 6576 2024 6580 2028
rect 6584 2024 6588 2081
rect 6611 2039 6615 2116
rect 6606 2027 6613 2039
rect 6351 1944 6355 1952
rect 6371 1948 6375 1952
rect 6381 1944 6385 1952
rect 6606 1984 6610 2027
rect 57 1940 61 1944
rect 65 1940 69 1944
rect 125 1940 129 1944
rect 145 1940 149 1944
rect 205 1940 209 1944
rect 225 1940 229 1944
rect 245 1940 249 1944
rect 305 1940 309 1944
rect 325 1940 329 1944
rect 345 1940 349 1944
rect 405 1940 409 1944
rect 425 1940 429 1944
rect 471 1940 475 1944
rect 491 1940 495 1944
rect 511 1940 515 1944
rect 597 1940 601 1944
rect 605 1940 609 1944
rect 656 1940 660 1944
rect 664 1940 668 1944
rect 686 1940 690 1944
rect 751 1940 755 1944
rect 771 1940 775 1944
rect 791 1940 795 1944
rect 851 1940 855 1944
rect 859 1940 863 1944
rect 945 1940 949 1944
rect 965 1940 969 1944
rect 1011 1940 1045 1944
rect 1061 1940 1065 1944
rect 1071 1940 1075 1944
rect 1135 1940 1139 1944
rect 1155 1940 1159 1944
rect 1169 1940 1173 1944
rect 1189 1940 1193 1944
rect 1201 1940 1205 1944
rect 1221 1940 1225 1944
rect 1267 1940 1271 1944
rect 1275 1940 1279 1944
rect 1295 1940 1299 1944
rect 1303 1940 1307 1944
rect 1325 1940 1329 1944
rect 1371 1940 1375 1944
rect 1431 1940 1435 1944
rect 1441 1940 1445 1944
rect 1471 1940 1475 1944
rect 1481 1940 1485 1944
rect 1570 1940 1574 1944
rect 1592 1940 1596 1944
rect 1600 1940 1604 1944
rect 1670 1940 1674 1944
rect 1692 1940 1696 1944
rect 1700 1940 1704 1944
rect 1777 1940 1781 1944
rect 1785 1940 1789 1944
rect 1850 1940 1854 1944
rect 1872 1940 1876 1944
rect 1880 1940 1884 1944
rect 1945 1940 1949 1944
rect 1955 1940 1959 1944
rect 1975 1940 2009 1944
rect 2065 1940 2069 1944
rect 2075 1940 2079 1944
rect 2095 1940 2129 1944
rect 2175 1940 2179 1944
rect 2195 1940 2199 1944
rect 2209 1940 2213 1944
rect 2229 1940 2233 1944
rect 2241 1940 2245 1944
rect 2261 1940 2265 1944
rect 2307 1940 2311 1944
rect 2315 1940 2319 1944
rect 2335 1940 2339 1944
rect 2343 1940 2347 1944
rect 2365 1940 2369 1944
rect 2430 1940 2434 1944
rect 2452 1940 2456 1944
rect 2460 1940 2464 1944
rect 2511 1940 2515 1944
rect 2519 1940 2523 1944
rect 2605 1940 2609 1944
rect 2625 1940 2629 1944
rect 2645 1940 2649 1944
rect 2691 1940 2725 1944
rect 2741 1940 2745 1944
rect 2751 1940 2755 1944
rect 2825 1940 2829 1944
rect 2835 1940 2839 1944
rect 2855 1940 2889 1944
rect 2931 1940 2935 1944
rect 2991 1940 2995 1944
rect 3001 1940 3005 1944
rect 3031 1940 3035 1944
rect 3041 1940 3045 1944
rect 3125 1940 3129 1944
rect 3145 1940 3149 1944
rect 3165 1940 3169 1944
rect 3211 1940 3215 1944
rect 3271 1940 3275 1944
rect 3281 1940 3285 1944
rect 3311 1940 3315 1944
rect 3321 1940 3325 1944
rect 3391 1940 3395 1944
rect 3399 1940 3403 1944
rect 3475 1940 3479 1944
rect 3495 1940 3499 1944
rect 3509 1940 3513 1944
rect 3529 1940 3533 1944
rect 3541 1940 3545 1944
rect 3561 1940 3565 1944
rect 3607 1940 3611 1944
rect 3615 1940 3619 1944
rect 3635 1940 3639 1944
rect 3643 1940 3647 1944
rect 3665 1940 3669 1944
rect 3737 1940 3741 1944
rect 3745 1940 3749 1944
rect 3815 1940 3819 1944
rect 3825 1940 3829 1944
rect 3855 1940 3859 1944
rect 3865 1940 3869 1944
rect 3925 1940 3929 1944
rect 3976 1940 3980 1944
rect 3984 1940 3988 1944
rect 4006 1940 4010 1944
rect 4071 1940 4075 1944
rect 4091 1940 4095 1944
rect 4177 1940 4181 1944
rect 4185 1940 4189 1944
rect 4235 1940 4239 1944
rect 4255 1940 4259 1944
rect 4269 1940 4273 1944
rect 4289 1940 4293 1944
rect 4301 1940 4305 1944
rect 4321 1940 4325 1944
rect 4367 1940 4371 1944
rect 4375 1940 4379 1944
rect 4395 1940 4399 1944
rect 4403 1940 4407 1944
rect 4425 1940 4429 1944
rect 4471 1940 4475 1944
rect 4531 1940 4535 1944
rect 4541 1940 4545 1944
rect 4571 1940 4575 1944
rect 4581 1940 4585 1944
rect 4651 1940 4655 1944
rect 4659 1940 4663 1944
rect 4750 1940 4754 1944
rect 4772 1940 4776 1944
rect 4780 1940 4784 1944
rect 4857 1940 4861 1944
rect 4865 1940 4869 1944
rect 4911 1940 4915 1944
rect 4921 1940 4925 1944
rect 4951 1940 4955 1944
rect 4961 1940 4965 1944
rect 5045 1940 5049 1944
rect 5065 1940 5069 1944
rect 5137 1940 5141 1944
rect 5145 1940 5149 1944
rect 5191 1940 5195 1944
rect 5201 1940 5205 1944
rect 5221 1940 5225 1944
rect 5315 1940 5319 1944
rect 5325 1940 5329 1944
rect 5355 1940 5359 1944
rect 5365 1940 5369 1944
rect 5411 1940 5415 1944
rect 5421 1940 5425 1944
rect 5451 1940 5455 1944
rect 5461 1940 5465 1944
rect 5557 1940 5561 1944
rect 5565 1940 5569 1944
rect 5635 1940 5639 1944
rect 5645 1940 5649 1944
rect 5675 1940 5679 1944
rect 5685 1940 5689 1944
rect 5745 1940 5749 1944
rect 5791 1940 5795 1944
rect 5811 1940 5815 1944
rect 5871 1940 5875 1944
rect 5893 1940 5897 1944
rect 5901 1940 5905 1944
rect 5921 1940 5925 1944
rect 5929 1940 5933 1944
rect 5975 1940 5979 1944
rect 5995 1940 5999 1944
rect 6007 1940 6011 1944
rect 6027 1940 6031 1944
rect 6041 1940 6045 1944
rect 6061 1940 6065 1944
rect 6115 1940 6119 1944
rect 6135 1940 6139 1944
rect 6149 1940 6153 1944
rect 6169 1940 6173 1944
rect 6181 1940 6185 1944
rect 6201 1940 6205 1944
rect 6247 1940 6251 1944
rect 6255 1940 6259 1944
rect 6275 1940 6279 1944
rect 6283 1940 6287 1944
rect 6305 1940 6309 1944
rect 6351 1940 6385 1944
rect 6401 1940 6405 1944
rect 6411 1940 6415 1944
rect 6471 1940 6475 1944
rect 6491 1940 6495 1944
rect 6511 1940 6515 1944
rect 6576 1940 6580 1944
rect 6584 1940 6588 1944
rect 6606 1940 6610 1944
rect 45 1916 49 1920
rect 91 1916 95 1920
rect 113 1916 117 1920
rect 121 1916 125 1920
rect 141 1916 145 1920
rect 149 1916 153 1920
rect 195 1916 199 1920
rect 215 1916 219 1920
rect 227 1916 231 1920
rect 247 1916 251 1920
rect 261 1916 265 1920
rect 281 1916 285 1920
rect 331 1916 335 1920
rect 339 1916 343 1920
rect 437 1916 441 1920
rect 445 1916 449 1920
rect 505 1916 509 1920
rect 570 1916 574 1920
rect 592 1916 596 1920
rect 600 1916 604 1920
rect 651 1916 655 1920
rect 673 1916 677 1920
rect 681 1916 685 1920
rect 701 1916 705 1920
rect 709 1916 713 1920
rect 755 1916 759 1920
rect 775 1916 779 1920
rect 787 1916 791 1920
rect 807 1916 811 1920
rect 821 1916 825 1920
rect 841 1916 845 1920
rect 905 1916 909 1920
rect 925 1916 929 1920
rect 945 1916 949 1920
rect 991 1916 995 1920
rect 1013 1916 1017 1920
rect 1035 1916 1039 1920
rect 1091 1916 1095 1920
rect 1156 1916 1160 1920
rect 1164 1916 1168 1920
rect 1186 1916 1190 1920
rect 1265 1916 1269 1920
rect 1285 1916 1289 1920
rect 1345 1916 1349 1920
rect 1365 1916 1369 1920
rect 1385 1916 1389 1920
rect 1431 1916 1435 1920
rect 1495 1916 1499 1920
rect 1515 1916 1519 1920
rect 1529 1916 1533 1920
rect 1549 1916 1553 1920
rect 1561 1916 1565 1920
rect 1581 1916 1585 1920
rect 1627 1916 1631 1920
rect 1635 1916 1639 1920
rect 1655 1916 1659 1920
rect 1663 1916 1667 1920
rect 1685 1916 1689 1920
rect 1731 1916 1735 1920
rect 1791 1916 1795 1920
rect 1801 1916 1805 1920
rect 1831 1916 1835 1920
rect 1841 1916 1845 1920
rect 1911 1916 1915 1920
rect 1919 1916 1923 1920
rect 1996 1916 2000 1920
rect 2004 1916 2008 1920
rect 2026 1916 2030 1920
rect 2091 1916 2095 1920
rect 2113 1916 2117 1920
rect 2121 1916 2125 1920
rect 2141 1916 2145 1920
rect 2149 1916 2153 1920
rect 2195 1916 2199 1920
rect 2215 1916 2219 1920
rect 2227 1916 2231 1920
rect 2247 1916 2251 1920
rect 2261 1916 2265 1920
rect 2281 1916 2285 1920
rect 2355 1916 2359 1920
rect 2365 1916 2369 1920
rect 2395 1916 2399 1920
rect 2405 1916 2409 1920
rect 2451 1916 2455 1920
rect 2511 1916 2515 1920
rect 2519 1916 2523 1920
rect 2591 1916 2595 1920
rect 2613 1916 2617 1920
rect 2621 1916 2625 1920
rect 2641 1916 2645 1920
rect 2649 1916 2653 1920
rect 2695 1916 2699 1920
rect 2715 1916 2719 1920
rect 2727 1916 2731 1920
rect 2747 1916 2751 1920
rect 2761 1916 2765 1920
rect 2781 1916 2785 1920
rect 2831 1916 2835 1920
rect 2851 1916 2855 1920
rect 2871 1916 2875 1920
rect 2950 1916 2954 1920
rect 2972 1916 2976 1920
rect 2980 1916 2984 1920
rect 3031 1916 3035 1920
rect 3039 1916 3043 1920
rect 3125 1916 3129 1920
rect 3145 1916 3149 1920
rect 3165 1916 3169 1920
rect 3225 1916 3229 1920
rect 3245 1916 3249 1920
rect 3265 1916 3269 1920
rect 3323 1916 3327 1920
rect 3345 1916 3349 1920
rect 3405 1916 3409 1920
rect 3425 1916 3429 1920
rect 3471 1916 3475 1920
rect 3479 1916 3483 1920
rect 3551 1916 3555 1920
rect 3571 1916 3575 1920
rect 3636 1916 3640 1920
rect 3644 1916 3648 1920
rect 3666 1916 3670 1920
rect 3745 1916 3749 1920
rect 3765 1916 3769 1920
rect 3825 1916 3829 1920
rect 3871 1916 3875 1920
rect 3891 1916 3895 1920
rect 3951 1916 3955 1920
rect 3959 1916 3963 1920
rect 4031 1916 4035 1920
rect 4041 1916 4045 1920
rect 4071 1916 4075 1920
rect 4081 1916 4085 1920
rect 4177 1916 4181 1920
rect 4185 1916 4189 1920
rect 4236 1916 4240 1920
rect 4244 1916 4248 1920
rect 4266 1916 4270 1920
rect 4331 1916 4335 1920
rect 4351 1916 4355 1920
rect 4416 1916 4420 1920
rect 4424 1916 4428 1920
rect 4446 1916 4450 1920
rect 4537 1916 4541 1920
rect 4545 1916 4549 1920
rect 4615 1916 4619 1920
rect 4625 1916 4629 1920
rect 4655 1916 4659 1920
rect 4665 1916 4669 1920
rect 4725 1916 4729 1920
rect 4771 1916 4775 1920
rect 4793 1916 4797 1920
rect 4801 1916 4805 1920
rect 4821 1916 4825 1920
rect 4829 1916 4833 1920
rect 4875 1916 4879 1920
rect 4895 1916 4899 1920
rect 4907 1916 4911 1920
rect 4927 1916 4931 1920
rect 4941 1916 4945 1920
rect 4961 1916 4965 1920
rect 5011 1916 5015 1920
rect 5031 1916 5035 1920
rect 5051 1916 5055 1920
rect 5111 1916 5115 1920
rect 5119 1916 5123 1920
rect 5196 1916 5200 1920
rect 5204 1916 5208 1920
rect 5226 1916 5230 1920
rect 5291 1916 5295 1920
rect 5311 1916 5315 1920
rect 5331 1916 5335 1920
rect 5391 1916 5395 1920
rect 5413 1916 5417 1920
rect 5485 1916 5489 1920
rect 5545 1916 5549 1920
rect 5610 1916 5614 1920
rect 5632 1916 5636 1920
rect 5640 1916 5644 1920
rect 5691 1916 5695 1920
rect 5711 1916 5715 1920
rect 5785 1916 5789 1920
rect 5805 1916 5809 1920
rect 5825 1916 5829 1920
rect 5845 1916 5849 1920
rect 5891 1916 5895 1920
rect 5913 1916 5917 1920
rect 5990 1916 5994 1920
rect 6012 1916 6016 1920
rect 6020 1916 6024 1920
rect 6095 1916 6099 1920
rect 6105 1916 6109 1920
rect 6135 1916 6139 1920
rect 6145 1916 6149 1920
rect 6191 1916 6225 1920
rect 6241 1916 6245 1920
rect 6251 1916 6255 1920
rect 6311 1916 6345 1920
rect 6361 1916 6365 1920
rect 6371 1916 6375 1920
rect 6431 1916 6435 1920
rect 6496 1916 6500 1920
rect 6504 1916 6508 1920
rect 6526 1916 6530 1920
rect 6605 1916 6609 1920
rect 6625 1916 6629 1920
rect 45 1793 49 1876
rect 113 1873 117 1896
rect 109 1866 117 1873
rect 109 1837 113 1866
rect 121 1856 125 1896
rect 141 1844 145 1876
rect 149 1872 153 1876
rect 149 1870 185 1872
rect 149 1868 173 1870
rect 91 1824 95 1836
rect 109 1831 117 1837
rect 91 1812 93 1824
rect 45 1781 54 1793
rect 45 1724 49 1781
rect 91 1744 95 1812
rect 113 1785 117 1831
rect 113 1724 117 1773
rect 141 1749 147 1844
rect 123 1745 147 1749
rect 123 1724 127 1745
rect 143 1740 161 1741
rect 143 1736 173 1740
rect 143 1724 147 1736
rect 181 1732 185 1858
rect 195 1850 199 1876
rect 215 1870 219 1876
rect 151 1728 185 1732
rect 151 1724 155 1728
rect 197 1724 201 1838
rect 213 1748 217 1858
rect 227 1836 231 1876
rect 222 1824 225 1836
rect 222 1760 226 1824
rect 247 1817 251 1876
rect 242 1809 251 1817
rect 242 1780 246 1809
rect 261 1794 265 1876
rect 281 1793 285 1836
rect 331 1813 335 1836
rect 326 1801 335 1813
rect 339 1813 343 1836
rect 437 1813 441 1836
rect 339 1801 354 1813
rect 426 1801 441 1813
rect 445 1813 449 1836
rect 445 1801 454 1813
rect 222 1756 255 1760
rect 221 1736 223 1748
rect 219 1724 223 1736
rect 229 1736 231 1748
rect 229 1724 233 1736
rect 251 1724 255 1756
rect 261 1724 265 1782
rect 281 1744 285 1781
rect 331 1724 335 1801
rect 351 1724 355 1801
rect 425 1724 429 1801
rect 445 1724 449 1801
rect 505 1793 509 1876
rect 570 1833 574 1876
rect 673 1873 677 1896
rect 669 1866 677 1873
rect 669 1837 673 1866
rect 681 1856 685 1896
rect 701 1844 705 1876
rect 709 1872 713 1876
rect 709 1870 745 1872
rect 709 1868 733 1870
rect 567 1821 574 1833
rect 505 1781 514 1793
rect 505 1724 509 1781
rect 565 1744 569 1821
rect 592 1779 596 1836
rect 600 1832 604 1836
rect 600 1824 618 1832
rect 614 1813 618 1824
rect 651 1824 655 1836
rect 669 1831 677 1837
rect 651 1812 653 1824
rect 585 1767 594 1779
rect 585 1744 589 1767
rect 614 1756 618 1801
rect 605 1749 618 1756
rect 605 1744 609 1749
rect 651 1744 655 1812
rect 673 1785 677 1831
rect 673 1724 677 1773
rect 701 1749 707 1844
rect 683 1745 707 1749
rect 683 1724 687 1745
rect 703 1740 721 1741
rect 703 1736 733 1740
rect 703 1724 707 1736
rect 741 1732 745 1858
rect 755 1850 759 1876
rect 775 1870 779 1876
rect 711 1728 745 1732
rect 711 1724 715 1728
rect 757 1724 761 1838
rect 773 1748 777 1858
rect 787 1836 791 1876
rect 782 1824 785 1836
rect 782 1760 786 1824
rect 807 1817 811 1876
rect 802 1809 811 1817
rect 802 1780 806 1809
rect 821 1794 825 1876
rect 841 1793 845 1836
rect 905 1833 909 1876
rect 925 1864 929 1876
rect 945 1868 949 1876
rect 945 1864 960 1868
rect 925 1860 940 1864
rect 934 1853 940 1860
rect 905 1821 913 1833
rect 925 1821 932 1833
rect 782 1756 815 1760
rect 781 1736 783 1748
rect 779 1724 783 1736
rect 789 1736 791 1748
rect 789 1724 793 1736
rect 811 1724 815 1756
rect 821 1724 825 1782
rect 841 1744 845 1781
rect 928 1764 932 1821
rect 936 1764 940 1841
rect 954 1833 960 1864
rect 944 1821 954 1833
rect 944 1764 948 1821
rect 991 1813 995 1876
rect 986 1801 995 1813
rect 991 1744 995 1801
rect 1013 1799 1017 1876
rect 1001 1787 1014 1799
rect 1001 1744 1005 1787
rect 1035 1762 1039 1836
rect 1091 1793 1095 1876
rect 1156 1832 1160 1836
rect 1142 1824 1160 1832
rect 1142 1813 1146 1824
rect 1086 1781 1095 1793
rect 1027 1750 1039 1762
rect 1021 1744 1025 1750
rect 1091 1724 1095 1781
rect 1142 1756 1146 1801
rect 1164 1779 1168 1836
rect 1186 1833 1190 1876
rect 1186 1821 1193 1833
rect 1166 1767 1175 1779
rect 1142 1749 1155 1756
rect 1151 1744 1155 1749
rect 1171 1744 1175 1767
rect 1191 1744 1195 1821
rect 1265 1799 1269 1876
rect 1266 1787 1269 1799
rect 1263 1771 1269 1787
rect 1285 1799 1289 1876
rect 1345 1833 1349 1876
rect 1365 1864 1369 1876
rect 1385 1868 1389 1876
rect 1385 1864 1400 1868
rect 1365 1860 1380 1864
rect 1374 1853 1380 1860
rect 1345 1821 1353 1833
rect 1365 1821 1372 1833
rect 1285 1787 1294 1799
rect 1285 1771 1291 1787
rect 1263 1764 1277 1771
rect 1273 1744 1277 1764
rect 1283 1764 1291 1771
rect 1368 1764 1372 1821
rect 1376 1764 1380 1841
rect 1394 1833 1400 1864
rect 1384 1821 1394 1833
rect 1384 1764 1388 1821
rect 1431 1793 1435 1876
rect 1495 1793 1499 1836
rect 1515 1794 1519 1876
rect 1529 1817 1533 1876
rect 1549 1836 1553 1876
rect 1561 1870 1565 1876
rect 1555 1824 1558 1836
rect 1529 1809 1538 1817
rect 1426 1781 1435 1793
rect 1283 1744 1287 1764
rect 1431 1724 1435 1781
rect 1495 1744 1499 1781
rect 1515 1724 1519 1782
rect 1534 1780 1538 1809
rect 1554 1760 1558 1824
rect 1525 1756 1558 1760
rect 1525 1724 1529 1756
rect 1563 1748 1567 1858
rect 1581 1850 1585 1876
rect 1627 1872 1631 1876
rect 1595 1870 1631 1872
rect 1607 1868 1631 1870
rect 1549 1736 1551 1748
rect 1547 1724 1551 1736
rect 1557 1736 1559 1748
rect 1557 1724 1561 1736
rect 1579 1724 1583 1838
rect 1595 1732 1599 1858
rect 1635 1844 1639 1876
rect 1655 1856 1659 1896
rect 1663 1873 1667 1896
rect 1663 1866 1671 1873
rect 1633 1749 1639 1844
rect 1667 1837 1671 1866
rect 1663 1831 1671 1837
rect 1663 1785 1667 1831
rect 1685 1824 1689 1836
rect 1687 1812 1689 1824
rect 1633 1745 1657 1749
rect 1619 1740 1637 1741
rect 1607 1736 1637 1740
rect 1595 1728 1629 1732
rect 1625 1724 1629 1728
rect 1633 1724 1637 1736
rect 1653 1724 1657 1745
rect 1663 1724 1667 1773
rect 1685 1744 1689 1812
rect 1731 1793 1735 1876
rect 1791 1832 1795 1836
rect 1781 1828 1795 1832
rect 1801 1832 1805 1836
rect 1801 1828 1815 1832
rect 1781 1813 1786 1828
rect 1726 1781 1735 1793
rect 1731 1724 1735 1781
rect 1780 1755 1786 1801
rect 1809 1779 1815 1828
rect 1831 1779 1835 1836
rect 1841 1832 1845 1836
rect 1841 1828 1855 1832
rect 1851 1813 1855 1828
rect 1911 1813 1915 1836
rect 1851 1801 1853 1813
rect 1906 1801 1915 1813
rect 1919 1813 1923 1836
rect 1996 1832 2000 1836
rect 1982 1824 2000 1832
rect 1982 1813 1986 1824
rect 1919 1801 1934 1813
rect 1806 1767 1815 1779
rect 1780 1751 1795 1755
rect 1791 1744 1795 1751
rect 1811 1744 1815 1767
rect 1831 1744 1835 1767
rect 1851 1744 1855 1801
rect 1911 1724 1915 1801
rect 1931 1724 1935 1801
rect 1982 1756 1986 1801
rect 2004 1779 2008 1836
rect 2026 1833 2030 1876
rect 2113 1873 2117 1896
rect 2109 1866 2117 1873
rect 2109 1837 2113 1866
rect 2121 1856 2125 1896
rect 2141 1844 2145 1876
rect 2149 1872 2153 1876
rect 2149 1870 2185 1872
rect 2149 1868 2173 1870
rect 2026 1821 2033 1833
rect 2091 1824 2095 1836
rect 2109 1831 2117 1837
rect 2006 1767 2015 1779
rect 1982 1749 1995 1756
rect 1991 1744 1995 1749
rect 2011 1744 2015 1767
rect 2031 1744 2035 1821
rect 2091 1812 2093 1824
rect 2091 1744 2095 1812
rect 2113 1785 2117 1831
rect 2113 1724 2117 1773
rect 2141 1749 2147 1844
rect 2123 1745 2147 1749
rect 2123 1724 2127 1745
rect 2143 1740 2161 1741
rect 2143 1736 2173 1740
rect 2143 1724 2147 1736
rect 2181 1732 2185 1858
rect 2195 1850 2199 1876
rect 2215 1870 2219 1876
rect 2151 1728 2185 1732
rect 2151 1724 2155 1728
rect 2197 1724 2201 1838
rect 2213 1748 2217 1858
rect 2227 1836 2231 1876
rect 2222 1824 2225 1836
rect 2222 1760 2226 1824
rect 2247 1817 2251 1876
rect 2242 1809 2251 1817
rect 2242 1780 2246 1809
rect 2261 1794 2265 1876
rect 2281 1793 2285 1836
rect 2355 1832 2359 1836
rect 2345 1828 2359 1832
rect 2345 1813 2349 1828
rect 2347 1801 2349 1813
rect 2222 1756 2255 1760
rect 2221 1736 2223 1748
rect 2219 1724 2223 1736
rect 2229 1736 2231 1748
rect 2229 1724 2233 1736
rect 2251 1724 2255 1756
rect 2261 1724 2265 1782
rect 2281 1744 2285 1781
rect 2345 1744 2349 1801
rect 2365 1779 2369 1836
rect 2395 1832 2399 1836
rect 2385 1828 2399 1832
rect 2405 1832 2409 1836
rect 2405 1828 2419 1832
rect 2385 1779 2391 1828
rect 2414 1813 2419 1828
rect 2385 1767 2394 1779
rect 2365 1744 2369 1767
rect 2385 1744 2389 1767
rect 2414 1755 2420 1801
rect 2451 1793 2455 1876
rect 2613 1873 2617 1896
rect 2609 1866 2617 1873
rect 2609 1837 2613 1866
rect 2621 1856 2625 1896
rect 2641 1844 2645 1876
rect 2649 1872 2653 1876
rect 2649 1870 2685 1872
rect 2649 1868 2673 1870
rect 2511 1813 2515 1836
rect 2506 1801 2515 1813
rect 2519 1813 2523 1836
rect 2591 1824 2595 1836
rect 2609 1831 2617 1837
rect 2519 1801 2534 1813
rect 2591 1812 2593 1824
rect 2446 1781 2455 1793
rect 2405 1751 2420 1755
rect 2405 1744 2409 1751
rect 2451 1724 2455 1781
rect 2511 1724 2515 1801
rect 2531 1724 2535 1801
rect 2591 1744 2595 1812
rect 2613 1785 2617 1831
rect 2613 1724 2617 1773
rect 2641 1749 2647 1844
rect 2623 1745 2647 1749
rect 2623 1724 2627 1745
rect 2643 1740 2661 1741
rect 2643 1736 2673 1740
rect 2643 1724 2647 1736
rect 2681 1732 2685 1858
rect 2695 1850 2699 1876
rect 2715 1870 2719 1876
rect 2651 1728 2685 1732
rect 2651 1724 2655 1728
rect 2697 1724 2701 1838
rect 2713 1748 2717 1858
rect 2727 1836 2731 1876
rect 2722 1824 2725 1836
rect 2722 1760 2726 1824
rect 2747 1817 2751 1876
rect 2742 1809 2751 1817
rect 2742 1780 2746 1809
rect 2761 1794 2765 1876
rect 2831 1868 2835 1876
rect 2820 1864 2835 1868
rect 2851 1864 2855 1876
rect 2781 1793 2785 1836
rect 2820 1833 2826 1864
rect 2840 1860 2855 1864
rect 2840 1853 2846 1860
rect 2826 1821 2836 1833
rect 2722 1756 2755 1760
rect 2721 1736 2723 1748
rect 2719 1724 2723 1736
rect 2729 1736 2731 1748
rect 2729 1724 2733 1736
rect 2751 1724 2755 1756
rect 2761 1724 2765 1782
rect 2781 1744 2785 1781
rect 2832 1764 2836 1821
rect 2840 1764 2844 1841
rect 2871 1833 2875 1876
rect 2950 1833 2954 1876
rect 2848 1821 2855 1833
rect 2867 1821 2875 1833
rect 2947 1821 2954 1833
rect 2848 1764 2852 1821
rect 2945 1744 2949 1821
rect 2972 1779 2976 1836
rect 2980 1832 2984 1836
rect 2980 1824 2998 1832
rect 2994 1813 2998 1824
rect 3031 1813 3035 1836
rect 3026 1801 3035 1813
rect 3039 1813 3043 1836
rect 3039 1801 3054 1813
rect 2965 1767 2974 1779
rect 2965 1744 2969 1767
rect 2994 1756 2998 1801
rect 2985 1749 2998 1756
rect 2985 1744 2989 1749
rect 3031 1724 3035 1801
rect 3051 1724 3055 1801
rect 3125 1779 3129 1836
rect 3145 1822 3149 1836
rect 3165 1822 3169 1836
rect 3145 1816 3160 1822
rect 3165 1816 3181 1822
rect 3154 1793 3160 1816
rect 3125 1767 3134 1779
rect 3132 1724 3136 1767
rect 3154 1744 3158 1781
rect 3174 1779 3181 1816
rect 3225 1779 3229 1836
rect 3245 1822 3249 1836
rect 3265 1822 3269 1836
rect 3323 1830 3327 1836
rect 3245 1816 3260 1822
rect 3265 1816 3281 1822
rect 3323 1818 3325 1830
rect 3254 1793 3260 1816
rect 3225 1767 3234 1779
rect 3174 1754 3181 1767
rect 3162 1748 3181 1754
rect 3162 1744 3166 1748
rect 3232 1724 3236 1767
rect 3254 1744 3258 1781
rect 3274 1779 3281 1816
rect 3345 1813 3349 1876
rect 3345 1801 3354 1813
rect 3274 1754 3281 1767
rect 3262 1748 3281 1754
rect 3323 1750 3325 1762
rect 3262 1744 3266 1748
rect 3323 1744 3327 1750
rect 3345 1724 3349 1801
rect 3405 1799 3409 1876
rect 3406 1787 3409 1799
rect 3403 1771 3409 1787
rect 3425 1799 3429 1876
rect 3471 1813 3475 1836
rect 3466 1801 3475 1813
rect 3479 1813 3483 1836
rect 3479 1801 3494 1813
rect 3425 1787 3434 1799
rect 3425 1771 3431 1787
rect 3403 1764 3417 1771
rect 3413 1744 3417 1764
rect 3423 1764 3431 1771
rect 3423 1744 3427 1764
rect 3471 1724 3475 1801
rect 3491 1724 3495 1801
rect 3551 1799 3555 1876
rect 3546 1787 3555 1799
rect 3549 1771 3555 1787
rect 3571 1799 3575 1876
rect 3636 1832 3640 1836
rect 3622 1824 3640 1832
rect 3622 1813 3626 1824
rect 3571 1787 3574 1799
rect 3571 1771 3577 1787
rect 3549 1764 3557 1771
rect 3553 1744 3557 1764
rect 3563 1764 3577 1771
rect 3563 1744 3567 1764
rect 3622 1756 3626 1801
rect 3644 1779 3648 1836
rect 3666 1833 3670 1876
rect 3666 1821 3673 1833
rect 3646 1767 3655 1779
rect 3622 1749 3635 1756
rect 3631 1744 3635 1749
rect 3651 1744 3655 1767
rect 3671 1744 3675 1821
rect 3745 1799 3749 1876
rect 3746 1787 3749 1799
rect 3743 1771 3749 1787
rect 3765 1799 3769 1876
rect 3765 1787 3774 1799
rect 3825 1793 3829 1876
rect 3871 1799 3875 1876
rect 3765 1771 3771 1787
rect 3743 1764 3757 1771
rect 3753 1744 3757 1764
rect 3763 1764 3771 1771
rect 3825 1781 3834 1793
rect 3866 1787 3875 1799
rect 3763 1744 3767 1764
rect 3825 1724 3829 1781
rect 3869 1771 3875 1787
rect 3891 1799 3895 1876
rect 3951 1813 3955 1836
rect 3946 1801 3955 1813
rect 3959 1813 3963 1836
rect 4031 1832 4035 1836
rect 4021 1828 4035 1832
rect 4041 1832 4045 1836
rect 4041 1828 4055 1832
rect 4021 1813 4026 1828
rect 3959 1801 3974 1813
rect 3891 1787 3894 1799
rect 3891 1771 3897 1787
rect 3869 1764 3877 1771
rect 3873 1744 3877 1764
rect 3883 1764 3897 1771
rect 3883 1744 3887 1764
rect 3951 1724 3955 1801
rect 3971 1724 3975 1801
rect 4020 1755 4026 1801
rect 4049 1779 4055 1828
rect 4071 1779 4075 1836
rect 4081 1832 4085 1836
rect 4081 1828 4095 1832
rect 4091 1813 4095 1828
rect 4177 1813 4181 1836
rect 4091 1801 4093 1813
rect 4166 1801 4181 1813
rect 4185 1813 4189 1836
rect 4236 1832 4240 1836
rect 4222 1824 4240 1832
rect 4222 1813 4226 1824
rect 4185 1801 4194 1813
rect 4046 1767 4055 1779
rect 4020 1751 4035 1755
rect 4031 1744 4035 1751
rect 4051 1744 4055 1767
rect 4071 1744 4075 1767
rect 4091 1744 4095 1801
rect 4165 1724 4169 1801
rect 4185 1724 4189 1801
rect 4222 1756 4226 1801
rect 4244 1779 4248 1836
rect 4266 1833 4270 1876
rect 4266 1821 4273 1833
rect 4331 1832 4335 1836
rect 4351 1832 4355 1836
rect 4416 1832 4420 1836
rect 4331 1828 4355 1832
rect 4246 1767 4255 1779
rect 4222 1749 4235 1756
rect 4231 1744 4235 1749
rect 4251 1744 4255 1767
rect 4271 1744 4275 1821
rect 4331 1779 4335 1828
rect 4402 1824 4420 1832
rect 4402 1813 4406 1824
rect 4326 1767 4335 1779
rect 4331 1752 4335 1767
rect 4402 1756 4406 1801
rect 4424 1779 4428 1836
rect 4446 1833 4450 1876
rect 4446 1821 4453 1833
rect 4426 1767 4435 1779
rect 4331 1748 4355 1752
rect 4402 1749 4415 1756
rect 4331 1744 4335 1748
rect 4351 1744 4355 1748
rect 4411 1744 4415 1749
rect 4431 1744 4435 1767
rect 4451 1744 4455 1821
rect 4537 1813 4541 1836
rect 4526 1801 4541 1813
rect 4545 1813 4549 1836
rect 4615 1832 4619 1836
rect 4605 1828 4619 1832
rect 4605 1813 4609 1828
rect 4545 1801 4554 1813
rect 4607 1801 4609 1813
rect 4525 1724 4529 1801
rect 4545 1724 4549 1801
rect 4605 1744 4609 1801
rect 4625 1779 4629 1836
rect 4655 1832 4659 1836
rect 4645 1828 4659 1832
rect 4665 1832 4669 1836
rect 4665 1828 4679 1832
rect 4645 1779 4651 1828
rect 4674 1813 4679 1828
rect 4645 1767 4654 1779
rect 4625 1744 4629 1767
rect 4645 1744 4649 1767
rect 4674 1755 4680 1801
rect 4665 1751 4680 1755
rect 4725 1793 4729 1876
rect 4793 1873 4797 1896
rect 4789 1866 4797 1873
rect 4789 1837 4793 1866
rect 4801 1856 4805 1896
rect 4821 1844 4825 1876
rect 4829 1872 4833 1876
rect 4829 1870 4865 1872
rect 4829 1868 4853 1870
rect 4771 1824 4775 1836
rect 4789 1831 4797 1837
rect 4771 1812 4773 1824
rect 4725 1781 4734 1793
rect 4665 1744 4669 1751
rect 4725 1724 4729 1781
rect 4771 1744 4775 1812
rect 4793 1785 4797 1831
rect 4793 1724 4797 1773
rect 4821 1749 4827 1844
rect 4803 1745 4827 1749
rect 4803 1724 4807 1745
rect 4823 1740 4841 1741
rect 4823 1736 4853 1740
rect 4823 1724 4827 1736
rect 4861 1732 4865 1858
rect 4875 1850 4879 1876
rect 4895 1870 4899 1876
rect 4831 1728 4865 1732
rect 4831 1724 4835 1728
rect 4877 1724 4881 1838
rect 4893 1748 4897 1858
rect 4907 1836 4911 1876
rect 4902 1824 4905 1836
rect 4902 1760 4906 1824
rect 4927 1817 4931 1876
rect 4922 1809 4931 1817
rect 4922 1780 4926 1809
rect 4941 1794 4945 1876
rect 4961 1793 4965 1836
rect 5011 1822 5015 1836
rect 5031 1822 5035 1836
rect 4999 1816 5015 1822
rect 5020 1816 5035 1822
rect 4902 1756 4935 1760
rect 4901 1736 4903 1748
rect 4899 1724 4903 1736
rect 4909 1736 4911 1748
rect 4909 1724 4913 1736
rect 4931 1724 4935 1756
rect 4941 1724 4945 1782
rect 4961 1744 4965 1781
rect 4999 1779 5006 1816
rect 5020 1793 5026 1816
rect 4999 1754 5006 1767
rect 4999 1748 5018 1754
rect 5014 1744 5018 1748
rect 5022 1744 5026 1781
rect 5051 1779 5055 1836
rect 5111 1813 5115 1836
rect 5106 1801 5115 1813
rect 5119 1813 5123 1836
rect 5196 1832 5200 1836
rect 5182 1824 5200 1832
rect 5182 1813 5186 1824
rect 5119 1801 5134 1813
rect 5046 1767 5055 1779
rect 5044 1724 5048 1767
rect 5111 1724 5115 1801
rect 5131 1724 5135 1801
rect 5182 1756 5186 1801
rect 5204 1779 5208 1836
rect 5226 1833 5230 1876
rect 5291 1868 5295 1876
rect 5280 1864 5295 1868
rect 5311 1864 5315 1876
rect 5280 1833 5286 1864
rect 5300 1860 5315 1864
rect 5300 1853 5306 1860
rect 5226 1821 5233 1833
rect 5286 1821 5296 1833
rect 5206 1767 5215 1779
rect 5182 1749 5195 1756
rect 5191 1744 5195 1749
rect 5211 1744 5215 1767
rect 5231 1744 5235 1821
rect 5292 1764 5296 1821
rect 5300 1764 5304 1841
rect 5331 1833 5335 1876
rect 5308 1821 5315 1833
rect 5327 1821 5335 1833
rect 5308 1764 5312 1821
rect 5391 1813 5395 1876
rect 5413 1830 5417 1836
rect 5415 1818 5417 1830
rect 5386 1801 5395 1813
rect 5391 1724 5395 1801
rect 5485 1793 5489 1876
rect 5485 1781 5494 1793
rect 5415 1750 5417 1762
rect 5413 1744 5417 1750
rect 5485 1724 5489 1781
rect 5545 1779 5549 1836
rect 5610 1833 5614 1876
rect 5607 1821 5614 1833
rect 5545 1767 5554 1779
rect 5545 1744 5549 1767
rect 5605 1744 5609 1821
rect 5632 1779 5636 1836
rect 5640 1832 5644 1836
rect 5640 1824 5658 1832
rect 5654 1813 5658 1824
rect 5625 1767 5634 1779
rect 5625 1744 5629 1767
rect 5654 1756 5658 1801
rect 5691 1799 5695 1876
rect 5686 1787 5695 1799
rect 5689 1771 5695 1787
rect 5711 1799 5715 1876
rect 5785 1813 5789 1836
rect 5786 1801 5789 1813
rect 5711 1787 5714 1799
rect 5711 1771 5717 1787
rect 5689 1764 5697 1771
rect 5645 1749 5658 1756
rect 5645 1744 5649 1749
rect 5693 1744 5697 1764
rect 5703 1764 5717 1771
rect 5703 1744 5707 1764
rect 5780 1753 5786 1801
rect 5805 1779 5809 1836
rect 5825 1814 5829 1836
rect 5845 1814 5849 1836
rect 5825 1808 5838 1814
rect 5845 1813 5865 1814
rect 5891 1813 5895 1876
rect 5913 1830 5917 1836
rect 5990 1833 5994 1876
rect 6191 1908 6195 1916
rect 6211 1908 6215 1912
rect 6221 1908 6225 1916
rect 6191 1864 6195 1868
rect 6183 1860 6195 1864
rect 5915 1818 5917 1830
rect 5987 1821 5994 1833
rect 5845 1808 5853 1813
rect 5834 1779 5838 1808
rect 5886 1801 5895 1813
rect 5807 1767 5809 1779
rect 5805 1765 5809 1767
rect 5805 1758 5818 1765
rect 5780 1749 5810 1753
rect 5806 1744 5810 1749
rect 5814 1744 5818 1758
rect 5834 1744 5838 1767
rect 5853 1759 5859 1801
rect 5842 1752 5859 1759
rect 5842 1744 5846 1752
rect 5891 1724 5895 1801
rect 5915 1750 5917 1762
rect 5913 1744 5917 1750
rect 5985 1744 5989 1821
rect 6012 1779 6016 1836
rect 6020 1832 6024 1836
rect 6095 1832 6099 1836
rect 6020 1824 6038 1832
rect 6034 1813 6038 1824
rect 6085 1828 6099 1832
rect 6085 1813 6089 1828
rect 6087 1801 6089 1813
rect 6005 1767 6014 1779
rect 6005 1744 6009 1767
rect 6034 1756 6038 1801
rect 6025 1749 6038 1756
rect 6025 1744 6029 1749
rect 6085 1744 6089 1801
rect 6105 1779 6109 1836
rect 6135 1832 6139 1836
rect 6125 1828 6139 1832
rect 6145 1832 6149 1836
rect 6145 1828 6159 1832
rect 6125 1779 6131 1828
rect 6154 1813 6159 1828
rect 6125 1767 6134 1779
rect 6105 1744 6109 1767
rect 6125 1744 6129 1767
rect 6154 1755 6160 1801
rect 6183 1779 6187 1860
rect 6311 1908 6315 1916
rect 6331 1908 6335 1912
rect 6341 1908 6345 1916
rect 6311 1864 6315 1868
rect 6303 1860 6315 1864
rect 6211 1823 6215 1828
rect 6221 1824 6225 1828
rect 6202 1819 6215 1823
rect 6202 1813 6207 1819
rect 6241 1814 6245 1836
rect 6215 1810 6245 1814
rect 6251 1813 6255 1836
rect 6145 1751 6160 1755
rect 6145 1744 6149 1751
rect 6183 1741 6187 1767
rect 6201 1770 6206 1801
rect 6251 1801 6254 1813
rect 6201 1764 6215 1770
rect 6211 1752 6215 1764
rect 6221 1752 6225 1798
rect 6241 1752 6245 1756
rect 6251 1752 6255 1801
rect 6303 1779 6307 1860
rect 6331 1823 6335 1828
rect 6341 1824 6345 1828
rect 6322 1819 6335 1823
rect 6322 1813 6327 1819
rect 6361 1814 6365 1836
rect 6335 1810 6365 1814
rect 6371 1813 6375 1836
rect 6183 1736 6195 1741
rect 6191 1732 6195 1736
rect 6303 1741 6307 1767
rect 6321 1770 6326 1801
rect 6371 1801 6374 1813
rect 6321 1764 6335 1770
rect 6331 1752 6335 1764
rect 6341 1752 6345 1798
rect 6361 1752 6365 1756
rect 6371 1752 6375 1801
rect 6431 1793 6435 1876
rect 6496 1832 6500 1836
rect 6482 1824 6500 1832
rect 6482 1813 6486 1824
rect 6426 1781 6435 1793
rect 6303 1736 6315 1741
rect 6311 1732 6315 1736
rect 6431 1724 6435 1781
rect 6482 1756 6486 1801
rect 6504 1779 6508 1836
rect 6526 1833 6530 1876
rect 6526 1821 6533 1833
rect 6506 1767 6515 1779
rect 6482 1749 6495 1756
rect 6491 1744 6495 1749
rect 6511 1744 6515 1767
rect 6531 1744 6535 1821
rect 6605 1799 6609 1876
rect 6606 1787 6609 1799
rect 6603 1771 6609 1787
rect 6625 1799 6629 1876
rect 6625 1787 6634 1799
rect 6625 1771 6631 1787
rect 6603 1764 6617 1771
rect 6613 1744 6617 1764
rect 6623 1764 6631 1771
rect 6623 1744 6627 1764
rect 6191 1704 6195 1712
rect 6211 1708 6215 1712
rect 6221 1708 6225 1712
rect 6241 1704 6245 1712
rect 6251 1708 6255 1712
rect 45 1700 49 1704
rect 91 1700 95 1704
rect 113 1700 117 1704
rect 123 1700 127 1704
rect 143 1700 147 1704
rect 151 1700 155 1704
rect 197 1700 201 1704
rect 219 1700 223 1704
rect 229 1700 233 1704
rect 251 1700 255 1704
rect 261 1700 265 1704
rect 281 1700 285 1704
rect 331 1700 335 1704
rect 351 1700 355 1704
rect 425 1700 429 1704
rect 445 1700 449 1704
rect 505 1700 509 1704
rect 565 1700 569 1704
rect 585 1700 589 1704
rect 605 1700 609 1704
rect 651 1700 655 1704
rect 673 1700 677 1704
rect 683 1700 687 1704
rect 703 1700 707 1704
rect 711 1700 715 1704
rect 757 1700 761 1704
rect 779 1700 783 1704
rect 789 1700 793 1704
rect 811 1700 815 1704
rect 821 1700 825 1704
rect 841 1700 845 1704
rect 928 1700 932 1704
rect 936 1700 940 1704
rect 944 1700 948 1704
rect 991 1700 995 1704
rect 1001 1700 1005 1704
rect 1021 1700 1025 1704
rect 1091 1700 1095 1704
rect 1151 1700 1155 1704
rect 1171 1700 1175 1704
rect 1191 1700 1195 1704
rect 1273 1700 1277 1704
rect 1283 1700 1287 1704
rect 1368 1700 1372 1704
rect 1376 1700 1380 1704
rect 1384 1700 1388 1704
rect 1431 1700 1435 1704
rect 1495 1700 1499 1704
rect 1515 1700 1519 1704
rect 1525 1700 1529 1704
rect 1547 1700 1551 1704
rect 1557 1700 1561 1704
rect 1579 1700 1583 1704
rect 1625 1700 1629 1704
rect 1633 1700 1637 1704
rect 1653 1700 1657 1704
rect 1663 1700 1667 1704
rect 1685 1700 1689 1704
rect 1731 1700 1735 1704
rect 1791 1700 1795 1704
rect 1811 1700 1815 1704
rect 1831 1700 1835 1704
rect 1851 1700 1855 1704
rect 1911 1700 1915 1704
rect 1931 1700 1935 1704
rect 1991 1700 1995 1704
rect 2011 1700 2015 1704
rect 2031 1700 2035 1704
rect 2091 1700 2095 1704
rect 2113 1700 2117 1704
rect 2123 1700 2127 1704
rect 2143 1700 2147 1704
rect 2151 1700 2155 1704
rect 2197 1700 2201 1704
rect 2219 1700 2223 1704
rect 2229 1700 2233 1704
rect 2251 1700 2255 1704
rect 2261 1700 2265 1704
rect 2281 1700 2285 1704
rect 2345 1700 2349 1704
rect 2365 1700 2369 1704
rect 2385 1700 2389 1704
rect 2405 1700 2409 1704
rect 2451 1700 2455 1704
rect 2511 1700 2515 1704
rect 2531 1700 2535 1704
rect 2591 1700 2595 1704
rect 2613 1700 2617 1704
rect 2623 1700 2627 1704
rect 2643 1700 2647 1704
rect 2651 1700 2655 1704
rect 2697 1700 2701 1704
rect 2719 1700 2723 1704
rect 2729 1700 2733 1704
rect 2751 1700 2755 1704
rect 2761 1700 2765 1704
rect 2781 1700 2785 1704
rect 2832 1700 2836 1704
rect 2840 1700 2844 1704
rect 2848 1700 2852 1704
rect 2945 1700 2949 1704
rect 2965 1700 2969 1704
rect 2985 1700 2989 1704
rect 3031 1700 3035 1704
rect 3051 1700 3055 1704
rect 3132 1700 3136 1704
rect 3154 1700 3158 1704
rect 3162 1700 3166 1704
rect 3232 1700 3236 1704
rect 3254 1700 3258 1704
rect 3262 1700 3266 1704
rect 3323 1700 3327 1704
rect 3345 1700 3349 1704
rect 3413 1700 3417 1704
rect 3423 1700 3427 1704
rect 3471 1700 3475 1704
rect 3491 1700 3495 1704
rect 3553 1700 3557 1704
rect 3563 1700 3567 1704
rect 3631 1700 3635 1704
rect 3651 1700 3655 1704
rect 3671 1700 3675 1704
rect 3753 1700 3757 1704
rect 3763 1700 3767 1704
rect 3825 1700 3829 1704
rect 3873 1700 3877 1704
rect 3883 1700 3887 1704
rect 3951 1700 3955 1704
rect 3971 1700 3975 1704
rect 4031 1700 4035 1704
rect 4051 1700 4055 1704
rect 4071 1700 4075 1704
rect 4091 1700 4095 1704
rect 4165 1700 4169 1704
rect 4185 1700 4189 1704
rect 4231 1700 4235 1704
rect 4251 1700 4255 1704
rect 4271 1700 4275 1704
rect 4331 1700 4335 1704
rect 4351 1700 4355 1704
rect 4411 1700 4415 1704
rect 4431 1700 4435 1704
rect 4451 1700 4455 1704
rect 4525 1700 4529 1704
rect 4545 1700 4549 1704
rect 4605 1700 4609 1704
rect 4625 1700 4629 1704
rect 4645 1700 4649 1704
rect 4665 1700 4669 1704
rect 4725 1700 4729 1704
rect 4771 1700 4775 1704
rect 4793 1700 4797 1704
rect 4803 1700 4807 1704
rect 4823 1700 4827 1704
rect 4831 1700 4835 1704
rect 4877 1700 4881 1704
rect 4899 1700 4903 1704
rect 4909 1700 4913 1704
rect 4931 1700 4935 1704
rect 4941 1700 4945 1704
rect 4961 1700 4965 1704
rect 5014 1700 5018 1704
rect 5022 1700 5026 1704
rect 5044 1700 5048 1704
rect 5111 1700 5115 1704
rect 5131 1700 5135 1704
rect 5191 1700 5195 1704
rect 5211 1700 5215 1704
rect 5231 1700 5235 1704
rect 5292 1700 5296 1704
rect 5300 1700 5304 1704
rect 5308 1700 5312 1704
rect 5391 1700 5395 1704
rect 5413 1700 5417 1704
rect 5485 1700 5489 1704
rect 5545 1700 5549 1704
rect 5605 1700 5609 1704
rect 5625 1700 5629 1704
rect 5645 1700 5649 1704
rect 5693 1700 5697 1704
rect 5703 1700 5707 1704
rect 5806 1700 5810 1704
rect 5814 1700 5818 1704
rect 5834 1700 5838 1704
rect 5842 1700 5846 1704
rect 5891 1700 5895 1704
rect 5913 1700 5917 1704
rect 5985 1700 5989 1704
rect 6005 1700 6009 1704
rect 6025 1700 6029 1704
rect 6085 1700 6089 1704
rect 6105 1700 6109 1704
rect 6125 1700 6129 1704
rect 6145 1700 6149 1704
rect 6191 1700 6245 1704
rect 6311 1704 6315 1712
rect 6331 1708 6335 1712
rect 6341 1708 6345 1712
rect 6361 1704 6365 1712
rect 6371 1708 6375 1712
rect 6311 1700 6365 1704
rect 6431 1700 6435 1704
rect 6491 1700 6495 1704
rect 6511 1700 6515 1704
rect 6531 1700 6535 1704
rect 6613 1700 6617 1704
rect 6623 1700 6627 1704
rect 45 1676 49 1680
rect 65 1676 69 1680
rect 125 1676 129 1680
rect 145 1676 149 1680
rect 165 1676 169 1680
rect 185 1676 189 1680
rect 205 1676 209 1680
rect 225 1676 229 1680
rect 245 1676 249 1680
rect 265 1676 269 1680
rect 315 1676 319 1680
rect 335 1676 339 1680
rect 345 1676 349 1680
rect 367 1676 371 1680
rect 377 1676 381 1680
rect 399 1676 403 1680
rect 445 1676 449 1680
rect 453 1676 457 1680
rect 473 1676 477 1680
rect 483 1676 487 1680
rect 505 1676 509 1680
rect 565 1676 569 1680
rect 612 1676 616 1680
rect 620 1676 624 1680
rect 628 1676 632 1680
rect 714 1676 718 1680
rect 722 1676 726 1680
rect 744 1676 748 1680
rect 815 1676 819 1680
rect 835 1676 839 1680
rect 845 1676 849 1680
rect 867 1676 871 1680
rect 877 1676 881 1680
rect 899 1676 903 1680
rect 945 1676 949 1680
rect 953 1676 957 1680
rect 973 1676 977 1680
rect 983 1676 987 1680
rect 1005 1676 1009 1680
rect 1065 1676 1069 1680
rect 1111 1676 1115 1680
rect 1131 1676 1135 1680
rect 1151 1676 1155 1680
rect 1171 1676 1175 1680
rect 1245 1676 1249 1680
rect 1265 1676 1269 1680
rect 1285 1676 1289 1680
rect 1345 1676 1349 1680
rect 1365 1676 1369 1680
rect 1435 1676 1489 1680
rect 45 1579 49 1656
rect 65 1579 69 1656
rect 125 1616 129 1636
rect 145 1616 149 1636
rect 165 1616 169 1636
rect 185 1616 189 1636
rect 205 1616 209 1636
rect 225 1616 229 1636
rect 125 1604 138 1616
rect 165 1604 178 1616
rect 205 1604 218 1616
rect 245 1613 249 1636
rect 265 1613 269 1636
rect 46 1567 61 1579
rect 57 1544 61 1567
rect 65 1567 74 1579
rect 65 1544 69 1567
rect 125 1544 129 1604
rect 145 1544 149 1604
rect 165 1544 169 1604
rect 185 1544 189 1604
rect 205 1544 209 1604
rect 225 1544 229 1604
rect 245 1601 254 1613
rect 266 1601 269 1613
rect 245 1544 249 1601
rect 265 1544 269 1601
rect 315 1599 319 1636
rect 335 1598 339 1656
rect 345 1624 349 1656
rect 367 1644 371 1656
rect 369 1632 371 1644
rect 377 1644 381 1656
rect 377 1632 379 1644
rect 345 1620 378 1624
rect 315 1544 319 1587
rect 335 1504 339 1586
rect 354 1571 358 1600
rect 349 1563 358 1571
rect 349 1504 353 1563
rect 374 1556 378 1620
rect 375 1544 378 1556
rect 369 1504 373 1544
rect 383 1522 387 1632
rect 399 1542 403 1656
rect 445 1652 449 1656
rect 415 1648 449 1652
rect 381 1504 385 1510
rect 401 1504 405 1530
rect 415 1522 419 1648
rect 453 1644 457 1656
rect 427 1640 457 1644
rect 439 1639 457 1640
rect 473 1635 477 1656
rect 453 1631 477 1635
rect 453 1536 459 1631
rect 483 1607 487 1656
rect 483 1549 487 1595
rect 505 1568 509 1636
rect 507 1556 509 1568
rect 483 1543 491 1549
rect 505 1544 509 1556
rect 565 1599 569 1656
rect 714 1632 718 1636
rect 699 1626 718 1632
rect 565 1587 574 1599
rect 427 1510 451 1512
rect 415 1508 451 1510
rect 447 1504 451 1508
rect 455 1504 459 1536
rect 475 1484 479 1524
rect 487 1514 491 1543
rect 483 1507 491 1514
rect 483 1484 487 1507
rect 565 1504 569 1587
rect 612 1559 616 1616
rect 606 1547 616 1559
rect 600 1516 606 1547
rect 620 1539 624 1616
rect 628 1559 632 1616
rect 699 1613 706 1626
rect 699 1564 706 1601
rect 722 1599 726 1636
rect 744 1613 748 1656
rect 746 1601 755 1613
rect 720 1564 726 1587
rect 628 1547 635 1559
rect 647 1547 655 1559
rect 699 1558 715 1564
rect 720 1558 735 1564
rect 620 1520 626 1527
rect 620 1516 635 1520
rect 600 1512 615 1516
rect 611 1504 615 1512
rect 631 1504 635 1516
rect 651 1504 655 1547
rect 711 1544 715 1558
rect 731 1544 735 1558
rect 751 1544 755 1601
rect 815 1599 819 1636
rect 835 1598 839 1656
rect 845 1624 849 1656
rect 867 1644 871 1656
rect 869 1632 871 1644
rect 877 1644 881 1656
rect 877 1632 879 1644
rect 845 1620 878 1624
rect 815 1544 819 1587
rect 835 1504 839 1586
rect 854 1571 858 1600
rect 849 1563 858 1571
rect 849 1504 853 1563
rect 874 1556 878 1620
rect 875 1544 878 1556
rect 869 1504 873 1544
rect 883 1522 887 1632
rect 899 1542 903 1656
rect 945 1652 949 1656
rect 915 1648 949 1652
rect 881 1504 885 1510
rect 901 1504 905 1530
rect 915 1522 919 1648
rect 953 1644 957 1656
rect 927 1640 957 1644
rect 939 1639 957 1640
rect 973 1635 977 1656
rect 953 1631 977 1635
rect 953 1536 959 1631
rect 983 1607 987 1656
rect 983 1549 987 1595
rect 1005 1568 1009 1636
rect 1007 1556 1009 1568
rect 983 1543 991 1549
rect 1005 1544 1009 1556
rect 1065 1599 1069 1656
rect 1425 1668 1429 1672
rect 1435 1668 1439 1676
rect 1455 1668 1459 1672
rect 1465 1668 1469 1672
rect 1485 1668 1489 1676
rect 1555 1676 1609 1680
rect 1545 1668 1549 1672
rect 1555 1668 1559 1676
rect 1575 1668 1579 1672
rect 1585 1668 1589 1672
rect 1605 1668 1609 1676
rect 1675 1676 1729 1680
rect 1771 1676 1775 1680
rect 1793 1676 1797 1680
rect 1803 1676 1807 1680
rect 1823 1676 1827 1680
rect 1831 1676 1835 1680
rect 1877 1676 1881 1680
rect 1899 1676 1903 1680
rect 1909 1676 1913 1680
rect 1931 1676 1935 1680
rect 1941 1676 1945 1680
rect 1961 1676 1965 1680
rect 2011 1676 2065 1680
rect 2131 1676 2135 1680
rect 2191 1676 2195 1680
rect 2211 1676 2215 1680
rect 2231 1676 2235 1680
rect 2251 1676 2255 1680
rect 2311 1676 2315 1680
rect 2331 1676 2335 1680
rect 2405 1676 2409 1680
rect 2425 1676 2429 1680
rect 2445 1676 2449 1680
rect 2503 1676 2507 1680
rect 2525 1676 2529 1680
rect 2571 1676 2575 1680
rect 2591 1676 2595 1680
rect 2673 1676 2677 1680
rect 2683 1676 2687 1680
rect 2733 1676 2737 1680
rect 2743 1676 2747 1680
rect 2835 1676 2889 1680
rect 2968 1676 2972 1680
rect 2976 1676 2980 1680
rect 2984 1676 2988 1680
rect 3045 1676 3049 1680
rect 3095 1676 3099 1680
rect 3115 1676 3119 1680
rect 3125 1676 3129 1680
rect 3147 1676 3151 1680
rect 3157 1676 3161 1680
rect 3179 1676 3183 1680
rect 3225 1676 3229 1680
rect 3233 1676 3237 1680
rect 3253 1676 3257 1680
rect 3263 1676 3267 1680
rect 3285 1676 3289 1680
rect 3353 1676 3357 1680
rect 3363 1676 3367 1680
rect 3425 1676 3429 1680
rect 3445 1676 3449 1680
rect 3465 1676 3469 1680
rect 3514 1676 3518 1680
rect 3522 1676 3526 1680
rect 3542 1676 3546 1680
rect 3550 1676 3554 1680
rect 3645 1676 3649 1680
rect 3665 1676 3669 1680
rect 3685 1676 3689 1680
rect 3745 1676 3749 1680
rect 3805 1676 3809 1680
rect 3825 1676 3829 1680
rect 3885 1676 3889 1680
rect 3905 1676 3909 1680
rect 3925 1676 3929 1680
rect 3945 1676 3949 1680
rect 4005 1676 4009 1680
rect 4055 1676 4059 1680
rect 4075 1676 4079 1680
rect 4085 1676 4089 1680
rect 4107 1676 4111 1680
rect 4117 1676 4121 1680
rect 4139 1676 4143 1680
rect 4185 1676 4189 1680
rect 4193 1676 4197 1680
rect 4213 1676 4217 1680
rect 4223 1676 4227 1680
rect 4245 1676 4249 1680
rect 4315 1676 4369 1680
rect 1665 1668 1669 1672
rect 1675 1668 1679 1676
rect 1695 1668 1699 1672
rect 1705 1668 1709 1672
rect 1725 1668 1729 1676
rect 1111 1629 1115 1636
rect 1100 1625 1115 1629
rect 1065 1587 1074 1599
rect 927 1510 951 1512
rect 915 1508 951 1510
rect 947 1504 951 1508
rect 955 1504 959 1536
rect 975 1484 979 1524
rect 987 1514 991 1543
rect 983 1507 991 1514
rect 983 1484 987 1507
rect 1065 1504 1069 1587
rect 1100 1579 1106 1625
rect 1131 1613 1135 1636
rect 1151 1613 1155 1636
rect 1126 1601 1135 1613
rect 1101 1552 1106 1567
rect 1129 1552 1135 1601
rect 1101 1548 1115 1552
rect 1111 1544 1115 1548
rect 1121 1548 1135 1552
rect 1121 1544 1125 1548
rect 1151 1544 1155 1601
rect 1171 1579 1175 1636
rect 1171 1567 1173 1579
rect 1171 1552 1175 1567
rect 1245 1559 1249 1636
rect 1265 1613 1269 1636
rect 1285 1631 1289 1636
rect 1285 1624 1298 1631
rect 1265 1601 1274 1613
rect 1161 1548 1175 1552
rect 1161 1544 1165 1548
rect 1247 1547 1254 1559
rect 1250 1504 1254 1547
rect 1272 1544 1276 1601
rect 1294 1579 1298 1624
rect 1345 1579 1349 1656
rect 1365 1579 1369 1656
rect 1485 1644 1489 1648
rect 1485 1639 1497 1644
rect 1425 1579 1429 1628
rect 1435 1624 1439 1628
rect 1455 1582 1459 1628
rect 1465 1616 1469 1628
rect 1465 1610 1479 1616
rect 1346 1567 1361 1579
rect 1294 1556 1298 1567
rect 1280 1548 1298 1556
rect 1280 1544 1284 1548
rect 1357 1544 1361 1567
rect 1365 1567 1374 1579
rect 1426 1567 1429 1579
rect 1474 1579 1479 1610
rect 1493 1613 1497 1639
rect 1605 1644 1609 1648
rect 1605 1639 1617 1644
rect 1365 1544 1369 1567
rect 1425 1544 1429 1567
rect 1435 1566 1465 1570
rect 1435 1544 1439 1566
rect 1473 1561 1478 1567
rect 1465 1557 1478 1561
rect 1455 1552 1459 1556
rect 1465 1552 1469 1557
rect 1493 1520 1497 1601
rect 1545 1579 1549 1628
rect 1555 1624 1559 1628
rect 1575 1582 1579 1628
rect 1585 1616 1589 1628
rect 1585 1610 1599 1616
rect 1546 1567 1549 1579
rect 1594 1579 1599 1610
rect 1613 1613 1617 1639
rect 1725 1644 1729 1648
rect 1725 1639 1737 1644
rect 1545 1544 1549 1567
rect 1555 1566 1585 1570
rect 1555 1544 1559 1566
rect 1593 1561 1598 1567
rect 1585 1557 1598 1561
rect 1575 1552 1579 1556
rect 1585 1552 1589 1557
rect 1485 1516 1497 1520
rect 1485 1512 1489 1516
rect 1455 1464 1459 1472
rect 1465 1468 1469 1472
rect 1485 1464 1489 1472
rect 1613 1520 1617 1601
rect 1665 1579 1669 1628
rect 1675 1624 1679 1628
rect 1695 1582 1699 1628
rect 1705 1616 1709 1628
rect 1705 1610 1719 1616
rect 1666 1567 1669 1579
rect 1714 1579 1719 1610
rect 1733 1613 1737 1639
rect 1665 1544 1669 1567
rect 1675 1566 1705 1570
rect 1675 1544 1679 1566
rect 1713 1561 1718 1567
rect 1705 1557 1718 1561
rect 1695 1552 1699 1556
rect 1705 1552 1709 1557
rect 1605 1516 1617 1520
rect 1605 1512 1609 1516
rect 1575 1464 1579 1472
rect 1585 1468 1589 1472
rect 1605 1464 1609 1472
rect 1733 1520 1737 1601
rect 1771 1568 1775 1636
rect 1793 1607 1797 1656
rect 1803 1635 1807 1656
rect 1823 1644 1827 1656
rect 1831 1652 1835 1656
rect 1831 1648 1865 1652
rect 1823 1640 1853 1644
rect 1823 1639 1841 1640
rect 1803 1631 1827 1635
rect 1771 1556 1773 1568
rect 1771 1544 1775 1556
rect 1793 1549 1797 1595
rect 1725 1516 1737 1520
rect 1725 1512 1729 1516
rect 1695 1464 1699 1472
rect 1705 1468 1709 1472
rect 1725 1464 1729 1472
rect 1789 1543 1797 1549
rect 1789 1514 1793 1543
rect 1821 1536 1827 1631
rect 1789 1507 1797 1514
rect 1793 1484 1797 1507
rect 1801 1484 1805 1524
rect 1821 1504 1825 1536
rect 1861 1522 1865 1648
rect 1877 1542 1881 1656
rect 1899 1644 1903 1656
rect 1901 1632 1903 1644
rect 1909 1644 1913 1656
rect 1909 1632 1911 1644
rect 1829 1510 1853 1512
rect 1829 1508 1865 1510
rect 1829 1504 1833 1508
rect 1875 1504 1879 1530
rect 1893 1522 1897 1632
rect 1931 1624 1935 1656
rect 1902 1620 1935 1624
rect 1902 1556 1906 1620
rect 1922 1571 1926 1600
rect 1941 1598 1945 1656
rect 2011 1668 2015 1676
rect 2031 1668 2035 1672
rect 2041 1668 2045 1672
rect 2061 1668 2065 1676
rect 2071 1668 2075 1672
rect 2011 1644 2015 1648
rect 2003 1639 2015 1644
rect 1961 1599 1965 1636
rect 2003 1613 2007 1639
rect 2031 1616 2035 1628
rect 1922 1563 1931 1571
rect 1902 1544 1905 1556
rect 1895 1504 1899 1510
rect 1907 1504 1911 1544
rect 1927 1504 1931 1563
rect 1941 1504 1945 1586
rect 1961 1544 1965 1587
rect 2003 1520 2007 1601
rect 2021 1610 2035 1616
rect 2021 1579 2026 1610
rect 2041 1582 2045 1628
rect 2061 1624 2065 1628
rect 2022 1561 2027 1567
rect 2071 1579 2075 1628
rect 2131 1599 2135 1656
rect 2191 1629 2195 1636
rect 2126 1587 2135 1599
rect 2035 1566 2065 1570
rect 2022 1557 2035 1561
rect 2031 1552 2035 1557
rect 2041 1552 2045 1556
rect 2003 1516 2015 1520
rect 2011 1512 2015 1516
rect 2061 1544 2065 1566
rect 2071 1567 2074 1579
rect 2071 1544 2075 1567
rect 2011 1464 2015 1472
rect 2031 1468 2035 1472
rect 2041 1464 2045 1472
rect 2131 1504 2135 1587
rect 2180 1625 2195 1629
rect 2180 1579 2186 1625
rect 2211 1613 2215 1636
rect 2231 1613 2235 1636
rect 2206 1601 2215 1613
rect 2181 1552 2186 1567
rect 2209 1552 2215 1601
rect 2181 1548 2195 1552
rect 2191 1544 2195 1548
rect 2201 1548 2215 1552
rect 2201 1544 2205 1548
rect 2231 1544 2235 1601
rect 2251 1579 2255 1636
rect 2311 1579 2315 1656
rect 2331 1579 2335 1656
rect 2251 1567 2253 1579
rect 2306 1567 2315 1579
rect 2251 1552 2255 1567
rect 2241 1548 2255 1552
rect 2241 1544 2245 1548
rect 2311 1544 2315 1567
rect 2319 1567 2334 1579
rect 2319 1544 2323 1567
rect 2405 1559 2409 1636
rect 2425 1613 2429 1636
rect 2445 1631 2449 1636
rect 2445 1624 2458 1631
rect 2425 1601 2434 1613
rect 2407 1547 2414 1559
rect 2410 1504 2414 1547
rect 2432 1544 2436 1601
rect 2454 1579 2458 1624
rect 2503 1630 2507 1636
rect 2503 1618 2505 1630
rect 2525 1579 2529 1656
rect 2571 1579 2575 1656
rect 2591 1579 2595 1656
rect 2825 1668 2829 1672
rect 2835 1668 2839 1676
rect 2855 1668 2859 1672
rect 2865 1668 2869 1672
rect 2885 1668 2889 1676
rect 2673 1616 2677 1636
rect 2663 1609 2677 1616
rect 2683 1616 2687 1636
rect 2733 1616 2737 1636
rect 2683 1609 2691 1616
rect 2663 1593 2669 1609
rect 2666 1581 2669 1593
rect 2525 1567 2534 1579
rect 2566 1567 2575 1579
rect 2454 1556 2458 1567
rect 2440 1548 2458 1556
rect 2503 1550 2505 1562
rect 2440 1544 2444 1548
rect 2503 1544 2507 1550
rect 2525 1504 2529 1567
rect 2571 1544 2575 1567
rect 2579 1567 2594 1579
rect 2579 1544 2583 1567
rect 2665 1504 2669 1581
rect 2685 1593 2691 1609
rect 2729 1609 2737 1616
rect 2743 1616 2747 1636
rect 2885 1644 2889 1648
rect 2885 1639 2897 1644
rect 2743 1609 2757 1616
rect 2729 1593 2735 1609
rect 2685 1581 2694 1593
rect 2726 1581 2735 1593
rect 2685 1504 2689 1581
rect 2731 1504 2735 1581
rect 2751 1593 2757 1609
rect 2751 1581 2754 1593
rect 2751 1504 2755 1581
rect 2825 1579 2829 1628
rect 2835 1624 2839 1628
rect 2855 1582 2859 1628
rect 2865 1616 2869 1628
rect 2865 1610 2879 1616
rect 2826 1567 2829 1579
rect 2874 1579 2879 1610
rect 2893 1613 2897 1639
rect 2825 1544 2829 1567
rect 2835 1566 2865 1570
rect 2835 1544 2839 1566
rect 2873 1561 2878 1567
rect 2865 1557 2878 1561
rect 2855 1552 2859 1556
rect 2865 1552 2869 1557
rect 2893 1520 2897 1601
rect 2968 1559 2972 1616
rect 2885 1516 2897 1520
rect 2945 1547 2953 1559
rect 2965 1547 2972 1559
rect 2885 1512 2889 1516
rect 2945 1504 2949 1547
rect 2976 1539 2980 1616
rect 2984 1559 2988 1616
rect 3045 1613 3049 1636
rect 3045 1601 3054 1613
rect 2984 1547 2994 1559
rect 2974 1520 2980 1527
rect 2965 1516 2980 1520
rect 2994 1516 3000 1547
rect 3045 1544 3049 1601
rect 3095 1599 3099 1636
rect 3115 1598 3119 1656
rect 3125 1624 3129 1656
rect 3147 1644 3151 1656
rect 3149 1632 3151 1644
rect 3157 1644 3161 1656
rect 3157 1632 3159 1644
rect 3125 1620 3158 1624
rect 3095 1544 3099 1587
rect 2965 1504 2969 1516
rect 2985 1512 3000 1516
rect 2985 1504 2989 1512
rect 2855 1464 2859 1472
rect 2865 1468 2869 1472
rect 2885 1464 2889 1472
rect 3115 1504 3119 1586
rect 3134 1571 3138 1600
rect 3129 1563 3138 1571
rect 3129 1504 3133 1563
rect 3154 1556 3158 1620
rect 3155 1544 3158 1556
rect 3149 1504 3153 1544
rect 3163 1522 3167 1632
rect 3179 1542 3183 1656
rect 3225 1652 3229 1656
rect 3195 1648 3229 1652
rect 3161 1504 3165 1510
rect 3181 1504 3185 1530
rect 3195 1522 3199 1648
rect 3233 1644 3237 1656
rect 3207 1640 3237 1644
rect 3219 1639 3237 1640
rect 3253 1635 3257 1656
rect 3233 1631 3257 1635
rect 3233 1536 3239 1631
rect 3263 1607 3267 1656
rect 3263 1549 3267 1595
rect 3285 1568 3289 1636
rect 3353 1616 3357 1636
rect 3343 1609 3357 1616
rect 3363 1616 3367 1636
rect 3363 1609 3371 1616
rect 3343 1593 3349 1609
rect 3346 1581 3349 1593
rect 3287 1556 3289 1568
rect 3263 1543 3271 1549
rect 3285 1544 3289 1556
rect 3207 1510 3231 1512
rect 3195 1508 3231 1510
rect 3227 1504 3231 1508
rect 3235 1504 3239 1536
rect 3255 1484 3259 1524
rect 3267 1514 3271 1543
rect 3263 1507 3271 1514
rect 3263 1484 3267 1507
rect 3345 1504 3349 1581
rect 3365 1593 3371 1609
rect 3365 1581 3374 1593
rect 3365 1504 3369 1581
rect 3425 1559 3429 1636
rect 3445 1613 3449 1636
rect 3465 1631 3469 1636
rect 3465 1624 3478 1631
rect 3514 1628 3518 1636
rect 3445 1601 3454 1613
rect 3427 1547 3434 1559
rect 3430 1504 3434 1547
rect 3452 1544 3456 1601
rect 3474 1579 3478 1624
rect 3501 1621 3518 1628
rect 3501 1579 3507 1621
rect 3522 1613 3526 1636
rect 3542 1622 3546 1636
rect 3550 1631 3554 1636
rect 3550 1627 3580 1631
rect 3542 1615 3555 1622
rect 3551 1613 3555 1615
rect 3551 1601 3553 1613
rect 3522 1572 3526 1601
rect 3507 1567 3515 1572
rect 3474 1556 3478 1567
rect 3495 1566 3515 1567
rect 3522 1566 3535 1572
rect 3460 1548 3478 1556
rect 3460 1544 3464 1548
rect 3511 1544 3515 1566
rect 3531 1544 3535 1566
rect 3551 1544 3555 1601
rect 3574 1579 3580 1627
rect 3571 1567 3574 1579
rect 3571 1544 3575 1567
rect 3645 1559 3649 1636
rect 3665 1613 3669 1636
rect 3685 1631 3689 1636
rect 3685 1624 3698 1631
rect 3665 1601 3674 1613
rect 3647 1547 3654 1559
rect 3650 1504 3654 1547
rect 3672 1544 3676 1601
rect 3694 1579 3698 1624
rect 3745 1599 3749 1656
rect 3745 1587 3754 1599
rect 3694 1556 3698 1567
rect 3680 1548 3698 1556
rect 3680 1544 3684 1548
rect 3745 1504 3749 1587
rect 3805 1579 3809 1656
rect 3825 1579 3829 1656
rect 3885 1579 3889 1636
rect 3905 1613 3909 1636
rect 3925 1613 3929 1636
rect 3945 1629 3949 1636
rect 3945 1625 3960 1629
rect 3925 1601 3934 1613
rect 3806 1567 3821 1579
rect 3817 1544 3821 1567
rect 3825 1567 3834 1579
rect 3887 1567 3889 1579
rect 3825 1544 3829 1567
rect 3885 1552 3889 1567
rect 3885 1548 3899 1552
rect 3895 1544 3899 1548
rect 3905 1544 3909 1601
rect 3925 1552 3931 1601
rect 3954 1579 3960 1625
rect 4005 1599 4009 1656
rect 4055 1599 4059 1636
rect 4005 1587 4014 1599
rect 4075 1598 4079 1656
rect 4085 1624 4089 1656
rect 4107 1644 4111 1656
rect 4109 1632 4111 1644
rect 4117 1644 4121 1656
rect 4117 1632 4119 1644
rect 4085 1620 4118 1624
rect 3954 1552 3959 1567
rect 3925 1548 3939 1552
rect 3935 1544 3939 1548
rect 3945 1548 3959 1552
rect 3945 1544 3949 1548
rect 4005 1504 4009 1587
rect 4055 1544 4059 1587
rect 4075 1504 4079 1586
rect 4094 1571 4098 1600
rect 4089 1563 4098 1571
rect 4089 1504 4093 1563
rect 4114 1556 4118 1620
rect 4115 1544 4118 1556
rect 4109 1504 4113 1544
rect 4123 1522 4127 1632
rect 4139 1542 4143 1656
rect 4185 1652 4189 1656
rect 4155 1648 4189 1652
rect 4121 1504 4125 1510
rect 4141 1504 4145 1530
rect 4155 1522 4159 1648
rect 4193 1644 4197 1656
rect 4167 1640 4197 1644
rect 4179 1639 4197 1640
rect 4213 1635 4217 1656
rect 4193 1631 4217 1635
rect 4193 1536 4199 1631
rect 4223 1607 4227 1656
rect 4305 1668 4309 1672
rect 4315 1668 4319 1676
rect 4335 1668 4339 1672
rect 4345 1668 4349 1672
rect 4365 1668 4369 1676
rect 4435 1676 4489 1680
rect 4425 1668 4429 1672
rect 4435 1668 4439 1676
rect 4455 1668 4459 1672
rect 4465 1668 4469 1672
rect 4485 1668 4489 1676
rect 4531 1676 4585 1680
rect 4531 1668 4535 1676
rect 4551 1668 4555 1672
rect 4561 1668 4565 1672
rect 4581 1668 4585 1676
rect 4651 1676 4705 1680
rect 4591 1668 4595 1672
rect 4651 1668 4655 1676
rect 4671 1668 4675 1672
rect 4681 1668 4685 1672
rect 4701 1668 4705 1676
rect 4771 1676 4825 1680
rect 4711 1668 4715 1672
rect 4771 1668 4775 1676
rect 4791 1668 4795 1672
rect 4801 1668 4805 1672
rect 4821 1668 4825 1676
rect 4891 1676 4945 1680
rect 5011 1676 5015 1680
rect 5033 1676 5037 1680
rect 5043 1676 5047 1680
rect 5063 1676 5067 1680
rect 5071 1676 5075 1680
rect 5117 1676 5121 1680
rect 5139 1676 5143 1680
rect 5149 1676 5153 1680
rect 5171 1676 5175 1680
rect 5181 1676 5185 1680
rect 5201 1676 5205 1680
rect 5251 1676 5255 1680
rect 5273 1676 5277 1680
rect 5283 1676 5287 1680
rect 5303 1676 5307 1680
rect 5311 1676 5315 1680
rect 5357 1676 5361 1680
rect 5379 1676 5383 1680
rect 5389 1676 5393 1680
rect 5411 1676 5415 1680
rect 5421 1676 5425 1680
rect 5441 1676 5445 1680
rect 5494 1676 5498 1680
rect 5502 1676 5506 1680
rect 5522 1676 5526 1680
rect 5530 1676 5534 1680
rect 5611 1676 5665 1680
rect 5745 1676 5749 1680
rect 5765 1676 5769 1680
rect 5785 1676 5789 1680
rect 5845 1676 5849 1680
rect 5865 1676 5869 1680
rect 5933 1676 5937 1680
rect 5943 1676 5947 1680
rect 6005 1676 6009 1680
rect 6025 1676 6029 1680
rect 6045 1676 6049 1680
rect 6105 1676 6109 1680
rect 6125 1676 6129 1680
rect 6185 1676 6189 1680
rect 6205 1676 6209 1680
rect 6225 1676 6229 1680
rect 6245 1676 6249 1680
rect 6315 1676 6369 1680
rect 6411 1676 6415 1680
rect 6471 1676 6475 1680
rect 6493 1676 6497 1680
rect 6503 1676 6507 1680
rect 6523 1676 6527 1680
rect 6531 1676 6535 1680
rect 6577 1676 6581 1680
rect 6599 1676 6603 1680
rect 6609 1676 6613 1680
rect 6631 1676 6635 1680
rect 6641 1676 6645 1680
rect 6661 1676 6665 1680
rect 4831 1668 4835 1672
rect 4891 1668 4895 1676
rect 4911 1668 4915 1672
rect 4921 1668 4925 1672
rect 4941 1668 4945 1676
rect 4951 1668 4955 1672
rect 4223 1549 4227 1595
rect 4245 1568 4249 1636
rect 4365 1644 4369 1648
rect 4365 1639 4377 1644
rect 4305 1579 4309 1628
rect 4315 1624 4319 1628
rect 4335 1582 4339 1628
rect 4345 1616 4349 1628
rect 4345 1610 4359 1616
rect 4247 1556 4249 1568
rect 4306 1567 4309 1579
rect 4354 1579 4359 1610
rect 4373 1613 4377 1639
rect 4485 1644 4489 1648
rect 4531 1644 4535 1648
rect 4485 1639 4497 1644
rect 4223 1543 4231 1549
rect 4245 1544 4249 1556
rect 4305 1544 4309 1567
rect 4315 1566 4345 1570
rect 4315 1544 4319 1566
rect 4353 1561 4358 1567
rect 4345 1557 4358 1561
rect 4335 1552 4339 1556
rect 4345 1552 4349 1557
rect 4167 1510 4191 1512
rect 4155 1508 4191 1510
rect 4187 1504 4191 1508
rect 4195 1504 4199 1536
rect 4215 1484 4219 1524
rect 4227 1514 4231 1543
rect 4223 1507 4231 1514
rect 4223 1484 4227 1507
rect 4373 1520 4377 1601
rect 4425 1579 4429 1628
rect 4435 1624 4439 1628
rect 4455 1582 4459 1628
rect 4465 1616 4469 1628
rect 4465 1610 4479 1616
rect 4426 1567 4429 1579
rect 4474 1579 4479 1610
rect 4493 1613 4497 1639
rect 4523 1639 4535 1644
rect 4523 1613 4527 1639
rect 4651 1644 4655 1648
rect 4643 1639 4655 1644
rect 4551 1616 4555 1628
rect 4425 1544 4429 1567
rect 4435 1566 4465 1570
rect 4435 1544 4439 1566
rect 4473 1561 4478 1567
rect 4465 1557 4478 1561
rect 4455 1552 4459 1556
rect 4465 1552 4469 1557
rect 4365 1516 4377 1520
rect 4365 1512 4369 1516
rect 4335 1464 4339 1472
rect 4345 1468 4349 1472
rect 4365 1464 4369 1472
rect 4493 1520 4497 1601
rect 4485 1516 4497 1520
rect 4523 1520 4527 1601
rect 4541 1610 4555 1616
rect 4541 1579 4546 1610
rect 4561 1582 4565 1628
rect 4581 1624 4585 1628
rect 4542 1561 4547 1567
rect 4591 1579 4595 1628
rect 4643 1613 4647 1639
rect 4771 1644 4775 1648
rect 4763 1639 4775 1644
rect 4671 1616 4675 1628
rect 4555 1566 4585 1570
rect 4542 1557 4555 1561
rect 4551 1552 4555 1557
rect 4561 1552 4565 1556
rect 4523 1516 4535 1520
rect 4485 1512 4489 1516
rect 4531 1512 4535 1516
rect 4581 1544 4585 1566
rect 4591 1567 4594 1579
rect 4591 1544 4595 1567
rect 4455 1464 4459 1472
rect 4465 1468 4469 1472
rect 4485 1464 4489 1472
rect 57 1460 61 1464
rect 65 1460 69 1464
rect 125 1460 129 1464
rect 145 1460 149 1464
rect 165 1460 169 1464
rect 185 1460 189 1464
rect 205 1460 209 1464
rect 225 1460 229 1464
rect 245 1460 249 1464
rect 265 1460 269 1464
rect 315 1460 319 1464
rect 335 1460 339 1464
rect 349 1460 353 1464
rect 369 1460 373 1464
rect 381 1460 385 1464
rect 401 1460 405 1464
rect 447 1460 451 1464
rect 455 1460 459 1464
rect 475 1460 479 1464
rect 483 1460 487 1464
rect 505 1460 509 1464
rect 565 1460 569 1464
rect 611 1460 615 1464
rect 631 1460 635 1464
rect 651 1460 655 1464
rect 711 1460 715 1464
rect 731 1460 735 1464
rect 751 1460 755 1464
rect 815 1460 819 1464
rect 835 1460 839 1464
rect 849 1460 853 1464
rect 869 1460 873 1464
rect 881 1460 885 1464
rect 901 1460 905 1464
rect 947 1460 951 1464
rect 955 1460 959 1464
rect 975 1460 979 1464
rect 983 1460 987 1464
rect 1005 1460 1009 1464
rect 1065 1460 1069 1464
rect 1111 1460 1115 1464
rect 1121 1460 1125 1464
rect 1151 1460 1155 1464
rect 1161 1460 1165 1464
rect 1250 1460 1254 1464
rect 1272 1460 1276 1464
rect 1280 1460 1284 1464
rect 1357 1460 1361 1464
rect 1365 1460 1369 1464
rect 1425 1460 1429 1464
rect 1435 1460 1439 1464
rect 1455 1460 1489 1464
rect 1545 1460 1549 1464
rect 1555 1460 1559 1464
rect 1575 1460 1609 1464
rect 1665 1460 1669 1464
rect 1675 1460 1679 1464
rect 1695 1460 1729 1464
rect 1771 1460 1775 1464
rect 1793 1460 1797 1464
rect 1801 1460 1805 1464
rect 1821 1460 1825 1464
rect 1829 1460 1833 1464
rect 1875 1460 1879 1464
rect 1895 1460 1899 1464
rect 1907 1460 1911 1464
rect 1927 1460 1931 1464
rect 1941 1460 1945 1464
rect 1961 1460 1965 1464
rect 2011 1460 2045 1464
rect 2061 1460 2065 1464
rect 2071 1460 2075 1464
rect 2131 1460 2135 1464
rect 2191 1460 2195 1464
rect 2201 1460 2205 1464
rect 2231 1460 2235 1464
rect 2241 1460 2245 1464
rect 2311 1460 2315 1464
rect 2319 1460 2323 1464
rect 2410 1460 2414 1464
rect 2432 1460 2436 1464
rect 2440 1460 2444 1464
rect 2503 1460 2507 1464
rect 2525 1460 2529 1464
rect 2571 1460 2575 1464
rect 2579 1460 2583 1464
rect 2665 1460 2669 1464
rect 2685 1460 2689 1464
rect 2731 1460 2735 1464
rect 2751 1460 2755 1464
rect 2825 1460 2829 1464
rect 2835 1460 2839 1464
rect 2855 1460 2889 1464
rect 2945 1460 2949 1464
rect 2965 1460 2969 1464
rect 2985 1460 2989 1464
rect 3045 1460 3049 1464
rect 3095 1460 3099 1464
rect 3115 1460 3119 1464
rect 3129 1460 3133 1464
rect 3149 1460 3153 1464
rect 3161 1460 3165 1464
rect 3181 1460 3185 1464
rect 3227 1460 3231 1464
rect 3235 1460 3239 1464
rect 3255 1460 3259 1464
rect 3263 1460 3267 1464
rect 3285 1460 3289 1464
rect 3345 1460 3349 1464
rect 3365 1460 3369 1464
rect 3430 1460 3434 1464
rect 3452 1460 3456 1464
rect 3460 1460 3464 1464
rect 3511 1460 3515 1464
rect 3531 1460 3535 1464
rect 3551 1460 3555 1464
rect 3571 1460 3575 1464
rect 3650 1460 3654 1464
rect 3672 1460 3676 1464
rect 3680 1460 3684 1464
rect 3745 1460 3749 1464
rect 3817 1460 3821 1464
rect 3825 1460 3829 1464
rect 3895 1460 3899 1464
rect 3905 1460 3909 1464
rect 3935 1460 3939 1464
rect 3945 1460 3949 1464
rect 4005 1460 4009 1464
rect 4055 1460 4059 1464
rect 4075 1460 4079 1464
rect 4089 1460 4093 1464
rect 4109 1460 4113 1464
rect 4121 1460 4125 1464
rect 4141 1460 4145 1464
rect 4187 1460 4191 1464
rect 4195 1460 4199 1464
rect 4215 1460 4219 1464
rect 4223 1460 4227 1464
rect 4245 1460 4249 1464
rect 4305 1460 4309 1464
rect 4315 1460 4319 1464
rect 4335 1460 4369 1464
rect 4425 1460 4429 1464
rect 4435 1460 4439 1464
rect 4455 1460 4489 1464
rect 4531 1464 4535 1472
rect 4551 1468 4555 1472
rect 4561 1464 4565 1472
rect 4643 1520 4647 1601
rect 4661 1610 4675 1616
rect 4661 1579 4666 1610
rect 4681 1582 4685 1628
rect 4701 1624 4705 1628
rect 4662 1561 4667 1567
rect 4711 1579 4715 1628
rect 4763 1613 4767 1639
rect 4891 1644 4895 1648
rect 4883 1639 4895 1644
rect 4791 1616 4795 1628
rect 4675 1566 4705 1570
rect 4662 1557 4675 1561
rect 4671 1552 4675 1557
rect 4681 1552 4685 1556
rect 4643 1516 4655 1520
rect 4651 1512 4655 1516
rect 4701 1544 4705 1566
rect 4711 1567 4714 1579
rect 4711 1544 4715 1567
rect 4651 1464 4655 1472
rect 4671 1468 4675 1472
rect 4681 1464 4685 1472
rect 4763 1520 4767 1601
rect 4781 1610 4795 1616
rect 4781 1579 4786 1610
rect 4801 1582 4805 1628
rect 4821 1624 4825 1628
rect 4782 1561 4787 1567
rect 4831 1579 4835 1628
rect 4883 1613 4887 1639
rect 4911 1616 4915 1628
rect 4795 1566 4825 1570
rect 4782 1557 4795 1561
rect 4791 1552 4795 1557
rect 4801 1552 4805 1556
rect 4763 1516 4775 1520
rect 4771 1512 4775 1516
rect 4821 1544 4825 1566
rect 4831 1567 4834 1579
rect 4831 1544 4835 1567
rect 4771 1464 4775 1472
rect 4791 1468 4795 1472
rect 4801 1464 4805 1472
rect 4883 1520 4887 1601
rect 4901 1610 4915 1616
rect 4901 1579 4906 1610
rect 4921 1582 4925 1628
rect 4941 1624 4945 1628
rect 4902 1561 4907 1567
rect 4951 1579 4955 1628
rect 4915 1566 4945 1570
rect 4902 1557 4915 1561
rect 4911 1552 4915 1557
rect 4921 1552 4925 1556
rect 4883 1516 4895 1520
rect 4891 1512 4895 1516
rect 4941 1544 4945 1566
rect 4951 1567 4954 1579
rect 5011 1568 5015 1636
rect 5033 1607 5037 1656
rect 5043 1635 5047 1656
rect 5063 1644 5067 1656
rect 5071 1652 5075 1656
rect 5071 1648 5105 1652
rect 5063 1640 5093 1644
rect 5063 1639 5081 1640
rect 5043 1631 5067 1635
rect 4951 1544 4955 1567
rect 5011 1556 5013 1568
rect 5011 1544 5015 1556
rect 5033 1549 5037 1595
rect 4891 1464 4895 1472
rect 4911 1468 4915 1472
rect 4921 1464 4925 1472
rect 5029 1543 5037 1549
rect 5029 1514 5033 1543
rect 5061 1536 5067 1631
rect 5029 1507 5037 1514
rect 5033 1484 5037 1507
rect 5041 1484 5045 1524
rect 5061 1504 5065 1536
rect 5101 1522 5105 1648
rect 5117 1542 5121 1656
rect 5139 1644 5143 1656
rect 5141 1632 5143 1644
rect 5149 1644 5153 1656
rect 5149 1632 5151 1644
rect 5069 1510 5093 1512
rect 5069 1508 5105 1510
rect 5069 1504 5073 1508
rect 5115 1504 5119 1530
rect 5133 1522 5137 1632
rect 5171 1624 5175 1656
rect 5142 1620 5175 1624
rect 5142 1556 5146 1620
rect 5162 1571 5166 1600
rect 5181 1598 5185 1656
rect 5201 1599 5205 1636
rect 5162 1563 5171 1571
rect 5142 1544 5145 1556
rect 5135 1504 5139 1510
rect 5147 1504 5151 1544
rect 5167 1504 5171 1563
rect 5181 1504 5185 1586
rect 5201 1544 5205 1587
rect 5251 1568 5255 1636
rect 5273 1607 5277 1656
rect 5283 1635 5287 1656
rect 5303 1644 5307 1656
rect 5311 1652 5315 1656
rect 5311 1648 5345 1652
rect 5303 1640 5333 1644
rect 5303 1639 5321 1640
rect 5283 1631 5307 1635
rect 5251 1556 5253 1568
rect 5251 1544 5255 1556
rect 5273 1549 5277 1595
rect 5269 1543 5277 1549
rect 5269 1514 5273 1543
rect 5301 1536 5307 1631
rect 5269 1507 5277 1514
rect 5273 1484 5277 1507
rect 5281 1484 5285 1524
rect 5301 1504 5305 1536
rect 5341 1522 5345 1648
rect 5357 1542 5361 1656
rect 5379 1644 5383 1656
rect 5381 1632 5383 1644
rect 5389 1644 5393 1656
rect 5389 1632 5391 1644
rect 5309 1510 5333 1512
rect 5309 1508 5345 1510
rect 5309 1504 5313 1508
rect 5355 1504 5359 1530
rect 5373 1522 5377 1632
rect 5411 1624 5415 1656
rect 5382 1620 5415 1624
rect 5382 1556 5386 1620
rect 5402 1571 5406 1600
rect 5421 1598 5425 1656
rect 5611 1668 5615 1676
rect 5631 1668 5635 1672
rect 5641 1668 5645 1672
rect 5661 1668 5665 1676
rect 5671 1668 5675 1672
rect 5611 1644 5615 1648
rect 5603 1639 5615 1644
rect 5441 1599 5445 1636
rect 5494 1628 5498 1636
rect 5481 1621 5498 1628
rect 5402 1563 5411 1571
rect 5382 1544 5385 1556
rect 5375 1504 5379 1510
rect 5387 1504 5391 1544
rect 5407 1504 5411 1563
rect 5421 1504 5425 1586
rect 5441 1544 5445 1587
rect 5481 1579 5487 1621
rect 5502 1613 5506 1636
rect 5522 1622 5526 1636
rect 5530 1631 5534 1636
rect 5530 1627 5560 1631
rect 5522 1615 5535 1622
rect 5531 1613 5535 1615
rect 5531 1601 5533 1613
rect 5502 1572 5506 1601
rect 5487 1567 5495 1572
rect 5475 1566 5495 1567
rect 5502 1566 5515 1572
rect 5491 1544 5495 1566
rect 5511 1544 5515 1566
rect 5531 1544 5535 1601
rect 5554 1579 5560 1627
rect 5603 1613 5607 1639
rect 5631 1616 5635 1628
rect 5551 1567 5554 1579
rect 5551 1544 5555 1567
rect 5603 1520 5607 1601
rect 5621 1610 5635 1616
rect 5621 1579 5626 1610
rect 5641 1582 5645 1628
rect 5661 1624 5665 1628
rect 5622 1561 5627 1567
rect 5671 1579 5675 1628
rect 5635 1566 5665 1570
rect 5622 1557 5635 1561
rect 5631 1552 5635 1557
rect 5641 1552 5645 1556
rect 5603 1516 5615 1520
rect 5611 1512 5615 1516
rect 5661 1544 5665 1566
rect 5671 1567 5674 1579
rect 5671 1544 5675 1567
rect 5745 1559 5749 1636
rect 5765 1613 5769 1636
rect 5785 1631 5789 1636
rect 5785 1624 5798 1631
rect 5765 1601 5774 1613
rect 5747 1547 5754 1559
rect 5611 1464 5615 1472
rect 5631 1468 5635 1472
rect 5641 1464 5645 1472
rect 5750 1504 5754 1547
rect 5772 1544 5776 1601
rect 5794 1579 5798 1624
rect 5845 1579 5849 1656
rect 5865 1579 5869 1656
rect 5933 1616 5937 1636
rect 5923 1609 5937 1616
rect 5943 1616 5947 1636
rect 5943 1609 5951 1616
rect 5923 1593 5929 1609
rect 5926 1581 5929 1593
rect 5846 1567 5861 1579
rect 5794 1556 5798 1567
rect 5780 1548 5798 1556
rect 5780 1544 5784 1548
rect 5857 1544 5861 1567
rect 5865 1567 5874 1579
rect 5865 1544 5869 1567
rect 5925 1504 5929 1581
rect 5945 1593 5951 1609
rect 5945 1581 5954 1593
rect 5945 1504 5949 1581
rect 6005 1559 6009 1636
rect 6025 1613 6029 1636
rect 6045 1631 6049 1636
rect 6045 1624 6058 1631
rect 6025 1601 6034 1613
rect 6007 1547 6014 1559
rect 6010 1504 6014 1547
rect 6032 1544 6036 1601
rect 6054 1579 6058 1624
rect 6105 1579 6109 1656
rect 6125 1579 6129 1656
rect 6305 1668 6309 1672
rect 6315 1668 6319 1676
rect 6335 1668 6339 1672
rect 6345 1668 6349 1672
rect 6365 1668 6369 1676
rect 6185 1579 6189 1636
rect 6205 1613 6209 1636
rect 6225 1613 6229 1636
rect 6245 1629 6249 1636
rect 6245 1625 6260 1629
rect 6365 1644 6369 1648
rect 6365 1639 6377 1644
rect 6225 1601 6234 1613
rect 6106 1567 6121 1579
rect 6054 1556 6058 1567
rect 6040 1548 6058 1556
rect 6040 1544 6044 1548
rect 6117 1544 6121 1567
rect 6125 1567 6134 1579
rect 6187 1567 6189 1579
rect 6125 1544 6129 1567
rect 6185 1552 6189 1567
rect 6185 1548 6199 1552
rect 6195 1544 6199 1548
rect 6205 1544 6209 1601
rect 6225 1552 6231 1601
rect 6254 1579 6260 1625
rect 6305 1579 6309 1628
rect 6315 1624 6319 1628
rect 6335 1582 6339 1628
rect 6345 1616 6349 1628
rect 6345 1610 6359 1616
rect 6306 1567 6309 1579
rect 6354 1579 6359 1610
rect 6373 1613 6377 1639
rect 6254 1552 6259 1567
rect 6225 1548 6239 1552
rect 6235 1544 6239 1548
rect 6245 1548 6259 1552
rect 6245 1544 6249 1548
rect 6305 1544 6309 1567
rect 6315 1566 6345 1570
rect 6315 1544 6319 1566
rect 6353 1561 6358 1567
rect 6345 1557 6358 1561
rect 6335 1552 6339 1556
rect 6345 1552 6349 1557
rect 6373 1520 6377 1601
rect 6411 1599 6415 1656
rect 6406 1587 6415 1599
rect 6365 1516 6377 1520
rect 6365 1512 6369 1516
rect 6411 1504 6415 1587
rect 6471 1568 6475 1636
rect 6493 1607 6497 1656
rect 6503 1635 6507 1656
rect 6523 1644 6527 1656
rect 6531 1652 6535 1656
rect 6531 1648 6565 1652
rect 6523 1640 6553 1644
rect 6523 1639 6541 1640
rect 6503 1631 6527 1635
rect 6471 1556 6473 1568
rect 6471 1544 6475 1556
rect 6493 1549 6497 1595
rect 6335 1464 6339 1472
rect 6345 1468 6349 1472
rect 6365 1464 6369 1472
rect 6489 1543 6497 1549
rect 6489 1514 6493 1543
rect 6521 1536 6527 1631
rect 6489 1507 6497 1514
rect 6493 1484 6497 1507
rect 6501 1484 6505 1524
rect 6521 1504 6525 1536
rect 6561 1522 6565 1648
rect 6577 1542 6581 1656
rect 6599 1644 6603 1656
rect 6601 1632 6603 1644
rect 6609 1644 6613 1656
rect 6609 1632 6611 1644
rect 6529 1510 6553 1512
rect 6529 1508 6565 1510
rect 6529 1504 6533 1508
rect 6575 1504 6579 1530
rect 6593 1522 6597 1632
rect 6631 1624 6635 1656
rect 6602 1620 6635 1624
rect 6602 1556 6606 1620
rect 6622 1571 6626 1600
rect 6641 1598 6645 1656
rect 6661 1599 6665 1636
rect 6622 1563 6631 1571
rect 6602 1544 6605 1556
rect 6595 1504 6599 1510
rect 6607 1504 6611 1544
rect 6627 1504 6631 1563
rect 6641 1504 6645 1586
rect 6661 1544 6665 1587
rect 4531 1460 4565 1464
rect 4581 1460 4585 1464
rect 4591 1460 4595 1464
rect 4651 1460 4685 1464
rect 4701 1460 4705 1464
rect 4711 1460 4715 1464
rect 4771 1460 4805 1464
rect 4821 1460 4825 1464
rect 4831 1460 4835 1464
rect 4891 1460 4925 1464
rect 4941 1460 4945 1464
rect 4951 1460 4955 1464
rect 5011 1460 5015 1464
rect 5033 1460 5037 1464
rect 5041 1460 5045 1464
rect 5061 1460 5065 1464
rect 5069 1460 5073 1464
rect 5115 1460 5119 1464
rect 5135 1460 5139 1464
rect 5147 1460 5151 1464
rect 5167 1460 5171 1464
rect 5181 1460 5185 1464
rect 5201 1460 5205 1464
rect 5251 1460 5255 1464
rect 5273 1460 5277 1464
rect 5281 1460 5285 1464
rect 5301 1460 5305 1464
rect 5309 1460 5313 1464
rect 5355 1460 5359 1464
rect 5375 1460 5379 1464
rect 5387 1460 5391 1464
rect 5407 1460 5411 1464
rect 5421 1460 5425 1464
rect 5441 1460 5445 1464
rect 5491 1460 5495 1464
rect 5511 1460 5515 1464
rect 5531 1460 5535 1464
rect 5551 1460 5555 1464
rect 5611 1460 5645 1464
rect 5661 1460 5665 1464
rect 5671 1460 5675 1464
rect 5750 1460 5754 1464
rect 5772 1460 5776 1464
rect 5780 1460 5784 1464
rect 5857 1460 5861 1464
rect 5865 1460 5869 1464
rect 5925 1460 5929 1464
rect 5945 1460 5949 1464
rect 6010 1460 6014 1464
rect 6032 1460 6036 1464
rect 6040 1460 6044 1464
rect 6117 1460 6121 1464
rect 6125 1460 6129 1464
rect 6195 1460 6199 1464
rect 6205 1460 6209 1464
rect 6235 1460 6239 1464
rect 6245 1460 6249 1464
rect 6305 1460 6309 1464
rect 6315 1460 6319 1464
rect 6335 1460 6369 1464
rect 6411 1460 6415 1464
rect 6471 1460 6475 1464
rect 6493 1460 6497 1464
rect 6501 1460 6505 1464
rect 6521 1460 6525 1464
rect 6529 1460 6533 1464
rect 6575 1460 6579 1464
rect 6595 1460 6599 1464
rect 6607 1460 6611 1464
rect 6627 1460 6631 1464
rect 6641 1460 6645 1464
rect 6661 1460 6665 1464
rect 31 1436 35 1440
rect 53 1436 57 1440
rect 75 1436 79 1440
rect 131 1436 135 1440
rect 139 1436 143 1440
rect 230 1436 234 1440
rect 252 1436 256 1440
rect 260 1436 264 1440
rect 337 1436 341 1440
rect 345 1436 349 1440
rect 391 1436 395 1440
rect 451 1436 455 1440
rect 525 1436 529 1440
rect 545 1436 549 1440
rect 591 1436 595 1440
rect 611 1436 615 1440
rect 631 1436 635 1440
rect 695 1436 699 1440
rect 715 1436 719 1440
rect 729 1436 733 1440
rect 749 1436 753 1440
rect 761 1436 765 1440
rect 781 1436 785 1440
rect 827 1436 831 1440
rect 835 1436 839 1440
rect 855 1436 859 1440
rect 863 1436 867 1440
rect 885 1436 889 1440
rect 945 1436 949 1440
rect 965 1436 969 1440
rect 1011 1436 1015 1440
rect 1031 1436 1035 1440
rect 1051 1436 1055 1440
rect 1111 1436 1115 1440
rect 1119 1436 1123 1440
rect 1195 1436 1199 1440
rect 1215 1436 1219 1440
rect 1229 1436 1233 1440
rect 1249 1436 1253 1440
rect 1261 1436 1265 1440
rect 1281 1436 1285 1440
rect 1327 1436 1331 1440
rect 1335 1436 1339 1440
rect 1355 1436 1359 1440
rect 1363 1436 1367 1440
rect 1385 1436 1389 1440
rect 1445 1436 1449 1440
rect 1465 1436 1469 1440
rect 1485 1436 1489 1440
rect 1505 1436 1509 1440
rect 1525 1436 1529 1440
rect 1545 1436 1549 1440
rect 1565 1436 1569 1440
rect 1585 1436 1589 1440
rect 1645 1436 1649 1440
rect 1655 1436 1659 1440
rect 1675 1436 1709 1440
rect 1777 1436 1781 1440
rect 1785 1436 1789 1440
rect 1855 1436 1859 1440
rect 1865 1436 1869 1440
rect 1895 1436 1899 1440
rect 1905 1436 1909 1440
rect 1970 1436 1974 1440
rect 1992 1436 1996 1440
rect 2000 1436 2004 1440
rect 2051 1436 2055 1440
rect 2116 1436 2120 1440
rect 2124 1436 2128 1440
rect 2146 1436 2150 1440
rect 2211 1436 2215 1440
rect 2231 1436 2235 1440
rect 2291 1436 2325 1440
rect 2341 1436 2345 1440
rect 2351 1436 2355 1440
rect 2425 1436 2429 1440
rect 2435 1436 2439 1440
rect 2455 1436 2489 1440
rect 2545 1436 2549 1440
rect 2565 1436 2569 1440
rect 2585 1436 2589 1440
rect 2605 1436 2609 1440
rect 2651 1436 2655 1440
rect 2671 1436 2675 1440
rect 2691 1436 2695 1440
rect 2711 1436 2715 1440
rect 2785 1436 2789 1440
rect 2805 1436 2809 1440
rect 2825 1436 2829 1440
rect 2845 1436 2849 1440
rect 2891 1436 2895 1440
rect 2913 1436 2917 1440
rect 2985 1436 2989 1440
rect 3005 1436 3009 1440
rect 3025 1436 3029 1440
rect 3045 1436 3049 1440
rect 3105 1436 3109 1440
rect 3165 1436 3169 1440
rect 3175 1436 3179 1440
rect 3195 1436 3229 1440
rect 3275 1436 3279 1440
rect 3295 1436 3299 1440
rect 3309 1436 3313 1440
rect 3329 1436 3333 1440
rect 3341 1436 3345 1440
rect 3361 1436 3365 1440
rect 3407 1436 3411 1440
rect 3415 1436 3419 1440
rect 3435 1436 3439 1440
rect 3443 1436 3447 1440
rect 3465 1436 3469 1440
rect 3537 1436 3541 1440
rect 3545 1436 3549 1440
rect 3615 1436 3619 1440
rect 3625 1436 3629 1440
rect 3655 1436 3659 1440
rect 3665 1436 3669 1440
rect 3730 1436 3734 1440
rect 3752 1436 3756 1440
rect 3760 1436 3764 1440
rect 3825 1436 3829 1440
rect 3871 1436 3875 1440
rect 3893 1436 3897 1440
rect 3901 1436 3905 1440
rect 3921 1436 3925 1440
rect 3929 1436 3933 1440
rect 3975 1436 3979 1440
rect 3995 1436 3999 1440
rect 4007 1436 4011 1440
rect 4027 1436 4031 1440
rect 4041 1436 4045 1440
rect 4061 1436 4065 1440
rect 4111 1436 4115 1440
rect 4133 1436 4137 1440
rect 4141 1436 4145 1440
rect 4161 1436 4165 1440
rect 4169 1436 4173 1440
rect 4215 1436 4219 1440
rect 4235 1436 4239 1440
rect 4247 1436 4251 1440
rect 4267 1436 4271 1440
rect 4281 1436 4285 1440
rect 4301 1436 4305 1440
rect 4365 1436 4369 1440
rect 4411 1436 4415 1440
rect 4431 1436 4435 1440
rect 4451 1436 4455 1440
rect 4471 1436 4475 1440
rect 4531 1436 4565 1440
rect 4581 1436 4585 1440
rect 4591 1436 4595 1440
rect 4665 1436 4669 1440
rect 4685 1436 4689 1440
rect 4705 1436 4709 1440
rect 4725 1436 4729 1440
rect 4783 1436 4787 1440
rect 4805 1436 4809 1440
rect 4865 1436 4869 1440
rect 4885 1436 4889 1440
rect 4945 1436 4949 1440
rect 4965 1436 4969 1440
rect 5035 1436 5039 1440
rect 5045 1436 5049 1440
rect 5075 1436 5079 1440
rect 5085 1436 5089 1440
rect 5155 1436 5159 1440
rect 5165 1436 5169 1440
rect 5195 1436 5199 1440
rect 5205 1436 5209 1440
rect 5251 1436 5255 1440
rect 5325 1436 5329 1440
rect 5345 1436 5349 1440
rect 5391 1436 5395 1440
rect 5401 1436 5405 1440
rect 5431 1436 5435 1440
rect 5441 1436 5445 1440
rect 5525 1436 5529 1440
rect 5545 1436 5549 1440
rect 5565 1436 5569 1440
rect 5611 1436 5615 1440
rect 5671 1436 5705 1440
rect 5721 1436 5725 1440
rect 5731 1436 5735 1440
rect 5805 1436 5809 1440
rect 5825 1436 5829 1440
rect 5890 1436 5894 1440
rect 5912 1436 5916 1440
rect 5920 1436 5924 1440
rect 5985 1436 5989 1440
rect 6036 1436 6040 1440
rect 6044 1436 6048 1440
rect 6066 1436 6070 1440
rect 6131 1436 6135 1440
rect 6141 1436 6145 1440
rect 6171 1436 6175 1440
rect 6181 1436 6185 1440
rect 6251 1436 6255 1440
rect 6273 1436 6277 1440
rect 6281 1436 6285 1440
rect 6301 1436 6305 1440
rect 6309 1436 6313 1440
rect 6355 1436 6359 1440
rect 6375 1436 6379 1440
rect 6387 1436 6391 1440
rect 6407 1436 6411 1440
rect 6421 1436 6425 1440
rect 6441 1436 6445 1440
rect 6491 1436 6495 1440
rect 6513 1436 6517 1440
rect 6521 1436 6525 1440
rect 6541 1436 6545 1440
rect 6549 1436 6553 1440
rect 6595 1436 6599 1440
rect 6615 1436 6619 1440
rect 6627 1436 6631 1440
rect 6647 1436 6651 1440
rect 6661 1436 6665 1440
rect 6681 1436 6685 1440
rect 31 1333 35 1396
rect 26 1321 35 1333
rect 31 1264 35 1321
rect 53 1319 57 1396
rect 41 1307 54 1319
rect 41 1264 45 1307
rect 75 1282 79 1356
rect 131 1333 135 1356
rect 126 1321 135 1333
rect 139 1333 143 1356
rect 230 1353 234 1396
rect 227 1341 234 1353
rect 139 1321 154 1333
rect 67 1270 79 1282
rect 61 1264 65 1270
rect 131 1244 135 1321
rect 151 1244 155 1321
rect 225 1264 229 1341
rect 252 1299 256 1356
rect 260 1352 264 1356
rect 260 1344 278 1352
rect 274 1333 278 1344
rect 337 1333 341 1356
rect 326 1321 341 1333
rect 345 1333 349 1356
rect 345 1321 354 1333
rect 245 1287 254 1299
rect 245 1264 249 1287
rect 274 1276 278 1321
rect 265 1269 278 1276
rect 265 1264 269 1269
rect 325 1244 329 1321
rect 345 1244 349 1321
rect 391 1313 395 1396
rect 451 1313 455 1396
rect 525 1319 529 1396
rect 386 1301 395 1313
rect 446 1301 455 1313
rect 526 1307 529 1319
rect 391 1244 395 1301
rect 451 1244 455 1301
rect 523 1291 529 1307
rect 545 1319 549 1396
rect 591 1342 595 1356
rect 611 1342 615 1356
rect 579 1336 595 1342
rect 600 1336 615 1342
rect 545 1307 554 1319
rect 545 1291 551 1307
rect 579 1299 586 1336
rect 600 1313 606 1336
rect 523 1284 537 1291
rect 533 1264 537 1284
rect 543 1284 551 1291
rect 543 1264 547 1284
rect 579 1274 586 1287
rect 579 1268 598 1274
rect 594 1264 598 1268
rect 602 1264 606 1301
rect 631 1299 635 1356
rect 695 1313 699 1356
rect 715 1314 719 1396
rect 729 1337 733 1396
rect 749 1356 753 1396
rect 761 1390 765 1396
rect 755 1344 758 1356
rect 729 1329 738 1337
rect 626 1287 635 1299
rect 624 1244 628 1287
rect 695 1264 699 1301
rect 715 1244 719 1302
rect 734 1300 738 1329
rect 754 1280 758 1344
rect 725 1276 758 1280
rect 725 1244 729 1276
rect 763 1268 767 1378
rect 781 1370 785 1396
rect 827 1392 831 1396
rect 795 1390 831 1392
rect 807 1388 831 1390
rect 749 1256 751 1268
rect 747 1244 751 1256
rect 757 1256 759 1268
rect 757 1244 761 1256
rect 779 1244 783 1358
rect 795 1252 799 1378
rect 835 1364 839 1396
rect 855 1376 859 1416
rect 863 1393 867 1416
rect 863 1386 871 1393
rect 833 1269 839 1364
rect 867 1357 871 1386
rect 863 1351 871 1357
rect 863 1305 867 1351
rect 885 1344 889 1356
rect 887 1332 889 1344
rect 833 1265 857 1269
rect 819 1260 837 1261
rect 807 1256 837 1260
rect 795 1248 829 1252
rect 825 1244 829 1248
rect 833 1244 837 1256
rect 853 1244 857 1265
rect 863 1244 867 1293
rect 885 1264 889 1332
rect 945 1319 949 1396
rect 946 1307 949 1319
rect 943 1291 949 1307
rect 965 1319 969 1396
rect 1011 1388 1015 1396
rect 1000 1384 1015 1388
rect 1031 1384 1035 1396
rect 1000 1353 1006 1384
rect 1020 1380 1035 1384
rect 1020 1373 1026 1380
rect 1006 1341 1016 1353
rect 965 1307 974 1319
rect 965 1291 971 1307
rect 943 1284 957 1291
rect 953 1264 957 1284
rect 963 1284 971 1291
rect 1012 1284 1016 1341
rect 1020 1284 1024 1361
rect 1051 1353 1055 1396
rect 1028 1341 1035 1353
rect 1047 1341 1055 1353
rect 1028 1284 1032 1341
rect 1111 1333 1115 1356
rect 1106 1321 1115 1333
rect 1119 1333 1123 1356
rect 1119 1321 1134 1333
rect 963 1264 967 1284
rect 1111 1244 1115 1321
rect 1131 1244 1135 1321
rect 1195 1313 1199 1356
rect 1215 1314 1219 1396
rect 1229 1337 1233 1396
rect 1249 1356 1253 1396
rect 1261 1390 1265 1396
rect 1255 1344 1258 1356
rect 1229 1329 1238 1337
rect 1195 1264 1199 1301
rect 1215 1244 1219 1302
rect 1234 1300 1238 1329
rect 1254 1280 1258 1344
rect 1225 1276 1258 1280
rect 1225 1244 1229 1276
rect 1263 1268 1267 1378
rect 1281 1370 1285 1396
rect 1327 1392 1331 1396
rect 1295 1390 1331 1392
rect 1307 1388 1331 1390
rect 1249 1256 1251 1268
rect 1247 1244 1251 1256
rect 1257 1256 1259 1268
rect 1257 1244 1261 1256
rect 1279 1244 1283 1358
rect 1295 1252 1299 1378
rect 1335 1364 1339 1396
rect 1355 1376 1359 1416
rect 1363 1393 1367 1416
rect 1363 1386 1371 1393
rect 1333 1269 1339 1364
rect 1367 1357 1371 1386
rect 1363 1351 1371 1357
rect 1675 1428 1679 1436
rect 1685 1428 1689 1432
rect 1705 1428 1709 1436
rect 1363 1305 1367 1351
rect 1385 1344 1389 1356
rect 1387 1332 1389 1344
rect 1333 1265 1357 1269
rect 1319 1260 1337 1261
rect 1307 1256 1337 1260
rect 1295 1248 1329 1252
rect 1325 1244 1329 1248
rect 1333 1244 1337 1256
rect 1353 1244 1357 1265
rect 1363 1244 1367 1293
rect 1385 1264 1389 1332
rect 1445 1296 1449 1356
rect 1465 1296 1469 1356
rect 1485 1296 1489 1356
rect 1505 1296 1509 1356
rect 1525 1296 1529 1356
rect 1545 1296 1549 1356
rect 1565 1299 1569 1356
rect 1585 1299 1589 1356
rect 1645 1333 1649 1356
rect 1646 1321 1649 1333
rect 1655 1334 1659 1356
rect 1705 1384 1709 1388
rect 1705 1380 1717 1384
rect 1675 1344 1679 1348
rect 1685 1343 1689 1348
rect 1685 1339 1698 1343
rect 1655 1330 1685 1334
rect 1445 1284 1458 1296
rect 1485 1284 1498 1296
rect 1525 1284 1538 1296
rect 1565 1287 1574 1299
rect 1586 1287 1589 1299
rect 1445 1264 1449 1284
rect 1465 1264 1469 1284
rect 1485 1264 1489 1284
rect 1505 1264 1509 1284
rect 1525 1264 1529 1284
rect 1545 1264 1549 1284
rect 1565 1264 1569 1287
rect 1585 1264 1589 1287
rect 1645 1272 1649 1321
rect 1693 1333 1698 1339
rect 1655 1272 1659 1276
rect 1675 1272 1679 1318
rect 1694 1290 1699 1321
rect 1685 1284 1699 1290
rect 1713 1299 1717 1380
rect 1777 1333 1781 1356
rect 1766 1321 1781 1333
rect 1785 1333 1789 1356
rect 1855 1352 1859 1356
rect 1845 1348 1859 1352
rect 1845 1333 1849 1348
rect 1785 1321 1794 1333
rect 1847 1321 1849 1333
rect 1685 1272 1689 1284
rect 1713 1261 1717 1287
rect 1705 1256 1717 1261
rect 1705 1252 1709 1256
rect 1765 1244 1769 1321
rect 1785 1244 1789 1321
rect 1845 1264 1849 1321
rect 1865 1299 1869 1356
rect 1895 1352 1899 1356
rect 1885 1348 1899 1352
rect 1905 1352 1909 1356
rect 1970 1353 1974 1396
rect 1905 1348 1919 1352
rect 1885 1299 1891 1348
rect 1914 1333 1919 1348
rect 1967 1341 1974 1353
rect 1885 1287 1894 1299
rect 1865 1264 1869 1287
rect 1885 1264 1889 1287
rect 1914 1275 1920 1321
rect 1905 1271 1920 1275
rect 1905 1264 1909 1271
rect 1965 1264 1969 1341
rect 1992 1299 1996 1356
rect 2000 1352 2004 1356
rect 2000 1344 2018 1352
rect 2014 1333 2018 1344
rect 1985 1287 1994 1299
rect 1985 1264 1989 1287
rect 2014 1276 2018 1321
rect 2051 1313 2055 1396
rect 2291 1428 2295 1436
rect 2311 1428 2315 1432
rect 2321 1428 2325 1436
rect 2116 1352 2120 1356
rect 2102 1344 2120 1352
rect 2102 1333 2106 1344
rect 2046 1301 2055 1313
rect 2005 1269 2018 1276
rect 2005 1264 2009 1269
rect 1645 1228 1649 1232
rect 1655 1224 1659 1232
rect 1675 1228 1679 1232
rect 1685 1228 1689 1232
rect 1705 1224 1709 1232
rect 2051 1244 2055 1301
rect 2102 1276 2106 1321
rect 2124 1299 2128 1356
rect 2146 1353 2150 1396
rect 2146 1341 2153 1353
rect 2126 1287 2135 1299
rect 2102 1269 2115 1276
rect 2111 1264 2115 1269
rect 2131 1264 2135 1287
rect 2151 1264 2155 1341
rect 2211 1319 2215 1396
rect 2206 1307 2215 1319
rect 2209 1291 2215 1307
rect 2231 1319 2235 1396
rect 2291 1384 2295 1388
rect 2283 1380 2295 1384
rect 2231 1307 2234 1319
rect 2231 1291 2237 1307
rect 2283 1299 2287 1380
rect 2455 1428 2459 1436
rect 2465 1428 2469 1432
rect 2485 1428 2489 1436
rect 2311 1343 2315 1348
rect 2321 1344 2325 1348
rect 2302 1339 2315 1343
rect 2302 1333 2307 1339
rect 2341 1334 2345 1356
rect 2315 1330 2345 1334
rect 2351 1333 2355 1356
rect 2425 1333 2429 1356
rect 2209 1284 2217 1291
rect 2213 1264 2217 1284
rect 2223 1284 2237 1291
rect 2223 1264 2227 1284
rect 2283 1261 2287 1287
rect 2301 1290 2306 1321
rect 2351 1321 2354 1333
rect 2426 1321 2429 1333
rect 2435 1334 2439 1356
rect 2485 1384 2489 1388
rect 2485 1380 2497 1384
rect 2455 1344 2459 1348
rect 2465 1343 2469 1348
rect 2465 1339 2478 1343
rect 2435 1330 2465 1334
rect 2301 1284 2315 1290
rect 2311 1272 2315 1284
rect 2321 1272 2325 1318
rect 2341 1272 2345 1276
rect 2351 1272 2355 1321
rect 2425 1272 2429 1321
rect 2473 1333 2478 1339
rect 2435 1272 2439 1276
rect 2455 1272 2459 1318
rect 2474 1290 2479 1321
rect 2465 1284 2479 1290
rect 2493 1299 2497 1380
rect 2545 1333 2549 1356
rect 2546 1321 2549 1333
rect 2465 1272 2469 1284
rect 2283 1256 2295 1261
rect 2291 1252 2295 1256
rect 2493 1261 2497 1287
rect 2540 1273 2546 1321
rect 2565 1299 2569 1356
rect 2585 1334 2589 1356
rect 2605 1334 2609 1356
rect 2651 1334 2655 1356
rect 2671 1334 2675 1356
rect 2585 1328 2598 1334
rect 2605 1333 2625 1334
rect 2605 1328 2613 1333
rect 2594 1299 2598 1328
rect 2635 1333 2655 1334
rect 2647 1328 2655 1333
rect 2662 1328 2675 1334
rect 2567 1287 2569 1299
rect 2565 1285 2569 1287
rect 2565 1278 2578 1285
rect 2540 1269 2570 1273
rect 2566 1264 2570 1269
rect 2574 1264 2578 1278
rect 2594 1264 2598 1287
rect 2613 1279 2619 1321
rect 2602 1272 2619 1279
rect 2641 1279 2647 1321
rect 2662 1299 2666 1328
rect 2691 1299 2695 1356
rect 2711 1333 2715 1356
rect 2785 1333 2789 1356
rect 2711 1321 2714 1333
rect 2786 1321 2789 1333
rect 2691 1287 2693 1299
rect 2641 1272 2658 1279
rect 2602 1264 2606 1272
rect 2654 1264 2658 1272
rect 2662 1264 2666 1287
rect 2691 1285 2695 1287
rect 2682 1278 2695 1285
rect 2682 1264 2686 1278
rect 2714 1273 2720 1321
rect 2690 1269 2720 1273
rect 2780 1273 2786 1321
rect 2805 1299 2809 1356
rect 2825 1334 2829 1356
rect 2845 1334 2849 1356
rect 2825 1328 2838 1334
rect 2845 1333 2865 1334
rect 2891 1333 2895 1396
rect 2913 1350 2917 1356
rect 2915 1338 2917 1350
rect 2985 1333 2989 1356
rect 2845 1328 2853 1333
rect 2834 1299 2838 1328
rect 2886 1321 2895 1333
rect 2986 1321 2989 1333
rect 2807 1287 2809 1299
rect 2805 1285 2809 1287
rect 2805 1278 2818 1285
rect 2780 1269 2810 1273
rect 2690 1264 2694 1269
rect 2806 1264 2810 1269
rect 2814 1264 2818 1278
rect 2834 1264 2838 1287
rect 2853 1279 2859 1321
rect 2842 1272 2859 1279
rect 2842 1264 2846 1272
rect 2485 1256 2497 1261
rect 2485 1252 2489 1256
rect 2291 1224 2295 1232
rect 2311 1228 2315 1232
rect 2321 1228 2325 1232
rect 2341 1224 2345 1232
rect 2351 1228 2355 1232
rect 2425 1228 2429 1232
rect 31 1220 35 1224
rect 41 1220 45 1224
rect 61 1220 65 1224
rect 131 1220 135 1224
rect 151 1220 155 1224
rect 225 1220 229 1224
rect 245 1220 249 1224
rect 265 1220 269 1224
rect 325 1220 329 1224
rect 345 1220 349 1224
rect 391 1220 395 1224
rect 451 1220 455 1224
rect 533 1220 537 1224
rect 543 1220 547 1224
rect 594 1220 598 1224
rect 602 1220 606 1224
rect 624 1220 628 1224
rect 695 1220 699 1224
rect 715 1220 719 1224
rect 725 1220 729 1224
rect 747 1220 751 1224
rect 757 1220 761 1224
rect 779 1220 783 1224
rect 825 1220 829 1224
rect 833 1220 837 1224
rect 853 1220 857 1224
rect 863 1220 867 1224
rect 885 1220 889 1224
rect 953 1220 957 1224
rect 963 1220 967 1224
rect 1012 1220 1016 1224
rect 1020 1220 1024 1224
rect 1028 1220 1032 1224
rect 1111 1220 1115 1224
rect 1131 1220 1135 1224
rect 1195 1220 1199 1224
rect 1215 1220 1219 1224
rect 1225 1220 1229 1224
rect 1247 1220 1251 1224
rect 1257 1220 1261 1224
rect 1279 1220 1283 1224
rect 1325 1220 1329 1224
rect 1333 1220 1337 1224
rect 1353 1220 1357 1224
rect 1363 1220 1367 1224
rect 1385 1220 1389 1224
rect 1445 1220 1449 1224
rect 1465 1220 1469 1224
rect 1485 1220 1489 1224
rect 1505 1220 1509 1224
rect 1525 1220 1529 1224
rect 1545 1220 1549 1224
rect 1565 1220 1569 1224
rect 1585 1220 1589 1224
rect 1655 1220 1709 1224
rect 1765 1220 1769 1224
rect 1785 1220 1789 1224
rect 1845 1220 1849 1224
rect 1865 1220 1869 1224
rect 1885 1220 1889 1224
rect 1905 1220 1909 1224
rect 1965 1220 1969 1224
rect 1985 1220 1989 1224
rect 2005 1220 2009 1224
rect 2051 1220 2055 1224
rect 2111 1220 2115 1224
rect 2131 1220 2135 1224
rect 2151 1220 2155 1224
rect 2213 1220 2217 1224
rect 2223 1220 2227 1224
rect 2291 1220 2345 1224
rect 2435 1224 2439 1232
rect 2455 1228 2459 1232
rect 2465 1228 2469 1232
rect 2485 1224 2489 1232
rect 2891 1244 2895 1321
rect 2915 1270 2917 1282
rect 2913 1264 2917 1270
rect 2980 1273 2986 1321
rect 3005 1299 3009 1356
rect 3025 1334 3029 1356
rect 3045 1334 3049 1356
rect 3025 1328 3038 1334
rect 3045 1333 3065 1334
rect 3045 1328 3053 1333
rect 3034 1299 3038 1328
rect 3007 1287 3009 1299
rect 3005 1285 3009 1287
rect 3005 1278 3018 1285
rect 2980 1269 3010 1273
rect 3006 1264 3010 1269
rect 3014 1264 3018 1278
rect 3034 1264 3038 1287
rect 3053 1279 3059 1321
rect 3042 1272 3059 1279
rect 3105 1313 3109 1396
rect 3195 1428 3199 1436
rect 3205 1428 3209 1432
rect 3225 1428 3229 1436
rect 3165 1333 3169 1356
rect 3166 1321 3169 1333
rect 3175 1334 3179 1356
rect 3225 1384 3229 1388
rect 3225 1380 3237 1384
rect 3195 1344 3199 1348
rect 3205 1343 3209 1348
rect 3205 1339 3218 1343
rect 3175 1330 3205 1334
rect 3105 1301 3114 1313
rect 3042 1264 3046 1272
rect 3105 1244 3109 1301
rect 3165 1272 3169 1321
rect 3213 1333 3218 1339
rect 3175 1272 3179 1276
rect 3195 1272 3199 1318
rect 3214 1290 3219 1321
rect 3205 1284 3219 1290
rect 3233 1299 3237 1380
rect 3275 1313 3279 1356
rect 3295 1314 3299 1396
rect 3309 1337 3313 1396
rect 3329 1356 3333 1396
rect 3341 1390 3345 1396
rect 3335 1344 3338 1356
rect 3309 1329 3318 1337
rect 3205 1272 3209 1284
rect 3233 1261 3237 1287
rect 3275 1264 3279 1301
rect 3225 1256 3237 1261
rect 3225 1252 3229 1256
rect 3165 1228 3169 1232
rect 3175 1224 3179 1232
rect 3195 1228 3199 1232
rect 3205 1228 3209 1232
rect 3225 1224 3229 1232
rect 3295 1244 3299 1302
rect 3314 1300 3318 1329
rect 3334 1280 3338 1344
rect 3305 1276 3338 1280
rect 3305 1244 3309 1276
rect 3343 1268 3347 1378
rect 3361 1370 3365 1396
rect 3407 1392 3411 1396
rect 3375 1390 3411 1392
rect 3387 1388 3411 1390
rect 3329 1256 3331 1268
rect 3327 1244 3331 1256
rect 3337 1256 3339 1268
rect 3337 1244 3341 1256
rect 3359 1244 3363 1358
rect 3375 1252 3379 1378
rect 3415 1364 3419 1396
rect 3435 1376 3439 1416
rect 3443 1393 3447 1416
rect 3443 1386 3451 1393
rect 3413 1269 3419 1364
rect 3447 1357 3451 1386
rect 3443 1351 3451 1357
rect 3443 1305 3447 1351
rect 3465 1344 3469 1356
rect 3467 1332 3469 1344
rect 3537 1333 3541 1356
rect 3413 1265 3437 1269
rect 3399 1260 3417 1261
rect 3387 1256 3417 1260
rect 3375 1248 3409 1252
rect 3405 1244 3409 1248
rect 3413 1244 3417 1256
rect 3433 1244 3437 1265
rect 3443 1244 3447 1293
rect 3465 1264 3469 1332
rect 3526 1321 3541 1333
rect 3545 1333 3549 1356
rect 3615 1352 3619 1356
rect 3605 1348 3619 1352
rect 3605 1333 3609 1348
rect 3545 1321 3554 1333
rect 3607 1321 3609 1333
rect 3525 1244 3529 1321
rect 3545 1244 3549 1321
rect 3605 1264 3609 1321
rect 3625 1299 3629 1356
rect 3655 1352 3659 1356
rect 3645 1348 3659 1352
rect 3665 1352 3669 1356
rect 3730 1353 3734 1396
rect 3665 1348 3679 1352
rect 3645 1299 3651 1348
rect 3674 1333 3679 1348
rect 3727 1341 3734 1353
rect 3645 1287 3654 1299
rect 3625 1264 3629 1287
rect 3645 1264 3649 1287
rect 3674 1275 3680 1321
rect 3665 1271 3680 1275
rect 3665 1264 3669 1271
rect 3725 1264 3729 1341
rect 3752 1299 3756 1356
rect 3760 1352 3764 1356
rect 3760 1344 3778 1352
rect 3774 1333 3778 1344
rect 3745 1287 3754 1299
rect 3745 1264 3749 1287
rect 3774 1276 3778 1321
rect 3765 1269 3778 1276
rect 3825 1313 3829 1396
rect 3893 1393 3897 1416
rect 3889 1386 3897 1393
rect 3889 1357 3893 1386
rect 3901 1376 3905 1416
rect 3921 1364 3925 1396
rect 3929 1392 3933 1396
rect 3929 1390 3965 1392
rect 3929 1388 3953 1390
rect 3871 1344 3875 1356
rect 3889 1351 3897 1357
rect 3871 1332 3873 1344
rect 3825 1301 3834 1313
rect 3765 1264 3769 1269
rect 3825 1244 3829 1301
rect 3871 1264 3875 1332
rect 3893 1305 3897 1351
rect 3893 1244 3897 1293
rect 3921 1269 3927 1364
rect 3903 1265 3927 1269
rect 3903 1244 3907 1265
rect 3923 1260 3941 1261
rect 3923 1256 3953 1260
rect 3923 1244 3927 1256
rect 3961 1252 3965 1378
rect 3975 1370 3979 1396
rect 3995 1390 3999 1396
rect 3931 1248 3965 1252
rect 3931 1244 3935 1248
rect 3977 1244 3981 1358
rect 3993 1268 3997 1378
rect 4007 1356 4011 1396
rect 4002 1344 4005 1356
rect 4002 1280 4006 1344
rect 4027 1337 4031 1396
rect 4022 1329 4031 1337
rect 4022 1300 4026 1329
rect 4041 1314 4045 1396
rect 4133 1393 4137 1416
rect 4129 1386 4137 1393
rect 4129 1357 4133 1386
rect 4141 1376 4145 1416
rect 4161 1364 4165 1396
rect 4169 1392 4173 1396
rect 4169 1390 4205 1392
rect 4169 1388 4193 1390
rect 4061 1313 4065 1356
rect 4111 1344 4115 1356
rect 4129 1351 4137 1357
rect 4111 1332 4113 1344
rect 4002 1276 4035 1280
rect 4001 1256 4003 1268
rect 3999 1244 4003 1256
rect 4009 1256 4011 1268
rect 4009 1244 4013 1256
rect 4031 1244 4035 1276
rect 4041 1244 4045 1302
rect 4061 1264 4065 1301
rect 4111 1264 4115 1332
rect 4133 1305 4137 1351
rect 4133 1244 4137 1293
rect 4161 1269 4167 1364
rect 4143 1265 4167 1269
rect 4143 1244 4147 1265
rect 4163 1260 4181 1261
rect 4163 1256 4193 1260
rect 4163 1244 4167 1256
rect 4201 1252 4205 1378
rect 4215 1370 4219 1396
rect 4235 1390 4239 1396
rect 4171 1248 4205 1252
rect 4171 1244 4175 1248
rect 4217 1244 4221 1358
rect 4233 1268 4237 1378
rect 4247 1356 4251 1396
rect 4242 1344 4245 1356
rect 4242 1280 4246 1344
rect 4267 1337 4271 1396
rect 4262 1329 4271 1337
rect 4262 1300 4266 1329
rect 4281 1314 4285 1396
rect 4301 1313 4305 1356
rect 4365 1313 4369 1396
rect 4531 1428 4535 1436
rect 4551 1428 4555 1432
rect 4561 1428 4565 1436
rect 4531 1384 4535 1388
rect 4523 1380 4535 1384
rect 4411 1334 4415 1356
rect 4431 1334 4435 1356
rect 4395 1333 4415 1334
rect 4407 1328 4415 1333
rect 4422 1328 4435 1334
rect 4242 1276 4275 1280
rect 4241 1256 4243 1268
rect 4239 1244 4243 1256
rect 4249 1256 4251 1268
rect 4249 1244 4253 1256
rect 4271 1244 4275 1276
rect 4281 1244 4285 1302
rect 4365 1301 4374 1313
rect 4301 1264 4305 1301
rect 4365 1244 4369 1301
rect 4401 1279 4407 1321
rect 4422 1299 4426 1328
rect 4451 1299 4455 1356
rect 4471 1333 4475 1356
rect 4471 1321 4474 1333
rect 4451 1287 4453 1299
rect 4401 1272 4418 1279
rect 4414 1264 4418 1272
rect 4422 1264 4426 1287
rect 4451 1285 4455 1287
rect 4442 1278 4455 1285
rect 4442 1264 4446 1278
rect 4474 1273 4480 1321
rect 4523 1299 4527 1380
rect 4551 1343 4555 1348
rect 4561 1344 4565 1348
rect 4542 1339 4555 1343
rect 4542 1333 4547 1339
rect 4581 1334 4585 1356
rect 4555 1330 4585 1334
rect 4591 1333 4595 1356
rect 4665 1333 4669 1356
rect 4450 1269 4480 1273
rect 4450 1264 4454 1269
rect 4523 1261 4527 1287
rect 4541 1290 4546 1321
rect 4591 1321 4594 1333
rect 4666 1321 4669 1333
rect 4541 1284 4555 1290
rect 4551 1272 4555 1284
rect 4561 1272 4565 1318
rect 4581 1272 4585 1276
rect 4591 1272 4595 1321
rect 4660 1273 4666 1321
rect 4685 1299 4689 1356
rect 4705 1334 4709 1356
rect 4725 1334 4729 1356
rect 4783 1350 4787 1356
rect 4783 1338 4785 1350
rect 4705 1328 4718 1334
rect 4725 1333 4745 1334
rect 4725 1328 4733 1333
rect 4714 1299 4718 1328
rect 4805 1333 4809 1396
rect 4805 1321 4814 1333
rect 4687 1287 4689 1299
rect 4685 1285 4689 1287
rect 4685 1278 4698 1285
rect 4523 1256 4535 1261
rect 4531 1252 4535 1256
rect 4660 1269 4690 1273
rect 4686 1264 4690 1269
rect 4694 1264 4698 1278
rect 4714 1264 4718 1287
rect 4733 1279 4739 1321
rect 4722 1272 4739 1279
rect 4722 1264 4726 1272
rect 4783 1270 4785 1282
rect 4783 1264 4787 1270
rect 4531 1224 4535 1232
rect 4551 1228 4555 1232
rect 4561 1228 4565 1232
rect 4581 1224 4585 1232
rect 4591 1228 4595 1232
rect 4805 1244 4809 1321
rect 4865 1319 4869 1396
rect 4866 1307 4869 1319
rect 4863 1291 4869 1307
rect 4885 1319 4889 1396
rect 4945 1319 4949 1396
rect 4885 1307 4894 1319
rect 4946 1307 4949 1319
rect 4885 1291 4891 1307
rect 4863 1284 4877 1291
rect 4873 1264 4877 1284
rect 4883 1284 4891 1291
rect 4943 1291 4949 1307
rect 4965 1319 4969 1396
rect 5035 1352 5039 1356
rect 5025 1348 5039 1352
rect 5025 1333 5029 1348
rect 5027 1321 5029 1333
rect 4965 1307 4974 1319
rect 4965 1291 4971 1307
rect 4943 1284 4957 1291
rect 4883 1264 4887 1284
rect 4953 1264 4957 1284
rect 4963 1284 4971 1291
rect 4963 1264 4967 1284
rect 5025 1264 5029 1321
rect 5045 1299 5049 1356
rect 5075 1352 5079 1356
rect 5065 1348 5079 1352
rect 5085 1352 5089 1356
rect 5155 1352 5159 1356
rect 5085 1348 5099 1352
rect 5065 1299 5071 1348
rect 5094 1333 5099 1348
rect 5145 1348 5159 1352
rect 5145 1333 5149 1348
rect 5147 1321 5149 1333
rect 5065 1287 5074 1299
rect 5045 1264 5049 1287
rect 5065 1264 5069 1287
rect 5094 1275 5100 1321
rect 5085 1271 5100 1275
rect 5085 1264 5089 1271
rect 5145 1264 5149 1321
rect 5165 1299 5169 1356
rect 5195 1352 5199 1356
rect 5185 1348 5199 1352
rect 5205 1352 5209 1356
rect 5205 1348 5219 1352
rect 5185 1299 5191 1348
rect 5214 1333 5219 1348
rect 5185 1287 5194 1299
rect 5165 1264 5169 1287
rect 5185 1264 5189 1287
rect 5214 1275 5220 1321
rect 5251 1299 5255 1356
rect 5325 1319 5329 1396
rect 5326 1307 5329 1319
rect 5246 1287 5255 1299
rect 5205 1271 5220 1275
rect 5205 1264 5209 1271
rect 5251 1264 5255 1287
rect 5323 1291 5329 1307
rect 5345 1319 5349 1396
rect 5671 1428 5675 1436
rect 5691 1428 5695 1432
rect 5701 1428 5705 1436
rect 5671 1384 5675 1388
rect 5663 1380 5675 1384
rect 5391 1352 5395 1356
rect 5381 1348 5395 1352
rect 5401 1352 5405 1356
rect 5401 1348 5415 1352
rect 5381 1333 5386 1348
rect 5345 1307 5354 1319
rect 5345 1291 5351 1307
rect 5323 1284 5337 1291
rect 5333 1264 5337 1284
rect 5343 1284 5351 1291
rect 5343 1264 5347 1284
rect 5380 1275 5386 1321
rect 5409 1299 5415 1348
rect 5431 1299 5435 1356
rect 5441 1352 5445 1356
rect 5441 1348 5455 1352
rect 5451 1333 5455 1348
rect 5451 1321 5453 1333
rect 5406 1287 5415 1299
rect 5380 1271 5395 1275
rect 5391 1264 5395 1271
rect 5411 1264 5415 1287
rect 5431 1264 5435 1287
rect 5451 1264 5455 1321
rect 5525 1299 5529 1356
rect 5545 1342 5549 1356
rect 5565 1342 5569 1356
rect 5545 1336 5560 1342
rect 5565 1336 5581 1342
rect 5554 1313 5560 1336
rect 5525 1287 5534 1299
rect 5532 1244 5536 1287
rect 5554 1264 5558 1301
rect 5574 1299 5581 1336
rect 5611 1299 5615 1356
rect 5663 1299 5667 1380
rect 5691 1343 5695 1348
rect 5701 1344 5705 1348
rect 5682 1339 5695 1343
rect 5682 1333 5687 1339
rect 5721 1334 5725 1356
rect 5695 1330 5725 1334
rect 5731 1333 5735 1356
rect 5606 1287 5615 1299
rect 5574 1274 5581 1287
rect 5562 1268 5581 1274
rect 5562 1264 5566 1268
rect 5611 1264 5615 1287
rect 5663 1261 5667 1287
rect 5681 1290 5686 1321
rect 5731 1321 5734 1333
rect 5681 1284 5695 1290
rect 5691 1272 5695 1284
rect 5701 1272 5705 1318
rect 5721 1272 5725 1276
rect 5731 1272 5735 1321
rect 5805 1319 5809 1396
rect 5806 1307 5809 1319
rect 5803 1291 5809 1307
rect 5825 1319 5829 1396
rect 5890 1353 5894 1396
rect 5887 1341 5894 1353
rect 5825 1307 5834 1319
rect 5825 1291 5831 1307
rect 5803 1284 5817 1291
rect 5663 1256 5675 1261
rect 5671 1252 5675 1256
rect 5813 1264 5817 1284
rect 5823 1284 5831 1291
rect 5823 1264 5827 1284
rect 5885 1264 5889 1341
rect 5912 1299 5916 1356
rect 5920 1352 5924 1356
rect 5920 1344 5938 1352
rect 5934 1333 5938 1344
rect 5905 1287 5914 1299
rect 5905 1264 5909 1287
rect 5934 1276 5938 1321
rect 5925 1269 5938 1276
rect 5985 1313 5989 1396
rect 6036 1352 6040 1356
rect 6022 1344 6040 1352
rect 6022 1333 6026 1344
rect 5985 1301 5994 1313
rect 5925 1264 5929 1269
rect 5671 1224 5675 1232
rect 5691 1228 5695 1232
rect 5701 1228 5705 1232
rect 5721 1224 5725 1232
rect 5731 1228 5735 1232
rect 5985 1244 5989 1301
rect 6022 1276 6026 1321
rect 6044 1299 6048 1356
rect 6066 1353 6070 1396
rect 6273 1393 6277 1416
rect 6269 1386 6277 1393
rect 6269 1357 6273 1386
rect 6281 1376 6285 1416
rect 6301 1364 6305 1396
rect 6309 1392 6313 1396
rect 6309 1390 6345 1392
rect 6309 1388 6333 1390
rect 6066 1341 6073 1353
rect 6131 1352 6135 1356
rect 6121 1348 6135 1352
rect 6141 1352 6145 1356
rect 6141 1348 6155 1352
rect 6046 1287 6055 1299
rect 6022 1269 6035 1276
rect 6031 1264 6035 1269
rect 6051 1264 6055 1287
rect 6071 1264 6075 1341
rect 6121 1333 6126 1348
rect 6120 1275 6126 1321
rect 6149 1299 6155 1348
rect 6171 1299 6175 1356
rect 6181 1352 6185 1356
rect 6181 1348 6195 1352
rect 6191 1333 6195 1348
rect 6251 1344 6255 1356
rect 6269 1351 6277 1357
rect 6191 1321 6193 1333
rect 6251 1332 6253 1344
rect 6146 1287 6155 1299
rect 6120 1271 6135 1275
rect 6131 1264 6135 1271
rect 6151 1264 6155 1287
rect 6171 1264 6175 1287
rect 6191 1264 6195 1321
rect 6251 1264 6255 1332
rect 6273 1305 6277 1351
rect 6273 1244 6277 1293
rect 6301 1269 6307 1364
rect 6283 1265 6307 1269
rect 6283 1244 6287 1265
rect 6303 1260 6321 1261
rect 6303 1256 6333 1260
rect 6303 1244 6307 1256
rect 6341 1252 6345 1378
rect 6355 1370 6359 1396
rect 6375 1390 6379 1396
rect 6311 1248 6345 1252
rect 6311 1244 6315 1248
rect 6357 1244 6361 1358
rect 6373 1268 6377 1378
rect 6387 1356 6391 1396
rect 6382 1344 6385 1356
rect 6382 1280 6386 1344
rect 6407 1337 6411 1396
rect 6402 1329 6411 1337
rect 6402 1300 6406 1329
rect 6421 1314 6425 1396
rect 6513 1393 6517 1416
rect 6509 1386 6517 1393
rect 6509 1357 6513 1386
rect 6521 1376 6525 1416
rect 6541 1364 6545 1396
rect 6549 1392 6553 1396
rect 6549 1390 6585 1392
rect 6549 1388 6573 1390
rect 6441 1313 6445 1356
rect 6491 1344 6495 1356
rect 6509 1351 6517 1357
rect 6491 1332 6493 1344
rect 6382 1276 6415 1280
rect 6381 1256 6383 1268
rect 6379 1244 6383 1256
rect 6389 1256 6391 1268
rect 6389 1244 6393 1256
rect 6411 1244 6415 1276
rect 6421 1244 6425 1302
rect 6441 1264 6445 1301
rect 6491 1264 6495 1332
rect 6513 1305 6517 1351
rect 6513 1244 6517 1293
rect 6541 1269 6547 1364
rect 6523 1265 6547 1269
rect 6523 1244 6527 1265
rect 6543 1260 6561 1261
rect 6543 1256 6573 1260
rect 6543 1244 6547 1256
rect 6581 1252 6585 1378
rect 6595 1370 6599 1396
rect 6615 1390 6619 1396
rect 6551 1248 6585 1252
rect 6551 1244 6555 1248
rect 6597 1244 6601 1358
rect 6613 1268 6617 1378
rect 6627 1356 6631 1396
rect 6622 1344 6625 1356
rect 6622 1280 6626 1344
rect 6647 1337 6651 1396
rect 6642 1329 6651 1337
rect 6642 1300 6646 1329
rect 6661 1314 6665 1396
rect 6681 1313 6685 1356
rect 6622 1276 6655 1280
rect 6621 1256 6623 1268
rect 6619 1244 6623 1256
rect 6629 1256 6631 1268
rect 6629 1244 6633 1256
rect 6651 1244 6655 1276
rect 6661 1244 6665 1302
rect 6681 1264 6685 1301
rect 2435 1220 2489 1224
rect 2566 1220 2570 1224
rect 2574 1220 2578 1224
rect 2594 1220 2598 1224
rect 2602 1220 2606 1224
rect 2654 1220 2658 1224
rect 2662 1220 2666 1224
rect 2682 1220 2686 1224
rect 2690 1220 2694 1224
rect 2806 1220 2810 1224
rect 2814 1220 2818 1224
rect 2834 1220 2838 1224
rect 2842 1220 2846 1224
rect 2891 1220 2895 1224
rect 2913 1220 2917 1224
rect 3006 1220 3010 1224
rect 3014 1220 3018 1224
rect 3034 1220 3038 1224
rect 3042 1220 3046 1224
rect 3105 1220 3109 1224
rect 3175 1220 3229 1224
rect 3275 1220 3279 1224
rect 3295 1220 3299 1224
rect 3305 1220 3309 1224
rect 3327 1220 3331 1224
rect 3337 1220 3341 1224
rect 3359 1220 3363 1224
rect 3405 1220 3409 1224
rect 3413 1220 3417 1224
rect 3433 1220 3437 1224
rect 3443 1220 3447 1224
rect 3465 1220 3469 1224
rect 3525 1220 3529 1224
rect 3545 1220 3549 1224
rect 3605 1220 3609 1224
rect 3625 1220 3629 1224
rect 3645 1220 3649 1224
rect 3665 1220 3669 1224
rect 3725 1220 3729 1224
rect 3745 1220 3749 1224
rect 3765 1220 3769 1224
rect 3825 1220 3829 1224
rect 3871 1220 3875 1224
rect 3893 1220 3897 1224
rect 3903 1220 3907 1224
rect 3923 1220 3927 1224
rect 3931 1220 3935 1224
rect 3977 1220 3981 1224
rect 3999 1220 4003 1224
rect 4009 1220 4013 1224
rect 4031 1220 4035 1224
rect 4041 1220 4045 1224
rect 4061 1220 4065 1224
rect 4111 1220 4115 1224
rect 4133 1220 4137 1224
rect 4143 1220 4147 1224
rect 4163 1220 4167 1224
rect 4171 1220 4175 1224
rect 4217 1220 4221 1224
rect 4239 1220 4243 1224
rect 4249 1220 4253 1224
rect 4271 1220 4275 1224
rect 4281 1220 4285 1224
rect 4301 1220 4305 1224
rect 4365 1220 4369 1224
rect 4414 1220 4418 1224
rect 4422 1220 4426 1224
rect 4442 1220 4446 1224
rect 4450 1220 4454 1224
rect 4531 1220 4585 1224
rect 4686 1220 4690 1224
rect 4694 1220 4698 1224
rect 4714 1220 4718 1224
rect 4722 1220 4726 1224
rect 4783 1220 4787 1224
rect 4805 1220 4809 1224
rect 4873 1220 4877 1224
rect 4883 1220 4887 1224
rect 4953 1220 4957 1224
rect 4963 1220 4967 1224
rect 5025 1220 5029 1224
rect 5045 1220 5049 1224
rect 5065 1220 5069 1224
rect 5085 1220 5089 1224
rect 5145 1220 5149 1224
rect 5165 1220 5169 1224
rect 5185 1220 5189 1224
rect 5205 1220 5209 1224
rect 5251 1220 5255 1224
rect 5333 1220 5337 1224
rect 5343 1220 5347 1224
rect 5391 1220 5395 1224
rect 5411 1220 5415 1224
rect 5431 1220 5435 1224
rect 5451 1220 5455 1224
rect 5532 1220 5536 1224
rect 5554 1220 5558 1224
rect 5562 1220 5566 1224
rect 5611 1220 5615 1224
rect 5671 1220 5725 1224
rect 5813 1220 5817 1224
rect 5823 1220 5827 1224
rect 5885 1220 5889 1224
rect 5905 1220 5909 1224
rect 5925 1220 5929 1224
rect 5985 1220 5989 1224
rect 6031 1220 6035 1224
rect 6051 1220 6055 1224
rect 6071 1220 6075 1224
rect 6131 1220 6135 1224
rect 6151 1220 6155 1224
rect 6171 1220 6175 1224
rect 6191 1220 6195 1224
rect 6251 1220 6255 1224
rect 6273 1220 6277 1224
rect 6283 1220 6287 1224
rect 6303 1220 6307 1224
rect 6311 1220 6315 1224
rect 6357 1220 6361 1224
rect 6379 1220 6383 1224
rect 6389 1220 6393 1224
rect 6411 1220 6415 1224
rect 6421 1220 6425 1224
rect 6441 1220 6445 1224
rect 6491 1220 6495 1224
rect 6513 1220 6517 1224
rect 6523 1220 6527 1224
rect 6543 1220 6547 1224
rect 6551 1220 6555 1224
rect 6597 1220 6601 1224
rect 6619 1220 6623 1224
rect 6629 1220 6633 1224
rect 6651 1220 6655 1224
rect 6661 1220 6665 1224
rect 6681 1220 6685 1224
rect 31 1196 35 1200
rect 53 1196 57 1200
rect 63 1196 67 1200
rect 83 1196 87 1200
rect 91 1196 95 1200
rect 137 1196 141 1200
rect 159 1196 163 1200
rect 169 1196 173 1200
rect 191 1196 195 1200
rect 201 1196 205 1200
rect 221 1196 225 1200
rect 285 1196 289 1200
rect 331 1196 335 1200
rect 353 1196 357 1200
rect 363 1196 367 1200
rect 383 1196 387 1200
rect 391 1196 395 1200
rect 437 1196 441 1200
rect 459 1196 463 1200
rect 469 1196 473 1200
rect 491 1196 495 1200
rect 501 1196 505 1200
rect 521 1196 525 1200
rect 571 1196 575 1200
rect 632 1196 636 1200
rect 640 1196 644 1200
rect 648 1196 652 1200
rect 731 1196 735 1200
rect 751 1196 755 1200
rect 812 1196 816 1200
rect 820 1196 824 1200
rect 828 1196 832 1200
rect 913 1196 917 1200
rect 923 1196 927 1200
rect 991 1196 995 1200
rect 1055 1196 1059 1200
rect 1075 1196 1079 1200
rect 1085 1196 1089 1200
rect 1107 1196 1111 1200
rect 1117 1196 1121 1200
rect 1139 1196 1143 1200
rect 1185 1196 1189 1200
rect 1193 1196 1197 1200
rect 1213 1196 1217 1200
rect 1223 1196 1227 1200
rect 1245 1196 1249 1200
rect 1291 1196 1295 1200
rect 1311 1196 1315 1200
rect 1331 1196 1335 1200
rect 1351 1196 1355 1200
rect 1371 1196 1375 1200
rect 1391 1196 1395 1200
rect 1411 1196 1415 1200
rect 1431 1196 1435 1200
rect 1495 1196 1499 1200
rect 1515 1196 1519 1200
rect 1525 1196 1529 1200
rect 1547 1196 1551 1200
rect 1557 1196 1561 1200
rect 1579 1196 1583 1200
rect 1625 1196 1629 1200
rect 1633 1196 1637 1200
rect 1653 1196 1657 1200
rect 1663 1196 1667 1200
rect 1685 1196 1689 1200
rect 1745 1196 1749 1200
rect 1765 1196 1769 1200
rect 1825 1196 1829 1200
rect 1845 1196 1849 1200
rect 1865 1196 1869 1200
rect 1885 1196 1889 1200
rect 1945 1196 1949 1200
rect 1965 1196 1969 1200
rect 1985 1196 1989 1200
rect 2045 1196 2049 1200
rect 2065 1196 2069 1200
rect 2085 1196 2089 1200
rect 2145 1196 2149 1200
rect 2165 1196 2169 1200
rect 2225 1196 2229 1200
rect 2245 1196 2249 1200
rect 2265 1196 2269 1200
rect 2285 1196 2289 1200
rect 2335 1196 2339 1200
rect 2355 1196 2359 1200
rect 2365 1196 2369 1200
rect 2387 1196 2391 1200
rect 2397 1196 2401 1200
rect 2419 1196 2423 1200
rect 2465 1196 2469 1200
rect 2473 1196 2477 1200
rect 2493 1196 2497 1200
rect 2503 1196 2507 1200
rect 2525 1196 2529 1200
rect 2585 1196 2589 1200
rect 2631 1196 2635 1200
rect 2651 1196 2655 1200
rect 2671 1196 2675 1200
rect 2743 1196 2747 1200
rect 2765 1196 2769 1200
rect 2811 1196 2815 1200
rect 2906 1196 2910 1200
rect 2914 1196 2918 1200
rect 2934 1196 2938 1200
rect 2942 1196 2946 1200
rect 2995 1196 2999 1200
rect 3015 1196 3019 1200
rect 3025 1196 3029 1200
rect 3047 1196 3051 1200
rect 3057 1196 3061 1200
rect 3079 1196 3083 1200
rect 3125 1196 3129 1200
rect 3133 1196 3137 1200
rect 3153 1196 3157 1200
rect 3163 1196 3167 1200
rect 3185 1196 3189 1200
rect 3233 1196 3237 1200
rect 3243 1196 3247 1200
rect 3335 1196 3389 1200
rect 31 1088 35 1156
rect 53 1127 57 1176
rect 63 1155 67 1176
rect 83 1164 87 1176
rect 91 1172 95 1176
rect 91 1168 125 1172
rect 83 1160 113 1164
rect 83 1159 101 1160
rect 63 1151 87 1155
rect 31 1076 33 1088
rect 31 1064 35 1076
rect 53 1069 57 1115
rect 49 1063 57 1069
rect 49 1034 53 1063
rect 81 1056 87 1151
rect 49 1027 57 1034
rect 53 1004 57 1027
rect 61 1004 65 1044
rect 81 1024 85 1056
rect 121 1042 125 1168
rect 137 1062 141 1176
rect 159 1164 163 1176
rect 161 1152 163 1164
rect 169 1164 173 1176
rect 169 1152 171 1164
rect 89 1030 113 1032
rect 89 1028 125 1030
rect 89 1024 93 1028
rect 135 1024 139 1050
rect 153 1042 157 1152
rect 191 1144 195 1176
rect 162 1140 195 1144
rect 162 1076 166 1140
rect 182 1091 186 1120
rect 201 1118 205 1176
rect 221 1119 225 1156
rect 285 1119 289 1176
rect 285 1107 294 1119
rect 182 1083 191 1091
rect 162 1064 165 1076
rect 155 1024 159 1030
rect 167 1024 171 1064
rect 187 1024 191 1083
rect 201 1024 205 1106
rect 221 1064 225 1107
rect 285 1024 289 1107
rect 331 1088 335 1156
rect 353 1127 357 1176
rect 363 1155 367 1176
rect 383 1164 387 1176
rect 391 1172 395 1176
rect 391 1168 425 1172
rect 383 1160 413 1164
rect 383 1159 401 1160
rect 363 1151 387 1155
rect 331 1076 333 1088
rect 331 1064 335 1076
rect 353 1069 357 1115
rect 349 1063 357 1069
rect 349 1034 353 1063
rect 381 1056 387 1151
rect 349 1027 357 1034
rect 353 1004 357 1027
rect 361 1004 365 1044
rect 381 1024 385 1056
rect 421 1042 425 1168
rect 437 1062 441 1176
rect 459 1164 463 1176
rect 461 1152 463 1164
rect 469 1164 473 1176
rect 469 1152 471 1164
rect 389 1030 413 1032
rect 389 1028 425 1030
rect 389 1024 393 1028
rect 435 1024 439 1050
rect 453 1042 457 1152
rect 491 1144 495 1176
rect 462 1140 495 1144
rect 462 1076 466 1140
rect 482 1091 486 1120
rect 501 1118 505 1176
rect 521 1119 525 1156
rect 571 1119 575 1176
rect 566 1107 575 1119
rect 482 1083 491 1091
rect 462 1064 465 1076
rect 455 1024 459 1030
rect 467 1024 471 1064
rect 487 1024 491 1083
rect 501 1024 505 1106
rect 521 1064 525 1107
rect 571 1024 575 1107
rect 632 1079 636 1136
rect 626 1067 636 1079
rect 620 1036 626 1067
rect 640 1059 644 1136
rect 648 1079 652 1136
rect 731 1099 735 1176
rect 751 1099 755 1176
rect 913 1136 917 1156
rect 726 1087 735 1099
rect 648 1067 655 1079
rect 667 1067 675 1079
rect 640 1040 646 1047
rect 640 1036 655 1040
rect 620 1032 635 1036
rect 631 1024 635 1032
rect 651 1024 655 1036
rect 671 1024 675 1067
rect 731 1064 735 1087
rect 739 1087 754 1099
rect 739 1064 743 1087
rect 812 1079 816 1136
rect 806 1067 816 1079
rect 800 1036 806 1067
rect 820 1059 824 1136
rect 828 1079 832 1136
rect 909 1129 917 1136
rect 923 1136 927 1156
rect 923 1129 937 1136
rect 909 1113 915 1129
rect 906 1101 915 1113
rect 828 1067 835 1079
rect 847 1067 855 1079
rect 820 1040 826 1047
rect 820 1036 835 1040
rect 800 1032 815 1036
rect 811 1024 815 1032
rect 831 1024 835 1036
rect 851 1024 855 1067
rect 911 1024 915 1101
rect 931 1113 937 1129
rect 991 1119 995 1176
rect 1055 1119 1059 1156
rect 931 1101 934 1113
rect 986 1107 995 1119
rect 1075 1118 1079 1176
rect 1085 1144 1089 1176
rect 1107 1164 1111 1176
rect 1109 1152 1111 1164
rect 1117 1164 1121 1176
rect 1117 1152 1119 1164
rect 1085 1140 1118 1144
rect 931 1024 935 1101
rect 991 1024 995 1107
rect 1055 1064 1059 1107
rect 1075 1024 1079 1106
rect 1094 1091 1098 1120
rect 1089 1083 1098 1091
rect 1089 1024 1093 1083
rect 1114 1076 1118 1140
rect 1115 1064 1118 1076
rect 1109 1024 1113 1064
rect 1123 1042 1127 1152
rect 1139 1062 1143 1176
rect 1185 1172 1189 1176
rect 1155 1168 1189 1172
rect 1121 1024 1125 1030
rect 1141 1024 1145 1050
rect 1155 1042 1159 1168
rect 1193 1164 1197 1176
rect 1167 1160 1197 1164
rect 1179 1159 1197 1160
rect 1213 1155 1217 1176
rect 1193 1151 1217 1155
rect 1193 1056 1199 1151
rect 1223 1127 1227 1176
rect 1223 1069 1227 1115
rect 1245 1088 1249 1156
rect 1247 1076 1249 1088
rect 1223 1063 1231 1069
rect 1245 1064 1249 1076
rect 1291 1133 1295 1156
rect 1311 1133 1315 1156
rect 1331 1136 1335 1156
rect 1351 1136 1355 1156
rect 1371 1136 1375 1156
rect 1391 1136 1395 1156
rect 1411 1136 1415 1156
rect 1431 1136 1435 1156
rect 1291 1121 1294 1133
rect 1306 1121 1315 1133
rect 1342 1124 1355 1136
rect 1382 1124 1395 1136
rect 1422 1124 1435 1136
rect 1291 1064 1295 1121
rect 1311 1064 1315 1121
rect 1331 1064 1335 1124
rect 1351 1064 1355 1124
rect 1371 1064 1375 1124
rect 1391 1064 1395 1124
rect 1411 1064 1415 1124
rect 1431 1064 1435 1124
rect 1495 1119 1499 1156
rect 1515 1118 1519 1176
rect 1525 1144 1529 1176
rect 1547 1164 1551 1176
rect 1549 1152 1551 1164
rect 1557 1164 1561 1176
rect 1557 1152 1559 1164
rect 1525 1140 1558 1144
rect 1495 1064 1499 1107
rect 1167 1030 1191 1032
rect 1155 1028 1191 1030
rect 1187 1024 1191 1028
rect 1195 1024 1199 1056
rect 1215 1004 1219 1044
rect 1227 1034 1231 1063
rect 1223 1027 1231 1034
rect 1223 1004 1227 1027
rect 1515 1024 1519 1106
rect 1534 1091 1538 1120
rect 1529 1083 1538 1091
rect 1529 1024 1533 1083
rect 1554 1076 1558 1140
rect 1555 1064 1558 1076
rect 1549 1024 1553 1064
rect 1563 1042 1567 1152
rect 1579 1062 1583 1176
rect 1625 1172 1629 1176
rect 1595 1168 1629 1172
rect 1561 1024 1565 1030
rect 1581 1024 1585 1050
rect 1595 1042 1599 1168
rect 1633 1164 1637 1176
rect 1607 1160 1637 1164
rect 1619 1159 1637 1160
rect 1653 1155 1657 1176
rect 1633 1151 1657 1155
rect 1633 1056 1639 1151
rect 1663 1127 1667 1176
rect 1663 1069 1667 1115
rect 1685 1088 1689 1156
rect 1745 1099 1749 1176
rect 1765 1099 1769 1176
rect 1825 1099 1829 1156
rect 1845 1133 1849 1156
rect 1865 1133 1869 1156
rect 1885 1149 1889 1156
rect 1885 1145 1900 1149
rect 1865 1121 1874 1133
rect 1687 1076 1689 1088
rect 1746 1087 1761 1099
rect 1663 1063 1671 1069
rect 1685 1064 1689 1076
rect 1757 1064 1761 1087
rect 1765 1087 1774 1099
rect 1827 1087 1829 1099
rect 1765 1064 1769 1087
rect 1825 1072 1829 1087
rect 1825 1068 1839 1072
rect 1835 1064 1839 1068
rect 1845 1064 1849 1121
rect 1865 1072 1871 1121
rect 1894 1099 1900 1145
rect 1894 1072 1899 1087
rect 1945 1079 1949 1156
rect 1965 1133 1969 1156
rect 1985 1151 1989 1156
rect 1985 1144 1998 1151
rect 1965 1121 1974 1133
rect 1865 1068 1879 1072
rect 1875 1064 1879 1068
rect 1885 1068 1899 1072
rect 1885 1064 1889 1068
rect 1947 1067 1954 1079
rect 1607 1030 1631 1032
rect 1595 1028 1631 1030
rect 1627 1024 1631 1028
rect 1635 1024 1639 1056
rect 1655 1004 1659 1044
rect 1667 1034 1671 1063
rect 1663 1027 1671 1034
rect 1663 1004 1667 1027
rect 1950 1024 1954 1067
rect 1972 1064 1976 1121
rect 1994 1099 1998 1144
rect 1994 1076 1998 1087
rect 2045 1079 2049 1156
rect 2065 1133 2069 1156
rect 2085 1151 2089 1156
rect 2085 1144 2098 1151
rect 2065 1121 2074 1133
rect 1980 1068 1998 1076
rect 1980 1064 1984 1068
rect 2047 1067 2054 1079
rect 2050 1024 2054 1067
rect 2072 1064 2076 1121
rect 2094 1099 2098 1144
rect 2145 1099 2149 1176
rect 2165 1099 2169 1176
rect 2225 1099 2229 1156
rect 2245 1133 2249 1156
rect 2265 1133 2269 1156
rect 2285 1149 2289 1156
rect 2285 1145 2300 1149
rect 2265 1121 2274 1133
rect 2146 1087 2161 1099
rect 2094 1076 2098 1087
rect 2080 1068 2098 1076
rect 2080 1064 2084 1068
rect 2157 1064 2161 1087
rect 2165 1087 2174 1099
rect 2227 1087 2229 1099
rect 2165 1064 2169 1087
rect 2225 1072 2229 1087
rect 2225 1068 2239 1072
rect 2235 1064 2239 1068
rect 2245 1064 2249 1121
rect 2265 1072 2271 1121
rect 2294 1099 2300 1145
rect 2335 1119 2339 1156
rect 2355 1118 2359 1176
rect 2365 1144 2369 1176
rect 2387 1164 2391 1176
rect 2389 1152 2391 1164
rect 2397 1164 2401 1176
rect 2397 1152 2399 1164
rect 2365 1140 2398 1144
rect 2294 1072 2299 1087
rect 2265 1068 2279 1072
rect 2275 1064 2279 1068
rect 2285 1068 2299 1072
rect 2285 1064 2289 1068
rect 2335 1064 2339 1107
rect 2355 1024 2359 1106
rect 2374 1091 2378 1120
rect 2369 1083 2378 1091
rect 2369 1024 2373 1083
rect 2394 1076 2398 1140
rect 2395 1064 2398 1076
rect 2389 1024 2393 1064
rect 2403 1042 2407 1152
rect 2419 1062 2423 1176
rect 2465 1172 2469 1176
rect 2435 1168 2469 1172
rect 2401 1024 2405 1030
rect 2421 1024 2425 1050
rect 2435 1042 2439 1168
rect 2473 1164 2477 1176
rect 2447 1160 2477 1164
rect 2459 1159 2477 1160
rect 2493 1155 2497 1176
rect 2473 1151 2497 1155
rect 2473 1056 2479 1151
rect 2503 1127 2507 1176
rect 2503 1069 2507 1115
rect 2525 1088 2529 1156
rect 2527 1076 2529 1088
rect 2503 1063 2511 1069
rect 2525 1064 2529 1076
rect 2585 1119 2589 1176
rect 2631 1151 2635 1156
rect 2622 1144 2635 1151
rect 2585 1107 2594 1119
rect 2447 1030 2471 1032
rect 2435 1028 2471 1030
rect 2467 1024 2471 1028
rect 2475 1024 2479 1056
rect 2495 1004 2499 1044
rect 2507 1034 2511 1063
rect 2503 1027 2511 1034
rect 2503 1004 2507 1027
rect 2585 1024 2589 1107
rect 2622 1099 2626 1144
rect 2651 1133 2655 1156
rect 2646 1121 2655 1133
rect 2622 1076 2626 1087
rect 2622 1068 2640 1076
rect 2636 1064 2640 1068
rect 2644 1064 2648 1121
rect 2671 1079 2675 1156
rect 2743 1150 2747 1156
rect 2743 1138 2745 1150
rect 2765 1099 2769 1176
rect 2811 1119 2815 1176
rect 2906 1151 2910 1156
rect 2806 1107 2815 1119
rect 2765 1087 2774 1099
rect 2666 1067 2673 1079
rect 2743 1070 2745 1082
rect 2666 1024 2670 1067
rect 2743 1064 2747 1070
rect 2765 1024 2769 1087
rect 2811 1024 2815 1107
rect 2880 1147 2910 1151
rect 2880 1099 2886 1147
rect 2914 1142 2918 1156
rect 2905 1135 2918 1142
rect 2905 1133 2909 1135
rect 2934 1133 2938 1156
rect 2942 1148 2946 1156
rect 2942 1141 2959 1148
rect 2907 1121 2909 1133
rect 2886 1087 2889 1099
rect 2885 1064 2889 1087
rect 2905 1064 2909 1121
rect 2934 1092 2938 1121
rect 2953 1099 2959 1141
rect 2995 1119 2999 1156
rect 3015 1118 3019 1176
rect 3025 1144 3029 1176
rect 3047 1164 3051 1176
rect 3049 1152 3051 1164
rect 3057 1164 3061 1176
rect 3057 1152 3059 1164
rect 3025 1140 3058 1144
rect 2925 1086 2938 1092
rect 2945 1087 2953 1092
rect 2945 1086 2965 1087
rect 2925 1064 2929 1086
rect 2945 1064 2949 1086
rect 2995 1064 2999 1107
rect 3015 1024 3019 1106
rect 3034 1091 3038 1120
rect 3029 1083 3038 1091
rect 3029 1024 3033 1083
rect 3054 1076 3058 1140
rect 3055 1064 3058 1076
rect 3049 1024 3053 1064
rect 3063 1042 3067 1152
rect 3079 1062 3083 1176
rect 3125 1172 3129 1176
rect 3095 1168 3129 1172
rect 3061 1024 3065 1030
rect 3081 1024 3085 1050
rect 3095 1042 3099 1168
rect 3133 1164 3137 1176
rect 3107 1160 3137 1164
rect 3119 1159 3137 1160
rect 3153 1155 3157 1176
rect 3133 1151 3157 1155
rect 3133 1056 3139 1151
rect 3163 1127 3167 1176
rect 3325 1188 3329 1192
rect 3335 1188 3339 1196
rect 3355 1188 3359 1192
rect 3365 1188 3369 1192
rect 3385 1188 3389 1196
rect 3431 1196 3485 1200
rect 3563 1196 3567 1200
rect 3585 1196 3589 1200
rect 3635 1196 3639 1200
rect 3655 1196 3659 1200
rect 3665 1196 3669 1200
rect 3687 1196 3691 1200
rect 3697 1196 3701 1200
rect 3719 1196 3723 1200
rect 3765 1196 3769 1200
rect 3773 1196 3777 1200
rect 3793 1196 3797 1200
rect 3803 1196 3807 1200
rect 3825 1196 3829 1200
rect 3871 1196 3925 1200
rect 3431 1188 3435 1196
rect 3451 1188 3455 1192
rect 3461 1188 3465 1192
rect 3481 1188 3485 1196
rect 3491 1188 3495 1192
rect 3163 1069 3167 1115
rect 3185 1088 3189 1156
rect 3233 1136 3237 1156
rect 3229 1129 3237 1136
rect 3243 1136 3247 1156
rect 3385 1164 3389 1168
rect 3431 1164 3435 1168
rect 3385 1159 3397 1164
rect 3243 1129 3257 1136
rect 3229 1113 3235 1129
rect 3226 1101 3235 1113
rect 3187 1076 3189 1088
rect 3163 1063 3171 1069
rect 3185 1064 3189 1076
rect 3107 1030 3131 1032
rect 3095 1028 3131 1030
rect 3127 1024 3131 1028
rect 3135 1024 3139 1056
rect 3155 1004 3159 1044
rect 3167 1034 3171 1063
rect 3163 1027 3171 1034
rect 3163 1004 3167 1027
rect 3231 1024 3235 1101
rect 3251 1113 3257 1129
rect 3251 1101 3254 1113
rect 3251 1024 3255 1101
rect 3325 1099 3329 1148
rect 3335 1144 3339 1148
rect 3355 1102 3359 1148
rect 3365 1136 3369 1148
rect 3365 1130 3379 1136
rect 3326 1087 3329 1099
rect 3374 1099 3379 1130
rect 3393 1133 3397 1159
rect 3423 1159 3435 1164
rect 3423 1133 3427 1159
rect 3563 1150 3567 1156
rect 3451 1136 3455 1148
rect 3325 1064 3329 1087
rect 3335 1086 3365 1090
rect 3335 1064 3339 1086
rect 3373 1081 3378 1087
rect 3365 1077 3378 1081
rect 3355 1072 3359 1076
rect 3365 1072 3369 1077
rect 3393 1040 3397 1121
rect 3385 1036 3397 1040
rect 3423 1040 3427 1121
rect 3441 1130 3455 1136
rect 3441 1099 3446 1130
rect 3461 1102 3465 1148
rect 3481 1144 3485 1148
rect 3442 1081 3447 1087
rect 3491 1099 3495 1148
rect 3563 1138 3565 1150
rect 3585 1099 3589 1176
rect 3635 1119 3639 1156
rect 3655 1118 3659 1176
rect 3665 1144 3669 1176
rect 3687 1164 3691 1176
rect 3689 1152 3691 1164
rect 3697 1164 3701 1176
rect 3697 1152 3699 1164
rect 3665 1140 3698 1144
rect 3455 1086 3485 1090
rect 3442 1077 3455 1081
rect 3451 1072 3455 1077
rect 3461 1072 3465 1076
rect 3423 1036 3435 1040
rect 3385 1032 3389 1036
rect 3431 1032 3435 1036
rect 3481 1064 3485 1086
rect 3491 1087 3494 1099
rect 3585 1087 3594 1099
rect 3491 1064 3495 1087
rect 3563 1070 3565 1082
rect 3563 1064 3567 1070
rect 3355 984 3359 992
rect 3365 988 3369 992
rect 3385 984 3389 992
rect 31 980 35 984
rect 53 980 57 984
rect 61 980 65 984
rect 81 980 85 984
rect 89 980 93 984
rect 135 980 139 984
rect 155 980 159 984
rect 167 980 171 984
rect 187 980 191 984
rect 201 980 205 984
rect 221 980 225 984
rect 285 980 289 984
rect 331 980 335 984
rect 353 980 357 984
rect 361 980 365 984
rect 381 980 385 984
rect 389 980 393 984
rect 435 980 439 984
rect 455 980 459 984
rect 467 980 471 984
rect 487 980 491 984
rect 501 980 505 984
rect 521 980 525 984
rect 571 980 575 984
rect 631 980 635 984
rect 651 980 655 984
rect 671 980 675 984
rect 731 980 735 984
rect 739 980 743 984
rect 811 980 815 984
rect 831 980 835 984
rect 851 980 855 984
rect 911 980 915 984
rect 931 980 935 984
rect 991 980 995 984
rect 1055 980 1059 984
rect 1075 980 1079 984
rect 1089 980 1093 984
rect 1109 980 1113 984
rect 1121 980 1125 984
rect 1141 980 1145 984
rect 1187 980 1191 984
rect 1195 980 1199 984
rect 1215 980 1219 984
rect 1223 980 1227 984
rect 1245 980 1249 984
rect 1291 980 1295 984
rect 1311 980 1315 984
rect 1331 980 1335 984
rect 1351 980 1355 984
rect 1371 980 1375 984
rect 1391 980 1395 984
rect 1411 980 1415 984
rect 1431 980 1435 984
rect 1495 980 1499 984
rect 1515 980 1519 984
rect 1529 980 1533 984
rect 1549 980 1553 984
rect 1561 980 1565 984
rect 1581 980 1585 984
rect 1627 980 1631 984
rect 1635 980 1639 984
rect 1655 980 1659 984
rect 1663 980 1667 984
rect 1685 980 1689 984
rect 1757 980 1761 984
rect 1765 980 1769 984
rect 1835 980 1839 984
rect 1845 980 1849 984
rect 1875 980 1879 984
rect 1885 980 1889 984
rect 1950 980 1954 984
rect 1972 980 1976 984
rect 1980 980 1984 984
rect 2050 980 2054 984
rect 2072 980 2076 984
rect 2080 980 2084 984
rect 2157 980 2161 984
rect 2165 980 2169 984
rect 2235 980 2239 984
rect 2245 980 2249 984
rect 2275 980 2279 984
rect 2285 980 2289 984
rect 2335 980 2339 984
rect 2355 980 2359 984
rect 2369 980 2373 984
rect 2389 980 2393 984
rect 2401 980 2405 984
rect 2421 980 2425 984
rect 2467 980 2471 984
rect 2475 980 2479 984
rect 2495 980 2499 984
rect 2503 980 2507 984
rect 2525 980 2529 984
rect 2585 980 2589 984
rect 2636 980 2640 984
rect 2644 980 2648 984
rect 2666 980 2670 984
rect 2743 980 2747 984
rect 2765 980 2769 984
rect 2811 980 2815 984
rect 2885 980 2889 984
rect 2905 980 2909 984
rect 2925 980 2929 984
rect 2945 980 2949 984
rect 2995 980 2999 984
rect 3015 980 3019 984
rect 3029 980 3033 984
rect 3049 980 3053 984
rect 3061 980 3065 984
rect 3081 980 3085 984
rect 3127 980 3131 984
rect 3135 980 3139 984
rect 3155 980 3159 984
rect 3163 980 3167 984
rect 3185 980 3189 984
rect 3231 980 3235 984
rect 3251 980 3255 984
rect 3325 980 3329 984
rect 3335 980 3339 984
rect 3355 980 3389 984
rect 3431 984 3435 992
rect 3451 988 3455 992
rect 3461 984 3465 992
rect 3585 1024 3589 1087
rect 3635 1064 3639 1107
rect 3655 1024 3659 1106
rect 3674 1091 3678 1120
rect 3669 1083 3678 1091
rect 3669 1024 3673 1083
rect 3694 1076 3698 1140
rect 3695 1064 3698 1076
rect 3689 1024 3693 1064
rect 3703 1042 3707 1152
rect 3719 1062 3723 1176
rect 3765 1172 3769 1176
rect 3735 1168 3769 1172
rect 3701 1024 3705 1030
rect 3721 1024 3725 1050
rect 3735 1042 3739 1168
rect 3773 1164 3777 1176
rect 3747 1160 3777 1164
rect 3759 1159 3777 1160
rect 3793 1155 3797 1176
rect 3773 1151 3797 1155
rect 3773 1056 3779 1151
rect 3803 1127 3807 1176
rect 3871 1188 3875 1196
rect 3891 1188 3895 1192
rect 3901 1188 3905 1192
rect 3921 1188 3925 1196
rect 4015 1196 4069 1200
rect 4111 1196 4115 1200
rect 4171 1196 4175 1200
rect 4191 1196 4195 1200
rect 4211 1196 4215 1200
rect 4231 1196 4235 1200
rect 4291 1196 4295 1200
rect 4311 1196 4315 1200
rect 4385 1196 4389 1200
rect 4405 1196 4409 1200
rect 4425 1196 4429 1200
rect 4492 1196 4496 1200
rect 4514 1196 4518 1200
rect 4522 1196 4526 1200
rect 4575 1196 4579 1200
rect 4595 1196 4599 1200
rect 4605 1196 4609 1200
rect 4627 1196 4631 1200
rect 4637 1196 4641 1200
rect 4659 1196 4663 1200
rect 4705 1196 4709 1200
rect 4713 1196 4717 1200
rect 4733 1196 4737 1200
rect 4743 1196 4747 1200
rect 4765 1196 4769 1200
rect 4811 1196 4815 1200
rect 4831 1196 4835 1200
rect 4851 1196 4855 1200
rect 4871 1196 4875 1200
rect 4945 1196 4949 1200
rect 4965 1196 4969 1200
rect 5025 1196 5029 1200
rect 5045 1196 5049 1200
rect 5065 1196 5069 1200
rect 5125 1196 5129 1200
rect 5145 1196 5149 1200
rect 5191 1196 5195 1200
rect 5211 1196 5215 1200
rect 5271 1196 5275 1200
rect 5291 1196 5295 1200
rect 5363 1196 5367 1200
rect 5385 1196 5389 1200
rect 5431 1196 5435 1200
rect 5451 1196 5455 1200
rect 5511 1196 5515 1200
rect 5531 1196 5535 1200
rect 5594 1196 5598 1200
rect 5602 1196 5606 1200
rect 5624 1196 5628 1200
rect 5691 1196 5695 1200
rect 5711 1196 5715 1200
rect 5731 1196 5735 1200
rect 5805 1196 5809 1200
rect 5825 1196 5829 1200
rect 5871 1196 5875 1200
rect 5891 1196 5895 1200
rect 5911 1196 5915 1200
rect 6008 1196 6012 1200
rect 6016 1196 6020 1200
rect 6024 1196 6028 1200
rect 6071 1196 6075 1200
rect 6091 1196 6095 1200
rect 6111 1196 6115 1200
rect 6185 1196 6189 1200
rect 6205 1196 6209 1200
rect 6251 1196 6255 1200
rect 6271 1196 6275 1200
rect 6331 1196 6335 1200
rect 6353 1196 6357 1200
rect 6363 1196 6367 1200
rect 6383 1196 6387 1200
rect 6391 1196 6395 1200
rect 6437 1196 6441 1200
rect 6459 1196 6463 1200
rect 6469 1196 6473 1200
rect 6491 1196 6495 1200
rect 6501 1196 6505 1200
rect 6521 1196 6525 1200
rect 6571 1196 6575 1200
rect 6591 1196 6595 1200
rect 6611 1196 6615 1200
rect 6631 1196 6635 1200
rect 3931 1188 3935 1192
rect 4005 1188 4009 1192
rect 4015 1188 4019 1196
rect 4035 1188 4039 1192
rect 4045 1188 4049 1192
rect 4065 1188 4069 1196
rect 3871 1164 3875 1168
rect 3863 1159 3875 1164
rect 3803 1069 3807 1115
rect 3825 1088 3829 1156
rect 3863 1133 3867 1159
rect 4065 1164 4069 1168
rect 4065 1159 4077 1164
rect 3891 1136 3895 1148
rect 3827 1076 3829 1088
rect 3803 1063 3811 1069
rect 3825 1064 3829 1076
rect 3747 1030 3771 1032
rect 3735 1028 3771 1030
rect 3767 1024 3771 1028
rect 3775 1024 3779 1056
rect 3795 1004 3799 1044
rect 3807 1034 3811 1063
rect 3803 1027 3811 1034
rect 3803 1004 3807 1027
rect 3863 1040 3867 1121
rect 3881 1130 3895 1136
rect 3881 1099 3886 1130
rect 3901 1102 3905 1148
rect 3921 1144 3925 1148
rect 3882 1081 3887 1087
rect 3931 1099 3935 1148
rect 4005 1099 4009 1148
rect 4015 1144 4019 1148
rect 4035 1102 4039 1148
rect 4045 1136 4049 1148
rect 4045 1130 4059 1136
rect 3895 1086 3925 1090
rect 3882 1077 3895 1081
rect 3891 1072 3895 1077
rect 3901 1072 3905 1076
rect 3863 1036 3875 1040
rect 3871 1032 3875 1036
rect 3921 1064 3925 1086
rect 3931 1087 3934 1099
rect 4006 1087 4009 1099
rect 4054 1099 4059 1130
rect 4073 1133 4077 1159
rect 3931 1064 3935 1087
rect 4005 1064 4009 1087
rect 4015 1086 4045 1090
rect 4015 1064 4019 1086
rect 4053 1081 4058 1087
rect 4045 1077 4058 1081
rect 4035 1072 4039 1076
rect 4045 1072 4049 1077
rect 3871 984 3875 992
rect 3891 988 3895 992
rect 3901 984 3905 992
rect 4073 1040 4077 1121
rect 4111 1119 4115 1176
rect 4171 1149 4175 1156
rect 4106 1107 4115 1119
rect 4065 1036 4077 1040
rect 4065 1032 4069 1036
rect 4111 1024 4115 1107
rect 4160 1145 4175 1149
rect 4160 1099 4166 1145
rect 4191 1133 4195 1156
rect 4211 1133 4215 1156
rect 4186 1121 4195 1133
rect 4161 1072 4166 1087
rect 4189 1072 4195 1121
rect 4161 1068 4175 1072
rect 4171 1064 4175 1068
rect 4181 1068 4195 1072
rect 4181 1064 4185 1068
rect 4211 1064 4215 1121
rect 4231 1099 4235 1156
rect 4291 1099 4295 1176
rect 4311 1099 4315 1176
rect 4231 1087 4233 1099
rect 4286 1087 4295 1099
rect 4231 1072 4235 1087
rect 4221 1068 4235 1072
rect 4221 1064 4225 1068
rect 4291 1064 4295 1087
rect 4299 1087 4314 1099
rect 4299 1064 4303 1087
rect 4385 1079 4389 1156
rect 4405 1133 4409 1156
rect 4425 1151 4429 1156
rect 4425 1144 4438 1151
rect 4405 1121 4414 1133
rect 4387 1067 4394 1079
rect 4035 984 4039 992
rect 4045 988 4049 992
rect 4065 984 4069 992
rect 4390 1024 4394 1067
rect 4412 1064 4416 1121
rect 4434 1099 4438 1144
rect 4492 1133 4496 1176
rect 4485 1121 4494 1133
rect 4434 1076 4438 1087
rect 4420 1068 4438 1076
rect 4420 1064 4424 1068
rect 4485 1064 4489 1121
rect 4514 1119 4518 1156
rect 4522 1152 4526 1156
rect 4522 1146 4541 1152
rect 4534 1133 4541 1146
rect 4514 1084 4520 1107
rect 4534 1084 4541 1121
rect 4575 1119 4579 1156
rect 4595 1118 4599 1176
rect 4605 1144 4609 1176
rect 4627 1164 4631 1176
rect 4629 1152 4631 1164
rect 4637 1164 4641 1176
rect 4637 1152 4639 1164
rect 4605 1140 4638 1144
rect 4505 1078 4520 1084
rect 4525 1078 4541 1084
rect 4505 1064 4509 1078
rect 4525 1064 4529 1078
rect 4575 1064 4579 1107
rect 4595 1024 4599 1106
rect 4614 1091 4618 1120
rect 4609 1083 4618 1091
rect 4609 1024 4613 1083
rect 4634 1076 4638 1140
rect 4635 1064 4638 1076
rect 4629 1024 4633 1064
rect 4643 1042 4647 1152
rect 4659 1062 4663 1176
rect 4705 1172 4709 1176
rect 4675 1168 4709 1172
rect 4641 1024 4645 1030
rect 4661 1024 4665 1050
rect 4675 1042 4679 1168
rect 4713 1164 4717 1176
rect 4687 1160 4717 1164
rect 4699 1159 4717 1160
rect 4733 1155 4737 1176
rect 4713 1151 4737 1155
rect 4713 1056 4719 1151
rect 4743 1127 4747 1176
rect 4743 1069 4747 1115
rect 4765 1088 4769 1156
rect 4811 1149 4815 1156
rect 4800 1145 4815 1149
rect 4800 1099 4806 1145
rect 4831 1133 4835 1156
rect 4851 1133 4855 1156
rect 4826 1121 4835 1133
rect 4767 1076 4769 1088
rect 4743 1063 4751 1069
rect 4765 1064 4769 1076
rect 4801 1072 4806 1087
rect 4829 1072 4835 1121
rect 4801 1068 4815 1072
rect 4811 1064 4815 1068
rect 4821 1068 4835 1072
rect 4821 1064 4825 1068
rect 4851 1064 4855 1121
rect 4871 1099 4875 1156
rect 4945 1099 4949 1176
rect 4965 1099 4969 1176
rect 4871 1087 4873 1099
rect 4946 1087 4961 1099
rect 4871 1072 4875 1087
rect 4861 1068 4875 1072
rect 4861 1064 4865 1068
rect 4957 1064 4961 1087
rect 4965 1087 4974 1099
rect 4965 1064 4969 1087
rect 5025 1079 5029 1156
rect 5045 1133 5049 1156
rect 5065 1151 5069 1156
rect 5065 1144 5078 1151
rect 5045 1121 5054 1133
rect 5027 1067 5034 1079
rect 4687 1030 4711 1032
rect 4675 1028 4711 1030
rect 4707 1024 4711 1028
rect 4715 1024 4719 1056
rect 4735 1004 4739 1044
rect 4747 1034 4751 1063
rect 4743 1027 4751 1034
rect 4743 1004 4747 1027
rect 5030 1024 5034 1067
rect 5052 1064 5056 1121
rect 5074 1099 5078 1144
rect 5125 1099 5129 1176
rect 5145 1099 5149 1176
rect 5191 1099 5195 1176
rect 5211 1099 5215 1176
rect 5271 1099 5275 1176
rect 5291 1099 5295 1176
rect 5363 1150 5367 1156
rect 5363 1138 5365 1150
rect 5385 1099 5389 1176
rect 5431 1099 5435 1176
rect 5451 1099 5455 1176
rect 5511 1099 5515 1176
rect 5531 1099 5535 1176
rect 5594 1152 5598 1156
rect 5579 1146 5598 1152
rect 5579 1133 5586 1146
rect 5126 1087 5141 1099
rect 5074 1076 5078 1087
rect 5060 1068 5078 1076
rect 5060 1064 5064 1068
rect 5137 1064 5141 1087
rect 5145 1087 5154 1099
rect 5186 1087 5195 1099
rect 5145 1064 5149 1087
rect 5191 1064 5195 1087
rect 5199 1087 5214 1099
rect 5266 1087 5275 1099
rect 5199 1064 5203 1087
rect 5271 1064 5275 1087
rect 5279 1087 5294 1099
rect 5385 1087 5394 1099
rect 5426 1087 5435 1099
rect 5279 1064 5283 1087
rect 5363 1070 5365 1082
rect 5363 1064 5367 1070
rect 5385 1024 5389 1087
rect 5431 1064 5435 1087
rect 5439 1087 5454 1099
rect 5506 1087 5515 1099
rect 5439 1064 5443 1087
rect 5511 1064 5515 1087
rect 5519 1087 5534 1099
rect 5519 1064 5523 1087
rect 5579 1084 5586 1121
rect 5602 1119 5606 1156
rect 5624 1133 5628 1176
rect 5691 1169 5695 1176
rect 5711 1169 5715 1176
rect 5682 1164 5695 1169
rect 5626 1121 5635 1133
rect 5600 1084 5606 1107
rect 5579 1078 5595 1084
rect 5600 1078 5615 1084
rect 5591 1064 5595 1078
rect 5611 1064 5615 1078
rect 5631 1064 5635 1121
rect 5682 1119 5686 1164
rect 5682 1073 5686 1107
rect 5701 1163 5715 1169
rect 5701 1099 5705 1163
rect 5731 1148 5735 1156
rect 5725 1136 5735 1148
rect 5805 1099 5809 1176
rect 5825 1099 5829 1176
rect 5871 1151 5875 1156
rect 5862 1144 5875 1151
rect 5862 1099 5866 1144
rect 5891 1133 5895 1156
rect 5886 1121 5895 1133
rect 5806 1087 5821 1099
rect 5682 1068 5695 1073
rect 5691 1064 5695 1068
rect 5701 1064 5705 1087
rect 5721 1064 5725 1069
rect 5817 1064 5821 1087
rect 5825 1087 5834 1099
rect 5825 1064 5829 1087
rect 5862 1076 5866 1087
rect 5862 1068 5880 1076
rect 5876 1064 5880 1068
rect 5884 1064 5888 1121
rect 5911 1079 5915 1156
rect 6071 1151 6075 1156
rect 6062 1144 6075 1151
rect 6008 1079 6012 1136
rect 5906 1067 5913 1079
rect 5985 1067 5993 1079
rect 6005 1067 6012 1079
rect 5906 1024 5910 1067
rect 5985 1024 5989 1067
rect 6016 1059 6020 1136
rect 6024 1079 6028 1136
rect 6062 1099 6066 1144
rect 6091 1133 6095 1156
rect 6086 1121 6095 1133
rect 6024 1067 6034 1079
rect 6062 1076 6066 1087
rect 6062 1068 6080 1076
rect 6014 1040 6020 1047
rect 6005 1036 6020 1040
rect 6034 1036 6040 1067
rect 6076 1064 6080 1068
rect 6084 1064 6088 1121
rect 6111 1079 6115 1156
rect 6185 1099 6189 1176
rect 6205 1099 6209 1176
rect 6251 1099 6255 1176
rect 6271 1099 6275 1176
rect 6186 1087 6201 1099
rect 6106 1067 6113 1079
rect 6005 1024 6009 1036
rect 6025 1032 6040 1036
rect 6025 1024 6029 1032
rect 6106 1024 6110 1067
rect 6197 1064 6201 1087
rect 6205 1087 6214 1099
rect 6246 1087 6255 1099
rect 6205 1064 6209 1087
rect 6251 1064 6255 1087
rect 6259 1087 6274 1099
rect 6331 1088 6335 1156
rect 6353 1127 6357 1176
rect 6363 1155 6367 1176
rect 6383 1164 6387 1176
rect 6391 1172 6395 1176
rect 6391 1168 6425 1172
rect 6383 1160 6413 1164
rect 6383 1159 6401 1160
rect 6363 1151 6387 1155
rect 6259 1064 6263 1087
rect 6331 1076 6333 1088
rect 6331 1064 6335 1076
rect 6353 1069 6357 1115
rect 6349 1063 6357 1069
rect 6349 1034 6353 1063
rect 6381 1056 6387 1151
rect 6349 1027 6357 1034
rect 6353 1004 6357 1027
rect 6361 1004 6365 1044
rect 6381 1024 6385 1056
rect 6421 1042 6425 1168
rect 6437 1062 6441 1176
rect 6459 1164 6463 1176
rect 6461 1152 6463 1164
rect 6469 1164 6473 1176
rect 6469 1152 6471 1164
rect 6389 1030 6413 1032
rect 6389 1028 6425 1030
rect 6389 1024 6393 1028
rect 6435 1024 6439 1050
rect 6453 1042 6457 1152
rect 6491 1144 6495 1176
rect 6462 1140 6495 1144
rect 6462 1076 6466 1140
rect 6482 1091 6486 1120
rect 6501 1118 6505 1176
rect 6521 1119 6525 1156
rect 6571 1149 6575 1156
rect 6560 1145 6575 1149
rect 6482 1083 6491 1091
rect 6462 1064 6465 1076
rect 6455 1024 6459 1030
rect 6467 1024 6471 1064
rect 6487 1024 6491 1083
rect 6501 1024 6505 1106
rect 6521 1064 6525 1107
rect 6560 1099 6566 1145
rect 6591 1133 6595 1156
rect 6611 1133 6615 1156
rect 6586 1121 6595 1133
rect 6561 1072 6566 1087
rect 6589 1072 6595 1121
rect 6561 1068 6575 1072
rect 6571 1064 6575 1068
rect 6581 1068 6595 1072
rect 6581 1064 6585 1068
rect 6611 1064 6615 1121
rect 6631 1099 6635 1156
rect 6631 1087 6633 1099
rect 6631 1072 6635 1087
rect 6621 1068 6635 1072
rect 6621 1064 6625 1068
rect 3431 980 3465 984
rect 3481 980 3485 984
rect 3491 980 3495 984
rect 3563 980 3567 984
rect 3585 980 3589 984
rect 3635 980 3639 984
rect 3655 980 3659 984
rect 3669 980 3673 984
rect 3689 980 3693 984
rect 3701 980 3705 984
rect 3721 980 3725 984
rect 3767 980 3771 984
rect 3775 980 3779 984
rect 3795 980 3799 984
rect 3803 980 3807 984
rect 3825 980 3829 984
rect 3871 980 3905 984
rect 3921 980 3925 984
rect 3931 980 3935 984
rect 4005 980 4009 984
rect 4015 980 4019 984
rect 4035 980 4069 984
rect 4111 980 4115 984
rect 4171 980 4175 984
rect 4181 980 4185 984
rect 4211 980 4215 984
rect 4221 980 4225 984
rect 4291 980 4295 984
rect 4299 980 4303 984
rect 4390 980 4394 984
rect 4412 980 4416 984
rect 4420 980 4424 984
rect 4485 980 4489 984
rect 4505 980 4509 984
rect 4525 980 4529 984
rect 4575 980 4579 984
rect 4595 980 4599 984
rect 4609 980 4613 984
rect 4629 980 4633 984
rect 4641 980 4645 984
rect 4661 980 4665 984
rect 4707 980 4711 984
rect 4715 980 4719 984
rect 4735 980 4739 984
rect 4743 980 4747 984
rect 4765 980 4769 984
rect 4811 980 4815 984
rect 4821 980 4825 984
rect 4851 980 4855 984
rect 4861 980 4865 984
rect 4957 980 4961 984
rect 4965 980 4969 984
rect 5030 980 5034 984
rect 5052 980 5056 984
rect 5060 980 5064 984
rect 5137 980 5141 984
rect 5145 980 5149 984
rect 5191 980 5195 984
rect 5199 980 5203 984
rect 5271 980 5275 984
rect 5279 980 5283 984
rect 5363 980 5367 984
rect 5385 980 5389 984
rect 5431 980 5435 984
rect 5439 980 5443 984
rect 5511 980 5515 984
rect 5519 980 5523 984
rect 5591 980 5595 984
rect 5611 980 5615 984
rect 5631 980 5635 984
rect 5691 980 5695 984
rect 5701 980 5705 984
rect 5721 980 5725 984
rect 5817 980 5821 984
rect 5825 980 5829 984
rect 5876 980 5880 984
rect 5884 980 5888 984
rect 5906 980 5910 984
rect 5985 980 5989 984
rect 6005 980 6009 984
rect 6025 980 6029 984
rect 6076 980 6080 984
rect 6084 980 6088 984
rect 6106 980 6110 984
rect 6197 980 6201 984
rect 6205 980 6209 984
rect 6251 980 6255 984
rect 6259 980 6263 984
rect 6331 980 6335 984
rect 6353 980 6357 984
rect 6361 980 6365 984
rect 6381 980 6385 984
rect 6389 980 6393 984
rect 6435 980 6439 984
rect 6455 980 6459 984
rect 6467 980 6471 984
rect 6487 980 6491 984
rect 6501 980 6505 984
rect 6521 980 6525 984
rect 6571 980 6575 984
rect 6581 980 6585 984
rect 6611 980 6615 984
rect 6621 980 6625 984
rect 31 956 35 960
rect 41 956 45 960
rect 61 956 65 960
rect 145 956 149 960
rect 165 956 169 960
rect 211 956 215 960
rect 233 956 237 960
rect 241 956 245 960
rect 261 956 265 960
rect 269 956 273 960
rect 315 956 319 960
rect 335 956 339 960
rect 347 956 351 960
rect 367 956 371 960
rect 381 956 385 960
rect 401 956 405 960
rect 465 956 469 960
rect 537 956 541 960
rect 545 956 549 960
rect 591 956 595 960
rect 599 956 603 960
rect 671 956 675 960
rect 691 956 695 960
rect 751 956 755 960
rect 771 956 775 960
rect 791 956 795 960
rect 851 956 855 960
rect 861 956 865 960
rect 891 956 895 960
rect 901 956 905 960
rect 976 956 980 960
rect 984 956 988 960
rect 1006 956 1010 960
rect 1076 956 1080 960
rect 1084 956 1088 960
rect 1106 956 1110 960
rect 1245 956 1249 960
rect 1265 956 1269 960
rect 1285 956 1289 960
rect 1305 956 1309 960
rect 1356 956 1360 960
rect 1364 956 1368 960
rect 1386 956 1390 960
rect 1465 956 1469 960
rect 1515 956 1519 960
rect 1535 956 1539 960
rect 1549 956 1553 960
rect 1569 956 1573 960
rect 1581 956 1585 960
rect 1601 956 1605 960
rect 1647 956 1651 960
rect 1655 956 1659 960
rect 1675 956 1679 960
rect 1683 956 1687 960
rect 1705 956 1709 960
rect 1751 956 1755 960
rect 1811 956 1845 960
rect 1861 956 1865 960
rect 1871 956 1875 960
rect 1936 956 1940 960
rect 1944 956 1948 960
rect 1966 956 1970 960
rect 2031 956 2035 960
rect 2051 956 2055 960
rect 2111 956 2115 960
rect 2133 956 2137 960
rect 2141 956 2145 960
rect 2161 956 2165 960
rect 2169 956 2173 960
rect 2215 956 2219 960
rect 2235 956 2239 960
rect 2247 956 2251 960
rect 2267 956 2271 960
rect 2281 956 2285 960
rect 2301 956 2305 960
rect 2351 956 2355 960
rect 2411 956 2415 960
rect 2421 956 2425 960
rect 2451 956 2455 960
rect 2461 956 2465 960
rect 2531 956 2535 960
rect 2539 956 2543 960
rect 2630 956 2634 960
rect 2652 956 2656 960
rect 2660 956 2664 960
rect 2725 956 2729 960
rect 2745 956 2749 960
rect 2765 956 2769 960
rect 2785 956 2789 960
rect 2805 956 2809 960
rect 2825 956 2829 960
rect 2845 956 2849 960
rect 2865 956 2869 960
rect 2911 956 2915 960
rect 2931 956 2935 960
rect 2951 956 2955 960
rect 3025 956 3029 960
rect 3045 956 3049 960
rect 3065 956 3069 960
rect 3125 956 3129 960
rect 3135 956 3139 960
rect 3155 956 3189 960
rect 3245 956 3249 960
rect 3255 956 3259 960
rect 3275 956 3309 960
rect 3370 956 3374 960
rect 3392 956 3396 960
rect 3400 956 3404 960
rect 3451 956 3455 960
rect 3471 956 3475 960
rect 3531 956 3565 960
rect 3581 956 3585 960
rect 3591 956 3595 960
rect 3665 956 3669 960
rect 3725 956 3729 960
rect 3735 956 3739 960
rect 3755 956 3789 960
rect 3835 956 3839 960
rect 3855 956 3859 960
rect 3869 956 3873 960
rect 3889 956 3893 960
rect 3901 956 3905 960
rect 3921 956 3925 960
rect 3967 956 3971 960
rect 3975 956 3979 960
rect 3995 956 3999 960
rect 4003 956 4007 960
rect 4025 956 4029 960
rect 4071 956 4105 960
rect 4121 956 4125 960
rect 4131 956 4135 960
rect 4191 956 4195 960
rect 4211 956 4215 960
rect 4231 956 4235 960
rect 4296 956 4300 960
rect 4304 956 4308 960
rect 4326 956 4330 960
rect 4405 956 4409 960
rect 4425 956 4429 960
rect 4445 956 4449 960
rect 4491 956 4495 960
rect 4556 956 4560 960
rect 4564 956 4568 960
rect 4586 956 4590 960
rect 4651 956 4655 960
rect 4671 956 4675 960
rect 4745 956 4749 960
rect 4796 956 4800 960
rect 4804 956 4808 960
rect 4826 956 4830 960
rect 4891 956 4895 960
rect 4911 956 4915 960
rect 4971 956 5005 960
rect 5021 956 5025 960
rect 5031 956 5035 960
rect 5105 956 5109 960
rect 5115 956 5119 960
rect 5135 956 5169 960
rect 5211 956 5215 960
rect 5231 956 5235 960
rect 5251 956 5255 960
rect 5271 956 5275 960
rect 5291 956 5295 960
rect 5311 956 5315 960
rect 5331 956 5335 960
rect 5351 956 5355 960
rect 5411 956 5415 960
rect 5431 956 5435 960
rect 5451 956 5455 960
rect 5525 956 5529 960
rect 5576 956 5580 960
rect 5584 956 5588 960
rect 5606 956 5610 960
rect 5671 956 5675 960
rect 5691 956 5695 960
rect 5756 956 5760 960
rect 5764 956 5768 960
rect 5786 956 5790 960
rect 5865 956 5869 960
rect 5885 956 5889 960
rect 5905 956 5909 960
rect 5955 956 5959 960
rect 5975 956 5979 960
rect 5989 956 5993 960
rect 6009 956 6013 960
rect 6021 956 6025 960
rect 6041 956 6045 960
rect 6087 956 6091 960
rect 6095 956 6099 960
rect 6115 956 6119 960
rect 6123 956 6127 960
rect 6145 956 6149 960
rect 6196 956 6200 960
rect 6204 956 6208 960
rect 6226 956 6230 960
rect 6296 956 6300 960
rect 6304 956 6308 960
rect 6326 956 6330 960
rect 6405 956 6409 960
rect 6425 956 6429 960
rect 6475 956 6479 960
rect 6495 956 6499 960
rect 6509 956 6513 960
rect 6529 956 6533 960
rect 6541 956 6545 960
rect 6561 956 6565 960
rect 6607 956 6611 960
rect 6615 956 6619 960
rect 6635 956 6639 960
rect 6643 956 6647 960
rect 6665 956 6669 960
rect 31 872 35 876
rect 22 867 35 872
rect 22 833 26 867
rect 41 853 45 876
rect 61 871 65 876
rect 22 776 26 821
rect 41 777 45 841
rect 145 839 149 916
rect 146 827 149 839
rect 143 811 149 827
rect 165 839 169 916
rect 233 913 237 936
rect 229 906 237 913
rect 229 877 233 906
rect 241 896 245 936
rect 261 884 265 916
rect 269 912 273 916
rect 269 910 305 912
rect 269 908 293 910
rect 211 864 215 876
rect 229 871 237 877
rect 211 852 213 864
rect 165 827 174 839
rect 165 811 171 827
rect 143 804 157 811
rect 65 792 75 804
rect 71 784 75 792
rect 153 784 157 804
rect 163 804 171 811
rect 163 784 167 804
rect 211 784 215 852
rect 233 825 237 871
rect 22 771 35 776
rect 41 771 55 777
rect 31 764 35 771
rect 51 764 55 771
rect 233 764 237 813
rect 261 789 267 884
rect 243 785 267 789
rect 243 764 247 785
rect 263 780 281 781
rect 263 776 293 780
rect 263 764 267 776
rect 301 772 305 898
rect 315 890 319 916
rect 335 910 339 916
rect 271 768 305 772
rect 271 764 275 768
rect 317 764 321 878
rect 333 788 337 898
rect 347 876 351 916
rect 342 864 345 876
rect 342 800 346 864
rect 367 857 371 916
rect 362 849 371 857
rect 362 820 366 849
rect 381 834 385 916
rect 401 833 405 876
rect 465 833 469 916
rect 537 853 541 876
rect 526 841 541 853
rect 545 853 549 876
rect 591 853 595 876
rect 545 841 554 853
rect 586 841 595 853
rect 599 853 603 876
rect 599 841 614 853
rect 342 796 375 800
rect 341 776 343 788
rect 339 764 343 776
rect 349 776 351 788
rect 349 764 353 776
rect 371 764 375 796
rect 381 764 385 822
rect 465 821 474 833
rect 401 784 405 821
rect 465 764 469 821
rect 525 764 529 841
rect 545 764 549 841
rect 591 764 595 841
rect 611 764 615 841
rect 671 839 675 916
rect 666 827 675 839
rect 669 811 675 827
rect 691 839 695 916
rect 751 908 755 916
rect 740 904 755 908
rect 771 904 775 916
rect 740 873 746 904
rect 760 900 775 904
rect 760 893 766 900
rect 746 861 756 873
rect 691 827 694 839
rect 691 811 697 827
rect 669 804 677 811
rect 673 784 677 804
rect 683 804 697 811
rect 752 804 756 861
rect 760 804 764 881
rect 791 873 795 916
rect 768 861 775 873
rect 787 861 795 873
rect 851 872 855 876
rect 841 868 855 872
rect 861 872 865 876
rect 861 868 875 872
rect 768 804 772 861
rect 841 853 846 868
rect 683 784 687 804
rect 840 795 846 841
rect 869 819 875 868
rect 891 819 895 876
rect 901 872 905 876
rect 976 872 980 876
rect 901 868 915 872
rect 911 853 915 868
rect 962 864 980 872
rect 962 853 966 864
rect 911 841 913 853
rect 866 807 875 819
rect 840 791 855 795
rect 851 784 855 791
rect 871 784 875 807
rect 891 784 895 807
rect 911 784 915 841
rect 962 796 966 841
rect 984 819 988 876
rect 1006 873 1010 916
rect 1181 948 1185 952
rect 1201 948 1205 952
rect 1006 861 1013 873
rect 1076 872 1080 876
rect 1062 864 1080 872
rect 986 807 995 819
rect 962 789 975 796
rect 971 784 975 789
rect 991 784 995 807
rect 1011 784 1015 861
rect 1062 853 1066 864
rect 1062 796 1066 841
rect 1084 819 1088 876
rect 1106 873 1110 916
rect 1245 892 1249 896
rect 1265 892 1269 896
rect 1245 888 1269 892
rect 1181 880 1185 888
rect 1201 880 1205 888
rect 1181 876 1231 880
rect 1106 861 1113 873
rect 1086 807 1095 819
rect 1062 789 1075 796
rect 1071 784 1075 789
rect 1091 784 1095 807
rect 1111 784 1115 861
rect 1225 853 1231 876
rect 1225 841 1234 853
rect 1225 786 1231 841
rect 1265 819 1269 888
rect 1266 807 1269 819
rect 1225 780 1249 786
rect 1245 764 1249 780
rect 1265 764 1269 807
rect 1285 892 1289 896
rect 1305 892 1309 896
rect 1285 888 1309 892
rect 1285 853 1289 888
rect 1356 872 1360 876
rect 1342 864 1360 872
rect 1342 853 1346 864
rect 1285 841 1294 853
rect 1285 764 1289 841
rect 1342 796 1346 841
rect 1364 819 1368 876
rect 1386 873 1390 916
rect 1386 861 1393 873
rect 1366 807 1375 819
rect 1342 789 1355 796
rect 1351 784 1355 789
rect 1371 784 1375 807
rect 1391 784 1395 861
rect 1465 833 1469 916
rect 1515 833 1519 876
rect 1535 834 1539 916
rect 1549 857 1553 916
rect 1569 876 1573 916
rect 1581 910 1585 916
rect 1575 864 1578 876
rect 1549 849 1558 857
rect 1465 821 1474 833
rect 1465 764 1469 821
rect 1515 784 1519 821
rect 1535 764 1539 822
rect 1554 820 1558 849
rect 1574 800 1578 864
rect 1545 796 1578 800
rect 1545 764 1549 796
rect 1583 788 1587 898
rect 1601 890 1605 916
rect 1647 912 1651 916
rect 1615 910 1651 912
rect 1627 908 1651 910
rect 1569 776 1571 788
rect 1567 764 1571 776
rect 1577 776 1579 788
rect 1577 764 1581 776
rect 1599 764 1603 878
rect 1615 772 1619 898
rect 1655 884 1659 916
rect 1675 896 1679 936
rect 1683 913 1687 936
rect 1683 906 1691 913
rect 1653 789 1659 884
rect 1687 877 1691 906
rect 1683 871 1691 877
rect 1811 948 1815 956
rect 1831 948 1835 952
rect 1841 948 1845 956
rect 1683 825 1687 871
rect 1705 864 1709 876
rect 1707 852 1709 864
rect 1653 785 1677 789
rect 1639 780 1657 781
rect 1627 776 1657 780
rect 1615 768 1649 772
rect 1645 764 1649 768
rect 1653 764 1657 776
rect 1673 764 1677 785
rect 1683 764 1687 813
rect 1705 784 1709 852
rect 1751 833 1755 916
rect 1811 904 1815 908
rect 1746 821 1755 833
rect 1751 764 1755 821
rect 1803 900 1815 904
rect 1803 819 1807 900
rect 1831 863 1835 868
rect 1841 864 1845 868
rect 1822 859 1835 863
rect 1822 853 1827 859
rect 1861 854 1865 876
rect 1835 850 1865 854
rect 1871 853 1875 876
rect 1936 872 1940 876
rect 1922 864 1940 872
rect 1922 853 1926 864
rect 1803 781 1807 807
rect 1821 810 1826 841
rect 1871 841 1874 853
rect 1821 804 1835 810
rect 1831 792 1835 804
rect 1841 792 1845 838
rect 1861 792 1865 796
rect 1871 792 1875 841
rect 1922 796 1926 841
rect 1944 819 1948 876
rect 1966 873 1970 916
rect 1966 861 1973 873
rect 1946 807 1955 819
rect 1803 776 1815 781
rect 1811 772 1815 776
rect 1922 789 1935 796
rect 1931 784 1935 789
rect 1951 784 1955 807
rect 1971 784 1975 861
rect 2031 839 2035 916
rect 2026 827 2035 839
rect 2029 811 2035 827
rect 2051 839 2055 916
rect 2133 913 2137 936
rect 2129 906 2137 913
rect 2129 877 2133 906
rect 2141 896 2145 936
rect 2161 884 2165 916
rect 2169 912 2173 916
rect 2169 910 2205 912
rect 2169 908 2193 910
rect 2111 864 2115 876
rect 2129 871 2137 877
rect 2111 852 2113 864
rect 2051 827 2054 839
rect 2051 811 2057 827
rect 2029 804 2037 811
rect 2033 784 2037 804
rect 2043 804 2057 811
rect 2043 784 2047 804
rect 2111 784 2115 852
rect 2133 825 2137 871
rect 1811 744 1815 752
rect 1831 748 1835 752
rect 1841 748 1845 752
rect 1861 744 1865 752
rect 1871 748 1875 752
rect 2133 764 2137 813
rect 2161 789 2167 884
rect 2143 785 2167 789
rect 2143 764 2147 785
rect 2163 780 2181 781
rect 2163 776 2193 780
rect 2163 764 2167 776
rect 2201 772 2205 898
rect 2215 890 2219 916
rect 2235 910 2239 916
rect 2171 768 2205 772
rect 2171 764 2175 768
rect 2217 764 2221 878
rect 2233 788 2237 898
rect 2247 876 2251 916
rect 2242 864 2245 876
rect 2242 800 2246 864
rect 2267 857 2271 916
rect 2262 849 2271 857
rect 2262 820 2266 849
rect 2281 834 2285 916
rect 2301 833 2305 876
rect 2351 833 2355 916
rect 2411 872 2415 876
rect 2401 868 2415 872
rect 2421 872 2425 876
rect 2421 868 2435 872
rect 2401 853 2406 868
rect 2242 796 2275 800
rect 2241 776 2243 788
rect 2239 764 2243 776
rect 2249 776 2251 788
rect 2249 764 2253 776
rect 2271 764 2275 796
rect 2281 764 2285 822
rect 2346 821 2355 833
rect 2301 784 2305 821
rect 2351 764 2355 821
rect 2400 795 2406 841
rect 2429 819 2435 868
rect 2451 819 2455 876
rect 2461 872 2465 876
rect 2461 868 2475 872
rect 2471 853 2475 868
rect 2531 853 2535 876
rect 2471 841 2473 853
rect 2526 841 2535 853
rect 2539 853 2543 876
rect 2630 873 2634 916
rect 3155 948 3159 956
rect 3165 948 3169 952
rect 3185 948 3189 956
rect 2627 861 2634 873
rect 2539 841 2554 853
rect 2426 807 2435 819
rect 2400 791 2415 795
rect 2411 784 2415 791
rect 2431 784 2435 807
rect 2451 784 2455 807
rect 2471 784 2475 841
rect 2531 764 2535 841
rect 2551 764 2555 841
rect 2625 784 2629 861
rect 2652 819 2656 876
rect 2660 872 2664 876
rect 2660 864 2678 872
rect 2674 853 2678 864
rect 2645 807 2654 819
rect 2645 784 2649 807
rect 2674 796 2678 841
rect 2665 789 2678 796
rect 2725 816 2729 876
rect 2745 816 2749 876
rect 2765 816 2769 876
rect 2785 816 2789 876
rect 2805 816 2809 876
rect 2825 816 2829 876
rect 2845 819 2849 876
rect 2865 819 2869 876
rect 2911 862 2915 876
rect 2931 862 2935 876
rect 2899 856 2915 862
rect 2920 856 2935 862
rect 2899 819 2906 856
rect 2920 833 2926 856
rect 2725 804 2738 816
rect 2765 804 2778 816
rect 2805 804 2818 816
rect 2845 807 2854 819
rect 2866 807 2869 819
rect 2665 784 2669 789
rect 2725 784 2729 804
rect 2745 784 2749 804
rect 2765 784 2769 804
rect 2785 784 2789 804
rect 2805 784 2809 804
rect 2825 784 2829 804
rect 2845 784 2849 807
rect 2865 784 2869 807
rect 2899 794 2906 807
rect 2899 788 2918 794
rect 2914 784 2918 788
rect 2922 784 2926 821
rect 2951 819 2955 876
rect 2946 807 2955 819
rect 3025 819 3029 876
rect 3045 862 3049 876
rect 3065 862 3069 876
rect 3045 856 3060 862
rect 3065 856 3081 862
rect 3054 833 3060 856
rect 3025 807 3034 819
rect 2944 764 2948 807
rect 3032 764 3036 807
rect 3054 784 3058 821
rect 3074 819 3081 856
rect 3125 853 3129 876
rect 3126 841 3129 853
rect 3135 854 3139 876
rect 3185 904 3189 908
rect 3185 900 3197 904
rect 3155 864 3159 868
rect 3165 863 3169 868
rect 3165 859 3178 863
rect 3135 850 3165 854
rect 3074 794 3081 807
rect 3062 788 3081 794
rect 3125 792 3129 841
rect 3173 853 3178 859
rect 3135 792 3139 796
rect 3155 792 3159 838
rect 3174 810 3179 841
rect 3165 804 3179 810
rect 3193 819 3197 900
rect 3275 948 3279 956
rect 3285 948 3289 952
rect 3305 948 3309 956
rect 3245 853 3249 876
rect 3246 841 3249 853
rect 3255 854 3259 876
rect 3305 904 3309 908
rect 3305 900 3317 904
rect 3275 864 3279 868
rect 3285 863 3289 868
rect 3285 859 3298 863
rect 3255 850 3285 854
rect 3165 792 3169 804
rect 3062 784 3066 788
rect 3193 781 3197 807
rect 3245 792 3249 841
rect 3293 853 3298 859
rect 3255 792 3259 796
rect 3275 792 3279 838
rect 3294 810 3299 841
rect 3285 804 3299 810
rect 3313 819 3317 900
rect 3370 873 3374 916
rect 3531 948 3535 956
rect 3551 948 3555 952
rect 3561 948 3565 956
rect 3367 861 3374 873
rect 3285 792 3289 804
rect 3185 776 3197 781
rect 3185 772 3189 776
rect 3313 781 3317 807
rect 3365 784 3369 861
rect 3392 819 3396 876
rect 3400 872 3404 876
rect 3400 864 3418 872
rect 3414 853 3418 864
rect 3385 807 3394 819
rect 3385 784 3389 807
rect 3414 796 3418 841
rect 3451 839 3455 916
rect 3446 827 3455 839
rect 3449 811 3455 827
rect 3471 839 3475 916
rect 3531 904 3535 908
rect 3523 900 3535 904
rect 3471 827 3474 839
rect 3471 811 3477 827
rect 3523 819 3527 900
rect 3551 863 3555 868
rect 3561 864 3565 868
rect 3542 859 3555 863
rect 3542 853 3547 859
rect 3581 854 3585 876
rect 3555 850 3585 854
rect 3591 853 3595 876
rect 3449 804 3457 811
rect 3405 789 3418 796
rect 3405 784 3409 789
rect 3453 784 3457 804
rect 3463 804 3477 811
rect 3463 784 3467 804
rect 3305 776 3317 781
rect 3305 772 3309 776
rect 3125 748 3129 752
rect 3135 744 3139 752
rect 3155 748 3159 752
rect 3165 748 3169 752
rect 3185 744 3189 752
rect 3245 748 3249 752
rect 31 740 35 744
rect 51 740 55 744
rect 71 740 75 744
rect 153 740 157 744
rect 163 740 167 744
rect 211 740 215 744
rect 233 740 237 744
rect 243 740 247 744
rect 263 740 267 744
rect 271 740 275 744
rect 317 740 321 744
rect 339 740 343 744
rect 349 740 353 744
rect 371 740 375 744
rect 381 740 385 744
rect 401 740 405 744
rect 465 740 469 744
rect 525 740 529 744
rect 545 740 549 744
rect 591 740 595 744
rect 611 740 615 744
rect 673 740 677 744
rect 683 740 687 744
rect 752 740 756 744
rect 760 740 764 744
rect 768 740 772 744
rect 851 740 855 744
rect 871 740 875 744
rect 891 740 895 744
rect 911 740 915 744
rect 971 740 975 744
rect 991 740 995 744
rect 1011 740 1015 744
rect 1071 740 1075 744
rect 1091 740 1095 744
rect 1111 740 1115 744
rect 1245 740 1249 744
rect 1265 740 1269 744
rect 1285 740 1289 744
rect 1351 740 1355 744
rect 1371 740 1375 744
rect 1391 740 1395 744
rect 1465 740 1469 744
rect 1515 740 1519 744
rect 1535 740 1539 744
rect 1545 740 1549 744
rect 1567 740 1571 744
rect 1577 740 1581 744
rect 1599 740 1603 744
rect 1645 740 1649 744
rect 1653 740 1657 744
rect 1673 740 1677 744
rect 1683 740 1687 744
rect 1705 740 1709 744
rect 1751 740 1755 744
rect 1811 740 1865 744
rect 1931 740 1935 744
rect 1951 740 1955 744
rect 1971 740 1975 744
rect 2033 740 2037 744
rect 2043 740 2047 744
rect 2111 740 2115 744
rect 2133 740 2137 744
rect 2143 740 2147 744
rect 2163 740 2167 744
rect 2171 740 2175 744
rect 2217 740 2221 744
rect 2239 740 2243 744
rect 2249 740 2253 744
rect 2271 740 2275 744
rect 2281 740 2285 744
rect 2301 740 2305 744
rect 2351 740 2355 744
rect 2411 740 2415 744
rect 2431 740 2435 744
rect 2451 740 2455 744
rect 2471 740 2475 744
rect 2531 740 2535 744
rect 2551 740 2555 744
rect 2625 740 2629 744
rect 2645 740 2649 744
rect 2665 740 2669 744
rect 2725 740 2729 744
rect 2745 740 2749 744
rect 2765 740 2769 744
rect 2785 740 2789 744
rect 2805 740 2809 744
rect 2825 740 2829 744
rect 2845 740 2849 744
rect 2865 740 2869 744
rect 2914 740 2918 744
rect 2922 740 2926 744
rect 2944 740 2948 744
rect 3032 740 3036 744
rect 3054 740 3058 744
rect 3062 740 3066 744
rect 3135 740 3189 744
rect 3255 744 3259 752
rect 3275 748 3279 752
rect 3285 748 3289 752
rect 3305 744 3309 752
rect 3523 781 3527 807
rect 3541 810 3546 841
rect 3591 841 3594 853
rect 3541 804 3555 810
rect 3551 792 3555 804
rect 3561 792 3565 838
rect 3581 792 3585 796
rect 3591 792 3595 841
rect 3665 833 3669 916
rect 3755 948 3759 956
rect 3765 948 3769 952
rect 3785 948 3789 956
rect 3725 853 3729 876
rect 3726 841 3729 853
rect 3735 854 3739 876
rect 3785 904 3789 908
rect 3785 900 3797 904
rect 3755 864 3759 868
rect 3765 863 3769 868
rect 3765 859 3778 863
rect 3735 850 3765 854
rect 3665 821 3674 833
rect 3523 776 3535 781
rect 3531 772 3535 776
rect 3665 764 3669 821
rect 3725 792 3729 841
rect 3773 853 3778 859
rect 3735 792 3739 796
rect 3755 792 3759 838
rect 3774 810 3779 841
rect 3765 804 3779 810
rect 3793 819 3797 900
rect 3835 833 3839 876
rect 3855 834 3859 916
rect 3869 857 3873 916
rect 3889 876 3893 916
rect 3901 910 3905 916
rect 3895 864 3898 876
rect 3869 849 3878 857
rect 3765 792 3769 804
rect 3531 744 3535 752
rect 3551 748 3555 752
rect 3561 748 3565 752
rect 3581 744 3585 752
rect 3591 748 3595 752
rect 3793 781 3797 807
rect 3835 784 3839 821
rect 3785 776 3797 781
rect 3785 772 3789 776
rect 3725 748 3729 752
rect 3735 744 3739 752
rect 3755 748 3759 752
rect 3765 748 3769 752
rect 3785 744 3789 752
rect 3855 764 3859 822
rect 3874 820 3878 849
rect 3894 800 3898 864
rect 3865 796 3898 800
rect 3865 764 3869 796
rect 3903 788 3907 898
rect 3921 890 3925 916
rect 3967 912 3971 916
rect 3935 910 3971 912
rect 3947 908 3971 910
rect 3889 776 3891 788
rect 3887 764 3891 776
rect 3897 776 3899 788
rect 3897 764 3901 776
rect 3919 764 3923 878
rect 3935 772 3939 898
rect 3975 884 3979 916
rect 3995 896 3999 936
rect 4003 913 4007 936
rect 4003 906 4011 913
rect 3973 789 3979 884
rect 4007 877 4011 906
rect 4003 871 4011 877
rect 4071 948 4075 956
rect 4091 948 4095 952
rect 4101 948 4105 956
rect 4071 904 4075 908
rect 4063 900 4075 904
rect 4003 825 4007 871
rect 4025 864 4029 876
rect 4027 852 4029 864
rect 3973 785 3997 789
rect 3959 780 3977 781
rect 3947 776 3977 780
rect 3935 768 3969 772
rect 3965 764 3969 768
rect 3973 764 3977 776
rect 3993 764 3997 785
rect 4003 764 4007 813
rect 4025 784 4029 852
rect 4063 819 4067 900
rect 4091 863 4095 868
rect 4101 864 4105 868
rect 4082 859 4095 863
rect 4082 853 4087 859
rect 4121 854 4125 876
rect 4095 850 4125 854
rect 4131 853 4135 876
rect 4191 862 4195 876
rect 4211 862 4215 876
rect 4179 856 4195 862
rect 4200 856 4215 862
rect 4063 781 4067 807
rect 4081 810 4086 841
rect 4131 841 4134 853
rect 4081 804 4095 810
rect 4091 792 4095 804
rect 4101 792 4105 838
rect 4121 792 4125 796
rect 4131 792 4135 841
rect 4179 819 4186 856
rect 4200 833 4206 856
rect 4179 794 4186 807
rect 4063 776 4075 781
rect 4071 772 4075 776
rect 4179 788 4198 794
rect 4194 784 4198 788
rect 4202 784 4206 821
rect 4231 819 4235 876
rect 4296 872 4300 876
rect 4282 864 4300 872
rect 4282 853 4286 864
rect 4226 807 4235 819
rect 4071 744 4075 752
rect 4091 748 4095 752
rect 4101 748 4105 752
rect 4121 744 4125 752
rect 4131 748 4135 752
rect 4224 764 4228 807
rect 4282 796 4286 841
rect 4304 819 4308 876
rect 4326 873 4330 916
rect 4405 873 4409 916
rect 4425 904 4429 916
rect 4445 908 4449 916
rect 4445 904 4460 908
rect 4425 900 4440 904
rect 4434 893 4440 900
rect 4326 861 4333 873
rect 4405 861 4413 873
rect 4425 861 4432 873
rect 4306 807 4315 819
rect 4282 789 4295 796
rect 4291 784 4295 789
rect 4311 784 4315 807
rect 4331 784 4335 861
rect 4428 804 4432 861
rect 4436 804 4440 881
rect 4454 873 4460 904
rect 4444 861 4454 873
rect 4444 804 4448 861
rect 4491 833 4495 916
rect 4556 872 4560 876
rect 4542 864 4560 872
rect 4542 853 4546 864
rect 4486 821 4495 833
rect 4491 764 4495 821
rect 4542 796 4546 841
rect 4564 819 4568 876
rect 4586 873 4590 916
rect 4586 861 4593 873
rect 4566 807 4575 819
rect 4542 789 4555 796
rect 4551 784 4555 789
rect 4571 784 4575 807
rect 4591 784 4595 861
rect 4651 839 4655 916
rect 4646 827 4655 839
rect 4649 811 4655 827
rect 4671 839 4675 916
rect 4671 827 4674 839
rect 4745 833 4749 916
rect 4971 948 4975 956
rect 4991 948 4995 952
rect 5001 948 5005 956
rect 4796 872 4800 876
rect 4782 864 4800 872
rect 4782 853 4786 864
rect 4671 811 4677 827
rect 4649 804 4657 811
rect 4653 784 4657 804
rect 4663 804 4677 811
rect 4745 821 4754 833
rect 4663 784 4667 804
rect 4745 764 4749 821
rect 4782 796 4786 841
rect 4804 819 4808 876
rect 4826 873 4830 916
rect 4826 861 4833 873
rect 4806 807 4815 819
rect 4782 789 4795 796
rect 4791 784 4795 789
rect 4811 784 4815 807
rect 4831 784 4835 861
rect 4891 839 4895 916
rect 4886 827 4895 839
rect 4889 811 4895 827
rect 4911 839 4915 916
rect 4971 904 4975 908
rect 4963 900 4975 904
rect 4911 827 4914 839
rect 4911 811 4917 827
rect 4963 819 4967 900
rect 5135 948 5139 956
rect 5145 948 5149 952
rect 5165 948 5169 956
rect 4991 863 4995 868
rect 5001 864 5005 868
rect 4982 859 4995 863
rect 4982 853 4987 859
rect 5021 854 5025 876
rect 4995 850 5025 854
rect 5031 853 5035 876
rect 5105 853 5109 876
rect 4889 804 4897 811
rect 4893 784 4897 804
rect 4903 804 4917 811
rect 4903 784 4907 804
rect 4963 781 4967 807
rect 4981 810 4986 841
rect 5031 841 5034 853
rect 5106 841 5109 853
rect 5115 854 5119 876
rect 5165 904 5169 908
rect 5165 900 5177 904
rect 5135 864 5139 868
rect 5145 863 5149 868
rect 5145 859 5158 863
rect 5115 850 5145 854
rect 4981 804 4995 810
rect 4991 792 4995 804
rect 5001 792 5005 838
rect 5021 792 5025 796
rect 5031 792 5035 841
rect 5105 792 5109 841
rect 5153 853 5158 859
rect 5115 792 5119 796
rect 5135 792 5139 838
rect 5154 810 5159 841
rect 5145 804 5159 810
rect 5173 819 5177 900
rect 5211 819 5215 876
rect 5231 819 5235 876
rect 5211 807 5214 819
rect 5226 807 5235 819
rect 5251 816 5255 876
rect 5271 816 5275 876
rect 5291 816 5295 876
rect 5311 816 5315 876
rect 5331 816 5335 876
rect 5351 816 5355 876
rect 5411 862 5415 876
rect 5431 862 5435 876
rect 5399 856 5415 862
rect 5420 856 5435 862
rect 5399 819 5406 856
rect 5420 833 5426 856
rect 5145 792 5149 804
rect 4963 776 4975 781
rect 4971 772 4975 776
rect 5173 781 5177 807
rect 5211 784 5215 807
rect 5231 784 5235 807
rect 5262 804 5275 816
rect 5302 804 5315 816
rect 5342 804 5355 816
rect 5251 784 5255 804
rect 5271 784 5275 804
rect 5291 784 5295 804
rect 5311 784 5315 804
rect 5331 784 5335 804
rect 5351 784 5355 804
rect 5399 794 5406 807
rect 5399 788 5418 794
rect 5414 784 5418 788
rect 5422 784 5426 821
rect 5451 819 5455 876
rect 5446 807 5455 819
rect 5525 833 5529 916
rect 5576 872 5580 876
rect 5562 864 5580 872
rect 5562 853 5566 864
rect 5525 821 5534 833
rect 5165 776 5177 781
rect 5165 772 5169 776
rect 4971 744 4975 752
rect 4991 748 4995 752
rect 5001 748 5005 752
rect 5021 744 5025 752
rect 5031 748 5035 752
rect 5105 748 5109 752
rect 3255 740 3309 744
rect 3365 740 3369 744
rect 3385 740 3389 744
rect 3405 740 3409 744
rect 3453 740 3457 744
rect 3463 740 3467 744
rect 3531 740 3585 744
rect 3665 740 3669 744
rect 3735 740 3789 744
rect 3835 740 3839 744
rect 3855 740 3859 744
rect 3865 740 3869 744
rect 3887 740 3891 744
rect 3897 740 3901 744
rect 3919 740 3923 744
rect 3965 740 3969 744
rect 3973 740 3977 744
rect 3993 740 3997 744
rect 4003 740 4007 744
rect 4025 740 4029 744
rect 4071 740 4125 744
rect 4194 740 4198 744
rect 4202 740 4206 744
rect 4224 740 4228 744
rect 4291 740 4295 744
rect 4311 740 4315 744
rect 4331 740 4335 744
rect 4428 740 4432 744
rect 4436 740 4440 744
rect 4444 740 4448 744
rect 4491 740 4495 744
rect 4551 740 4555 744
rect 4571 740 4575 744
rect 4591 740 4595 744
rect 4653 740 4657 744
rect 4663 740 4667 744
rect 4745 740 4749 744
rect 4791 740 4795 744
rect 4811 740 4815 744
rect 4831 740 4835 744
rect 4893 740 4897 744
rect 4903 740 4907 744
rect 4971 740 5025 744
rect 5115 744 5119 752
rect 5135 748 5139 752
rect 5145 748 5149 752
rect 5165 744 5169 752
rect 5444 764 5448 807
rect 5525 764 5529 821
rect 5562 796 5566 841
rect 5584 819 5588 876
rect 5606 873 5610 916
rect 5606 861 5613 873
rect 5586 807 5595 819
rect 5562 789 5575 796
rect 5571 784 5575 789
rect 5591 784 5595 807
rect 5611 784 5615 861
rect 5671 839 5675 916
rect 5666 827 5675 839
rect 5669 811 5675 827
rect 5691 839 5695 916
rect 5756 872 5760 876
rect 5742 864 5760 872
rect 5742 853 5746 864
rect 5691 827 5694 839
rect 5691 811 5697 827
rect 5669 804 5677 811
rect 5673 784 5677 804
rect 5683 804 5697 811
rect 5683 784 5687 804
rect 5742 796 5746 841
rect 5764 819 5768 876
rect 5786 873 5790 916
rect 5865 873 5869 916
rect 5885 904 5889 916
rect 5905 908 5909 916
rect 5905 904 5920 908
rect 5885 900 5900 904
rect 5894 893 5900 900
rect 5786 861 5793 873
rect 5865 861 5873 873
rect 5885 861 5892 873
rect 5766 807 5775 819
rect 5742 789 5755 796
rect 5751 784 5755 789
rect 5771 784 5775 807
rect 5791 784 5795 861
rect 5888 804 5892 861
rect 5896 804 5900 881
rect 5914 873 5920 904
rect 5904 861 5914 873
rect 5904 804 5908 861
rect 5955 833 5959 876
rect 5975 834 5979 916
rect 5989 857 5993 916
rect 6009 876 6013 916
rect 6021 910 6025 916
rect 6015 864 6018 876
rect 5989 849 5998 857
rect 5955 784 5959 821
rect 5975 764 5979 822
rect 5994 820 5998 849
rect 6014 800 6018 864
rect 5985 796 6018 800
rect 5985 764 5989 796
rect 6023 788 6027 898
rect 6041 890 6045 916
rect 6087 912 6091 916
rect 6055 910 6091 912
rect 6067 908 6091 910
rect 6009 776 6011 788
rect 6007 764 6011 776
rect 6017 776 6019 788
rect 6017 764 6021 776
rect 6039 764 6043 878
rect 6055 772 6059 898
rect 6095 884 6099 916
rect 6115 896 6119 936
rect 6123 913 6127 936
rect 6123 906 6131 913
rect 6093 789 6099 884
rect 6127 877 6131 906
rect 6123 871 6131 877
rect 6123 825 6127 871
rect 6145 864 6149 876
rect 6196 872 6200 876
rect 6147 852 6149 864
rect 6182 864 6200 872
rect 6182 853 6186 864
rect 6093 785 6117 789
rect 6079 780 6097 781
rect 6067 776 6097 780
rect 6055 768 6089 772
rect 6085 764 6089 768
rect 6093 764 6097 776
rect 6113 764 6117 785
rect 6123 764 6127 813
rect 6145 784 6149 852
rect 6182 796 6186 841
rect 6204 819 6208 876
rect 6226 873 6230 916
rect 6226 861 6233 873
rect 6296 872 6300 876
rect 6282 864 6300 872
rect 6206 807 6215 819
rect 6182 789 6195 796
rect 6191 784 6195 789
rect 6211 784 6215 807
rect 6231 784 6235 861
rect 6282 853 6286 864
rect 6282 796 6286 841
rect 6304 819 6308 876
rect 6326 873 6330 916
rect 6326 861 6333 873
rect 6306 807 6315 819
rect 6282 789 6295 796
rect 6291 784 6295 789
rect 6311 784 6315 807
rect 6331 784 6335 861
rect 6405 839 6409 916
rect 6406 827 6409 839
rect 6403 811 6409 827
rect 6425 839 6429 916
rect 6425 827 6434 839
rect 6475 833 6479 876
rect 6495 834 6499 916
rect 6509 857 6513 916
rect 6529 876 6533 916
rect 6541 910 6545 916
rect 6535 864 6538 876
rect 6509 849 6518 857
rect 6425 811 6431 827
rect 6403 804 6417 811
rect 6413 784 6417 804
rect 6423 804 6431 811
rect 6423 784 6427 804
rect 6475 784 6479 821
rect 6495 764 6499 822
rect 6514 820 6518 849
rect 6534 800 6538 864
rect 6505 796 6538 800
rect 6505 764 6509 796
rect 6543 788 6547 898
rect 6561 890 6565 916
rect 6607 912 6611 916
rect 6575 910 6611 912
rect 6587 908 6611 910
rect 6529 776 6531 788
rect 6527 764 6531 776
rect 6537 776 6539 788
rect 6537 764 6541 776
rect 6559 764 6563 878
rect 6575 772 6579 898
rect 6615 884 6619 916
rect 6635 896 6639 936
rect 6643 913 6647 936
rect 6643 906 6651 913
rect 6613 789 6619 884
rect 6647 877 6651 906
rect 6643 871 6651 877
rect 6643 825 6647 871
rect 6665 864 6669 876
rect 6667 852 6669 864
rect 6613 785 6637 789
rect 6599 780 6617 781
rect 6587 776 6617 780
rect 6575 768 6609 772
rect 6605 764 6609 768
rect 6613 764 6617 776
rect 6633 764 6637 785
rect 6643 764 6647 813
rect 6665 784 6669 852
rect 5115 740 5169 744
rect 5211 740 5215 744
rect 5231 740 5235 744
rect 5251 740 5255 744
rect 5271 740 5275 744
rect 5291 740 5295 744
rect 5311 740 5315 744
rect 5331 740 5335 744
rect 5351 740 5355 744
rect 5414 740 5418 744
rect 5422 740 5426 744
rect 5444 740 5448 744
rect 5525 740 5529 744
rect 5571 740 5575 744
rect 5591 740 5595 744
rect 5611 740 5615 744
rect 5673 740 5677 744
rect 5683 740 5687 744
rect 5751 740 5755 744
rect 5771 740 5775 744
rect 5791 740 5795 744
rect 5888 740 5892 744
rect 5896 740 5900 744
rect 5904 740 5908 744
rect 5955 740 5959 744
rect 5975 740 5979 744
rect 5985 740 5989 744
rect 6007 740 6011 744
rect 6017 740 6021 744
rect 6039 740 6043 744
rect 6085 740 6089 744
rect 6093 740 6097 744
rect 6113 740 6117 744
rect 6123 740 6127 744
rect 6145 740 6149 744
rect 6191 740 6195 744
rect 6211 740 6215 744
rect 6231 740 6235 744
rect 6291 740 6295 744
rect 6311 740 6315 744
rect 6331 740 6335 744
rect 6413 740 6417 744
rect 6423 740 6427 744
rect 6475 740 6479 744
rect 6495 740 6499 744
rect 6505 740 6509 744
rect 6527 740 6531 744
rect 6537 740 6541 744
rect 6559 740 6563 744
rect 6605 740 6609 744
rect 6613 740 6617 744
rect 6633 740 6637 744
rect 6643 740 6647 744
rect 6665 740 6669 744
rect 31 716 35 720
rect 93 716 97 720
rect 103 716 107 720
rect 174 716 178 720
rect 182 716 186 720
rect 204 716 208 720
rect 271 716 275 720
rect 352 716 356 720
rect 374 716 378 720
rect 382 716 386 720
rect 432 716 436 720
rect 440 716 444 720
rect 448 716 452 720
rect 553 716 557 720
rect 563 716 567 720
rect 648 716 652 720
rect 656 716 660 720
rect 664 716 668 720
rect 711 716 715 720
rect 771 716 775 720
rect 845 716 849 720
rect 865 716 869 720
rect 985 716 989 720
rect 1005 716 1009 720
rect 1025 716 1029 720
rect 1095 716 1099 720
rect 1115 716 1119 720
rect 1125 716 1129 720
rect 1147 716 1151 720
rect 1157 716 1161 720
rect 1179 716 1183 720
rect 1225 716 1229 720
rect 1233 716 1237 720
rect 1253 716 1257 720
rect 1263 716 1267 720
rect 1285 716 1289 720
rect 1331 716 1335 720
rect 1353 716 1357 720
rect 1413 716 1417 720
rect 1423 716 1427 720
rect 1495 716 1499 720
rect 1515 716 1519 720
rect 1525 716 1529 720
rect 1547 716 1551 720
rect 1557 716 1561 720
rect 1579 716 1583 720
rect 1625 716 1629 720
rect 1633 716 1637 720
rect 1653 716 1657 720
rect 1663 716 1667 720
rect 1685 716 1689 720
rect 1735 716 1739 720
rect 1755 716 1759 720
rect 1765 716 1769 720
rect 1787 716 1791 720
rect 1797 716 1801 720
rect 1819 716 1823 720
rect 1865 716 1869 720
rect 1873 716 1877 720
rect 1893 716 1897 720
rect 1903 716 1907 720
rect 1925 716 1929 720
rect 1975 716 1979 720
rect 1995 716 1999 720
rect 2005 716 2009 720
rect 2027 716 2031 720
rect 2037 716 2041 720
rect 2059 716 2063 720
rect 2105 716 2109 720
rect 2113 716 2117 720
rect 2133 716 2137 720
rect 2143 716 2147 720
rect 2165 716 2169 720
rect 2215 716 2219 720
rect 2235 716 2239 720
rect 2245 716 2249 720
rect 2267 716 2271 720
rect 2277 716 2281 720
rect 2299 716 2303 720
rect 2345 716 2349 720
rect 2353 716 2357 720
rect 2373 716 2377 720
rect 2383 716 2387 720
rect 2405 716 2409 720
rect 2451 716 2455 720
rect 2473 716 2477 720
rect 2483 716 2487 720
rect 2503 716 2507 720
rect 2511 716 2515 720
rect 2557 716 2561 720
rect 2579 716 2583 720
rect 2589 716 2593 720
rect 2611 716 2615 720
rect 2621 716 2625 720
rect 2641 716 2645 720
rect 2726 716 2730 720
rect 2734 716 2738 720
rect 2754 716 2758 720
rect 2762 716 2766 720
rect 2825 716 2829 720
rect 2892 716 2896 720
rect 2914 716 2918 720
rect 2922 716 2926 720
rect 2971 716 2975 720
rect 3031 716 3035 720
rect 3051 716 3055 720
rect 3071 716 3075 720
rect 3133 716 3137 720
rect 3143 716 3147 720
rect 3212 716 3216 720
rect 3220 716 3224 720
rect 3228 716 3232 720
rect 3311 716 3315 720
rect 3371 716 3375 720
rect 3391 716 3395 720
rect 3411 716 3415 720
rect 3473 716 3477 720
rect 3483 716 3487 720
rect 3554 716 3558 720
rect 3562 716 3566 720
rect 3584 716 3588 720
rect 3651 716 3655 720
rect 3671 716 3675 720
rect 3731 716 3735 720
rect 3751 716 3755 720
rect 3771 716 3775 720
rect 3868 716 3872 720
rect 3876 716 3880 720
rect 3884 716 3888 720
rect 3931 716 3935 720
rect 3953 716 3957 720
rect 3963 716 3967 720
rect 3983 716 3987 720
rect 3991 716 3995 720
rect 4037 716 4041 720
rect 4059 716 4063 720
rect 4069 716 4073 720
rect 4091 716 4095 720
rect 4101 716 4105 720
rect 4121 716 4125 720
rect 4185 716 4189 720
rect 4205 716 4209 720
rect 4251 716 4255 720
rect 4273 716 4277 720
rect 4283 716 4287 720
rect 4303 716 4307 720
rect 4311 716 4315 720
rect 4357 716 4361 720
rect 4379 716 4383 720
rect 4389 716 4393 720
rect 4411 716 4415 720
rect 4421 716 4425 720
rect 4441 716 4445 720
rect 4491 716 4495 720
rect 4554 716 4558 720
rect 4562 716 4566 720
rect 4582 716 4586 720
rect 4590 716 4594 720
rect 4692 716 4696 720
rect 4714 716 4718 720
rect 4722 716 4726 720
rect 4785 716 4789 720
rect 4805 716 4809 720
rect 4825 716 4829 720
rect 4873 716 4877 720
rect 4883 716 4887 720
rect 4965 716 4969 720
rect 5035 716 5089 720
rect 5132 716 5136 720
rect 5140 716 5144 720
rect 5148 716 5152 720
rect 5231 716 5235 720
rect 5253 716 5257 720
rect 5263 716 5267 720
rect 5283 716 5287 720
rect 5291 716 5295 720
rect 5337 716 5341 720
rect 5359 716 5363 720
rect 5369 716 5373 720
rect 5391 716 5395 720
rect 5401 716 5405 720
rect 5421 716 5425 720
rect 5471 716 5475 720
rect 5531 716 5585 720
rect 5665 716 5669 720
rect 5685 716 5689 720
rect 5745 716 5749 720
rect 5765 716 5769 720
rect 5825 716 5829 720
rect 5845 716 5849 720
rect 5891 716 5895 720
rect 5911 716 5915 720
rect 5985 716 5989 720
rect 6005 716 6009 720
rect 6051 716 6055 720
rect 6071 716 6075 720
rect 6091 716 6095 720
rect 6151 716 6155 720
rect 6171 716 6175 720
rect 6191 716 6195 720
rect 6273 716 6277 720
rect 6283 716 6287 720
rect 6335 716 6339 720
rect 6355 716 6359 720
rect 6365 716 6369 720
rect 6387 716 6391 720
rect 6397 716 6401 720
rect 6419 716 6423 720
rect 6465 716 6469 720
rect 6473 716 6477 720
rect 6493 716 6497 720
rect 6503 716 6507 720
rect 6525 716 6529 720
rect 6571 716 6575 720
rect 6631 716 6635 720
rect 31 639 35 696
rect 93 656 97 676
rect 26 627 35 639
rect 89 649 97 656
rect 103 656 107 676
rect 174 672 178 676
rect 159 666 178 672
rect 103 649 117 656
rect 159 653 166 666
rect 89 633 95 649
rect 31 544 35 627
rect 86 621 95 633
rect 91 544 95 621
rect 111 633 117 649
rect 111 621 114 633
rect 111 544 115 621
rect 159 604 166 641
rect 182 639 186 676
rect 204 653 208 696
rect 206 641 215 653
rect 180 604 186 627
rect 159 598 175 604
rect 180 598 195 604
rect 171 584 175 598
rect 191 584 195 598
rect 211 584 215 641
rect 271 639 275 696
rect 352 653 356 696
rect 266 627 275 639
rect 271 544 275 627
rect 345 641 354 653
rect 345 584 349 641
rect 374 639 378 676
rect 382 672 386 676
rect 382 666 401 672
rect 394 653 401 666
rect 553 656 557 676
rect 374 604 380 627
rect 394 604 401 641
rect 365 598 380 604
rect 385 598 401 604
rect 432 599 436 656
rect 365 584 369 598
rect 385 584 389 598
rect 426 587 436 599
rect 420 556 426 587
rect 440 579 444 656
rect 448 599 452 656
rect 543 649 557 656
rect 563 656 567 676
rect 563 649 571 656
rect 543 633 549 649
rect 546 621 549 633
rect 448 587 455 599
rect 467 587 475 599
rect 440 560 446 567
rect 440 556 455 560
rect 420 552 435 556
rect 431 544 435 552
rect 451 544 455 556
rect 471 544 475 587
rect 545 544 549 621
rect 565 633 571 649
rect 565 621 574 633
rect 565 544 569 621
rect 648 599 652 656
rect 625 587 633 599
rect 645 587 652 599
rect 625 544 629 587
rect 656 579 660 656
rect 664 599 668 656
rect 711 639 715 696
rect 771 639 775 696
rect 706 627 715 639
rect 766 627 775 639
rect 664 587 674 599
rect 654 560 660 567
rect 645 556 660 560
rect 674 556 680 587
rect 645 544 649 556
rect 665 552 680 556
rect 665 544 669 552
rect 711 544 715 627
rect 771 544 775 627
rect 845 619 849 696
rect 865 619 869 696
rect 985 680 989 696
rect 965 674 989 680
rect 965 619 971 674
rect 1005 653 1009 696
rect 1006 641 1009 653
rect 846 607 861 619
rect 857 584 861 607
rect 865 607 874 619
rect 965 607 974 619
rect 865 584 869 607
rect 965 584 971 607
rect 921 580 971 584
rect 921 572 925 580
rect 941 572 945 580
rect 1005 572 1009 641
rect 985 568 1009 572
rect 985 564 989 568
rect 1005 564 1009 568
rect 1025 619 1029 696
rect 1095 639 1099 676
rect 1115 638 1119 696
rect 1125 664 1129 696
rect 1147 684 1151 696
rect 1149 672 1151 684
rect 1157 684 1161 696
rect 1157 672 1159 684
rect 1125 660 1158 664
rect 1025 607 1034 619
rect 1025 572 1029 607
rect 1095 584 1099 627
rect 1025 568 1049 572
rect 1025 564 1029 568
rect 1045 564 1049 568
rect 921 508 925 512
rect 941 508 945 512
rect 1115 544 1119 626
rect 1134 611 1138 640
rect 1129 603 1138 611
rect 1129 544 1133 603
rect 1154 596 1158 660
rect 1155 584 1158 596
rect 1149 544 1153 584
rect 1163 562 1167 672
rect 1179 582 1183 696
rect 1225 692 1229 696
rect 1195 688 1229 692
rect 1161 544 1165 550
rect 1181 544 1185 570
rect 1195 562 1199 688
rect 1233 684 1237 696
rect 1207 680 1237 684
rect 1219 679 1237 680
rect 1253 675 1257 696
rect 1233 671 1257 675
rect 1233 576 1239 671
rect 1263 647 1267 696
rect 1263 589 1267 635
rect 1285 608 1289 676
rect 1331 619 1335 696
rect 1353 670 1357 676
rect 1355 658 1357 670
rect 1413 656 1417 676
rect 1409 649 1417 656
rect 1423 656 1427 676
rect 1423 649 1437 656
rect 1409 633 1415 649
rect 1406 621 1415 633
rect 1287 596 1289 608
rect 1326 607 1335 619
rect 1263 583 1271 589
rect 1285 584 1289 596
rect 1207 550 1231 552
rect 1195 548 1231 550
rect 1227 544 1231 548
rect 1235 544 1239 576
rect 1255 524 1259 564
rect 1267 554 1271 583
rect 1263 547 1271 554
rect 1263 524 1267 547
rect 1331 544 1335 607
rect 1355 590 1357 602
rect 1353 584 1357 590
rect 1411 544 1415 621
rect 1431 633 1437 649
rect 1495 639 1499 676
rect 1431 621 1434 633
rect 1515 638 1519 696
rect 1525 664 1529 696
rect 1547 684 1551 696
rect 1549 672 1551 684
rect 1557 684 1561 696
rect 1557 672 1559 684
rect 1525 660 1558 664
rect 1431 544 1435 621
rect 1495 584 1499 627
rect 1515 544 1519 626
rect 1534 611 1538 640
rect 1529 603 1538 611
rect 1529 544 1533 603
rect 1554 596 1558 660
rect 1555 584 1558 596
rect 1549 544 1553 584
rect 1563 562 1567 672
rect 1579 582 1583 696
rect 1625 692 1629 696
rect 1595 688 1629 692
rect 1561 544 1565 550
rect 1581 544 1585 570
rect 1595 562 1599 688
rect 1633 684 1637 696
rect 1607 680 1637 684
rect 1619 679 1637 680
rect 1653 675 1657 696
rect 1633 671 1657 675
rect 1633 576 1639 671
rect 1663 647 1667 696
rect 1663 589 1667 635
rect 1685 608 1689 676
rect 1735 639 1739 676
rect 1755 638 1759 696
rect 1765 664 1769 696
rect 1787 684 1791 696
rect 1789 672 1791 684
rect 1797 684 1801 696
rect 1797 672 1799 684
rect 1765 660 1798 664
rect 1687 596 1689 608
rect 1663 583 1671 589
rect 1685 584 1689 596
rect 1735 584 1739 627
rect 1607 550 1631 552
rect 1595 548 1631 550
rect 1627 544 1631 548
rect 1635 544 1639 576
rect 1655 524 1659 564
rect 1667 554 1671 583
rect 1663 547 1671 554
rect 1663 524 1667 547
rect 1755 544 1759 626
rect 1774 611 1778 640
rect 1769 603 1778 611
rect 1769 544 1773 603
rect 1794 596 1798 660
rect 1795 584 1798 596
rect 1789 544 1793 584
rect 1803 562 1807 672
rect 1819 582 1823 696
rect 1865 692 1869 696
rect 1835 688 1869 692
rect 1801 544 1805 550
rect 1821 544 1825 570
rect 1835 562 1839 688
rect 1873 684 1877 696
rect 1847 680 1877 684
rect 1859 679 1877 680
rect 1893 675 1897 696
rect 1873 671 1897 675
rect 1873 576 1879 671
rect 1903 647 1907 696
rect 1903 589 1907 635
rect 1925 608 1929 676
rect 1975 639 1979 676
rect 1995 638 1999 696
rect 2005 664 2009 696
rect 2027 684 2031 696
rect 2029 672 2031 684
rect 2037 684 2041 696
rect 2037 672 2039 684
rect 2005 660 2038 664
rect 1927 596 1929 608
rect 1903 583 1911 589
rect 1925 584 1929 596
rect 1975 584 1979 627
rect 1847 550 1871 552
rect 1835 548 1871 550
rect 1867 544 1871 548
rect 1875 544 1879 576
rect 1895 524 1899 564
rect 1907 554 1911 583
rect 1903 547 1911 554
rect 1903 524 1907 547
rect 1995 544 1999 626
rect 2014 611 2018 640
rect 2009 603 2018 611
rect 2009 544 2013 603
rect 2034 596 2038 660
rect 2035 584 2038 596
rect 2029 544 2033 584
rect 2043 562 2047 672
rect 2059 582 2063 696
rect 2105 692 2109 696
rect 2075 688 2109 692
rect 2041 544 2045 550
rect 2061 544 2065 570
rect 2075 562 2079 688
rect 2113 684 2117 696
rect 2087 680 2117 684
rect 2099 679 2117 680
rect 2133 675 2137 696
rect 2113 671 2137 675
rect 2113 576 2119 671
rect 2143 647 2147 696
rect 2143 589 2147 635
rect 2165 608 2169 676
rect 2215 639 2219 676
rect 2235 638 2239 696
rect 2245 664 2249 696
rect 2267 684 2271 696
rect 2269 672 2271 684
rect 2277 684 2281 696
rect 2277 672 2279 684
rect 2245 660 2278 664
rect 2167 596 2169 608
rect 2143 583 2151 589
rect 2165 584 2169 596
rect 2215 584 2219 627
rect 2087 550 2111 552
rect 2075 548 2111 550
rect 2107 544 2111 548
rect 2115 544 2119 576
rect 2135 524 2139 564
rect 2147 554 2151 583
rect 2143 547 2151 554
rect 2143 524 2147 547
rect 2235 544 2239 626
rect 2254 611 2258 640
rect 2249 603 2258 611
rect 2249 544 2253 603
rect 2274 596 2278 660
rect 2275 584 2278 596
rect 2269 544 2273 584
rect 2283 562 2287 672
rect 2299 582 2303 696
rect 2345 692 2349 696
rect 2315 688 2349 692
rect 2281 544 2285 550
rect 2301 544 2305 570
rect 2315 562 2319 688
rect 2353 684 2357 696
rect 2327 680 2357 684
rect 2339 679 2357 680
rect 2373 675 2377 696
rect 2353 671 2377 675
rect 2353 576 2359 671
rect 2383 647 2387 696
rect 2383 589 2387 635
rect 2405 608 2409 676
rect 2407 596 2409 608
rect 2383 583 2391 589
rect 2405 584 2409 596
rect 2451 608 2455 676
rect 2473 647 2477 696
rect 2483 675 2487 696
rect 2503 684 2507 696
rect 2511 692 2515 696
rect 2511 688 2545 692
rect 2503 680 2533 684
rect 2503 679 2521 680
rect 2483 671 2507 675
rect 2451 596 2453 608
rect 2451 584 2455 596
rect 2473 589 2477 635
rect 2327 550 2351 552
rect 2315 548 2351 550
rect 2347 544 2351 548
rect 2355 544 2359 576
rect 2375 524 2379 564
rect 2387 554 2391 583
rect 2383 547 2391 554
rect 2383 524 2387 547
rect 2469 583 2477 589
rect 2469 554 2473 583
rect 2501 576 2507 671
rect 2469 547 2477 554
rect 2473 524 2477 547
rect 2481 524 2485 564
rect 2501 544 2505 576
rect 2541 562 2545 688
rect 2557 582 2561 696
rect 2579 684 2583 696
rect 2581 672 2583 684
rect 2589 684 2593 696
rect 2589 672 2591 684
rect 2509 550 2533 552
rect 2509 548 2545 550
rect 2509 544 2513 548
rect 2555 544 2559 570
rect 2573 562 2577 672
rect 2611 664 2615 696
rect 2582 660 2615 664
rect 2582 596 2586 660
rect 2602 611 2606 640
rect 2621 638 2625 696
rect 2641 639 2645 676
rect 2726 671 2730 676
rect 2700 667 2730 671
rect 2602 603 2611 611
rect 2582 584 2585 596
rect 2575 544 2579 550
rect 2587 544 2591 584
rect 2607 544 2611 603
rect 2621 544 2625 626
rect 2641 584 2645 627
rect 2700 619 2706 667
rect 2734 662 2738 676
rect 2725 655 2738 662
rect 2725 653 2729 655
rect 2754 653 2758 676
rect 2762 668 2766 676
rect 2762 661 2779 668
rect 2727 641 2729 653
rect 2706 607 2709 619
rect 2705 584 2709 607
rect 2725 584 2729 641
rect 2754 612 2758 641
rect 2773 619 2779 661
rect 2825 639 2829 696
rect 2892 653 2896 696
rect 2885 641 2894 653
rect 2825 627 2834 639
rect 2745 606 2758 612
rect 2765 607 2773 612
rect 2765 606 2785 607
rect 2745 584 2749 606
rect 2765 584 2769 606
rect 2825 544 2829 627
rect 2885 584 2889 641
rect 2914 639 2918 676
rect 2922 672 2926 676
rect 2922 666 2941 672
rect 2934 653 2941 666
rect 2914 604 2920 627
rect 2934 604 2941 641
rect 2971 639 2975 696
rect 3031 671 3035 676
rect 2966 627 2975 639
rect 2905 598 2920 604
rect 2925 598 2941 604
rect 2905 584 2909 598
rect 2925 584 2929 598
rect 2971 544 2975 627
rect 3022 664 3035 671
rect 3022 619 3026 664
rect 3051 653 3055 676
rect 3046 641 3055 653
rect 3022 596 3026 607
rect 3022 588 3040 596
rect 3036 584 3040 588
rect 3044 584 3048 641
rect 3071 599 3075 676
rect 3133 656 3137 676
rect 3129 649 3137 656
rect 3143 656 3147 676
rect 3143 649 3157 656
rect 3129 633 3135 649
rect 3126 621 3135 633
rect 3066 587 3073 599
rect 3066 544 3070 587
rect 3131 544 3135 621
rect 3151 633 3157 649
rect 3151 621 3154 633
rect 3151 544 3155 621
rect 3212 599 3216 656
rect 3206 587 3216 599
rect 3200 556 3206 587
rect 3220 579 3224 656
rect 3228 599 3232 656
rect 3311 639 3315 696
rect 3371 671 3375 676
rect 3306 627 3315 639
rect 3228 587 3235 599
rect 3247 587 3255 599
rect 3220 560 3226 567
rect 3220 556 3235 560
rect 3200 552 3215 556
rect 3211 544 3215 552
rect 3231 544 3235 556
rect 3251 544 3255 587
rect 3311 544 3315 627
rect 3362 664 3375 671
rect 3362 619 3366 664
rect 3391 653 3395 676
rect 3386 641 3395 653
rect 3362 596 3366 607
rect 3362 588 3380 596
rect 3376 584 3380 588
rect 3384 584 3388 641
rect 3411 599 3415 676
rect 3473 656 3477 676
rect 3469 649 3477 656
rect 3483 656 3487 676
rect 3554 672 3558 676
rect 3539 666 3558 672
rect 3483 649 3497 656
rect 3539 653 3546 666
rect 3469 633 3475 649
rect 3466 621 3475 633
rect 3406 587 3413 599
rect 3406 544 3410 587
rect 3471 544 3475 621
rect 3491 633 3497 649
rect 3491 621 3494 633
rect 3491 544 3495 621
rect 3539 604 3546 641
rect 3562 639 3566 676
rect 3584 653 3588 696
rect 3586 641 3595 653
rect 3560 604 3566 627
rect 3539 598 3555 604
rect 3560 598 3575 604
rect 3551 584 3555 598
rect 3571 584 3575 598
rect 3591 584 3595 641
rect 3651 619 3655 696
rect 3671 619 3675 696
rect 3731 671 3735 676
rect 3722 664 3735 671
rect 3722 619 3726 664
rect 3751 653 3755 676
rect 3746 641 3755 653
rect 3646 607 3655 619
rect 3651 584 3655 607
rect 3659 607 3674 619
rect 3659 584 3663 607
rect 3722 596 3726 607
rect 3722 588 3740 596
rect 3736 584 3740 588
rect 3744 584 3748 641
rect 3771 599 3775 676
rect 3868 599 3872 656
rect 3766 587 3773 599
rect 3845 587 3853 599
rect 3865 587 3872 599
rect 3766 544 3770 587
rect 3845 544 3849 587
rect 3876 579 3880 656
rect 3884 599 3888 656
rect 3931 608 3935 676
rect 3953 647 3957 696
rect 3963 675 3967 696
rect 3983 684 3987 696
rect 3991 692 3995 696
rect 3991 688 4025 692
rect 3983 680 4013 684
rect 3983 679 4001 680
rect 3963 671 3987 675
rect 3884 587 3894 599
rect 3931 596 3933 608
rect 3874 560 3880 567
rect 3865 556 3880 560
rect 3894 556 3900 587
rect 3931 584 3935 596
rect 3953 589 3957 635
rect 3865 544 3869 556
rect 3885 552 3900 556
rect 3885 544 3889 552
rect 3949 583 3957 589
rect 3949 554 3953 583
rect 3981 576 3987 671
rect 3949 547 3957 554
rect 3953 524 3957 547
rect 3961 524 3965 564
rect 3981 544 3985 576
rect 4021 562 4025 688
rect 4037 582 4041 696
rect 4059 684 4063 696
rect 4061 672 4063 684
rect 4069 684 4073 696
rect 4069 672 4071 684
rect 3989 550 4013 552
rect 3989 548 4025 550
rect 3989 544 3993 548
rect 4035 544 4039 570
rect 4053 562 4057 672
rect 4091 664 4095 696
rect 4062 660 4095 664
rect 4062 596 4066 660
rect 4082 611 4086 640
rect 4101 638 4105 696
rect 4121 639 4125 676
rect 4082 603 4091 611
rect 4062 584 4065 596
rect 4055 544 4059 550
rect 4067 544 4071 584
rect 4087 544 4091 603
rect 4101 544 4105 626
rect 4121 584 4125 627
rect 4185 619 4189 696
rect 4205 619 4209 696
rect 4186 607 4201 619
rect 4197 584 4201 607
rect 4205 607 4214 619
rect 4251 608 4255 676
rect 4273 647 4277 696
rect 4283 675 4287 696
rect 4303 684 4307 696
rect 4311 692 4315 696
rect 4311 688 4345 692
rect 4303 680 4333 684
rect 4303 679 4321 680
rect 4283 671 4307 675
rect 4205 584 4209 607
rect 4251 596 4253 608
rect 4251 584 4255 596
rect 4273 589 4277 635
rect 4269 583 4277 589
rect 4269 554 4273 583
rect 4301 576 4307 671
rect 4269 547 4277 554
rect 4273 524 4277 547
rect 4281 524 4285 564
rect 4301 544 4305 576
rect 4341 562 4345 688
rect 4357 582 4361 696
rect 4379 684 4383 696
rect 4381 672 4383 684
rect 4389 684 4393 696
rect 4389 672 4391 684
rect 4309 550 4333 552
rect 4309 548 4345 550
rect 4309 544 4313 548
rect 4355 544 4359 570
rect 4373 562 4377 672
rect 4411 664 4415 696
rect 4382 660 4415 664
rect 4382 596 4386 660
rect 4402 611 4406 640
rect 4421 638 4425 696
rect 4441 639 4445 676
rect 4491 639 4495 696
rect 4554 668 4558 676
rect 4486 627 4495 639
rect 4402 603 4411 611
rect 4382 584 4385 596
rect 4375 544 4379 550
rect 4387 544 4391 584
rect 4407 544 4411 603
rect 4421 544 4425 626
rect 4441 584 4445 627
rect 4491 544 4495 627
rect 4541 661 4558 668
rect 4541 619 4547 661
rect 4562 653 4566 676
rect 4582 662 4586 676
rect 4590 671 4594 676
rect 4590 667 4620 671
rect 4582 655 4595 662
rect 4591 653 4595 655
rect 4591 641 4593 653
rect 4562 612 4566 641
rect 4547 607 4555 612
rect 4535 606 4555 607
rect 4562 606 4575 612
rect 4551 584 4555 606
rect 4571 584 4575 606
rect 4591 584 4595 641
rect 4614 619 4620 667
rect 4692 653 4696 696
rect 5025 708 5029 712
rect 5035 708 5039 716
rect 5055 708 5059 712
rect 5065 708 5069 712
rect 5085 708 5089 716
rect 4685 641 4694 653
rect 4611 607 4614 619
rect 4611 584 4615 607
rect 4685 584 4689 641
rect 4714 639 4718 676
rect 4722 672 4726 676
rect 4722 666 4741 672
rect 4734 653 4741 666
rect 4714 604 4720 627
rect 4734 604 4741 641
rect 4705 598 4720 604
rect 4725 598 4741 604
rect 4785 599 4789 676
rect 4805 653 4809 676
rect 4825 671 4829 676
rect 4825 664 4838 671
rect 4805 641 4814 653
rect 4705 584 4709 598
rect 4725 584 4729 598
rect 4787 587 4794 599
rect 4790 544 4794 587
rect 4812 584 4816 641
rect 4834 619 4838 664
rect 4873 656 4877 676
rect 4869 649 4877 656
rect 4883 656 4887 676
rect 4883 649 4897 656
rect 4869 633 4875 649
rect 4866 621 4875 633
rect 4834 596 4838 607
rect 4820 588 4838 596
rect 4820 584 4824 588
rect 4871 544 4875 621
rect 4891 633 4897 649
rect 4965 639 4969 696
rect 5085 684 5089 688
rect 5085 679 5097 684
rect 4891 621 4894 633
rect 4965 627 4974 639
rect 4891 544 4895 621
rect 4965 544 4969 627
rect 5025 619 5029 668
rect 5035 664 5039 668
rect 5055 622 5059 668
rect 5065 656 5069 668
rect 5065 650 5079 656
rect 5026 607 5029 619
rect 5074 619 5079 650
rect 5093 653 5097 679
rect 5025 584 5029 607
rect 5035 606 5065 610
rect 5035 584 5039 606
rect 5073 601 5078 607
rect 5065 597 5078 601
rect 5055 592 5059 596
rect 5065 592 5069 597
rect 5093 560 5097 641
rect 5132 599 5136 656
rect 5126 587 5136 599
rect 5085 556 5097 560
rect 5120 556 5126 587
rect 5140 579 5144 656
rect 5148 599 5152 656
rect 5231 608 5235 676
rect 5253 647 5257 696
rect 5263 675 5267 696
rect 5283 684 5287 696
rect 5291 692 5295 696
rect 5291 688 5325 692
rect 5283 680 5313 684
rect 5283 679 5301 680
rect 5263 671 5287 675
rect 5148 587 5155 599
rect 5167 587 5175 599
rect 5140 560 5146 567
rect 5140 556 5155 560
rect 5085 552 5089 556
rect 5120 552 5135 556
rect 5131 544 5135 552
rect 5151 544 5155 556
rect 5171 544 5175 587
rect 5231 596 5233 608
rect 5231 584 5235 596
rect 5253 589 5257 635
rect 5055 504 5059 512
rect 5065 508 5069 512
rect 5085 504 5089 512
rect 5249 583 5257 589
rect 5249 554 5253 583
rect 5281 576 5287 671
rect 5249 547 5257 554
rect 5253 524 5257 547
rect 5261 524 5265 564
rect 5281 544 5285 576
rect 5321 562 5325 688
rect 5337 582 5341 696
rect 5359 684 5363 696
rect 5361 672 5363 684
rect 5369 684 5373 696
rect 5369 672 5371 684
rect 5289 550 5313 552
rect 5289 548 5325 550
rect 5289 544 5293 548
rect 5335 544 5339 570
rect 5353 562 5357 672
rect 5391 664 5395 696
rect 5362 660 5395 664
rect 5362 596 5366 660
rect 5382 611 5386 640
rect 5401 638 5405 696
rect 5531 708 5535 716
rect 5551 708 5555 712
rect 5561 708 5565 712
rect 5581 708 5585 716
rect 5591 708 5595 712
rect 5531 684 5535 688
rect 5523 679 5535 684
rect 5421 639 5425 676
rect 5471 653 5475 676
rect 5523 653 5527 679
rect 5551 656 5555 668
rect 5466 641 5475 653
rect 5382 603 5391 611
rect 5362 584 5365 596
rect 5355 544 5359 550
rect 5367 544 5371 584
rect 5387 544 5391 603
rect 5401 544 5405 626
rect 5421 584 5425 627
rect 5471 584 5475 641
rect 5523 560 5527 641
rect 5541 650 5555 656
rect 5541 619 5546 650
rect 5561 622 5565 668
rect 5581 664 5585 668
rect 5542 601 5547 607
rect 5591 619 5595 668
rect 5665 619 5669 696
rect 5685 619 5689 696
rect 5745 619 5749 696
rect 5765 619 5769 696
rect 5825 619 5829 696
rect 5845 619 5849 696
rect 5891 619 5895 696
rect 5911 619 5915 696
rect 5985 619 5989 696
rect 6005 619 6009 696
rect 6051 671 6055 676
rect 6042 664 6055 671
rect 6042 619 6046 664
rect 6071 653 6075 676
rect 6066 641 6075 653
rect 5555 606 5585 610
rect 5542 597 5555 601
rect 5551 592 5555 597
rect 5561 592 5565 596
rect 5523 556 5535 560
rect 5531 552 5535 556
rect 5581 584 5585 606
rect 5591 607 5594 619
rect 5666 607 5681 619
rect 5591 584 5595 607
rect 5677 584 5681 607
rect 5685 607 5694 619
rect 5746 607 5761 619
rect 5685 584 5689 607
rect 5757 584 5761 607
rect 5765 607 5774 619
rect 5826 607 5841 619
rect 5765 584 5769 607
rect 5837 584 5841 607
rect 5845 607 5854 619
rect 5886 607 5895 619
rect 5845 584 5849 607
rect 5891 584 5895 607
rect 5899 607 5914 619
rect 5986 607 6001 619
rect 5899 584 5903 607
rect 5997 584 6001 607
rect 6005 607 6014 619
rect 6005 584 6009 607
rect 6042 596 6046 607
rect 6042 588 6060 596
rect 6056 584 6060 588
rect 6064 584 6068 641
rect 6091 599 6095 676
rect 6151 671 6155 676
rect 6142 664 6155 671
rect 6142 619 6146 664
rect 6171 653 6175 676
rect 6166 641 6175 653
rect 6086 587 6093 599
rect 6142 596 6146 607
rect 6142 588 6160 596
rect 5531 504 5535 512
rect 5551 508 5555 512
rect 5561 504 5565 512
rect 6086 544 6090 587
rect 6156 584 6160 588
rect 6164 584 6168 641
rect 6191 599 6195 676
rect 6273 656 6277 676
rect 6263 649 6277 656
rect 6283 656 6287 676
rect 6283 649 6291 656
rect 6263 633 6269 649
rect 6266 621 6269 633
rect 6186 587 6193 599
rect 6186 544 6190 587
rect 6265 544 6269 621
rect 6285 633 6291 649
rect 6335 639 6339 676
rect 6285 621 6294 633
rect 6355 638 6359 696
rect 6365 664 6369 696
rect 6387 684 6391 696
rect 6389 672 6391 684
rect 6397 684 6401 696
rect 6397 672 6399 684
rect 6365 660 6398 664
rect 6285 544 6289 621
rect 6335 584 6339 627
rect 6355 544 6359 626
rect 6374 611 6378 640
rect 6369 603 6378 611
rect 6369 544 6373 603
rect 6394 596 6398 660
rect 6395 584 6398 596
rect 6389 544 6393 584
rect 6403 562 6407 672
rect 6419 582 6423 696
rect 6465 692 6469 696
rect 6435 688 6469 692
rect 6401 544 6405 550
rect 6421 544 6425 570
rect 6435 562 6439 688
rect 6473 684 6477 696
rect 6447 680 6477 684
rect 6459 679 6477 680
rect 6493 675 6497 696
rect 6473 671 6497 675
rect 6473 576 6479 671
rect 6503 647 6507 696
rect 6503 589 6507 635
rect 6525 608 6529 676
rect 6571 639 6575 696
rect 6631 639 6635 696
rect 6566 627 6575 639
rect 6626 627 6635 639
rect 6527 596 6529 608
rect 6503 583 6511 589
rect 6525 584 6529 596
rect 6447 550 6471 552
rect 6435 548 6471 550
rect 6467 544 6471 548
rect 6475 544 6479 576
rect 6495 524 6499 564
rect 6507 554 6511 583
rect 6503 547 6511 554
rect 6503 524 6507 547
rect 6571 544 6575 627
rect 6631 544 6635 627
rect 31 500 35 504
rect 91 500 95 504
rect 111 500 115 504
rect 171 500 175 504
rect 191 500 195 504
rect 211 500 215 504
rect 271 500 275 504
rect 345 500 349 504
rect 365 500 369 504
rect 385 500 389 504
rect 431 500 435 504
rect 451 500 455 504
rect 471 500 475 504
rect 545 500 549 504
rect 565 500 569 504
rect 625 500 629 504
rect 645 500 649 504
rect 665 500 669 504
rect 711 500 715 504
rect 771 500 775 504
rect 857 500 861 504
rect 865 500 869 504
rect 985 500 989 504
rect 1005 500 1009 504
rect 1025 500 1029 504
rect 1045 500 1049 504
rect 1095 500 1099 504
rect 1115 500 1119 504
rect 1129 500 1133 504
rect 1149 500 1153 504
rect 1161 500 1165 504
rect 1181 500 1185 504
rect 1227 500 1231 504
rect 1235 500 1239 504
rect 1255 500 1259 504
rect 1263 500 1267 504
rect 1285 500 1289 504
rect 1331 500 1335 504
rect 1353 500 1357 504
rect 1411 500 1415 504
rect 1431 500 1435 504
rect 1495 500 1499 504
rect 1515 500 1519 504
rect 1529 500 1533 504
rect 1549 500 1553 504
rect 1561 500 1565 504
rect 1581 500 1585 504
rect 1627 500 1631 504
rect 1635 500 1639 504
rect 1655 500 1659 504
rect 1663 500 1667 504
rect 1685 500 1689 504
rect 1735 500 1739 504
rect 1755 500 1759 504
rect 1769 500 1773 504
rect 1789 500 1793 504
rect 1801 500 1805 504
rect 1821 500 1825 504
rect 1867 500 1871 504
rect 1875 500 1879 504
rect 1895 500 1899 504
rect 1903 500 1907 504
rect 1925 500 1929 504
rect 1975 500 1979 504
rect 1995 500 1999 504
rect 2009 500 2013 504
rect 2029 500 2033 504
rect 2041 500 2045 504
rect 2061 500 2065 504
rect 2107 500 2111 504
rect 2115 500 2119 504
rect 2135 500 2139 504
rect 2143 500 2147 504
rect 2165 500 2169 504
rect 2215 500 2219 504
rect 2235 500 2239 504
rect 2249 500 2253 504
rect 2269 500 2273 504
rect 2281 500 2285 504
rect 2301 500 2305 504
rect 2347 500 2351 504
rect 2355 500 2359 504
rect 2375 500 2379 504
rect 2383 500 2387 504
rect 2405 500 2409 504
rect 2451 500 2455 504
rect 2473 500 2477 504
rect 2481 500 2485 504
rect 2501 500 2505 504
rect 2509 500 2513 504
rect 2555 500 2559 504
rect 2575 500 2579 504
rect 2587 500 2591 504
rect 2607 500 2611 504
rect 2621 500 2625 504
rect 2641 500 2645 504
rect 2705 500 2709 504
rect 2725 500 2729 504
rect 2745 500 2749 504
rect 2765 500 2769 504
rect 2825 500 2829 504
rect 2885 500 2889 504
rect 2905 500 2909 504
rect 2925 500 2929 504
rect 2971 500 2975 504
rect 3036 500 3040 504
rect 3044 500 3048 504
rect 3066 500 3070 504
rect 3131 500 3135 504
rect 3151 500 3155 504
rect 3211 500 3215 504
rect 3231 500 3235 504
rect 3251 500 3255 504
rect 3311 500 3315 504
rect 3376 500 3380 504
rect 3384 500 3388 504
rect 3406 500 3410 504
rect 3471 500 3475 504
rect 3491 500 3495 504
rect 3551 500 3555 504
rect 3571 500 3575 504
rect 3591 500 3595 504
rect 3651 500 3655 504
rect 3659 500 3663 504
rect 3736 500 3740 504
rect 3744 500 3748 504
rect 3766 500 3770 504
rect 3845 500 3849 504
rect 3865 500 3869 504
rect 3885 500 3889 504
rect 3931 500 3935 504
rect 3953 500 3957 504
rect 3961 500 3965 504
rect 3981 500 3985 504
rect 3989 500 3993 504
rect 4035 500 4039 504
rect 4055 500 4059 504
rect 4067 500 4071 504
rect 4087 500 4091 504
rect 4101 500 4105 504
rect 4121 500 4125 504
rect 4197 500 4201 504
rect 4205 500 4209 504
rect 4251 500 4255 504
rect 4273 500 4277 504
rect 4281 500 4285 504
rect 4301 500 4305 504
rect 4309 500 4313 504
rect 4355 500 4359 504
rect 4375 500 4379 504
rect 4387 500 4391 504
rect 4407 500 4411 504
rect 4421 500 4425 504
rect 4441 500 4445 504
rect 4491 500 4495 504
rect 4551 500 4555 504
rect 4571 500 4575 504
rect 4591 500 4595 504
rect 4611 500 4615 504
rect 4685 500 4689 504
rect 4705 500 4709 504
rect 4725 500 4729 504
rect 4790 500 4794 504
rect 4812 500 4816 504
rect 4820 500 4824 504
rect 4871 500 4875 504
rect 4891 500 4895 504
rect 4965 500 4969 504
rect 5025 500 5029 504
rect 5035 500 5039 504
rect 5055 500 5089 504
rect 5131 500 5135 504
rect 5151 500 5155 504
rect 5171 500 5175 504
rect 5231 500 5235 504
rect 5253 500 5257 504
rect 5261 500 5265 504
rect 5281 500 5285 504
rect 5289 500 5293 504
rect 5335 500 5339 504
rect 5355 500 5359 504
rect 5367 500 5371 504
rect 5387 500 5391 504
rect 5401 500 5405 504
rect 5421 500 5425 504
rect 5471 500 5475 504
rect 5531 500 5565 504
rect 5581 500 5585 504
rect 5591 500 5595 504
rect 5677 500 5681 504
rect 5685 500 5689 504
rect 5757 500 5761 504
rect 5765 500 5769 504
rect 5837 500 5841 504
rect 5845 500 5849 504
rect 5891 500 5895 504
rect 5899 500 5903 504
rect 5997 500 6001 504
rect 6005 500 6009 504
rect 6056 500 6060 504
rect 6064 500 6068 504
rect 6086 500 6090 504
rect 6156 500 6160 504
rect 6164 500 6168 504
rect 6186 500 6190 504
rect 6265 500 6269 504
rect 6285 500 6289 504
rect 6335 500 6339 504
rect 6355 500 6359 504
rect 6369 500 6373 504
rect 6389 500 6393 504
rect 6401 500 6405 504
rect 6421 500 6425 504
rect 6467 500 6471 504
rect 6475 500 6479 504
rect 6495 500 6499 504
rect 6503 500 6507 504
rect 6525 500 6529 504
rect 6571 500 6575 504
rect 6631 500 6635 504
rect 31 476 35 480
rect 53 476 57 480
rect 61 476 65 480
rect 81 476 85 480
rect 89 476 93 480
rect 135 476 139 480
rect 155 476 159 480
rect 167 476 171 480
rect 187 476 191 480
rect 201 476 205 480
rect 221 476 225 480
rect 275 476 279 480
rect 295 476 299 480
rect 309 476 313 480
rect 329 476 333 480
rect 341 476 345 480
rect 361 476 365 480
rect 407 476 411 480
rect 415 476 419 480
rect 435 476 439 480
rect 443 476 447 480
rect 465 476 469 480
rect 511 476 515 480
rect 531 476 535 480
rect 551 476 555 480
rect 611 476 615 480
rect 619 476 623 480
rect 717 476 721 480
rect 725 476 729 480
rect 771 476 775 480
rect 791 476 795 480
rect 865 476 869 480
rect 915 476 919 480
rect 935 476 939 480
rect 949 476 953 480
rect 969 476 973 480
rect 981 476 985 480
rect 1001 476 1005 480
rect 1047 476 1051 480
rect 1055 476 1059 480
rect 1075 476 1079 480
rect 1083 476 1087 480
rect 1105 476 1109 480
rect 1163 476 1167 480
rect 1185 476 1189 480
rect 1231 476 1235 480
rect 1253 476 1257 480
rect 1311 476 1315 480
rect 1333 476 1337 480
rect 1405 476 1409 480
rect 1456 476 1460 480
rect 1464 476 1468 480
rect 1486 476 1490 480
rect 1565 476 1569 480
rect 1616 476 1620 480
rect 1624 476 1628 480
rect 1646 476 1650 480
rect 1715 476 1719 480
rect 1735 476 1739 480
rect 1749 476 1753 480
rect 1769 476 1773 480
rect 1781 476 1785 480
rect 1801 476 1805 480
rect 1847 476 1851 480
rect 1855 476 1859 480
rect 1875 476 1879 480
rect 1883 476 1887 480
rect 1905 476 1909 480
rect 1965 476 1969 480
rect 2025 476 2029 480
rect 2076 476 2080 480
rect 2084 476 2088 480
rect 2106 476 2110 480
rect 2171 476 2175 480
rect 2231 476 2235 480
rect 2241 476 2245 480
rect 2271 476 2275 480
rect 2281 476 2285 480
rect 2370 476 2374 480
rect 2392 476 2396 480
rect 2400 476 2404 480
rect 2451 476 2455 480
rect 2459 476 2463 480
rect 2535 476 2539 480
rect 2555 476 2559 480
rect 2569 476 2573 480
rect 2589 476 2593 480
rect 2601 476 2605 480
rect 2621 476 2625 480
rect 2667 476 2671 480
rect 2675 476 2679 480
rect 2695 476 2699 480
rect 2703 476 2707 480
rect 2725 476 2729 480
rect 2790 476 2794 480
rect 2812 476 2816 480
rect 2820 476 2824 480
rect 2871 476 2875 480
rect 2879 476 2883 480
rect 2955 476 2959 480
rect 2975 476 2979 480
rect 2989 476 2993 480
rect 3009 476 3013 480
rect 3021 476 3025 480
rect 3041 476 3045 480
rect 3087 476 3091 480
rect 3095 476 3099 480
rect 3115 476 3119 480
rect 3123 476 3127 480
rect 3145 476 3149 480
rect 3191 476 3195 480
rect 3211 476 3215 480
rect 3290 476 3294 480
rect 3312 476 3316 480
rect 3320 476 3324 480
rect 3371 476 3375 480
rect 3379 476 3383 480
rect 3465 476 3469 480
rect 3485 476 3489 480
rect 3505 476 3509 480
rect 3556 476 3560 480
rect 3564 476 3568 480
rect 3586 476 3590 480
rect 3651 476 3655 480
rect 3659 476 3663 480
rect 3731 476 3735 480
rect 3751 476 3755 480
rect 3771 476 3775 480
rect 3857 476 3861 480
rect 3865 476 3869 480
rect 3916 476 3920 480
rect 3924 476 3928 480
rect 3946 476 3950 480
rect 4025 476 4029 480
rect 4045 476 4049 480
rect 4065 476 4069 480
rect 4111 476 4115 480
rect 4119 476 4123 480
rect 4191 476 4195 480
rect 4213 476 4217 480
rect 4221 476 4225 480
rect 4241 476 4245 480
rect 4249 476 4253 480
rect 4295 476 4299 480
rect 4315 476 4319 480
rect 4327 476 4331 480
rect 4347 476 4351 480
rect 4361 476 4365 480
rect 4381 476 4385 480
rect 4431 476 4435 480
rect 4439 476 4443 480
rect 4530 476 4534 480
rect 4552 476 4556 480
rect 4560 476 4564 480
rect 4611 476 4615 480
rect 4619 476 4623 480
rect 4715 476 4719 480
rect 4725 476 4729 480
rect 4755 476 4759 480
rect 4765 476 4769 480
rect 4825 476 4829 480
rect 4875 476 4879 480
rect 4895 476 4899 480
rect 4909 476 4913 480
rect 4929 476 4933 480
rect 4941 476 4945 480
rect 4961 476 4965 480
rect 5007 476 5011 480
rect 5015 476 5019 480
rect 5035 476 5039 480
rect 5043 476 5047 480
rect 5065 476 5069 480
rect 5125 476 5129 480
rect 5145 476 5149 480
rect 5165 476 5169 480
rect 5211 476 5215 480
rect 5219 476 5223 480
rect 5310 476 5314 480
rect 5332 476 5336 480
rect 5340 476 5344 480
rect 5391 476 5395 480
rect 5399 476 5403 480
rect 5471 476 5475 480
rect 5491 476 5495 480
rect 5511 476 5515 480
rect 5571 476 5575 480
rect 5591 476 5595 480
rect 5611 476 5615 480
rect 5676 476 5680 480
rect 5684 476 5688 480
rect 5706 476 5710 480
rect 5785 476 5789 480
rect 5805 476 5809 480
rect 5870 476 5874 480
rect 5892 476 5896 480
rect 5900 476 5904 480
rect 5956 476 5960 480
rect 5964 476 5968 480
rect 5986 476 5990 480
rect 6056 476 6060 480
rect 6064 476 6068 480
rect 6086 476 6090 480
rect 6177 476 6181 480
rect 6185 476 6189 480
rect 6257 476 6261 480
rect 6265 476 6269 480
rect 6335 476 6339 480
rect 6345 476 6349 480
rect 6375 476 6379 480
rect 6385 476 6389 480
rect 6435 476 6439 480
rect 6455 476 6459 480
rect 6469 476 6473 480
rect 6489 476 6493 480
rect 6501 476 6505 480
rect 6521 476 6525 480
rect 6567 476 6571 480
rect 6575 476 6579 480
rect 6595 476 6599 480
rect 6603 476 6607 480
rect 6625 476 6629 480
rect 53 433 57 456
rect 49 426 57 433
rect 49 397 53 426
rect 61 416 65 456
rect 81 404 85 436
rect 89 432 93 436
rect 89 430 125 432
rect 89 428 113 430
rect 31 384 35 396
rect 49 391 57 397
rect 31 372 33 384
rect 31 304 35 372
rect 53 345 57 391
rect 53 284 57 333
rect 81 309 87 404
rect 63 305 87 309
rect 63 284 67 305
rect 83 300 101 301
rect 83 296 113 300
rect 83 284 87 296
rect 121 292 125 418
rect 135 410 139 436
rect 155 430 159 436
rect 91 288 125 292
rect 91 284 95 288
rect 137 284 141 398
rect 153 308 157 418
rect 167 396 171 436
rect 162 384 165 396
rect 162 320 166 384
rect 187 377 191 436
rect 182 369 191 377
rect 182 340 186 369
rect 201 354 205 436
rect 221 353 225 396
rect 275 353 279 396
rect 295 354 299 436
rect 309 377 313 436
rect 329 396 333 436
rect 341 430 345 436
rect 335 384 338 396
rect 309 369 318 377
rect 162 316 195 320
rect 161 296 163 308
rect 159 284 163 296
rect 169 296 171 308
rect 169 284 173 296
rect 191 284 195 316
rect 201 284 205 342
rect 221 304 225 341
rect 275 304 279 341
rect 295 284 299 342
rect 314 340 318 369
rect 334 320 338 384
rect 305 316 338 320
rect 305 284 309 316
rect 343 308 347 418
rect 361 410 365 436
rect 407 432 411 436
rect 375 430 411 432
rect 387 428 411 430
rect 329 296 331 308
rect 327 284 331 296
rect 337 296 339 308
rect 337 284 341 296
rect 359 284 363 398
rect 375 292 379 418
rect 415 404 419 436
rect 435 416 439 456
rect 443 433 447 456
rect 443 426 451 433
rect 413 309 419 404
rect 447 397 451 426
rect 443 391 451 397
rect 511 428 515 436
rect 500 424 515 428
rect 531 424 535 436
rect 443 345 447 391
rect 465 384 469 396
rect 500 393 506 424
rect 520 420 535 424
rect 520 413 526 420
rect 467 372 469 384
rect 506 381 516 393
rect 413 305 437 309
rect 399 300 417 301
rect 387 296 417 300
rect 375 288 409 292
rect 405 284 409 288
rect 413 284 417 296
rect 433 284 437 305
rect 443 284 447 333
rect 465 304 469 372
rect 512 324 516 381
rect 520 324 524 401
rect 551 393 555 436
rect 528 381 535 393
rect 547 381 555 393
rect 528 324 532 381
rect 611 373 615 396
rect 606 361 615 373
rect 619 373 623 396
rect 717 373 721 396
rect 619 361 634 373
rect 706 361 721 373
rect 725 373 729 396
rect 725 361 734 373
rect 611 284 615 361
rect 631 284 635 361
rect 705 284 709 361
rect 725 284 729 361
rect 771 359 775 436
rect 766 347 775 359
rect 769 331 775 347
rect 791 359 795 436
rect 791 347 794 359
rect 865 353 869 436
rect 915 353 919 396
rect 935 354 939 436
rect 949 377 953 436
rect 969 396 973 436
rect 981 430 985 436
rect 975 384 978 396
rect 949 369 958 377
rect 791 331 797 347
rect 769 324 777 331
rect 773 304 777 324
rect 783 324 797 331
rect 865 341 874 353
rect 783 304 787 324
rect 865 284 869 341
rect 915 304 919 341
rect 935 284 939 342
rect 954 340 958 369
rect 974 320 978 384
rect 945 316 978 320
rect 945 284 949 316
rect 983 308 987 418
rect 1001 410 1005 436
rect 1047 432 1051 436
rect 1015 430 1051 432
rect 1027 428 1051 430
rect 969 296 971 308
rect 967 284 971 296
rect 977 296 979 308
rect 977 284 981 296
rect 999 284 1003 398
rect 1015 292 1019 418
rect 1055 404 1059 436
rect 1075 416 1079 456
rect 1083 433 1087 456
rect 1083 426 1091 433
rect 1053 309 1059 404
rect 1087 397 1091 426
rect 1083 391 1091 397
rect 1083 345 1087 391
rect 1105 384 1109 396
rect 1107 372 1109 384
rect 1163 390 1167 396
rect 1163 378 1165 390
rect 1053 305 1077 309
rect 1039 300 1057 301
rect 1027 296 1057 300
rect 1015 288 1049 292
rect 1045 284 1049 288
rect 1053 284 1057 296
rect 1073 284 1077 305
rect 1083 284 1087 333
rect 1105 304 1109 372
rect 1185 373 1189 436
rect 1231 373 1235 436
rect 1253 390 1257 396
rect 1255 378 1257 390
rect 1311 373 1315 436
rect 1333 390 1337 396
rect 1335 378 1337 390
rect 1185 361 1194 373
rect 1226 361 1235 373
rect 1306 361 1315 373
rect 1163 310 1165 322
rect 1163 304 1167 310
rect 1185 284 1189 361
rect 1231 284 1235 361
rect 1255 310 1257 322
rect 1253 304 1257 310
rect 1311 284 1315 361
rect 1405 353 1409 436
rect 1456 392 1460 396
rect 1442 384 1460 392
rect 1442 373 1446 384
rect 1405 341 1414 353
rect 1335 310 1337 322
rect 1333 304 1337 310
rect 1405 284 1409 341
rect 1442 316 1446 361
rect 1464 339 1468 396
rect 1486 393 1490 436
rect 1486 381 1493 393
rect 1466 327 1475 339
rect 1442 309 1455 316
rect 1451 304 1455 309
rect 1471 304 1475 327
rect 1491 304 1495 381
rect 1565 353 1569 436
rect 1616 392 1620 396
rect 1602 384 1620 392
rect 1602 373 1606 384
rect 1565 341 1574 353
rect 1565 284 1569 341
rect 1602 316 1606 361
rect 1624 339 1628 396
rect 1646 393 1650 436
rect 1646 381 1653 393
rect 1626 327 1635 339
rect 1602 309 1615 316
rect 1611 304 1615 309
rect 1631 304 1635 327
rect 1651 304 1655 381
rect 1715 353 1719 396
rect 1735 354 1739 436
rect 1749 377 1753 436
rect 1769 396 1773 436
rect 1781 430 1785 436
rect 1775 384 1778 396
rect 1749 369 1758 377
rect 1715 304 1719 341
rect 1735 284 1739 342
rect 1754 340 1758 369
rect 1774 320 1778 384
rect 1745 316 1778 320
rect 1745 284 1749 316
rect 1783 308 1787 418
rect 1801 410 1805 436
rect 1847 432 1851 436
rect 1815 430 1851 432
rect 1827 428 1851 430
rect 1769 296 1771 308
rect 1767 284 1771 296
rect 1777 296 1779 308
rect 1777 284 1781 296
rect 1799 284 1803 398
rect 1815 292 1819 418
rect 1855 404 1859 436
rect 1875 416 1879 456
rect 1883 433 1887 456
rect 1883 426 1891 433
rect 1853 309 1859 404
rect 1887 397 1891 426
rect 1883 391 1891 397
rect 1883 345 1887 391
rect 1905 384 1909 396
rect 1907 372 1909 384
rect 1853 305 1877 309
rect 1839 300 1857 301
rect 1827 296 1857 300
rect 1815 288 1849 292
rect 1845 284 1849 288
rect 1853 284 1857 296
rect 1873 284 1877 305
rect 1883 284 1887 333
rect 1905 304 1909 372
rect 1965 353 1969 436
rect 2025 353 2029 436
rect 2076 392 2080 396
rect 2062 384 2080 392
rect 2062 373 2066 384
rect 1965 341 1974 353
rect 2025 341 2034 353
rect 1965 284 1969 341
rect 2025 284 2029 341
rect 2062 316 2066 361
rect 2084 339 2088 396
rect 2106 393 2110 436
rect 2106 381 2113 393
rect 2086 327 2095 339
rect 2062 309 2075 316
rect 2071 304 2075 309
rect 2091 304 2095 327
rect 2111 304 2115 381
rect 2171 353 2175 436
rect 2231 392 2235 396
rect 2221 388 2235 392
rect 2241 392 2245 396
rect 2241 388 2255 392
rect 2221 373 2226 388
rect 2166 341 2175 353
rect 2171 284 2175 341
rect 2220 315 2226 361
rect 2249 339 2255 388
rect 2271 339 2275 396
rect 2281 392 2285 396
rect 2370 393 2374 436
rect 2281 388 2295 392
rect 2291 373 2295 388
rect 2367 381 2374 393
rect 2291 361 2293 373
rect 2246 327 2255 339
rect 2220 311 2235 315
rect 2231 304 2235 311
rect 2251 304 2255 327
rect 2271 304 2275 327
rect 2291 304 2295 361
rect 2365 304 2369 381
rect 2392 339 2396 396
rect 2400 392 2404 396
rect 2400 384 2418 392
rect 2414 373 2418 384
rect 2451 373 2455 396
rect 2446 361 2455 373
rect 2459 373 2463 396
rect 2459 361 2474 373
rect 2385 327 2394 339
rect 2385 304 2389 327
rect 2414 316 2418 361
rect 2405 309 2418 316
rect 2405 304 2409 309
rect 2451 284 2455 361
rect 2471 284 2475 361
rect 2535 353 2539 396
rect 2555 354 2559 436
rect 2569 377 2573 436
rect 2589 396 2593 436
rect 2601 430 2605 436
rect 2595 384 2598 396
rect 2569 369 2578 377
rect 2535 304 2539 341
rect 2555 284 2559 342
rect 2574 340 2578 369
rect 2594 320 2598 384
rect 2565 316 2598 320
rect 2565 284 2569 316
rect 2603 308 2607 418
rect 2621 410 2625 436
rect 2667 432 2671 436
rect 2635 430 2671 432
rect 2647 428 2671 430
rect 2589 296 2591 308
rect 2587 284 2591 296
rect 2597 296 2599 308
rect 2597 284 2601 296
rect 2619 284 2623 398
rect 2635 292 2639 418
rect 2675 404 2679 436
rect 2695 416 2699 456
rect 2703 433 2707 456
rect 2703 426 2711 433
rect 2673 309 2679 404
rect 2707 397 2711 426
rect 2703 391 2711 397
rect 2703 345 2707 391
rect 2725 384 2729 396
rect 2790 393 2794 436
rect 2727 372 2729 384
rect 2787 381 2794 393
rect 2673 305 2697 309
rect 2659 300 2677 301
rect 2647 296 2677 300
rect 2635 288 2669 292
rect 2665 284 2669 288
rect 2673 284 2677 296
rect 2693 284 2697 305
rect 2703 284 2707 333
rect 2725 304 2729 372
rect 2785 304 2789 381
rect 2812 339 2816 396
rect 2820 392 2824 396
rect 2820 384 2838 392
rect 2834 373 2838 384
rect 2871 373 2875 396
rect 2866 361 2875 373
rect 2879 373 2883 396
rect 2879 361 2894 373
rect 2805 327 2814 339
rect 2805 304 2809 327
rect 2834 316 2838 361
rect 2825 309 2838 316
rect 2825 304 2829 309
rect 2871 284 2875 361
rect 2891 284 2895 361
rect 2955 353 2959 396
rect 2975 354 2979 436
rect 2989 377 2993 436
rect 3009 396 3013 436
rect 3021 430 3025 436
rect 3015 384 3018 396
rect 2989 369 2998 377
rect 2955 304 2959 341
rect 2975 284 2979 342
rect 2994 340 2998 369
rect 3014 320 3018 384
rect 2985 316 3018 320
rect 2985 284 2989 316
rect 3023 308 3027 418
rect 3041 410 3045 436
rect 3087 432 3091 436
rect 3055 430 3091 432
rect 3067 428 3091 430
rect 3009 296 3011 308
rect 3007 284 3011 296
rect 3017 296 3019 308
rect 3017 284 3021 296
rect 3039 284 3043 398
rect 3055 292 3059 418
rect 3095 404 3099 436
rect 3115 416 3119 456
rect 3123 433 3127 456
rect 3123 426 3131 433
rect 3093 309 3099 404
rect 3127 397 3131 426
rect 3123 391 3131 397
rect 3123 345 3127 391
rect 3145 384 3149 396
rect 3147 372 3149 384
rect 3093 305 3117 309
rect 3079 300 3097 301
rect 3067 296 3097 300
rect 3055 288 3089 292
rect 3085 284 3089 288
rect 3093 284 3097 296
rect 3113 284 3117 305
rect 3123 284 3127 333
rect 3145 304 3149 372
rect 3191 359 3195 436
rect 3186 347 3195 359
rect 3189 331 3195 347
rect 3211 359 3215 436
rect 3290 393 3294 436
rect 3287 381 3294 393
rect 3211 347 3214 359
rect 3211 331 3217 347
rect 3189 324 3197 331
rect 3193 304 3197 324
rect 3203 324 3217 331
rect 3203 304 3207 324
rect 3285 304 3289 381
rect 3312 339 3316 396
rect 3320 392 3324 396
rect 3320 384 3338 392
rect 3334 373 3338 384
rect 3371 373 3375 396
rect 3366 361 3375 373
rect 3379 373 3383 396
rect 3379 361 3394 373
rect 3305 327 3314 339
rect 3305 304 3309 327
rect 3334 316 3338 361
rect 3325 309 3338 316
rect 3325 304 3329 309
rect 3371 284 3375 361
rect 3391 284 3395 361
rect 3465 339 3469 396
rect 3485 382 3489 396
rect 3505 382 3509 396
rect 3556 392 3560 396
rect 3542 384 3560 392
rect 3485 376 3500 382
rect 3505 376 3521 382
rect 3494 353 3500 376
rect 3465 327 3474 339
rect 3472 284 3476 327
rect 3494 304 3498 341
rect 3514 339 3521 376
rect 3542 373 3546 384
rect 3514 314 3521 327
rect 3502 308 3521 314
rect 3542 316 3546 361
rect 3564 339 3568 396
rect 3586 393 3590 436
rect 3586 381 3593 393
rect 3566 327 3575 339
rect 3542 309 3555 316
rect 3502 304 3506 308
rect 3551 304 3555 309
rect 3571 304 3575 327
rect 3591 304 3595 381
rect 3651 373 3655 396
rect 3646 361 3655 373
rect 3659 373 3663 396
rect 3731 382 3735 396
rect 3751 382 3755 396
rect 3719 376 3735 382
rect 3740 376 3755 382
rect 3659 361 3674 373
rect 3651 284 3655 361
rect 3671 284 3675 361
rect 3719 339 3726 376
rect 3740 353 3746 376
rect 3719 314 3726 327
rect 3719 308 3738 314
rect 3734 304 3738 308
rect 3742 304 3746 341
rect 3771 339 3775 396
rect 3857 373 3861 396
rect 3846 361 3861 373
rect 3865 373 3869 396
rect 3916 392 3920 396
rect 3902 384 3920 392
rect 3902 373 3906 384
rect 3865 361 3874 373
rect 3766 327 3775 339
rect 3764 284 3768 327
rect 3845 284 3849 361
rect 3865 284 3869 361
rect 3902 316 3906 361
rect 3924 339 3928 396
rect 3946 393 3950 436
rect 4025 393 4029 436
rect 4045 424 4049 436
rect 4065 428 4069 436
rect 4065 424 4080 428
rect 4045 420 4060 424
rect 4054 413 4060 420
rect 3946 381 3953 393
rect 4025 381 4033 393
rect 4045 381 4052 393
rect 3926 327 3935 339
rect 3902 309 3915 316
rect 3911 304 3915 309
rect 3931 304 3935 327
rect 3951 304 3955 381
rect 4048 324 4052 381
rect 4056 324 4060 401
rect 4074 393 4080 424
rect 4213 433 4217 456
rect 4209 426 4217 433
rect 4209 397 4213 426
rect 4221 416 4225 456
rect 4241 404 4245 436
rect 4249 432 4253 436
rect 4249 430 4285 432
rect 4249 428 4273 430
rect 4064 381 4074 393
rect 4064 324 4068 381
rect 4111 373 4115 396
rect 4106 361 4115 373
rect 4119 373 4123 396
rect 4191 384 4195 396
rect 4209 391 4217 397
rect 4119 361 4134 373
rect 4191 372 4193 384
rect 4111 284 4115 361
rect 4131 284 4135 361
rect 4191 304 4195 372
rect 4213 345 4217 391
rect 4213 284 4217 333
rect 4241 309 4247 404
rect 4223 305 4247 309
rect 4223 284 4227 305
rect 4243 300 4261 301
rect 4243 296 4273 300
rect 4243 284 4247 296
rect 4281 292 4285 418
rect 4295 410 4299 436
rect 4315 430 4319 436
rect 4251 288 4285 292
rect 4251 284 4255 288
rect 4297 284 4301 398
rect 4313 308 4317 418
rect 4327 396 4331 436
rect 4322 384 4325 396
rect 4322 320 4326 384
rect 4347 377 4351 436
rect 4342 369 4351 377
rect 4342 340 4346 369
rect 4361 354 4365 436
rect 4381 353 4385 396
rect 4431 373 4435 396
rect 4426 361 4435 373
rect 4439 373 4443 396
rect 4530 393 4534 436
rect 4527 381 4534 393
rect 4439 361 4454 373
rect 4322 316 4355 320
rect 4321 296 4323 308
rect 4319 284 4323 296
rect 4329 296 4331 308
rect 4329 284 4333 296
rect 4351 284 4355 316
rect 4361 284 4365 342
rect 4381 304 4385 341
rect 4431 284 4435 361
rect 4451 284 4455 361
rect 4525 304 4529 381
rect 4552 339 4556 396
rect 4560 392 4564 396
rect 4560 384 4578 392
rect 4574 373 4578 384
rect 4611 373 4615 396
rect 4606 361 4615 373
rect 4619 373 4623 396
rect 4715 392 4719 396
rect 4705 388 4719 392
rect 4705 373 4709 388
rect 4619 361 4634 373
rect 4707 361 4709 373
rect 4545 327 4554 339
rect 4545 304 4549 327
rect 4574 316 4578 361
rect 4565 309 4578 316
rect 4565 304 4569 309
rect 4611 284 4615 361
rect 4631 284 4635 361
rect 4705 304 4709 361
rect 4725 339 4729 396
rect 4755 392 4759 396
rect 4745 388 4759 392
rect 4765 392 4769 396
rect 4765 388 4779 392
rect 4745 339 4751 388
rect 4774 373 4779 388
rect 4745 327 4754 339
rect 4725 304 4729 327
rect 4745 304 4749 327
rect 4774 315 4780 361
rect 4765 311 4780 315
rect 4825 353 4829 436
rect 4875 353 4879 396
rect 4895 354 4899 436
rect 4909 377 4913 436
rect 4929 396 4933 436
rect 4941 430 4945 436
rect 4935 384 4938 396
rect 4909 369 4918 377
rect 4825 341 4834 353
rect 4765 304 4769 311
rect 4825 284 4829 341
rect 4875 304 4879 341
rect 4895 284 4899 342
rect 4914 340 4918 369
rect 4934 320 4938 384
rect 4905 316 4938 320
rect 4905 284 4909 316
rect 4943 308 4947 418
rect 4961 410 4965 436
rect 5007 432 5011 436
rect 4975 430 5011 432
rect 4987 428 5011 430
rect 4929 296 4931 308
rect 4927 284 4931 296
rect 4937 296 4939 308
rect 4937 284 4941 296
rect 4959 284 4963 398
rect 4975 292 4979 418
rect 5015 404 5019 436
rect 5035 416 5039 456
rect 5043 433 5047 456
rect 5043 426 5051 433
rect 5013 309 5019 404
rect 5047 397 5051 426
rect 5043 391 5051 397
rect 5043 345 5047 391
rect 5065 384 5069 396
rect 5067 372 5069 384
rect 5013 305 5037 309
rect 4999 300 5017 301
rect 4987 296 5017 300
rect 4975 288 5009 292
rect 5005 284 5009 288
rect 5013 284 5017 296
rect 5033 284 5037 305
rect 5043 284 5047 333
rect 5065 304 5069 372
rect 5125 339 5129 396
rect 5145 382 5149 396
rect 5165 382 5169 396
rect 5145 376 5160 382
rect 5165 376 5181 382
rect 5154 353 5160 376
rect 5125 327 5134 339
rect 5132 284 5136 327
rect 5154 304 5158 341
rect 5174 339 5181 376
rect 5211 373 5215 396
rect 5206 361 5215 373
rect 5219 373 5223 396
rect 5310 393 5314 436
rect 5571 428 5575 436
rect 5560 424 5575 428
rect 5591 424 5595 436
rect 5307 381 5314 393
rect 5219 361 5234 373
rect 5174 314 5181 327
rect 5162 308 5181 314
rect 5162 304 5166 308
rect 5211 284 5215 361
rect 5231 284 5235 361
rect 5305 304 5309 381
rect 5332 339 5336 396
rect 5340 392 5344 396
rect 5340 384 5358 392
rect 5354 373 5358 384
rect 5391 373 5395 396
rect 5386 361 5395 373
rect 5399 373 5403 396
rect 5471 382 5475 396
rect 5491 382 5495 396
rect 5459 376 5475 382
rect 5480 376 5495 382
rect 5399 361 5414 373
rect 5325 327 5334 339
rect 5325 304 5329 327
rect 5354 316 5358 361
rect 5345 309 5358 316
rect 5345 304 5349 309
rect 5391 284 5395 361
rect 5411 284 5415 361
rect 5459 339 5466 376
rect 5480 353 5486 376
rect 5459 314 5466 327
rect 5459 308 5478 314
rect 5474 304 5478 308
rect 5482 304 5486 341
rect 5511 339 5515 396
rect 5560 393 5566 424
rect 5580 420 5595 424
rect 5580 413 5586 420
rect 5566 381 5576 393
rect 5506 327 5515 339
rect 5504 284 5508 327
rect 5572 324 5576 381
rect 5580 324 5584 401
rect 5611 393 5615 436
rect 5588 381 5595 393
rect 5607 381 5615 393
rect 5676 392 5680 396
rect 5662 384 5680 392
rect 5588 324 5592 381
rect 5662 373 5666 384
rect 5662 316 5666 361
rect 5684 339 5688 396
rect 5706 393 5710 436
rect 5706 381 5713 393
rect 5686 327 5695 339
rect 5662 309 5675 316
rect 5671 304 5675 309
rect 5691 304 5695 327
rect 5711 304 5715 381
rect 5785 359 5789 436
rect 5786 347 5789 359
rect 5783 331 5789 347
rect 5805 359 5809 436
rect 5870 393 5874 436
rect 5867 381 5874 393
rect 5805 347 5814 359
rect 5805 331 5811 347
rect 5783 324 5797 331
rect 5793 304 5797 324
rect 5803 324 5811 331
rect 5803 304 5807 324
rect 5865 304 5869 381
rect 5892 339 5896 396
rect 5900 392 5904 396
rect 5956 392 5960 396
rect 5900 384 5918 392
rect 5914 373 5918 384
rect 5942 384 5960 392
rect 5942 373 5946 384
rect 5885 327 5894 339
rect 5885 304 5889 327
rect 5914 316 5918 361
rect 5905 309 5918 316
rect 5942 316 5946 361
rect 5964 339 5968 396
rect 5986 393 5990 436
rect 5986 381 5993 393
rect 6056 392 6060 396
rect 6042 384 6060 392
rect 5966 327 5975 339
rect 5942 309 5955 316
rect 5905 304 5909 309
rect 5951 304 5955 309
rect 5971 304 5975 327
rect 5991 304 5995 381
rect 6042 373 6046 384
rect 6042 316 6046 361
rect 6064 339 6068 396
rect 6086 393 6090 436
rect 6086 381 6093 393
rect 6066 327 6075 339
rect 6042 309 6055 316
rect 6051 304 6055 309
rect 6071 304 6075 327
rect 6091 304 6095 381
rect 6177 373 6181 396
rect 6166 361 6181 373
rect 6185 373 6189 396
rect 6257 373 6261 396
rect 6185 361 6194 373
rect 6246 361 6261 373
rect 6265 373 6269 396
rect 6335 392 6339 396
rect 6325 388 6339 392
rect 6325 373 6329 388
rect 6265 361 6274 373
rect 6327 361 6329 373
rect 6165 284 6169 361
rect 6185 284 6189 361
rect 6245 284 6249 361
rect 6265 284 6269 361
rect 6325 304 6329 361
rect 6345 339 6349 396
rect 6375 392 6379 396
rect 6365 388 6379 392
rect 6385 392 6389 396
rect 6385 388 6399 392
rect 6365 339 6371 388
rect 6394 373 6399 388
rect 6365 327 6374 339
rect 6345 304 6349 327
rect 6365 304 6369 327
rect 6394 315 6400 361
rect 6435 353 6439 396
rect 6455 354 6459 436
rect 6469 377 6473 436
rect 6489 396 6493 436
rect 6501 430 6505 436
rect 6495 384 6498 396
rect 6469 369 6478 377
rect 6385 311 6400 315
rect 6385 304 6389 311
rect 6435 304 6439 341
rect 6455 284 6459 342
rect 6474 340 6478 369
rect 6494 320 6498 384
rect 6465 316 6498 320
rect 6465 284 6469 316
rect 6503 308 6507 418
rect 6521 410 6525 436
rect 6567 432 6571 436
rect 6535 430 6571 432
rect 6547 428 6571 430
rect 6489 296 6491 308
rect 6487 284 6491 296
rect 6497 296 6499 308
rect 6497 284 6501 296
rect 6519 284 6523 398
rect 6535 292 6539 418
rect 6575 404 6579 436
rect 6595 416 6599 456
rect 6603 433 6607 456
rect 6603 426 6611 433
rect 6573 309 6579 404
rect 6607 397 6611 426
rect 6603 391 6611 397
rect 6603 345 6607 391
rect 6625 384 6629 396
rect 6627 372 6629 384
rect 6573 305 6597 309
rect 6559 300 6577 301
rect 6547 296 6577 300
rect 6535 288 6569 292
rect 6565 284 6569 288
rect 6573 284 6577 296
rect 6593 284 6597 305
rect 6603 284 6607 333
rect 6625 304 6629 372
rect 31 260 35 264
rect 53 260 57 264
rect 63 260 67 264
rect 83 260 87 264
rect 91 260 95 264
rect 137 260 141 264
rect 159 260 163 264
rect 169 260 173 264
rect 191 260 195 264
rect 201 260 205 264
rect 221 260 225 264
rect 275 260 279 264
rect 295 260 299 264
rect 305 260 309 264
rect 327 260 331 264
rect 337 260 341 264
rect 359 260 363 264
rect 405 260 409 264
rect 413 260 417 264
rect 433 260 437 264
rect 443 260 447 264
rect 465 260 469 264
rect 512 260 516 264
rect 520 260 524 264
rect 528 260 532 264
rect 611 260 615 264
rect 631 260 635 264
rect 705 260 709 264
rect 725 260 729 264
rect 773 260 777 264
rect 783 260 787 264
rect 865 260 869 264
rect 915 260 919 264
rect 935 260 939 264
rect 945 260 949 264
rect 967 260 971 264
rect 977 260 981 264
rect 999 260 1003 264
rect 1045 260 1049 264
rect 1053 260 1057 264
rect 1073 260 1077 264
rect 1083 260 1087 264
rect 1105 260 1109 264
rect 1163 260 1167 264
rect 1185 260 1189 264
rect 1231 260 1235 264
rect 1253 260 1257 264
rect 1311 260 1315 264
rect 1333 260 1337 264
rect 1405 260 1409 264
rect 1451 260 1455 264
rect 1471 260 1475 264
rect 1491 260 1495 264
rect 1565 260 1569 264
rect 1611 260 1615 264
rect 1631 260 1635 264
rect 1651 260 1655 264
rect 1715 260 1719 264
rect 1735 260 1739 264
rect 1745 260 1749 264
rect 1767 260 1771 264
rect 1777 260 1781 264
rect 1799 260 1803 264
rect 1845 260 1849 264
rect 1853 260 1857 264
rect 1873 260 1877 264
rect 1883 260 1887 264
rect 1905 260 1909 264
rect 1965 260 1969 264
rect 2025 260 2029 264
rect 2071 260 2075 264
rect 2091 260 2095 264
rect 2111 260 2115 264
rect 2171 260 2175 264
rect 2231 260 2235 264
rect 2251 260 2255 264
rect 2271 260 2275 264
rect 2291 260 2295 264
rect 2365 260 2369 264
rect 2385 260 2389 264
rect 2405 260 2409 264
rect 2451 260 2455 264
rect 2471 260 2475 264
rect 2535 260 2539 264
rect 2555 260 2559 264
rect 2565 260 2569 264
rect 2587 260 2591 264
rect 2597 260 2601 264
rect 2619 260 2623 264
rect 2665 260 2669 264
rect 2673 260 2677 264
rect 2693 260 2697 264
rect 2703 260 2707 264
rect 2725 260 2729 264
rect 2785 260 2789 264
rect 2805 260 2809 264
rect 2825 260 2829 264
rect 2871 260 2875 264
rect 2891 260 2895 264
rect 2955 260 2959 264
rect 2975 260 2979 264
rect 2985 260 2989 264
rect 3007 260 3011 264
rect 3017 260 3021 264
rect 3039 260 3043 264
rect 3085 260 3089 264
rect 3093 260 3097 264
rect 3113 260 3117 264
rect 3123 260 3127 264
rect 3145 260 3149 264
rect 3193 260 3197 264
rect 3203 260 3207 264
rect 3285 260 3289 264
rect 3305 260 3309 264
rect 3325 260 3329 264
rect 3371 260 3375 264
rect 3391 260 3395 264
rect 3472 260 3476 264
rect 3494 260 3498 264
rect 3502 260 3506 264
rect 3551 260 3555 264
rect 3571 260 3575 264
rect 3591 260 3595 264
rect 3651 260 3655 264
rect 3671 260 3675 264
rect 3734 260 3738 264
rect 3742 260 3746 264
rect 3764 260 3768 264
rect 3845 260 3849 264
rect 3865 260 3869 264
rect 3911 260 3915 264
rect 3931 260 3935 264
rect 3951 260 3955 264
rect 4048 260 4052 264
rect 4056 260 4060 264
rect 4064 260 4068 264
rect 4111 260 4115 264
rect 4131 260 4135 264
rect 4191 260 4195 264
rect 4213 260 4217 264
rect 4223 260 4227 264
rect 4243 260 4247 264
rect 4251 260 4255 264
rect 4297 260 4301 264
rect 4319 260 4323 264
rect 4329 260 4333 264
rect 4351 260 4355 264
rect 4361 260 4365 264
rect 4381 260 4385 264
rect 4431 260 4435 264
rect 4451 260 4455 264
rect 4525 260 4529 264
rect 4545 260 4549 264
rect 4565 260 4569 264
rect 4611 260 4615 264
rect 4631 260 4635 264
rect 4705 260 4709 264
rect 4725 260 4729 264
rect 4745 260 4749 264
rect 4765 260 4769 264
rect 4825 260 4829 264
rect 4875 260 4879 264
rect 4895 260 4899 264
rect 4905 260 4909 264
rect 4927 260 4931 264
rect 4937 260 4941 264
rect 4959 260 4963 264
rect 5005 260 5009 264
rect 5013 260 5017 264
rect 5033 260 5037 264
rect 5043 260 5047 264
rect 5065 260 5069 264
rect 5132 260 5136 264
rect 5154 260 5158 264
rect 5162 260 5166 264
rect 5211 260 5215 264
rect 5231 260 5235 264
rect 5305 260 5309 264
rect 5325 260 5329 264
rect 5345 260 5349 264
rect 5391 260 5395 264
rect 5411 260 5415 264
rect 5474 260 5478 264
rect 5482 260 5486 264
rect 5504 260 5508 264
rect 5572 260 5576 264
rect 5580 260 5584 264
rect 5588 260 5592 264
rect 5671 260 5675 264
rect 5691 260 5695 264
rect 5711 260 5715 264
rect 5793 260 5797 264
rect 5803 260 5807 264
rect 5865 260 5869 264
rect 5885 260 5889 264
rect 5905 260 5909 264
rect 5951 260 5955 264
rect 5971 260 5975 264
rect 5991 260 5995 264
rect 6051 260 6055 264
rect 6071 260 6075 264
rect 6091 260 6095 264
rect 6165 260 6169 264
rect 6185 260 6189 264
rect 6245 260 6249 264
rect 6265 260 6269 264
rect 6325 260 6329 264
rect 6345 260 6349 264
rect 6365 260 6369 264
rect 6385 260 6389 264
rect 6435 260 6439 264
rect 6455 260 6459 264
rect 6465 260 6469 264
rect 6487 260 6491 264
rect 6497 260 6501 264
rect 6519 260 6523 264
rect 6565 260 6569 264
rect 6573 260 6577 264
rect 6593 260 6597 264
rect 6603 260 6607 264
rect 6625 260 6629 264
rect 31 236 35 240
rect 53 236 57 240
rect 63 236 67 240
rect 83 236 87 240
rect 91 236 95 240
rect 137 236 141 240
rect 159 236 163 240
rect 169 236 173 240
rect 191 236 195 240
rect 201 236 205 240
rect 221 236 225 240
rect 271 236 275 240
rect 293 236 297 240
rect 303 236 307 240
rect 323 236 327 240
rect 331 236 335 240
rect 377 236 381 240
rect 399 236 403 240
rect 409 236 413 240
rect 431 236 435 240
rect 441 236 445 240
rect 461 236 465 240
rect 523 236 527 240
rect 545 236 549 240
rect 591 236 595 240
rect 613 236 617 240
rect 683 236 687 240
rect 705 236 709 240
rect 751 236 755 240
rect 773 236 777 240
rect 783 236 787 240
rect 803 236 807 240
rect 811 236 815 240
rect 857 236 861 240
rect 879 236 883 240
rect 889 236 893 240
rect 911 236 915 240
rect 921 236 925 240
rect 941 236 945 240
rect 991 236 995 240
rect 1013 236 1017 240
rect 1093 236 1097 240
rect 1103 236 1107 240
rect 1165 236 1169 240
rect 1185 236 1189 240
rect 1205 236 1209 240
rect 1255 236 1259 240
rect 1275 236 1279 240
rect 1285 236 1289 240
rect 1307 236 1311 240
rect 1317 236 1321 240
rect 1339 236 1343 240
rect 1385 236 1389 240
rect 1393 236 1397 240
rect 1413 236 1417 240
rect 1423 236 1427 240
rect 1445 236 1449 240
rect 1505 236 1509 240
rect 1553 236 1557 240
rect 1563 236 1567 240
rect 1645 236 1649 240
rect 1665 236 1669 240
rect 1685 236 1689 240
rect 1731 236 1735 240
rect 1793 236 1797 240
rect 1803 236 1807 240
rect 1873 236 1877 240
rect 1883 236 1887 240
rect 1953 236 1957 240
rect 1963 236 1967 240
rect 2045 236 2049 240
rect 2065 236 2069 240
rect 2085 236 2089 240
rect 2135 236 2139 240
rect 2155 236 2159 240
rect 2165 236 2169 240
rect 2187 236 2191 240
rect 2197 236 2201 240
rect 2219 236 2223 240
rect 2265 236 2269 240
rect 2273 236 2277 240
rect 2293 236 2297 240
rect 2303 236 2307 240
rect 2325 236 2329 240
rect 2373 236 2377 240
rect 2383 236 2387 240
rect 2473 236 2477 240
rect 2483 236 2487 240
rect 2545 236 2549 240
rect 2565 236 2569 240
rect 2585 236 2589 240
rect 2645 236 2649 240
rect 2695 236 2699 240
rect 2715 236 2719 240
rect 2725 236 2729 240
rect 2747 236 2751 240
rect 2757 236 2761 240
rect 2779 236 2783 240
rect 2825 236 2829 240
rect 2833 236 2837 240
rect 2853 236 2857 240
rect 2863 236 2867 240
rect 2885 236 2889 240
rect 2945 236 2949 240
rect 2965 236 2969 240
rect 2985 236 2989 240
rect 3045 236 3049 240
rect 3065 236 3069 240
rect 3125 236 3129 240
rect 3145 236 3149 240
rect 3165 236 3169 240
rect 3185 236 3189 240
rect 3245 236 3249 240
rect 3291 236 3295 240
rect 3313 236 3317 240
rect 3323 236 3327 240
rect 3343 236 3347 240
rect 3351 236 3355 240
rect 3397 236 3401 240
rect 3419 236 3423 240
rect 3429 236 3433 240
rect 3451 236 3455 240
rect 3461 236 3465 240
rect 3481 236 3485 240
rect 3553 236 3557 240
rect 3563 236 3567 240
rect 3625 236 3629 240
rect 3645 236 3649 240
rect 3665 236 3669 240
rect 3711 236 3715 240
rect 3731 236 3735 240
rect 3751 236 3755 240
rect 3811 236 3815 240
rect 3833 236 3837 240
rect 3843 236 3847 240
rect 3863 236 3867 240
rect 3871 236 3875 240
rect 3917 236 3921 240
rect 3939 236 3943 240
rect 3949 236 3953 240
rect 3971 236 3975 240
rect 3981 236 3985 240
rect 4001 236 4005 240
rect 4051 236 4055 240
rect 4071 236 4075 240
rect 4091 236 4095 240
rect 4151 236 4155 240
rect 4171 236 4175 240
rect 4191 236 4195 240
rect 4253 236 4257 240
rect 4263 236 4267 240
rect 4331 236 4335 240
rect 4353 236 4357 240
rect 4363 236 4367 240
rect 4383 236 4387 240
rect 4391 236 4395 240
rect 4437 236 4441 240
rect 4459 236 4463 240
rect 4469 236 4473 240
rect 4491 236 4495 240
rect 4501 236 4505 240
rect 4521 236 4525 240
rect 4571 236 4575 240
rect 4591 236 4595 240
rect 4611 236 4615 240
rect 4671 236 4675 240
rect 4691 236 4695 240
rect 4711 236 4715 240
rect 4773 236 4777 240
rect 4783 236 4787 240
rect 4851 236 4855 240
rect 4873 236 4877 240
rect 4883 236 4887 240
rect 4903 236 4907 240
rect 4911 236 4915 240
rect 4957 236 4961 240
rect 4979 236 4983 240
rect 4989 236 4993 240
rect 5011 236 5015 240
rect 5021 236 5025 240
rect 5041 236 5045 240
rect 5105 236 5109 240
rect 5125 236 5129 240
rect 5145 236 5149 240
rect 5191 236 5195 240
rect 5211 236 5215 240
rect 5231 236 5235 240
rect 5293 236 5297 240
rect 5303 236 5307 240
rect 5371 236 5375 240
rect 5393 236 5397 240
rect 5403 236 5407 240
rect 5423 236 5427 240
rect 5431 236 5435 240
rect 5477 236 5481 240
rect 5499 236 5503 240
rect 5509 236 5513 240
rect 5531 236 5535 240
rect 5541 236 5545 240
rect 5561 236 5565 240
rect 5611 236 5615 240
rect 5633 236 5637 240
rect 5643 236 5647 240
rect 5663 236 5667 240
rect 5671 236 5675 240
rect 5717 236 5721 240
rect 5739 236 5743 240
rect 5749 236 5753 240
rect 5771 236 5775 240
rect 5781 236 5785 240
rect 5801 236 5805 240
rect 5851 236 5855 240
rect 5873 236 5877 240
rect 5883 236 5887 240
rect 5903 236 5907 240
rect 5911 236 5915 240
rect 5957 236 5961 240
rect 5979 236 5983 240
rect 5989 236 5993 240
rect 6011 236 6015 240
rect 6021 236 6025 240
rect 6041 236 6045 240
rect 6105 236 6109 240
rect 6151 236 6155 240
rect 6171 236 6175 240
rect 6191 236 6195 240
rect 6265 236 6269 240
rect 6285 236 6289 240
rect 6305 236 6309 240
rect 6325 236 6329 240
rect 6385 236 6389 240
rect 6431 236 6435 240
rect 6453 236 6457 240
rect 6463 236 6467 240
rect 6483 236 6487 240
rect 6491 236 6495 240
rect 6537 236 6541 240
rect 6559 236 6563 240
rect 6569 236 6573 240
rect 6591 236 6595 240
rect 6601 236 6605 240
rect 6621 236 6625 240
rect 31 128 35 196
rect 53 167 57 216
rect 63 195 67 216
rect 83 204 87 216
rect 91 212 95 216
rect 91 208 125 212
rect 83 200 113 204
rect 83 199 101 200
rect 63 191 87 195
rect 31 116 33 128
rect 31 104 35 116
rect 53 109 57 155
rect 49 103 57 109
rect 49 74 53 103
rect 81 96 87 191
rect 49 67 57 74
rect 53 44 57 67
rect 61 44 65 84
rect 81 64 85 96
rect 121 82 125 208
rect 137 102 141 216
rect 159 204 163 216
rect 161 192 163 204
rect 169 204 173 216
rect 169 192 171 204
rect 89 70 113 72
rect 89 68 125 70
rect 89 64 93 68
rect 135 64 139 90
rect 153 82 157 192
rect 191 184 195 216
rect 162 180 195 184
rect 162 116 166 180
rect 182 131 186 160
rect 201 158 205 216
rect 221 159 225 196
rect 182 123 191 131
rect 162 104 165 116
rect 155 64 159 70
rect 167 64 171 104
rect 187 64 191 123
rect 201 64 205 146
rect 221 104 225 147
rect 271 128 275 196
rect 293 167 297 216
rect 303 195 307 216
rect 323 204 327 216
rect 331 212 335 216
rect 331 208 365 212
rect 323 200 353 204
rect 323 199 341 200
rect 303 191 327 195
rect 271 116 273 128
rect 271 104 275 116
rect 293 109 297 155
rect 289 103 297 109
rect 289 74 293 103
rect 321 96 327 191
rect 289 67 297 74
rect 293 44 297 67
rect 301 44 305 84
rect 321 64 325 96
rect 361 82 365 208
rect 377 102 381 216
rect 399 204 403 216
rect 401 192 403 204
rect 409 204 413 216
rect 409 192 411 204
rect 329 70 353 72
rect 329 68 365 70
rect 329 64 333 68
rect 375 64 379 90
rect 393 82 397 192
rect 431 184 435 216
rect 402 180 435 184
rect 402 116 406 180
rect 422 131 426 160
rect 441 158 445 216
rect 461 159 465 196
rect 523 190 527 196
rect 523 178 525 190
rect 422 123 431 131
rect 402 104 405 116
rect 395 64 399 70
rect 407 64 411 104
rect 427 64 431 123
rect 441 64 445 146
rect 461 104 465 147
rect 545 139 549 216
rect 591 139 595 216
rect 613 190 617 196
rect 615 178 617 190
rect 683 190 687 196
rect 683 178 685 190
rect 545 127 554 139
rect 586 127 595 139
rect 523 110 525 122
rect 523 104 527 110
rect 545 64 549 127
rect 591 64 595 127
rect 705 139 709 216
rect 705 127 714 139
rect 751 128 755 196
rect 773 167 777 216
rect 783 195 787 216
rect 803 204 807 216
rect 811 212 815 216
rect 811 208 845 212
rect 803 200 833 204
rect 803 199 821 200
rect 783 191 807 195
rect 615 110 617 122
rect 613 104 617 110
rect 683 110 685 122
rect 683 104 687 110
rect 705 64 709 127
rect 751 116 753 128
rect 751 104 755 116
rect 773 109 777 155
rect 769 103 777 109
rect 769 74 773 103
rect 801 96 807 191
rect 769 67 777 74
rect 773 44 777 67
rect 781 44 785 84
rect 801 64 805 96
rect 841 82 845 208
rect 857 102 861 216
rect 879 204 883 216
rect 881 192 883 204
rect 889 204 893 216
rect 889 192 891 204
rect 809 70 833 72
rect 809 68 845 70
rect 809 64 813 68
rect 855 64 859 90
rect 873 82 877 192
rect 911 184 915 216
rect 882 180 915 184
rect 882 116 886 180
rect 902 131 906 160
rect 921 158 925 216
rect 941 159 945 196
rect 902 123 911 131
rect 882 104 885 116
rect 875 64 879 70
rect 887 64 891 104
rect 907 64 911 123
rect 921 64 925 146
rect 941 104 945 147
rect 991 139 995 216
rect 1013 190 1017 196
rect 1015 178 1017 190
rect 1093 176 1097 196
rect 1083 169 1097 176
rect 1103 176 1107 196
rect 1103 169 1111 176
rect 1083 153 1089 169
rect 1086 141 1089 153
rect 986 127 995 139
rect 991 64 995 127
rect 1015 110 1017 122
rect 1013 104 1017 110
rect 1085 64 1089 141
rect 1105 153 1111 169
rect 1105 141 1114 153
rect 1105 64 1109 141
rect 1165 119 1169 196
rect 1185 173 1189 196
rect 1205 191 1209 196
rect 1205 184 1218 191
rect 1185 161 1194 173
rect 1167 107 1174 119
rect 1170 64 1174 107
rect 1192 104 1196 161
rect 1214 139 1218 184
rect 1255 159 1259 196
rect 1275 158 1279 216
rect 1285 184 1289 216
rect 1307 204 1311 216
rect 1309 192 1311 204
rect 1317 204 1321 216
rect 1317 192 1319 204
rect 1285 180 1318 184
rect 1214 116 1218 127
rect 1200 108 1218 116
rect 1200 104 1204 108
rect 1255 104 1259 147
rect 1275 64 1279 146
rect 1294 131 1298 160
rect 1289 123 1298 131
rect 1289 64 1293 123
rect 1314 116 1318 180
rect 1315 104 1318 116
rect 1309 64 1313 104
rect 1323 82 1327 192
rect 1339 102 1343 216
rect 1385 212 1389 216
rect 1355 208 1389 212
rect 1321 64 1325 70
rect 1341 64 1345 90
rect 1355 82 1359 208
rect 1393 204 1397 216
rect 1367 200 1397 204
rect 1379 199 1397 200
rect 1413 195 1417 216
rect 1393 191 1417 195
rect 1393 96 1399 191
rect 1423 167 1427 216
rect 1423 109 1427 155
rect 1445 128 1449 196
rect 1447 116 1449 128
rect 1423 103 1431 109
rect 1445 104 1449 116
rect 1505 159 1509 216
rect 1553 176 1557 196
rect 1549 169 1557 176
rect 1563 176 1567 196
rect 1563 169 1577 176
rect 1505 147 1514 159
rect 1549 153 1555 169
rect 1367 70 1391 72
rect 1355 68 1391 70
rect 1387 64 1391 68
rect 1395 64 1399 96
rect 1415 44 1419 84
rect 1427 74 1431 103
rect 1423 67 1431 74
rect 1423 44 1427 67
rect 1505 64 1509 147
rect 1546 141 1555 153
rect 1551 64 1555 141
rect 1571 153 1577 169
rect 1571 141 1574 153
rect 1571 64 1575 141
rect 1645 119 1649 196
rect 1665 173 1669 196
rect 1685 191 1689 196
rect 1685 184 1698 191
rect 1665 161 1674 173
rect 1647 107 1654 119
rect 1650 64 1654 107
rect 1672 104 1676 161
rect 1694 139 1698 184
rect 1731 159 1735 216
rect 1793 176 1797 196
rect 1726 147 1735 159
rect 1789 169 1797 176
rect 1803 176 1807 196
rect 1873 176 1877 196
rect 1803 169 1817 176
rect 1789 153 1795 169
rect 1694 116 1698 127
rect 1680 108 1698 116
rect 1680 104 1684 108
rect 1731 64 1735 147
rect 1786 141 1795 153
rect 1791 64 1795 141
rect 1811 153 1817 169
rect 1869 169 1877 176
rect 1883 176 1887 196
rect 1953 176 1957 196
rect 1883 169 1897 176
rect 1869 153 1875 169
rect 1811 141 1814 153
rect 1866 141 1875 153
rect 1811 64 1815 141
rect 1871 64 1875 141
rect 1891 153 1897 169
rect 1949 169 1957 176
rect 1963 176 1967 196
rect 1963 169 1977 176
rect 1949 153 1955 169
rect 1891 141 1894 153
rect 1946 141 1955 153
rect 1891 64 1895 141
rect 1951 64 1955 141
rect 1971 153 1977 169
rect 1971 141 1974 153
rect 1971 64 1975 141
rect 2045 119 2049 196
rect 2065 173 2069 196
rect 2085 191 2089 196
rect 2085 184 2098 191
rect 2065 161 2074 173
rect 2047 107 2054 119
rect 2050 64 2054 107
rect 2072 104 2076 161
rect 2094 139 2098 184
rect 2135 159 2139 196
rect 2155 158 2159 216
rect 2165 184 2169 216
rect 2187 204 2191 216
rect 2189 192 2191 204
rect 2197 204 2201 216
rect 2197 192 2199 204
rect 2165 180 2198 184
rect 2094 116 2098 127
rect 2080 108 2098 116
rect 2080 104 2084 108
rect 2135 104 2139 147
rect 2155 64 2159 146
rect 2174 131 2178 160
rect 2169 123 2178 131
rect 2169 64 2173 123
rect 2194 116 2198 180
rect 2195 104 2198 116
rect 2189 64 2193 104
rect 2203 82 2207 192
rect 2219 102 2223 216
rect 2265 212 2269 216
rect 2235 208 2269 212
rect 2201 64 2205 70
rect 2221 64 2225 90
rect 2235 82 2239 208
rect 2273 204 2277 216
rect 2247 200 2277 204
rect 2259 199 2277 200
rect 2293 195 2297 216
rect 2273 191 2297 195
rect 2273 96 2279 191
rect 2303 167 2307 216
rect 2303 109 2307 155
rect 2325 128 2329 196
rect 2373 176 2377 196
rect 2369 169 2377 176
rect 2383 176 2387 196
rect 2473 176 2477 196
rect 2383 169 2397 176
rect 2369 153 2375 169
rect 2366 141 2375 153
rect 2327 116 2329 128
rect 2303 103 2311 109
rect 2325 104 2329 116
rect 2247 70 2271 72
rect 2235 68 2271 70
rect 2267 64 2271 68
rect 2275 64 2279 96
rect 2295 44 2299 84
rect 2307 74 2311 103
rect 2303 67 2311 74
rect 2303 44 2307 67
rect 2371 64 2375 141
rect 2391 153 2397 169
rect 2463 169 2477 176
rect 2483 176 2487 196
rect 2483 169 2491 176
rect 2463 153 2469 169
rect 2391 141 2394 153
rect 2466 141 2469 153
rect 2391 64 2395 141
rect 2465 64 2469 141
rect 2485 153 2491 169
rect 2485 141 2494 153
rect 2485 64 2489 141
rect 2545 119 2549 196
rect 2565 173 2569 196
rect 2585 191 2589 196
rect 2585 184 2598 191
rect 2565 161 2574 173
rect 2547 107 2554 119
rect 2550 64 2554 107
rect 2572 104 2576 161
rect 2594 139 2598 184
rect 2645 159 2649 216
rect 2695 159 2699 196
rect 2645 147 2654 159
rect 2715 158 2719 216
rect 2725 184 2729 216
rect 2747 204 2751 216
rect 2749 192 2751 204
rect 2757 204 2761 216
rect 2757 192 2759 204
rect 2725 180 2758 184
rect 2594 116 2598 127
rect 2580 108 2598 116
rect 2580 104 2584 108
rect 2645 64 2649 147
rect 2695 104 2699 147
rect 2715 64 2719 146
rect 2734 131 2738 160
rect 2729 123 2738 131
rect 2729 64 2733 123
rect 2754 116 2758 180
rect 2755 104 2758 116
rect 2749 64 2753 104
rect 2763 82 2767 192
rect 2779 102 2783 216
rect 2825 212 2829 216
rect 2795 208 2829 212
rect 2761 64 2765 70
rect 2781 64 2785 90
rect 2795 82 2799 208
rect 2833 204 2837 216
rect 2807 200 2837 204
rect 2819 199 2837 200
rect 2853 195 2857 216
rect 2833 191 2857 195
rect 2833 96 2839 191
rect 2863 167 2867 216
rect 2863 109 2867 155
rect 2885 128 2889 196
rect 2887 116 2889 128
rect 2945 119 2949 196
rect 2965 173 2969 196
rect 2985 191 2989 196
rect 2985 184 2998 191
rect 2965 161 2974 173
rect 2863 103 2871 109
rect 2885 104 2889 116
rect 2947 107 2954 119
rect 2807 70 2831 72
rect 2795 68 2831 70
rect 2827 64 2831 68
rect 2835 64 2839 96
rect 2855 44 2859 84
rect 2867 74 2871 103
rect 2863 67 2871 74
rect 2863 44 2867 67
rect 2950 64 2954 107
rect 2972 104 2976 161
rect 2994 139 2998 184
rect 3045 139 3049 216
rect 3065 139 3069 216
rect 3125 139 3129 196
rect 3145 173 3149 196
rect 3165 173 3169 196
rect 3185 189 3189 196
rect 3185 185 3200 189
rect 3165 161 3174 173
rect 3046 127 3061 139
rect 2994 116 2998 127
rect 2980 108 2998 116
rect 2980 104 2984 108
rect 3057 104 3061 127
rect 3065 127 3074 139
rect 3127 127 3129 139
rect 3065 104 3069 127
rect 3125 112 3129 127
rect 3125 108 3139 112
rect 3135 104 3139 108
rect 3145 104 3149 161
rect 3165 112 3171 161
rect 3194 139 3200 185
rect 3245 159 3249 216
rect 3245 147 3254 159
rect 3194 112 3199 127
rect 3165 108 3179 112
rect 3175 104 3179 108
rect 3185 108 3199 112
rect 3185 104 3189 108
rect 3245 64 3249 147
rect 3291 128 3295 196
rect 3313 167 3317 216
rect 3323 195 3327 216
rect 3343 204 3347 216
rect 3351 212 3355 216
rect 3351 208 3385 212
rect 3343 200 3373 204
rect 3343 199 3361 200
rect 3323 191 3347 195
rect 3291 116 3293 128
rect 3291 104 3295 116
rect 3313 109 3317 155
rect 3309 103 3317 109
rect 3309 74 3313 103
rect 3341 96 3347 191
rect 3309 67 3317 74
rect 3313 44 3317 67
rect 3321 44 3325 84
rect 3341 64 3345 96
rect 3381 82 3385 208
rect 3397 102 3401 216
rect 3419 204 3423 216
rect 3421 192 3423 204
rect 3429 204 3433 216
rect 3429 192 3431 204
rect 3349 70 3373 72
rect 3349 68 3385 70
rect 3349 64 3353 68
rect 3395 64 3399 90
rect 3413 82 3417 192
rect 3451 184 3455 216
rect 3422 180 3455 184
rect 3422 116 3426 180
rect 3442 131 3446 160
rect 3461 158 3465 216
rect 3481 159 3485 196
rect 3553 176 3557 196
rect 3543 169 3557 176
rect 3563 176 3567 196
rect 3563 169 3571 176
rect 3543 153 3549 169
rect 3442 123 3451 131
rect 3422 104 3425 116
rect 3415 64 3419 70
rect 3427 64 3431 104
rect 3447 64 3451 123
rect 3461 64 3465 146
rect 3481 104 3485 147
rect 3546 141 3549 153
rect 3545 64 3549 141
rect 3565 153 3571 169
rect 3565 141 3574 153
rect 3565 64 3569 141
rect 3625 119 3629 196
rect 3645 173 3649 196
rect 3665 191 3669 196
rect 3711 191 3715 196
rect 3665 184 3678 191
rect 3645 161 3654 173
rect 3627 107 3634 119
rect 3630 64 3634 107
rect 3652 104 3656 161
rect 3674 139 3678 184
rect 3702 184 3715 191
rect 3702 139 3706 184
rect 3731 173 3735 196
rect 3726 161 3735 173
rect 3674 116 3678 127
rect 3660 108 3678 116
rect 3702 116 3706 127
rect 3702 108 3720 116
rect 3660 104 3664 108
rect 3716 104 3720 108
rect 3724 104 3728 161
rect 3751 119 3755 196
rect 3811 128 3815 196
rect 3833 167 3837 216
rect 3843 195 3847 216
rect 3863 204 3867 216
rect 3871 212 3875 216
rect 3871 208 3905 212
rect 3863 200 3893 204
rect 3863 199 3881 200
rect 3843 191 3867 195
rect 3746 107 3753 119
rect 3811 116 3813 128
rect 3746 64 3750 107
rect 3811 104 3815 116
rect 3833 109 3837 155
rect 3829 103 3837 109
rect 3829 74 3833 103
rect 3861 96 3867 191
rect 3829 67 3837 74
rect 3833 44 3837 67
rect 3841 44 3845 84
rect 3861 64 3865 96
rect 3901 82 3905 208
rect 3917 102 3921 216
rect 3939 204 3943 216
rect 3941 192 3943 204
rect 3949 204 3953 216
rect 3949 192 3951 204
rect 3869 70 3893 72
rect 3869 68 3905 70
rect 3869 64 3873 68
rect 3915 64 3919 90
rect 3933 82 3937 192
rect 3971 184 3975 216
rect 3942 180 3975 184
rect 3942 116 3946 180
rect 3962 131 3966 160
rect 3981 158 3985 216
rect 4001 159 4005 196
rect 4051 191 4055 196
rect 4042 184 4055 191
rect 3962 123 3971 131
rect 3942 104 3945 116
rect 3935 64 3939 70
rect 3947 64 3951 104
rect 3967 64 3971 123
rect 3981 64 3985 146
rect 4001 104 4005 147
rect 4042 139 4046 184
rect 4071 173 4075 196
rect 4066 161 4075 173
rect 4042 116 4046 127
rect 4042 108 4060 116
rect 4056 104 4060 108
rect 4064 104 4068 161
rect 4091 119 4095 196
rect 4151 191 4155 196
rect 4142 184 4155 191
rect 4142 139 4146 184
rect 4171 173 4175 196
rect 4166 161 4175 173
rect 4086 107 4093 119
rect 4142 116 4146 127
rect 4142 108 4160 116
rect 4086 64 4090 107
rect 4156 104 4160 108
rect 4164 104 4168 161
rect 4191 119 4195 196
rect 4253 176 4257 196
rect 4249 169 4257 176
rect 4263 176 4267 196
rect 4263 169 4277 176
rect 4249 153 4255 169
rect 4246 141 4255 153
rect 4186 107 4193 119
rect 4186 64 4190 107
rect 4251 64 4255 141
rect 4271 153 4277 169
rect 4271 141 4274 153
rect 4271 64 4275 141
rect 4331 128 4335 196
rect 4353 167 4357 216
rect 4363 195 4367 216
rect 4383 204 4387 216
rect 4391 212 4395 216
rect 4391 208 4425 212
rect 4383 200 4413 204
rect 4383 199 4401 200
rect 4363 191 4387 195
rect 4331 116 4333 128
rect 4331 104 4335 116
rect 4353 109 4357 155
rect 4349 103 4357 109
rect 4349 74 4353 103
rect 4381 96 4387 191
rect 4349 67 4357 74
rect 4353 44 4357 67
rect 4361 44 4365 84
rect 4381 64 4385 96
rect 4421 82 4425 208
rect 4437 102 4441 216
rect 4459 204 4463 216
rect 4461 192 4463 204
rect 4469 204 4473 216
rect 4469 192 4471 204
rect 4389 70 4413 72
rect 4389 68 4425 70
rect 4389 64 4393 68
rect 4435 64 4439 90
rect 4453 82 4457 192
rect 4491 184 4495 216
rect 4462 180 4495 184
rect 4462 116 4466 180
rect 4482 131 4486 160
rect 4501 158 4505 216
rect 4521 159 4525 196
rect 4571 191 4575 196
rect 4562 184 4575 191
rect 4482 123 4491 131
rect 4462 104 4465 116
rect 4455 64 4459 70
rect 4467 64 4471 104
rect 4487 64 4491 123
rect 4501 64 4505 146
rect 4521 104 4525 147
rect 4562 139 4566 184
rect 4591 173 4595 196
rect 4586 161 4595 173
rect 4562 116 4566 127
rect 4562 108 4580 116
rect 4576 104 4580 108
rect 4584 104 4588 161
rect 4611 119 4615 196
rect 4671 191 4675 196
rect 4662 184 4675 191
rect 4662 139 4666 184
rect 4691 173 4695 196
rect 4686 161 4695 173
rect 4606 107 4613 119
rect 4662 116 4666 127
rect 4662 108 4680 116
rect 4606 64 4610 107
rect 4676 104 4680 108
rect 4684 104 4688 161
rect 4711 119 4715 196
rect 4773 176 4777 196
rect 4769 169 4777 176
rect 4783 176 4787 196
rect 4783 169 4797 176
rect 4769 153 4775 169
rect 4766 141 4775 153
rect 4706 107 4713 119
rect 4706 64 4710 107
rect 4771 64 4775 141
rect 4791 153 4797 169
rect 4791 141 4794 153
rect 4791 64 4795 141
rect 4851 128 4855 196
rect 4873 167 4877 216
rect 4883 195 4887 216
rect 4903 204 4907 216
rect 4911 212 4915 216
rect 4911 208 4945 212
rect 4903 200 4933 204
rect 4903 199 4921 200
rect 4883 191 4907 195
rect 4851 116 4853 128
rect 4851 104 4855 116
rect 4873 109 4877 155
rect 4869 103 4877 109
rect 4869 74 4873 103
rect 4901 96 4907 191
rect 4869 67 4877 74
rect 4873 44 4877 67
rect 4881 44 4885 84
rect 4901 64 4905 96
rect 4941 82 4945 208
rect 4957 102 4961 216
rect 4979 204 4983 216
rect 4981 192 4983 204
rect 4989 204 4993 216
rect 4989 192 4991 204
rect 4909 70 4933 72
rect 4909 68 4945 70
rect 4909 64 4913 68
rect 4955 64 4959 90
rect 4973 82 4977 192
rect 5011 184 5015 216
rect 4982 180 5015 184
rect 4982 116 4986 180
rect 5002 131 5006 160
rect 5021 158 5025 216
rect 5041 159 5045 196
rect 5002 123 5011 131
rect 4982 104 4985 116
rect 4975 64 4979 70
rect 4987 64 4991 104
rect 5007 64 5011 123
rect 5021 64 5025 146
rect 5041 104 5045 147
rect 5105 119 5109 196
rect 5125 173 5129 196
rect 5145 191 5149 196
rect 5191 191 5195 196
rect 5145 184 5158 191
rect 5125 161 5134 173
rect 5107 107 5114 119
rect 5110 64 5114 107
rect 5132 104 5136 161
rect 5154 139 5158 184
rect 5182 184 5195 191
rect 5182 139 5186 184
rect 5211 173 5215 196
rect 5206 161 5215 173
rect 5154 116 5158 127
rect 5140 108 5158 116
rect 5182 116 5186 127
rect 5182 108 5200 116
rect 5140 104 5144 108
rect 5196 104 5200 108
rect 5204 104 5208 161
rect 5231 119 5235 196
rect 5293 176 5297 196
rect 5289 169 5297 176
rect 5303 176 5307 196
rect 5303 169 5317 176
rect 5289 153 5295 169
rect 5286 141 5295 153
rect 5226 107 5233 119
rect 5226 64 5230 107
rect 5291 64 5295 141
rect 5311 153 5317 169
rect 5311 141 5314 153
rect 5311 64 5315 141
rect 5371 128 5375 196
rect 5393 167 5397 216
rect 5403 195 5407 216
rect 5423 204 5427 216
rect 5431 212 5435 216
rect 5431 208 5465 212
rect 5423 200 5453 204
rect 5423 199 5441 200
rect 5403 191 5427 195
rect 5371 116 5373 128
rect 5371 104 5375 116
rect 5393 109 5397 155
rect 5389 103 5397 109
rect 5389 74 5393 103
rect 5421 96 5427 191
rect 5389 67 5397 74
rect 5393 44 5397 67
rect 5401 44 5405 84
rect 5421 64 5425 96
rect 5461 82 5465 208
rect 5477 102 5481 216
rect 5499 204 5503 216
rect 5501 192 5503 204
rect 5509 204 5513 216
rect 5509 192 5511 204
rect 5429 70 5453 72
rect 5429 68 5465 70
rect 5429 64 5433 68
rect 5475 64 5479 90
rect 5493 82 5497 192
rect 5531 184 5535 216
rect 5502 180 5535 184
rect 5502 116 5506 180
rect 5522 131 5526 160
rect 5541 158 5545 216
rect 5561 159 5565 196
rect 5522 123 5531 131
rect 5502 104 5505 116
rect 5495 64 5499 70
rect 5507 64 5511 104
rect 5527 64 5531 123
rect 5541 64 5545 146
rect 5561 104 5565 147
rect 5611 128 5615 196
rect 5633 167 5637 216
rect 5643 195 5647 216
rect 5663 204 5667 216
rect 5671 212 5675 216
rect 5671 208 5705 212
rect 5663 200 5693 204
rect 5663 199 5681 200
rect 5643 191 5667 195
rect 5611 116 5613 128
rect 5611 104 5615 116
rect 5633 109 5637 155
rect 5629 103 5637 109
rect 5629 74 5633 103
rect 5661 96 5667 191
rect 5629 67 5637 74
rect 5633 44 5637 67
rect 5641 44 5645 84
rect 5661 64 5665 96
rect 5701 82 5705 208
rect 5717 102 5721 216
rect 5739 204 5743 216
rect 5741 192 5743 204
rect 5749 204 5753 216
rect 5749 192 5751 204
rect 5669 70 5693 72
rect 5669 68 5705 70
rect 5669 64 5673 68
rect 5715 64 5719 90
rect 5733 82 5737 192
rect 5771 184 5775 216
rect 5742 180 5775 184
rect 5742 116 5746 180
rect 5762 131 5766 160
rect 5781 158 5785 216
rect 5801 159 5805 196
rect 5762 123 5771 131
rect 5742 104 5745 116
rect 5735 64 5739 70
rect 5747 64 5751 104
rect 5767 64 5771 123
rect 5781 64 5785 146
rect 5801 104 5805 147
rect 5851 128 5855 196
rect 5873 167 5877 216
rect 5883 195 5887 216
rect 5903 204 5907 216
rect 5911 212 5915 216
rect 5911 208 5945 212
rect 5903 200 5933 204
rect 5903 199 5921 200
rect 5883 191 5907 195
rect 5851 116 5853 128
rect 5851 104 5855 116
rect 5873 109 5877 155
rect 5869 103 5877 109
rect 5869 74 5873 103
rect 5901 96 5907 191
rect 5869 67 5877 74
rect 5873 44 5877 67
rect 5881 44 5885 84
rect 5901 64 5905 96
rect 5941 82 5945 208
rect 5957 102 5961 216
rect 5979 204 5983 216
rect 5981 192 5983 204
rect 5989 204 5993 216
rect 5989 192 5991 204
rect 5909 70 5933 72
rect 5909 68 5945 70
rect 5909 64 5913 68
rect 5955 64 5959 90
rect 5973 82 5977 192
rect 6011 184 6015 216
rect 5982 180 6015 184
rect 5982 116 5986 180
rect 6002 131 6006 160
rect 6021 158 6025 216
rect 6041 159 6045 196
rect 6105 173 6109 196
rect 6151 191 6155 196
rect 6142 184 6155 191
rect 6105 161 6114 173
rect 6002 123 6011 131
rect 5982 104 5985 116
rect 5975 64 5979 70
rect 5987 64 5991 104
rect 6007 64 6011 123
rect 6021 64 6025 146
rect 6041 104 6045 147
rect 6105 104 6109 161
rect 6142 139 6146 184
rect 6171 173 6175 196
rect 6166 161 6175 173
rect 6142 116 6146 127
rect 6142 108 6160 116
rect 6156 104 6160 108
rect 6164 104 6168 161
rect 6191 119 6195 196
rect 6265 139 6269 196
rect 6285 173 6289 196
rect 6305 173 6309 196
rect 6325 189 6329 196
rect 6325 185 6340 189
rect 6305 161 6314 173
rect 6267 127 6269 139
rect 6186 107 6193 119
rect 6265 112 6269 127
rect 6265 108 6279 112
rect 6186 64 6190 107
rect 6275 104 6279 108
rect 6285 104 6289 161
rect 6305 112 6311 161
rect 6334 139 6340 185
rect 6385 159 6389 216
rect 6385 147 6394 159
rect 6334 112 6339 127
rect 6305 108 6319 112
rect 6315 104 6319 108
rect 6325 108 6339 112
rect 6325 104 6329 108
rect 6385 64 6389 147
rect 6431 128 6435 196
rect 6453 167 6457 216
rect 6463 195 6467 216
rect 6483 204 6487 216
rect 6491 212 6495 216
rect 6491 208 6525 212
rect 6483 200 6513 204
rect 6483 199 6501 200
rect 6463 191 6487 195
rect 6431 116 6433 128
rect 6431 104 6435 116
rect 6453 109 6457 155
rect 6449 103 6457 109
rect 6449 74 6453 103
rect 6481 96 6487 191
rect 6449 67 6457 74
rect 6453 44 6457 67
rect 6461 44 6465 84
rect 6481 64 6485 96
rect 6521 82 6525 208
rect 6537 102 6541 216
rect 6559 204 6563 216
rect 6561 192 6563 204
rect 6569 204 6573 216
rect 6569 192 6571 204
rect 6489 70 6513 72
rect 6489 68 6525 70
rect 6489 64 6493 68
rect 6535 64 6539 90
rect 6553 82 6557 192
rect 6591 184 6595 216
rect 6562 180 6595 184
rect 6562 116 6566 180
rect 6582 131 6586 160
rect 6601 158 6605 216
rect 6621 159 6625 196
rect 6582 123 6591 131
rect 6562 104 6565 116
rect 6555 64 6559 70
rect 6567 64 6571 104
rect 6587 64 6591 123
rect 6601 64 6605 146
rect 6621 104 6625 147
rect 31 20 35 24
rect 53 20 57 24
rect 61 20 65 24
rect 81 20 85 24
rect 89 20 93 24
rect 135 20 139 24
rect 155 20 159 24
rect 167 20 171 24
rect 187 20 191 24
rect 201 20 205 24
rect 221 20 225 24
rect 271 20 275 24
rect 293 20 297 24
rect 301 20 305 24
rect 321 20 325 24
rect 329 20 333 24
rect 375 20 379 24
rect 395 20 399 24
rect 407 20 411 24
rect 427 20 431 24
rect 441 20 445 24
rect 461 20 465 24
rect 523 20 527 24
rect 545 20 549 24
rect 591 20 595 24
rect 613 20 617 24
rect 683 20 687 24
rect 705 20 709 24
rect 751 20 755 24
rect 773 20 777 24
rect 781 20 785 24
rect 801 20 805 24
rect 809 20 813 24
rect 855 20 859 24
rect 875 20 879 24
rect 887 20 891 24
rect 907 20 911 24
rect 921 20 925 24
rect 941 20 945 24
rect 991 20 995 24
rect 1013 20 1017 24
rect 1085 20 1089 24
rect 1105 20 1109 24
rect 1170 20 1174 24
rect 1192 20 1196 24
rect 1200 20 1204 24
rect 1255 20 1259 24
rect 1275 20 1279 24
rect 1289 20 1293 24
rect 1309 20 1313 24
rect 1321 20 1325 24
rect 1341 20 1345 24
rect 1387 20 1391 24
rect 1395 20 1399 24
rect 1415 20 1419 24
rect 1423 20 1427 24
rect 1445 20 1449 24
rect 1505 20 1509 24
rect 1551 20 1555 24
rect 1571 20 1575 24
rect 1650 20 1654 24
rect 1672 20 1676 24
rect 1680 20 1684 24
rect 1731 20 1735 24
rect 1791 20 1795 24
rect 1811 20 1815 24
rect 1871 20 1875 24
rect 1891 20 1895 24
rect 1951 20 1955 24
rect 1971 20 1975 24
rect 2050 20 2054 24
rect 2072 20 2076 24
rect 2080 20 2084 24
rect 2135 20 2139 24
rect 2155 20 2159 24
rect 2169 20 2173 24
rect 2189 20 2193 24
rect 2201 20 2205 24
rect 2221 20 2225 24
rect 2267 20 2271 24
rect 2275 20 2279 24
rect 2295 20 2299 24
rect 2303 20 2307 24
rect 2325 20 2329 24
rect 2371 20 2375 24
rect 2391 20 2395 24
rect 2465 20 2469 24
rect 2485 20 2489 24
rect 2550 20 2554 24
rect 2572 20 2576 24
rect 2580 20 2584 24
rect 2645 20 2649 24
rect 2695 20 2699 24
rect 2715 20 2719 24
rect 2729 20 2733 24
rect 2749 20 2753 24
rect 2761 20 2765 24
rect 2781 20 2785 24
rect 2827 20 2831 24
rect 2835 20 2839 24
rect 2855 20 2859 24
rect 2863 20 2867 24
rect 2885 20 2889 24
rect 2950 20 2954 24
rect 2972 20 2976 24
rect 2980 20 2984 24
rect 3057 20 3061 24
rect 3065 20 3069 24
rect 3135 20 3139 24
rect 3145 20 3149 24
rect 3175 20 3179 24
rect 3185 20 3189 24
rect 3245 20 3249 24
rect 3291 20 3295 24
rect 3313 20 3317 24
rect 3321 20 3325 24
rect 3341 20 3345 24
rect 3349 20 3353 24
rect 3395 20 3399 24
rect 3415 20 3419 24
rect 3427 20 3431 24
rect 3447 20 3451 24
rect 3461 20 3465 24
rect 3481 20 3485 24
rect 3545 20 3549 24
rect 3565 20 3569 24
rect 3630 20 3634 24
rect 3652 20 3656 24
rect 3660 20 3664 24
rect 3716 20 3720 24
rect 3724 20 3728 24
rect 3746 20 3750 24
rect 3811 20 3815 24
rect 3833 20 3837 24
rect 3841 20 3845 24
rect 3861 20 3865 24
rect 3869 20 3873 24
rect 3915 20 3919 24
rect 3935 20 3939 24
rect 3947 20 3951 24
rect 3967 20 3971 24
rect 3981 20 3985 24
rect 4001 20 4005 24
rect 4056 20 4060 24
rect 4064 20 4068 24
rect 4086 20 4090 24
rect 4156 20 4160 24
rect 4164 20 4168 24
rect 4186 20 4190 24
rect 4251 20 4255 24
rect 4271 20 4275 24
rect 4331 20 4335 24
rect 4353 20 4357 24
rect 4361 20 4365 24
rect 4381 20 4385 24
rect 4389 20 4393 24
rect 4435 20 4439 24
rect 4455 20 4459 24
rect 4467 20 4471 24
rect 4487 20 4491 24
rect 4501 20 4505 24
rect 4521 20 4525 24
rect 4576 20 4580 24
rect 4584 20 4588 24
rect 4606 20 4610 24
rect 4676 20 4680 24
rect 4684 20 4688 24
rect 4706 20 4710 24
rect 4771 20 4775 24
rect 4791 20 4795 24
rect 4851 20 4855 24
rect 4873 20 4877 24
rect 4881 20 4885 24
rect 4901 20 4905 24
rect 4909 20 4913 24
rect 4955 20 4959 24
rect 4975 20 4979 24
rect 4987 20 4991 24
rect 5007 20 5011 24
rect 5021 20 5025 24
rect 5041 20 5045 24
rect 5110 20 5114 24
rect 5132 20 5136 24
rect 5140 20 5144 24
rect 5196 20 5200 24
rect 5204 20 5208 24
rect 5226 20 5230 24
rect 5291 20 5295 24
rect 5311 20 5315 24
rect 5371 20 5375 24
rect 5393 20 5397 24
rect 5401 20 5405 24
rect 5421 20 5425 24
rect 5429 20 5433 24
rect 5475 20 5479 24
rect 5495 20 5499 24
rect 5507 20 5511 24
rect 5527 20 5531 24
rect 5541 20 5545 24
rect 5561 20 5565 24
rect 5611 20 5615 24
rect 5633 20 5637 24
rect 5641 20 5645 24
rect 5661 20 5665 24
rect 5669 20 5673 24
rect 5715 20 5719 24
rect 5735 20 5739 24
rect 5747 20 5751 24
rect 5767 20 5771 24
rect 5781 20 5785 24
rect 5801 20 5805 24
rect 5851 20 5855 24
rect 5873 20 5877 24
rect 5881 20 5885 24
rect 5901 20 5905 24
rect 5909 20 5913 24
rect 5955 20 5959 24
rect 5975 20 5979 24
rect 5987 20 5991 24
rect 6007 20 6011 24
rect 6021 20 6025 24
rect 6041 20 6045 24
rect 6105 20 6109 24
rect 6156 20 6160 24
rect 6164 20 6168 24
rect 6186 20 6190 24
rect 6275 20 6279 24
rect 6285 20 6289 24
rect 6315 20 6319 24
rect 6325 20 6329 24
rect 6385 20 6389 24
rect 6431 20 6435 24
rect 6453 20 6457 24
rect 6461 20 6465 24
rect 6481 20 6485 24
rect 6489 20 6493 24
rect 6535 20 6539 24
rect 6555 20 6559 24
rect 6567 20 6571 24
rect 6587 20 6591 24
rect 6601 20 6605 24
rect 6621 20 6625 24
<< polycontact >>
rect 34 6387 46 6399
rect 77 6432 89 6444
rect 99 6432 111 6444
rect 74 6400 86 6412
rect 54 6386 66 6398
rect 83 6344 95 6356
rect 115 6330 127 6342
rect 101 6310 113 6322
rect 147 6428 159 6440
rect 201 6395 213 6407
rect 215 6356 227 6368
rect 314 6401 326 6413
rect 275 6347 287 6359
rect 163 6324 175 6336
rect 135 6310 147 6322
rect 187 6324 199 6336
rect 354 6381 366 6393
rect 334 6367 346 6379
rect 394 6381 406 6393
rect 454 6381 466 6393
rect 494 6381 506 6393
rect 514 6381 526 6393
rect 554 6381 566 6393
rect 627 6395 639 6407
rect 613 6356 625 6368
rect 681 6428 693 6440
rect 641 6324 653 6336
rect 665 6324 677 6336
rect 729 6432 741 6444
rect 751 6432 763 6444
rect 713 6330 725 6342
rect 693 6310 705 6322
rect 754 6400 766 6412
rect 774 6386 786 6398
rect 794 6387 806 6399
rect 834 6387 846 6399
rect 745 6344 757 6356
rect 727 6310 739 6322
rect 915 6401 927 6413
rect 953 6401 965 6413
rect 895 6367 907 6379
rect 1054 6387 1066 6399
rect 974 6367 986 6379
rect 1107 6395 1119 6407
rect 1093 6356 1105 6368
rect 1161 6428 1173 6440
rect 1121 6324 1133 6336
rect 1145 6324 1157 6336
rect 1209 6432 1221 6444
rect 1231 6432 1243 6444
rect 1193 6330 1205 6342
rect 1173 6310 1185 6322
rect 1234 6400 1246 6412
rect 1254 6386 1266 6398
rect 1274 6387 1286 6399
rect 1225 6344 1237 6356
rect 1207 6310 1219 6322
rect 1334 6401 1346 6413
rect 1370 6401 1382 6413
rect 1314 6367 1326 6379
rect 1393 6367 1405 6379
rect 1494 6401 1506 6413
rect 1455 6347 1467 6359
rect 1573 6418 1585 6430
rect 1514 6367 1526 6379
rect 1574 6381 1586 6393
rect 1674 6387 1686 6399
rect 1614 6367 1626 6379
rect 1727 6395 1739 6407
rect 1713 6356 1725 6368
rect 1781 6428 1793 6440
rect 1741 6324 1753 6336
rect 1765 6324 1777 6336
rect 1829 6432 1841 6444
rect 1851 6432 1863 6444
rect 1813 6330 1825 6342
rect 1793 6310 1805 6322
rect 1854 6400 1866 6412
rect 1874 6386 1886 6398
rect 1894 6387 1906 6399
rect 1845 6344 1857 6356
rect 1827 6310 1839 6322
rect 1954 6401 1966 6413
rect 1934 6367 1946 6379
rect 2034 6381 2046 6393
rect 1993 6347 2005 6359
rect 2074 6381 2086 6393
rect 2174 6401 2186 6413
rect 2135 6347 2147 6359
rect 2254 6401 2266 6413
rect 2194 6367 2206 6379
rect 2294 6401 2306 6413
rect 2274 6387 2286 6399
rect 2334 6381 2346 6393
rect 2374 6381 2386 6393
rect 2554 6381 2566 6393
rect 2414 6367 2426 6379
rect 2454 6367 2466 6379
rect 2474 6367 2486 6379
rect 2514 6367 2526 6379
rect 2594 6381 2606 6393
rect 2673 6347 2685 6359
rect 2734 6381 2746 6393
rect 2714 6347 2726 6359
rect 2694 6327 2706 6339
rect 2774 6381 2786 6393
rect 2853 6347 2865 6359
rect 2974 6401 2986 6413
rect 2894 6347 2906 6359
rect 2935 6347 2947 6359
rect 2874 6327 2886 6339
rect 2994 6367 3006 6379
rect 3074 6401 3086 6413
rect 3035 6347 3047 6359
rect 3234 6401 3246 6413
rect 3154 6387 3166 6399
rect 3214 6387 3226 6399
rect 3094 6367 3106 6379
rect 3274 6401 3286 6413
rect 3254 6387 3266 6399
rect 3354 6401 3366 6413
rect 3334 6367 3346 6379
rect 3474 6401 3486 6413
rect 3393 6347 3405 6359
rect 3514 6401 3526 6413
rect 3574 6401 3586 6413
rect 3494 6387 3506 6399
rect 3614 6401 3626 6413
rect 3594 6387 3606 6399
rect 3634 6347 3646 6359
rect 3794 6401 3806 6413
rect 3675 6347 3687 6359
rect 3755 6347 3767 6359
rect 3654 6327 3666 6339
rect 3854 6401 3866 6413
rect 3814 6367 3826 6379
rect 3834 6367 3846 6379
rect 3934 6387 3946 6399
rect 4113 6418 4125 6430
rect 3893 6347 3905 6359
rect 3994 6381 4006 6393
rect 4034 6381 4046 6393
rect 4114 6381 4126 6393
rect 4174 6381 4186 6393
rect 4154 6367 4166 6379
rect 4214 6381 4226 6393
rect 4293 6347 4305 6359
rect 4334 6347 4346 6359
rect 4393 6347 4405 6359
rect 4314 6327 4326 6339
rect 4434 6347 4446 6359
rect 4493 6347 4505 6359
rect 4414 6327 4426 6339
rect 4614 6401 4626 6413
rect 4554 6387 4566 6399
rect 4534 6347 4546 6359
rect 4514 6327 4526 6339
rect 4654 6401 4666 6413
rect 4714 6401 4726 6413
rect 4634 6387 4646 6399
rect 4754 6401 4766 6413
rect 4734 6387 4746 6399
rect 4834 6401 4846 6413
rect 4814 6367 4826 6379
rect 4974 6401 4986 6413
rect 4873 6347 4885 6359
rect 4935 6347 4947 6359
rect 5034 6401 5046 6413
rect 4994 6367 5006 6379
rect 5014 6367 5026 6379
rect 5073 6347 5085 6359
rect 5153 6347 5165 6359
rect 5194 6347 5206 6359
rect 5253 6347 5265 6359
rect 5174 6327 5186 6339
rect 5294 6347 5306 6359
rect 5353 6347 5365 6359
rect 5274 6327 5286 6339
rect 5414 6401 5426 6413
rect 5454 6401 5466 6413
rect 5434 6387 5446 6399
rect 5394 6347 5406 6359
rect 5374 6327 5386 6339
rect 5554 6401 5566 6413
rect 5594 6401 5606 6413
rect 5574 6387 5586 6399
rect 5674 6401 5686 6413
rect 5654 6387 5666 6399
rect 5714 6401 5726 6413
rect 5694 6387 5706 6399
rect 5774 6347 5786 6359
rect 5914 6401 5926 6413
rect 5815 6347 5827 6359
rect 5794 6327 5806 6339
rect 5954 6401 5966 6413
rect 5934 6387 5946 6399
rect 6074 6401 6086 6413
rect 6014 6387 6026 6399
rect 6114 6401 6126 6413
rect 6094 6387 6106 6399
rect 6194 6401 6206 6413
rect 6155 6347 6167 6359
rect 6274 6401 6286 6413
rect 6214 6367 6226 6379
rect 6314 6401 6326 6413
rect 6294 6387 6306 6399
rect 6334 6347 6346 6359
rect 6375 6347 6387 6359
rect 6354 6327 6366 6339
rect 6473 6347 6485 6359
rect 6534 6387 6546 6399
rect 6514 6347 6526 6359
rect 6494 6327 6506 6339
rect 6615 6401 6627 6413
rect 6653 6401 6665 6413
rect 6595 6367 6607 6379
rect 6674 6367 6686 6379
rect 61 6164 73 6176
rect 113 6178 125 6190
rect 85 6164 97 6176
rect 33 6132 45 6144
rect 47 6093 59 6105
rect 101 6060 113 6072
rect 147 6178 159 6190
rect 133 6158 145 6170
rect 165 6144 177 6156
rect 194 6102 206 6114
rect 174 6088 186 6100
rect 149 6056 161 6068
rect 171 6056 183 6068
rect 214 6101 226 6113
rect 314 6101 326 6113
rect 294 6087 306 6099
rect 374 6107 386 6119
rect 334 6087 346 6099
rect 434 6121 446 6133
rect 474 6121 486 6133
rect 414 6107 426 6119
rect 534 6107 546 6119
rect 594 6121 606 6133
rect 574 6107 586 6119
rect 653 6141 665 6153
rect 715 6141 727 6153
rect 614 6087 626 6099
rect 774 6121 786 6133
rect 794 6121 806 6133
rect 834 6121 846 6133
rect 754 6087 766 6099
rect 934 6101 946 6113
rect 914 6087 926 6099
rect 1013 6139 1025 6151
rect 994 6121 1006 6133
rect 974 6101 986 6113
rect 954 6087 966 6099
rect 1134 6121 1146 6133
rect 1235 6141 1247 6153
rect 1174 6121 1186 6133
rect 1114 6101 1126 6113
rect 1013 6072 1025 6084
rect 1294 6121 1306 6133
rect 1274 6087 1286 6099
rect 1434 6121 1446 6133
rect 1474 6121 1486 6133
rect 1514 6121 1526 6133
rect 1554 6121 1566 6133
rect 1354 6101 1366 6113
rect 1414 6101 1426 6113
rect 1654 6121 1666 6133
rect 1694 6121 1706 6133
rect 1734 6121 1746 6133
rect 1774 6121 1786 6133
rect 1814 6121 1826 6133
rect 1594 6101 1606 6113
rect 1873 6141 1885 6153
rect 1834 6087 1846 6099
rect 1914 6101 1926 6113
rect 2034 6101 2046 6113
rect 2014 6087 2026 6099
rect 2155 6141 2167 6153
rect 2074 6101 2086 6113
rect 2054 6087 2066 6099
rect 2214 6121 2226 6133
rect 2194 6087 2206 6099
rect 2315 6141 2327 6153
rect 2234 6101 2246 6113
rect 2454 6161 2466 6173
rect 2433 6141 2445 6153
rect 2374 6121 2386 6133
rect 2354 6087 2366 6099
rect 2474 6141 2486 6153
rect 2554 6101 2566 6113
rect 2534 6087 2546 6099
rect 2614 6121 2626 6133
rect 2734 6161 2746 6173
rect 2713 6141 2725 6153
rect 2654 6121 2666 6133
rect 2574 6087 2586 6099
rect 2754 6141 2766 6153
rect 2794 6121 2806 6133
rect 2873 6121 2885 6133
rect 2815 6087 2827 6099
rect 2853 6087 2865 6099
rect 2974 6161 2986 6173
rect 2954 6141 2966 6153
rect 2934 6101 2946 6113
rect 2995 6141 3007 6153
rect 3214 6161 3226 6173
rect 3193 6141 3205 6153
rect 3114 6101 3126 6113
rect 3094 6087 3106 6099
rect 3134 6087 3146 6099
rect 3234 6141 3246 6153
rect 3314 6101 3326 6113
rect 3294 6087 3306 6099
rect 3474 6161 3486 6173
rect 3453 6141 3465 6153
rect 3394 6101 3406 6113
rect 3334 6087 3346 6099
rect 3534 6161 3546 6173
rect 3494 6141 3506 6153
rect 3514 6141 3526 6153
rect 3555 6141 3567 6153
rect 3614 6101 3626 6113
rect 3694 6101 3706 6113
rect 3674 6087 3686 6099
rect 3794 6107 3806 6119
rect 3714 6087 3726 6099
rect 3834 6107 3846 6119
rect 3854 6107 3866 6119
rect 3955 6141 3967 6153
rect 3894 6107 3906 6119
rect 4014 6121 4026 6133
rect 4034 6121 4046 6133
rect 3994 6087 4006 6099
rect 4093 6141 4105 6153
rect 4054 6087 4066 6099
rect 4154 6121 4166 6133
rect 4194 6121 4206 6133
rect 4214 6101 4226 6113
rect 4294 6107 4306 6119
rect 4354 6121 4366 6133
rect 4334 6107 4346 6119
rect 4394 6107 4406 6119
rect 4475 6141 4487 6153
rect 4395 6070 4407 6082
rect 4534 6121 4546 6133
rect 4514 6087 4526 6099
rect 4674 6161 4686 6173
rect 4654 6141 4666 6153
rect 4614 6101 4626 6113
rect 4594 6087 4606 6099
rect 4634 6087 4646 6099
rect 4695 6141 4707 6153
rect 4914 6161 4926 6173
rect 4893 6141 4905 6153
rect 4814 6101 4826 6113
rect 4794 6087 4806 6099
rect 4834 6087 4846 6099
rect 4974 6161 4986 6173
rect 4934 6141 4946 6153
rect 4954 6141 4966 6153
rect 4995 6141 5007 6153
rect 5075 6141 5087 6153
rect 5134 6121 5146 6133
rect 5114 6087 5126 6099
rect 5174 6107 5186 6119
rect 5234 6121 5246 6133
rect 5214 6107 5226 6119
rect 5274 6107 5286 6119
rect 5334 6121 5346 6133
rect 5275 6070 5287 6082
rect 5393 6141 5405 6153
rect 5354 6087 5366 6099
rect 5594 6161 5606 6173
rect 5573 6141 5585 6153
rect 5494 6101 5506 6113
rect 5474 6087 5486 6099
rect 5514 6087 5526 6099
rect 5654 6161 5666 6173
rect 5614 6141 5626 6153
rect 5634 6141 5646 6153
rect 5675 6141 5687 6153
rect 5854 6161 5866 6173
rect 5834 6141 5846 6153
rect 5794 6101 5806 6113
rect 5774 6087 5786 6099
rect 5814 6087 5826 6099
rect 5875 6141 5887 6153
rect 5934 6121 5946 6133
rect 5993 6141 6005 6153
rect 5954 6087 5966 6099
rect 6034 6121 6046 6133
rect 6154 6161 6166 6173
rect 6093 6141 6105 6153
rect 6134 6141 6146 6153
rect 6054 6087 6066 6099
rect 6254 6161 6266 6173
rect 6175 6141 6187 6153
rect 6234 6141 6246 6153
rect 6275 6141 6287 6153
rect 6394 6161 6406 6173
rect 6373 6141 6385 6153
rect 6414 6141 6426 6153
rect 6494 6101 6506 6113
rect 6474 6087 6486 6099
rect 6534 6101 6546 6113
rect 6594 6101 6606 6113
rect 6514 6087 6526 6099
rect 45 5938 57 5950
rect 94 5901 106 5913
rect 74 5887 86 5899
rect 45 5870 57 5882
rect 134 5901 146 5913
rect 174 5901 186 5913
rect 294 5921 306 5933
rect 214 5901 226 5913
rect 334 5921 346 5933
rect 314 5907 326 5919
rect 374 5901 386 5913
rect 414 5901 426 5913
rect 434 5907 446 5919
rect 674 5921 686 5933
rect 514 5887 526 5899
rect 554 5887 566 5899
rect 574 5887 586 5899
rect 614 5887 626 5899
rect 654 5887 666 5899
rect 794 5907 806 5919
rect 713 5867 725 5879
rect 914 5901 926 5913
rect 814 5887 826 5899
rect 854 5887 866 5899
rect 954 5901 966 5913
rect 1034 5921 1046 5933
rect 995 5867 1007 5879
rect 1194 5907 1206 5919
rect 1054 5887 1066 5899
rect 1074 5887 1086 5899
rect 1114 5887 1126 5899
rect 1247 5915 1259 5927
rect 1233 5876 1245 5888
rect 1301 5948 1313 5960
rect 1261 5844 1273 5856
rect 1285 5844 1297 5856
rect 1349 5952 1361 5964
rect 1371 5952 1383 5964
rect 1333 5850 1345 5862
rect 1313 5830 1325 5842
rect 1374 5920 1386 5932
rect 1394 5906 1406 5918
rect 1414 5907 1426 5919
rect 1365 5864 1377 5876
rect 1347 5830 1359 5842
rect 1454 5901 1466 5913
rect 1494 5901 1506 5913
rect 1573 5867 1585 5879
rect 1694 5921 1706 5933
rect 1614 5867 1626 5879
rect 1655 5867 1667 5879
rect 1594 5847 1606 5859
rect 1714 5887 1726 5899
rect 1754 5887 1766 5899
rect 1794 5887 1806 5899
rect 1853 5867 1865 5879
rect 1914 5907 1926 5919
rect 1894 5867 1906 5879
rect 1874 5847 1886 5859
rect 2034 5921 2046 5933
rect 1995 5867 2007 5879
rect 2054 5887 2066 5899
rect 2074 5867 2086 5879
rect 2214 5921 2226 5933
rect 2115 5867 2127 5879
rect 2094 5847 2106 5859
rect 2254 5921 2266 5933
rect 2234 5907 2246 5919
rect 2294 5921 2306 5933
rect 2274 5887 2286 5899
rect 2394 5901 2406 5913
rect 2333 5867 2345 5879
rect 2434 5901 2446 5913
rect 2493 5867 2505 5879
rect 2594 5921 2606 5933
rect 2534 5867 2546 5879
rect 2514 5847 2526 5859
rect 2634 5921 2646 5933
rect 2614 5907 2626 5919
rect 2654 5901 2666 5913
rect 2694 5901 2706 5913
rect 2773 5867 2785 5879
rect 2814 5867 2826 5879
rect 2873 5867 2885 5879
rect 2794 5847 2806 5859
rect 2914 5867 2926 5879
rect 2973 5867 2985 5879
rect 2894 5847 2906 5859
rect 3014 5867 3026 5879
rect 3073 5867 3085 5879
rect 2994 5847 3006 5859
rect 3114 5867 3126 5879
rect 3134 5867 3146 5879
rect 3094 5847 3106 5859
rect 3294 5921 3306 5933
rect 3175 5867 3187 5879
rect 3255 5867 3267 5879
rect 3154 5847 3166 5859
rect 3354 5921 3366 5933
rect 3314 5887 3326 5899
rect 3334 5887 3346 5899
rect 3474 5921 3486 5933
rect 3393 5867 3405 5879
rect 3514 5921 3526 5933
rect 3494 5907 3506 5919
rect 3594 5921 3606 5933
rect 3555 5867 3567 5879
rect 3614 5887 3626 5899
rect 3673 5867 3685 5879
rect 3734 5921 3746 5933
rect 3774 5921 3786 5933
rect 3754 5907 3766 5919
rect 3714 5867 3726 5879
rect 3694 5847 3706 5859
rect 3873 5867 3885 5879
rect 3974 5921 3986 5933
rect 3914 5867 3926 5879
rect 3894 5847 3906 5859
rect 4014 5921 4026 5933
rect 3994 5907 4006 5919
rect 4073 5867 4085 5879
rect 4174 5921 4186 5933
rect 4114 5867 4126 5879
rect 4094 5847 4106 5859
rect 4214 5921 4226 5933
rect 4194 5907 4206 5919
rect 4234 5867 4246 5879
rect 4334 5901 4346 5913
rect 4275 5867 4287 5879
rect 4254 5847 4266 5859
rect 4374 5901 4386 5913
rect 4474 5921 4486 5933
rect 4435 5867 4447 5879
rect 4635 5938 4647 5950
rect 4634 5901 4646 5913
rect 4494 5887 4506 5899
rect 4534 5887 4546 5899
rect 4574 5887 4586 5899
rect 4594 5887 4606 5899
rect 4734 5921 4746 5933
rect 4774 5921 4786 5933
rect 4754 5907 4766 5919
rect 4794 5901 4806 5913
rect 4834 5901 4846 5913
rect 4914 5907 4926 5919
rect 4973 5867 4985 5879
rect 5034 5921 5046 5933
rect 5074 5921 5086 5933
rect 5054 5907 5066 5919
rect 5014 5867 5026 5879
rect 4994 5847 5006 5859
rect 5154 5921 5166 5933
rect 5134 5887 5146 5899
rect 5254 5921 5266 5933
rect 5234 5887 5246 5899
rect 5193 5867 5205 5879
rect 5355 5921 5367 5933
rect 5393 5921 5405 5933
rect 5335 5887 5347 5899
rect 5293 5867 5305 5879
rect 5474 5901 5486 5913
rect 5414 5887 5426 5899
rect 5514 5901 5526 5913
rect 5534 5907 5546 5919
rect 5633 5867 5645 5879
rect 5694 5921 5706 5933
rect 5734 5921 5746 5933
rect 5714 5907 5726 5919
rect 5674 5867 5686 5879
rect 5654 5847 5666 5859
rect 5854 5921 5866 5933
rect 5815 5867 5827 5879
rect 5914 5921 5926 5933
rect 5874 5887 5886 5899
rect 5894 5887 5906 5899
rect 6054 5921 6066 5933
rect 5953 5867 5965 5879
rect 6015 5867 6027 5879
rect 6115 5921 6127 5933
rect 6153 5921 6165 5933
rect 6074 5887 6086 5899
rect 6095 5887 6107 5899
rect 6234 5901 6246 5913
rect 6174 5887 6186 5899
rect 6274 5901 6286 5913
rect 6335 5938 6347 5950
rect 6334 5901 6346 5913
rect 6294 5887 6306 5899
rect 6414 5921 6426 5933
rect 6394 5887 6406 5899
rect 6453 5867 6465 5879
rect 6494 5867 6506 5879
rect 6594 5901 6606 5913
rect 6535 5867 6547 5879
rect 6514 5847 6526 5859
rect 6634 5901 6646 5913
rect 45 5658 57 5670
rect 125 5658 137 5670
rect 221 5684 233 5696
rect 273 5698 285 5710
rect 245 5684 257 5696
rect 74 5641 86 5653
rect 154 5641 166 5653
rect 193 5652 205 5664
rect 45 5590 57 5602
rect 125 5590 137 5602
rect 207 5613 219 5625
rect 261 5580 273 5592
rect 307 5698 319 5710
rect 293 5678 305 5690
rect 325 5664 337 5676
rect 354 5622 366 5634
rect 434 5641 446 5653
rect 474 5641 486 5653
rect 334 5608 346 5620
rect 309 5576 321 5588
rect 331 5576 343 5588
rect 374 5621 386 5633
rect 514 5621 526 5633
rect 494 5607 506 5619
rect 594 5627 606 5639
rect 534 5607 546 5619
rect 674 5641 686 5653
rect 634 5627 646 5639
rect 714 5627 726 5639
rect 774 5627 786 5639
rect 814 5627 826 5639
rect 854 5627 866 5639
rect 715 5590 727 5602
rect 934 5641 946 5653
rect 974 5641 986 5653
rect 894 5627 906 5639
rect 1113 5659 1125 5671
rect 1094 5641 1106 5653
rect 1174 5641 1186 5653
rect 1214 5641 1226 5653
rect 1014 5621 1026 5633
rect 1074 5621 1086 5633
rect 1113 5592 1125 5604
rect 1314 5641 1326 5653
rect 1354 5641 1366 5653
rect 1254 5621 1266 5633
rect 1501 5684 1513 5696
rect 1553 5698 1565 5710
rect 1525 5684 1537 5696
rect 1394 5621 1406 5633
rect 1473 5652 1485 5664
rect 1487 5613 1499 5625
rect 1541 5580 1553 5592
rect 1587 5698 1599 5710
rect 1573 5678 1585 5690
rect 1605 5664 1617 5676
rect 1634 5622 1646 5634
rect 1694 5641 1706 5653
rect 1614 5608 1626 5620
rect 1589 5576 1601 5588
rect 1611 5576 1623 5588
rect 1654 5621 1666 5633
rect 1835 5661 1847 5673
rect 1773 5641 1785 5653
rect 1714 5607 1726 5619
rect 1750 5607 1762 5619
rect 1894 5641 1906 5653
rect 1874 5607 1886 5619
rect 1934 5627 1946 5639
rect 1974 5627 1986 5639
rect 1994 5621 2006 5633
rect 2114 5621 2126 5633
rect 2094 5607 2106 5619
rect 2154 5641 2166 5653
rect 2194 5641 2206 5653
rect 2134 5607 2146 5619
rect 2234 5627 2246 5639
rect 2394 5641 2406 5653
rect 2274 5627 2286 5639
rect 2414 5607 2426 5619
rect 2454 5641 2466 5653
rect 2514 5627 2526 5639
rect 2634 5681 2646 5693
rect 2613 5661 2625 5673
rect 2554 5627 2566 5639
rect 2734 5681 2746 5693
rect 2654 5661 2666 5673
rect 2713 5661 2725 5673
rect 2754 5661 2766 5673
rect 2774 5627 2786 5639
rect 2854 5641 2866 5653
rect 2814 5627 2826 5639
rect 3014 5681 3026 5693
rect 2913 5661 2925 5673
rect 2993 5661 3005 5673
rect 2874 5607 2886 5619
rect 3034 5661 3046 5673
rect 3074 5621 3086 5633
rect 3054 5607 3066 5619
rect 3175 5661 3187 5673
rect 3094 5607 3106 5619
rect 3234 5641 3246 5653
rect 3214 5607 3226 5619
rect 3334 5681 3346 5693
rect 3314 5661 3326 5673
rect 3294 5621 3306 5633
rect 3355 5661 3367 5673
rect 3474 5681 3486 5693
rect 3453 5661 3465 5673
rect 3574 5681 3586 5693
rect 3494 5661 3506 5673
rect 3553 5661 3565 5673
rect 3594 5661 3606 5673
rect 3695 5661 3707 5673
rect 3654 5621 3666 5633
rect 3754 5641 3766 5653
rect 3794 5641 3806 5653
rect 3834 5641 3846 5653
rect 3854 5641 3866 5653
rect 3734 5607 3746 5619
rect 3913 5661 3925 5673
rect 3874 5607 3886 5619
rect 4034 5641 4046 5653
rect 3994 5621 4006 5633
rect 4155 5661 4167 5673
rect 4113 5641 4125 5653
rect 4055 5607 4067 5619
rect 4093 5607 4105 5619
rect 4294 5681 4306 5693
rect 4273 5661 4285 5673
rect 4214 5641 4226 5653
rect 4194 5607 4206 5619
rect 4314 5661 4326 5673
rect 4415 5661 4427 5673
rect 4334 5621 4346 5633
rect 4474 5641 4486 5653
rect 4454 5607 4466 5619
rect 4574 5641 4586 5653
rect 4534 5627 4546 5639
rect 4533 5590 4545 5602
rect 4594 5627 4606 5639
rect 4695 5661 4707 5673
rect 4634 5627 4646 5639
rect 4754 5641 4766 5653
rect 4774 5641 4786 5653
rect 4734 5607 4746 5619
rect 4934 5681 4946 5693
rect 4833 5661 4845 5673
rect 4913 5661 4925 5673
rect 4794 5607 4806 5619
rect 4954 5661 4966 5673
rect 4994 5621 5006 5633
rect 4974 5607 4986 5619
rect 5074 5641 5086 5653
rect 5014 5607 5026 5619
rect 5194 5681 5206 5693
rect 5133 5661 5145 5673
rect 5174 5661 5186 5673
rect 5094 5607 5106 5619
rect 5215 5661 5227 5673
rect 5274 5627 5286 5639
rect 5374 5681 5386 5693
rect 5354 5661 5366 5673
rect 5314 5627 5326 5639
rect 5395 5661 5407 5673
rect 5474 5621 5486 5633
rect 5454 5607 5466 5619
rect 5554 5627 5566 5639
rect 5494 5607 5506 5619
rect 5594 5627 5606 5639
rect 5654 5627 5666 5639
rect 5715 5641 5727 5653
rect 5694 5627 5706 5639
rect 5855 5661 5867 5673
rect 5794 5641 5806 5653
rect 5735 5607 5747 5619
rect 5773 5607 5785 5619
rect 5914 5641 5926 5653
rect 5894 5607 5906 5619
rect 5995 5641 6007 5653
rect 5934 5621 5946 5633
rect 6134 5681 6146 5693
rect 6114 5661 6126 5673
rect 6074 5641 6086 5653
rect 6015 5607 6027 5619
rect 6053 5607 6065 5619
rect 6155 5661 6167 5673
rect 6254 5621 6266 5633
rect 6294 5621 6306 5633
rect 6274 5607 6286 5619
rect 6394 5681 6406 5693
rect 6374 5661 6386 5673
rect 6314 5607 6326 5619
rect 6494 5681 6506 5693
rect 6415 5661 6427 5673
rect 6474 5661 6486 5673
rect 6594 5681 6606 5693
rect 6515 5661 6527 5673
rect 6574 5661 6586 5673
rect 6615 5661 6627 5673
rect 47 5435 59 5447
rect 33 5396 45 5408
rect 101 5468 113 5480
rect 61 5364 73 5376
rect 85 5364 97 5376
rect 149 5472 161 5484
rect 171 5472 183 5484
rect 133 5370 145 5382
rect 113 5350 125 5362
rect 174 5440 186 5452
rect 194 5426 206 5438
rect 214 5427 226 5439
rect 165 5384 177 5396
rect 147 5350 159 5362
rect 254 5421 266 5433
rect 374 5441 386 5453
rect 294 5421 306 5433
rect 414 5441 426 5453
rect 553 5458 565 5470
rect 394 5427 406 5439
rect 454 5421 466 5433
rect 494 5421 506 5433
rect 554 5421 566 5433
rect 774 5421 786 5433
rect 594 5407 606 5419
rect 614 5407 626 5419
rect 654 5407 666 5419
rect 694 5407 706 5419
rect 734 5407 746 5419
rect 814 5421 826 5433
rect 854 5421 866 5433
rect 994 5441 1006 5453
rect 894 5421 906 5433
rect 934 5427 946 5439
rect 1034 5441 1046 5453
rect 1014 5427 1026 5439
rect 1135 5441 1147 5453
rect 1173 5441 1185 5453
rect 1114 5407 1126 5419
rect 1193 5407 1205 5419
rect 1247 5435 1259 5447
rect 1233 5396 1245 5408
rect 1301 5468 1313 5480
rect 1261 5364 1273 5376
rect 1285 5364 1297 5376
rect 1349 5472 1361 5484
rect 1371 5472 1383 5484
rect 1333 5370 1345 5382
rect 1313 5350 1325 5362
rect 1374 5440 1386 5452
rect 1394 5426 1406 5438
rect 1414 5427 1426 5439
rect 1365 5384 1377 5396
rect 1347 5350 1359 5362
rect 1493 5387 1505 5399
rect 1534 5387 1546 5399
rect 1593 5387 1605 5399
rect 1514 5367 1526 5379
rect 1694 5427 1706 5439
rect 1634 5387 1646 5399
rect 1614 5367 1626 5379
rect 1774 5441 1786 5453
rect 1735 5387 1747 5399
rect 1853 5458 1865 5470
rect 1794 5407 1806 5419
rect 1854 5421 1866 5433
rect 1934 5421 1946 5433
rect 1894 5407 1906 5419
rect 1974 5421 1986 5433
rect 2054 5441 2066 5453
rect 2015 5387 2027 5399
rect 2094 5421 2106 5433
rect 2074 5407 2086 5419
rect 2134 5421 2146 5433
rect 2214 5427 2226 5439
rect 2294 5441 2306 5453
rect 2255 5387 2267 5399
rect 2514 5441 2526 5453
rect 2454 5427 2466 5439
rect 2314 5407 2326 5419
rect 2334 5407 2346 5419
rect 2374 5407 2386 5419
rect 2554 5441 2566 5453
rect 2534 5427 2546 5439
rect 2594 5441 2606 5453
rect 2574 5407 2586 5419
rect 2674 5421 2686 5433
rect 2633 5387 2645 5399
rect 2714 5421 2726 5433
rect 2793 5387 2805 5399
rect 2874 5421 2886 5433
rect 2834 5387 2846 5399
rect 2814 5367 2826 5379
rect 2914 5421 2926 5433
rect 3034 5441 3046 5453
rect 2954 5407 2966 5419
rect 2994 5407 3006 5419
rect 3014 5407 3026 5419
rect 3134 5421 3146 5433
rect 3073 5387 3085 5399
rect 3174 5421 3186 5433
rect 3214 5441 3226 5453
rect 3194 5407 3206 5419
rect 3333 5458 3345 5470
rect 3253 5387 3265 5399
rect 3334 5421 3346 5433
rect 3474 5427 3486 5439
rect 3374 5407 3386 5419
rect 3394 5407 3406 5419
rect 3434 5407 3446 5419
rect 3513 5456 3525 5468
rect 3594 5441 3606 5453
rect 3494 5407 3506 5419
rect 3574 5407 3586 5419
rect 3513 5389 3525 5401
rect 3774 5441 3786 5453
rect 3810 5441 3822 5453
rect 3694 5407 3706 5419
rect 3633 5387 3645 5399
rect 3734 5407 3746 5419
rect 3754 5407 3766 5419
rect 3974 5441 3986 5453
rect 3833 5407 3845 5419
rect 3894 5407 3906 5419
rect 3934 5407 3946 5419
rect 3954 5407 3966 5419
rect 4013 5387 4025 5399
rect 4093 5387 4105 5399
rect 4174 5421 4186 5433
rect 4134 5387 4146 5399
rect 4114 5367 4126 5379
rect 4214 5421 4226 5433
rect 4234 5427 4246 5439
rect 4354 5441 4366 5453
rect 4315 5387 4327 5399
rect 4414 5421 4426 5433
rect 4374 5407 4386 5419
rect 4454 5421 4466 5433
rect 4474 5421 4486 5433
rect 4514 5421 4526 5433
rect 4614 5441 4626 5453
rect 4575 5387 4587 5399
rect 4634 5407 4646 5419
rect 4714 5441 4726 5453
rect 4675 5387 4687 5399
rect 4793 5458 4805 5470
rect 4734 5407 4746 5419
rect 4794 5421 4806 5433
rect 4834 5407 4846 5419
rect 4914 5441 4926 5453
rect 4875 5387 4887 5399
rect 5073 5458 5085 5470
rect 4974 5421 4986 5433
rect 4934 5407 4946 5419
rect 5014 5421 5026 5433
rect 5074 5421 5086 5433
rect 5134 5421 5146 5433
rect 5114 5407 5126 5419
rect 5174 5421 5186 5433
rect 5234 5441 5246 5453
rect 5214 5407 5226 5419
rect 5353 5458 5365 5470
rect 5273 5387 5285 5399
rect 5354 5421 5366 5433
rect 5434 5441 5446 5453
rect 5394 5407 5406 5419
rect 5414 5407 5426 5419
rect 5733 5458 5745 5470
rect 5514 5421 5526 5433
rect 5473 5387 5485 5399
rect 5554 5421 5566 5433
rect 5594 5387 5606 5399
rect 5635 5387 5647 5399
rect 5614 5367 5626 5379
rect 5734 5421 5746 5433
rect 5835 5441 5847 5453
rect 5873 5441 5885 5453
rect 5774 5407 5786 5419
rect 5814 5407 5826 5419
rect 5914 5421 5926 5433
rect 5893 5407 5905 5419
rect 5954 5421 5966 5433
rect 5994 5387 6006 5399
rect 6094 5441 6106 5453
rect 6134 5441 6146 5453
rect 6114 5427 6126 5439
rect 6035 5387 6047 5399
rect 6014 5367 6026 5379
rect 6254 5441 6266 5453
rect 6215 5387 6227 5399
rect 6314 5441 6326 5453
rect 6274 5407 6286 5419
rect 6294 5407 6306 5419
rect 6454 5441 6466 5453
rect 6353 5387 6365 5399
rect 6415 5387 6427 5399
rect 6474 5407 6486 5419
rect 6533 5387 6545 5399
rect 6634 5441 6646 5453
rect 6574 5387 6586 5399
rect 6554 5367 6566 5379
rect 6674 5441 6686 5453
rect 6654 5427 6666 5439
rect 45 5178 57 5190
rect 141 5204 153 5216
rect 193 5218 205 5230
rect 165 5204 177 5216
rect 74 5161 86 5173
rect 113 5172 125 5184
rect 45 5110 57 5122
rect 127 5133 139 5145
rect 181 5100 193 5112
rect 227 5218 239 5230
rect 213 5198 225 5210
rect 245 5184 257 5196
rect 274 5142 286 5154
rect 254 5128 266 5140
rect 229 5096 241 5108
rect 251 5096 263 5108
rect 294 5141 306 5153
rect 334 5147 346 5159
rect 374 5147 386 5159
rect 474 5141 486 5153
rect 454 5127 466 5139
rect 534 5147 546 5159
rect 494 5127 506 5139
rect 574 5147 586 5159
rect 681 5218 693 5230
rect 663 5184 675 5196
rect 614 5141 626 5153
rect 634 5142 646 5154
rect 654 5128 666 5140
rect 715 5218 727 5230
rect 695 5198 707 5210
rect 657 5096 669 5108
rect 679 5096 691 5108
rect 743 5204 755 5216
rect 767 5204 779 5216
rect 727 5100 739 5112
rect 795 5172 807 5184
rect 781 5133 793 5145
rect 834 5147 846 5159
rect 935 5181 947 5193
rect 874 5147 886 5159
rect 1035 5181 1047 5193
rect 994 5161 1006 5173
rect 974 5127 986 5139
rect 1094 5161 1106 5173
rect 1074 5127 1086 5139
rect 1261 5204 1273 5216
rect 1313 5218 1325 5230
rect 1285 5204 1297 5216
rect 1194 5161 1206 5173
rect 1233 5172 1245 5184
rect 1154 5147 1166 5159
rect 1153 5110 1165 5122
rect 1247 5133 1259 5145
rect 1301 5100 1313 5112
rect 1347 5218 1359 5230
rect 1333 5198 1345 5210
rect 1365 5184 1377 5196
rect 1394 5142 1406 5154
rect 1374 5128 1386 5140
rect 1349 5096 1361 5108
rect 1371 5096 1383 5108
rect 1414 5141 1426 5153
rect 1474 5147 1486 5159
rect 1514 5147 1526 5159
rect 1534 5147 1546 5159
rect 1661 5204 1673 5216
rect 1713 5218 1725 5230
rect 1685 5204 1697 5216
rect 1633 5172 1645 5184
rect 1574 5147 1586 5159
rect 1647 5133 1659 5145
rect 1701 5100 1713 5112
rect 1747 5218 1759 5230
rect 1733 5198 1745 5210
rect 1765 5184 1777 5196
rect 1794 5142 1806 5154
rect 1874 5161 1886 5173
rect 1774 5128 1786 5140
rect 1749 5096 1761 5108
rect 1771 5096 1783 5108
rect 1814 5141 1826 5153
rect 1953 5161 1965 5173
rect 1895 5127 1907 5139
rect 1933 5127 1945 5139
rect 1974 5141 1986 5153
rect 2114 5161 2126 5173
rect 2074 5147 2086 5159
rect 2073 5110 2085 5122
rect 2134 5147 2146 5159
rect 2255 5179 2267 5191
rect 2274 5161 2286 5173
rect 2174 5147 2186 5159
rect 2255 5112 2267 5124
rect 2294 5141 2306 5153
rect 2334 5147 2346 5159
rect 2454 5201 2466 5213
rect 2433 5181 2445 5193
rect 2374 5147 2386 5159
rect 2474 5181 2486 5193
rect 2514 5161 2526 5173
rect 2554 5161 2566 5173
rect 2574 5141 2586 5153
rect 2714 5161 2726 5173
rect 2734 5161 2746 5173
rect 2774 5161 2786 5173
rect 2674 5147 2686 5159
rect 2673 5110 2685 5122
rect 2834 5147 2846 5159
rect 2874 5147 2886 5159
rect 2914 5147 2926 5159
rect 2954 5147 2966 5159
rect 3013 5179 3025 5191
rect 2994 5161 3006 5173
rect 2974 5141 2986 5153
rect 3013 5112 3025 5124
rect 3154 5161 3166 5173
rect 3114 5147 3126 5159
rect 3113 5110 3125 5122
rect 3174 5147 3186 5159
rect 3314 5201 3326 5213
rect 3293 5181 3305 5193
rect 3214 5147 3226 5159
rect 3334 5181 3346 5193
rect 3394 5141 3406 5153
rect 3474 5141 3486 5153
rect 3454 5127 3466 5139
rect 3534 5161 3546 5173
rect 3574 5161 3586 5173
rect 3594 5161 3606 5173
rect 3494 5127 3506 5139
rect 3653 5181 3665 5193
rect 3715 5181 3727 5193
rect 3614 5127 3626 5139
rect 3774 5161 3786 5173
rect 3794 5161 3806 5173
rect 3834 5161 3846 5173
rect 3754 5127 3766 5139
rect 3874 5147 3886 5159
rect 3914 5147 3926 5159
rect 3974 5147 3986 5159
rect 4034 5161 4046 5173
rect 4014 5147 4026 5159
rect 4093 5181 4105 5193
rect 4054 5127 4066 5139
rect 4154 5147 4166 5159
rect 4194 5147 4206 5159
rect 4294 5161 4306 5173
rect 4254 5147 4266 5159
rect 4253 5110 4265 5122
rect 4334 5147 4346 5159
rect 4415 5181 4427 5193
rect 4374 5147 4386 5159
rect 4515 5181 4527 5193
rect 4474 5161 4486 5173
rect 4454 5127 4466 5139
rect 4574 5161 4586 5173
rect 4554 5127 4566 5139
rect 4594 5147 4606 5159
rect 4634 5147 4646 5159
rect 4674 5147 4686 5159
rect 4714 5147 4726 5159
rect 4874 5201 4886 5213
rect 4853 5181 4865 5193
rect 4754 5141 4766 5153
rect 4894 5181 4906 5193
rect 4914 5161 4926 5173
rect 4973 5181 4985 5193
rect 4934 5127 4946 5139
rect 5074 5147 5086 5159
rect 5014 5127 5026 5139
rect 5114 5147 5126 5159
rect 5234 5147 5246 5159
rect 5154 5127 5166 5139
rect 5314 5161 5326 5173
rect 5274 5147 5286 5159
rect 5434 5201 5446 5213
rect 5373 5181 5385 5193
rect 5414 5181 5426 5193
rect 5334 5127 5346 5139
rect 5534 5201 5546 5213
rect 5455 5181 5467 5193
rect 5514 5181 5526 5193
rect 5555 5181 5567 5193
rect 5694 5201 5706 5213
rect 5674 5181 5686 5193
rect 5614 5141 5626 5153
rect 5715 5181 5727 5193
rect 5774 5161 5786 5173
rect 5833 5181 5845 5193
rect 5794 5127 5806 5139
rect 5894 5147 5906 5159
rect 5974 5201 5986 5213
rect 5954 5181 5966 5193
rect 5934 5147 5946 5159
rect 5995 5181 6007 5193
rect 6054 5147 6066 5159
rect 6094 5147 6106 5159
rect 6194 5141 6206 5153
rect 6174 5127 6186 5139
rect 6354 5201 6366 5213
rect 6333 5181 6345 5193
rect 6274 5141 6286 5153
rect 6214 5127 6226 5139
rect 6454 5201 6466 5213
rect 6374 5181 6386 5193
rect 6433 5181 6445 5193
rect 6474 5181 6486 5193
rect 6614 5201 6626 5213
rect 6593 5181 6605 5193
rect 6494 5141 6506 5153
rect 6634 5181 6646 5193
rect 6654 5147 6666 5159
rect 6694 5147 6706 5159
rect 45 4978 57 4990
rect 125 4978 137 4990
rect 194 4941 206 4953
rect 74 4927 86 4939
rect 154 4927 166 4939
rect 45 4910 57 4922
rect 125 4910 137 4922
rect 234 4941 246 4953
rect 287 4955 299 4967
rect 273 4916 285 4928
rect 341 4988 353 5000
rect 301 4884 313 4896
rect 325 4884 337 4896
rect 389 4992 401 5004
rect 411 4992 423 5004
rect 373 4890 385 4902
rect 353 4870 365 4882
rect 414 4960 426 4972
rect 534 4961 546 4973
rect 434 4946 446 4958
rect 454 4947 466 4959
rect 405 4904 417 4916
rect 387 4870 399 4882
rect 574 4961 586 4973
rect 554 4947 566 4959
rect 614 4941 626 4953
rect 654 4941 666 4953
rect 674 4941 686 4953
rect 714 4941 726 4953
rect 774 4941 786 4953
rect 814 4941 826 4953
rect 867 4955 879 4967
rect 853 4916 865 4928
rect 921 4988 933 5000
rect 881 4884 893 4896
rect 905 4884 917 4896
rect 969 4992 981 5004
rect 991 4992 1003 5004
rect 953 4890 965 4902
rect 933 4870 945 4882
rect 994 4960 1006 4972
rect 1105 4978 1117 4990
rect 1014 4946 1026 4958
rect 1034 4947 1046 4959
rect 985 4904 997 4916
rect 967 4870 979 4882
rect 1194 4961 1206 4973
rect 1134 4927 1146 4939
rect 1105 4910 1117 4922
rect 1234 4961 1246 4973
rect 1365 4978 1377 4990
rect 1214 4947 1226 4959
rect 1274 4941 1286 4953
rect 1314 4941 1326 4953
rect 1414 4941 1426 4953
rect 1394 4927 1406 4939
rect 1365 4910 1377 4922
rect 1454 4941 1466 4953
rect 1514 4941 1526 4953
rect 1554 4941 1566 4953
rect 1634 4961 1646 4973
rect 1595 4907 1607 4919
rect 1694 4941 1706 4953
rect 1654 4927 1666 4939
rect 1734 4941 1746 4953
rect 1814 4961 1826 4973
rect 1775 4907 1787 4919
rect 1854 4941 1866 4953
rect 1834 4927 1846 4939
rect 1894 4941 1906 4953
rect 1994 4961 2006 4973
rect 1955 4907 1967 4919
rect 2014 4927 2026 4939
rect 2094 4961 2106 4973
rect 2055 4907 2067 4919
rect 2173 4978 2185 4990
rect 2114 4927 2126 4939
rect 2174 4941 2186 4953
rect 2234 4947 2246 4959
rect 2214 4927 2226 4939
rect 2415 4976 2427 4988
rect 2454 4947 2466 4959
rect 2314 4927 2326 4939
rect 2354 4927 2366 4939
rect 2434 4927 2446 4939
rect 2415 4909 2427 4921
rect 2494 4941 2506 4953
rect 2534 4941 2546 4953
rect 2614 4961 2626 4973
rect 2575 4907 2587 4919
rect 2634 4927 2646 4939
rect 2714 4961 2726 4973
rect 2675 4907 2687 4919
rect 2794 4947 2806 4959
rect 2734 4927 2746 4939
rect 2834 4961 2846 4973
rect 2814 4927 2826 4939
rect 2974 4961 2986 4973
rect 2873 4907 2885 4919
rect 2935 4907 2947 4919
rect 2994 4927 3006 4939
rect 3074 4961 3086 4973
rect 3035 4907 3047 4919
rect 3234 4961 3246 4973
rect 3094 4927 3106 4939
rect 3134 4927 3146 4939
rect 3174 4927 3186 4939
rect 3274 4941 3286 4953
rect 3314 4941 3326 4953
rect 3394 4961 3406 4973
rect 3355 4907 3367 4919
rect 3454 4947 3466 4959
rect 3497 4992 3509 5004
rect 3519 4992 3531 5004
rect 3494 4960 3506 4972
rect 3414 4927 3426 4939
rect 3474 4946 3486 4958
rect 3503 4904 3515 4916
rect 3535 4890 3547 4902
rect 3521 4870 3533 4882
rect 3567 4988 3579 5000
rect 3621 4955 3633 4967
rect 3694 4961 3706 4973
rect 3635 4916 3647 4928
rect 3674 4927 3686 4939
rect 3814 4961 3826 4973
rect 3733 4907 3745 4919
rect 3583 4884 3595 4896
rect 3555 4870 3567 4882
rect 3607 4884 3619 4896
rect 3854 4961 3866 4973
rect 3834 4947 3846 4959
rect 3913 4907 3925 4919
rect 4014 4961 4026 4973
rect 3954 4907 3966 4919
rect 3934 4887 3946 4899
rect 4173 4978 4185 4990
rect 4054 4961 4066 4973
rect 4114 4961 4126 4973
rect 4034 4947 4046 4959
rect 4174 4941 4186 4953
rect 4254 4941 4266 4953
rect 4214 4927 4226 4939
rect 4294 4941 4306 4953
rect 4355 4978 4367 4990
rect 4354 4941 4366 4953
rect 4314 4927 4326 4939
rect 4474 4961 4486 4973
rect 4435 4907 4447 4919
rect 4494 4927 4506 4939
rect 4514 4907 4526 4919
rect 4634 4961 4646 4973
rect 4614 4927 4626 4939
rect 4555 4907 4567 4919
rect 4534 4887 4546 4899
rect 4833 4978 4845 4990
rect 4734 4941 4746 4953
rect 4673 4907 4685 4919
rect 4774 4941 4786 4953
rect 4834 4941 4846 4953
rect 4914 4941 4926 4953
rect 4874 4927 4886 4939
rect 4954 4941 4966 4953
rect 4974 4941 4986 4953
rect 5014 4941 5026 4953
rect 5095 4978 5107 4990
rect 5094 4941 5106 4953
rect 5054 4927 5066 4939
rect 5273 4978 5285 4990
rect 5174 4941 5186 4953
rect 5214 4941 5226 4953
rect 5274 4941 5286 4953
rect 5375 4978 5387 4990
rect 5374 4941 5386 4953
rect 5314 4927 5326 4939
rect 5334 4927 5346 4939
rect 5475 4961 5487 4973
rect 5513 4961 5525 4973
rect 5454 4927 5466 4939
rect 5574 4941 5586 4953
rect 5533 4927 5545 4939
rect 5614 4941 5626 4953
rect 5634 4907 5646 4919
rect 5774 4961 5786 4973
rect 5675 4907 5687 4919
rect 5654 4887 5666 4899
rect 5814 4961 5826 4973
rect 5794 4947 5806 4959
rect 5873 4907 5885 4919
rect 5954 4941 5966 4953
rect 5914 4907 5926 4919
rect 5894 4887 5906 4899
rect 5994 4941 6006 4953
rect 6035 4961 6047 4973
rect 6073 4961 6085 4973
rect 6015 4927 6027 4939
rect 6094 4927 6106 4939
rect 6173 4907 6185 4919
rect 6254 4961 6266 4973
rect 6234 4927 6246 4939
rect 6214 4907 6226 4919
rect 6194 4887 6206 4899
rect 6293 4907 6305 4919
rect 6373 4907 6385 4919
rect 6414 4907 6426 4919
rect 6473 4907 6485 4919
rect 6394 4887 6406 4899
rect 6534 4941 6546 4953
rect 6514 4907 6526 4919
rect 6494 4887 6506 4899
rect 6574 4941 6586 4953
rect 6654 4947 6666 4959
rect 34 4647 46 4659
rect 234 4681 246 4693
rect 274 4681 286 4693
rect 70 4644 82 4656
rect 110 4644 122 4656
rect 150 4644 162 4656
rect 334 4661 346 4673
rect 414 4661 426 4673
rect 394 4647 406 4659
rect 534 4681 546 4693
rect 574 4681 586 4693
rect 494 4661 506 4673
rect 434 4647 446 4659
rect 674 4681 686 4693
rect 694 4681 706 4693
rect 805 4698 817 4710
rect 734 4681 746 4693
rect 834 4681 846 4693
rect 634 4667 646 4679
rect 633 4630 645 4642
rect 805 4630 817 4642
rect 874 4667 886 4679
rect 981 4724 993 4736
rect 1033 4738 1045 4750
rect 1005 4724 1017 4736
rect 953 4692 965 4704
rect 914 4667 926 4679
rect 967 4653 979 4665
rect 1021 4620 1033 4632
rect 1067 4738 1079 4750
rect 1053 4718 1065 4730
rect 1085 4704 1097 4716
rect 1114 4662 1126 4674
rect 1195 4701 1207 4713
rect 1094 4648 1106 4660
rect 1069 4616 1081 4628
rect 1091 4616 1103 4628
rect 1134 4661 1146 4673
rect 1254 4681 1266 4693
rect 1234 4647 1246 4659
rect 1294 4667 1306 4679
rect 1334 4667 1346 4679
rect 1354 4667 1366 4679
rect 1455 4701 1467 4713
rect 1394 4667 1406 4679
rect 1514 4681 1526 4693
rect 1534 4681 1546 4693
rect 1574 4681 1586 4693
rect 1614 4681 1626 4693
rect 1654 4681 1666 4693
rect 1494 4647 1506 4659
rect 1754 4681 1766 4693
rect 1794 4681 1806 4693
rect 1834 4681 1846 4693
rect 1694 4661 1706 4673
rect 1981 4724 1993 4736
rect 2033 4738 2045 4750
rect 2005 4724 2017 4736
rect 1893 4701 1905 4713
rect 1854 4647 1866 4659
rect 1953 4692 1965 4704
rect 1967 4653 1979 4665
rect 2021 4620 2033 4632
rect 2067 4738 2079 4750
rect 2053 4718 2065 4730
rect 2085 4704 2097 4716
rect 2114 4662 2126 4674
rect 2094 4648 2106 4660
rect 2069 4616 2081 4628
rect 2091 4616 2103 4628
rect 2134 4661 2146 4673
rect 2194 4667 2206 4679
rect 2295 4699 2307 4711
rect 2314 4681 2326 4693
rect 2234 4667 2246 4679
rect 2295 4632 2307 4644
rect 2334 4661 2346 4673
rect 2354 4667 2366 4679
rect 2434 4681 2446 4693
rect 2474 4681 2486 4693
rect 2394 4667 2406 4679
rect 2534 4661 2546 4673
rect 2514 4647 2526 4659
rect 2554 4647 2566 4659
rect 2721 4724 2733 4736
rect 2773 4738 2785 4750
rect 2745 4724 2757 4736
rect 2693 4692 2705 4704
rect 2654 4661 2666 4673
rect 2707 4653 2719 4665
rect 2761 4620 2773 4632
rect 2807 4738 2819 4750
rect 2793 4718 2805 4730
rect 2825 4704 2837 4716
rect 2854 4662 2866 4674
rect 2914 4681 2926 4693
rect 2834 4648 2846 4660
rect 2809 4616 2821 4628
rect 2831 4616 2843 4628
rect 2874 4661 2886 4673
rect 3061 4724 3073 4736
rect 3113 4738 3125 4750
rect 3085 4724 3097 4736
rect 2973 4701 2985 4713
rect 2934 4647 2946 4659
rect 3033 4692 3045 4704
rect 3047 4653 3059 4665
rect 3101 4620 3113 4632
rect 3147 4738 3159 4750
rect 3133 4718 3145 4730
rect 3165 4704 3177 4716
rect 3301 4724 3313 4736
rect 3353 4738 3365 4750
rect 3325 4724 3337 4736
rect 3194 4662 3206 4674
rect 3273 4692 3285 4704
rect 3174 4648 3186 4660
rect 3149 4616 3161 4628
rect 3171 4616 3183 4628
rect 3214 4661 3226 4673
rect 3287 4653 3299 4665
rect 3341 4620 3353 4632
rect 3387 4738 3399 4750
rect 3373 4718 3385 4730
rect 3405 4704 3417 4716
rect 3434 4662 3446 4674
rect 3515 4701 3527 4713
rect 3414 4648 3426 4660
rect 3389 4616 3401 4628
rect 3411 4616 3423 4628
rect 3454 4661 3466 4673
rect 3574 4681 3586 4693
rect 3554 4647 3566 4659
rect 3674 4667 3686 4679
rect 3634 4647 3646 4659
rect 3755 4701 3767 4713
rect 3714 4667 3726 4679
rect 3814 4681 3826 4693
rect 3794 4647 3806 4659
rect 3921 4738 3933 4750
rect 3903 4704 3915 4716
rect 3854 4661 3866 4673
rect 3874 4662 3886 4674
rect 3894 4648 3906 4660
rect 3955 4738 3967 4750
rect 3935 4718 3947 4730
rect 3897 4616 3909 4628
rect 3919 4616 3931 4628
rect 3983 4724 3995 4736
rect 4007 4724 4019 4736
rect 3967 4620 3979 4632
rect 4035 4692 4047 4704
rect 4021 4653 4033 4665
rect 4154 4667 4166 4679
rect 4114 4647 4126 4659
rect 4261 4724 4273 4736
rect 4313 4738 4325 4750
rect 4285 4724 4297 4736
rect 4233 4692 4245 4704
rect 4194 4667 4206 4679
rect 4247 4653 4259 4665
rect 4301 4620 4313 4632
rect 4347 4738 4359 4750
rect 4333 4718 4345 4730
rect 4365 4704 4377 4716
rect 4394 4662 4406 4674
rect 4514 4721 4526 4733
rect 4493 4701 4505 4713
rect 4374 4648 4386 4660
rect 4349 4616 4361 4628
rect 4371 4616 4383 4628
rect 4414 4661 4426 4673
rect 4534 4701 4546 4713
rect 4554 4661 4566 4673
rect 4614 4647 4626 4659
rect 4734 4681 4746 4693
rect 4714 4661 4726 4673
rect 4793 4701 4805 4713
rect 4754 4647 4766 4659
rect 4834 4681 4846 4693
rect 4874 4681 4886 4693
rect 4914 4667 4926 4679
rect 4954 4667 4966 4679
rect 4994 4667 5006 4679
rect 5034 4667 5046 4679
rect 5094 4667 5106 4679
rect 5154 4681 5166 4693
rect 5134 4667 5146 4679
rect 5213 4701 5225 4713
rect 5174 4647 5186 4659
rect 5275 4681 5287 4693
rect 5354 4681 5366 4693
rect 5298 4647 5310 4659
rect 5334 4647 5346 4659
rect 5374 4667 5386 4679
rect 5414 4667 5426 4679
rect 5474 4667 5486 4679
rect 5554 4721 5566 4733
rect 5534 4701 5546 4713
rect 5514 4667 5526 4679
rect 5575 4701 5587 4713
rect 5654 4667 5666 4679
rect 5734 4721 5746 4733
rect 5714 4701 5726 4713
rect 5694 4667 5706 4679
rect 5755 4701 5767 4713
rect 5894 4721 5906 4733
rect 5874 4701 5886 4713
rect 5854 4661 5866 4673
rect 5915 4701 5927 4713
rect 6054 4681 6066 4693
rect 6074 4681 6086 4693
rect 6014 4667 6026 4679
rect 6013 4630 6025 4642
rect 6133 4701 6145 4713
rect 6094 4647 6106 4659
rect 6194 4667 6206 4679
rect 6234 4667 6246 4679
rect 6274 4661 6286 4673
rect 6254 4647 6266 4659
rect 6374 4721 6386 4733
rect 6354 4701 6366 4713
rect 6294 4647 6306 4659
rect 6395 4701 6407 4713
rect 6614 4721 6626 4733
rect 6593 4701 6605 4713
rect 6534 4681 6546 4693
rect 6494 4667 6506 4679
rect 6493 4630 6505 4642
rect 6634 4701 6646 4713
rect 54 4467 66 4479
rect 194 4467 206 4479
rect 94 4447 106 4459
rect 134 4447 146 4459
rect 234 4481 246 4493
rect 214 4447 226 4459
rect 414 4481 426 4493
rect 334 4447 346 4459
rect 273 4427 285 4439
rect 374 4447 386 4459
rect 394 4447 406 4459
rect 494 4467 506 4479
rect 453 4427 465 4439
rect 533 4496 545 4508
rect 594 4481 606 4493
rect 514 4447 526 4459
rect 634 4481 646 4493
rect 614 4467 626 4479
rect 533 4429 545 4441
rect 734 4467 746 4479
rect 834 4467 846 4479
rect 754 4447 766 4459
rect 794 4447 806 4459
rect 974 4467 986 4479
rect 894 4447 906 4459
rect 934 4447 946 4459
rect 1054 4481 1066 4493
rect 1090 4484 1102 4496
rect 1130 4484 1142 4496
rect 1170 4484 1182 4496
rect 1263 4498 1275 4510
rect 1234 4447 1246 4459
rect 1354 4467 1366 4479
rect 1263 4430 1275 4442
rect 1474 4461 1486 4473
rect 1394 4447 1406 4459
rect 1434 4447 1446 4459
rect 1514 4461 1526 4473
rect 1534 4461 1546 4473
rect 1574 4461 1586 4473
rect 1754 4467 1766 4479
rect 1797 4512 1809 4524
rect 1819 4512 1831 4524
rect 1794 4480 1806 4492
rect 1694 4447 1706 4459
rect 1774 4466 1786 4478
rect 1803 4424 1815 4436
rect 1835 4410 1847 4422
rect 1821 4390 1833 4402
rect 1867 4508 1879 4520
rect 1921 4475 1933 4487
rect 1974 4461 1986 4473
rect 1935 4436 1947 4448
rect 1883 4404 1895 4416
rect 1855 4390 1867 4402
rect 1907 4404 1919 4416
rect 2014 4461 2026 4473
rect 2087 4475 2099 4487
rect 2073 4436 2085 4448
rect 2141 4508 2153 4520
rect 2101 4404 2113 4416
rect 2125 4404 2137 4416
rect 2189 4512 2201 4524
rect 2211 4512 2223 4524
rect 2173 4410 2185 4422
rect 2153 4390 2165 4402
rect 2214 4480 2226 4492
rect 2234 4466 2246 4478
rect 2254 4467 2266 4479
rect 2294 4467 2306 4479
rect 2205 4424 2217 4436
rect 2187 4390 2199 4402
rect 2514 4467 2526 4479
rect 2354 4447 2366 4459
rect 2394 4447 2406 4459
rect 2434 4447 2446 4459
rect 2474 4447 2486 4459
rect 2607 4475 2619 4487
rect 2593 4436 2605 4448
rect 2661 4508 2673 4520
rect 2621 4404 2633 4416
rect 2645 4404 2657 4416
rect 2709 4512 2721 4524
rect 2731 4512 2743 4524
rect 2693 4410 2705 4422
rect 2673 4390 2685 4402
rect 2734 4480 2746 4492
rect 2754 4466 2766 4478
rect 2774 4467 2786 4479
rect 2725 4424 2737 4436
rect 2707 4390 2719 4402
rect 2834 4481 2846 4493
rect 2814 4447 2826 4459
rect 2914 4461 2926 4473
rect 2873 4427 2885 4439
rect 2954 4461 2966 4473
rect 3034 4467 3046 4479
rect 3074 4481 3086 4493
rect 3054 4447 3066 4459
rect 3187 4475 3199 4487
rect 3113 4427 3125 4439
rect 3173 4436 3185 4448
rect 3241 4508 3253 4520
rect 3201 4404 3213 4416
rect 3225 4404 3237 4416
rect 3289 4512 3301 4524
rect 3311 4512 3323 4524
rect 3273 4410 3285 4422
rect 3253 4390 3265 4402
rect 3314 4480 3326 4492
rect 3334 4466 3346 4478
rect 3354 4467 3366 4479
rect 3305 4424 3317 4436
rect 3287 4390 3299 4402
rect 3414 4481 3426 4493
rect 3394 4447 3406 4459
rect 3554 4481 3566 4493
rect 3453 4427 3465 4439
rect 3515 4427 3527 4439
rect 3614 4467 3626 4479
rect 3657 4512 3669 4524
rect 3679 4512 3691 4524
rect 3654 4480 3666 4492
rect 3574 4447 3586 4459
rect 3634 4466 3646 4478
rect 3663 4424 3675 4436
rect 3695 4410 3707 4422
rect 3681 4390 3693 4402
rect 3727 4508 3739 4520
rect 3781 4475 3793 4487
rect 3854 4481 3866 4493
rect 3795 4436 3807 4448
rect 3834 4447 3846 4459
rect 3954 4467 3966 4479
rect 3997 4512 4009 4524
rect 4019 4512 4031 4524
rect 3994 4480 4006 4492
rect 3893 4427 3905 4439
rect 3743 4404 3755 4416
rect 3715 4390 3727 4402
rect 3767 4404 3779 4416
rect 3974 4466 3986 4478
rect 4003 4424 4015 4436
rect 4035 4410 4047 4422
rect 4021 4390 4033 4402
rect 4067 4508 4079 4520
rect 4121 4475 4133 4487
rect 4135 4436 4147 4448
rect 4213 4427 4225 4439
rect 4083 4404 4095 4416
rect 4055 4390 4067 4402
rect 4107 4404 4119 4416
rect 4294 4481 4306 4493
rect 4274 4447 4286 4459
rect 4254 4427 4266 4439
rect 4234 4407 4246 4419
rect 4494 4481 4506 4493
rect 4394 4447 4406 4459
rect 4333 4427 4345 4439
rect 4434 4447 4446 4459
rect 4534 4481 4546 4493
rect 4514 4467 4526 4479
rect 4554 4427 4566 4439
rect 4694 4467 4706 4479
rect 4595 4427 4607 4439
rect 4574 4407 4586 4419
rect 4734 4481 4746 4493
rect 4714 4447 4726 4459
rect 4855 4496 4867 4508
rect 4894 4467 4906 4479
rect 4874 4447 4886 4459
rect 4773 4427 4785 4439
rect 4855 4429 4867 4441
rect 4934 4461 4946 4473
rect 4974 4461 4986 4473
rect 5033 4427 5045 4439
rect 5114 4481 5126 4493
rect 5094 4447 5106 4459
rect 5074 4427 5086 4439
rect 5054 4407 5066 4419
rect 5235 4496 5247 4508
rect 5274 4467 5286 4479
rect 5254 4447 5266 4459
rect 5153 4427 5165 4439
rect 5235 4429 5247 4441
rect 5314 4481 5326 4493
rect 5294 4447 5306 4459
rect 5394 4467 5406 4479
rect 5353 4427 5365 4439
rect 5493 4427 5505 4439
rect 5554 4461 5566 4473
rect 5534 4427 5546 4439
rect 5514 4407 5526 4419
rect 5594 4461 5606 4473
rect 5654 4481 5666 4493
rect 5634 4447 5646 4459
rect 5754 4461 5766 4473
rect 5693 4427 5705 4439
rect 5794 4461 5806 4473
rect 5853 4427 5865 4439
rect 5974 4481 5986 4493
rect 5894 4427 5906 4439
rect 5935 4427 5947 4439
rect 5874 4407 5886 4419
rect 6014 4467 6026 4479
rect 5994 4447 6006 4459
rect 6114 4467 6126 4479
rect 6134 4427 6146 4439
rect 6294 4481 6306 4493
rect 6175 4427 6187 4439
rect 6255 4427 6267 4439
rect 6154 4407 6166 4419
rect 6314 4447 6326 4459
rect 6334 4427 6346 4439
rect 6375 4427 6387 4439
rect 6434 4427 6446 4439
rect 6354 4407 6366 4419
rect 6554 4481 6566 4493
rect 6534 4447 6546 4459
rect 6475 4427 6487 4439
rect 6454 4407 6466 4419
rect 6634 4467 6646 4479
rect 6593 4427 6605 4439
rect 45 4218 57 4230
rect 115 4221 127 4233
rect 74 4201 86 4213
rect 45 4150 57 4162
rect 174 4201 186 4213
rect 194 4201 206 4213
rect 154 4167 166 4179
rect 253 4221 265 4233
rect 214 4167 226 4179
rect 381 4258 393 4270
rect 363 4224 375 4236
rect 314 4181 326 4193
rect 334 4182 346 4194
rect 354 4168 366 4180
rect 415 4258 427 4270
rect 395 4238 407 4250
rect 357 4136 369 4148
rect 379 4136 391 4148
rect 443 4244 455 4256
rect 467 4244 479 4256
rect 427 4140 439 4152
rect 495 4212 507 4224
rect 481 4173 493 4185
rect 534 4187 546 4199
rect 634 4201 646 4213
rect 574 4187 586 4199
rect 713 4201 725 4213
rect 655 4167 667 4179
rect 693 4167 705 4179
rect 841 4244 853 4256
rect 893 4258 905 4270
rect 865 4244 877 4256
rect 813 4212 825 4224
rect 774 4181 786 4193
rect 827 4173 839 4185
rect 881 4140 893 4152
rect 927 4258 939 4270
rect 913 4238 925 4250
rect 945 4224 957 4236
rect 974 4182 986 4194
rect 954 4168 966 4180
rect 929 4136 941 4148
rect 951 4136 963 4148
rect 994 4181 1006 4193
rect 1034 4187 1046 4199
rect 1161 4244 1173 4256
rect 1213 4258 1225 4270
rect 1185 4244 1197 4256
rect 1133 4212 1145 4224
rect 1074 4187 1086 4199
rect 1147 4173 1159 4185
rect 1201 4140 1213 4152
rect 1247 4258 1259 4270
rect 1233 4238 1245 4250
rect 1265 4224 1277 4236
rect 1294 4182 1306 4194
rect 1274 4168 1286 4180
rect 1249 4136 1261 4148
rect 1271 4136 1283 4148
rect 1314 4181 1326 4193
rect 1354 4187 1366 4199
rect 1394 4187 1406 4199
rect 1515 4221 1527 4233
rect 1434 4181 1446 4193
rect 1574 4201 1586 4213
rect 1554 4167 1566 4179
rect 1654 4181 1666 4193
rect 1634 4167 1646 4179
rect 1714 4187 1726 4199
rect 1674 4167 1686 4179
rect 1754 4187 1766 4199
rect 1774 4187 1786 4199
rect 1901 4244 1913 4256
rect 1953 4258 1965 4270
rect 1925 4244 1937 4256
rect 1873 4212 1885 4224
rect 1814 4187 1826 4199
rect 1887 4173 1899 4185
rect 1941 4140 1953 4152
rect 1987 4258 1999 4270
rect 1973 4238 1985 4250
rect 2005 4224 2017 4236
rect 2034 4182 2046 4194
rect 2014 4168 2026 4180
rect 1989 4136 2001 4148
rect 2011 4136 2023 4148
rect 2054 4181 2066 4193
rect 2094 4187 2106 4199
rect 2195 4221 2207 4233
rect 2134 4187 2146 4199
rect 2254 4201 2266 4213
rect 2234 4167 2246 4179
rect 2361 4258 2373 4270
rect 2343 4224 2355 4236
rect 2294 4181 2306 4193
rect 2314 4182 2326 4194
rect 2334 4168 2346 4180
rect 2395 4258 2407 4270
rect 2375 4238 2387 4250
rect 2337 4136 2349 4148
rect 2359 4136 2371 4148
rect 2423 4244 2435 4256
rect 2447 4244 2459 4256
rect 2407 4140 2419 4152
rect 2475 4212 2487 4224
rect 2461 4173 2473 4185
rect 2534 4201 2546 4213
rect 2574 4201 2586 4213
rect 2654 4201 2666 4213
rect 2594 4181 2606 4193
rect 2713 4221 2725 4233
rect 2674 4167 2686 4179
rect 2754 4187 2766 4199
rect 2855 4221 2867 4233
rect 2794 4187 2806 4199
rect 2914 4201 2926 4213
rect 2894 4167 2906 4179
rect 2994 4201 3006 4213
rect 3034 4201 3046 4213
rect 2934 4181 2946 4193
rect 3181 4244 3193 4256
rect 3233 4258 3245 4270
rect 3205 4244 3217 4256
rect 3153 4212 3165 4224
rect 3114 4181 3126 4193
rect 3167 4173 3179 4185
rect 3221 4140 3233 4152
rect 3267 4258 3279 4270
rect 3253 4238 3265 4250
rect 3285 4224 3297 4236
rect 3314 4182 3326 4194
rect 3374 4201 3386 4213
rect 3294 4168 3306 4180
rect 3269 4136 3281 4148
rect 3291 4136 3303 4148
rect 3334 4181 3346 4193
rect 3453 4201 3465 4213
rect 3394 4167 3406 4179
rect 3430 4167 3442 4179
rect 3494 4187 3506 4199
rect 3534 4187 3546 4199
rect 3594 4167 3606 4179
rect 3774 4187 3786 4199
rect 3630 4164 3642 4176
rect 3670 4164 3682 4176
rect 3710 4164 3722 4176
rect 3814 4187 3826 4199
rect 3854 4187 3866 4199
rect 3894 4187 3906 4199
rect 3954 4187 3966 4199
rect 3994 4187 4006 4199
rect 4095 4221 4107 4233
rect 4014 4181 4026 4193
rect 4154 4201 4166 4213
rect 4174 4201 4186 4213
rect 4134 4167 4146 4179
rect 4233 4221 4245 4233
rect 4194 4167 4206 4179
rect 4361 4258 4373 4270
rect 4343 4224 4355 4236
rect 4294 4181 4306 4193
rect 4314 4182 4326 4194
rect 4334 4168 4346 4180
rect 4395 4258 4407 4270
rect 4375 4238 4387 4250
rect 4337 4136 4349 4148
rect 4359 4136 4371 4148
rect 4423 4244 4435 4256
rect 4447 4244 4459 4256
rect 4407 4140 4419 4152
rect 4475 4212 4487 4224
rect 4535 4221 4547 4233
rect 4461 4173 4473 4185
rect 4594 4201 4606 4213
rect 4574 4167 4586 4179
rect 4701 4258 4713 4270
rect 4683 4224 4695 4236
rect 4634 4181 4646 4193
rect 4654 4182 4666 4194
rect 4674 4168 4686 4180
rect 4735 4258 4747 4270
rect 4715 4238 4727 4250
rect 4677 4136 4689 4148
rect 4699 4136 4711 4148
rect 4763 4244 4775 4256
rect 4787 4244 4799 4256
rect 4747 4140 4759 4152
rect 4815 4212 4827 4224
rect 4801 4173 4813 4185
rect 5034 4241 5046 4253
rect 5014 4221 5026 4233
rect 4974 4181 4986 4193
rect 4894 4167 4906 4179
rect 4954 4167 4966 4179
rect 4994 4167 5006 4179
rect 5055 4221 5067 4233
rect 5174 4201 5186 4213
rect 5154 4181 5166 4193
rect 5233 4221 5245 4233
rect 5194 4167 5206 4179
rect 5361 4258 5373 4270
rect 5343 4224 5355 4236
rect 5294 4181 5306 4193
rect 5314 4182 5326 4194
rect 5334 4168 5346 4180
rect 5395 4258 5407 4270
rect 5375 4238 5387 4250
rect 5337 4136 5349 4148
rect 5359 4136 5371 4148
rect 5423 4244 5435 4256
rect 5447 4244 5459 4256
rect 5407 4140 5419 4152
rect 5475 4212 5487 4224
rect 5461 4173 5473 4185
rect 5514 4187 5526 4199
rect 5554 4187 5566 4199
rect 5654 4201 5666 4213
rect 5594 4181 5606 4193
rect 5713 4221 5725 4233
rect 5674 4167 5686 4179
rect 5874 4241 5886 4253
rect 5854 4221 5866 4233
rect 5834 4201 5846 4213
rect 5794 4187 5806 4199
rect 5793 4150 5805 4162
rect 5895 4221 5907 4233
rect 6014 4201 6026 4213
rect 5994 4167 6006 4179
rect 6073 4221 6085 4233
rect 6034 4167 6046 4179
rect 6143 4218 6155 4230
rect 6114 4201 6126 4213
rect 6194 4187 6206 4199
rect 6234 4187 6246 4199
rect 6143 4150 6155 4162
rect 6354 4201 6366 4213
rect 6314 4187 6326 4199
rect 6313 4150 6325 4162
rect 6374 4187 6386 4199
rect 6414 4187 6426 4199
rect 6454 4181 6466 4193
rect 6634 4241 6646 4253
rect 6614 4221 6626 4233
rect 6574 4181 6586 4193
rect 6554 4167 6566 4179
rect 6594 4167 6606 4179
rect 6655 4221 6667 4233
rect 45 4018 57 4030
rect 74 3967 86 3979
rect 127 3995 139 4007
rect 45 3950 57 3962
rect 113 3956 125 3968
rect 181 4028 193 4040
rect 141 3924 153 3936
rect 165 3924 177 3936
rect 229 4032 241 4044
rect 251 4032 263 4044
rect 213 3930 225 3942
rect 193 3910 205 3922
rect 254 4000 266 4012
rect 274 3986 286 3998
rect 294 3987 306 3999
rect 245 3944 257 3956
rect 227 3910 239 3922
rect 334 3981 346 3993
rect 454 4001 466 4013
rect 374 3981 386 3993
rect 494 4001 506 4013
rect 474 3987 486 3999
rect 534 3981 546 3993
rect 705 4018 717 4030
rect 574 3981 586 3993
rect 614 3981 626 3993
rect 654 3981 666 3993
rect 734 3967 746 3979
rect 787 3995 799 4007
rect 705 3950 717 3962
rect 773 3956 785 3968
rect 841 4028 853 4040
rect 801 3924 813 3936
rect 825 3924 837 3936
rect 889 4032 901 4044
rect 911 4032 923 4044
rect 873 3930 885 3942
rect 853 3910 865 3922
rect 914 4000 926 4012
rect 934 3986 946 3998
rect 954 3987 966 3999
rect 905 3944 917 3956
rect 887 3910 899 3922
rect 1014 3981 1026 3993
rect 1054 3981 1066 3993
rect 1074 3981 1086 3993
rect 1114 3981 1126 3993
rect 1154 3981 1166 3993
rect 1274 4001 1286 4013
rect 1194 3981 1206 3993
rect 1314 4001 1326 4013
rect 1294 3987 1306 3999
rect 1367 3995 1379 4007
rect 1353 3956 1365 3968
rect 1421 4028 1433 4040
rect 1381 3924 1393 3936
rect 1405 3924 1417 3936
rect 1469 4032 1481 4044
rect 1491 4032 1503 4044
rect 1453 3930 1465 3942
rect 1433 3910 1445 3922
rect 1494 4000 1506 4012
rect 1514 3986 1526 3998
rect 1534 3987 1546 3999
rect 1485 3944 1497 3956
rect 1467 3910 1479 3922
rect 1594 3981 1606 3993
rect 1634 3981 1646 3993
rect 1683 4018 1695 4030
rect 1734 3981 1746 3993
rect 1654 3967 1666 3979
rect 1683 3950 1695 3962
rect 1774 3981 1786 3993
rect 1847 3995 1859 4007
rect 1833 3956 1845 3968
rect 1901 4028 1913 4040
rect 1861 3924 1873 3936
rect 1885 3924 1897 3936
rect 1949 4032 1961 4044
rect 1971 4032 1983 4044
rect 1933 3930 1945 3942
rect 1913 3910 1925 3922
rect 1974 4000 1986 4012
rect 1994 3986 2006 3998
rect 2014 3987 2026 3999
rect 1965 3944 1977 3956
rect 1947 3910 1959 3922
rect 2054 3981 2066 3993
rect 2094 3981 2106 3993
rect 2194 4001 2206 4013
rect 2155 3947 2167 3959
rect 2254 3981 2266 3993
rect 2214 3967 2226 3979
rect 2294 3981 2306 3993
rect 2314 3981 2326 3993
rect 2354 3981 2366 3993
rect 2434 3987 2446 3999
rect 2514 4001 2526 4013
rect 2475 3947 2487 3959
rect 2714 3987 2726 3999
rect 2534 3967 2546 3979
rect 2554 3967 2566 3979
rect 2594 3967 2606 3979
rect 2654 3967 2666 3979
rect 2694 3967 2706 3979
rect 2814 3987 2826 3999
rect 2854 3981 2866 3993
rect 2894 3981 2906 3993
rect 3014 4001 3026 4013
rect 2914 3967 2926 3979
rect 2954 3967 2966 3979
rect 2994 3967 3006 3979
rect 3094 3987 3106 3999
rect 3053 3947 3065 3959
rect 3254 3981 3266 3993
rect 3154 3967 3166 3979
rect 3194 3967 3206 3979
rect 3294 3981 3306 3993
rect 3334 3981 3346 3993
rect 3374 3981 3386 3993
rect 3414 3987 3426 3999
rect 3457 4032 3469 4044
rect 3479 4032 3491 4044
rect 3454 4000 3466 4012
rect 3434 3986 3446 3998
rect 3463 3944 3475 3956
rect 3495 3930 3507 3942
rect 3481 3910 3493 3922
rect 3527 4028 3539 4040
rect 3581 3995 3593 4007
rect 3595 3956 3607 3968
rect 3674 3987 3686 3999
rect 3714 3987 3726 3999
rect 3757 4032 3769 4044
rect 3779 4032 3791 4044
rect 3754 4000 3766 4012
rect 3543 3924 3555 3936
rect 3515 3910 3527 3922
rect 3567 3924 3579 3936
rect 3734 3986 3746 3998
rect 3763 3944 3775 3956
rect 3795 3930 3807 3942
rect 3781 3910 3793 3922
rect 3827 4028 3839 4040
rect 3881 3995 3893 4007
rect 3895 3956 3907 3968
rect 3973 3947 3985 3959
rect 3843 3924 3855 3936
rect 3815 3910 3827 3922
rect 3867 3924 3879 3936
rect 4034 3981 4046 3993
rect 4014 3947 4026 3959
rect 3994 3927 4006 3939
rect 4074 3981 4086 3993
rect 4174 4001 4186 4013
rect 4135 3947 4147 3959
rect 4334 3987 4346 3999
rect 4194 3967 4206 3979
rect 4214 3967 4226 3979
rect 4254 3967 4266 3979
rect 4374 3981 4386 3993
rect 4414 3981 4426 3993
rect 4494 4001 4506 4013
rect 4455 3947 4467 3959
rect 4554 3987 4566 3999
rect 4597 4032 4609 4044
rect 4619 4032 4631 4044
rect 4594 4000 4606 4012
rect 4514 3967 4526 3979
rect 4574 3986 4586 3998
rect 4603 3944 4615 3956
rect 4635 3930 4647 3942
rect 4621 3910 4633 3922
rect 4667 4028 4679 4040
rect 4721 3995 4733 4007
rect 4794 3981 4806 3993
rect 4735 3956 4747 3968
rect 4683 3924 4695 3936
rect 4655 3910 4667 3922
rect 4707 3924 4719 3936
rect 4834 3981 4846 3993
rect 4914 4001 4926 4013
rect 4875 3947 4887 3959
rect 4974 3987 4986 3999
rect 5017 4032 5029 4044
rect 5039 4032 5051 4044
rect 5014 4000 5026 4012
rect 4934 3967 4946 3979
rect 4994 3986 5006 3998
rect 5023 3944 5035 3956
rect 5055 3930 5067 3942
rect 5041 3910 5053 3922
rect 5087 4028 5099 4040
rect 5141 3995 5153 4007
rect 5214 3981 5226 3993
rect 5155 3956 5167 3968
rect 5103 3924 5115 3936
rect 5075 3910 5087 3922
rect 5127 3924 5139 3936
rect 5254 3981 5266 3993
rect 5334 4001 5346 4013
rect 5295 3947 5307 3959
rect 5394 3981 5406 3993
rect 5354 3967 5366 3979
rect 5434 3981 5446 3993
rect 5474 4001 5486 4013
rect 5454 3967 5466 3979
rect 5594 3987 5606 3999
rect 5634 3987 5646 3999
rect 5677 4032 5689 4044
rect 5699 4032 5711 4044
rect 5674 4000 5686 4012
rect 5513 3947 5525 3959
rect 5654 3986 5666 3998
rect 5683 3944 5695 3956
rect 5715 3930 5727 3942
rect 5701 3910 5713 3922
rect 5747 4028 5759 4040
rect 5801 3995 5813 4007
rect 5854 3987 5866 3999
rect 5815 3956 5827 3968
rect 5763 3924 5775 3936
rect 5735 3910 5747 3922
rect 5787 3924 5799 3936
rect 5953 3947 5965 3959
rect 6047 3995 6059 4007
rect 5994 3947 6006 3959
rect 6033 3956 6045 3968
rect 5974 3927 5986 3939
rect 6101 4028 6113 4040
rect 6061 3924 6073 3936
rect 6085 3924 6097 3936
rect 6149 4032 6161 4044
rect 6171 4032 6183 4044
rect 6133 3930 6145 3942
rect 6113 3910 6125 3922
rect 6174 4000 6186 4012
rect 6194 3986 6206 3998
rect 6214 3987 6226 3999
rect 6165 3944 6177 3956
rect 6147 3910 6159 3922
rect 6287 3995 6299 4007
rect 6273 3956 6285 3968
rect 6341 4028 6353 4040
rect 6301 3924 6313 3936
rect 6325 3924 6337 3936
rect 6389 4032 6401 4044
rect 6411 4032 6423 4044
rect 6373 3930 6385 3942
rect 6353 3910 6365 3922
rect 6414 4000 6426 4012
rect 6434 3986 6446 3998
rect 6454 3987 6466 3999
rect 6405 3944 6417 3956
rect 6387 3910 6399 3922
rect 6527 3995 6539 4007
rect 6513 3956 6525 3968
rect 6581 4028 6593 4040
rect 6541 3924 6553 3936
rect 6565 3924 6577 3936
rect 6629 4032 6641 4044
rect 6651 4032 6663 4044
rect 6613 3930 6625 3942
rect 6593 3910 6605 3922
rect 6654 4000 6666 4012
rect 6674 3986 6686 3998
rect 6694 3987 6706 3999
rect 6645 3944 6657 3956
rect 6627 3910 6639 3922
rect 45 3738 57 3750
rect 125 3738 137 3750
rect 74 3721 86 3733
rect 154 3721 166 3733
rect 45 3670 57 3682
rect 125 3670 137 3682
rect 194 3707 206 3719
rect 301 3764 313 3776
rect 353 3778 365 3790
rect 325 3764 337 3776
rect 273 3732 285 3744
rect 234 3707 246 3719
rect 287 3693 299 3705
rect 341 3660 353 3672
rect 387 3778 399 3790
rect 373 3758 385 3770
rect 405 3744 417 3756
rect 434 3702 446 3714
rect 414 3688 426 3700
rect 389 3656 401 3668
rect 411 3656 423 3668
rect 454 3701 466 3713
rect 554 3701 566 3713
rect 534 3687 546 3699
rect 614 3707 626 3719
rect 574 3687 586 3699
rect 654 3707 666 3719
rect 674 3707 686 3719
rect 714 3707 726 3719
rect 774 3707 786 3719
rect 881 3764 893 3776
rect 933 3778 945 3790
rect 905 3764 917 3776
rect 853 3732 865 3744
rect 814 3707 826 3719
rect 867 3693 879 3705
rect 921 3660 933 3672
rect 967 3778 979 3790
rect 953 3758 965 3770
rect 985 3744 997 3756
rect 1014 3702 1026 3714
rect 994 3688 1006 3700
rect 969 3656 981 3668
rect 991 3656 1003 3668
rect 1034 3701 1046 3713
rect 1094 3701 1106 3713
rect 1074 3687 1086 3699
rect 1194 3707 1206 3719
rect 1114 3687 1126 3699
rect 1283 3738 1295 3750
rect 1254 3721 1266 3733
rect 1234 3707 1246 3719
rect 1394 3701 1406 3713
rect 1374 3687 1386 3699
rect 1283 3670 1295 3682
rect 1454 3707 1466 3719
rect 1414 3687 1426 3699
rect 1494 3707 1506 3719
rect 1514 3707 1526 3719
rect 1721 3764 1733 3776
rect 1773 3778 1785 3790
rect 1745 3764 1757 3776
rect 1594 3721 1606 3733
rect 1634 3721 1646 3733
rect 1693 3732 1705 3744
rect 1554 3707 1566 3719
rect 1707 3693 1719 3705
rect 1761 3660 1773 3672
rect 1807 3778 1819 3790
rect 1793 3758 1805 3770
rect 1825 3744 1837 3756
rect 1854 3702 1866 3714
rect 1834 3688 1846 3700
rect 1809 3656 1821 3668
rect 1831 3656 1843 3668
rect 1874 3701 1886 3713
rect 1934 3707 1946 3719
rect 1994 3721 2006 3733
rect 2034 3721 2046 3733
rect 1974 3707 1986 3719
rect 2134 3721 2146 3733
rect 2074 3701 2086 3713
rect 2193 3741 2205 3753
rect 2255 3741 2267 3753
rect 2154 3687 2166 3699
rect 2314 3721 2326 3733
rect 2294 3687 2306 3699
rect 2394 3701 2406 3713
rect 2374 3687 2386 3699
rect 2434 3701 2446 3713
rect 2414 3687 2426 3699
rect 2554 3721 2566 3733
rect 2534 3701 2546 3713
rect 2674 3761 2686 3773
rect 2613 3741 2625 3753
rect 2654 3741 2666 3753
rect 2574 3687 2586 3699
rect 2695 3741 2707 3753
rect 2794 3701 2806 3713
rect 2834 3707 2846 3719
rect 2894 3721 2906 3733
rect 2874 3707 2886 3719
rect 2953 3741 2965 3753
rect 2914 3687 2926 3699
rect 2994 3721 3006 3733
rect 3053 3741 3065 3753
rect 3014 3687 3026 3699
rect 3114 3701 3126 3713
rect 3094 3687 3106 3699
rect 3214 3721 3226 3733
rect 3134 3687 3146 3699
rect 3293 3721 3305 3733
rect 3235 3687 3247 3699
rect 3273 3687 3285 3699
rect 3334 3707 3346 3719
rect 3374 3707 3386 3719
rect 3414 3707 3426 3719
rect 3454 3707 3466 3719
rect 3561 3778 3573 3790
rect 3543 3744 3555 3756
rect 3494 3701 3506 3713
rect 3514 3702 3526 3714
rect 3534 3688 3546 3700
rect 3595 3778 3607 3790
rect 3575 3758 3587 3770
rect 3537 3656 3549 3668
rect 3559 3656 3571 3668
rect 3623 3764 3635 3776
rect 3647 3764 3659 3776
rect 3607 3660 3619 3672
rect 3675 3732 3687 3744
rect 3661 3693 3673 3705
rect 3734 3707 3746 3719
rect 3814 3721 3826 3733
rect 3774 3707 3786 3719
rect 3893 3721 3905 3733
rect 3835 3687 3847 3699
rect 3873 3687 3885 3699
rect 3914 3701 3926 3713
rect 3974 3707 3986 3719
rect 4054 3721 4066 3733
rect 4014 3707 4026 3719
rect 4113 3741 4125 3753
rect 4074 3687 4086 3699
rect 4241 3778 4253 3790
rect 4223 3744 4235 3756
rect 4174 3701 4186 3713
rect 4194 3702 4206 3714
rect 4214 3688 4226 3700
rect 4275 3778 4287 3790
rect 4255 3758 4267 3770
rect 4217 3656 4229 3668
rect 4239 3656 4251 3668
rect 4303 3764 4315 3776
rect 4327 3764 4339 3776
rect 4287 3660 4299 3672
rect 4355 3732 4367 3744
rect 4341 3693 4353 3705
rect 4394 3707 4406 3719
rect 4434 3707 4446 3719
rect 4494 3707 4506 3719
rect 4534 3707 4546 3719
rect 4841 3778 4853 3790
rect 4823 3744 4835 3756
rect 4774 3701 4786 3713
rect 4794 3702 4806 3714
rect 4598 3684 4610 3696
rect 4638 3684 4650 3696
rect 4678 3684 4690 3696
rect 4714 3687 4726 3699
rect 4814 3688 4826 3700
rect 4875 3778 4887 3790
rect 4855 3758 4867 3770
rect 4817 3656 4829 3668
rect 4839 3656 4851 3668
rect 4903 3764 4915 3776
rect 4927 3764 4939 3776
rect 4887 3660 4899 3672
rect 4955 3732 4967 3744
rect 4941 3693 4953 3705
rect 4994 3721 5006 3733
rect 5053 3741 5065 3753
rect 5014 3687 5026 3699
rect 5114 3707 5126 3719
rect 5154 3707 5166 3719
rect 5194 3707 5206 3719
rect 5234 3707 5246 3719
rect 5561 3764 5573 3776
rect 5613 3778 5625 3790
rect 5585 3764 5597 3776
rect 5294 3701 5306 3713
rect 5334 3687 5346 3699
rect 5370 3684 5382 3696
rect 5410 3684 5422 3696
rect 5450 3684 5462 3696
rect 5533 3732 5545 3744
rect 5547 3693 5559 3705
rect 5601 3660 5613 3672
rect 5647 3778 5659 3790
rect 5633 3758 5645 3770
rect 5665 3744 5677 3756
rect 5694 3702 5706 3714
rect 5674 3688 5686 3700
rect 5649 3656 5661 3668
rect 5671 3656 5683 3668
rect 5714 3701 5726 3713
rect 5794 3701 5806 3713
rect 5814 3707 5826 3719
rect 5854 3707 5866 3719
rect 5894 3707 5906 3719
rect 5934 3707 5946 3719
rect 6341 3764 6353 3776
rect 6393 3778 6405 3790
rect 6365 3764 6377 3776
rect 6034 3721 6046 3733
rect 6074 3721 6086 3733
rect 6134 3721 6146 3733
rect 6174 3721 6186 3733
rect 6014 3701 6026 3713
rect 6214 3701 6226 3713
rect 6194 3687 6206 3699
rect 6234 3687 6246 3699
rect 6313 3732 6325 3744
rect 6327 3693 6339 3705
rect 6381 3660 6393 3672
rect 6427 3778 6439 3790
rect 6413 3758 6425 3770
rect 6445 3744 6457 3756
rect 6474 3702 6486 3714
rect 6534 3721 6546 3733
rect 6454 3688 6466 3700
rect 6429 3656 6441 3668
rect 6451 3656 6463 3668
rect 6494 3701 6506 3713
rect 6593 3741 6605 3753
rect 6554 3687 6566 3699
rect 6634 3707 6646 3719
rect 6674 3707 6686 3719
rect 45 3538 57 3550
rect 74 3487 86 3499
rect 127 3515 139 3527
rect 45 3470 57 3482
rect 113 3476 125 3488
rect 181 3548 193 3560
rect 141 3444 153 3456
rect 165 3444 177 3456
rect 229 3552 241 3564
rect 251 3552 263 3564
rect 213 3450 225 3462
rect 193 3430 205 3442
rect 254 3520 266 3532
rect 274 3506 286 3518
rect 294 3507 306 3519
rect 245 3464 257 3476
rect 227 3430 239 3442
rect 334 3501 346 3513
rect 374 3501 386 3513
rect 443 3538 455 3550
rect 414 3487 426 3499
rect 534 3521 546 3533
rect 443 3470 455 3482
rect 574 3521 586 3533
rect 705 3538 717 3550
rect 554 3507 566 3519
rect 614 3501 626 3513
rect 654 3501 666 3513
rect 783 3538 795 3550
rect 945 3538 957 3550
rect 834 3501 846 3513
rect 734 3487 746 3499
rect 754 3487 766 3499
rect 705 3470 717 3482
rect 783 3470 795 3482
rect 874 3501 886 3513
rect 1085 3538 1097 3550
rect 1034 3507 1046 3519
rect 974 3487 986 3499
rect 945 3470 957 3482
rect 1165 3538 1177 3550
rect 1114 3487 1126 3499
rect 1194 3487 1206 3499
rect 1247 3515 1259 3527
rect 1085 3470 1097 3482
rect 1165 3470 1177 3482
rect 1233 3476 1245 3488
rect 1301 3548 1313 3560
rect 1261 3444 1273 3456
rect 1285 3444 1297 3456
rect 1349 3552 1361 3564
rect 1371 3552 1383 3564
rect 1333 3450 1345 3462
rect 1313 3430 1325 3442
rect 1374 3520 1386 3532
rect 1394 3506 1406 3518
rect 1414 3507 1426 3519
rect 1365 3464 1377 3476
rect 1347 3430 1359 3442
rect 1474 3487 1486 3499
rect 1514 3487 1526 3499
rect 1567 3515 1579 3527
rect 1553 3476 1565 3488
rect 1621 3548 1633 3560
rect 1581 3444 1593 3456
rect 1605 3444 1617 3456
rect 1669 3552 1681 3564
rect 1691 3552 1703 3564
rect 1653 3450 1665 3462
rect 1633 3430 1645 3442
rect 1694 3520 1706 3532
rect 1813 3538 1825 3550
rect 1714 3506 1726 3518
rect 1734 3507 1746 3519
rect 1685 3464 1697 3476
rect 1667 3430 1679 3442
rect 1814 3501 1826 3513
rect 1914 3507 1926 3519
rect 1854 3487 1866 3499
rect 1994 3521 2006 3533
rect 1955 3467 1967 3479
rect 2213 3538 2225 3550
rect 2154 3507 2166 3519
rect 2014 3487 2026 3499
rect 2034 3487 2046 3499
rect 2074 3487 2086 3499
rect 2214 3501 2226 3513
rect 2254 3487 2266 3499
rect 2294 3487 2306 3499
rect 2334 3487 2346 3499
rect 2387 3515 2399 3527
rect 2373 3476 2385 3488
rect 2441 3548 2453 3560
rect 2401 3444 2413 3456
rect 2425 3444 2437 3456
rect 2489 3552 2501 3564
rect 2511 3552 2523 3564
rect 2473 3450 2485 3462
rect 2453 3430 2465 3442
rect 2514 3520 2526 3532
rect 2534 3506 2546 3518
rect 2554 3507 2566 3519
rect 2505 3464 2517 3476
rect 2487 3430 2499 3442
rect 2694 3521 2706 3533
rect 2594 3487 2606 3499
rect 2634 3487 2646 3499
rect 2674 3487 2686 3499
rect 2814 3507 2826 3519
rect 2733 3467 2745 3479
rect 2854 3501 2866 3513
rect 2894 3501 2906 3513
rect 2934 3521 2946 3533
rect 2914 3487 2926 3499
rect 3014 3521 3026 3533
rect 3054 3521 3066 3533
rect 3114 3521 3126 3533
rect 3034 3507 3046 3519
rect 2973 3467 2985 3479
rect 3215 3521 3227 3533
rect 3253 3521 3265 3533
rect 3194 3487 3206 3499
rect 3334 3507 3346 3519
rect 3273 3487 3285 3499
rect 3387 3515 3399 3527
rect 3373 3476 3385 3488
rect 3441 3548 3453 3560
rect 3401 3444 3413 3456
rect 3425 3444 3437 3456
rect 3489 3552 3501 3564
rect 3511 3552 3523 3564
rect 3473 3450 3485 3462
rect 3453 3430 3465 3442
rect 3514 3520 3526 3532
rect 3534 3506 3546 3518
rect 3554 3507 3566 3519
rect 3505 3464 3517 3476
rect 3487 3430 3499 3442
rect 3635 3521 3647 3533
rect 3673 3521 3685 3533
rect 3614 3487 3626 3499
rect 3693 3487 3705 3499
rect 3747 3515 3759 3527
rect 3733 3476 3745 3488
rect 3801 3548 3813 3560
rect 3761 3444 3773 3456
rect 3785 3444 3797 3456
rect 3849 3552 3861 3564
rect 3871 3552 3883 3564
rect 3833 3450 3845 3462
rect 3813 3430 3825 3442
rect 3874 3520 3886 3532
rect 3894 3506 3906 3518
rect 3914 3507 3926 3519
rect 3994 3507 4006 3519
rect 3865 3464 3877 3476
rect 3847 3430 3859 3442
rect 4047 3515 4059 3527
rect 4033 3476 4045 3488
rect 4101 3548 4113 3560
rect 4061 3444 4073 3456
rect 4085 3444 4097 3456
rect 4149 3552 4161 3564
rect 4171 3552 4183 3564
rect 4133 3450 4145 3462
rect 4113 3430 4125 3442
rect 4174 3520 4186 3532
rect 4194 3506 4206 3518
rect 4214 3507 4226 3519
rect 4294 3507 4306 3519
rect 4354 3507 4366 3519
rect 4165 3464 4177 3476
rect 4147 3430 4159 3442
rect 4374 3501 4386 3513
rect 4414 3501 4426 3513
rect 4474 3507 4486 3519
rect 4517 3552 4529 3564
rect 4539 3552 4551 3564
rect 4514 3520 4526 3532
rect 4494 3506 4506 3518
rect 4523 3464 4535 3476
rect 4555 3450 4567 3462
rect 4541 3430 4553 3442
rect 4587 3548 4599 3560
rect 4641 3515 4653 3527
rect 4655 3476 4667 3488
rect 4734 3507 4746 3519
rect 4603 3444 4615 3456
rect 4575 3430 4587 3442
rect 4627 3444 4639 3456
rect 4787 3515 4799 3527
rect 4773 3476 4785 3488
rect 4841 3548 4853 3560
rect 4801 3444 4813 3456
rect 4825 3444 4837 3456
rect 4889 3552 4901 3564
rect 4911 3552 4923 3564
rect 4873 3450 4885 3462
rect 4853 3430 4865 3442
rect 4914 3520 4926 3532
rect 4934 3506 4946 3518
rect 4954 3507 4966 3519
rect 4905 3464 4917 3476
rect 4887 3430 4899 3442
rect 5035 3521 5047 3533
rect 5073 3521 5085 3533
rect 5014 3487 5026 3499
rect 5154 3507 5166 3519
rect 5093 3487 5105 3499
rect 5207 3515 5219 3527
rect 5193 3476 5205 3488
rect 5261 3548 5273 3560
rect 5221 3444 5233 3456
rect 5245 3444 5257 3456
rect 5309 3552 5321 3564
rect 5331 3552 5343 3564
rect 5293 3450 5305 3462
rect 5273 3430 5285 3442
rect 5334 3520 5346 3532
rect 5354 3506 5366 3518
rect 5374 3507 5386 3519
rect 5325 3464 5337 3476
rect 5307 3430 5319 3442
rect 5447 3515 5459 3527
rect 5433 3476 5445 3488
rect 5501 3548 5513 3560
rect 5461 3444 5473 3456
rect 5485 3444 5497 3456
rect 5549 3552 5561 3564
rect 5571 3552 5583 3564
rect 5533 3450 5545 3462
rect 5513 3430 5525 3442
rect 5574 3520 5586 3532
rect 5594 3506 5606 3518
rect 5614 3507 5626 3519
rect 5565 3464 5577 3476
rect 5547 3430 5559 3442
rect 5674 3521 5686 3533
rect 5654 3487 5666 3499
rect 5774 3521 5786 3533
rect 5754 3487 5766 3499
rect 5713 3467 5725 3479
rect 5894 3507 5906 3519
rect 5813 3467 5825 3479
rect 5955 3521 5967 3533
rect 5993 3521 6005 3533
rect 5934 3487 5946 3499
rect 6034 3501 6046 3513
rect 6013 3487 6025 3499
rect 6074 3501 6086 3513
rect 6154 3507 6166 3519
rect 6194 3487 6206 3499
rect 6234 3521 6246 3533
rect 6254 3487 6266 3499
rect 6394 3507 6406 3519
rect 6447 3515 6459 3527
rect 6433 3476 6445 3488
rect 6501 3548 6513 3560
rect 6461 3444 6473 3456
rect 6485 3444 6497 3456
rect 6549 3552 6561 3564
rect 6571 3552 6583 3564
rect 6533 3450 6545 3462
rect 6513 3430 6525 3442
rect 6574 3520 6586 3532
rect 6594 3506 6606 3518
rect 6614 3507 6626 3519
rect 6565 3464 6577 3476
rect 6547 3430 6559 3442
rect 45 3258 57 3270
rect 141 3284 153 3296
rect 193 3298 205 3310
rect 165 3284 177 3296
rect 74 3241 86 3253
rect 113 3252 125 3264
rect 45 3190 57 3202
rect 127 3213 139 3225
rect 181 3180 193 3192
rect 227 3298 239 3310
rect 213 3278 225 3290
rect 245 3264 257 3276
rect 274 3222 286 3234
rect 254 3208 266 3220
rect 229 3176 241 3188
rect 251 3176 263 3188
rect 294 3221 306 3233
rect 334 3227 346 3239
rect 374 3227 386 3239
rect 474 3221 486 3233
rect 454 3207 466 3219
rect 534 3227 546 3239
rect 494 3207 506 3219
rect 574 3227 586 3239
rect 674 3281 686 3293
rect 654 3261 666 3273
rect 594 3221 606 3233
rect 695 3261 707 3273
rect 754 3227 766 3239
rect 855 3261 867 3273
rect 794 3227 806 3239
rect 914 3241 926 3253
rect 894 3207 906 3219
rect 994 3241 1006 3253
rect 1034 3241 1046 3253
rect 1074 3241 1086 3253
rect 934 3221 946 3233
rect 1133 3261 1145 3273
rect 1094 3207 1106 3219
rect 1174 3241 1186 3253
rect 1233 3261 1245 3273
rect 1194 3207 1206 3219
rect 1274 3227 1286 3239
rect 1401 3284 1413 3296
rect 1453 3298 1465 3310
rect 1425 3284 1437 3296
rect 1373 3252 1385 3264
rect 1314 3227 1326 3239
rect 1387 3213 1399 3225
rect 1441 3180 1453 3192
rect 1487 3298 1499 3310
rect 1473 3278 1485 3290
rect 1505 3264 1517 3276
rect 1534 3222 1546 3234
rect 1514 3208 1526 3220
rect 1489 3176 1501 3188
rect 1511 3176 1523 3188
rect 1554 3221 1566 3233
rect 1674 3241 1686 3253
rect 1634 3227 1646 3239
rect 1633 3190 1645 3202
rect 1854 3281 1866 3293
rect 1833 3261 1845 3273
rect 1754 3221 1766 3233
rect 1734 3207 1746 3219
rect 1774 3207 1786 3219
rect 1874 3261 1886 3273
rect 1914 3221 1926 3233
rect 1894 3207 1906 3219
rect 2081 3298 2093 3310
rect 2063 3264 2075 3276
rect 2014 3221 2026 3233
rect 2034 3222 2046 3234
rect 1934 3207 1946 3219
rect 2054 3208 2066 3220
rect 2115 3298 2127 3310
rect 2095 3278 2107 3290
rect 2057 3176 2069 3188
rect 2079 3176 2091 3188
rect 2143 3284 2155 3296
rect 2167 3284 2179 3296
rect 2127 3180 2139 3192
rect 2195 3252 2207 3264
rect 2181 3213 2193 3225
rect 2234 3227 2246 3239
rect 2314 3241 2326 3253
rect 2354 3241 2366 3253
rect 2414 3241 2426 3253
rect 2495 3261 2507 3273
rect 2454 3241 2466 3253
rect 2274 3227 2286 3239
rect 2554 3241 2566 3253
rect 2534 3207 2546 3219
rect 2721 3298 2733 3310
rect 2703 3264 2715 3276
rect 2574 3221 2586 3233
rect 2654 3221 2666 3233
rect 2674 3222 2686 3234
rect 2694 3208 2706 3220
rect 2755 3298 2767 3310
rect 2735 3278 2747 3290
rect 2697 3176 2709 3188
rect 2719 3176 2731 3188
rect 2783 3284 2795 3296
rect 2807 3284 2819 3296
rect 2767 3180 2779 3192
rect 2835 3252 2847 3264
rect 2821 3213 2833 3225
rect 2874 3227 2886 3239
rect 2914 3227 2926 3239
rect 2974 3227 2986 3239
rect 3055 3261 3067 3273
rect 3014 3227 3026 3239
rect 3114 3241 3126 3253
rect 3094 3207 3106 3219
rect 3154 3227 3166 3239
rect 3194 3227 3206 3239
rect 3295 3261 3307 3273
rect 3254 3221 3266 3233
rect 3354 3241 3366 3253
rect 3334 3207 3346 3219
rect 3741 3284 3753 3296
rect 3793 3298 3805 3310
rect 3765 3284 3777 3296
rect 3454 3241 3466 3253
rect 3494 3241 3506 3253
rect 3374 3221 3386 3233
rect 3574 3221 3586 3233
rect 3554 3207 3566 3219
rect 3634 3241 3646 3253
rect 3674 3241 3686 3253
rect 3713 3252 3725 3264
rect 3594 3207 3606 3219
rect 3727 3213 3739 3225
rect 3781 3180 3793 3192
rect 3827 3298 3839 3310
rect 3813 3278 3825 3290
rect 3845 3264 3857 3276
rect 3874 3222 3886 3234
rect 3935 3241 3947 3253
rect 3854 3208 3866 3220
rect 3829 3176 3841 3188
rect 3851 3176 3863 3188
rect 3894 3221 3906 3233
rect 4014 3241 4026 3253
rect 4074 3241 4086 3253
rect 3955 3207 3967 3219
rect 3993 3207 4005 3219
rect 4153 3241 4165 3253
rect 4095 3207 4107 3219
rect 4133 3207 4145 3219
rect 4261 3298 4273 3310
rect 4243 3264 4255 3276
rect 4194 3221 4206 3233
rect 4214 3222 4226 3234
rect 4234 3208 4246 3220
rect 4295 3298 4307 3310
rect 4275 3278 4287 3290
rect 4237 3176 4249 3188
rect 4259 3176 4271 3188
rect 4323 3284 4335 3296
rect 4347 3284 4359 3296
rect 4307 3180 4319 3192
rect 4375 3252 4387 3264
rect 4361 3213 4373 3225
rect 4414 3241 4426 3253
rect 4454 3241 4466 3253
rect 4495 3241 4507 3253
rect 4574 3241 4586 3253
rect 4614 3241 4626 3253
rect 4654 3241 4666 3253
rect 4694 3241 4706 3253
rect 4734 3241 4746 3253
rect 4515 3207 4527 3219
rect 4553 3207 4565 3219
rect 5101 3284 5113 3296
rect 5153 3298 5165 3310
rect 5125 3284 5137 3296
rect 4835 3241 4847 3253
rect 4774 3221 4786 3233
rect 4914 3241 4926 3253
rect 4855 3207 4867 3219
rect 4893 3207 4905 3219
rect 4974 3221 4986 3233
rect 4954 3207 4966 3219
rect 4994 3207 5006 3219
rect 5073 3252 5085 3264
rect 5087 3213 5099 3225
rect 5141 3180 5153 3192
rect 5187 3298 5199 3310
rect 5173 3278 5185 3290
rect 5205 3264 5217 3276
rect 5234 3222 5246 3234
rect 5214 3208 5226 3220
rect 5189 3176 5201 3188
rect 5211 3176 5223 3188
rect 5254 3221 5266 3233
rect 5334 3221 5346 3233
rect 5375 3241 5387 3253
rect 5355 3207 5367 3219
rect 5395 3238 5407 3250
rect 5434 3241 5446 3253
rect 5621 3298 5633 3310
rect 5603 3264 5615 3276
rect 5514 3221 5526 3233
rect 5554 3221 5566 3233
rect 5574 3222 5586 3234
rect 5594 3208 5606 3220
rect 5655 3298 5667 3310
rect 5635 3278 5647 3290
rect 5597 3176 5609 3188
rect 5619 3176 5631 3188
rect 5683 3284 5695 3296
rect 5707 3284 5719 3296
rect 5667 3180 5679 3192
rect 5735 3252 5747 3264
rect 5795 3261 5807 3273
rect 5721 3213 5733 3225
rect 5854 3241 5866 3253
rect 5834 3207 5846 3219
rect 5914 3221 5926 3233
rect 5994 3221 6006 3233
rect 5974 3207 5986 3219
rect 6034 3241 6046 3253
rect 6014 3207 6026 3219
rect 6093 3261 6105 3273
rect 6054 3207 6066 3219
rect 6154 3227 6166 3239
rect 6194 3227 6206 3239
rect 6274 3221 6286 3233
rect 6254 3207 6266 3219
rect 6334 3227 6346 3239
rect 6294 3207 6306 3219
rect 6394 3241 6406 3253
rect 6374 3227 6386 3239
rect 6541 3284 6553 3296
rect 6593 3298 6605 3310
rect 6565 3284 6577 3296
rect 6453 3261 6465 3273
rect 6414 3207 6426 3219
rect 6513 3252 6525 3264
rect 6527 3213 6539 3225
rect 6581 3180 6593 3192
rect 6627 3298 6639 3310
rect 6613 3278 6625 3290
rect 6645 3264 6657 3276
rect 6674 3222 6686 3234
rect 6654 3208 6666 3220
rect 6629 3176 6641 3188
rect 6651 3176 6663 3188
rect 6694 3221 6706 3233
rect 245 3058 257 3070
rect 34 3041 46 3053
rect 70 3044 82 3056
rect 110 3044 122 3056
rect 150 3044 162 3056
rect 314 3027 326 3039
rect 357 3072 369 3084
rect 379 3072 391 3084
rect 354 3040 366 3052
rect 274 3007 286 3019
rect 245 2990 257 3002
rect 334 3026 346 3038
rect 363 2984 375 2996
rect 395 2970 407 2982
rect 381 2950 393 2962
rect 427 3068 439 3080
rect 481 3035 493 3047
rect 554 3021 566 3033
rect 495 2996 507 3008
rect 443 2964 455 2976
rect 415 2950 427 2962
rect 467 2964 479 2976
rect 594 3021 606 3033
rect 614 3021 626 3033
rect 654 3021 666 3033
rect 754 3041 766 3053
rect 715 2987 727 2999
rect 814 3021 826 3033
rect 774 3007 786 3019
rect 854 3021 866 3033
rect 894 3021 906 3033
rect 954 3041 966 3053
rect 934 3021 946 3033
rect 994 3041 1006 3053
rect 974 3027 986 3039
rect 1087 3035 1099 3047
rect 1073 2996 1085 3008
rect 1141 3068 1153 3080
rect 1101 2964 1113 2976
rect 1125 2964 1137 2976
rect 1189 3072 1201 3084
rect 1211 3072 1223 3084
rect 1173 2970 1185 2982
rect 1153 2950 1165 2962
rect 1214 3040 1226 3052
rect 1234 3026 1246 3038
rect 1254 3027 1266 3039
rect 1205 2984 1217 2996
rect 1187 2950 1199 2962
rect 1314 3021 1326 3033
rect 1354 3021 1366 3033
rect 1407 3035 1419 3047
rect 1393 2996 1405 3008
rect 1461 3068 1473 3080
rect 1421 2964 1433 2976
rect 1445 2964 1457 2976
rect 1509 3072 1521 3084
rect 1531 3072 1543 3084
rect 1493 2970 1505 2982
rect 1473 2950 1485 2962
rect 1534 3040 1546 3052
rect 1554 3026 1566 3038
rect 1574 3027 1586 3039
rect 1654 3027 1666 3039
rect 1525 2984 1537 2996
rect 1507 2950 1519 2962
rect 1734 3041 1746 3053
rect 1695 2987 1707 2999
rect 1893 3058 1905 3070
rect 1754 3007 1766 3019
rect 1794 3007 1806 3019
rect 1834 3007 1846 3019
rect 1894 3021 1906 3033
rect 1974 3041 1986 3053
rect 1934 3007 1946 3019
rect 1954 3007 1966 3019
rect 2094 3041 2106 3053
rect 2013 2987 2025 2999
rect 2134 3041 2146 3053
rect 2114 3027 2126 3039
rect 2154 3021 2166 3033
rect 2194 3021 2206 3033
rect 2274 3027 2286 3039
rect 2335 3058 2347 3070
rect 2334 3021 2346 3033
rect 2294 3007 2306 3019
rect 2414 3027 2426 3039
rect 2457 3072 2469 3084
rect 2479 3072 2491 3084
rect 2454 3040 2466 3052
rect 2434 3026 2446 3038
rect 2463 2984 2475 2996
rect 2495 2970 2507 2982
rect 2481 2950 2493 2962
rect 2527 3068 2539 3080
rect 2581 3035 2593 3047
rect 2634 3027 2646 3039
rect 2595 2996 2607 3008
rect 2543 2964 2555 2976
rect 2515 2950 2527 2962
rect 2567 2964 2579 2976
rect 2814 3027 2826 3039
rect 2694 3007 2706 3019
rect 2734 3007 2746 3019
rect 2894 3041 2906 3053
rect 2855 2987 2867 2999
rect 2934 3041 2946 3053
rect 2914 3007 2926 3019
rect 3033 2987 3045 2999
rect 3114 3021 3126 3033
rect 3074 2987 3086 2999
rect 3054 2967 3066 2979
rect 3154 3021 3166 3033
rect 3234 3041 3246 3053
rect 3195 2987 3207 2999
rect 3274 3021 3286 3033
rect 3254 3007 3266 3019
rect 3314 3021 3326 3033
rect 3354 3021 3366 3033
rect 3394 3021 3406 3033
rect 3454 3041 3466 3053
rect 3434 3007 3446 3019
rect 3575 3058 3587 3070
rect 3574 3021 3586 3033
rect 3534 3007 3546 3019
rect 3493 2987 3505 2999
rect 3675 3041 3687 3053
rect 3713 3041 3725 3053
rect 3654 3007 3666 3019
rect 3814 3041 3826 3053
rect 3733 3007 3745 3019
rect 3854 3027 3866 3039
rect 3897 3072 3909 3084
rect 3919 3072 3931 3084
rect 3894 3040 3906 3052
rect 3874 3026 3886 3038
rect 3903 2984 3915 2996
rect 3935 2970 3947 2982
rect 3921 2950 3933 2962
rect 3967 3068 3979 3080
rect 4021 3035 4033 3047
rect 4094 3041 4106 3053
rect 4035 2996 4047 3008
rect 4074 3007 4086 3019
rect 4133 2987 4145 2999
rect 4213 2987 4225 2999
rect 3983 2964 3995 2976
rect 3955 2950 3967 2962
rect 4007 2964 4019 2976
rect 4294 3027 4306 3039
rect 4337 3072 4349 3084
rect 4359 3072 4371 3084
rect 4334 3040 4346 3052
rect 4254 2987 4266 2999
rect 4234 2967 4246 2979
rect 4314 3026 4326 3038
rect 4343 2984 4355 2996
rect 4375 2970 4387 2982
rect 4361 2950 4373 2962
rect 4407 3068 4419 3080
rect 4461 3035 4473 3047
rect 4558 3041 4570 3053
rect 4594 3041 4606 3053
rect 4475 2996 4487 3008
rect 4535 3007 4547 3019
rect 4674 3027 4686 3039
rect 4614 3007 4626 3019
rect 4423 2964 4435 2976
rect 4395 2950 4407 2962
rect 4447 2964 4459 2976
rect 4714 3007 4726 3019
rect 4753 3010 4765 3022
rect 4793 3041 4805 3053
rect 4773 3007 4785 3019
rect 4835 3041 4847 3053
rect 4873 3041 4885 3053
rect 4815 3007 4827 3019
rect 4974 3027 4986 3039
rect 4894 3007 4906 3019
rect 5015 3041 5027 3053
rect 5053 3041 5065 3053
rect 4995 3007 5007 3019
rect 5114 3027 5126 3039
rect 5074 3007 5086 3019
rect 5274 3027 5286 3039
rect 5317 3072 5329 3084
rect 5339 3072 5351 3084
rect 5314 3040 5326 3052
rect 5174 3007 5186 3019
rect 5214 3007 5226 3019
rect 5294 3026 5306 3038
rect 5323 2984 5335 2996
rect 5355 2970 5367 2982
rect 5341 2950 5353 2962
rect 5387 3068 5399 3080
rect 5441 3035 5453 3047
rect 5594 3041 5606 3053
rect 5455 2996 5467 3008
rect 5514 3007 5526 3019
rect 5554 3007 5566 3019
rect 5574 3007 5586 3019
rect 5633 2987 5645 2999
rect 5713 2987 5725 2999
rect 5403 2964 5415 2976
rect 5375 2950 5387 2962
rect 5427 2964 5439 2976
rect 5818 3041 5830 3053
rect 5854 3041 5866 3053
rect 5795 3007 5807 3019
rect 5754 2987 5766 2999
rect 5734 2967 5746 2979
rect 5955 3041 5967 3053
rect 5894 3027 5906 3039
rect 5874 3007 5886 3019
rect 5975 3007 5987 3019
rect 5995 3010 6007 3022
rect 6114 3041 6126 3053
rect 6034 3007 6046 3019
rect 6154 3041 6166 3053
rect 6134 3027 6146 3039
rect 6254 3027 6266 3039
rect 6194 3007 6206 3019
rect 6234 3007 6246 3019
rect 6355 3041 6367 3053
rect 6393 3041 6405 3053
rect 6334 3007 6346 3019
rect 6474 3027 6486 3039
rect 6494 3027 6506 3039
rect 6413 3007 6425 3019
rect 6574 3041 6586 3053
rect 6554 3007 6566 3019
rect 6613 2987 6625 2999
rect 94 2761 106 2773
rect 134 2761 146 2773
rect 14 2741 26 2753
rect 241 2818 253 2830
rect 223 2784 235 2796
rect 174 2741 186 2753
rect 194 2742 206 2754
rect 214 2728 226 2740
rect 275 2818 287 2830
rect 255 2798 267 2810
rect 217 2696 229 2708
rect 239 2696 251 2708
rect 303 2804 315 2816
rect 327 2804 339 2816
rect 287 2700 299 2712
rect 355 2772 367 2784
rect 341 2733 353 2745
rect 474 2761 486 2773
rect 514 2761 526 2773
rect 394 2741 406 2753
rect 621 2818 633 2830
rect 603 2784 615 2796
rect 554 2741 566 2753
rect 574 2742 586 2754
rect 594 2728 606 2740
rect 655 2818 667 2830
rect 635 2798 647 2810
rect 597 2696 609 2708
rect 619 2696 631 2708
rect 683 2804 695 2816
rect 707 2804 719 2816
rect 667 2700 679 2712
rect 735 2772 747 2784
rect 805 2778 817 2790
rect 721 2733 733 2745
rect 834 2761 846 2773
rect 805 2710 817 2722
rect 934 2747 946 2759
rect 854 2727 866 2739
rect 974 2747 986 2759
rect 1014 2747 1026 2759
rect 1054 2747 1066 2759
rect 1155 2761 1167 2773
rect 1094 2741 1106 2753
rect 1234 2761 1246 2773
rect 1175 2727 1187 2739
rect 1213 2727 1225 2739
rect 1334 2741 1346 2753
rect 1314 2727 1326 2739
rect 1455 2781 1467 2793
rect 1414 2741 1426 2753
rect 1354 2727 1366 2739
rect 1514 2761 1526 2773
rect 1534 2761 1546 2773
rect 1574 2761 1586 2773
rect 1494 2727 1506 2739
rect 1614 2747 1626 2759
rect 1694 2761 1706 2773
rect 1795 2781 1807 2793
rect 1734 2761 1746 2773
rect 1654 2747 1666 2759
rect 1854 2761 1866 2773
rect 1834 2727 1846 2739
rect 1913 2779 1925 2791
rect 1894 2761 1906 2773
rect 1974 2761 1986 2773
rect 1874 2741 1886 2753
rect 1913 2712 1925 2724
rect 2033 2781 2045 2793
rect 1994 2727 2006 2739
rect 2134 2741 2146 2753
rect 2114 2727 2126 2739
rect 2261 2818 2273 2830
rect 2243 2784 2255 2796
rect 2194 2741 2206 2753
rect 2214 2742 2226 2754
rect 2154 2727 2166 2739
rect 2234 2728 2246 2740
rect 2295 2818 2307 2830
rect 2275 2798 2287 2810
rect 2237 2696 2249 2708
rect 2259 2696 2271 2708
rect 2323 2804 2335 2816
rect 2347 2804 2359 2816
rect 2307 2700 2319 2712
rect 2375 2772 2387 2784
rect 2361 2733 2373 2745
rect 2414 2747 2426 2759
rect 2454 2747 2466 2759
rect 2494 2741 2506 2753
rect 2701 2818 2713 2830
rect 2683 2784 2695 2796
rect 2594 2741 2606 2753
rect 2634 2741 2646 2753
rect 2654 2742 2666 2754
rect 2674 2728 2686 2740
rect 2735 2818 2747 2830
rect 2715 2798 2727 2810
rect 2677 2696 2689 2708
rect 2699 2696 2711 2708
rect 2763 2804 2775 2816
rect 2787 2804 2799 2816
rect 2747 2700 2759 2712
rect 2815 2772 2827 2784
rect 2801 2733 2813 2745
rect 2854 2761 2866 2773
rect 3101 2804 3113 2816
rect 3153 2818 3165 2830
rect 3125 2804 3137 2816
rect 2913 2781 2925 2793
rect 2874 2727 2886 2739
rect 3014 2741 3026 2753
rect 2994 2727 3006 2739
rect 3073 2772 3085 2784
rect 3034 2727 3046 2739
rect 3087 2733 3099 2745
rect 3141 2700 3153 2712
rect 3187 2818 3199 2830
rect 3173 2798 3185 2810
rect 3205 2784 3217 2796
rect 3234 2742 3246 2754
rect 3354 2761 3366 2773
rect 3214 2728 3226 2740
rect 3189 2696 3201 2708
rect 3211 2696 3223 2708
rect 3254 2741 3266 2753
rect 3294 2741 3306 2753
rect 3433 2761 3445 2773
rect 3474 2761 3486 2773
rect 3374 2727 3386 2739
rect 3410 2727 3422 2739
rect 3533 2781 3545 2793
rect 3494 2727 3506 2739
rect 3595 2761 3607 2773
rect 3674 2761 3686 2773
rect 3694 2761 3706 2773
rect 3618 2727 3630 2739
rect 3654 2727 3666 2739
rect 3753 2781 3765 2793
rect 3714 2727 3726 2739
rect 3815 2761 3827 2773
rect 3894 2761 3906 2773
rect 3838 2727 3850 2739
rect 3874 2727 3886 2739
rect 3974 2761 3986 2773
rect 4014 2761 4026 2773
rect 4054 2761 4066 2773
rect 4094 2761 4106 2773
rect 3954 2741 3966 2753
rect 4194 2741 4206 2753
rect 4174 2727 4186 2739
rect 4234 2761 4246 2773
rect 4214 2727 4226 2739
rect 4394 2801 4406 2813
rect 4293 2781 4305 2793
rect 4373 2781 4385 2793
rect 4254 2727 4266 2739
rect 4414 2781 4426 2793
rect 4521 2818 4533 2830
rect 4503 2784 4515 2796
rect 4454 2741 4466 2753
rect 4474 2742 4486 2754
rect 4494 2728 4506 2740
rect 4555 2818 4567 2830
rect 4535 2798 4547 2810
rect 4497 2696 4509 2708
rect 4519 2696 4531 2708
rect 4583 2804 4595 2816
rect 4607 2804 4619 2816
rect 4567 2700 4579 2712
rect 4635 2772 4647 2784
rect 4621 2733 4633 2745
rect 4734 2761 4746 2773
rect 4774 2761 4786 2773
rect 4814 2761 4826 2773
rect 4674 2741 4686 2753
rect 4873 2781 4885 2793
rect 4834 2727 4846 2739
rect 4934 2761 4946 2773
rect 4974 2761 4986 2773
rect 5015 2761 5027 2773
rect 5094 2761 5106 2773
rect 5038 2727 5050 2739
rect 5074 2727 5086 2739
rect 5134 2741 5146 2753
rect 5114 2727 5126 2739
rect 5243 2778 5255 2790
rect 5214 2761 5226 2773
rect 5294 2761 5306 2773
rect 5154 2727 5166 2739
rect 5243 2710 5255 2722
rect 5353 2781 5365 2793
rect 5314 2727 5326 2739
rect 5415 2761 5427 2773
rect 5494 2761 5506 2773
rect 5438 2727 5450 2739
rect 5474 2727 5486 2739
rect 5661 2818 5673 2830
rect 5643 2784 5655 2796
rect 5554 2741 5566 2753
rect 5594 2741 5606 2753
rect 5614 2742 5626 2754
rect 5634 2728 5646 2740
rect 5695 2818 5707 2830
rect 5675 2798 5687 2810
rect 5637 2696 5649 2708
rect 5659 2696 5671 2708
rect 5723 2804 5735 2816
rect 5747 2804 5759 2816
rect 5707 2700 5719 2712
rect 5775 2772 5787 2784
rect 5761 2733 5773 2745
rect 5835 2761 5847 2773
rect 5815 2727 5827 2739
rect 5855 2758 5867 2770
rect 5894 2761 5906 2773
rect 5955 2761 5967 2773
rect 5935 2727 5947 2739
rect 5975 2758 5987 2770
rect 6014 2761 6026 2773
rect 6075 2761 6087 2773
rect 6055 2727 6067 2739
rect 6095 2758 6107 2770
rect 6134 2761 6146 2773
rect 6254 2761 6266 2773
rect 6214 2747 6226 2759
rect 6213 2710 6225 2722
rect 6354 2761 6366 2773
rect 6334 2727 6346 2739
rect 6501 2804 6513 2816
rect 6553 2818 6565 2830
rect 6525 2804 6537 2816
rect 6394 2747 6406 2759
rect 6395 2710 6407 2722
rect 6473 2772 6485 2784
rect 6487 2733 6499 2745
rect 6541 2700 6553 2712
rect 6587 2818 6599 2830
rect 6573 2798 6585 2810
rect 6605 2784 6617 2796
rect 6634 2742 6646 2754
rect 6614 2728 6626 2740
rect 6589 2696 6601 2708
rect 6611 2696 6623 2708
rect 6654 2741 6666 2753
rect 47 2555 59 2567
rect 33 2516 45 2528
rect 101 2588 113 2600
rect 61 2484 73 2496
rect 85 2484 97 2496
rect 149 2592 161 2604
rect 171 2592 183 2604
rect 133 2490 145 2502
rect 113 2470 125 2482
rect 174 2560 186 2572
rect 285 2578 297 2590
rect 194 2546 206 2558
rect 214 2547 226 2559
rect 165 2504 177 2516
rect 147 2470 159 2482
rect 314 2527 326 2539
rect 367 2555 379 2567
rect 285 2510 297 2522
rect 353 2516 365 2528
rect 421 2588 433 2600
rect 381 2484 393 2496
rect 405 2484 417 2496
rect 469 2592 481 2604
rect 491 2592 503 2604
rect 453 2490 465 2502
rect 433 2470 445 2482
rect 494 2560 506 2572
rect 614 2561 626 2573
rect 514 2546 526 2558
rect 534 2547 546 2559
rect 485 2504 497 2516
rect 467 2470 479 2482
rect 654 2561 666 2573
rect 634 2547 646 2559
rect 674 2541 686 2553
rect 714 2541 726 2553
rect 774 2541 786 2553
rect 878 2564 890 2576
rect 918 2564 930 2576
rect 958 2564 970 2576
rect 814 2541 826 2553
rect 994 2561 1006 2573
rect 1067 2555 1079 2567
rect 1053 2516 1065 2528
rect 1121 2588 1133 2600
rect 1081 2484 1093 2496
rect 1105 2484 1117 2496
rect 1169 2592 1181 2604
rect 1191 2592 1203 2604
rect 1153 2490 1165 2502
rect 1133 2470 1145 2482
rect 1194 2560 1206 2572
rect 1214 2546 1226 2558
rect 1234 2547 1246 2559
rect 1185 2504 1197 2516
rect 1167 2470 1179 2482
rect 1294 2541 1306 2553
rect 1334 2541 1346 2553
rect 1434 2547 1446 2559
rect 1354 2527 1366 2539
rect 1394 2527 1406 2539
rect 1554 2561 1566 2573
rect 1515 2507 1527 2519
rect 1614 2547 1626 2559
rect 1657 2592 1669 2604
rect 1679 2592 1691 2604
rect 1654 2560 1666 2572
rect 1574 2527 1586 2539
rect 1634 2546 1646 2558
rect 1663 2504 1675 2516
rect 1695 2490 1707 2502
rect 1681 2470 1693 2482
rect 1727 2588 1739 2600
rect 1781 2555 1793 2567
rect 1834 2547 1846 2559
rect 1894 2547 1906 2559
rect 1795 2516 1807 2528
rect 1743 2484 1755 2496
rect 1715 2470 1727 2482
rect 1767 2484 1779 2496
rect 1974 2561 1986 2573
rect 2010 2561 2022 2573
rect 1954 2527 1966 2539
rect 2155 2561 2167 2573
rect 2033 2527 2045 2539
rect 2074 2527 2086 2539
rect 2114 2527 2126 2539
rect 2175 2527 2187 2539
rect 2195 2530 2207 2542
rect 2275 2561 2287 2573
rect 2234 2527 2246 2539
rect 2295 2527 2307 2539
rect 2315 2530 2327 2542
rect 2414 2547 2426 2559
rect 2457 2592 2469 2604
rect 2479 2592 2491 2604
rect 2454 2560 2466 2572
rect 2354 2527 2366 2539
rect 2434 2546 2446 2558
rect 2463 2504 2475 2516
rect 2495 2490 2507 2502
rect 2481 2470 2493 2482
rect 2527 2588 2539 2600
rect 2581 2555 2593 2567
rect 2635 2561 2647 2573
rect 2595 2516 2607 2528
rect 2543 2484 2555 2496
rect 2515 2470 2527 2482
rect 2567 2484 2579 2496
rect 2655 2527 2667 2539
rect 2675 2530 2687 2542
rect 2714 2527 2726 2539
rect 2774 2527 2786 2539
rect 2814 2527 2826 2539
rect 2854 2527 2866 2539
rect 2893 2530 2905 2542
rect 2933 2561 2945 2573
rect 2913 2527 2925 2539
rect 2998 2561 3010 2573
rect 3034 2561 3046 2573
rect 2975 2527 2987 2539
rect 3114 2547 3126 2559
rect 3154 2547 3166 2559
rect 3197 2592 3209 2604
rect 3219 2592 3231 2604
rect 3194 2560 3206 2572
rect 3054 2527 3066 2539
rect 3174 2546 3186 2558
rect 3203 2504 3215 2516
rect 3235 2490 3247 2502
rect 3221 2470 3233 2482
rect 3267 2588 3279 2600
rect 3321 2555 3333 2567
rect 3474 2541 3486 2553
rect 3335 2516 3347 2528
rect 3374 2527 3386 2539
rect 3414 2527 3426 2539
rect 3283 2484 3295 2496
rect 3255 2470 3267 2482
rect 3307 2484 3319 2496
rect 3514 2541 3526 2553
rect 3534 2547 3546 2559
rect 3594 2507 3606 2519
rect 3635 2507 3647 2519
rect 3694 2507 3706 2519
rect 3614 2487 3626 2499
rect 3735 2507 3747 2519
rect 3714 2487 3726 2499
rect 3833 2507 3845 2519
rect 3914 2561 3926 2573
rect 3894 2527 3906 2539
rect 3874 2507 3886 2519
rect 3854 2487 3866 2499
rect 3994 2561 4006 2573
rect 4034 2561 4046 2573
rect 4014 2547 4026 2559
rect 3953 2507 3965 2519
rect 4218 2561 4230 2573
rect 4254 2561 4266 2573
rect 4114 2527 4126 2539
rect 4154 2527 4166 2539
rect 4195 2527 4207 2539
rect 4314 2547 4326 2559
rect 4357 2592 4369 2604
rect 4379 2592 4391 2604
rect 4354 2560 4366 2572
rect 4274 2527 4286 2539
rect 4334 2546 4346 2558
rect 4363 2504 4375 2516
rect 4395 2490 4407 2502
rect 4381 2470 4393 2482
rect 4427 2588 4439 2600
rect 4481 2555 4493 2567
rect 4495 2516 4507 2528
rect 4574 2547 4586 2559
rect 4443 2484 4455 2496
rect 4415 2470 4427 2482
rect 4467 2484 4479 2496
rect 4638 2561 4650 2573
rect 4674 2561 4686 2573
rect 4615 2527 4627 2539
rect 4715 2561 4727 2573
rect 4694 2527 4706 2539
rect 4735 2527 4747 2539
rect 4755 2530 4767 2542
rect 4794 2527 4806 2539
rect 4867 2555 4879 2567
rect 4853 2516 4865 2528
rect 4921 2588 4933 2600
rect 4881 2484 4893 2496
rect 4905 2484 4917 2496
rect 4969 2592 4981 2604
rect 4991 2592 5003 2604
rect 4953 2490 4965 2502
rect 4933 2470 4945 2482
rect 4994 2560 5006 2572
rect 5014 2546 5026 2558
rect 5034 2547 5046 2559
rect 5074 2547 5086 2559
rect 4985 2504 4997 2516
rect 4967 2470 4979 2482
rect 5154 2561 5166 2573
rect 5190 2561 5202 2573
rect 5134 2527 5146 2539
rect 5274 2561 5286 2573
rect 5213 2527 5225 2539
rect 5254 2527 5266 2539
rect 5534 2561 5546 2573
rect 5570 2564 5582 2576
rect 5610 2564 5622 2576
rect 5650 2564 5662 2576
rect 5354 2527 5366 2539
rect 5313 2507 5325 2519
rect 5394 2527 5406 2539
rect 5454 2527 5466 2539
rect 5494 2527 5506 2539
rect 5814 2561 5826 2573
rect 5734 2527 5746 2539
rect 5774 2527 5786 2539
rect 5794 2527 5806 2539
rect 5938 2561 5950 2573
rect 5974 2561 5986 2573
rect 5915 2527 5927 2539
rect 5853 2507 5865 2519
rect 6054 2547 6066 2559
rect 5994 2527 6006 2539
rect 6107 2555 6119 2567
rect 6093 2516 6105 2528
rect 6161 2588 6173 2600
rect 6121 2484 6133 2496
rect 6145 2484 6157 2496
rect 6209 2592 6221 2604
rect 6231 2592 6243 2604
rect 6193 2490 6205 2502
rect 6173 2470 6185 2482
rect 6234 2560 6246 2572
rect 6254 2546 6266 2558
rect 6274 2547 6286 2559
rect 6225 2504 6237 2516
rect 6207 2470 6219 2482
rect 6355 2561 6367 2573
rect 6393 2561 6405 2573
rect 6334 2527 6346 2539
rect 6434 2561 6446 2573
rect 6413 2527 6425 2539
rect 6514 2547 6526 2559
rect 6595 2561 6607 2573
rect 6633 2561 6645 2573
rect 6575 2527 6587 2539
rect 6654 2527 6666 2539
rect 101 2338 113 2350
rect 83 2304 95 2316
rect 34 2261 46 2273
rect 54 2262 66 2274
rect 74 2248 86 2260
rect 135 2338 147 2350
rect 115 2318 127 2330
rect 77 2216 89 2228
rect 99 2216 111 2228
rect 163 2324 175 2336
rect 187 2324 199 2336
rect 147 2220 159 2232
rect 215 2292 227 2304
rect 285 2298 297 2310
rect 201 2253 213 2265
rect 314 2281 326 2293
rect 285 2230 297 2242
rect 474 2281 486 2293
rect 514 2281 526 2293
rect 534 2281 546 2293
rect 434 2261 446 2273
rect 374 2247 386 2259
rect 593 2301 605 2313
rect 554 2247 566 2259
rect 754 2321 766 2333
rect 734 2301 746 2313
rect 714 2281 726 2293
rect 674 2267 686 2279
rect 673 2230 685 2242
rect 775 2301 787 2313
rect 834 2267 846 2279
rect 961 2324 973 2336
rect 1013 2338 1025 2350
rect 985 2324 997 2336
rect 933 2292 945 2304
rect 874 2267 886 2279
rect 947 2253 959 2265
rect 1001 2220 1013 2232
rect 1047 2338 1059 2350
rect 1033 2318 1045 2330
rect 1065 2304 1077 2316
rect 1094 2262 1106 2274
rect 1301 2338 1313 2350
rect 1283 2304 1295 2316
rect 1074 2248 1086 2260
rect 1049 2216 1061 2228
rect 1071 2216 1083 2228
rect 1114 2261 1126 2273
rect 1154 2261 1166 2273
rect 1234 2261 1246 2273
rect 1254 2262 1266 2274
rect 1274 2248 1286 2260
rect 1335 2338 1347 2350
rect 1315 2318 1327 2330
rect 1277 2216 1289 2228
rect 1299 2216 1311 2228
rect 1363 2324 1375 2336
rect 1387 2324 1399 2336
rect 1347 2220 1359 2232
rect 1415 2292 1427 2304
rect 1401 2253 1413 2265
rect 1514 2281 1526 2293
rect 1494 2261 1506 2273
rect 1593 2281 1605 2293
rect 1634 2281 1646 2293
rect 1534 2247 1546 2259
rect 1570 2247 1582 2259
rect 1693 2301 1705 2313
rect 1654 2247 1666 2259
rect 1754 2281 1766 2293
rect 1794 2281 1806 2293
rect 1834 2281 1846 2293
rect 1874 2281 1886 2293
rect 1915 2281 1927 2293
rect 1994 2281 2006 2293
rect 1938 2247 1950 2259
rect 1974 2247 1986 2259
rect 2161 2338 2173 2350
rect 2143 2304 2155 2316
rect 2054 2261 2066 2273
rect 2094 2261 2106 2273
rect 2114 2262 2126 2274
rect 2134 2248 2146 2260
rect 2195 2338 2207 2350
rect 2175 2318 2187 2330
rect 2137 2216 2149 2228
rect 2159 2216 2171 2228
rect 2223 2324 2235 2336
rect 2247 2324 2259 2336
rect 2207 2220 2219 2232
rect 2275 2292 2287 2304
rect 2261 2253 2273 2265
rect 2334 2281 2346 2293
rect 2374 2281 2386 2293
rect 2394 2281 2406 2293
rect 2554 2321 2566 2333
rect 2453 2301 2465 2313
rect 2533 2301 2545 2313
rect 2414 2247 2426 2259
rect 2574 2301 2586 2313
rect 2654 2261 2666 2273
rect 2634 2247 2646 2259
rect 2694 2281 2706 2293
rect 2674 2247 2686 2259
rect 2921 2324 2933 2336
rect 2973 2338 2985 2350
rect 2945 2324 2957 2336
rect 2753 2301 2765 2313
rect 2714 2247 2726 2259
rect 2814 2281 2826 2293
rect 2854 2281 2866 2293
rect 2893 2292 2905 2304
rect 2907 2253 2919 2265
rect 2961 2220 2973 2232
rect 3007 2338 3019 2350
rect 2993 2318 3005 2330
rect 3025 2304 3037 2316
rect 3054 2262 3066 2274
rect 3114 2281 3126 2293
rect 3034 2248 3046 2260
rect 3009 2216 3021 2228
rect 3031 2216 3043 2228
rect 3074 2261 3086 2273
rect 3173 2301 3185 2313
rect 3134 2247 3146 2259
rect 3235 2281 3247 2293
rect 3314 2281 3326 2293
rect 3354 2281 3366 2293
rect 3394 2281 3406 2293
rect 3258 2247 3270 2259
rect 3294 2247 3306 2259
rect 3494 2281 3506 2293
rect 3534 2281 3546 2293
rect 3454 2261 3466 2273
rect 3641 2338 3653 2350
rect 3623 2304 3635 2316
rect 3574 2261 3586 2273
rect 3594 2262 3606 2274
rect 3614 2248 3626 2260
rect 3675 2338 3687 2350
rect 3655 2318 3667 2330
rect 3617 2216 3629 2228
rect 3639 2216 3651 2228
rect 3703 2324 3715 2336
rect 3727 2324 3739 2336
rect 3687 2220 3699 2232
rect 3755 2292 3767 2304
rect 3741 2253 3753 2265
rect 3794 2267 3806 2279
rect 3894 2321 3906 2333
rect 3874 2301 3886 2313
rect 3834 2267 3846 2279
rect 3915 2301 3927 2313
rect 3995 2281 4007 2293
rect 3975 2247 3987 2259
rect 4015 2278 4027 2290
rect 4054 2281 4066 2293
rect 4115 2281 4127 2293
rect 4095 2247 4107 2259
rect 4135 2278 4147 2290
rect 4174 2281 4186 2293
rect 4235 2281 4247 2293
rect 4363 2298 4375 2310
rect 4215 2247 4227 2259
rect 4255 2278 4267 2290
rect 4294 2281 4306 2293
rect 4334 2281 4346 2293
rect 4434 2281 4446 2293
rect 4474 2281 4486 2293
rect 4363 2230 4375 2242
rect 4515 2281 4527 2293
rect 4495 2247 4507 2259
rect 4535 2278 4547 2290
rect 4574 2281 4586 2293
rect 4634 2281 4646 2293
rect 4673 2278 4685 2290
rect 4693 2281 4705 2293
rect 4755 2281 4767 2293
rect 4713 2247 4725 2259
rect 4735 2247 4747 2259
rect 4775 2278 4787 2290
rect 4814 2281 4826 2293
rect 4854 2281 4866 2293
rect 4894 2281 4906 2293
rect 4955 2281 4967 2293
rect 4935 2247 4947 2259
rect 4975 2278 4987 2290
rect 5014 2281 5026 2293
rect 5114 2261 5126 2273
rect 5094 2247 5106 2259
rect 5214 2281 5226 2293
rect 5154 2261 5166 2273
rect 5134 2247 5146 2259
rect 5293 2281 5305 2293
rect 5354 2281 5366 2293
rect 5234 2247 5246 2259
rect 5270 2247 5282 2259
rect 5393 2278 5405 2290
rect 5413 2281 5425 2293
rect 5475 2281 5487 2293
rect 5433 2247 5445 2259
rect 5455 2247 5467 2259
rect 5495 2278 5507 2290
rect 5534 2281 5546 2293
rect 5595 2281 5607 2293
rect 5754 2321 5766 2333
rect 5733 2301 5745 2313
rect 5575 2247 5587 2259
rect 5615 2278 5627 2290
rect 5654 2281 5666 2293
rect 5854 2321 5866 2333
rect 5774 2301 5786 2313
rect 5833 2301 5845 2313
rect 5874 2301 5886 2313
rect 5974 2281 5986 2293
rect 5934 2261 5946 2273
rect 6053 2281 6065 2293
rect 6094 2281 6106 2293
rect 5995 2247 6007 2259
rect 6033 2247 6045 2259
rect 6133 2278 6145 2290
rect 6153 2281 6165 2293
rect 6214 2281 6226 2293
rect 6173 2247 6185 2259
rect 6253 2278 6265 2290
rect 6273 2281 6285 2293
rect 6374 2281 6386 2293
rect 6314 2261 6326 2273
rect 6293 2247 6305 2259
rect 6433 2301 6445 2313
rect 6394 2247 6406 2259
rect 6474 2267 6486 2279
rect 6514 2267 6526 2279
rect 6574 2261 6586 2273
rect 6554 2247 6566 2259
rect 6654 2261 6666 2273
rect 6594 2247 6606 2259
rect 114 2061 126 2073
rect 34 2047 46 2059
rect 74 2047 86 2059
rect 154 2061 166 2073
rect 213 2027 225 2039
rect 254 2027 266 2039
rect 313 2027 325 2039
rect 234 2007 246 2019
rect 394 2061 406 2073
rect 354 2027 366 2039
rect 334 2007 346 2019
rect 434 2061 446 2073
rect 454 2027 466 2039
rect 654 2081 666 2093
rect 574 2047 586 2059
rect 495 2027 507 2039
rect 474 2007 486 2019
rect 614 2047 626 2059
rect 634 2047 646 2059
rect 693 2027 705 2039
rect 734 2027 746 2039
rect 934 2061 946 2073
rect 834 2047 846 2059
rect 775 2027 787 2039
rect 754 2007 766 2019
rect 874 2047 886 2059
rect 995 2081 1007 2093
rect 974 2061 986 2073
rect 1015 2047 1027 2059
rect 1035 2050 1047 2062
rect 1134 2067 1146 2079
rect 1177 2112 1189 2124
rect 1199 2112 1211 2124
rect 1174 2080 1186 2092
rect 1074 2047 1086 2059
rect 1154 2066 1166 2078
rect 1183 2024 1195 2036
rect 1215 2010 1227 2022
rect 1201 1990 1213 2002
rect 1247 2108 1259 2120
rect 1301 2075 1313 2087
rect 1354 2067 1366 2079
rect 1315 2036 1327 2048
rect 1263 2004 1275 2016
rect 1235 1990 1247 2002
rect 1287 2004 1299 2016
rect 1434 2081 1446 2093
rect 1470 2081 1482 2093
rect 1414 2047 1426 2059
rect 1493 2047 1505 2059
rect 1594 2081 1606 2093
rect 1555 2027 1567 2039
rect 1614 2047 1626 2059
rect 1694 2081 1706 2093
rect 1655 2027 1667 2039
rect 1714 2047 1726 2059
rect 1754 2047 1766 2059
rect 1794 2047 1806 2059
rect 1874 2081 1886 2093
rect 1835 2027 1847 2039
rect 1894 2047 1906 2059
rect 1934 2047 1946 2059
rect 1973 2050 1985 2062
rect 2013 2081 2025 2093
rect 1993 2047 2005 2059
rect 2054 2047 2066 2059
rect 2093 2050 2105 2062
rect 2133 2081 2145 2093
rect 2113 2047 2125 2059
rect 2174 2067 2186 2079
rect 2217 2112 2229 2124
rect 2239 2112 2251 2124
rect 2214 2080 2226 2092
rect 2194 2066 2206 2078
rect 2223 2024 2235 2036
rect 2255 2010 2267 2022
rect 2241 1990 2253 2002
rect 2287 2108 2299 2120
rect 2341 2075 2353 2087
rect 2355 2036 2367 2048
rect 2454 2081 2466 2093
rect 2415 2027 2427 2039
rect 2303 2004 2315 2016
rect 2275 1990 2287 2002
rect 2327 2004 2339 2016
rect 2474 2047 2486 2059
rect 2494 2047 2506 2059
rect 2534 2047 2546 2059
rect 2613 2027 2625 2039
rect 2675 2081 2687 2093
rect 2654 2027 2666 2039
rect 2634 2007 2646 2019
rect 2695 2047 2707 2059
rect 2715 2050 2727 2062
rect 2754 2047 2766 2059
rect 2814 2047 2826 2059
rect 2853 2050 2865 2062
rect 2893 2081 2905 2093
rect 2873 2047 2885 2059
rect 2914 2067 2926 2079
rect 2994 2081 3006 2093
rect 3030 2081 3042 2093
rect 2974 2047 2986 2059
rect 3134 2081 3146 2093
rect 3053 2047 3065 2059
rect 3174 2081 3186 2093
rect 3154 2067 3166 2079
rect 3194 2067 3206 2079
rect 3274 2081 3286 2093
rect 3310 2081 3322 2093
rect 3254 2047 3266 2059
rect 3474 2067 3486 2079
rect 3517 2112 3529 2124
rect 3539 2112 3551 2124
rect 3514 2080 3526 2092
rect 3333 2047 3345 2059
rect 3374 2047 3386 2059
rect 3414 2047 3426 2059
rect 3494 2066 3506 2078
rect 3523 2024 3535 2036
rect 3555 2010 3567 2022
rect 3541 1990 3553 2002
rect 3587 2108 3599 2120
rect 3641 2075 3653 2087
rect 3818 2081 3830 2093
rect 3854 2081 3866 2093
rect 3655 2036 3667 2048
rect 3714 2047 3726 2059
rect 3754 2047 3766 2059
rect 3795 2047 3807 2059
rect 3934 2067 3946 2079
rect 3874 2047 3886 2059
rect 3603 2004 3615 2016
rect 3575 1990 3587 2002
rect 3627 2004 3639 2016
rect 3974 2081 3986 2093
rect 3954 2047 3966 2059
rect 4054 2061 4066 2073
rect 4013 2027 4025 2039
rect 4094 2061 4106 2073
rect 4234 2067 4246 2079
rect 4277 2112 4289 2124
rect 4299 2112 4311 2124
rect 4274 2080 4286 2092
rect 4154 2047 4166 2059
rect 4194 2047 4206 2059
rect 4254 2066 4266 2078
rect 4283 2024 4295 2036
rect 4315 2010 4327 2022
rect 4301 1990 4313 2002
rect 4347 2108 4359 2120
rect 4401 2075 4413 2087
rect 4454 2067 4466 2079
rect 4415 2036 4427 2048
rect 4363 2004 4375 2016
rect 4335 1990 4347 2002
rect 4387 2004 4399 2016
rect 4534 2081 4546 2093
rect 4570 2081 4582 2093
rect 4514 2047 4526 2059
rect 4593 2047 4605 2059
rect 4634 2047 4646 2059
rect 4674 2047 4686 2059
rect 4774 2081 4786 2093
rect 4735 2027 4747 2039
rect 4914 2081 4926 2093
rect 4950 2081 4962 2093
rect 4794 2047 4806 2059
rect 4834 2047 4846 2059
rect 4874 2047 4886 2059
rect 4894 2047 4906 2059
rect 5034 2061 5046 2073
rect 4973 2047 4985 2059
rect 5074 2061 5086 2073
rect 5174 2067 5186 2079
rect 5114 2047 5126 2059
rect 5154 2047 5166 2059
rect 5213 2096 5225 2108
rect 5318 2081 5330 2093
rect 5354 2081 5366 2093
rect 5194 2047 5206 2059
rect 5295 2047 5307 2059
rect 5213 2029 5225 2041
rect 5414 2081 5426 2093
rect 5450 2081 5462 2093
rect 5374 2047 5386 2059
rect 5394 2047 5406 2059
rect 5638 2081 5650 2093
rect 5674 2081 5686 2093
rect 5473 2047 5485 2059
rect 5534 2047 5546 2059
rect 5574 2047 5586 2059
rect 5615 2047 5627 2059
rect 5754 2067 5766 2079
rect 5694 2047 5706 2059
rect 5774 2061 5786 2073
rect 5814 2061 5826 2073
rect 5887 2075 5899 2087
rect 5873 2036 5885 2048
rect 5941 2108 5953 2120
rect 5901 2004 5913 2016
rect 5925 2004 5937 2016
rect 5989 2112 6001 2124
rect 6011 2112 6023 2124
rect 5973 2010 5985 2022
rect 5953 1990 5965 2002
rect 6014 2080 6026 2092
rect 6034 2066 6046 2078
rect 6054 2067 6066 2079
rect 6114 2067 6126 2079
rect 6157 2112 6169 2124
rect 6179 2112 6191 2124
rect 6154 2080 6166 2092
rect 6005 2024 6017 2036
rect 5987 1990 5999 2002
rect 6134 2066 6146 2078
rect 6163 2024 6175 2036
rect 6195 2010 6207 2022
rect 6181 1990 6193 2002
rect 6227 2108 6239 2120
rect 6281 2075 6293 2087
rect 6335 2081 6347 2093
rect 6295 2036 6307 2048
rect 6243 2004 6255 2016
rect 6215 1990 6227 2002
rect 6267 2004 6279 2016
rect 6355 2047 6367 2059
rect 6375 2050 6387 2062
rect 6454 2081 6466 2093
rect 6414 2047 6426 2059
rect 6494 2081 6506 2093
rect 6474 2067 6486 2079
rect 6574 2081 6586 2093
rect 6554 2047 6566 2059
rect 6613 2027 6625 2039
rect 121 1844 133 1856
rect 173 1858 185 1870
rect 145 1844 157 1856
rect 93 1812 105 1824
rect 54 1781 66 1793
rect 107 1773 119 1785
rect 161 1740 173 1752
rect 207 1858 219 1870
rect 193 1838 205 1850
rect 225 1824 237 1836
rect 254 1782 266 1794
rect 314 1801 326 1813
rect 354 1801 366 1813
rect 414 1801 426 1813
rect 454 1801 466 1813
rect 234 1768 246 1780
rect 209 1736 221 1748
rect 231 1736 243 1748
rect 274 1781 286 1793
rect 681 1844 693 1856
rect 733 1858 745 1870
rect 705 1844 717 1856
rect 555 1821 567 1833
rect 514 1781 526 1793
rect 614 1801 626 1813
rect 653 1812 665 1824
rect 594 1767 606 1779
rect 667 1773 679 1785
rect 721 1740 733 1752
rect 767 1858 779 1870
rect 753 1838 765 1850
rect 785 1824 797 1836
rect 814 1782 826 1794
rect 934 1841 946 1853
rect 913 1821 925 1833
rect 794 1768 806 1780
rect 769 1736 781 1748
rect 791 1736 803 1748
rect 834 1781 846 1793
rect 954 1821 966 1833
rect 974 1801 986 1813
rect 1014 1787 1026 1799
rect 1134 1801 1146 1813
rect 1074 1781 1086 1793
rect 1015 1750 1027 1762
rect 1193 1821 1205 1833
rect 1154 1767 1166 1779
rect 1254 1787 1266 1799
rect 1374 1841 1386 1853
rect 1353 1821 1365 1833
rect 1294 1787 1306 1799
rect 1394 1821 1406 1833
rect 1561 1858 1573 1870
rect 1543 1824 1555 1836
rect 1414 1781 1426 1793
rect 1494 1781 1506 1793
rect 1514 1782 1526 1794
rect 1534 1768 1546 1780
rect 1595 1858 1607 1870
rect 1575 1838 1587 1850
rect 1537 1736 1549 1748
rect 1559 1736 1571 1748
rect 1623 1844 1635 1856
rect 1647 1844 1659 1856
rect 1607 1740 1619 1752
rect 1675 1812 1687 1824
rect 1661 1773 1673 1785
rect 1774 1801 1786 1813
rect 1714 1781 1726 1793
rect 1853 1801 1865 1813
rect 1894 1801 1906 1813
rect 1934 1801 1946 1813
rect 1974 1801 1986 1813
rect 1794 1767 1806 1779
rect 1830 1767 1842 1779
rect 2121 1844 2133 1856
rect 2173 1858 2185 1870
rect 2145 1844 2157 1856
rect 2033 1821 2045 1833
rect 1994 1767 2006 1779
rect 2093 1812 2105 1824
rect 2107 1773 2119 1785
rect 2161 1740 2173 1752
rect 2207 1858 2219 1870
rect 2193 1838 2205 1850
rect 2225 1824 2237 1836
rect 2254 1782 2266 1794
rect 2335 1801 2347 1813
rect 2234 1768 2246 1780
rect 2209 1736 2221 1748
rect 2231 1736 2243 1748
rect 2274 1781 2286 1793
rect 2414 1801 2426 1813
rect 2358 1767 2370 1779
rect 2394 1767 2406 1779
rect 2621 1844 2633 1856
rect 2673 1858 2685 1870
rect 2645 1844 2657 1856
rect 2494 1801 2506 1813
rect 2534 1801 2546 1813
rect 2593 1812 2605 1824
rect 2434 1781 2446 1793
rect 2607 1773 2619 1785
rect 2661 1740 2673 1752
rect 2707 1858 2719 1870
rect 2693 1838 2705 1850
rect 2725 1824 2737 1836
rect 2754 1782 2766 1794
rect 2834 1841 2846 1853
rect 2814 1821 2826 1833
rect 2734 1768 2746 1780
rect 2709 1736 2721 1748
rect 2731 1736 2743 1748
rect 2774 1781 2786 1793
rect 2855 1821 2867 1833
rect 2935 1821 2947 1833
rect 2994 1801 3006 1813
rect 3014 1801 3026 1813
rect 3054 1801 3066 1813
rect 2974 1767 2986 1779
rect 3154 1781 3166 1793
rect 3134 1767 3146 1779
rect 3325 1818 3337 1830
rect 3254 1781 3266 1793
rect 3174 1767 3186 1779
rect 3234 1767 3246 1779
rect 3354 1801 3366 1813
rect 3274 1767 3286 1779
rect 3325 1750 3337 1762
rect 3394 1787 3406 1799
rect 3454 1801 3466 1813
rect 3494 1801 3506 1813
rect 3434 1787 3446 1799
rect 3534 1787 3546 1799
rect 3614 1801 3626 1813
rect 3574 1787 3586 1799
rect 3673 1821 3685 1833
rect 3634 1767 3646 1779
rect 3734 1787 3746 1799
rect 3774 1787 3786 1799
rect 3834 1781 3846 1793
rect 3854 1787 3866 1799
rect 3934 1801 3946 1813
rect 3974 1801 3986 1813
rect 4014 1801 4026 1813
rect 3894 1787 3906 1799
rect 4093 1801 4105 1813
rect 4154 1801 4166 1813
rect 4194 1801 4206 1813
rect 4214 1801 4226 1813
rect 4034 1767 4046 1779
rect 4070 1767 4082 1779
rect 4273 1821 4285 1833
rect 4234 1767 4246 1779
rect 4394 1801 4406 1813
rect 4314 1767 4326 1779
rect 4453 1821 4465 1833
rect 4414 1767 4426 1779
rect 4514 1801 4526 1813
rect 4554 1801 4566 1813
rect 4595 1801 4607 1813
rect 4674 1801 4686 1813
rect 4618 1767 4630 1779
rect 4654 1767 4666 1779
rect 4801 1844 4813 1856
rect 4853 1858 4865 1870
rect 4825 1844 4837 1856
rect 4773 1812 4785 1824
rect 4734 1781 4746 1793
rect 4787 1773 4799 1785
rect 4841 1740 4853 1752
rect 4887 1858 4899 1870
rect 4873 1838 4885 1850
rect 4905 1824 4917 1836
rect 4934 1782 4946 1794
rect 4914 1768 4926 1780
rect 4889 1736 4901 1748
rect 4911 1736 4923 1748
rect 4954 1781 4966 1793
rect 5014 1781 5026 1793
rect 4994 1767 5006 1779
rect 5094 1801 5106 1813
rect 5134 1801 5146 1813
rect 5174 1801 5186 1813
rect 5034 1767 5046 1779
rect 5294 1841 5306 1853
rect 5233 1821 5245 1833
rect 5274 1821 5286 1833
rect 5194 1767 5206 1779
rect 5315 1821 5327 1833
rect 5403 1818 5415 1830
rect 5374 1801 5386 1813
rect 5494 1781 5506 1793
rect 5403 1750 5415 1762
rect 5595 1821 5607 1833
rect 5554 1767 5566 1779
rect 5654 1801 5666 1813
rect 5634 1767 5646 1779
rect 5674 1787 5686 1799
rect 5774 1801 5786 1813
rect 5714 1787 5726 1799
rect 5903 1818 5915 1830
rect 5975 1821 5987 1833
rect 5853 1801 5865 1813
rect 5874 1801 5886 1813
rect 5795 1767 5807 1779
rect 5833 1767 5845 1779
rect 5903 1750 5915 1762
rect 6034 1801 6046 1813
rect 6075 1801 6087 1813
rect 6014 1767 6026 1779
rect 6154 1801 6166 1813
rect 6098 1767 6110 1779
rect 6134 1767 6146 1779
rect 6195 1801 6207 1813
rect 6175 1767 6187 1779
rect 6215 1798 6227 1810
rect 6254 1801 6266 1813
rect 6315 1801 6327 1813
rect 6295 1767 6307 1779
rect 6335 1798 6347 1810
rect 6374 1801 6386 1813
rect 6474 1801 6486 1813
rect 6414 1781 6426 1793
rect 6533 1821 6545 1833
rect 6494 1767 6506 1779
rect 6594 1787 6606 1799
rect 6634 1787 6646 1799
rect 138 1604 150 1616
rect 178 1604 190 1616
rect 218 1604 230 1616
rect 34 1567 46 1579
rect 74 1567 86 1579
rect 254 1601 266 1613
rect 314 1587 326 1599
rect 357 1632 369 1644
rect 379 1632 391 1644
rect 354 1600 366 1612
rect 334 1586 346 1598
rect 363 1544 375 1556
rect 395 1530 407 1542
rect 381 1510 393 1522
rect 427 1628 439 1640
rect 481 1595 493 1607
rect 495 1556 507 1568
rect 574 1587 586 1599
rect 443 1524 455 1536
rect 415 1510 427 1522
rect 467 1524 479 1536
rect 594 1547 606 1559
rect 694 1601 706 1613
rect 734 1601 746 1613
rect 714 1587 726 1599
rect 635 1547 647 1559
rect 614 1527 626 1539
rect 814 1587 826 1599
rect 857 1632 869 1644
rect 879 1632 891 1644
rect 854 1600 866 1612
rect 834 1586 846 1598
rect 863 1544 875 1556
rect 895 1530 907 1542
rect 881 1510 893 1522
rect 927 1628 939 1640
rect 981 1595 993 1607
rect 995 1556 1007 1568
rect 1074 1587 1086 1599
rect 943 1524 955 1536
rect 915 1510 927 1522
rect 967 1524 979 1536
rect 1114 1601 1126 1613
rect 1150 1601 1162 1613
rect 1094 1567 1106 1579
rect 1173 1567 1185 1579
rect 1274 1601 1286 1613
rect 1235 1547 1247 1559
rect 1294 1567 1306 1579
rect 1334 1567 1346 1579
rect 1374 1567 1386 1579
rect 1414 1567 1426 1579
rect 1453 1570 1465 1582
rect 1493 1601 1505 1613
rect 1473 1567 1485 1579
rect 1534 1567 1546 1579
rect 1573 1570 1585 1582
rect 1613 1601 1625 1613
rect 1593 1567 1605 1579
rect 1654 1567 1666 1579
rect 1693 1570 1705 1582
rect 1733 1601 1745 1613
rect 1713 1567 1725 1579
rect 1787 1595 1799 1607
rect 1773 1556 1785 1568
rect 1841 1628 1853 1640
rect 1801 1524 1813 1536
rect 1825 1524 1837 1536
rect 1889 1632 1901 1644
rect 1911 1632 1923 1644
rect 1873 1530 1885 1542
rect 1853 1510 1865 1522
rect 1914 1600 1926 1612
rect 1995 1601 2007 1613
rect 1934 1586 1946 1598
rect 1954 1587 1966 1599
rect 1905 1544 1917 1556
rect 1887 1510 1899 1522
rect 2015 1567 2027 1579
rect 2035 1570 2047 1582
rect 2114 1587 2126 1599
rect 2074 1567 2086 1579
rect 2194 1601 2206 1613
rect 2230 1601 2242 1613
rect 2174 1567 2186 1579
rect 2253 1567 2265 1579
rect 2294 1567 2306 1579
rect 2334 1567 2346 1579
rect 2434 1601 2446 1613
rect 2395 1547 2407 1559
rect 2505 1618 2517 1630
rect 2654 1581 2666 1593
rect 2454 1567 2466 1579
rect 2534 1567 2546 1579
rect 2554 1567 2566 1579
rect 2505 1550 2517 1562
rect 2594 1567 2606 1579
rect 2694 1581 2706 1593
rect 2714 1581 2726 1593
rect 2754 1581 2766 1593
rect 2814 1567 2826 1579
rect 2853 1570 2865 1582
rect 2893 1601 2905 1613
rect 2873 1567 2885 1579
rect 2953 1547 2965 1559
rect 3054 1601 3066 1613
rect 2994 1547 3006 1559
rect 2974 1527 2986 1539
rect 3094 1587 3106 1599
rect 3137 1632 3149 1644
rect 3159 1632 3171 1644
rect 3134 1600 3146 1612
rect 3114 1586 3126 1598
rect 3143 1544 3155 1556
rect 3175 1530 3187 1542
rect 3161 1510 3173 1522
rect 3207 1628 3219 1640
rect 3261 1595 3273 1607
rect 3334 1581 3346 1593
rect 3275 1556 3287 1568
rect 3223 1524 3235 1536
rect 3195 1510 3207 1522
rect 3247 1524 3259 1536
rect 3374 1581 3386 1593
rect 3454 1601 3466 1613
rect 3415 1547 3427 1559
rect 3515 1601 3527 1613
rect 3553 1601 3565 1613
rect 3474 1567 3486 1579
rect 3495 1567 3507 1579
rect 3574 1567 3586 1579
rect 3674 1601 3686 1613
rect 3635 1547 3647 1559
rect 3754 1587 3766 1599
rect 3694 1567 3706 1579
rect 3898 1601 3910 1613
rect 3934 1601 3946 1613
rect 3794 1567 3806 1579
rect 3834 1567 3846 1579
rect 3875 1567 3887 1579
rect 4014 1587 4026 1599
rect 4054 1587 4066 1599
rect 4097 1632 4109 1644
rect 4119 1632 4131 1644
rect 4094 1600 4106 1612
rect 3954 1567 3966 1579
rect 4074 1586 4086 1598
rect 4103 1544 4115 1556
rect 4135 1530 4147 1542
rect 4121 1510 4133 1522
rect 4167 1628 4179 1640
rect 4221 1595 4233 1607
rect 4235 1556 4247 1568
rect 4294 1567 4306 1579
rect 4333 1570 4345 1582
rect 4373 1601 4385 1613
rect 4353 1567 4365 1579
rect 4183 1524 4195 1536
rect 4155 1510 4167 1522
rect 4207 1524 4219 1536
rect 4414 1567 4426 1579
rect 4453 1570 4465 1582
rect 4493 1601 4505 1613
rect 4515 1601 4527 1613
rect 4473 1567 4485 1579
rect 4535 1567 4547 1579
rect 4555 1570 4567 1582
rect 4635 1601 4647 1613
rect 4594 1567 4606 1579
rect 4655 1567 4667 1579
rect 4675 1570 4687 1582
rect 4755 1601 4767 1613
rect 4714 1567 4726 1579
rect 4775 1567 4787 1579
rect 4795 1570 4807 1582
rect 4875 1601 4887 1613
rect 4834 1567 4846 1579
rect 4895 1567 4907 1579
rect 4915 1570 4927 1582
rect 4954 1567 4966 1579
rect 5027 1595 5039 1607
rect 5013 1556 5025 1568
rect 5081 1628 5093 1640
rect 5041 1524 5053 1536
rect 5065 1524 5077 1536
rect 5129 1632 5141 1644
rect 5151 1632 5163 1644
rect 5113 1530 5125 1542
rect 5093 1510 5105 1522
rect 5154 1600 5166 1612
rect 5174 1586 5186 1598
rect 5194 1587 5206 1599
rect 5145 1544 5157 1556
rect 5127 1510 5139 1522
rect 5267 1595 5279 1607
rect 5253 1556 5265 1568
rect 5321 1628 5333 1640
rect 5281 1524 5293 1536
rect 5305 1524 5317 1536
rect 5369 1632 5381 1644
rect 5391 1632 5403 1644
rect 5353 1530 5365 1542
rect 5333 1510 5345 1522
rect 5394 1600 5406 1612
rect 5414 1586 5426 1598
rect 5434 1587 5446 1599
rect 5385 1544 5397 1556
rect 5367 1510 5379 1522
rect 5495 1601 5507 1613
rect 5533 1601 5545 1613
rect 5475 1567 5487 1579
rect 5595 1601 5607 1613
rect 5554 1567 5566 1579
rect 5615 1567 5627 1579
rect 5635 1570 5647 1582
rect 5674 1567 5686 1579
rect 5774 1601 5786 1613
rect 5735 1547 5747 1559
rect 5914 1581 5926 1593
rect 5794 1567 5806 1579
rect 5834 1567 5846 1579
rect 5874 1567 5886 1579
rect 5954 1581 5966 1593
rect 6034 1601 6046 1613
rect 5995 1547 6007 1559
rect 6198 1601 6210 1613
rect 6234 1601 6246 1613
rect 6054 1567 6066 1579
rect 6094 1567 6106 1579
rect 6134 1567 6146 1579
rect 6175 1567 6187 1579
rect 6254 1567 6266 1579
rect 6294 1567 6306 1579
rect 6333 1570 6345 1582
rect 6373 1601 6385 1613
rect 6353 1567 6365 1579
rect 6394 1587 6406 1599
rect 6487 1595 6499 1607
rect 6473 1556 6485 1568
rect 6541 1628 6553 1640
rect 6501 1524 6513 1536
rect 6525 1524 6537 1536
rect 6589 1632 6601 1644
rect 6611 1632 6623 1644
rect 6573 1530 6585 1542
rect 6553 1510 6565 1522
rect 6614 1600 6626 1612
rect 6634 1586 6646 1598
rect 6654 1587 6666 1599
rect 6605 1544 6617 1556
rect 6587 1510 6599 1522
rect 14 1321 26 1333
rect 54 1307 66 1319
rect 114 1321 126 1333
rect 215 1341 227 1353
rect 154 1321 166 1333
rect 55 1270 67 1282
rect 274 1321 286 1333
rect 314 1321 326 1333
rect 354 1321 366 1333
rect 254 1287 266 1299
rect 374 1301 386 1313
rect 434 1301 446 1313
rect 514 1307 526 1319
rect 554 1307 566 1319
rect 594 1301 606 1313
rect 574 1287 586 1299
rect 761 1378 773 1390
rect 743 1344 755 1356
rect 694 1301 706 1313
rect 714 1302 726 1314
rect 614 1287 626 1299
rect 734 1288 746 1300
rect 795 1378 807 1390
rect 775 1358 787 1370
rect 737 1256 749 1268
rect 759 1256 771 1268
rect 823 1364 835 1376
rect 847 1364 859 1376
rect 807 1260 819 1272
rect 875 1332 887 1344
rect 861 1293 873 1305
rect 934 1307 946 1319
rect 1014 1361 1026 1373
rect 994 1341 1006 1353
rect 974 1307 986 1319
rect 1035 1341 1047 1353
rect 1094 1321 1106 1333
rect 1134 1321 1146 1333
rect 1261 1378 1273 1390
rect 1243 1344 1255 1356
rect 1194 1301 1206 1313
rect 1214 1302 1226 1314
rect 1234 1288 1246 1300
rect 1295 1378 1307 1390
rect 1275 1358 1287 1370
rect 1237 1256 1249 1268
rect 1259 1256 1271 1268
rect 1323 1364 1335 1376
rect 1347 1364 1359 1376
rect 1307 1260 1319 1272
rect 1375 1332 1387 1344
rect 1361 1293 1373 1305
rect 1634 1321 1646 1333
rect 1458 1284 1470 1296
rect 1498 1284 1510 1296
rect 1538 1284 1550 1296
rect 1574 1287 1586 1299
rect 1673 1318 1685 1330
rect 1693 1321 1705 1333
rect 1754 1321 1766 1333
rect 1794 1321 1806 1333
rect 1835 1321 1847 1333
rect 1713 1287 1725 1299
rect 1955 1341 1967 1353
rect 1914 1321 1926 1333
rect 1858 1287 1870 1299
rect 1894 1287 1906 1299
rect 2014 1321 2026 1333
rect 1994 1287 2006 1299
rect 2094 1321 2106 1333
rect 2034 1301 2046 1313
rect 2153 1341 2165 1353
rect 2114 1287 2126 1299
rect 2194 1307 2206 1319
rect 2234 1307 2246 1319
rect 2295 1321 2307 1333
rect 2275 1287 2287 1299
rect 2315 1318 2327 1330
rect 2354 1321 2366 1333
rect 2414 1321 2426 1333
rect 2453 1318 2465 1330
rect 2473 1321 2485 1333
rect 2534 1321 2546 1333
rect 2493 1287 2505 1299
rect 2613 1321 2625 1333
rect 2635 1321 2647 1333
rect 2555 1287 2567 1299
rect 2593 1287 2605 1299
rect 2714 1321 2726 1333
rect 2774 1321 2786 1333
rect 2655 1287 2667 1299
rect 2693 1287 2705 1299
rect 2903 1338 2915 1350
rect 2853 1321 2865 1333
rect 2874 1321 2886 1333
rect 2974 1321 2986 1333
rect 2795 1287 2807 1299
rect 2833 1287 2845 1299
rect 2903 1270 2915 1282
rect 3053 1321 3065 1333
rect 2995 1287 3007 1299
rect 3033 1287 3045 1299
rect 3154 1321 3166 1333
rect 3114 1301 3126 1313
rect 3193 1318 3205 1330
rect 3213 1321 3225 1333
rect 3341 1378 3353 1390
rect 3323 1344 3335 1356
rect 3274 1301 3286 1313
rect 3294 1302 3306 1314
rect 3233 1287 3245 1299
rect 3314 1288 3326 1300
rect 3375 1378 3387 1390
rect 3355 1358 3367 1370
rect 3317 1256 3329 1268
rect 3339 1256 3351 1268
rect 3403 1364 3415 1376
rect 3427 1364 3439 1376
rect 3387 1260 3399 1272
rect 3455 1332 3467 1344
rect 3441 1293 3453 1305
rect 3514 1321 3526 1333
rect 3554 1321 3566 1333
rect 3595 1321 3607 1333
rect 3715 1341 3727 1353
rect 3674 1321 3686 1333
rect 3618 1287 3630 1299
rect 3654 1287 3666 1299
rect 3774 1321 3786 1333
rect 3754 1287 3766 1299
rect 3901 1364 3913 1376
rect 3953 1378 3965 1390
rect 3925 1364 3937 1376
rect 3873 1332 3885 1344
rect 3834 1301 3846 1313
rect 3887 1293 3899 1305
rect 3941 1260 3953 1272
rect 3987 1378 3999 1390
rect 3973 1358 3985 1370
rect 4005 1344 4017 1356
rect 4141 1364 4153 1376
rect 4193 1378 4205 1390
rect 4165 1364 4177 1376
rect 4034 1302 4046 1314
rect 4113 1332 4125 1344
rect 4014 1288 4026 1300
rect 3989 1256 4001 1268
rect 4011 1256 4023 1268
rect 4054 1301 4066 1313
rect 4127 1293 4139 1305
rect 4181 1260 4193 1272
rect 4227 1378 4239 1390
rect 4213 1358 4225 1370
rect 4245 1344 4257 1356
rect 4274 1302 4286 1314
rect 4395 1321 4407 1333
rect 4254 1288 4266 1300
rect 4229 1256 4241 1268
rect 4251 1256 4263 1268
rect 4294 1301 4306 1313
rect 4374 1301 4386 1313
rect 4474 1321 4486 1333
rect 4415 1287 4427 1299
rect 4453 1287 4465 1299
rect 4535 1321 4547 1333
rect 4515 1287 4527 1299
rect 4555 1318 4567 1330
rect 4594 1321 4606 1333
rect 4654 1321 4666 1333
rect 4785 1338 4797 1350
rect 4733 1321 4745 1333
rect 4814 1321 4826 1333
rect 4675 1287 4687 1299
rect 4713 1287 4725 1299
rect 4785 1270 4797 1282
rect 4854 1307 4866 1319
rect 4894 1307 4906 1319
rect 4934 1307 4946 1319
rect 5015 1321 5027 1333
rect 4974 1307 4986 1319
rect 5094 1321 5106 1333
rect 5135 1321 5147 1333
rect 5038 1287 5050 1299
rect 5074 1287 5086 1299
rect 5214 1321 5226 1333
rect 5158 1287 5170 1299
rect 5194 1287 5206 1299
rect 5314 1307 5326 1319
rect 5234 1287 5246 1299
rect 5374 1321 5386 1333
rect 5354 1307 5366 1319
rect 5453 1321 5465 1333
rect 5394 1287 5406 1299
rect 5430 1287 5442 1299
rect 5554 1301 5566 1313
rect 5534 1287 5546 1299
rect 5675 1321 5687 1333
rect 5574 1287 5586 1299
rect 5594 1287 5606 1299
rect 5655 1287 5667 1299
rect 5695 1318 5707 1330
rect 5734 1321 5746 1333
rect 5794 1307 5806 1319
rect 5875 1341 5887 1353
rect 5834 1307 5846 1319
rect 5934 1321 5946 1333
rect 5914 1287 5926 1299
rect 6014 1321 6026 1333
rect 5994 1301 6006 1313
rect 6281 1364 6293 1376
rect 6333 1378 6345 1390
rect 6305 1364 6317 1376
rect 6073 1341 6085 1353
rect 6034 1287 6046 1299
rect 6114 1321 6126 1333
rect 6193 1321 6205 1333
rect 6253 1332 6265 1344
rect 6134 1287 6146 1299
rect 6170 1287 6182 1299
rect 6267 1293 6279 1305
rect 6321 1260 6333 1272
rect 6367 1378 6379 1390
rect 6353 1358 6365 1370
rect 6385 1344 6397 1356
rect 6521 1364 6533 1376
rect 6573 1378 6585 1390
rect 6545 1364 6557 1376
rect 6414 1302 6426 1314
rect 6493 1332 6505 1344
rect 6394 1288 6406 1300
rect 6369 1256 6381 1268
rect 6391 1256 6403 1268
rect 6434 1301 6446 1313
rect 6507 1293 6519 1305
rect 6561 1260 6573 1272
rect 6607 1378 6619 1390
rect 6593 1358 6605 1370
rect 6625 1344 6637 1356
rect 6654 1302 6666 1314
rect 6634 1288 6646 1300
rect 6609 1256 6621 1268
rect 6631 1256 6643 1268
rect 6674 1301 6686 1313
rect 47 1115 59 1127
rect 33 1076 45 1088
rect 101 1148 113 1160
rect 61 1044 73 1056
rect 85 1044 97 1056
rect 149 1152 161 1164
rect 171 1152 183 1164
rect 133 1050 145 1062
rect 113 1030 125 1042
rect 174 1120 186 1132
rect 194 1106 206 1118
rect 214 1107 226 1119
rect 294 1107 306 1119
rect 165 1064 177 1076
rect 147 1030 159 1042
rect 347 1115 359 1127
rect 333 1076 345 1088
rect 401 1148 413 1160
rect 361 1044 373 1056
rect 385 1044 397 1056
rect 449 1152 461 1164
rect 471 1152 483 1164
rect 433 1050 445 1062
rect 413 1030 425 1042
rect 474 1120 486 1132
rect 494 1106 506 1118
rect 514 1107 526 1119
rect 554 1107 566 1119
rect 465 1064 477 1076
rect 447 1030 459 1042
rect 614 1067 626 1079
rect 714 1087 726 1099
rect 655 1067 667 1079
rect 634 1047 646 1059
rect 754 1087 766 1099
rect 794 1067 806 1079
rect 894 1101 906 1113
rect 835 1067 847 1079
rect 814 1047 826 1059
rect 934 1101 946 1113
rect 974 1107 986 1119
rect 1054 1107 1066 1119
rect 1097 1152 1109 1164
rect 1119 1152 1131 1164
rect 1094 1120 1106 1132
rect 1074 1106 1086 1118
rect 1103 1064 1115 1076
rect 1135 1050 1147 1062
rect 1121 1030 1133 1042
rect 1167 1148 1179 1160
rect 1221 1115 1233 1127
rect 1235 1076 1247 1088
rect 1294 1121 1306 1133
rect 1330 1124 1342 1136
rect 1370 1124 1382 1136
rect 1410 1124 1422 1136
rect 1494 1107 1506 1119
rect 1537 1152 1549 1164
rect 1559 1152 1571 1164
rect 1534 1120 1546 1132
rect 1514 1106 1526 1118
rect 1183 1044 1195 1056
rect 1155 1030 1167 1042
rect 1207 1044 1219 1056
rect 1543 1064 1555 1076
rect 1575 1050 1587 1062
rect 1561 1030 1573 1042
rect 1607 1148 1619 1160
rect 1661 1115 1673 1127
rect 1838 1121 1850 1133
rect 1874 1121 1886 1133
rect 1675 1076 1687 1088
rect 1734 1087 1746 1099
rect 1774 1087 1786 1099
rect 1815 1087 1827 1099
rect 1894 1087 1906 1099
rect 1974 1121 1986 1133
rect 1935 1067 1947 1079
rect 1623 1044 1635 1056
rect 1595 1030 1607 1042
rect 1647 1044 1659 1056
rect 1994 1087 2006 1099
rect 2074 1121 2086 1133
rect 2035 1067 2047 1079
rect 2238 1121 2250 1133
rect 2274 1121 2286 1133
rect 2094 1087 2106 1099
rect 2134 1087 2146 1099
rect 2174 1087 2186 1099
rect 2215 1087 2227 1099
rect 2334 1107 2346 1119
rect 2377 1152 2389 1164
rect 2399 1152 2411 1164
rect 2374 1120 2386 1132
rect 2294 1087 2306 1099
rect 2354 1106 2366 1118
rect 2383 1064 2395 1076
rect 2415 1050 2427 1062
rect 2401 1030 2413 1042
rect 2447 1148 2459 1160
rect 2501 1115 2513 1127
rect 2515 1076 2527 1088
rect 2594 1107 2606 1119
rect 2463 1044 2475 1056
rect 2435 1030 2447 1042
rect 2487 1044 2499 1056
rect 2634 1121 2646 1133
rect 2614 1087 2626 1099
rect 2745 1138 2757 1150
rect 2794 1107 2806 1119
rect 2774 1087 2786 1099
rect 2673 1067 2685 1079
rect 2745 1070 2757 1082
rect 2895 1121 2907 1133
rect 2933 1121 2945 1133
rect 2874 1087 2886 1099
rect 2994 1107 3006 1119
rect 3037 1152 3049 1164
rect 3059 1152 3071 1164
rect 3034 1120 3046 1132
rect 2953 1087 2965 1099
rect 3014 1106 3026 1118
rect 3043 1064 3055 1076
rect 3075 1050 3087 1062
rect 3061 1030 3073 1042
rect 3107 1148 3119 1160
rect 3161 1115 3173 1127
rect 3214 1101 3226 1113
rect 3175 1076 3187 1088
rect 3123 1044 3135 1056
rect 3095 1030 3107 1042
rect 3147 1044 3159 1056
rect 3254 1101 3266 1113
rect 3314 1087 3326 1099
rect 3353 1090 3365 1102
rect 3393 1121 3405 1133
rect 3415 1121 3427 1133
rect 3373 1087 3385 1099
rect 3435 1087 3447 1099
rect 3455 1090 3467 1102
rect 3565 1138 3577 1150
rect 3634 1107 3646 1119
rect 3677 1152 3689 1164
rect 3699 1152 3711 1164
rect 3674 1120 3686 1132
rect 3494 1087 3506 1099
rect 3594 1087 3606 1099
rect 3565 1070 3577 1082
rect 3654 1106 3666 1118
rect 3683 1064 3695 1076
rect 3715 1050 3727 1062
rect 3701 1030 3713 1042
rect 3747 1148 3759 1160
rect 3801 1115 3813 1127
rect 3855 1121 3867 1133
rect 3815 1076 3827 1088
rect 3763 1044 3775 1056
rect 3735 1030 3747 1042
rect 3787 1044 3799 1056
rect 3875 1087 3887 1099
rect 3895 1090 3907 1102
rect 3934 1087 3946 1099
rect 3994 1087 4006 1099
rect 4033 1090 4045 1102
rect 4073 1121 4085 1133
rect 4053 1087 4065 1099
rect 4094 1107 4106 1119
rect 4174 1121 4186 1133
rect 4210 1121 4222 1133
rect 4154 1087 4166 1099
rect 4233 1087 4245 1099
rect 4274 1087 4286 1099
rect 4314 1087 4326 1099
rect 4414 1121 4426 1133
rect 4375 1067 4387 1079
rect 4494 1121 4506 1133
rect 4434 1087 4446 1099
rect 4534 1121 4546 1133
rect 4514 1107 4526 1119
rect 4574 1107 4586 1119
rect 4617 1152 4629 1164
rect 4639 1152 4651 1164
rect 4614 1120 4626 1132
rect 4594 1106 4606 1118
rect 4623 1064 4635 1076
rect 4655 1050 4667 1062
rect 4641 1030 4653 1042
rect 4687 1148 4699 1160
rect 4741 1115 4753 1127
rect 4814 1121 4826 1133
rect 4850 1121 4862 1133
rect 4755 1076 4767 1088
rect 4794 1087 4806 1099
rect 4873 1087 4885 1099
rect 4934 1087 4946 1099
rect 4974 1087 4986 1099
rect 5054 1121 5066 1133
rect 5015 1067 5027 1079
rect 4703 1044 4715 1056
rect 4675 1030 4687 1042
rect 4727 1044 4739 1056
rect 5365 1138 5377 1150
rect 5574 1121 5586 1133
rect 5074 1087 5086 1099
rect 5114 1087 5126 1099
rect 5154 1087 5166 1099
rect 5174 1087 5186 1099
rect 5214 1087 5226 1099
rect 5254 1087 5266 1099
rect 5294 1087 5306 1099
rect 5394 1087 5406 1099
rect 5414 1087 5426 1099
rect 5365 1070 5377 1082
rect 5454 1087 5466 1099
rect 5494 1087 5506 1099
rect 5534 1087 5546 1099
rect 5614 1121 5626 1133
rect 5594 1107 5606 1119
rect 5674 1107 5686 1119
rect 5713 1136 5725 1148
rect 5874 1121 5886 1133
rect 5694 1087 5706 1099
rect 5794 1087 5806 1099
rect 5713 1069 5725 1081
rect 5834 1087 5846 1099
rect 5854 1087 5866 1099
rect 5913 1067 5925 1079
rect 5993 1067 6005 1079
rect 6074 1121 6086 1133
rect 6054 1087 6066 1099
rect 6034 1067 6046 1079
rect 6014 1047 6026 1059
rect 6174 1087 6186 1099
rect 6113 1067 6125 1079
rect 6214 1087 6226 1099
rect 6234 1087 6246 1099
rect 6274 1087 6286 1099
rect 6347 1115 6359 1127
rect 6333 1076 6345 1088
rect 6401 1148 6413 1160
rect 6361 1044 6373 1056
rect 6385 1044 6397 1056
rect 6449 1152 6461 1164
rect 6471 1152 6483 1164
rect 6433 1050 6445 1062
rect 6413 1030 6425 1042
rect 6474 1120 6486 1132
rect 6494 1106 6506 1118
rect 6514 1107 6526 1119
rect 6465 1064 6477 1076
rect 6447 1030 6459 1042
rect 6574 1121 6586 1133
rect 6610 1121 6622 1133
rect 6554 1087 6566 1099
rect 6633 1087 6645 1099
rect 53 859 65 871
rect 34 841 46 853
rect 14 821 26 833
rect 134 827 146 839
rect 241 884 253 896
rect 293 898 305 910
rect 265 884 277 896
rect 213 852 225 864
rect 174 827 186 839
rect 53 792 65 804
rect 227 813 239 825
rect 281 780 293 792
rect 327 898 339 910
rect 313 878 325 890
rect 345 864 357 876
rect 374 822 386 834
rect 514 841 526 853
rect 554 841 566 853
rect 574 841 586 853
rect 614 841 626 853
rect 354 808 366 820
rect 329 776 341 788
rect 351 776 363 788
rect 394 821 406 833
rect 474 821 486 833
rect 654 827 666 839
rect 754 881 766 893
rect 734 861 746 873
rect 694 827 706 839
rect 775 861 787 873
rect 834 841 846 853
rect 913 841 925 853
rect 954 841 966 853
rect 854 807 866 819
rect 890 807 902 819
rect 1013 861 1025 873
rect 974 807 986 819
rect 1054 841 1066 853
rect 1113 861 1125 873
rect 1074 807 1086 819
rect 1234 841 1246 853
rect 1254 807 1266 819
rect 1294 841 1306 853
rect 1334 841 1346 853
rect 1393 861 1405 873
rect 1354 807 1366 819
rect 1581 898 1593 910
rect 1563 864 1575 876
rect 1474 821 1486 833
rect 1514 821 1526 833
rect 1534 822 1546 834
rect 1554 808 1566 820
rect 1615 898 1627 910
rect 1595 878 1607 890
rect 1557 776 1569 788
rect 1579 776 1591 788
rect 1643 884 1655 896
rect 1667 884 1679 896
rect 1627 780 1639 792
rect 1695 852 1707 864
rect 1681 813 1693 825
rect 1734 821 1746 833
rect 1815 841 1827 853
rect 1795 807 1807 819
rect 1835 838 1847 850
rect 1874 841 1886 853
rect 1914 841 1926 853
rect 1973 861 1985 873
rect 1934 807 1946 819
rect 2014 827 2026 839
rect 2141 884 2153 896
rect 2193 898 2205 910
rect 2165 884 2177 896
rect 2113 852 2125 864
rect 2054 827 2066 839
rect 2127 813 2139 825
rect 2181 780 2193 792
rect 2227 898 2239 910
rect 2213 878 2225 890
rect 2245 864 2257 876
rect 2274 822 2286 834
rect 2394 841 2406 853
rect 2254 808 2266 820
rect 2229 776 2241 788
rect 2251 776 2263 788
rect 2294 821 2306 833
rect 2334 821 2346 833
rect 2473 841 2485 853
rect 2514 841 2526 853
rect 2615 861 2627 873
rect 2554 841 2566 853
rect 2414 807 2426 819
rect 2450 807 2462 819
rect 2674 841 2686 853
rect 2654 807 2666 819
rect 2914 821 2926 833
rect 2738 804 2750 816
rect 2778 804 2790 816
rect 2818 804 2830 816
rect 2854 807 2866 819
rect 2894 807 2906 819
rect 2934 807 2946 819
rect 3054 821 3066 833
rect 3034 807 3046 819
rect 3114 841 3126 853
rect 3074 807 3086 819
rect 3153 838 3165 850
rect 3173 841 3185 853
rect 3234 841 3246 853
rect 3193 807 3205 819
rect 3273 838 3285 850
rect 3293 841 3305 853
rect 3355 861 3367 873
rect 3313 807 3325 819
rect 3414 841 3426 853
rect 3394 807 3406 819
rect 3434 827 3446 839
rect 3474 827 3486 839
rect 3535 841 3547 853
rect 3515 807 3527 819
rect 3555 838 3567 850
rect 3594 841 3606 853
rect 3714 841 3726 853
rect 3674 821 3686 833
rect 3753 838 3765 850
rect 3773 841 3785 853
rect 3901 898 3913 910
rect 3883 864 3895 876
rect 3834 821 3846 833
rect 3854 822 3866 834
rect 3793 807 3805 819
rect 3874 808 3886 820
rect 3935 898 3947 910
rect 3915 878 3927 890
rect 3877 776 3889 788
rect 3899 776 3911 788
rect 3963 884 3975 896
rect 3987 884 3999 896
rect 3947 780 3959 792
rect 4015 852 4027 864
rect 4001 813 4013 825
rect 4075 841 4087 853
rect 4055 807 4067 819
rect 4095 838 4107 850
rect 4134 841 4146 853
rect 4194 821 4206 833
rect 4174 807 4186 819
rect 4274 841 4286 853
rect 4214 807 4226 819
rect 4434 881 4446 893
rect 4333 861 4345 873
rect 4413 861 4425 873
rect 4294 807 4306 819
rect 4454 861 4466 873
rect 4534 841 4546 853
rect 4474 821 4486 833
rect 4593 861 4605 873
rect 4554 807 4566 819
rect 4634 827 4646 839
rect 4674 827 4686 839
rect 4774 841 4786 853
rect 4754 821 4766 833
rect 4833 861 4845 873
rect 4794 807 4806 819
rect 4874 827 4886 839
rect 4914 827 4926 839
rect 4975 841 4987 853
rect 4955 807 4967 819
rect 4995 838 5007 850
rect 5034 841 5046 853
rect 5094 841 5106 853
rect 5133 838 5145 850
rect 5153 841 5165 853
rect 5173 807 5185 819
rect 5214 807 5226 819
rect 5414 821 5426 833
rect 5250 804 5262 816
rect 5290 804 5302 816
rect 5330 804 5342 816
rect 5394 807 5406 819
rect 5434 807 5446 819
rect 5554 841 5566 853
rect 5534 821 5546 833
rect 5613 861 5625 873
rect 5574 807 5586 819
rect 5654 827 5666 839
rect 5734 841 5746 853
rect 5694 827 5706 839
rect 5894 881 5906 893
rect 5793 861 5805 873
rect 5873 861 5885 873
rect 5754 807 5766 819
rect 5914 861 5926 873
rect 6021 898 6033 910
rect 6003 864 6015 876
rect 5954 821 5966 833
rect 5974 822 5986 834
rect 5994 808 6006 820
rect 6055 898 6067 910
rect 6035 878 6047 890
rect 5997 776 6009 788
rect 6019 776 6031 788
rect 6083 884 6095 896
rect 6107 884 6119 896
rect 6067 780 6079 792
rect 6135 852 6147 864
rect 6121 813 6133 825
rect 6174 841 6186 853
rect 6233 861 6245 873
rect 6194 807 6206 819
rect 6274 841 6286 853
rect 6333 861 6345 873
rect 6294 807 6306 819
rect 6394 827 6406 839
rect 6434 827 6446 839
rect 6541 898 6553 910
rect 6523 864 6535 876
rect 6474 821 6486 833
rect 6494 822 6506 834
rect 6514 808 6526 820
rect 6575 898 6587 910
rect 6555 878 6567 890
rect 6517 776 6529 788
rect 6539 776 6551 788
rect 6603 884 6615 896
rect 6627 884 6639 896
rect 6587 780 6599 792
rect 6655 852 6667 864
rect 6641 813 6653 825
rect 14 627 26 639
rect 74 621 86 633
rect 154 641 166 653
rect 114 621 126 633
rect 194 641 206 653
rect 174 627 186 639
rect 254 627 266 639
rect 354 641 366 653
rect 394 641 406 653
rect 374 627 386 639
rect 414 587 426 599
rect 534 621 546 633
rect 455 587 467 599
rect 434 567 446 579
rect 574 621 586 633
rect 633 587 645 599
rect 694 627 706 639
rect 754 627 766 639
rect 674 587 686 599
rect 654 567 666 579
rect 994 641 1006 653
rect 834 607 846 619
rect 874 607 886 619
rect 974 607 986 619
rect 1094 627 1106 639
rect 1137 672 1149 684
rect 1159 672 1171 684
rect 1134 640 1146 652
rect 1034 607 1046 619
rect 1114 626 1126 638
rect 1143 584 1155 596
rect 1175 570 1187 582
rect 1161 550 1173 562
rect 1207 668 1219 680
rect 1261 635 1273 647
rect 1343 658 1355 670
rect 1394 621 1406 633
rect 1275 596 1287 608
rect 1314 607 1326 619
rect 1223 564 1235 576
rect 1195 550 1207 562
rect 1247 564 1259 576
rect 1343 590 1355 602
rect 1434 621 1446 633
rect 1494 627 1506 639
rect 1537 672 1549 684
rect 1559 672 1571 684
rect 1534 640 1546 652
rect 1514 626 1526 638
rect 1543 584 1555 596
rect 1575 570 1587 582
rect 1561 550 1573 562
rect 1607 668 1619 680
rect 1661 635 1673 647
rect 1734 627 1746 639
rect 1777 672 1789 684
rect 1799 672 1811 684
rect 1774 640 1786 652
rect 1675 596 1687 608
rect 1754 626 1766 638
rect 1623 564 1635 576
rect 1595 550 1607 562
rect 1647 564 1659 576
rect 1783 584 1795 596
rect 1815 570 1827 582
rect 1801 550 1813 562
rect 1847 668 1859 680
rect 1901 635 1913 647
rect 1974 627 1986 639
rect 2017 672 2029 684
rect 2039 672 2051 684
rect 2014 640 2026 652
rect 1915 596 1927 608
rect 1994 626 2006 638
rect 1863 564 1875 576
rect 1835 550 1847 562
rect 1887 564 1899 576
rect 2023 584 2035 596
rect 2055 570 2067 582
rect 2041 550 2053 562
rect 2087 668 2099 680
rect 2141 635 2153 647
rect 2214 627 2226 639
rect 2257 672 2269 684
rect 2279 672 2291 684
rect 2254 640 2266 652
rect 2155 596 2167 608
rect 2234 626 2246 638
rect 2103 564 2115 576
rect 2075 550 2087 562
rect 2127 564 2139 576
rect 2263 584 2275 596
rect 2295 570 2307 582
rect 2281 550 2293 562
rect 2327 668 2339 680
rect 2381 635 2393 647
rect 2395 596 2407 608
rect 2467 635 2479 647
rect 2453 596 2465 608
rect 2343 564 2355 576
rect 2315 550 2327 562
rect 2367 564 2379 576
rect 2521 668 2533 680
rect 2481 564 2493 576
rect 2505 564 2517 576
rect 2569 672 2581 684
rect 2591 672 2603 684
rect 2553 570 2565 582
rect 2533 550 2545 562
rect 2594 640 2606 652
rect 2614 626 2626 638
rect 2634 627 2646 639
rect 2585 584 2597 596
rect 2567 550 2579 562
rect 2715 641 2727 653
rect 2753 641 2765 653
rect 2694 607 2706 619
rect 2894 641 2906 653
rect 2834 627 2846 639
rect 2773 607 2785 619
rect 2934 641 2946 653
rect 2914 627 2926 639
rect 2954 627 2966 639
rect 3034 641 3046 653
rect 3014 607 3026 619
rect 3114 621 3126 633
rect 3073 587 3085 599
rect 3154 621 3166 633
rect 3194 587 3206 599
rect 3294 627 3306 639
rect 3235 587 3247 599
rect 3214 567 3226 579
rect 3374 641 3386 653
rect 3354 607 3366 619
rect 3454 621 3466 633
rect 3413 587 3425 599
rect 3534 641 3546 653
rect 3494 621 3506 633
rect 3574 641 3586 653
rect 3554 627 3566 639
rect 3734 641 3746 653
rect 3634 607 3646 619
rect 3674 607 3686 619
rect 3714 607 3726 619
rect 3773 587 3785 599
rect 3853 587 3865 599
rect 3947 635 3959 647
rect 3894 587 3906 599
rect 3933 596 3945 608
rect 3874 567 3886 579
rect 4001 668 4013 680
rect 3961 564 3973 576
rect 3985 564 3997 576
rect 4049 672 4061 684
rect 4071 672 4083 684
rect 4033 570 4045 582
rect 4013 550 4025 562
rect 4074 640 4086 652
rect 4094 626 4106 638
rect 4114 627 4126 639
rect 4065 584 4077 596
rect 4047 550 4059 562
rect 4174 607 4186 619
rect 4214 607 4226 619
rect 4267 635 4279 647
rect 4253 596 4265 608
rect 4321 668 4333 680
rect 4281 564 4293 576
rect 4305 564 4317 576
rect 4369 672 4381 684
rect 4391 672 4403 684
rect 4353 570 4365 582
rect 4333 550 4345 562
rect 4394 640 4406 652
rect 4414 626 4426 638
rect 4434 627 4446 639
rect 4474 627 4486 639
rect 4385 584 4397 596
rect 4367 550 4379 562
rect 4555 641 4567 653
rect 4593 641 4605 653
rect 4535 607 4547 619
rect 4694 641 4706 653
rect 4614 607 4626 619
rect 4734 641 4746 653
rect 4714 627 4726 639
rect 4814 641 4826 653
rect 4775 587 4787 599
rect 4854 621 4866 633
rect 4834 607 4846 619
rect 4894 621 4906 633
rect 4974 627 4986 639
rect 5014 607 5026 619
rect 5053 610 5065 622
rect 5093 641 5105 653
rect 5073 607 5085 619
rect 5114 587 5126 599
rect 5247 635 5259 647
rect 5155 587 5167 599
rect 5134 567 5146 579
rect 5233 596 5245 608
rect 5301 668 5313 680
rect 5261 564 5273 576
rect 5285 564 5297 576
rect 5349 672 5361 684
rect 5371 672 5383 684
rect 5333 570 5345 582
rect 5313 550 5325 562
rect 5374 640 5386 652
rect 5454 641 5466 653
rect 5515 641 5527 653
rect 5394 626 5406 638
rect 5414 627 5426 639
rect 5365 584 5377 596
rect 5347 550 5359 562
rect 5535 607 5547 619
rect 5555 610 5567 622
rect 6054 641 6066 653
rect 5594 607 5606 619
rect 5654 607 5666 619
rect 5694 607 5706 619
rect 5734 607 5746 619
rect 5774 607 5786 619
rect 5814 607 5826 619
rect 5854 607 5866 619
rect 5874 607 5886 619
rect 5914 607 5926 619
rect 5974 607 5986 619
rect 6014 607 6026 619
rect 6034 607 6046 619
rect 6154 641 6166 653
rect 6134 607 6146 619
rect 6093 587 6105 599
rect 6254 621 6266 633
rect 6193 587 6205 599
rect 6294 621 6306 633
rect 6334 627 6346 639
rect 6377 672 6389 684
rect 6399 672 6411 684
rect 6374 640 6386 652
rect 6354 626 6366 638
rect 6383 584 6395 596
rect 6415 570 6427 582
rect 6401 550 6413 562
rect 6447 668 6459 680
rect 6501 635 6513 647
rect 6554 627 6566 639
rect 6614 627 6626 639
rect 6515 596 6527 608
rect 6463 564 6475 576
rect 6435 550 6447 562
rect 6487 564 6499 576
rect 61 404 73 416
rect 113 418 125 430
rect 85 404 97 416
rect 33 372 45 384
rect 47 333 59 345
rect 101 300 113 312
rect 147 418 159 430
rect 133 398 145 410
rect 165 384 177 396
rect 194 342 206 354
rect 341 418 353 430
rect 323 384 335 396
rect 174 328 186 340
rect 149 296 161 308
rect 171 296 183 308
rect 214 341 226 353
rect 274 341 286 353
rect 294 342 306 354
rect 314 328 326 340
rect 375 418 387 430
rect 355 398 367 410
rect 317 296 329 308
rect 339 296 351 308
rect 403 404 415 416
rect 427 404 439 416
rect 387 300 399 312
rect 514 401 526 413
rect 455 372 467 384
rect 494 381 506 393
rect 441 333 453 345
rect 535 381 547 393
rect 594 361 606 373
rect 634 361 646 373
rect 694 361 706 373
rect 734 361 746 373
rect 754 347 766 359
rect 794 347 806 359
rect 981 418 993 430
rect 963 384 975 396
rect 874 341 886 353
rect 914 341 926 353
rect 934 342 946 354
rect 954 328 966 340
rect 1015 418 1027 430
rect 995 398 1007 410
rect 957 296 969 308
rect 979 296 991 308
rect 1043 404 1055 416
rect 1067 404 1079 416
rect 1027 300 1039 312
rect 1095 372 1107 384
rect 1165 378 1177 390
rect 1081 333 1093 345
rect 1243 378 1255 390
rect 1323 378 1335 390
rect 1194 361 1206 373
rect 1214 361 1226 373
rect 1294 361 1306 373
rect 1165 310 1177 322
rect 1243 310 1255 322
rect 1434 361 1446 373
rect 1414 341 1426 353
rect 1323 310 1335 322
rect 1493 381 1505 393
rect 1454 327 1466 339
rect 1594 361 1606 373
rect 1574 341 1586 353
rect 1653 381 1665 393
rect 1614 327 1626 339
rect 1781 418 1793 430
rect 1763 384 1775 396
rect 1714 341 1726 353
rect 1734 342 1746 354
rect 1754 328 1766 340
rect 1815 418 1827 430
rect 1795 398 1807 410
rect 1757 296 1769 308
rect 1779 296 1791 308
rect 1843 404 1855 416
rect 1867 404 1879 416
rect 1827 300 1839 312
rect 1895 372 1907 384
rect 1881 333 1893 345
rect 2054 361 2066 373
rect 1974 341 1986 353
rect 2034 341 2046 353
rect 2113 381 2125 393
rect 2074 327 2086 339
rect 2214 361 2226 373
rect 2154 341 2166 353
rect 2355 381 2367 393
rect 2293 361 2305 373
rect 2234 327 2246 339
rect 2270 327 2282 339
rect 2414 361 2426 373
rect 2434 361 2446 373
rect 2474 361 2486 373
rect 2394 327 2406 339
rect 2601 418 2613 430
rect 2583 384 2595 396
rect 2534 341 2546 353
rect 2554 342 2566 354
rect 2574 328 2586 340
rect 2635 418 2647 430
rect 2615 398 2627 410
rect 2577 296 2589 308
rect 2599 296 2611 308
rect 2663 404 2675 416
rect 2687 404 2699 416
rect 2647 300 2659 312
rect 2715 372 2727 384
rect 2775 381 2787 393
rect 2701 333 2713 345
rect 2834 361 2846 373
rect 2854 361 2866 373
rect 2894 361 2906 373
rect 2814 327 2826 339
rect 3021 418 3033 430
rect 3003 384 3015 396
rect 2954 341 2966 353
rect 2974 342 2986 354
rect 2994 328 3006 340
rect 3055 418 3067 430
rect 3035 398 3047 410
rect 2997 296 3009 308
rect 3019 296 3031 308
rect 3083 404 3095 416
rect 3107 404 3119 416
rect 3067 300 3079 312
rect 3135 372 3147 384
rect 3121 333 3133 345
rect 3174 347 3186 359
rect 3275 381 3287 393
rect 3214 347 3226 359
rect 3334 361 3346 373
rect 3354 361 3366 373
rect 3394 361 3406 373
rect 3314 327 3326 339
rect 3494 341 3506 353
rect 3474 327 3486 339
rect 3534 361 3546 373
rect 3514 327 3526 339
rect 3593 381 3605 393
rect 3554 327 3566 339
rect 3634 361 3646 373
rect 3674 361 3686 373
rect 3734 341 3746 353
rect 3714 327 3726 339
rect 3834 361 3846 373
rect 3874 361 3886 373
rect 3894 361 3906 373
rect 3754 327 3766 339
rect 4054 401 4066 413
rect 3953 381 3965 393
rect 4033 381 4045 393
rect 3914 327 3926 339
rect 4221 404 4233 416
rect 4273 418 4285 430
rect 4245 404 4257 416
rect 4074 381 4086 393
rect 4094 361 4106 373
rect 4134 361 4146 373
rect 4193 372 4205 384
rect 4207 333 4219 345
rect 4261 300 4273 312
rect 4307 418 4319 430
rect 4293 398 4305 410
rect 4325 384 4337 396
rect 4354 342 4366 354
rect 4414 361 4426 373
rect 4515 381 4527 393
rect 4454 361 4466 373
rect 4334 328 4346 340
rect 4309 296 4321 308
rect 4331 296 4343 308
rect 4374 341 4386 353
rect 4574 361 4586 373
rect 4594 361 4606 373
rect 4634 361 4646 373
rect 4695 361 4707 373
rect 4554 327 4566 339
rect 4774 361 4786 373
rect 4718 327 4730 339
rect 4754 327 4766 339
rect 4941 418 4953 430
rect 4923 384 4935 396
rect 4834 341 4846 353
rect 4874 341 4886 353
rect 4894 342 4906 354
rect 4914 328 4926 340
rect 4975 418 4987 430
rect 4955 398 4967 410
rect 4917 296 4929 308
rect 4939 296 4951 308
rect 5003 404 5015 416
rect 5027 404 5039 416
rect 4987 300 4999 312
rect 5055 372 5067 384
rect 5041 333 5053 345
rect 5154 341 5166 353
rect 5134 327 5146 339
rect 5194 361 5206 373
rect 5295 381 5307 393
rect 5234 361 5246 373
rect 5174 327 5186 339
rect 5354 361 5366 373
rect 5374 361 5386 373
rect 5414 361 5426 373
rect 5334 327 5346 339
rect 5474 341 5486 353
rect 5454 327 5466 339
rect 5574 401 5586 413
rect 5554 381 5566 393
rect 5494 327 5506 339
rect 5595 381 5607 393
rect 5654 361 5666 373
rect 5713 381 5725 393
rect 5674 327 5686 339
rect 5774 347 5786 359
rect 5855 381 5867 393
rect 5814 347 5826 359
rect 5914 361 5926 373
rect 5934 361 5946 373
rect 5894 327 5906 339
rect 5993 381 6005 393
rect 5954 327 5966 339
rect 6034 361 6046 373
rect 6093 381 6105 393
rect 6054 327 6066 339
rect 6154 361 6166 373
rect 6194 361 6206 373
rect 6234 361 6246 373
rect 6274 361 6286 373
rect 6315 361 6327 373
rect 6394 361 6406 373
rect 6338 327 6350 339
rect 6374 327 6386 339
rect 6501 418 6513 430
rect 6483 384 6495 396
rect 6434 341 6446 353
rect 6454 342 6466 354
rect 6474 328 6486 340
rect 6535 418 6547 430
rect 6515 398 6527 410
rect 6477 296 6489 308
rect 6499 296 6511 308
rect 6563 404 6575 416
rect 6587 404 6599 416
rect 6547 300 6559 312
rect 6615 372 6627 384
rect 6601 333 6613 345
rect 47 155 59 167
rect 33 116 45 128
rect 101 188 113 200
rect 61 84 73 96
rect 85 84 97 96
rect 149 192 161 204
rect 171 192 183 204
rect 133 90 145 102
rect 113 70 125 82
rect 174 160 186 172
rect 194 146 206 158
rect 214 147 226 159
rect 165 104 177 116
rect 147 70 159 82
rect 287 155 299 167
rect 273 116 285 128
rect 341 188 353 200
rect 301 84 313 96
rect 325 84 337 96
rect 389 192 401 204
rect 411 192 423 204
rect 373 90 385 102
rect 353 70 365 82
rect 414 160 426 172
rect 525 178 537 190
rect 434 146 446 158
rect 454 147 466 159
rect 405 104 417 116
rect 387 70 399 82
rect 603 178 615 190
rect 685 178 697 190
rect 554 127 566 139
rect 574 127 586 139
rect 525 110 537 122
rect 714 127 726 139
rect 767 155 779 167
rect 603 110 615 122
rect 685 110 697 122
rect 753 116 765 128
rect 821 188 833 200
rect 781 84 793 96
rect 805 84 817 96
rect 869 192 881 204
rect 891 192 903 204
rect 853 90 865 102
rect 833 70 845 82
rect 894 160 906 172
rect 914 146 926 158
rect 934 147 946 159
rect 885 104 897 116
rect 867 70 879 82
rect 1003 178 1015 190
rect 1074 141 1086 153
rect 974 127 986 139
rect 1003 110 1015 122
rect 1114 141 1126 153
rect 1194 161 1206 173
rect 1155 107 1167 119
rect 1254 147 1266 159
rect 1297 192 1309 204
rect 1319 192 1331 204
rect 1294 160 1306 172
rect 1214 127 1226 139
rect 1274 146 1286 158
rect 1303 104 1315 116
rect 1335 90 1347 102
rect 1321 70 1333 82
rect 1367 188 1379 200
rect 1421 155 1433 167
rect 1435 116 1447 128
rect 1514 147 1526 159
rect 1383 84 1395 96
rect 1355 70 1367 82
rect 1407 84 1419 96
rect 1534 141 1546 153
rect 1574 141 1586 153
rect 1674 161 1686 173
rect 1635 107 1647 119
rect 1714 147 1726 159
rect 1694 127 1706 139
rect 1774 141 1786 153
rect 1814 141 1826 153
rect 1854 141 1866 153
rect 1894 141 1906 153
rect 1934 141 1946 153
rect 1974 141 1986 153
rect 2074 161 2086 173
rect 2035 107 2047 119
rect 2134 147 2146 159
rect 2177 192 2189 204
rect 2199 192 2211 204
rect 2174 160 2186 172
rect 2094 127 2106 139
rect 2154 146 2166 158
rect 2183 104 2195 116
rect 2215 90 2227 102
rect 2201 70 2213 82
rect 2247 188 2259 200
rect 2301 155 2313 167
rect 2354 141 2366 153
rect 2315 116 2327 128
rect 2263 84 2275 96
rect 2235 70 2247 82
rect 2287 84 2299 96
rect 2394 141 2406 153
rect 2454 141 2466 153
rect 2494 141 2506 153
rect 2574 161 2586 173
rect 2535 107 2547 119
rect 2654 147 2666 159
rect 2694 147 2706 159
rect 2737 192 2749 204
rect 2759 192 2771 204
rect 2734 160 2746 172
rect 2594 127 2606 139
rect 2714 146 2726 158
rect 2743 104 2755 116
rect 2775 90 2787 102
rect 2761 70 2773 82
rect 2807 188 2819 200
rect 2861 155 2873 167
rect 2875 116 2887 128
rect 2974 161 2986 173
rect 2935 107 2947 119
rect 2823 84 2835 96
rect 2795 70 2807 82
rect 2847 84 2859 96
rect 3138 161 3150 173
rect 3174 161 3186 173
rect 2994 127 3006 139
rect 3034 127 3046 139
rect 3074 127 3086 139
rect 3115 127 3127 139
rect 3254 147 3266 159
rect 3194 127 3206 139
rect 3307 155 3319 167
rect 3293 116 3305 128
rect 3361 188 3373 200
rect 3321 84 3333 96
rect 3345 84 3357 96
rect 3409 192 3421 204
rect 3431 192 3443 204
rect 3393 90 3405 102
rect 3373 70 3385 82
rect 3434 160 3446 172
rect 3454 146 3466 158
rect 3474 147 3486 159
rect 3425 104 3437 116
rect 3407 70 3419 82
rect 3534 141 3546 153
rect 3574 141 3586 153
rect 3654 161 3666 173
rect 3615 107 3627 119
rect 3714 161 3726 173
rect 3674 127 3686 139
rect 3694 127 3706 139
rect 3827 155 3839 167
rect 3753 107 3765 119
rect 3813 116 3825 128
rect 3881 188 3893 200
rect 3841 84 3853 96
rect 3865 84 3877 96
rect 3929 192 3941 204
rect 3951 192 3963 204
rect 3913 90 3925 102
rect 3893 70 3905 82
rect 3954 160 3966 172
rect 3974 146 3986 158
rect 3994 147 4006 159
rect 3945 104 3957 116
rect 3927 70 3939 82
rect 4054 161 4066 173
rect 4034 127 4046 139
rect 4154 161 4166 173
rect 4134 127 4146 139
rect 4093 107 4105 119
rect 4234 141 4246 153
rect 4193 107 4205 119
rect 4274 141 4286 153
rect 4347 155 4359 167
rect 4333 116 4345 128
rect 4401 188 4413 200
rect 4361 84 4373 96
rect 4385 84 4397 96
rect 4449 192 4461 204
rect 4471 192 4483 204
rect 4433 90 4445 102
rect 4413 70 4425 82
rect 4474 160 4486 172
rect 4494 146 4506 158
rect 4514 147 4526 159
rect 4465 104 4477 116
rect 4447 70 4459 82
rect 4574 161 4586 173
rect 4554 127 4566 139
rect 4674 161 4686 173
rect 4654 127 4666 139
rect 4613 107 4625 119
rect 4754 141 4766 153
rect 4713 107 4725 119
rect 4794 141 4806 153
rect 4867 155 4879 167
rect 4853 116 4865 128
rect 4921 188 4933 200
rect 4881 84 4893 96
rect 4905 84 4917 96
rect 4969 192 4981 204
rect 4991 192 5003 204
rect 4953 90 4965 102
rect 4933 70 4945 82
rect 4994 160 5006 172
rect 5014 146 5026 158
rect 5034 147 5046 159
rect 4985 104 4997 116
rect 4967 70 4979 82
rect 5134 161 5146 173
rect 5095 107 5107 119
rect 5194 161 5206 173
rect 5154 127 5166 139
rect 5174 127 5186 139
rect 5274 141 5286 153
rect 5233 107 5245 119
rect 5314 141 5326 153
rect 5387 155 5399 167
rect 5373 116 5385 128
rect 5441 188 5453 200
rect 5401 84 5413 96
rect 5425 84 5437 96
rect 5489 192 5501 204
rect 5511 192 5523 204
rect 5473 90 5485 102
rect 5453 70 5465 82
rect 5514 160 5526 172
rect 5534 146 5546 158
rect 5554 147 5566 159
rect 5505 104 5517 116
rect 5487 70 5499 82
rect 5627 155 5639 167
rect 5613 116 5625 128
rect 5681 188 5693 200
rect 5641 84 5653 96
rect 5665 84 5677 96
rect 5729 192 5741 204
rect 5751 192 5763 204
rect 5713 90 5725 102
rect 5693 70 5705 82
rect 5754 160 5766 172
rect 5774 146 5786 158
rect 5794 147 5806 159
rect 5745 104 5757 116
rect 5727 70 5739 82
rect 5867 155 5879 167
rect 5853 116 5865 128
rect 5921 188 5933 200
rect 5881 84 5893 96
rect 5905 84 5917 96
rect 5969 192 5981 204
rect 5991 192 6003 204
rect 5953 90 5965 102
rect 5933 70 5945 82
rect 5994 160 6006 172
rect 6114 161 6126 173
rect 6014 146 6026 158
rect 6034 147 6046 159
rect 5985 104 5997 116
rect 5967 70 5979 82
rect 6154 161 6166 173
rect 6134 127 6146 139
rect 6278 161 6290 173
rect 6314 161 6326 173
rect 6255 127 6267 139
rect 6193 107 6205 119
rect 6394 147 6406 159
rect 6334 127 6346 139
rect 6447 155 6459 167
rect 6433 116 6445 128
rect 6501 188 6513 200
rect 6461 84 6473 96
rect 6485 84 6497 96
rect 6549 192 6561 204
rect 6571 192 6583 204
rect 6533 90 6545 102
rect 6513 70 6525 82
rect 6574 160 6586 172
rect 6594 146 6606 158
rect 6614 147 6626 159
rect 6565 104 6577 116
rect 6547 70 6559 82
<< metal1 >>
rect -62 6258 -2 6498
rect 4 6496 6802 6498
rect 6736 6484 6802 6496
rect 4 6482 6802 6484
rect 41 6476 53 6482
rect 103 6476 115 6482
rect 151 6476 163 6482
rect 209 6476 221 6482
rect 311 6476 323 6482
rect 359 6476 371 6482
rect 489 6476 501 6482
rect 60 6456 73 6462
rect 60 6450 67 6456
rect 125 6444 132 6456
rect 21 6352 27 6436
rect 111 6437 132 6444
rect 182 6450 189 6456
rect 182 6442 193 6450
rect 79 6426 86 6432
rect 147 6426 153 6428
rect 79 6420 153 6426
rect 235 6421 243 6436
rect 79 6412 86 6420
rect 40 6404 74 6412
rect 40 6399 46 6404
rect 66 6386 93 6393
rect 21 6344 83 6352
rect 95 6348 139 6354
rect 77 6330 115 6338
rect 133 6334 139 6348
rect 147 6348 153 6420
rect 227 6407 243 6421
rect 275 6422 283 6436
rect 303 6436 331 6442
rect 291 6433 343 6436
rect 389 6428 401 6436
rect 377 6422 401 6428
rect 519 6476 531 6482
rect 619 6476 631 6482
rect 677 6476 689 6482
rect 725 6476 737 6482
rect 787 6476 799 6482
rect 837 6476 849 6482
rect 900 6476 912 6482
rect 956 6476 968 6482
rect 1051 6476 1063 6482
rect 1099 6476 1111 6482
rect 1157 6476 1169 6482
rect 1205 6476 1217 6482
rect 1267 6476 1279 6482
rect 1337 6476 1349 6482
rect 1491 6476 1503 6482
rect 1581 6476 1593 6482
rect 1671 6476 1683 6482
rect 1719 6476 1731 6482
rect 1777 6476 1789 6482
rect 1825 6476 1837 6482
rect 1887 6476 1899 6482
rect 1957 6476 1969 6482
rect 2039 6476 2051 6482
rect 2171 6476 2183 6482
rect 2238 6476 2250 6482
rect 2288 6476 2300 6482
rect 2369 6476 2381 6482
rect 459 6428 471 6436
rect 549 6428 561 6436
rect 275 6415 300 6422
rect 213 6393 227 6407
rect 147 6342 187 6348
rect 207 6348 221 6356
rect 235 6344 243 6407
rect 293 6393 301 6415
rect 299 6344 307 6379
rect 377 6373 385 6422
rect 417 6417 433 6423
rect 77 6324 85 6330
rect 133 6328 163 6334
rect 181 6324 187 6342
rect 67 6310 85 6324
rect 113 6310 135 6322
rect 77 6304 85 6310
rect 127 6304 139 6310
rect 181 6284 193 6318
rect 377 6304 385 6359
rect 417 6343 423 6417
rect 459 6422 483 6428
rect 475 6373 483 6422
rect 537 6422 561 6428
rect 767 6456 780 6462
rect 651 6450 658 6456
rect 647 6442 658 6450
rect 708 6444 715 6456
rect 773 6450 780 6456
rect 537 6373 545 6422
rect 597 6421 605 6436
rect 708 6437 729 6444
rect 687 6426 693 6428
rect 754 6426 761 6432
rect 597 6407 613 6421
rect 687 6420 761 6426
rect 397 6337 423 6343
rect 397 6327 403 6337
rect 475 6304 483 6359
rect 537 6304 545 6359
rect 597 6344 605 6407
rect 613 6393 627 6407
rect 619 6348 633 6356
rect 41 6258 53 6264
rect 107 6258 119 6264
rect 153 6258 165 6264
rect 211 6258 223 6264
rect 276 6258 288 6264
rect 326 6258 338 6264
rect 357 6258 369 6264
rect 397 6258 409 6264
rect 451 6258 463 6264
rect 491 6258 503 6264
rect 687 6348 693 6420
rect 754 6412 761 6420
rect 766 6404 800 6412
rect 794 6399 800 6404
rect 747 6386 774 6393
rect 653 6342 693 6348
rect 701 6348 745 6354
rect 653 6324 659 6342
rect 701 6334 707 6348
rect 813 6352 819 6436
rect 856 6401 864 6456
rect 757 6344 819 6352
rect 677 6328 707 6334
rect 725 6330 763 6338
rect 755 6324 763 6330
rect 647 6284 659 6318
rect 705 6310 727 6322
rect 755 6310 773 6324
rect 701 6304 713 6310
rect 755 6304 763 6310
rect 856 6304 864 6387
rect 933 6393 940 6436
rect 1036 6401 1044 6456
rect 1247 6456 1260 6462
rect 1131 6450 1138 6456
rect 1127 6442 1138 6450
rect 1188 6444 1195 6456
rect 1253 6450 1260 6456
rect 1077 6421 1085 6436
rect 1188 6437 1209 6444
rect 1167 6426 1173 6428
rect 1234 6426 1241 6432
rect 1077 6407 1093 6421
rect 1167 6420 1241 6426
rect 941 6356 947 6379
rect 941 6350 968 6356
rect 956 6344 968 6350
rect 909 6336 937 6342
rect 949 6264 977 6270
rect 1036 6304 1044 6387
rect 1077 6344 1085 6407
rect 1093 6393 1107 6407
rect 1099 6348 1113 6356
rect 1167 6348 1173 6420
rect 1234 6412 1241 6420
rect 1246 6404 1280 6412
rect 1274 6399 1280 6404
rect 1227 6386 1254 6393
rect 1133 6342 1173 6348
rect 1181 6348 1225 6354
rect 1133 6324 1139 6342
rect 1181 6334 1187 6348
rect 1293 6352 1299 6436
rect 1329 6436 1357 6440
rect 1369 6470 1397 6476
rect 1317 6434 1369 6436
rect 1379 6426 1385 6436
rect 1356 6419 1385 6426
rect 1455 6422 1463 6436
rect 1483 6436 1511 6442
rect 1471 6433 1523 6436
rect 1551 6436 1561 6446
rect 1356 6393 1364 6419
rect 1455 6415 1480 6422
rect 1427 6397 1453 6403
rect 1473 6393 1481 6415
rect 1551 6393 1559 6436
rect 1611 6426 1623 6436
rect 1585 6418 1623 6426
rect 1551 6379 1553 6393
rect 1237 6344 1299 6352
rect 1357 6344 1365 6379
rect 1479 6344 1487 6379
rect 1551 6344 1559 6379
rect 1157 6328 1187 6334
rect 1205 6330 1243 6338
rect 1235 6324 1243 6330
rect 1127 6284 1139 6318
rect 1185 6310 1207 6322
rect 1235 6310 1253 6324
rect 1181 6304 1193 6310
rect 1235 6304 1243 6310
rect 517 6258 529 6264
rect 557 6258 569 6264
rect 617 6258 629 6264
rect 675 6258 687 6264
rect 721 6258 733 6264
rect 787 6258 799 6264
rect 837 6258 849 6264
rect 917 6258 929 6264
rect 1051 6258 1063 6264
rect 1097 6258 1109 6264
rect 1155 6258 1167 6264
rect 1201 6258 1213 6264
rect 1267 6258 1279 6264
rect 1317 6258 1329 6264
rect 1387 6258 1399 6264
rect -62 6256 1433 6258
rect 1594 6304 1602 6418
rect 1656 6401 1664 6456
rect 1867 6456 1880 6462
rect 1751 6450 1758 6456
rect 1747 6442 1758 6450
rect 1808 6444 1815 6456
rect 1873 6450 1880 6456
rect 1697 6421 1705 6436
rect 1808 6437 1829 6444
rect 1787 6426 1793 6428
rect 1854 6426 1861 6432
rect 1697 6407 1713 6421
rect 1787 6420 1861 6426
rect 1656 6304 1664 6387
rect 1697 6344 1705 6407
rect 1713 6393 1727 6407
rect 1719 6348 1733 6356
rect 1787 6348 1793 6420
rect 1854 6412 1861 6420
rect 1866 6404 1900 6412
rect 1894 6399 1900 6404
rect 1847 6386 1874 6393
rect 1753 6342 1793 6348
rect 1801 6348 1845 6354
rect 1753 6324 1759 6342
rect 1801 6334 1807 6348
rect 1913 6352 1919 6436
rect 1949 6436 1977 6442
rect 1937 6433 1989 6436
rect 1997 6422 2005 6436
rect 2069 6428 2081 6436
rect 1980 6415 2005 6422
rect 2057 6422 2081 6428
rect 2135 6422 2143 6436
rect 2163 6436 2191 6442
rect 2151 6433 2203 6436
rect 2234 6436 2260 6447
rect 2411 6476 2423 6482
rect 2451 6476 2463 6482
rect 2477 6476 2489 6482
rect 2517 6476 2529 6482
rect 2559 6476 2571 6482
rect 2710 6476 2722 6482
rect 1979 6393 1987 6415
rect 1857 6344 1919 6352
rect 1973 6344 1981 6379
rect 2057 6373 2065 6422
rect 2135 6415 2160 6422
rect 2153 6393 2161 6415
rect 2234 6393 2242 6436
rect 2339 6428 2351 6436
rect 2339 6422 2363 6428
rect 1777 6328 1807 6334
rect 1825 6330 1863 6338
rect 1855 6324 1863 6330
rect 1747 6284 1759 6318
rect 1805 6310 1827 6322
rect 1855 6310 1873 6324
rect 1801 6304 1813 6310
rect 1855 6304 1863 6310
rect 2057 6304 2065 6359
rect 2159 6344 2167 6379
rect 2234 6344 2242 6379
rect 2355 6373 2363 6422
rect 2433 6413 2440 6456
rect 2500 6413 2507 6456
rect 2589 6428 2601 6436
rect 1456 6258 1468 6264
rect 1506 6258 1518 6264
rect 1567 6258 1579 6264
rect 1611 6258 1623 6264
rect 1671 6258 1683 6264
rect 1717 6258 1729 6264
rect 1775 6258 1787 6264
rect 1821 6258 1833 6264
rect 1887 6258 1899 6264
rect 1942 6258 1954 6264
rect 1992 6258 2004 6264
rect 2037 6258 2049 6264
rect 2077 6258 2089 6264
rect 1447 6256 2113 6258
rect 2263 6338 2303 6344
rect 2291 6336 2303 6338
rect 2355 6304 2363 6359
rect 2433 6351 2440 6399
rect 2423 6344 2440 6351
rect 2500 6351 2507 6399
rect 2577 6422 2601 6428
rect 2577 6373 2585 6422
rect 2656 6418 2674 6420
rect 2656 6409 2686 6418
rect 2739 6476 2751 6482
rect 2890 6476 2902 6482
rect 2971 6476 2983 6482
rect 3071 6476 3083 6482
rect 3151 6476 3163 6482
rect 3211 6476 3223 6482
rect 2769 6428 2781 6436
rect 2757 6422 2781 6428
rect 2656 6381 2664 6409
rect 2500 6344 2517 6351
rect 2136 6258 2148 6264
rect 2186 6258 2198 6264
rect 2271 6258 2283 6264
rect 2331 6258 2343 6264
rect 2371 6258 2383 6264
rect 2451 6258 2463 6264
rect 2577 6304 2585 6359
rect 2655 6312 2662 6367
rect 2757 6373 2765 6422
rect 2836 6418 2854 6420
rect 2836 6409 2866 6418
rect 2935 6422 2943 6436
rect 2963 6436 2991 6442
rect 2951 6433 3003 6436
rect 3035 6422 3043 6436
rect 3063 6436 3091 6442
rect 3240 6476 3252 6482
rect 3290 6476 3302 6482
rect 3357 6476 3369 6482
rect 3458 6476 3470 6482
rect 3508 6476 3520 6482
rect 3051 6433 3103 6436
rect 2935 6415 2960 6422
rect 3035 6415 3060 6422
rect 2836 6381 2844 6409
rect 2953 6393 2961 6415
rect 3053 6393 3061 6415
rect 3136 6401 3144 6456
rect 3196 6401 3204 6456
rect 3280 6436 3306 6447
rect 3298 6393 3306 6436
rect 3349 6436 3377 6442
rect 3337 6433 3389 6436
rect 3454 6436 3480 6447
rect 3558 6476 3570 6482
rect 3608 6476 3620 6482
rect 3554 6436 3580 6447
rect 3638 6476 3650 6482
rect 3791 6476 3803 6482
rect 3857 6476 3869 6482
rect 3937 6476 3949 6482
rect 3999 6476 4011 6482
rect 4121 6476 4133 6482
rect 4179 6476 4191 6482
rect 4330 6476 4342 6482
rect 4430 6476 4442 6482
rect 4530 6476 4542 6482
rect 3397 6422 3405 6436
rect 3380 6415 3405 6422
rect 2655 6306 2702 6312
rect 2655 6304 2663 6306
rect 2691 6304 2702 6306
rect 2757 6304 2765 6359
rect 2835 6312 2842 6367
rect 2959 6344 2967 6379
rect 3059 6344 3067 6379
rect 2835 6306 2882 6312
rect 2835 6304 2843 6306
rect 2477 6258 2489 6264
rect 2557 6258 2569 6264
rect 2597 6258 2609 6264
rect 2671 6258 2683 6264
rect 2711 6258 2723 6264
rect 2871 6304 2882 6306
rect 2737 6258 2749 6264
rect 2777 6258 2789 6264
rect 2851 6258 2863 6264
rect 2891 6258 2903 6264
rect 2936 6258 2948 6264
rect 2986 6258 2998 6264
rect 3136 6304 3144 6387
rect 3196 6304 3204 6387
rect 3379 6393 3387 6415
rect 3454 6393 3462 6436
rect 3554 6393 3562 6436
rect 3755 6422 3763 6436
rect 3783 6436 3811 6442
rect 3771 6433 3823 6436
rect 3849 6436 3877 6442
rect 3837 6433 3889 6436
rect 3897 6422 3905 6436
rect 3686 6418 3704 6420
rect 3674 6409 3704 6418
rect 3755 6415 3780 6422
rect 3880 6415 3905 6422
rect 3696 6381 3704 6409
rect 3773 6393 3781 6415
rect 3298 6344 3306 6379
rect 3373 6344 3381 6379
rect 3454 6344 3462 6379
rect 3554 6344 3562 6379
rect 3879 6393 3887 6415
rect 3956 6401 3964 6456
rect 4029 6428 4041 6436
rect 4017 6422 4041 6428
rect 4091 6436 4101 6446
rect 3237 6338 3277 6344
rect 3237 6336 3249 6338
rect 3483 6338 3523 6344
rect 3511 6336 3523 6338
rect 3583 6338 3623 6344
rect 3611 6336 3623 6338
rect 3698 6312 3705 6367
rect 3779 6344 3787 6379
rect 3873 6344 3881 6379
rect 3658 6306 3705 6312
rect 3658 6304 3669 6306
rect 3697 6304 3705 6306
rect 3036 6258 3048 6264
rect 3086 6258 3098 6264
rect 3151 6258 3163 6264
rect 3211 6258 3223 6264
rect 3257 6258 3269 6264
rect 3342 6258 3354 6264
rect 3392 6258 3404 6264
rect 3491 6258 3503 6264
rect 3591 6258 3603 6264
rect 3637 6258 3649 6264
rect 3677 6258 3689 6264
rect 3756 6258 3768 6264
rect 3806 6258 3818 6264
rect 3956 6304 3964 6387
rect 4017 6373 4025 6422
rect 4091 6393 4099 6436
rect 4151 6426 4163 6436
rect 4209 6428 4221 6436
rect 4125 6418 4163 6426
rect 4197 6422 4221 6428
rect 4091 6379 4093 6393
rect 4017 6304 4025 6359
rect 4091 6344 4099 6379
rect 3842 6258 3854 6264
rect 3892 6258 3904 6264
rect 4134 6304 4142 6418
rect 4197 6373 4205 6422
rect 4276 6418 4294 6420
rect 4276 6409 4306 6418
rect 4376 6418 4394 6420
rect 4376 6409 4406 6418
rect 4476 6418 4494 6420
rect 4476 6409 4506 6418
rect 4557 6476 4569 6482
rect 4620 6476 4632 6482
rect 4670 6476 4682 6482
rect 4276 6381 4284 6409
rect 4376 6381 4384 6409
rect 4476 6381 4484 6409
rect 4576 6401 4584 6456
rect 4720 6476 4732 6482
rect 4770 6476 4782 6482
rect 4837 6476 4849 6482
rect 4971 6476 4983 6482
rect 5037 6476 5049 6482
rect 5190 6476 5202 6482
rect 5290 6476 5302 6482
rect 5390 6476 5402 6482
rect 4660 6436 4686 6447
rect 4760 6436 4786 6447
rect 4678 6393 4686 6436
rect 4197 6304 4205 6359
rect 4275 6312 4282 6367
rect 4375 6312 4382 6367
rect 4475 6312 4482 6367
rect 4275 6306 4322 6312
rect 4275 6304 4283 6306
rect 3937 6258 3949 6264
rect 3997 6258 4009 6264
rect 4037 6258 4049 6264
rect 4107 6258 4119 6264
rect 4151 6258 4163 6264
rect 4311 6304 4322 6306
rect 4375 6306 4422 6312
rect 4375 6304 4383 6306
rect 4411 6304 4422 6306
rect 4475 6306 4522 6312
rect 4475 6304 4483 6306
rect 4511 6304 4522 6306
rect 4576 6304 4584 6387
rect 4607 6357 4633 6363
rect 4678 6344 4686 6379
rect 4697 6363 4703 6413
rect 4778 6393 4786 6436
rect 4829 6436 4857 6442
rect 4817 6433 4869 6436
rect 4877 6422 4885 6436
rect 4860 6415 4885 6422
rect 4935 6422 4943 6436
rect 4963 6436 4991 6442
rect 4951 6433 5003 6436
rect 5029 6436 5057 6442
rect 5017 6433 5069 6436
rect 5077 6422 5085 6436
rect 4935 6415 4960 6422
rect 5060 6415 5085 6422
rect 5136 6418 5154 6420
rect 4859 6393 4867 6415
rect 4887 6397 4893 6403
rect 4953 6393 4961 6415
rect 5059 6393 5067 6415
rect 5136 6409 5166 6418
rect 5136 6381 5144 6409
rect 4697 6357 4713 6363
rect 4778 6344 4786 6379
rect 4853 6344 4861 6379
rect 4959 6344 4967 6379
rect 5053 6344 5061 6379
rect 4617 6338 4657 6344
rect 4617 6336 4629 6338
rect 4177 6258 4189 6264
rect 4217 6258 4229 6264
rect 4291 6258 4303 6264
rect 4331 6258 4343 6264
rect 4391 6258 4403 6264
rect 4431 6258 4443 6264
rect 4491 6258 4503 6264
rect 4531 6258 4543 6264
rect 4717 6338 4757 6344
rect 4717 6336 4729 6338
rect 4887 6317 4913 6323
rect 4557 6258 4569 6264
rect 4637 6258 4649 6264
rect 4737 6258 4749 6264
rect 4822 6258 4834 6264
rect 4872 6258 4884 6264
rect 4936 6258 4948 6264
rect 4986 6258 4998 6264
rect 5135 6312 5142 6367
rect 5217 6323 5223 6433
rect 5236 6418 5254 6420
rect 5236 6409 5266 6418
rect 5336 6418 5354 6420
rect 5336 6409 5366 6418
rect 5420 6476 5432 6482
rect 5470 6476 5482 6482
rect 5538 6476 5550 6482
rect 5588 6476 5600 6482
rect 5651 6476 5663 6482
rect 5460 6436 5486 6447
rect 5236 6381 5244 6409
rect 5287 6397 5313 6403
rect 5336 6381 5344 6409
rect 5478 6393 5486 6436
rect 5534 6436 5560 6447
rect 5680 6476 5692 6482
rect 5730 6476 5742 6482
rect 5534 6393 5542 6436
rect 5207 6317 5223 6323
rect 5235 6312 5242 6367
rect 5636 6401 5644 6456
rect 5778 6476 5790 6482
rect 5898 6476 5910 6482
rect 5948 6476 5960 6482
rect 6011 6476 6023 6482
rect 5720 6436 5746 6447
rect 5738 6393 5746 6436
rect 5894 6436 5920 6447
rect 6058 6476 6070 6482
rect 6108 6476 6120 6482
rect 6191 6476 6203 6482
rect 6258 6476 6270 6482
rect 6308 6476 6320 6482
rect 5826 6418 5844 6420
rect 5814 6409 5844 6418
rect 5335 6312 5342 6367
rect 5478 6344 5486 6379
rect 5534 6344 5542 6379
rect 5417 6338 5457 6344
rect 5417 6336 5429 6338
rect 5135 6306 5182 6312
rect 5135 6304 5143 6306
rect 5171 6304 5182 6306
rect 5235 6306 5282 6312
rect 5235 6304 5243 6306
rect 5271 6304 5282 6306
rect 5335 6306 5382 6312
rect 5335 6304 5343 6306
rect 5371 6304 5382 6306
rect 5563 6338 5603 6344
rect 5591 6336 5603 6338
rect 5636 6304 5644 6387
rect 5836 6381 5844 6409
rect 5894 6393 5902 6436
rect 5738 6344 5746 6379
rect 5996 6401 6004 6456
rect 6027 6437 6043 6443
rect 5677 6338 5717 6344
rect 5677 6336 5689 6338
rect 5838 6312 5845 6367
rect 5894 6344 5902 6379
rect 5798 6306 5845 6312
rect 5798 6304 5809 6306
rect 5837 6304 5845 6306
rect 5923 6338 5963 6344
rect 5951 6336 5963 6338
rect 5996 6304 6004 6387
rect 6037 6363 6043 6437
rect 6054 6436 6080 6447
rect 6054 6393 6062 6436
rect 6155 6422 6163 6436
rect 6183 6436 6211 6442
rect 6171 6433 6223 6436
rect 6254 6436 6280 6447
rect 6338 6476 6350 6482
rect 6510 6476 6522 6482
rect 6155 6415 6180 6422
rect 6137 6397 6153 6403
rect 6027 6357 6043 6363
rect 6054 6344 6062 6379
rect 6083 6338 6123 6344
rect 6111 6336 6123 6338
rect 6137 6323 6143 6397
rect 6173 6393 6181 6415
rect 6254 6393 6262 6436
rect 6386 6418 6404 6420
rect 6374 6409 6404 6418
rect 6396 6381 6404 6409
rect 6456 6418 6474 6420
rect 6456 6409 6486 6418
rect 6537 6476 6549 6482
rect 6600 6476 6612 6482
rect 6656 6476 6668 6482
rect 6456 6381 6464 6409
rect 6556 6401 6564 6456
rect 6179 6344 6187 6379
rect 6254 6344 6262 6379
rect 6137 6317 6153 6323
rect 6283 6338 6323 6344
rect 6311 6336 6323 6338
rect 6398 6312 6405 6367
rect 6358 6306 6405 6312
rect 6358 6304 6369 6306
rect 6397 6304 6405 6306
rect 6455 6312 6462 6367
rect 6455 6306 6502 6312
rect 6455 6304 6463 6306
rect 6491 6304 6502 6306
rect 6556 6304 6564 6387
rect 6633 6393 6640 6436
rect 6641 6356 6647 6379
rect 6641 6350 6668 6356
rect 6656 6344 6668 6350
rect 5022 6258 5034 6264
rect 5072 6258 5084 6264
rect 5151 6258 5163 6264
rect 5191 6258 5203 6264
rect 5251 6258 5263 6264
rect 5291 6258 5303 6264
rect 5351 6258 5363 6264
rect 5391 6258 5403 6264
rect 5437 6258 5449 6264
rect 5571 6258 5583 6264
rect 5651 6258 5663 6264
rect 5697 6258 5709 6264
rect 5777 6258 5789 6264
rect 5817 6258 5829 6264
rect 5931 6258 5943 6264
rect 6011 6258 6023 6264
rect 6091 6258 6103 6264
rect 6156 6258 6168 6264
rect 6206 6258 6218 6264
rect 6291 6258 6303 6264
rect 6337 6258 6349 6264
rect 6377 6258 6389 6264
rect 6471 6258 6483 6264
rect 6511 6258 6523 6264
rect 6609 6336 6637 6342
rect 6649 6264 6677 6270
rect 6537 6258 6549 6264
rect 6617 6258 6629 6264
rect 2127 6256 6736 6258
rect -62 6244 4 6256
rect -62 6242 1893 6244
rect -62 5778 -2 6242
rect 37 6236 49 6242
rect 95 6236 107 6242
rect 141 6236 153 6242
rect 207 6236 219 6242
rect 311 6236 323 6242
rect 371 6236 383 6242
rect 411 6236 423 6242
rect 67 6182 79 6216
rect 121 6190 133 6196
rect 175 6190 183 6196
rect 125 6178 147 6190
rect 175 6176 193 6190
rect 73 6158 79 6176
rect 97 6166 127 6172
rect 175 6170 183 6176
rect 17 6093 25 6156
rect 39 6144 53 6152
rect 73 6152 113 6158
rect 33 6093 47 6107
rect 17 6079 33 6093
rect 107 6080 113 6152
rect 121 6152 127 6166
rect 145 6162 183 6170
rect 437 6236 449 6242
rect 531 6236 543 6242
rect 571 6236 583 6242
rect 331 6162 343 6164
rect 303 6156 343 6162
rect 121 6146 165 6152
rect 177 6148 239 6156
rect 167 6107 194 6114
rect 214 6096 220 6101
rect 186 6088 220 6096
rect 174 6080 181 6088
rect 17 6064 25 6079
rect 107 6074 181 6080
rect 107 6072 113 6074
rect 174 6068 181 6074
rect 67 6050 78 6058
rect 71 6044 78 6050
rect 128 6056 149 6063
rect 233 6064 239 6148
rect 274 6121 282 6156
rect 395 6141 403 6196
rect 602 6236 614 6242
rect 652 6236 664 6242
rect 460 6149 477 6156
rect 128 6044 135 6056
rect 193 6044 200 6050
rect 187 6038 200 6044
rect 274 6064 282 6107
rect 395 6078 403 6127
rect 460 6101 467 6149
rect 555 6141 563 6196
rect 716 6236 728 6242
rect 766 6236 778 6242
rect 797 6236 809 6242
rect 931 6236 943 6242
rect 1007 6236 1019 6242
rect 1111 6236 1123 6242
rect 951 6162 963 6164
rect 923 6156 963 6162
rect 1137 6236 1149 6242
rect 1236 6236 1248 6242
rect 1286 6236 1298 6242
rect 1351 6236 1363 6242
rect 1411 6236 1423 6242
rect 1039 6157 1043 6166
rect 379 6072 403 6078
rect 379 6064 391 6072
rect 274 6053 300 6064
rect 460 6044 467 6087
rect 555 6078 563 6127
rect 633 6121 641 6156
rect 739 6121 747 6156
rect 820 6149 837 6156
rect 639 6085 647 6107
rect 733 6085 741 6107
rect 820 6101 827 6149
rect 894 6121 902 6156
rect 977 6148 985 6156
rect 977 6140 1013 6148
rect 640 6078 665 6085
rect 539 6072 563 6078
rect 539 6064 551 6072
rect 597 6064 649 6067
rect 39 6018 51 6024
rect 97 6018 109 6024
rect 145 6018 157 6024
rect 207 6018 219 6024
rect 278 6018 290 6024
rect 328 6018 340 6024
rect 409 6018 421 6024
rect 609 6058 637 6064
rect 657 6064 665 6078
rect 715 6078 740 6085
rect 715 6064 723 6078
rect 731 6064 783 6067
rect 743 6058 771 6064
rect 820 6044 827 6087
rect 894 6064 902 6107
rect 1018 6084 1024 6139
rect 1034 6113 1043 6157
rect 1096 6113 1104 6196
rect 1437 6236 1449 6242
rect 1517 6236 1529 6242
rect 1597 6236 1609 6242
rect 1657 6236 1669 6242
rect 1737 6236 1749 6242
rect 1822 6236 1834 6242
rect 1872 6236 1884 6242
rect 1160 6149 1177 6156
rect 1160 6101 1167 6149
rect 1259 6121 1267 6156
rect 1003 6072 1013 6078
rect 894 6053 920 6064
rect 437 6018 449 6024
rect 477 6018 489 6024
rect 569 6018 581 6024
rect 617 6018 629 6024
rect 751 6018 763 6024
rect 797 6018 809 6024
rect 837 6018 849 6024
rect 1003 6044 1009 6072
rect 1040 6064 1047 6099
rect 898 6018 910 6024
rect 948 6018 960 6024
rect 1096 6044 1104 6099
rect 1160 6044 1167 6087
rect 1253 6085 1261 6107
rect 1336 6113 1344 6196
rect 1396 6113 1404 6196
rect 1460 6149 1477 6156
rect 1540 6149 1557 6156
rect 1235 6078 1260 6085
rect 1235 6064 1243 6078
rect 977 6018 985 6024
rect 1017 6018 1029 6024
rect 1111 6018 1123 6024
rect 1251 6064 1303 6067
rect 1263 6058 1291 6064
rect 1336 6044 1344 6099
rect 1460 6101 1467 6149
rect 1540 6101 1547 6149
rect 1616 6113 1624 6196
rect 1907 6242 6736 6244
rect 1917 6236 1929 6242
rect 2031 6236 2043 6242
rect 2077 6236 2089 6242
rect 2156 6236 2168 6242
rect 2206 6236 2218 6242
rect 1680 6149 1697 6156
rect 1760 6149 1777 6156
rect 1396 6044 1404 6099
rect 1680 6101 1687 6149
rect 1460 6044 1467 6087
rect 1540 6044 1547 6087
rect 1616 6044 1624 6099
rect 1680 6044 1687 6087
rect 1717 6083 1723 6113
rect 1760 6101 1767 6149
rect 1707 6077 1723 6083
rect 1760 6044 1767 6087
rect 1797 6083 1803 6133
rect 1853 6121 1861 6156
rect 1936 6113 1944 6196
rect 2051 6162 2063 6164
rect 2023 6156 2063 6162
rect 1994 6121 2002 6156
rect 1859 6085 1867 6107
rect 2096 6113 2104 6196
rect 2237 6236 2249 6242
rect 2316 6236 2328 6242
rect 2366 6236 2378 6242
rect 2431 6236 2443 6242
rect 2471 6236 2483 6242
rect 2551 6236 2563 6242
rect 2651 6236 2663 6242
rect 2711 6236 2723 6242
rect 2751 6236 2763 6242
rect 2851 6236 2863 6242
rect 2931 6236 2943 6242
rect 1777 6077 1803 6083
rect 1860 6078 1885 6085
rect 1777 6067 1783 6077
rect 1817 6064 1869 6067
rect 1137 6018 1149 6024
rect 1177 6018 1189 6024
rect 1271 6018 1283 6024
rect 1351 6018 1363 6024
rect 1411 6018 1423 6024
rect 1437 6018 1449 6024
rect 1477 6018 1489 6024
rect 1517 6018 1529 6024
rect 1557 6018 1569 6024
rect 1597 6018 1609 6024
rect 1657 6018 1669 6024
rect 1697 6018 1709 6024
rect 1829 6058 1857 6064
rect 1877 6064 1885 6078
rect 1936 6044 1944 6099
rect 1994 6064 2002 6107
rect 1994 6053 2020 6064
rect 2096 6044 2104 6099
rect 2137 6087 2143 6153
rect 2179 6121 2187 6156
rect 2173 6085 2181 6107
rect 2256 6113 2264 6196
rect 2297 6177 2313 6183
rect 2297 6103 2303 6177
rect 2415 6194 2423 6196
rect 2451 6194 2462 6196
rect 2415 6188 2462 6194
rect 2339 6121 2347 6156
rect 2415 6133 2422 6188
rect 2571 6162 2583 6164
rect 2543 6156 2583 6162
rect 2695 6194 2703 6196
rect 2731 6194 2742 6196
rect 2695 6188 2742 6194
rect 2155 6078 2180 6085
rect 2155 6064 2163 6078
rect 1737 6018 1749 6024
rect 1777 6018 1789 6024
rect 1837 6018 1849 6024
rect 1917 6018 1929 6024
rect 1998 6018 2010 6024
rect 2048 6018 2060 6024
rect 2171 6064 2223 6067
rect 2183 6058 2211 6064
rect 2256 6044 2264 6099
rect 2297 6097 2313 6103
rect 2333 6085 2341 6107
rect 2514 6121 2522 6156
rect 2623 6149 2640 6156
rect 2416 6091 2424 6119
rect 2315 6078 2340 6085
rect 2416 6082 2446 6091
rect 2416 6080 2434 6082
rect 2315 6064 2323 6078
rect 2331 6064 2383 6067
rect 2343 6058 2371 6064
rect 2514 6064 2522 6107
rect 2633 6101 2640 6149
rect 2695 6133 2702 6188
rect 2803 6230 2831 6236
rect 2843 6158 2871 6164
rect 2957 6236 2969 6242
rect 2997 6236 3009 6242
rect 3111 6236 3123 6242
rect 3191 6236 3203 6242
rect 3231 6236 3243 6242
rect 3311 6236 3323 6242
rect 3391 6236 3403 6242
rect 3451 6236 3463 6242
rect 3491 6236 3503 6242
rect 2812 6150 2824 6156
rect 2812 6144 2839 6150
rect 2833 6121 2839 6144
rect 2696 6091 2704 6119
rect 2514 6053 2540 6064
rect 2077 6018 2089 6024
rect 2191 6018 2203 6024
rect 2237 6018 2249 6024
rect 2351 6018 2363 6024
rect 2470 6018 2482 6024
rect 2633 6044 2640 6087
rect 2696 6082 2726 6091
rect 2696 6080 2714 6082
rect 2518 6018 2530 6024
rect 2568 6018 2580 6024
rect 2840 6064 2847 6107
rect 2916 6113 2924 6196
rect 2978 6194 2989 6196
rect 3017 6194 3025 6196
rect 2978 6188 3025 6194
rect 3018 6133 3025 6188
rect 3131 6162 3143 6164
rect 3103 6156 3143 6162
rect 3175 6194 3183 6196
rect 3211 6194 3222 6196
rect 3175 6188 3222 6194
rect 3074 6121 3082 6156
rect 3175 6133 3182 6188
rect 3331 6162 3343 6164
rect 3303 6156 3343 6162
rect 2611 6018 2623 6024
rect 2651 6018 2663 6024
rect 2750 6018 2762 6024
rect 2916 6044 2924 6099
rect 3016 6091 3024 6119
rect 3274 6121 3282 6156
rect 2812 6018 2824 6024
rect 2868 6018 2880 6024
rect 2931 6018 2943 6024
rect 2994 6082 3024 6091
rect 3006 6080 3024 6082
rect 3074 6064 3082 6107
rect 3176 6091 3184 6119
rect 3376 6113 3384 6196
rect 3435 6194 3443 6196
rect 3517 6236 3529 6242
rect 3557 6236 3569 6242
rect 3617 6236 3629 6242
rect 3697 6236 3709 6242
rect 3791 6236 3803 6242
rect 3831 6236 3843 6242
rect 3471 6194 3482 6196
rect 3435 6188 3482 6194
rect 3538 6194 3549 6196
rect 3577 6194 3585 6196
rect 3538 6188 3585 6194
rect 3435 6133 3442 6188
rect 3578 6133 3585 6188
rect 3176 6082 3206 6091
rect 3176 6080 3194 6082
rect 3074 6053 3100 6064
rect 3274 6064 3282 6107
rect 3274 6053 3300 6064
rect 2958 6018 2970 6024
rect 3078 6018 3090 6024
rect 3128 6018 3140 6024
rect 3230 6018 3242 6024
rect 3376 6044 3384 6099
rect 3436 6091 3444 6119
rect 3576 6091 3584 6119
rect 3436 6082 3466 6091
rect 3436 6080 3454 6082
rect 3278 6018 3290 6024
rect 3328 6018 3340 6024
rect 3391 6018 3403 6024
rect 3490 6018 3502 6024
rect 3554 6082 3584 6091
rect 3597 6087 3603 6153
rect 3636 6113 3644 6196
rect 3677 6162 3689 6164
rect 3677 6156 3717 6162
rect 3857 6236 3869 6242
rect 3897 6236 3909 6242
rect 3956 6236 3968 6242
rect 4006 6236 4018 6242
rect 3738 6121 3746 6156
rect 3815 6141 3823 6196
rect 3877 6141 3885 6196
rect 4042 6236 4054 6242
rect 4092 6236 4104 6242
rect 4191 6236 4203 6242
rect 4217 6236 4229 6242
rect 4291 6236 4303 6242
rect 4331 6236 4343 6242
rect 4357 6236 4369 6242
rect 4401 6236 4413 6242
rect 4476 6236 4488 6242
rect 4526 6236 4538 6242
rect 4611 6236 4623 6242
rect 4657 6236 4669 6242
rect 4697 6236 4709 6242
rect 4811 6236 4823 6242
rect 4891 6236 4903 6242
rect 4931 6236 4943 6242
rect 3566 6080 3584 6082
rect 3636 6044 3644 6099
rect 3738 6064 3746 6107
rect 3815 6078 3823 6127
rect 3720 6053 3746 6064
rect 3799 6072 3823 6078
rect 3877 6078 3885 6127
rect 3979 6121 3987 6156
rect 4073 6121 4081 6156
rect 4163 6149 4180 6156
rect 3973 6085 3981 6107
rect 4079 6085 4087 6107
rect 4173 6101 4180 6149
rect 4236 6113 4244 6196
rect 4315 6141 4323 6196
rect 3955 6078 3980 6085
rect 4080 6078 4105 6085
rect 3877 6072 3901 6078
rect 3799 6064 3811 6072
rect 3889 6064 3901 6072
rect 3955 6064 3963 6078
rect 3518 6018 3530 6024
rect 3617 6018 3629 6024
rect 3680 6018 3692 6024
rect 3730 6018 3742 6024
rect 3829 6018 3841 6024
rect 3971 6064 4023 6067
rect 3983 6058 4011 6064
rect 4037 6064 4089 6067
rect 4049 6058 4077 6064
rect 4097 6064 4105 6078
rect 4173 6044 4180 6087
rect 4236 6044 4244 6099
rect 4315 6078 4323 6127
rect 4378 6082 4386 6196
rect 4678 6194 4689 6196
rect 4717 6194 4725 6196
rect 4678 6188 4725 6194
rect 4631 6162 4643 6164
rect 4603 6156 4643 6162
rect 4421 6121 4429 6156
rect 4499 6121 4507 6156
rect 4574 6121 4582 6156
rect 4718 6133 4725 6188
rect 4831 6162 4843 6164
rect 4803 6156 4843 6162
rect 4875 6194 4883 6196
rect 4957 6236 4969 6242
rect 4997 6236 5009 6242
rect 5076 6236 5088 6242
rect 5126 6236 5138 6242
rect 4911 6194 4922 6196
rect 4875 6188 4922 6194
rect 4978 6194 4989 6196
rect 5017 6194 5025 6196
rect 4978 6188 5025 6194
rect 4427 6107 4429 6121
rect 4299 6072 4323 6078
rect 4357 6074 4395 6082
rect 4299 6064 4311 6072
rect 4357 6064 4369 6074
rect 4421 6064 4429 6107
rect 4493 6085 4501 6107
rect 4774 6121 4782 6156
rect 4875 6133 4882 6188
rect 4475 6078 4500 6085
rect 4475 6064 4483 6078
rect 3859 6018 3871 6024
rect 3991 6018 4003 6024
rect 4057 6018 4069 6024
rect 4151 6018 4163 6024
rect 4191 6018 4203 6024
rect 4419 6054 4429 6064
rect 4491 6064 4543 6067
rect 4503 6058 4531 6064
rect 4574 6064 4582 6107
rect 4716 6091 4724 6119
rect 5018 6133 5025 6188
rect 5171 6236 5183 6242
rect 5211 6236 5223 6242
rect 5237 6236 5249 6242
rect 5281 6236 5293 6242
rect 5342 6236 5354 6242
rect 5392 6236 5404 6242
rect 5491 6236 5503 6242
rect 5571 6236 5583 6242
rect 5611 6236 5623 6242
rect 5099 6121 5107 6156
rect 5195 6141 5203 6196
rect 4574 6053 4600 6064
rect 4217 6018 4229 6024
rect 4329 6018 4341 6024
rect 4387 6018 4399 6024
rect 4511 6018 4523 6024
rect 4578 6018 4590 6024
rect 4628 6018 4640 6024
rect 4694 6082 4724 6091
rect 4706 6080 4724 6082
rect 4774 6064 4782 6107
rect 4876 6091 4884 6119
rect 5016 6091 5024 6119
rect 4876 6082 4906 6091
rect 4876 6080 4894 6082
rect 4774 6053 4800 6064
rect 4658 6018 4670 6024
rect 4778 6018 4790 6024
rect 4828 6018 4840 6024
rect 4930 6018 4942 6024
rect 4994 6082 5024 6091
rect 5093 6085 5101 6107
rect 5006 6080 5024 6082
rect 5075 6078 5100 6085
rect 5195 6078 5203 6127
rect 5258 6082 5266 6196
rect 5511 6162 5523 6164
rect 5483 6156 5523 6162
rect 5555 6194 5563 6196
rect 5637 6236 5649 6242
rect 5677 6236 5689 6242
rect 5791 6236 5803 6242
rect 5837 6236 5849 6242
rect 5877 6236 5889 6242
rect 5942 6236 5954 6242
rect 5992 6236 6004 6242
rect 5591 6194 5602 6196
rect 5555 6188 5602 6194
rect 5658 6194 5669 6196
rect 5697 6194 5705 6196
rect 5658 6188 5705 6194
rect 5301 6121 5309 6156
rect 5373 6121 5381 6156
rect 5454 6121 5462 6156
rect 5555 6133 5562 6188
rect 5307 6107 5309 6121
rect 5075 6064 5083 6078
rect 5179 6072 5203 6078
rect 5237 6074 5275 6082
rect 5091 6064 5143 6067
rect 5103 6058 5131 6064
rect 5179 6064 5191 6072
rect 5237 6064 5249 6074
rect 5301 6064 5309 6107
rect 5698 6133 5705 6188
rect 5858 6194 5869 6196
rect 5897 6194 5905 6196
rect 5858 6188 5905 6194
rect 5811 6162 5823 6164
rect 5783 6156 5823 6162
rect 5754 6121 5762 6156
rect 5898 6133 5905 6188
rect 6042 6236 6054 6242
rect 6092 6236 6104 6242
rect 6137 6236 6149 6242
rect 6177 6236 6189 6242
rect 6237 6236 6249 6242
rect 6277 6236 6289 6242
rect 6371 6236 6383 6242
rect 6411 6236 6423 6242
rect 6491 6236 6503 6242
rect 6537 6236 6549 6242
rect 6597 6236 6609 6242
rect 6158 6194 6169 6196
rect 6197 6194 6205 6196
rect 6158 6188 6205 6194
rect 6258 6194 6269 6196
rect 6297 6194 6305 6196
rect 6258 6188 6305 6194
rect 5379 6085 5387 6107
rect 5380 6078 5405 6085
rect 5299 6054 5309 6064
rect 5337 6064 5389 6067
rect 5349 6058 5377 6064
rect 5397 6064 5405 6078
rect 5454 6064 5462 6107
rect 5556 6091 5564 6119
rect 5696 6091 5704 6119
rect 5973 6121 5981 6156
rect 6073 6121 6081 6156
rect 6198 6133 6205 6188
rect 6217 6177 6233 6183
rect 5556 6082 5586 6091
rect 5556 6080 5574 6082
rect 5454 6053 5480 6064
rect 4958 6018 4970 6024
rect 5111 6018 5123 6024
rect 5209 6018 5221 6024
rect 5267 6018 5279 6024
rect 5357 6018 5369 6024
rect 5458 6018 5470 6024
rect 5508 6018 5520 6024
rect 5610 6018 5622 6024
rect 5674 6082 5704 6091
rect 5686 6080 5704 6082
rect 5754 6064 5762 6107
rect 5896 6091 5904 6119
rect 5754 6053 5780 6064
rect 5638 6018 5650 6024
rect 5758 6018 5770 6024
rect 5808 6018 5820 6024
rect 5874 6082 5904 6091
rect 5979 6085 5987 6107
rect 6079 6085 6087 6107
rect 6196 6091 6204 6119
rect 6217 6103 6223 6177
rect 6298 6133 6305 6188
rect 6355 6194 6363 6196
rect 6391 6194 6402 6196
rect 6355 6188 6402 6194
rect 6355 6133 6362 6188
rect 6511 6162 6523 6164
rect 6483 6156 6523 6162
rect 6454 6121 6462 6156
rect 6217 6097 6233 6103
rect 6296 6091 6304 6119
rect 5886 6080 5904 6082
rect 5980 6078 6005 6085
rect 6080 6078 6105 6085
rect 5937 6064 5989 6067
rect 5949 6058 5977 6064
rect 5997 6064 6005 6078
rect 6037 6064 6089 6067
rect 6049 6058 6077 6064
rect 6097 6064 6105 6078
rect 6174 6082 6204 6091
rect 6186 6080 6204 6082
rect 6274 6082 6304 6091
rect 6286 6080 6304 6082
rect 6356 6091 6364 6119
rect 6556 6113 6564 6196
rect 6616 6113 6624 6196
rect 6356 6082 6386 6091
rect 6356 6080 6374 6082
rect 6454 6064 6462 6107
rect 6454 6053 6480 6064
rect 5838 6018 5850 6024
rect 5957 6018 5969 6024
rect 6057 6018 6069 6024
rect 6138 6018 6150 6024
rect 6238 6018 6250 6024
rect 6410 6018 6422 6024
rect 6556 6044 6564 6099
rect 6616 6044 6624 6099
rect 6458 6018 6470 6024
rect 6508 6018 6520 6024
rect 6537 6018 6549 6024
rect 6597 6018 6609 6024
rect 6742 6018 6802 6482
rect 4 6016 6802 6018
rect 6736 6004 6802 6016
rect 4 6002 6802 6004
rect 49 5996 61 6002
rect 99 5996 111 6002
rect 179 5996 191 6002
rect 278 5996 290 6002
rect 328 5996 340 6002
rect 409 5996 421 6002
rect 31 5913 39 5956
rect 71 5950 79 5976
rect 57 5944 79 5950
rect 129 5948 141 5956
rect 209 5948 221 5956
rect 57 5938 60 5944
rect 31 5899 33 5913
rect 31 5864 39 5899
rect 53 5882 60 5938
rect 117 5942 141 5948
rect 197 5942 221 5948
rect 274 5956 300 5967
rect 437 5996 449 6002
rect 511 5996 523 6002
rect 551 5996 563 6002
rect 577 5996 589 6002
rect 617 5996 629 6002
rect 677 5996 689 6002
rect 791 5996 803 6002
rect 117 5893 125 5942
rect 57 5876 60 5882
rect 197 5893 205 5942
rect 274 5913 282 5956
rect 379 5948 391 5956
rect 379 5942 403 5948
rect 57 5870 83 5876
rect 75 5824 83 5870
rect 117 5824 125 5879
rect 197 5824 205 5879
rect 274 5864 282 5899
rect 395 5893 403 5942
rect 456 5921 464 5976
rect 533 5933 540 5976
rect 600 5933 607 5976
rect 669 5956 697 5962
rect 657 5953 709 5956
rect 817 5996 829 6002
rect 857 5996 869 6002
rect 949 5996 961 6002
rect 1031 5996 1043 6002
rect 1077 5996 1089 6002
rect 1117 5996 1129 6002
rect 1191 5996 1203 6002
rect 1239 5996 1251 6002
rect 1297 5996 1309 6002
rect 1345 5996 1357 6002
rect 1407 5996 1419 6002
rect 1459 5996 1471 6002
rect 1610 5996 1622 6002
rect 1691 5996 1703 6002
rect 1751 5996 1763 6002
rect 1791 5996 1803 6002
rect 1890 5996 1902 6002
rect 49 5778 61 5784
rect 97 5778 109 5784
rect 137 5778 149 5784
rect 303 5858 343 5864
rect 331 5856 343 5858
rect 395 5824 403 5879
rect 456 5824 464 5907
rect 533 5871 540 5919
rect 523 5864 540 5871
rect 600 5871 607 5919
rect 637 5937 653 5943
rect 600 5864 617 5871
rect 637 5867 643 5937
rect 717 5942 725 5956
rect 700 5935 725 5942
rect 699 5913 707 5935
rect 776 5921 784 5976
rect 840 5933 847 5976
rect 919 5948 931 5956
rect 919 5942 943 5948
rect 177 5778 189 5784
rect 217 5778 229 5784
rect 311 5778 323 5784
rect 371 5778 383 5784
rect 411 5778 423 5784
rect 437 5778 449 5784
rect 551 5778 563 5784
rect 693 5864 701 5899
rect 776 5824 784 5907
rect 840 5871 847 5919
rect 935 5893 943 5942
rect 995 5942 1003 5956
rect 1023 5956 1051 5962
rect 1011 5953 1063 5956
rect 995 5935 1020 5942
rect 1013 5913 1021 5935
rect 1100 5933 1107 5976
rect 1176 5921 1184 5976
rect 1387 5976 1400 5982
rect 1271 5970 1278 5976
rect 1267 5962 1278 5970
rect 1328 5964 1335 5976
rect 1393 5970 1400 5976
rect 1217 5941 1225 5956
rect 1328 5957 1349 5964
rect 1307 5946 1313 5948
rect 1374 5946 1381 5952
rect 840 5864 857 5871
rect 577 5778 589 5784
rect 662 5778 674 5784
rect 712 5778 724 5784
rect 791 5778 803 5784
rect 935 5824 943 5879
rect 1019 5864 1027 5899
rect 1100 5871 1107 5919
rect 1217 5927 1233 5941
rect 1307 5940 1381 5946
rect 1100 5864 1117 5871
rect 817 5778 829 5784
rect 911 5778 923 5784
rect 951 5778 963 5784
rect 996 5778 1008 5784
rect 1046 5778 1058 5784
rect 1176 5824 1184 5907
rect 1217 5864 1225 5927
rect 1233 5913 1247 5927
rect 1239 5868 1253 5876
rect 1307 5868 1313 5940
rect 1374 5932 1381 5940
rect 1386 5924 1420 5932
rect 1414 5919 1420 5924
rect 1367 5906 1394 5913
rect 1273 5862 1313 5868
rect 1321 5868 1365 5874
rect 1273 5844 1279 5862
rect 1321 5854 1327 5868
rect 1433 5872 1439 5956
rect 1489 5948 1501 5956
rect 1477 5942 1501 5948
rect 1477 5893 1485 5942
rect 1556 5938 1574 5940
rect 1556 5929 1586 5938
rect 1655 5942 1663 5956
rect 1683 5956 1711 5962
rect 1671 5953 1723 5956
rect 1655 5935 1680 5942
rect 1556 5901 1564 5929
rect 1673 5913 1681 5935
rect 1773 5933 1780 5976
rect 1836 5938 1854 5940
rect 1377 5864 1439 5872
rect 1297 5848 1327 5854
rect 1345 5850 1383 5858
rect 1375 5844 1383 5850
rect 1267 5804 1279 5838
rect 1325 5830 1347 5842
rect 1375 5830 1393 5844
rect 1321 5824 1333 5830
rect 1375 5824 1383 5830
rect 1477 5824 1485 5879
rect 1555 5832 1562 5887
rect 1637 5843 1643 5913
rect 1836 5929 1866 5938
rect 1917 5996 1929 6002
rect 2031 5996 2043 6002
rect 2078 5996 2090 6002
rect 2198 5996 2210 6002
rect 2248 5996 2260 6002
rect 2297 5996 2309 6002
rect 2429 5996 2441 6002
rect 2530 5996 2542 6002
rect 1679 5864 1687 5899
rect 1773 5871 1780 5919
rect 1836 5901 1844 5929
rect 1936 5921 1944 5976
rect 1995 5942 2003 5956
rect 2023 5956 2051 5962
rect 2011 5953 2063 5956
rect 1995 5935 2020 5942
rect 2194 5956 2220 5967
rect 2289 5956 2317 5962
rect 2126 5938 2144 5940
rect 1977 5917 1993 5923
rect 1763 5864 1780 5871
rect 1627 5837 1643 5843
rect 1555 5826 1602 5832
rect 1555 5824 1563 5826
rect 1591 5824 1602 5826
rect 1077 5778 1089 5784
rect 1191 5778 1203 5784
rect 1237 5778 1249 5784
rect 1295 5778 1307 5784
rect 1341 5778 1353 5784
rect 1407 5778 1419 5784
rect 1457 5778 1469 5784
rect 1497 5778 1509 5784
rect 1571 5778 1583 5784
rect 1611 5778 1623 5784
rect -62 5776 1633 5778
rect 1656 5778 1668 5784
rect 1706 5778 1718 5784
rect 1647 5776 1733 5778
rect 1835 5832 1842 5887
rect 1835 5826 1882 5832
rect 1835 5824 1843 5826
rect 1871 5824 1882 5826
rect 1936 5824 1944 5907
rect 1957 5847 1963 5913
rect 1977 5843 1983 5917
rect 2013 5913 2021 5935
rect 2114 5929 2144 5938
rect 2136 5901 2144 5929
rect 2194 5913 2202 5956
rect 2277 5953 2329 5956
rect 2337 5942 2345 5956
rect 2399 5948 2411 5956
rect 2399 5942 2423 5948
rect 2320 5935 2345 5942
rect 2019 5864 2027 5899
rect 2319 5913 2327 5935
rect 1977 5837 1993 5843
rect 1791 5778 1803 5784
rect 1851 5778 1863 5784
rect 1891 5778 1903 5784
rect 2138 5832 2145 5887
rect 2194 5864 2202 5899
rect 2313 5864 2321 5899
rect 2415 5893 2423 5942
rect 2476 5938 2494 5940
rect 2476 5929 2506 5938
rect 2578 5996 2590 6002
rect 2628 5996 2640 6002
rect 2574 5956 2600 5967
rect 2659 5996 2671 6002
rect 2810 5996 2822 6002
rect 2910 5996 2922 6002
rect 3010 5996 3022 6002
rect 3110 5996 3122 6002
rect 2476 5901 2484 5929
rect 2574 5913 2582 5956
rect 2689 5948 2701 5956
rect 2677 5942 2701 5948
rect 2098 5826 2145 5832
rect 2098 5824 2109 5826
rect 1917 5778 1929 5784
rect 1996 5778 2008 5784
rect 2046 5778 2058 5784
rect 2137 5824 2145 5826
rect 2223 5858 2263 5864
rect 2251 5856 2263 5858
rect 2415 5824 2423 5879
rect 2475 5832 2482 5887
rect 2574 5864 2582 5899
rect 2677 5893 2685 5942
rect 2756 5938 2774 5940
rect 2756 5929 2786 5938
rect 2856 5938 2874 5940
rect 2856 5929 2886 5938
rect 2937 5957 2953 5963
rect 2756 5901 2764 5929
rect 2856 5901 2864 5929
rect 2937 5923 2943 5957
rect 2897 5917 2943 5923
rect 2956 5938 2974 5940
rect 2956 5929 2986 5938
rect 3056 5938 3074 5940
rect 3056 5929 3086 5938
rect 3138 5996 3150 6002
rect 3291 5996 3303 6002
rect 3357 5996 3369 6002
rect 3458 5996 3470 6002
rect 3508 5996 3520 6002
rect 3591 5996 3603 6002
rect 3710 5996 3722 6002
rect 3255 5942 3263 5956
rect 3283 5956 3311 5962
rect 3271 5953 3323 5956
rect 3349 5956 3377 5962
rect 3337 5953 3389 5956
rect 3454 5956 3480 5967
rect 3397 5942 3405 5956
rect 3186 5938 3204 5940
rect 3174 5929 3204 5938
rect 3255 5935 3280 5942
rect 3380 5935 3405 5942
rect 2897 5907 2903 5917
rect 2475 5826 2522 5832
rect 2475 5824 2483 5826
rect 2077 5778 2089 5784
rect 2117 5778 2129 5784
rect 2231 5778 2243 5784
rect 2282 5778 2294 5784
rect 2332 5778 2344 5784
rect 2511 5824 2522 5826
rect 2603 5858 2643 5864
rect 2631 5856 2643 5858
rect 2677 5824 2685 5879
rect 2755 5832 2762 5887
rect 2956 5901 2964 5929
rect 3056 5901 3064 5929
rect 3107 5917 3133 5923
rect 3196 5901 3204 5929
rect 3273 5913 3281 5935
rect 2855 5832 2862 5887
rect 2955 5832 2962 5887
rect 3055 5832 3062 5887
rect 3379 5913 3387 5935
rect 3454 5913 3462 5956
rect 3555 5942 3563 5956
rect 3583 5956 3611 5962
rect 3571 5953 3623 5956
rect 3555 5935 3580 5942
rect 3656 5938 3674 5940
rect 3573 5913 3581 5935
rect 3656 5929 3686 5938
rect 3740 5996 3752 6002
rect 3790 5996 3802 6002
rect 3910 5996 3922 6002
rect 3780 5956 3806 5967
rect 3656 5901 3664 5929
rect 3798 5913 3806 5956
rect 3856 5938 3874 5940
rect 3856 5929 3886 5938
rect 3958 5996 3970 6002
rect 4008 5996 4020 6002
rect 4110 5996 4122 6002
rect 3954 5956 3980 5967
rect 3198 5832 3205 5887
rect 3279 5864 3287 5899
rect 3373 5864 3381 5899
rect 3454 5864 3462 5899
rect 3579 5864 3587 5899
rect 3856 5901 3864 5929
rect 3954 5913 3962 5956
rect 4056 5938 4074 5940
rect 2755 5826 2802 5832
rect 2755 5824 2763 5826
rect 2791 5824 2802 5826
rect 2855 5826 2902 5832
rect 2855 5824 2863 5826
rect 2891 5824 2902 5826
rect 2955 5826 3002 5832
rect 2955 5824 2963 5826
rect 2991 5824 3002 5826
rect 3055 5826 3102 5832
rect 3055 5824 3063 5826
rect 3091 5824 3102 5826
rect 3158 5826 3205 5832
rect 3158 5824 3169 5826
rect 2391 5778 2403 5784
rect 2431 5778 2443 5784
rect 2491 5778 2503 5784
rect 2531 5778 2543 5784
rect 2611 5778 2623 5784
rect 2657 5778 2669 5784
rect 2697 5778 2709 5784
rect 2771 5778 2783 5784
rect 2811 5778 2823 5784
rect 2871 5778 2883 5784
rect 2911 5778 2923 5784
rect 2971 5778 2983 5784
rect 3011 5778 3023 5784
rect 3071 5778 3083 5784
rect 3111 5778 3123 5784
rect 3197 5824 3205 5826
rect 3137 5778 3149 5784
rect 3177 5778 3189 5784
rect 3256 5778 3268 5784
rect 3306 5778 3318 5784
rect 3483 5858 3523 5864
rect 3511 5856 3523 5858
rect 3655 5832 3662 5887
rect 3798 5864 3806 5899
rect 4056 5929 4086 5938
rect 4158 5996 4170 6002
rect 4208 5996 4220 6002
rect 4154 5956 4180 5967
rect 4238 5996 4250 6002
rect 4339 5996 4351 6002
rect 4471 5996 4483 6002
rect 4531 5996 4543 6002
rect 4571 5996 4583 6002
rect 4627 5996 4639 6002
rect 4718 5996 4730 6002
rect 4768 5996 4780 6002
rect 4056 5901 4064 5929
rect 4154 5913 4162 5956
rect 4369 5948 4381 5956
rect 4357 5942 4381 5948
rect 4435 5942 4443 5956
rect 4463 5956 4491 5962
rect 4451 5953 4503 5956
rect 4286 5938 4304 5940
rect 4097 5907 4103 5913
rect 3737 5858 3777 5864
rect 3737 5856 3749 5858
rect 3655 5826 3702 5832
rect 3655 5824 3663 5826
rect 3691 5824 3702 5826
rect 3855 5832 3862 5887
rect 3954 5864 3962 5899
rect 4274 5929 4304 5938
rect 4296 5901 4304 5929
rect 3987 5877 4013 5883
rect 3855 5826 3902 5832
rect 3855 5824 3863 5826
rect 3891 5824 3902 5826
rect 3983 5858 4023 5864
rect 4011 5856 4023 5858
rect 4055 5832 4062 5887
rect 4154 5864 4162 5899
rect 4357 5893 4365 5942
rect 4435 5935 4460 5942
rect 4453 5913 4461 5935
rect 4553 5933 4560 5976
rect 4659 5956 4669 5966
rect 4597 5946 4609 5956
rect 4597 5938 4635 5946
rect 4055 5826 4102 5832
rect 4055 5824 4063 5826
rect 4091 5824 4102 5826
rect 4183 5858 4223 5864
rect 4211 5856 4223 5858
rect 4298 5832 4305 5887
rect 4258 5826 4305 5832
rect 4258 5824 4269 5826
rect 4297 5824 4305 5826
rect 4357 5824 4365 5879
rect 4459 5864 4467 5899
rect 4553 5871 4560 5919
rect 4543 5864 4560 5871
rect 3342 5778 3354 5784
rect 3392 5778 3404 5784
rect 3491 5778 3503 5784
rect 3556 5778 3568 5784
rect 3606 5778 3618 5784
rect 3671 5778 3683 5784
rect 3711 5778 3723 5784
rect 3757 5778 3769 5784
rect 3871 5778 3883 5784
rect 3911 5778 3923 5784
rect 3991 5778 4003 5784
rect 4071 5778 4083 5784
rect 4111 5778 4123 5784
rect 4191 5778 4203 5784
rect 4237 5778 4249 5784
rect 4277 5778 4289 5784
rect 4337 5778 4349 5784
rect 4377 5778 4389 5784
rect 4618 5824 4626 5938
rect 4661 5913 4669 5956
rect 4714 5956 4740 5967
rect 4799 5996 4811 6002
rect 4911 5996 4923 6002
rect 5010 5996 5022 6002
rect 4714 5913 4722 5956
rect 4829 5948 4841 5956
rect 4817 5942 4841 5948
rect 4667 5899 4669 5913
rect 4661 5864 4669 5899
rect 4714 5864 4722 5899
rect 4817 5893 4825 5942
rect 4896 5921 4904 5976
rect 4956 5938 4974 5940
rect 4956 5929 4986 5938
rect 5040 5996 5052 6002
rect 5090 5996 5102 6002
rect 5157 5996 5169 6002
rect 5257 5996 5269 6002
rect 5340 5996 5352 6002
rect 5396 5996 5408 6002
rect 5509 5996 5521 6002
rect 5080 5956 5106 5967
rect 4436 5778 4448 5784
rect 4486 5778 4498 5784
rect 4571 5778 4583 5784
rect 4743 5858 4783 5864
rect 4771 5856 4783 5858
rect 4817 5824 4825 5879
rect 4896 5824 4904 5907
rect 4956 5901 4964 5929
rect 5098 5913 5106 5956
rect 5149 5956 5177 5962
rect 5137 5953 5189 5956
rect 5249 5956 5277 5962
rect 5197 5942 5205 5956
rect 5237 5953 5289 5956
rect 5537 5996 5549 6002
rect 5670 5996 5682 6002
rect 5297 5942 5305 5956
rect 5180 5935 5205 5942
rect 5280 5935 5305 5942
rect 5179 5913 5187 5935
rect 5279 5913 5287 5935
rect 5373 5913 5380 5956
rect 5479 5948 5491 5956
rect 5479 5942 5503 5948
rect 4955 5832 4962 5887
rect 5098 5864 5106 5899
rect 5173 5864 5181 5899
rect 5273 5864 5281 5899
rect 5381 5876 5387 5899
rect 5495 5893 5503 5942
rect 5556 5921 5564 5976
rect 5597 5957 5613 5963
rect 5381 5870 5408 5876
rect 5396 5864 5408 5870
rect 5037 5858 5077 5864
rect 5037 5856 5049 5858
rect 4955 5826 5002 5832
rect 4955 5824 4963 5826
rect 4991 5824 5002 5826
rect 4597 5778 4609 5784
rect 4641 5778 4653 5784
rect 4751 5778 4763 5784
rect 4797 5778 4809 5784
rect 4837 5778 4849 5784
rect 4911 5778 4923 5784
rect 4971 5778 4983 5784
rect 5011 5778 5023 5784
rect 5057 5778 5069 5784
rect 5142 5778 5154 5784
rect 5192 5778 5204 5784
rect 5349 5856 5377 5862
rect 5389 5784 5417 5790
rect 5495 5824 5503 5879
rect 5556 5824 5564 5907
rect 5577 5847 5583 5933
rect 5597 5867 5603 5957
rect 5616 5938 5634 5940
rect 5616 5929 5646 5938
rect 5700 5996 5712 6002
rect 5750 5996 5762 6002
rect 5851 5996 5863 6002
rect 5917 5996 5929 6002
rect 6051 5996 6063 6002
rect 6100 5996 6112 6002
rect 6156 5996 6168 6002
rect 6269 5996 6281 6002
rect 6327 5996 6339 6002
rect 6417 5996 6429 6002
rect 6498 5996 6510 6002
rect 6599 5996 6611 6002
rect 5740 5956 5766 5967
rect 5616 5901 5624 5929
rect 5758 5913 5766 5956
rect 5815 5942 5823 5956
rect 5843 5956 5871 5962
rect 5831 5953 5883 5956
rect 5909 5956 5937 5962
rect 5897 5953 5949 5956
rect 5957 5942 5965 5956
rect 5815 5935 5840 5942
rect 5940 5935 5965 5942
rect 6015 5942 6023 5956
rect 6043 5956 6071 5962
rect 6359 5956 6369 5966
rect 6031 5953 6083 5956
rect 6015 5935 6040 5942
rect 5833 5913 5841 5935
rect 5939 5913 5947 5935
rect 6033 5913 6041 5935
rect 6133 5913 6140 5956
rect 6239 5948 6251 5956
rect 6239 5942 6263 5948
rect 5615 5832 5622 5887
rect 5707 5877 5733 5883
rect 5758 5864 5766 5899
rect 5839 5864 5847 5899
rect 5933 5864 5941 5899
rect 6039 5864 6047 5899
rect 6141 5876 6147 5899
rect 6255 5893 6263 5942
rect 6297 5946 6309 5956
rect 6297 5938 6335 5946
rect 6141 5870 6168 5876
rect 6156 5864 6168 5870
rect 5697 5858 5737 5864
rect 5697 5856 5709 5858
rect 5615 5826 5662 5832
rect 5615 5824 5623 5826
rect 5242 5778 5254 5784
rect 5292 5778 5304 5784
rect 5357 5778 5369 5784
rect 5471 5778 5483 5784
rect 5511 5778 5523 5784
rect 5651 5824 5662 5826
rect 5537 5778 5549 5784
rect 5631 5778 5643 5784
rect 5671 5778 5683 5784
rect 5717 5778 5729 5784
rect 5816 5778 5828 5784
rect 5866 5778 5878 5784
rect 5902 5778 5914 5784
rect 5952 5778 5964 5784
rect 6109 5856 6137 5862
rect 6149 5784 6177 5790
rect 6255 5824 6263 5879
rect 6318 5824 6326 5938
rect 6361 5913 6369 5956
rect 6409 5956 6437 5962
rect 6397 5953 6449 5956
rect 6457 5942 6465 5956
rect 6440 5935 6465 5942
rect 6629 5948 6641 5956
rect 6617 5942 6641 5948
rect 6546 5938 6564 5940
rect 6367 5899 6369 5913
rect 6439 5913 6447 5935
rect 6534 5929 6564 5938
rect 6361 5864 6369 5899
rect 6433 5864 6441 5899
rect 6016 5778 6028 5784
rect 6066 5778 6078 5784
rect 6117 5778 6129 5784
rect 6231 5778 6243 5784
rect 6271 5778 6283 5784
rect 6477 5843 6483 5913
rect 6556 5901 6564 5929
rect 6477 5837 6493 5843
rect 6558 5832 6565 5887
rect 6577 5863 6583 5893
rect 6617 5893 6625 5942
rect 6577 5857 6593 5863
rect 6518 5826 6565 5832
rect 6518 5824 6529 5826
rect 6297 5778 6309 5784
rect 6341 5778 6353 5784
rect 6402 5778 6414 5784
rect 6452 5778 6464 5784
rect 6557 5824 6565 5826
rect 6617 5824 6625 5879
rect 6497 5778 6509 5784
rect 6537 5778 6549 5784
rect 6597 5778 6609 5784
rect 6637 5778 6649 5784
rect 1747 5776 6736 5778
rect -62 5764 4 5776
rect -62 5762 6736 5764
rect -62 5298 -2 5762
rect 49 5756 61 5762
rect 129 5756 141 5762
rect 197 5756 209 5762
rect 255 5756 267 5762
rect 301 5756 313 5762
rect 367 5756 379 5762
rect 471 5756 483 5762
rect 517 5756 529 5762
rect 597 5756 609 5762
rect 637 5756 649 5762
rect 31 5641 39 5676
rect 75 5670 83 5716
rect 57 5664 83 5670
rect 57 5658 60 5664
rect 31 5627 33 5641
rect 31 5584 39 5627
rect 53 5602 60 5658
rect 111 5641 119 5676
rect 155 5670 163 5716
rect 137 5664 163 5670
rect 227 5702 239 5736
rect 281 5710 293 5716
rect 335 5710 343 5716
rect 285 5698 307 5710
rect 335 5696 353 5710
rect 233 5678 239 5696
rect 257 5686 287 5692
rect 335 5690 343 5696
rect 137 5658 140 5664
rect 111 5627 113 5641
rect 57 5596 60 5602
rect 57 5590 79 5596
rect 71 5564 79 5590
rect 111 5584 119 5627
rect 133 5602 140 5658
rect 137 5596 140 5602
rect 177 5613 185 5676
rect 199 5664 213 5672
rect 233 5672 273 5678
rect 193 5613 207 5627
rect 177 5599 193 5613
rect 267 5600 273 5672
rect 281 5672 287 5686
rect 305 5682 343 5690
rect 281 5666 325 5672
rect 337 5668 399 5676
rect 497 5682 509 5684
rect 497 5676 537 5682
rect 677 5756 689 5762
rect 721 5756 733 5762
rect 777 5756 789 5762
rect 817 5756 829 5762
rect 443 5669 460 5676
rect 327 5627 354 5634
rect 374 5616 380 5621
rect 346 5608 380 5616
rect 334 5600 341 5608
rect 137 5590 159 5596
rect 151 5564 159 5590
rect 177 5584 185 5599
rect 267 5594 341 5600
rect 267 5592 273 5594
rect 334 5588 341 5594
rect 227 5570 238 5578
rect 231 5564 238 5570
rect 288 5576 309 5583
rect 393 5584 399 5668
rect 288 5564 295 5576
rect 353 5564 360 5570
rect 347 5558 360 5564
rect 453 5621 460 5669
rect 558 5641 566 5676
rect 617 5661 625 5716
rect 453 5564 460 5607
rect 558 5584 566 5627
rect 617 5598 625 5647
rect 698 5602 706 5716
rect 857 5756 869 5762
rect 897 5756 909 5762
rect 937 5756 949 5762
rect 1017 5756 1029 5762
rect 1107 5756 1119 5762
rect 1177 5756 1189 5762
rect 1257 5756 1269 5762
rect 1317 5756 1329 5762
rect 1397 5756 1409 5762
rect 1477 5756 1489 5762
rect 1535 5756 1547 5762
rect 1581 5756 1593 5762
rect 1647 5756 1659 5762
rect 1697 5756 1709 5762
rect 1767 5756 1779 5762
rect 741 5641 749 5676
rect 797 5661 805 5716
rect 877 5661 885 5716
rect 960 5669 977 5676
rect 747 5627 749 5641
rect 617 5592 641 5598
rect 629 5584 641 5592
rect 49 5538 61 5544
rect 129 5538 141 5544
rect 199 5538 211 5544
rect 257 5538 269 5544
rect 305 5538 317 5544
rect 367 5538 379 5544
rect 431 5538 443 5544
rect 471 5538 483 5544
rect 540 5573 566 5584
rect 500 5538 512 5544
rect 550 5538 562 5544
rect 677 5594 715 5602
rect 677 5584 689 5594
rect 741 5584 749 5627
rect 797 5598 805 5647
rect 877 5598 885 5647
rect 960 5621 967 5669
rect 1036 5633 1044 5716
rect 1139 5677 1143 5686
rect 1077 5668 1085 5676
rect 1077 5660 1113 5668
rect 797 5592 821 5598
rect 877 5592 901 5598
rect 809 5584 821 5592
rect 889 5584 901 5592
rect 739 5574 749 5584
rect 960 5564 967 5607
rect 1036 5564 1044 5619
rect 1118 5604 1124 5659
rect 1134 5633 1143 5677
rect 1200 5669 1217 5676
rect 1200 5621 1207 5669
rect 1276 5633 1284 5716
rect 1340 5669 1357 5676
rect 1103 5592 1113 5598
rect 1103 5564 1109 5592
rect 1140 5584 1147 5619
rect 1340 5621 1347 5669
rect 1416 5633 1424 5716
rect 1507 5702 1519 5736
rect 1561 5710 1573 5716
rect 1615 5710 1623 5716
rect 1565 5698 1587 5710
rect 1615 5696 1633 5710
rect 1513 5678 1519 5696
rect 1537 5686 1567 5692
rect 1615 5690 1623 5696
rect 599 5538 611 5544
rect 707 5538 719 5544
rect 779 5538 791 5544
rect 859 5538 871 5544
rect 937 5538 949 5544
rect 977 5538 989 5544
rect 1200 5564 1207 5607
rect 1276 5564 1284 5619
rect 1340 5564 1347 5607
rect 1416 5564 1424 5619
rect 1457 5613 1465 5676
rect 1479 5664 1493 5672
rect 1513 5672 1553 5678
rect 1473 5613 1487 5627
rect 1457 5599 1473 5613
rect 1547 5600 1553 5672
rect 1561 5672 1567 5686
rect 1585 5682 1623 5690
rect 1836 5756 1848 5762
rect 1886 5756 1898 5762
rect 1931 5756 1943 5762
rect 1971 5756 1983 5762
rect 1997 5756 2009 5762
rect 2111 5756 2123 5762
rect 2157 5756 2169 5762
rect 2237 5756 2249 5762
rect 2277 5756 2289 5762
rect 2451 5756 2463 5762
rect 2511 5756 2523 5762
rect 2551 5756 2563 5762
rect 2611 5756 2623 5762
rect 2651 5756 2663 5762
rect 2711 5756 2723 5762
rect 2751 5756 2763 5762
rect 1561 5666 1605 5672
rect 1617 5668 1679 5676
rect 1607 5627 1634 5634
rect 1654 5616 1660 5621
rect 1626 5608 1660 5616
rect 1614 5600 1621 5608
rect 1457 5584 1465 5599
rect 1547 5594 1621 5600
rect 1547 5592 1553 5594
rect 1017 5538 1029 5544
rect 1077 5538 1085 5544
rect 1117 5538 1129 5544
rect 1177 5538 1189 5544
rect 1217 5538 1229 5544
rect 1257 5538 1269 5544
rect 1317 5538 1329 5544
rect 1357 5538 1369 5544
rect 1614 5588 1621 5594
rect 1507 5570 1518 5578
rect 1511 5564 1518 5570
rect 1568 5576 1589 5583
rect 1673 5584 1679 5668
rect 1737 5641 1745 5676
rect 1859 5641 1867 5676
rect 1955 5661 1963 5716
rect 1736 5601 1744 5627
rect 1853 5605 1861 5627
rect 1736 5594 1765 5601
rect 1568 5564 1575 5576
rect 1633 5564 1640 5570
rect 1627 5558 1640 5564
rect 1697 5584 1749 5586
rect 1759 5584 1765 5594
rect 1835 5598 1860 5605
rect 1955 5598 1963 5647
rect 2016 5633 2024 5716
rect 2131 5682 2143 5684
rect 2103 5676 2143 5682
rect 2327 5750 2379 5756
rect 2327 5748 2339 5750
rect 2074 5641 2082 5676
rect 2180 5669 2197 5676
rect 1835 5584 1843 5598
rect 1939 5592 1963 5598
rect 1709 5580 1737 5584
rect 1749 5544 1777 5550
rect 1851 5584 1903 5587
rect 1863 5578 1891 5584
rect 1939 5584 1951 5592
rect 2016 5564 2024 5619
rect 2074 5584 2082 5627
rect 2180 5621 2187 5669
rect 2257 5661 2265 5716
rect 2367 5748 2379 5750
rect 2351 5676 2359 5692
rect 2403 5750 2431 5756
rect 2411 5692 2423 5696
rect 2379 5688 2423 5692
rect 2367 5686 2423 5688
rect 2431 5690 2443 5696
rect 2471 5690 2483 5696
rect 2431 5684 2483 5690
rect 2351 5668 2374 5676
rect 2074 5573 2100 5584
rect 1397 5538 1409 5544
rect 1479 5538 1491 5544
rect 1537 5538 1549 5544
rect 1585 5538 1597 5544
rect 1647 5538 1659 5544
rect 1717 5538 1729 5544
rect 1871 5538 1883 5544
rect 1969 5538 1981 5544
rect 2180 5564 2187 5607
rect 2257 5598 2265 5647
rect 2366 5633 2374 5668
rect 2535 5661 2543 5716
rect 2595 5714 2603 5716
rect 2631 5714 2642 5716
rect 2595 5708 2642 5714
rect 2695 5714 2703 5716
rect 2777 5756 2789 5762
rect 2817 5756 2829 5762
rect 2862 5756 2874 5762
rect 2912 5756 2924 5762
rect 2991 5756 3003 5762
rect 3031 5756 3043 5762
rect 3077 5756 3089 5762
rect 3176 5756 3188 5762
rect 3226 5756 3238 5762
rect 3291 5756 3303 5762
rect 2731 5714 2742 5716
rect 2695 5708 2742 5714
rect 2367 5619 2374 5633
rect 2257 5592 2281 5598
rect 2269 5584 2281 5592
rect 1997 5538 2009 5544
rect 2078 5538 2090 5544
rect 2128 5538 2140 5544
rect 2157 5538 2169 5544
rect 2197 5538 2209 5544
rect 2366 5576 2374 5619
rect 2535 5598 2543 5647
rect 2519 5592 2543 5598
rect 2577 5603 2583 5673
rect 2595 5653 2602 5708
rect 2567 5597 2583 5603
rect 2596 5611 2604 5639
rect 2677 5627 2683 5673
rect 2695 5653 2702 5708
rect 2797 5661 2805 5716
rect 2975 5714 2983 5716
rect 3011 5714 3022 5716
rect 2975 5708 3022 5714
rect 2696 5611 2704 5639
rect 2596 5602 2626 5611
rect 2596 5600 2614 5602
rect 2519 5584 2531 5592
rect 2366 5570 2438 5576
rect 2391 5564 2398 5570
rect 2431 5564 2438 5570
rect 2696 5602 2726 5611
rect 2696 5600 2714 5602
rect 2797 5598 2805 5647
rect 2893 5641 2901 5676
rect 2975 5653 2982 5708
rect 3057 5682 3069 5684
rect 3057 5676 3097 5682
rect 3317 5756 3329 5762
rect 3357 5756 3369 5762
rect 3451 5756 3463 5762
rect 3491 5756 3503 5762
rect 3551 5756 3563 5762
rect 3591 5756 3603 5762
rect 3651 5756 3663 5762
rect 3118 5641 3126 5676
rect 3199 5641 3207 5676
rect 2899 5605 2907 5627
rect 2976 5611 2984 5639
rect 2900 5598 2925 5605
rect 2976 5602 3006 5611
rect 2976 5600 2994 5602
rect 2797 5592 2821 5598
rect 2809 5584 2821 5592
rect 2239 5538 2251 5544
rect 2411 5538 2423 5544
rect 2451 5538 2465 5544
rect 2549 5538 2561 5544
rect 2650 5538 2662 5544
rect 2750 5538 2762 5544
rect 2857 5584 2909 5587
rect 2869 5578 2897 5584
rect 2917 5584 2925 5598
rect 3118 5584 3126 5627
rect 3193 5605 3201 5627
rect 3276 5633 3284 5716
rect 3338 5714 3349 5716
rect 3377 5714 3385 5716
rect 3338 5708 3385 5714
rect 3378 5653 3385 5708
rect 3435 5714 3443 5716
rect 3471 5714 3482 5716
rect 3435 5708 3482 5714
rect 3535 5714 3543 5716
rect 3696 5756 3708 5762
rect 3746 5756 3758 5762
rect 3831 5756 3843 5762
rect 3571 5714 3582 5716
rect 3535 5708 3582 5714
rect 3435 5653 3442 5708
rect 3535 5653 3542 5708
rect 3175 5598 3200 5605
rect 3175 5584 3183 5598
rect 2779 5538 2791 5544
rect 2877 5538 2889 5544
rect 3030 5538 3042 5544
rect 3100 5573 3126 5584
rect 3191 5584 3243 5587
rect 3203 5578 3231 5584
rect 3276 5564 3284 5619
rect 3376 5611 3384 5639
rect 3060 5538 3072 5544
rect 3110 5538 3122 5544
rect 3211 5538 3223 5544
rect 3291 5538 3303 5544
rect 3354 5602 3384 5611
rect 3366 5600 3384 5602
rect 3436 5611 3444 5639
rect 3487 5617 3513 5623
rect 3536 5611 3544 5639
rect 3636 5633 3644 5716
rect 3862 5756 3874 5762
rect 3912 5756 3924 5762
rect 3991 5756 4003 5762
rect 4091 5756 4103 5762
rect 4156 5756 4168 5762
rect 4206 5756 4218 5762
rect 4271 5756 4283 5762
rect 4311 5756 4323 5762
rect 3719 5641 3727 5676
rect 3803 5669 3820 5676
rect 3436 5602 3466 5611
rect 3436 5600 3454 5602
rect 3536 5602 3566 5611
rect 3536 5600 3554 5602
rect 3636 5564 3644 5619
rect 3713 5605 3721 5627
rect 3813 5621 3820 5669
rect 3893 5641 3901 5676
rect 3976 5633 3984 5716
rect 4043 5750 4071 5756
rect 4083 5678 4111 5684
rect 4137 5697 4153 5703
rect 4052 5670 4064 5676
rect 4052 5664 4079 5670
rect 4073 5641 4079 5664
rect 3695 5598 3720 5605
rect 3695 5584 3703 5598
rect 3711 5584 3763 5587
rect 3723 5578 3751 5584
rect 3813 5564 3820 5607
rect 3899 5605 3907 5627
rect 3900 5598 3925 5605
rect 3857 5584 3909 5587
rect 3869 5578 3897 5584
rect 3917 5584 3925 5598
rect 3976 5564 3984 5619
rect 4080 5584 4087 5627
rect 4137 5623 4143 5697
rect 4255 5714 4263 5716
rect 4337 5756 4349 5762
rect 4416 5756 4428 5762
rect 4466 5756 4478 5762
rect 4527 5756 4539 5762
rect 4571 5756 4583 5762
rect 4291 5714 4302 5716
rect 4255 5708 4302 5714
rect 4179 5641 4187 5676
rect 4255 5653 4262 5708
rect 4137 5617 4153 5623
rect 4173 5605 4181 5627
rect 4256 5611 4264 5639
rect 4356 5633 4364 5716
rect 4597 5756 4609 5762
rect 4637 5756 4649 5762
rect 4696 5756 4708 5762
rect 4746 5756 4758 5762
rect 4439 5641 4447 5676
rect 4511 5641 4519 5676
rect 4155 5598 4180 5605
rect 4256 5602 4286 5611
rect 4256 5600 4274 5602
rect 4155 5584 4163 5598
rect 3318 5538 3330 5544
rect 3490 5538 3502 5544
rect 3590 5538 3602 5544
rect 3651 5538 3663 5544
rect 3731 5538 3743 5544
rect 3791 5538 3803 5544
rect 3831 5538 3843 5544
rect 3877 5538 3889 5544
rect 3991 5538 4003 5544
rect 4171 5584 4223 5587
rect 4183 5578 4211 5584
rect 4356 5564 4364 5619
rect 4433 5605 4441 5627
rect 4511 5627 4513 5641
rect 4415 5598 4440 5605
rect 4415 5584 4423 5598
rect 4052 5538 4064 5544
rect 4108 5538 4120 5544
rect 4191 5538 4203 5544
rect 4310 5538 4322 5544
rect 4431 5584 4483 5587
rect 4443 5578 4471 5584
rect 4511 5584 4519 5627
rect 4554 5602 4562 5716
rect 4617 5661 4625 5716
rect 4782 5756 4794 5762
rect 4832 5756 4844 5762
rect 4911 5756 4923 5762
rect 4951 5756 4963 5762
rect 4997 5756 5009 5762
rect 5082 5756 5094 5762
rect 5132 5756 5144 5762
rect 4895 5714 4903 5716
rect 4931 5714 4942 5716
rect 4545 5594 4583 5602
rect 4571 5584 4583 5594
rect 4617 5598 4625 5647
rect 4719 5641 4727 5676
rect 4813 5641 4821 5676
rect 4713 5605 4721 5627
rect 4819 5605 4827 5627
rect 4857 5623 4863 5713
rect 4895 5708 4942 5714
rect 4895 5653 4902 5708
rect 4977 5682 4989 5684
rect 4977 5676 5017 5682
rect 5177 5756 5189 5762
rect 5217 5756 5229 5762
rect 5277 5756 5289 5762
rect 5317 5756 5329 5762
rect 5198 5714 5209 5716
rect 5357 5756 5369 5762
rect 5397 5756 5409 5762
rect 5477 5756 5489 5762
rect 5557 5756 5569 5762
rect 5597 5756 5609 5762
rect 5237 5714 5245 5716
rect 5198 5708 5245 5714
rect 5157 5697 5173 5703
rect 5038 5641 5046 5676
rect 4847 5617 4883 5623
rect 4695 5598 4720 5605
rect 4820 5598 4845 5605
rect 4617 5592 4641 5598
rect 4629 5584 4641 5592
rect 4695 5584 4703 5598
rect 4511 5574 4521 5584
rect 4711 5584 4763 5587
rect 4723 5578 4751 5584
rect 4777 5584 4829 5587
rect 4789 5578 4817 5584
rect 4837 5584 4845 5598
rect 4877 5583 4883 5617
rect 4896 5611 4904 5639
rect 4896 5602 4926 5611
rect 4896 5600 4914 5602
rect 4877 5577 4893 5583
rect 5038 5584 5046 5627
rect 5057 5587 5063 5653
rect 5113 5641 5121 5676
rect 5119 5605 5127 5627
rect 5157 5623 5163 5697
rect 5238 5653 5245 5708
rect 5157 5617 5193 5623
rect 5236 5611 5244 5639
rect 5120 5598 5145 5605
rect 4337 5538 4349 5544
rect 4451 5538 4463 5544
rect 4541 5538 4553 5544
rect 4599 5538 4611 5544
rect 4731 5538 4743 5544
rect 4797 5538 4809 5544
rect 4950 5538 4962 5544
rect 5020 5573 5046 5584
rect 5077 5584 5129 5587
rect 5089 5578 5117 5584
rect 5137 5584 5145 5598
rect 5214 5602 5244 5611
rect 5226 5600 5244 5602
rect 5257 5583 5263 5673
rect 5297 5661 5305 5716
rect 5378 5714 5389 5716
rect 5417 5714 5425 5716
rect 5378 5708 5425 5714
rect 5297 5598 5305 5647
rect 5418 5653 5425 5708
rect 5457 5682 5469 5684
rect 5457 5676 5497 5682
rect 5651 5756 5663 5762
rect 5691 5756 5703 5762
rect 5737 5756 5749 5762
rect 5856 5756 5868 5762
rect 5906 5756 5918 5762
rect 5518 5641 5526 5676
rect 5577 5661 5585 5716
rect 5637 5677 5653 5683
rect 5416 5611 5424 5639
rect 5297 5592 5321 5598
rect 5309 5584 5321 5592
rect 5247 5577 5263 5583
rect 5394 5602 5424 5611
rect 5406 5600 5424 5602
rect 5518 5584 5526 5627
rect 5577 5598 5585 5647
rect 5577 5592 5601 5598
rect 5589 5584 5601 5592
rect 5500 5573 5526 5584
rect 4980 5538 4992 5544
rect 5030 5538 5042 5544
rect 5097 5538 5109 5544
rect 5178 5538 5190 5544
rect 5279 5538 5291 5544
rect 5358 5538 5370 5544
rect 5460 5538 5472 5544
rect 5510 5538 5522 5544
rect 5637 5567 5643 5677
rect 5675 5661 5683 5716
rect 5729 5678 5757 5684
rect 5769 5750 5797 5756
rect 5937 5756 5949 5762
rect 6017 5756 6029 5762
rect 6117 5756 6129 5762
rect 6157 5756 6169 5762
rect 6251 5756 6263 5762
rect 6297 5756 6309 5762
rect 6377 5756 6389 5762
rect 6417 5756 6429 5762
rect 6477 5756 6489 5762
rect 6517 5756 6529 5762
rect 6577 5756 6589 5762
rect 6617 5756 6629 5762
rect 5776 5670 5788 5676
rect 5761 5664 5788 5670
rect 5675 5598 5683 5647
rect 5761 5641 5767 5664
rect 5879 5641 5887 5676
rect 5659 5592 5683 5598
rect 5659 5584 5671 5592
rect 5753 5584 5760 5627
rect 5873 5605 5881 5627
rect 5956 5633 5964 5716
rect 6009 5678 6037 5684
rect 6049 5750 6077 5756
rect 6138 5714 6149 5716
rect 6177 5714 6185 5716
rect 6138 5708 6185 5714
rect 6056 5670 6068 5676
rect 6041 5664 6068 5670
rect 6041 5641 6047 5664
rect 6178 5653 6185 5708
rect 5855 5598 5880 5605
rect 5855 5584 5863 5598
rect 5559 5538 5571 5544
rect 5689 5538 5701 5544
rect 5871 5584 5923 5587
rect 5883 5578 5911 5584
rect 5956 5564 5964 5619
rect 6033 5584 6040 5627
rect 6176 5611 6184 5639
rect 6236 5633 6244 5716
rect 6277 5682 6289 5684
rect 6277 5676 6317 5682
rect 6398 5714 6409 5716
rect 6437 5714 6445 5716
rect 6398 5708 6445 5714
rect 6498 5714 6509 5716
rect 6537 5714 6545 5716
rect 6498 5708 6545 5714
rect 6598 5714 6609 5716
rect 6637 5714 6645 5716
rect 6598 5708 6645 5714
rect 6338 5641 6346 5676
rect 5720 5538 5732 5544
rect 5776 5538 5788 5544
rect 5891 5538 5903 5544
rect 5937 5538 5949 5544
rect 6000 5538 6012 5544
rect 6056 5538 6068 5544
rect 6154 5602 6184 5611
rect 6166 5600 6184 5602
rect 6236 5564 6244 5619
rect 6338 5584 6346 5627
rect 6357 5607 6363 5653
rect 6438 5653 6445 5708
rect 6436 5611 6444 5639
rect 6457 5627 6463 5693
rect 6538 5653 6545 5708
rect 6638 5653 6645 5708
rect 6536 5611 6544 5639
rect 6636 5611 6644 5639
rect 6118 5538 6130 5544
rect 6251 5538 6263 5544
rect 6320 5573 6346 5584
rect 6280 5538 6292 5544
rect 6330 5538 6342 5544
rect 6414 5602 6444 5611
rect 6426 5600 6444 5602
rect 6514 5602 6544 5611
rect 6526 5600 6544 5602
rect 6614 5602 6644 5611
rect 6626 5600 6644 5602
rect 6378 5538 6390 5544
rect 6478 5538 6490 5544
rect 6578 5538 6590 5544
rect 6742 5538 6802 6002
rect 4 5536 6802 5538
rect 6736 5524 6802 5536
rect 4 5522 6802 5524
rect 39 5516 51 5522
rect 97 5516 109 5522
rect 145 5516 157 5522
rect 207 5516 219 5522
rect 259 5516 271 5522
rect 358 5516 370 5522
rect 408 5516 420 5522
rect 489 5516 501 5522
rect 561 5516 573 5522
rect 617 5516 629 5522
rect 657 5516 669 5522
rect 187 5496 200 5502
rect 71 5490 78 5496
rect 67 5482 78 5490
rect 128 5484 135 5496
rect 193 5490 200 5496
rect 17 5461 25 5476
rect 128 5477 149 5484
rect 107 5466 113 5468
rect 174 5466 181 5472
rect 17 5447 33 5461
rect 107 5460 181 5466
rect 17 5384 25 5447
rect 33 5433 47 5447
rect 39 5388 53 5396
rect 107 5388 113 5460
rect 174 5452 181 5460
rect 186 5444 220 5452
rect 214 5439 220 5444
rect 167 5426 194 5433
rect 73 5382 113 5388
rect 121 5388 165 5394
rect 73 5364 79 5382
rect 121 5374 127 5388
rect 233 5392 239 5476
rect 289 5468 301 5476
rect 277 5462 301 5468
rect 354 5476 380 5487
rect 531 5476 541 5486
rect 697 5516 709 5522
rect 737 5516 749 5522
rect 779 5516 791 5522
rect 859 5516 871 5522
rect 937 5516 949 5522
rect 1000 5516 1012 5522
rect 1050 5516 1062 5522
rect 277 5413 285 5462
rect 354 5433 362 5476
rect 459 5468 471 5476
rect 459 5462 483 5468
rect 177 5384 239 5392
rect 97 5368 127 5374
rect 145 5370 183 5378
rect 175 5364 183 5370
rect 67 5324 79 5358
rect 125 5350 147 5362
rect 175 5350 193 5364
rect 121 5344 133 5350
rect 175 5344 183 5350
rect 277 5344 285 5399
rect 354 5384 362 5419
rect 475 5413 483 5462
rect 531 5433 539 5476
rect 591 5466 603 5476
rect 565 5458 603 5466
rect 531 5419 533 5433
rect 383 5378 423 5384
rect 411 5376 423 5378
rect 475 5344 483 5399
rect 531 5384 539 5419
rect 574 5344 582 5458
rect 640 5453 647 5496
rect 720 5453 727 5496
rect 809 5468 821 5476
rect 889 5468 901 5476
rect 640 5391 647 5439
rect 720 5391 727 5439
rect 797 5462 821 5468
rect 877 5462 901 5468
rect 797 5413 805 5462
rect 877 5413 885 5462
rect 917 5403 923 5473
rect 956 5441 964 5496
rect 1132 5516 1144 5522
rect 1188 5516 1200 5522
rect 1239 5516 1251 5522
rect 1297 5516 1309 5522
rect 1345 5516 1357 5522
rect 1407 5516 1419 5522
rect 1530 5516 1542 5522
rect 1630 5516 1642 5522
rect 1691 5516 1703 5522
rect 1771 5516 1783 5522
rect 1861 5516 1873 5522
rect 1969 5516 1981 5522
rect 2051 5516 2063 5522
rect 2099 5516 2111 5522
rect 2211 5516 2223 5522
rect 2291 5516 2303 5522
rect 2337 5516 2349 5522
rect 2377 5516 2389 5522
rect 2451 5516 2463 5522
rect 1040 5476 1066 5487
rect 1387 5496 1400 5502
rect 1271 5490 1278 5496
rect 1267 5482 1278 5490
rect 1328 5484 1335 5496
rect 1393 5490 1400 5496
rect 1058 5433 1066 5476
rect 640 5384 657 5391
rect 720 5384 737 5391
rect 37 5298 49 5304
rect 95 5298 107 5304
rect 141 5298 153 5304
rect 207 5298 219 5304
rect 257 5298 269 5304
rect 297 5298 309 5304
rect 391 5298 403 5304
rect 451 5298 463 5304
rect 491 5298 503 5304
rect 547 5298 559 5304
rect 591 5298 603 5304
rect 797 5344 805 5399
rect 877 5344 885 5399
rect 917 5397 933 5403
rect 956 5344 964 5427
rect 1160 5433 1167 5476
rect 1217 5461 1225 5476
rect 1328 5477 1349 5484
rect 1307 5466 1313 5468
rect 1374 5466 1381 5472
rect 1217 5447 1233 5461
rect 1307 5460 1381 5466
rect 987 5397 1013 5403
rect 1058 5384 1066 5419
rect 1153 5396 1159 5419
rect 1132 5390 1159 5396
rect 1132 5384 1144 5390
rect 1217 5384 1225 5447
rect 1233 5433 1247 5447
rect 1239 5388 1253 5396
rect 997 5378 1037 5384
rect 997 5376 1009 5378
rect 617 5298 629 5304
rect 697 5298 709 5304
rect 777 5298 789 5304
rect 817 5298 829 5304
rect 857 5298 869 5304
rect 897 5298 909 5304
rect 1123 5304 1151 5310
rect 1163 5376 1191 5382
rect 1307 5388 1313 5460
rect 1374 5452 1381 5460
rect 1386 5444 1420 5452
rect 1414 5439 1420 5444
rect 1367 5426 1394 5433
rect 1273 5382 1313 5388
rect 1321 5388 1365 5394
rect 1273 5364 1279 5382
rect 1321 5374 1327 5388
rect 1433 5392 1439 5476
rect 1476 5458 1494 5460
rect 1476 5449 1506 5458
rect 1576 5458 1594 5460
rect 1576 5449 1606 5458
rect 1476 5421 1484 5449
rect 1576 5421 1584 5449
rect 1627 5437 1653 5443
rect 1676 5441 1684 5496
rect 1735 5462 1743 5476
rect 1763 5476 1791 5482
rect 1751 5473 1803 5476
rect 1831 5476 1841 5486
rect 1735 5455 1760 5462
rect 1717 5437 1733 5443
rect 1377 5384 1439 5392
rect 1297 5368 1327 5374
rect 1345 5370 1383 5378
rect 1375 5364 1383 5370
rect 1267 5324 1279 5358
rect 1325 5350 1347 5362
rect 1375 5350 1393 5364
rect 1321 5344 1333 5350
rect 1375 5344 1383 5350
rect 1475 5352 1482 5407
rect 1575 5352 1582 5407
rect 1475 5346 1522 5352
rect 1475 5344 1483 5346
rect 1511 5344 1522 5346
rect 1575 5346 1622 5352
rect 1575 5344 1583 5346
rect 1611 5344 1622 5346
rect 1676 5344 1684 5427
rect 1717 5403 1723 5437
rect 1753 5433 1761 5455
rect 1831 5433 1839 5476
rect 1891 5466 1903 5476
rect 1865 5458 1903 5466
rect 1939 5468 1951 5476
rect 1939 5462 1963 5468
rect 1831 5419 1833 5433
rect 1707 5397 1723 5403
rect 1759 5384 1767 5419
rect 1831 5384 1839 5419
rect 937 5298 949 5304
rect 1017 5298 1029 5304
rect 1171 5298 1183 5304
rect 1237 5298 1249 5304
rect 1295 5298 1307 5304
rect 1341 5298 1353 5304
rect 1407 5298 1419 5304
rect 1491 5298 1503 5304
rect 1531 5298 1543 5304
rect 1591 5298 1603 5304
rect 1631 5298 1643 5304
rect 1691 5298 1703 5304
rect -62 5296 1713 5298
rect 1874 5344 1882 5458
rect 1955 5413 1963 5462
rect 2015 5462 2023 5476
rect 2043 5476 2071 5482
rect 2031 5473 2083 5476
rect 2129 5468 2141 5476
rect 2117 5462 2141 5468
rect 2015 5455 2040 5462
rect 2033 5433 2041 5455
rect 1955 5344 1963 5399
rect 2039 5384 2047 5419
rect 2117 5413 2125 5462
rect 2196 5441 2204 5496
rect 2255 5462 2263 5476
rect 2283 5476 2311 5482
rect 2498 5516 2510 5522
rect 2548 5516 2560 5522
rect 2597 5516 2609 5522
rect 2679 5516 2691 5522
rect 2830 5516 2842 5522
rect 2909 5516 2921 5522
rect 2271 5473 2323 5476
rect 2255 5455 2280 5462
rect 2273 5433 2281 5455
rect 2360 5453 2367 5496
rect 1736 5298 1748 5304
rect 1786 5298 1798 5304
rect 1847 5298 1859 5304
rect 1891 5298 1903 5304
rect 1931 5298 1943 5304
rect 1971 5298 1983 5304
rect 2117 5344 2125 5399
rect 2196 5344 2204 5427
rect 2436 5441 2444 5496
rect 2494 5476 2520 5487
rect 2589 5476 2617 5482
rect 2279 5384 2287 5419
rect 2360 5391 2367 5439
rect 2494 5433 2502 5476
rect 2577 5473 2629 5476
rect 2637 5462 2645 5476
rect 2709 5468 2721 5476
rect 2620 5455 2645 5462
rect 2697 5462 2721 5468
rect 2360 5384 2377 5391
rect 2016 5298 2028 5304
rect 2066 5298 2078 5304
rect 2097 5298 2109 5304
rect 2137 5298 2149 5304
rect 2211 5298 2223 5304
rect 2256 5298 2268 5304
rect 2306 5298 2318 5304
rect 2436 5344 2444 5427
rect 2619 5433 2627 5455
rect 2494 5384 2502 5419
rect 2613 5384 2621 5419
rect 2697 5413 2705 5462
rect 2776 5458 2794 5460
rect 2776 5449 2806 5458
rect 2951 5516 2963 5522
rect 2991 5516 3003 5522
rect 3037 5516 3049 5522
rect 3169 5516 3181 5522
rect 3217 5516 3229 5522
rect 3341 5516 3353 5522
rect 3397 5516 3409 5522
rect 3437 5516 3449 5522
rect 2879 5468 2891 5476
rect 2879 5462 2903 5468
rect 2776 5421 2784 5449
rect 2523 5378 2563 5384
rect 2551 5376 2563 5378
rect 2697 5344 2705 5399
rect 2775 5352 2782 5407
rect 2895 5413 2903 5462
rect 2973 5453 2980 5496
rect 3029 5476 3057 5482
rect 3017 5473 3069 5476
rect 3209 5476 3237 5482
rect 3077 5462 3085 5476
rect 3139 5468 3151 5476
rect 3197 5473 3249 5476
rect 3311 5476 3321 5486
rect 3477 5516 3485 5522
rect 3517 5516 3529 5522
rect 3597 5516 3609 5522
rect 3691 5516 3703 5522
rect 3731 5516 3743 5522
rect 3777 5516 3789 5522
rect 3891 5516 3903 5522
rect 3931 5516 3943 5522
rect 3977 5516 3989 5522
rect 4130 5516 4142 5522
rect 4209 5516 4221 5522
rect 3139 5462 3163 5468
rect 3257 5462 3265 5476
rect 3060 5455 3085 5462
rect 2775 5346 2822 5352
rect 2775 5344 2783 5346
rect 2337 5298 2349 5304
rect 2451 5298 2463 5304
rect 2531 5298 2543 5304
rect 2582 5298 2594 5304
rect 2632 5298 2644 5304
rect 2811 5344 2822 5346
rect 2895 5344 2903 5399
rect 2973 5391 2980 5439
rect 3059 5433 3067 5455
rect 2963 5384 2980 5391
rect 3053 5384 3061 5419
rect 3155 5413 3163 5462
rect 3240 5455 3265 5462
rect 3239 5433 3247 5455
rect 3311 5433 3319 5476
rect 3371 5466 3383 5476
rect 3345 5458 3383 5466
rect 3311 5419 3313 5433
rect 2677 5298 2689 5304
rect 2717 5298 2729 5304
rect 2791 5298 2803 5304
rect 2831 5298 2843 5304
rect 2871 5298 2883 5304
rect 2911 5298 2923 5304
rect 1727 5296 2933 5298
rect 2991 5298 3003 5304
rect 3155 5344 3163 5399
rect 3233 5384 3241 5419
rect 3311 5384 3319 5419
rect 3022 5298 3034 5304
rect 3072 5298 3084 5304
rect 3131 5298 3143 5304
rect 3171 5298 3183 5304
rect 3354 5344 3362 5458
rect 3420 5453 3427 5496
rect 3503 5468 3509 5496
rect 3589 5476 3617 5482
rect 3503 5462 3513 5468
rect 3420 5391 3427 5439
rect 3518 5401 3524 5456
rect 3540 5441 3547 5476
rect 3577 5473 3629 5476
rect 3637 5462 3645 5476
rect 3620 5455 3645 5462
rect 3477 5392 3513 5400
rect 3420 5384 3437 5391
rect 3202 5298 3214 5304
rect 3252 5298 3264 5304
rect 3327 5298 3339 5304
rect 3371 5298 3383 5304
rect 3477 5384 3485 5392
rect 3534 5383 3543 5427
rect 3619 5433 3627 5455
rect 3713 5453 3720 5496
rect 3769 5476 3797 5480
rect 3809 5510 3837 5516
rect 3757 5474 3809 5476
rect 3819 5466 3825 5476
rect 3796 5459 3825 5466
rect 3613 5384 3621 5419
rect 3713 5391 3720 5439
rect 3796 5433 3804 5459
rect 3913 5453 3920 5496
rect 3969 5476 3997 5482
rect 3957 5473 4009 5476
rect 4017 5462 4025 5476
rect 4000 5455 4025 5462
rect 4076 5458 4094 5460
rect 3703 5384 3720 5391
rect 3797 5384 3805 5419
rect 3913 5391 3920 5439
rect 3999 5433 4007 5455
rect 4076 5449 4106 5458
rect 4237 5516 4249 5522
rect 4351 5516 4363 5522
rect 4449 5516 4461 5522
rect 4179 5468 4191 5476
rect 4179 5462 4203 5468
rect 4076 5421 4084 5449
rect 3903 5384 3920 5391
rect 3993 5384 4001 5419
rect 3539 5374 3543 5383
rect 3397 5298 3409 5304
rect 3507 5298 3519 5304
rect 3582 5298 3594 5304
rect 3632 5298 3644 5304
rect 3731 5298 3743 5304
rect 3757 5298 3769 5304
rect 3827 5298 3839 5304
rect 3931 5298 3943 5304
rect 4075 5352 4082 5407
rect 4195 5413 4203 5462
rect 4256 5441 4264 5496
rect 4315 5462 4323 5476
rect 4343 5476 4371 5482
rect 4331 5473 4383 5476
rect 4479 5516 4491 5522
rect 4611 5516 4623 5522
rect 4711 5516 4723 5522
rect 4801 5516 4813 5522
rect 4911 5516 4923 5522
rect 5009 5516 5021 5522
rect 5081 5516 5093 5522
rect 5139 5516 5151 5522
rect 5237 5516 5249 5522
rect 5361 5516 5373 5522
rect 5437 5516 5449 5522
rect 5519 5516 5531 5522
rect 5598 5516 5610 5522
rect 5741 5516 5753 5522
rect 5832 5516 5844 5522
rect 5888 5516 5900 5522
rect 4419 5468 4431 5476
rect 4509 5468 4521 5476
rect 4419 5462 4443 5468
rect 4315 5455 4340 5462
rect 4333 5433 4341 5455
rect 4075 5346 4122 5352
rect 4075 5344 4083 5346
rect 4111 5344 4122 5346
rect 4195 5344 4203 5399
rect 4256 5344 4264 5427
rect 4339 5384 4347 5419
rect 4435 5413 4443 5462
rect 4497 5462 4521 5468
rect 4575 5462 4583 5476
rect 4603 5476 4631 5482
rect 4591 5473 4643 5476
rect 4675 5462 4683 5476
rect 4703 5476 4731 5482
rect 4691 5473 4743 5476
rect 4771 5476 4781 5486
rect 4497 5413 4505 5462
rect 4575 5455 4600 5462
rect 4675 5455 4700 5462
rect 4557 5437 4573 5443
rect 3962 5298 3974 5304
rect 4012 5298 4024 5304
rect 4091 5298 4103 5304
rect 4131 5298 4143 5304
rect 4171 5298 4183 5304
rect 4211 5298 4223 5304
rect 4435 5344 4443 5399
rect 4497 5344 4505 5399
rect 4557 5363 4563 5437
rect 4593 5433 4601 5455
rect 4693 5433 4701 5455
rect 4599 5384 4607 5419
rect 4657 5387 4663 5433
rect 4771 5433 4779 5476
rect 4831 5466 4843 5476
rect 4805 5458 4843 5466
rect 4875 5462 4883 5476
rect 4903 5476 4931 5482
rect 4891 5473 4943 5476
rect 5051 5476 5061 5486
rect 4979 5468 4991 5476
rect 4979 5462 5003 5468
rect 4771 5419 4773 5433
rect 4557 5357 4573 5363
rect 4237 5298 4249 5304
rect 4316 5298 4328 5304
rect 4366 5298 4378 5304
rect 4411 5298 4423 5304
rect 4451 5298 4463 5304
rect 4477 5298 4489 5304
rect 4517 5298 4529 5304
rect 4699 5384 4707 5419
rect 4771 5384 4779 5419
rect 4576 5298 4588 5304
rect 4626 5298 4638 5304
rect 4814 5344 4822 5458
rect 4875 5455 4900 5462
rect 4893 5433 4901 5455
rect 4899 5384 4907 5419
rect 4995 5413 5003 5462
rect 5051 5433 5059 5476
rect 5111 5466 5123 5476
rect 5169 5468 5181 5476
rect 5229 5476 5257 5482
rect 5217 5473 5269 5476
rect 5331 5476 5341 5486
rect 5085 5458 5123 5466
rect 5157 5462 5181 5468
rect 5277 5462 5285 5476
rect 5051 5419 5053 5433
rect 4676 5298 4688 5304
rect 4726 5298 4738 5304
rect 4787 5298 4799 5304
rect 4831 5298 4843 5304
rect 4995 5344 5003 5399
rect 5051 5384 5059 5419
rect 4876 5298 4888 5304
rect 4926 5298 4938 5304
rect 5094 5344 5102 5458
rect 5157 5413 5165 5462
rect 5260 5455 5285 5462
rect 5259 5433 5267 5455
rect 5331 5433 5339 5476
rect 5391 5466 5403 5476
rect 5429 5476 5457 5482
rect 5417 5473 5469 5476
rect 5365 5458 5403 5466
rect 5477 5462 5485 5476
rect 5549 5468 5561 5476
rect 5331 5419 5333 5433
rect 5157 5344 5165 5399
rect 5253 5384 5261 5419
rect 5331 5384 5339 5419
rect 4971 5298 4983 5304
rect 5011 5298 5023 5304
rect 5067 5298 5079 5304
rect 5111 5298 5123 5304
rect 5137 5298 5149 5304
rect 5177 5298 5189 5304
rect 5374 5344 5382 5458
rect 5460 5455 5485 5462
rect 5537 5462 5561 5468
rect 5459 5433 5467 5455
rect 5487 5437 5503 5443
rect 5453 5384 5461 5419
rect 5222 5298 5234 5304
rect 5272 5298 5284 5304
rect 5347 5298 5359 5304
rect 5391 5298 5403 5304
rect 5497 5363 5503 5437
rect 5537 5413 5545 5462
rect 5711 5476 5721 5486
rect 5919 5516 5931 5522
rect 5998 5516 6010 5522
rect 6100 5516 6112 5522
rect 6150 5516 6162 5522
rect 6251 5516 6263 5522
rect 6317 5516 6329 5522
rect 6451 5516 6463 5522
rect 6570 5516 6582 5522
rect 5646 5458 5664 5460
rect 5634 5449 5664 5458
rect 5577 5437 5613 5443
rect 5487 5357 5503 5363
rect 5537 5344 5545 5399
rect 5577 5367 5583 5437
rect 5656 5421 5664 5449
rect 5711 5433 5719 5476
rect 5771 5466 5783 5476
rect 5745 5458 5783 5466
rect 5711 5419 5713 5433
rect 5658 5352 5665 5407
rect 5711 5384 5719 5419
rect 5618 5346 5665 5352
rect 5618 5344 5629 5346
rect 5422 5298 5434 5304
rect 5472 5298 5484 5304
rect 5517 5298 5529 5304
rect 5557 5298 5569 5304
rect 5657 5344 5665 5346
rect 5754 5344 5762 5458
rect 5860 5433 5867 5476
rect 5949 5468 5961 5476
rect 5937 5462 5961 5468
rect 5853 5396 5859 5419
rect 5937 5413 5945 5462
rect 6140 5476 6166 5487
rect 6046 5458 6064 5460
rect 6034 5449 6064 5458
rect 6056 5421 6064 5449
rect 6158 5433 6166 5476
rect 6215 5462 6223 5476
rect 6243 5476 6271 5482
rect 6231 5473 6283 5476
rect 6309 5476 6337 5482
rect 6297 5473 6349 5476
rect 6357 5462 6365 5476
rect 6215 5455 6240 5462
rect 6340 5455 6365 5462
rect 6415 5462 6423 5476
rect 6443 5476 6471 5482
rect 6431 5473 6483 5476
rect 6415 5455 6440 5462
rect 6516 5458 6534 5460
rect 6233 5433 6241 5455
rect 6339 5433 6347 5455
rect 6377 5437 6413 5443
rect 5832 5390 5859 5396
rect 5832 5384 5844 5390
rect 5823 5304 5851 5310
rect 5863 5376 5891 5382
rect 5937 5344 5945 5399
rect 6058 5352 6065 5407
rect 6158 5384 6166 5419
rect 6239 5384 6247 5419
rect 6333 5384 6341 5419
rect 6018 5346 6065 5352
rect 6018 5344 6029 5346
rect 5597 5298 5609 5304
rect 5637 5298 5649 5304
rect 5727 5298 5739 5304
rect 5771 5298 5783 5304
rect 5871 5298 5883 5304
rect 5917 5298 5929 5304
rect 5957 5298 5969 5304
rect 6057 5344 6065 5346
rect 6097 5378 6137 5384
rect 6097 5376 6109 5378
rect 5997 5298 6009 5304
rect 6037 5298 6049 5304
rect 6117 5298 6129 5304
rect 6216 5298 6228 5304
rect 6266 5298 6278 5304
rect 6377 5363 6383 5437
rect 6433 5433 6441 5455
rect 6516 5449 6546 5458
rect 6618 5516 6630 5522
rect 6668 5516 6680 5522
rect 6614 5476 6640 5487
rect 6516 5421 6524 5449
rect 6567 5437 6573 5443
rect 6614 5433 6622 5476
rect 6367 5357 6383 5363
rect 6397 5363 6403 5413
rect 6439 5384 6447 5419
rect 6397 5357 6413 5363
rect 6302 5298 6314 5304
rect 6352 5298 6364 5304
rect 6515 5352 6522 5407
rect 6614 5384 6622 5419
rect 6515 5346 6562 5352
rect 6515 5344 6523 5346
rect 6551 5344 6562 5346
rect 6643 5378 6683 5384
rect 6671 5376 6683 5378
rect 6416 5298 6428 5304
rect 6466 5298 6478 5304
rect 6531 5298 6543 5304
rect 6571 5298 6583 5304
rect 6651 5298 6663 5304
rect 2947 5296 6736 5298
rect -62 5284 4 5296
rect -62 5282 1013 5284
rect -62 4818 -2 5282
rect 49 5276 61 5282
rect 117 5276 129 5282
rect 175 5276 187 5282
rect 221 5276 233 5282
rect 287 5276 299 5282
rect 337 5276 349 5282
rect 377 5276 389 5282
rect 471 5276 483 5282
rect 531 5276 543 5282
rect 571 5276 583 5282
rect 621 5276 633 5282
rect 687 5276 699 5282
rect 733 5276 745 5282
rect 791 5276 803 5282
rect 837 5276 849 5282
rect 877 5276 889 5282
rect 31 5161 39 5196
rect 75 5190 83 5236
rect 57 5184 83 5190
rect 147 5222 159 5256
rect 201 5230 213 5236
rect 255 5230 263 5236
rect 205 5218 227 5230
rect 255 5216 273 5230
rect 153 5198 159 5216
rect 177 5206 207 5212
rect 255 5210 263 5216
rect 57 5178 60 5184
rect 31 5147 33 5161
rect 31 5104 39 5147
rect 53 5122 60 5178
rect 57 5116 60 5122
rect 97 5133 105 5196
rect 119 5184 133 5192
rect 153 5192 193 5198
rect 113 5133 127 5147
rect 97 5119 113 5133
rect 187 5120 193 5192
rect 201 5192 207 5206
rect 225 5202 263 5210
rect 201 5186 245 5192
rect 257 5188 319 5196
rect 247 5147 274 5154
rect 294 5136 300 5141
rect 266 5128 300 5136
rect 254 5120 261 5128
rect 57 5110 79 5116
rect 71 5084 79 5110
rect 97 5104 105 5119
rect 187 5114 261 5120
rect 187 5112 193 5114
rect 254 5108 261 5114
rect 147 5090 158 5098
rect 151 5084 158 5090
rect 208 5096 229 5103
rect 313 5104 319 5188
rect 357 5181 365 5236
rect 491 5202 503 5204
rect 463 5196 503 5202
rect 357 5118 365 5167
rect 434 5161 442 5196
rect 555 5181 563 5236
rect 657 5230 665 5236
rect 707 5230 719 5236
rect 647 5216 665 5230
rect 693 5218 715 5230
rect 761 5222 773 5256
rect 657 5210 665 5216
rect 657 5202 695 5210
rect 713 5206 743 5212
rect 601 5188 663 5196
rect 357 5112 381 5118
rect 369 5104 381 5112
rect 208 5084 215 5096
rect 273 5084 280 5090
rect 267 5078 280 5084
rect 434 5104 442 5147
rect 555 5118 563 5167
rect 539 5112 563 5118
rect 539 5104 551 5112
rect 601 5104 607 5188
rect 713 5192 719 5206
rect 761 5198 767 5216
rect 675 5186 719 5192
rect 727 5192 767 5198
rect 646 5147 673 5154
rect 620 5136 626 5141
rect 620 5128 654 5136
rect 659 5120 666 5128
rect 727 5120 733 5192
rect 936 5276 948 5282
rect 986 5276 998 5282
rect 787 5184 801 5192
rect 793 5133 807 5147
rect 815 5133 823 5196
rect 857 5181 865 5236
rect 1027 5282 3673 5284
rect 1036 5276 1048 5282
rect 1086 5276 1098 5282
rect 1147 5276 1159 5282
rect 1191 5276 1203 5282
rect 1237 5276 1249 5282
rect 1295 5276 1307 5282
rect 1341 5276 1353 5282
rect 1407 5276 1419 5282
rect 1471 5276 1483 5282
rect 1511 5276 1523 5282
rect 659 5114 733 5120
rect 807 5119 823 5133
rect 659 5108 666 5114
rect 727 5112 733 5114
rect 434 5093 460 5104
rect 691 5096 712 5103
rect 815 5104 823 5119
rect 857 5118 865 5167
rect 959 5161 967 5196
rect 1059 5161 1067 5196
rect 1131 5161 1139 5196
rect 953 5125 961 5147
rect 1053 5125 1061 5147
rect 1131 5147 1133 5161
rect 935 5118 960 5125
rect 1035 5118 1060 5125
rect 857 5112 881 5118
rect 869 5104 881 5112
rect 935 5104 943 5118
rect 640 5084 647 5090
rect 705 5084 712 5096
rect 762 5090 773 5098
rect 762 5084 769 5090
rect 640 5078 653 5084
rect 951 5104 1003 5107
rect 1035 5104 1043 5118
rect 963 5098 991 5104
rect 1051 5104 1103 5107
rect 1063 5098 1091 5104
rect 1131 5104 1139 5147
rect 1174 5122 1182 5236
rect 1267 5222 1279 5256
rect 1321 5230 1333 5236
rect 1375 5230 1383 5236
rect 1325 5218 1347 5230
rect 1375 5216 1393 5230
rect 1273 5198 1279 5216
rect 1297 5206 1327 5212
rect 1375 5210 1383 5216
rect 1217 5133 1225 5196
rect 1239 5184 1253 5192
rect 1273 5192 1313 5198
rect 1233 5133 1247 5147
rect 1165 5114 1203 5122
rect 1191 5104 1203 5114
rect 1131 5094 1141 5104
rect 1217 5119 1233 5133
rect 1307 5120 1313 5192
rect 1321 5192 1327 5206
rect 1345 5202 1383 5210
rect 1537 5276 1549 5282
rect 1577 5276 1589 5282
rect 1637 5276 1649 5282
rect 1695 5276 1707 5282
rect 1741 5276 1753 5282
rect 1807 5276 1819 5282
rect 1931 5276 1943 5282
rect 1977 5276 1989 5282
rect 2067 5276 2079 5282
rect 2111 5276 2123 5282
rect 1321 5186 1365 5192
rect 1377 5188 1439 5196
rect 1367 5147 1394 5154
rect 1414 5136 1420 5141
rect 1386 5128 1420 5136
rect 1374 5120 1381 5128
rect 1217 5104 1225 5119
rect 1307 5114 1381 5120
rect 1307 5112 1313 5114
rect 1374 5108 1381 5114
rect 1267 5090 1278 5098
rect 1271 5084 1278 5090
rect 1328 5096 1349 5103
rect 1433 5104 1439 5188
rect 1495 5181 1503 5236
rect 1557 5181 1565 5236
rect 1667 5222 1679 5256
rect 1721 5230 1733 5236
rect 1775 5230 1783 5236
rect 1725 5218 1747 5230
rect 1775 5216 1793 5230
rect 1673 5198 1679 5216
rect 1697 5206 1727 5212
rect 1775 5210 1783 5216
rect 1495 5118 1503 5167
rect 1328 5084 1335 5096
rect 1393 5084 1400 5090
rect 1387 5078 1400 5084
rect 1479 5112 1503 5118
rect 1557 5118 1565 5167
rect 1617 5133 1625 5196
rect 1639 5184 1653 5192
rect 1673 5192 1713 5198
rect 1633 5133 1647 5147
rect 1617 5119 1633 5133
rect 1707 5120 1713 5192
rect 1721 5192 1727 5206
rect 1745 5202 1783 5210
rect 1883 5270 1911 5276
rect 1923 5198 1951 5204
rect 1721 5186 1765 5192
rect 1777 5188 1839 5196
rect 1767 5147 1794 5154
rect 1814 5136 1820 5141
rect 1786 5128 1820 5136
rect 1774 5120 1781 5128
rect 1557 5112 1581 5118
rect 1479 5104 1491 5112
rect 1569 5104 1581 5112
rect 49 5058 61 5064
rect 119 5058 131 5064
rect 177 5058 189 5064
rect 225 5058 237 5064
rect 287 5058 299 5064
rect 339 5058 351 5064
rect 438 5058 450 5064
rect 488 5058 500 5064
rect 569 5058 581 5064
rect 621 5058 633 5064
rect 683 5058 695 5064
rect 731 5058 743 5064
rect 789 5058 801 5064
rect 839 5058 851 5064
rect 971 5058 983 5064
rect 1071 5058 1083 5064
rect 1161 5058 1173 5064
rect 1239 5058 1251 5064
rect 1297 5058 1309 5064
rect 1345 5058 1357 5064
rect 1407 5058 1419 5064
rect 1509 5058 1521 5064
rect 1617 5104 1625 5119
rect 1707 5114 1781 5120
rect 1707 5112 1713 5114
rect 1774 5108 1781 5114
rect 1667 5090 1678 5098
rect 1671 5084 1678 5090
rect 1728 5096 1749 5103
rect 1833 5104 1839 5188
rect 1892 5190 1904 5196
rect 1892 5184 1919 5190
rect 1913 5161 1919 5184
rect 1920 5104 1927 5147
rect 1996 5153 2004 5236
rect 2137 5276 2149 5282
rect 2177 5276 2189 5282
rect 2261 5276 2273 5282
rect 2331 5276 2343 5282
rect 2371 5276 2383 5282
rect 2431 5276 2443 5282
rect 2471 5276 2483 5282
rect 2551 5276 2563 5282
rect 2051 5161 2059 5196
rect 2051 5147 2053 5161
rect 1728 5084 1735 5096
rect 1793 5084 1800 5090
rect 1787 5078 1800 5084
rect 1996 5084 2004 5139
rect 2051 5104 2059 5147
rect 2094 5122 2102 5236
rect 2157 5181 2165 5236
rect 2237 5197 2241 5206
rect 2085 5114 2123 5122
rect 2111 5104 2123 5114
rect 2157 5118 2165 5167
rect 2237 5153 2246 5197
rect 2295 5188 2303 5196
rect 2267 5180 2303 5188
rect 2355 5181 2363 5236
rect 2415 5234 2423 5236
rect 2451 5234 2462 5236
rect 2415 5228 2462 5234
rect 2157 5112 2181 5118
rect 2169 5104 2181 5112
rect 2233 5104 2240 5139
rect 2256 5124 2262 5179
rect 2415 5173 2422 5228
rect 2577 5276 2589 5282
rect 2667 5276 2679 5282
rect 2711 5276 2723 5282
rect 2523 5189 2540 5196
rect 2355 5118 2363 5167
rect 2416 5131 2424 5159
rect 2533 5141 2540 5189
rect 2596 5153 2604 5236
rect 2737 5276 2749 5282
rect 2831 5276 2843 5282
rect 2871 5276 2883 5282
rect 2651 5161 2659 5196
rect 2416 5122 2446 5131
rect 2651 5147 2653 5161
rect 2416 5120 2434 5122
rect 2267 5112 2277 5118
rect 2051 5094 2061 5104
rect 1539 5058 1551 5064
rect 1639 5058 1651 5064
rect 1697 5058 1709 5064
rect 1745 5058 1757 5064
rect 1807 5058 1819 5064
rect 1892 5058 1904 5064
rect 1948 5058 1960 5064
rect 2271 5084 2277 5112
rect 2339 5112 2363 5118
rect 2339 5104 2351 5112
rect 2533 5084 2540 5127
rect 2596 5084 2604 5139
rect 2651 5104 2659 5147
rect 2694 5122 2702 5236
rect 2911 5276 2923 5282
rect 2951 5276 2963 5282
rect 3007 5276 3019 5282
rect 3107 5276 3119 5282
rect 3151 5276 3163 5282
rect 2760 5189 2777 5196
rect 2760 5141 2767 5189
rect 2855 5181 2863 5236
rect 2935 5181 2943 5236
rect 3039 5197 3043 5206
rect 2977 5188 2985 5196
rect 2685 5114 2723 5122
rect 2711 5104 2723 5114
rect 2651 5094 2661 5104
rect 1977 5058 1989 5064
rect 2081 5058 2093 5064
rect 2139 5058 2151 5064
rect 2251 5058 2263 5064
rect 2295 5058 2303 5064
rect 2369 5058 2381 5064
rect 2470 5058 2482 5064
rect 2511 5058 2523 5064
rect 2551 5058 2563 5064
rect 2760 5084 2767 5127
rect 2855 5118 2863 5167
rect 2977 5180 3013 5188
rect 2935 5118 2943 5167
rect 3018 5124 3024 5179
rect 3034 5153 3043 5197
rect 3177 5276 3189 5282
rect 3217 5276 3229 5282
rect 3291 5276 3303 5282
rect 3331 5276 3343 5282
rect 3391 5276 3403 5282
rect 3471 5276 3483 5282
rect 3571 5276 3583 5282
rect 3091 5161 3099 5196
rect 2839 5112 2863 5118
rect 2919 5112 2943 5118
rect 3003 5112 3013 5118
rect 2839 5104 2851 5112
rect 2919 5104 2931 5112
rect 3003 5084 3009 5112
rect 3040 5104 3047 5139
rect 3091 5147 3093 5161
rect 3091 5104 3099 5147
rect 3134 5122 3142 5236
rect 3197 5181 3205 5236
rect 3275 5234 3283 5236
rect 3311 5234 3322 5236
rect 3275 5228 3322 5234
rect 3275 5173 3282 5228
rect 3125 5114 3163 5122
rect 3151 5104 3163 5114
rect 3197 5118 3205 5167
rect 3276 5131 3284 5159
rect 3376 5153 3384 5236
rect 3491 5202 3503 5204
rect 3463 5196 3503 5202
rect 3602 5276 3614 5282
rect 3652 5276 3664 5282
rect 3687 5282 4113 5284
rect 3716 5276 3728 5282
rect 3766 5276 3778 5282
rect 3667 5217 3683 5223
rect 3434 5161 3442 5196
rect 3543 5189 3560 5196
rect 3276 5122 3306 5131
rect 3276 5120 3294 5122
rect 3197 5112 3221 5118
rect 3209 5104 3221 5112
rect 2577 5058 2589 5064
rect 2681 5058 2693 5064
rect 2737 5058 2749 5064
rect 2777 5058 2789 5064
rect 2869 5058 2881 5064
rect 2949 5058 2961 5064
rect 3091 5094 3101 5104
rect 3376 5084 3384 5139
rect 3434 5104 3442 5147
rect 3553 5141 3560 5189
rect 3633 5161 3641 5196
rect 3434 5093 3460 5104
rect 2977 5058 2985 5064
rect 3017 5058 3029 5064
rect 3121 5058 3133 5064
rect 3179 5058 3191 5064
rect 3330 5058 3342 5064
rect 3391 5058 3403 5064
rect 3553 5084 3560 5127
rect 3639 5125 3647 5147
rect 3677 5143 3683 5217
rect 3797 5276 3809 5282
rect 3877 5276 3889 5282
rect 3917 5276 3929 5282
rect 3971 5276 3983 5282
rect 4011 5276 4023 5282
rect 4042 5276 4054 5282
rect 4092 5276 4104 5282
rect 3739 5161 3747 5196
rect 3820 5189 3837 5196
rect 3857 5197 3873 5203
rect 3667 5137 3683 5143
rect 3733 5125 3741 5147
rect 3820 5141 3827 5189
rect 3640 5118 3665 5125
rect 3597 5104 3649 5107
rect 3438 5058 3450 5064
rect 3488 5058 3500 5064
rect 3609 5098 3637 5104
rect 3657 5104 3665 5118
rect 3715 5118 3740 5125
rect 3715 5104 3723 5118
rect 3731 5104 3783 5107
rect 3743 5098 3771 5104
rect 3820 5084 3827 5127
rect 3857 5123 3863 5197
rect 3897 5181 3905 5236
rect 3927 5197 3943 5203
rect 3857 5117 3873 5123
rect 3897 5118 3905 5167
rect 3897 5112 3921 5118
rect 3909 5104 3921 5112
rect 3531 5058 3543 5064
rect 3571 5058 3583 5064
rect 3617 5058 3629 5064
rect 3751 5058 3763 5064
rect 3797 5058 3809 5064
rect 3837 5058 3849 5064
rect 3937 5083 3943 5197
rect 3995 5181 4003 5236
rect 4127 5282 6736 5284
rect 4151 5276 4163 5282
rect 4191 5276 4203 5282
rect 4247 5276 4259 5282
rect 4291 5276 4303 5282
rect 4107 5217 4153 5223
rect 3995 5118 4003 5167
rect 4073 5161 4081 5196
rect 4175 5181 4183 5236
rect 4331 5276 4343 5282
rect 4371 5276 4383 5282
rect 4416 5276 4428 5282
rect 4466 5276 4478 5282
rect 4079 5125 4087 5147
rect 4080 5118 4105 5125
rect 4175 5118 4183 5167
rect 4231 5161 4239 5196
rect 4231 5147 4233 5161
rect 3979 5112 4003 5118
rect 3979 5104 3991 5112
rect 4037 5104 4089 5107
rect 3937 5077 3953 5083
rect 4049 5098 4077 5104
rect 4097 5104 4105 5118
rect 4159 5112 4183 5118
rect 4159 5104 4171 5112
rect 4231 5104 4239 5147
rect 4274 5122 4282 5236
rect 4307 5197 4333 5203
rect 4355 5181 4363 5236
rect 4516 5276 4528 5282
rect 4566 5276 4578 5282
rect 4497 5217 4513 5223
rect 4265 5114 4303 5122
rect 4355 5118 4363 5167
rect 4439 5161 4447 5196
rect 4433 5125 4441 5147
rect 4497 5143 4503 5217
rect 4597 5276 4609 5282
rect 4637 5276 4649 5282
rect 4677 5276 4689 5282
rect 4717 5276 4729 5282
rect 4757 5276 4769 5282
rect 4851 5276 4863 5282
rect 4891 5276 4903 5282
rect 4539 5161 4547 5196
rect 4617 5181 4625 5236
rect 4647 5197 4663 5203
rect 4497 5137 4513 5143
rect 4533 5125 4541 5147
rect 4291 5104 4303 5114
rect 4231 5094 4241 5104
rect 4339 5112 4363 5118
rect 4415 5118 4440 5125
rect 4515 5118 4540 5125
rect 4617 5118 4625 5167
rect 4657 5127 4663 5197
rect 4697 5181 4705 5236
rect 4727 5197 4753 5203
rect 4737 5177 4753 5183
rect 4339 5104 4351 5112
rect 4415 5104 4423 5118
rect 4431 5104 4483 5107
rect 4515 5104 4523 5118
rect 4617 5112 4641 5118
rect 4697 5118 4705 5167
rect 4737 5147 4743 5177
rect 4776 5153 4784 5236
rect 4835 5234 4843 5236
rect 4922 5276 4934 5282
rect 4972 5276 4984 5282
rect 4871 5234 4882 5236
rect 4835 5228 4882 5234
rect 4697 5112 4721 5118
rect 4443 5098 4471 5104
rect 4531 5104 4583 5107
rect 4629 5104 4641 5112
rect 4709 5104 4721 5112
rect 4543 5098 4571 5104
rect 4776 5084 4784 5139
rect 4797 5127 4803 5193
rect 4835 5173 4842 5228
rect 5017 5276 5029 5282
rect 5077 5276 5089 5282
rect 5117 5276 5129 5282
rect 4987 5217 5003 5223
rect 4953 5161 4961 5196
rect 4817 5127 4823 5153
rect 4836 5131 4844 5159
rect 4836 5122 4866 5131
rect 4959 5125 4967 5147
rect 4997 5143 5003 5217
rect 5157 5274 5169 5282
rect 5197 5276 5209 5282
rect 5036 5161 5044 5196
rect 5097 5181 5105 5236
rect 5237 5276 5249 5282
rect 5277 5276 5289 5282
rect 5322 5276 5334 5282
rect 5372 5276 5384 5282
rect 4987 5137 5003 5143
rect 4836 5120 4854 5122
rect 4960 5118 4985 5125
rect 4917 5104 4969 5107
rect 4929 5098 4957 5104
rect 4977 5104 4985 5118
rect 5036 5104 5044 5147
rect 5097 5118 5105 5167
rect 5179 5153 5188 5196
rect 5257 5181 5265 5236
rect 5287 5217 5303 5223
rect 5179 5139 5193 5153
rect 5097 5112 5121 5118
rect 5109 5104 5121 5112
rect 5179 5104 5188 5139
rect 5257 5118 5265 5167
rect 5297 5123 5303 5217
rect 5417 5276 5429 5282
rect 5457 5276 5469 5282
rect 5517 5276 5529 5282
rect 5557 5276 5569 5282
rect 5617 5276 5629 5282
rect 5677 5276 5689 5282
rect 5717 5276 5729 5282
rect 5782 5276 5794 5282
rect 5832 5276 5844 5282
rect 5438 5234 5449 5236
rect 5477 5234 5485 5236
rect 5438 5228 5485 5234
rect 5538 5234 5549 5236
rect 5577 5234 5585 5236
rect 5538 5228 5585 5234
rect 5353 5161 5361 5196
rect 5478 5173 5485 5228
rect 5257 5112 5281 5118
rect 5297 5117 5313 5123
rect 5359 5125 5367 5147
rect 5387 5137 5413 5143
rect 5476 5131 5484 5159
rect 5497 5143 5503 5193
rect 5578 5173 5585 5228
rect 5597 5177 5613 5183
rect 5497 5137 5533 5143
rect 5576 5131 5584 5159
rect 5360 5118 5385 5125
rect 5269 5104 5281 5112
rect 3879 5058 3891 5064
rect 4009 5058 4021 5064
rect 4057 5058 4069 5064
rect 4189 5058 4201 5064
rect 4261 5058 4273 5064
rect 4369 5058 4381 5064
rect 4451 5058 4463 5064
rect 4551 5058 4563 5064
rect 4599 5058 4611 5064
rect 4679 5058 4691 5064
rect 4757 5058 4769 5064
rect 4890 5058 4902 5064
rect 4937 5058 4949 5064
rect 5017 5058 5029 5064
rect 5079 5058 5091 5064
rect 5157 5058 5169 5064
rect 5197 5058 5209 5064
rect 5317 5104 5369 5107
rect 5329 5098 5357 5104
rect 5377 5104 5385 5118
rect 5454 5122 5484 5131
rect 5466 5120 5484 5122
rect 5554 5122 5584 5131
rect 5566 5120 5584 5122
rect 5597 5103 5603 5177
rect 5636 5153 5644 5236
rect 5698 5234 5709 5236
rect 5737 5234 5745 5236
rect 5698 5228 5745 5234
rect 5738 5173 5745 5228
rect 5891 5276 5903 5282
rect 5931 5276 5943 5282
rect 5957 5276 5969 5282
rect 5997 5276 6009 5282
rect 6057 5276 6069 5282
rect 6097 5276 6109 5282
rect 6191 5276 6203 5282
rect 6271 5276 6283 5282
rect 6331 5276 6343 5282
rect 6371 5276 6383 5282
rect 6431 5276 6443 5282
rect 6471 5276 6483 5282
rect 5813 5161 5821 5196
rect 5915 5181 5923 5236
rect 5978 5234 5989 5236
rect 6017 5234 6025 5236
rect 5978 5228 6025 5234
rect 5587 5097 5603 5103
rect 5636 5084 5644 5139
rect 5736 5131 5744 5159
rect 5714 5122 5744 5131
rect 5819 5125 5827 5147
rect 5857 5143 5863 5173
rect 5847 5137 5863 5143
rect 5726 5120 5744 5122
rect 5820 5118 5845 5125
rect 5915 5118 5923 5167
rect 6018 5173 6025 5228
rect 6077 5181 6085 5236
rect 6107 5197 6123 5203
rect 6016 5131 6024 5159
rect 5777 5104 5829 5107
rect 5789 5098 5817 5104
rect 5837 5104 5845 5118
rect 5899 5112 5923 5118
rect 5899 5104 5911 5112
rect 5239 5058 5251 5064
rect 5337 5058 5349 5064
rect 5418 5058 5430 5064
rect 5518 5058 5530 5064
rect 5617 5058 5629 5064
rect 5678 5058 5690 5064
rect 5797 5058 5809 5064
rect 5929 5058 5941 5064
rect 5994 5122 6024 5131
rect 6006 5120 6024 5122
rect 6077 5118 6085 5167
rect 6077 5112 6101 5118
rect 6089 5104 6101 5112
rect 6117 5107 6123 5197
rect 6211 5202 6223 5204
rect 6183 5196 6223 5202
rect 6154 5161 6162 5196
rect 6207 5177 6243 5183
rect 6154 5104 6162 5147
rect 6237 5127 6243 5177
rect 6256 5153 6264 5236
rect 6315 5234 6323 5236
rect 6351 5234 6362 5236
rect 6315 5228 6362 5234
rect 6415 5234 6423 5236
rect 6497 5276 6509 5282
rect 6591 5276 6603 5282
rect 6631 5276 6643 5282
rect 6451 5234 6462 5236
rect 6415 5228 6462 5234
rect 6287 5177 6303 5183
rect 6154 5093 6180 5104
rect 6256 5084 6264 5139
rect 6297 5103 6303 5177
rect 6315 5173 6322 5228
rect 6387 5217 6403 5223
rect 6397 5167 6403 5217
rect 6415 5173 6422 5228
rect 6316 5131 6324 5159
rect 6416 5131 6424 5159
rect 6516 5153 6524 5236
rect 6575 5234 6583 5236
rect 6657 5276 6669 5282
rect 6697 5276 6709 5282
rect 6611 5234 6622 5236
rect 6575 5228 6622 5234
rect 6316 5122 6346 5131
rect 6316 5120 6334 5122
rect 6287 5097 6303 5103
rect 6416 5122 6446 5131
rect 6416 5120 6434 5122
rect 6516 5084 6524 5139
rect 6557 5103 6563 5213
rect 6575 5173 6582 5228
rect 6677 5181 6685 5236
rect 6576 5131 6584 5159
rect 6576 5122 6606 5131
rect 6576 5120 6594 5122
rect 6557 5097 6573 5103
rect 5958 5058 5970 5064
rect 6059 5058 6071 5064
rect 6158 5058 6170 5064
rect 6208 5058 6220 5064
rect 6271 5058 6283 5064
rect 6370 5058 6382 5064
rect 6470 5058 6482 5064
rect 6677 5118 6685 5167
rect 6717 5127 6723 5193
rect 6677 5112 6701 5118
rect 6689 5104 6701 5112
rect 6497 5058 6509 5064
rect 6630 5058 6642 5064
rect 6659 5058 6671 5064
rect 6742 5058 6802 5522
rect 4 5056 6802 5058
rect 6736 5044 6802 5056
rect 4 5042 6802 5044
rect 49 5036 61 5042
rect 129 5036 141 5042
rect 229 5036 241 5042
rect 279 5036 291 5042
rect 337 5036 349 5042
rect 385 5036 397 5042
rect 447 5036 459 5042
rect 518 5036 530 5042
rect 568 5036 580 5042
rect 649 5036 661 5042
rect 31 4953 39 4996
rect 71 4990 79 5016
rect 57 4984 79 4990
rect 57 4978 60 4984
rect 31 4939 33 4953
rect 31 4904 39 4939
rect 53 4922 60 4978
rect 111 4953 119 4996
rect 151 4990 159 5016
rect 137 4984 159 4990
rect 427 5016 440 5022
rect 311 5010 318 5016
rect 307 5002 318 5010
rect 368 5004 375 5016
rect 433 5010 440 5016
rect 199 4988 211 4996
rect 137 4978 140 4984
rect 199 4982 223 4988
rect 111 4939 113 4953
rect 57 4916 60 4922
rect 57 4910 83 4916
rect 75 4864 83 4910
rect 111 4904 119 4939
rect 133 4922 140 4978
rect 215 4933 223 4982
rect 257 4981 265 4996
rect 368 4997 389 5004
rect 347 4986 353 4988
rect 414 4986 421 4992
rect 257 4967 273 4981
rect 347 4980 421 4986
rect 137 4916 140 4922
rect 137 4910 163 4916
rect 155 4864 163 4910
rect 215 4864 223 4919
rect 257 4904 265 4967
rect 273 4953 287 4967
rect 279 4908 293 4916
rect 347 4908 353 4980
rect 414 4972 421 4980
rect 426 4964 460 4972
rect 454 4959 460 4964
rect 407 4946 434 4953
rect 313 4902 353 4908
rect 361 4908 405 4914
rect 313 4884 319 4902
rect 361 4894 367 4908
rect 473 4912 479 4996
rect 514 4996 540 5007
rect 679 5036 691 5042
rect 809 5036 821 5042
rect 859 5036 871 5042
rect 917 5036 929 5042
rect 965 5036 977 5042
rect 1027 5036 1039 5042
rect 1109 5036 1121 5042
rect 1178 5036 1190 5042
rect 1228 5036 1240 5042
rect 1309 5036 1321 5042
rect 1369 5036 1381 5042
rect 1419 5036 1431 5042
rect 1549 5036 1561 5042
rect 1631 5036 1643 5042
rect 1729 5036 1741 5042
rect 1811 5036 1823 5042
rect 1859 5036 1871 5042
rect 1991 5036 2003 5042
rect 2091 5036 2103 5042
rect 2181 5036 2193 5042
rect 2237 5036 2249 5042
rect 2311 5036 2323 5042
rect 2351 5036 2363 5042
rect 2411 5036 2423 5042
rect 2455 5036 2463 5042
rect 2529 5036 2541 5042
rect 2611 5036 2623 5042
rect 2711 5036 2723 5042
rect 2791 5036 2803 5042
rect 2837 5036 2849 5042
rect 2971 5036 2983 5042
rect 3071 5036 3083 5042
rect 3131 5036 3143 5042
rect 3171 5036 3183 5042
rect 3231 5036 3243 5042
rect 3309 5036 3321 5042
rect 3391 5036 3403 5042
rect 3461 5036 3473 5042
rect 3523 5036 3535 5042
rect 3571 5036 3583 5042
rect 3629 5036 3641 5042
rect 3697 5036 3709 5042
rect 3798 5036 3810 5042
rect 3848 5036 3860 5042
rect 3950 5036 3962 5042
rect 514 4953 522 4996
rect 619 4988 631 4996
rect 709 4988 721 4996
rect 619 4982 643 4988
rect 417 4904 479 4912
rect 514 4904 522 4939
rect 635 4933 643 4982
rect 697 4982 721 4988
rect 1007 5016 1020 5022
rect 891 5010 898 5016
rect 887 5002 898 5010
rect 948 5004 955 5016
rect 1013 5010 1020 5016
rect 779 4988 791 4996
rect 779 4982 803 4988
rect 567 4917 603 4923
rect 697 4933 705 4982
rect 337 4888 367 4894
rect 385 4890 423 4898
rect 415 4884 423 4890
rect 307 4844 319 4878
rect 365 4870 387 4882
rect 415 4870 433 4884
rect 361 4864 373 4870
rect 415 4864 423 4870
rect 543 4898 583 4904
rect 571 4896 583 4898
rect 597 4903 603 4917
rect 597 4897 613 4903
rect 635 4864 643 4919
rect 697 4864 705 4919
rect 737 4887 743 4953
rect 795 4933 803 4982
rect 837 4981 845 4996
rect 948 4997 969 5004
rect 927 4986 933 4988
rect 994 4986 1001 4992
rect 837 4967 853 4981
rect 927 4980 1001 4986
rect 795 4864 803 4919
rect 837 4904 845 4967
rect 853 4953 867 4967
rect 859 4908 873 4916
rect 49 4818 61 4824
rect 129 4818 141 4824
rect 191 4818 203 4824
rect 231 4818 243 4824
rect 277 4818 289 4824
rect 335 4818 347 4824
rect 381 4818 393 4824
rect 447 4818 459 4824
rect 551 4818 563 4824
rect 611 4818 623 4824
rect 651 4818 663 4824
rect 677 4818 689 4824
rect 717 4818 729 4824
rect 927 4908 933 4980
rect 994 4972 1001 4980
rect 1006 4964 1040 4972
rect 1034 4959 1040 4964
rect 987 4946 1014 4953
rect 893 4902 933 4908
rect 941 4908 985 4914
rect 893 4884 899 4902
rect 941 4894 947 4908
rect 1053 4912 1059 4996
rect 997 4904 1059 4912
rect 1091 4953 1099 4996
rect 1131 4990 1139 5016
rect 1117 4984 1139 4990
rect 1174 4996 1200 5007
rect 1117 4978 1120 4984
rect 1091 4939 1093 4953
rect 1091 4904 1099 4939
rect 1113 4922 1120 4978
rect 1174 4953 1182 4996
rect 1117 4916 1120 4922
rect 1117 4910 1143 4916
rect 917 4888 947 4894
rect 965 4890 1003 4898
rect 995 4884 1003 4890
rect 887 4844 899 4878
rect 945 4870 967 4882
rect 995 4870 1013 4884
rect 941 4864 953 4870
rect 995 4864 1003 4870
rect 1135 4864 1143 4910
rect 1174 4904 1182 4939
rect 1257 4923 1263 4993
rect 1279 4988 1291 4996
rect 1279 4982 1303 4988
rect 1295 4933 1303 4982
rect 1351 4953 1359 4996
rect 1391 4990 1399 5016
rect 1377 4984 1399 4990
rect 1449 4988 1461 4996
rect 1377 4978 1380 4984
rect 1227 4917 1263 4923
rect 1351 4939 1353 4953
rect 1203 4898 1243 4904
rect 1231 4896 1243 4898
rect 1295 4864 1303 4919
rect 1351 4904 1359 4939
rect 1373 4922 1380 4978
rect 1437 4982 1461 4988
rect 1519 4988 1531 4996
rect 1519 4982 1543 4988
rect 1437 4933 1445 4982
rect 1377 4916 1380 4922
rect 1535 4933 1543 4982
rect 1595 4982 1603 4996
rect 1623 4996 1651 5002
rect 1611 4993 1663 4996
rect 1595 4975 1620 4982
rect 1613 4953 1621 4975
rect 1377 4910 1403 4916
rect 1395 4864 1403 4910
rect 1437 4864 1445 4919
rect 1535 4864 1543 4919
rect 1619 4904 1627 4939
rect 1677 4907 1683 4993
rect 1699 4988 1711 4996
rect 1699 4982 1723 4988
rect 1715 4933 1723 4982
rect 1775 4982 1783 4996
rect 1803 4996 1831 5002
rect 1791 4993 1843 4996
rect 1889 4988 1901 4996
rect 1877 4982 1901 4988
rect 1955 4982 1963 4996
rect 1983 4996 2011 5002
rect 1971 4993 2023 4996
rect 2055 4982 2063 4996
rect 2083 4996 2111 5002
rect 2071 4993 2123 4996
rect 2151 4996 2161 5006
rect 1775 4975 1800 4982
rect 1793 4953 1801 4975
rect 771 4818 783 4824
rect 811 4818 823 4824
rect 857 4818 869 4824
rect 915 4818 927 4824
rect 961 4818 973 4824
rect 1027 4818 1039 4824
rect 1109 4818 1121 4824
rect 1211 4818 1223 4824
rect 1271 4818 1283 4824
rect 1311 4818 1323 4824
rect 1369 4818 1381 4824
rect 1417 4818 1429 4824
rect 1457 4818 1469 4824
rect 1511 4818 1523 4824
rect 1551 4818 1563 4824
rect 1715 4864 1723 4919
rect 1799 4904 1807 4939
rect 1877 4933 1885 4982
rect 1955 4975 1980 4982
rect 2055 4975 2080 4982
rect 1973 4953 1981 4975
rect 2073 4953 2081 4975
rect 1596 4818 1608 4824
rect 1646 4818 1658 4824
rect 1691 4818 1703 4824
rect 1731 4818 1743 4824
rect 1877 4864 1885 4919
rect 1917 4903 1923 4913
rect 1979 4904 1987 4939
rect 1907 4897 1923 4903
rect 1776 4818 1788 4824
rect 1826 4818 1838 4824
rect 1857 4818 1869 4824
rect 1897 4818 1909 4824
rect 2037 4883 2043 4953
rect 2151 4953 2159 4996
rect 2211 4986 2223 4996
rect 2185 4978 2223 4986
rect 2151 4939 2153 4953
rect 2079 4904 2087 4939
rect 2151 4904 2159 4939
rect 2037 4877 2053 4883
rect 1956 4818 1968 4824
rect 2006 4818 2018 4824
rect -62 4816 2033 4818
rect 2194 4864 2202 4978
rect 2256 4961 2264 5016
rect 2333 4973 2340 5016
rect 2393 4961 2400 4996
rect 2431 4988 2437 5016
rect 2427 4982 2437 4988
rect 2499 4988 2511 4996
rect 2499 4982 2523 4988
rect 2256 4864 2264 4947
rect 2333 4911 2340 4959
rect 2323 4904 2340 4911
rect 2056 4818 2068 4824
rect 2106 4818 2118 4824
rect 2167 4818 2179 4824
rect 2211 4818 2223 4824
rect 2397 4903 2406 4947
rect 2416 4921 2422 4976
rect 2515 4933 2523 4982
rect 2575 4982 2583 4996
rect 2603 4996 2631 5002
rect 2591 4993 2643 4996
rect 2675 4982 2683 4996
rect 2703 4996 2731 5002
rect 2691 4993 2743 4996
rect 2575 4975 2600 4982
rect 2675 4975 2700 4982
rect 2593 4953 2601 4975
rect 2427 4912 2463 4920
rect 2693 4953 2701 4975
rect 2776 4961 2784 5016
rect 2829 4996 2857 5002
rect 2817 4993 2869 4996
rect 2877 4982 2885 4996
rect 2860 4975 2885 4982
rect 2935 4982 2943 4996
rect 2963 4996 2991 5002
rect 2951 4993 3003 4996
rect 3035 4982 3043 4996
rect 3063 4996 3091 5002
rect 3051 4993 3103 4996
rect 2935 4975 2960 4982
rect 3035 4975 3060 4982
rect 2455 4904 2463 4912
rect 2397 4894 2401 4903
rect 2515 4864 2523 4919
rect 2599 4904 2607 4939
rect 2699 4904 2707 4939
rect 2237 4818 2249 4824
rect 2351 4818 2363 4824
rect 2421 4818 2433 4824
rect 2491 4818 2503 4824
rect 2531 4818 2543 4824
rect 2047 4816 2553 4818
rect 2576 4818 2588 4824
rect 2626 4818 2638 4824
rect 2776 4864 2784 4947
rect 2859 4953 2867 4975
rect 2953 4953 2961 4975
rect 3053 4953 3061 4975
rect 3153 4973 3160 5016
rect 2853 4904 2861 4939
rect 2959 4904 2967 4939
rect 3059 4904 3067 4939
rect 3153 4911 3160 4959
rect 3216 4953 3224 4996
rect 3279 4988 3291 4996
rect 3279 4982 3303 4988
rect 3143 4904 3160 4911
rect 3216 4904 3224 4939
rect 3295 4933 3303 4982
rect 3355 4982 3363 4996
rect 3383 4996 3411 5002
rect 3371 4993 3423 4996
rect 3480 5016 3493 5022
rect 3480 5010 3487 5016
rect 3545 5004 3552 5016
rect 3355 4975 3380 4982
rect 3373 4953 3381 4975
rect 2676 4818 2688 4824
rect 2726 4818 2738 4824
rect 2791 4818 2803 4824
rect 2822 4818 2834 4824
rect 2872 4818 2884 4824
rect 2567 4816 2913 4818
rect 2936 4818 2948 4824
rect 2986 4818 2998 4824
rect 3295 4864 3303 4919
rect 3379 4904 3387 4939
rect 3441 4912 3447 4996
rect 3531 4997 3552 5004
rect 3602 5010 3609 5016
rect 3602 5002 3613 5010
rect 3499 4986 3506 4992
rect 3567 4986 3573 4988
rect 3499 4980 3573 4986
rect 3655 4981 3663 4996
rect 3689 4996 3717 5002
rect 3677 4993 3729 4996
rect 3794 4996 3820 5007
rect 3877 4997 3893 5003
rect 3737 4982 3745 4996
rect 3499 4972 3506 4980
rect 3460 4964 3494 4972
rect 3460 4959 3466 4964
rect 3486 4946 3513 4953
rect 3441 4904 3503 4912
rect 3515 4908 3559 4914
rect 3036 4818 3048 4824
rect 3086 4818 3098 4824
rect 3171 4818 3183 4824
rect 3231 4818 3243 4824
rect 3271 4818 3283 4824
rect 3311 4818 3323 4824
rect 3497 4890 3535 4898
rect 3553 4894 3559 4908
rect 3567 4908 3573 4980
rect 3647 4967 3663 4981
rect 3720 4975 3745 4982
rect 3633 4953 3647 4967
rect 3567 4902 3607 4908
rect 3627 4908 3641 4916
rect 3655 4904 3663 4967
rect 3719 4953 3727 4975
rect 3794 4953 3802 4996
rect 3713 4904 3721 4939
rect 3794 4904 3802 4939
rect 3877 4923 3883 4997
rect 3896 4978 3914 4980
rect 3896 4969 3926 4978
rect 3998 5036 4010 5042
rect 4048 5036 4060 5042
rect 4111 5036 4123 5042
rect 4181 5036 4193 5042
rect 4289 5036 4301 5042
rect 4347 5036 4359 5042
rect 4471 5036 4483 5042
rect 4518 5036 4530 5042
rect 4637 5036 4649 5042
rect 4769 5036 4781 5042
rect 4841 5036 4853 5042
rect 4949 5036 4961 5042
rect 3994 4996 4020 5007
rect 4151 4996 4161 5006
rect 3896 4941 3904 4969
rect 3994 4953 4002 4996
rect 4096 4953 4104 4996
rect 4151 4953 4159 4996
rect 4211 4986 4223 4996
rect 4185 4978 4223 4986
rect 4379 4996 4389 5006
rect 4259 4988 4271 4996
rect 4259 4982 4283 4988
rect 4151 4939 4153 4953
rect 3847 4917 3883 4923
rect 3497 4884 3505 4890
rect 3553 4888 3583 4894
rect 3601 4884 3607 4902
rect 3487 4870 3505 4884
rect 3533 4870 3555 4882
rect 3497 4864 3505 4870
rect 3547 4864 3559 4870
rect 3601 4844 3613 4878
rect 3823 4898 3863 4904
rect 3851 4896 3863 4898
rect 3895 4872 3902 4927
rect 3994 4904 4002 4939
rect 4027 4917 4073 4923
rect 4096 4904 4104 4939
rect 4151 4904 4159 4939
rect 3895 4866 3942 4872
rect 3895 4864 3903 4866
rect 3931 4864 3942 4866
rect 4023 4898 4063 4904
rect 4051 4896 4063 4898
rect 4194 4864 4202 4978
rect 4275 4933 4283 4982
rect 4317 4986 4329 4996
rect 4317 4978 4355 4986
rect 4275 4864 4283 4919
rect 4338 4864 4346 4978
rect 4381 4953 4389 4996
rect 4435 4982 4443 4996
rect 4463 4996 4491 5002
rect 4451 4993 4503 4996
rect 4435 4975 4460 4982
rect 4629 4996 4657 5002
rect 4617 4993 4669 4996
rect 4811 4996 4821 5006
rect 4677 4982 4685 4996
rect 4739 4988 4751 4996
rect 4739 4982 4763 4988
rect 4566 4978 4584 4980
rect 4387 4939 4389 4953
rect 4453 4953 4461 4975
rect 4554 4969 4584 4978
rect 4660 4975 4685 4982
rect 4576 4941 4584 4969
rect 4381 4904 4389 4939
rect 4459 4904 4467 4939
rect 4659 4953 4667 4975
rect 4687 4957 4703 4963
rect 3356 4818 3368 4824
rect 3406 4818 3418 4824
rect 3461 4818 3473 4824
rect 3527 4818 3539 4824
rect 3573 4818 3585 4824
rect 3631 4818 3643 4824
rect 3682 4818 3694 4824
rect 3732 4818 3744 4824
rect 3831 4818 3843 4824
rect 3911 4818 3923 4824
rect 3951 4818 3963 4824
rect 4031 4818 4043 4824
rect 4111 4818 4123 4824
rect 4167 4818 4179 4824
rect 4211 4818 4223 4824
rect 4251 4818 4263 4824
rect 4291 4818 4303 4824
rect 4317 4818 4329 4824
rect 4361 4818 4373 4824
rect 2927 4816 4413 4818
rect 4578 4872 4585 4927
rect 4653 4904 4661 4939
rect 4538 4866 4585 4872
rect 4538 4864 4549 4866
rect 4436 4818 4448 4824
rect 4486 4818 4498 4824
rect 4577 4864 4585 4866
rect 4697 4883 4703 4957
rect 4755 4933 4763 4982
rect 4811 4953 4819 4996
rect 4871 4986 4883 4996
rect 4979 5036 4991 5042
rect 5087 5036 5099 5042
rect 5209 5036 5221 5042
rect 5281 5036 5293 5042
rect 5367 5036 5379 5042
rect 5472 5036 5484 5042
rect 5528 5036 5540 5042
rect 5609 5036 5621 5042
rect 4919 4988 4931 4996
rect 5009 4988 5021 4996
rect 4845 4978 4883 4986
rect 4811 4939 4813 4953
rect 4717 4903 4723 4913
rect 4717 4897 4733 4903
rect 4687 4877 4703 4883
rect 4755 4864 4763 4919
rect 4811 4904 4819 4939
rect 4517 4818 4529 4824
rect 4557 4818 4569 4824
rect 4622 4818 4634 4824
rect 4672 4818 4684 4824
rect 4854 4864 4862 4978
rect 4919 4982 4943 4988
rect 4897 4903 4903 4973
rect 4935 4933 4943 4982
rect 4997 4982 5021 4988
rect 5119 4996 5129 5006
rect 5057 4986 5069 4996
rect 4997 4933 5005 4982
rect 5057 4978 5095 4986
rect 4897 4897 4913 4903
rect 4935 4864 4943 4919
rect 4997 4864 5005 4919
rect 5078 4864 5086 4978
rect 5121 4953 5129 4996
rect 5251 4996 5261 5006
rect 5179 4988 5191 4996
rect 5179 4982 5203 4988
rect 5127 4939 5129 4953
rect 5121 4904 5129 4939
rect 5195 4933 5203 4982
rect 5251 4953 5259 4996
rect 5311 4986 5323 4996
rect 5285 4978 5323 4986
rect 5399 4996 5409 5006
rect 5638 5036 5650 5042
rect 5758 5036 5770 5042
rect 5808 5036 5820 5042
rect 5910 5036 5922 5042
rect 5989 5036 6001 5042
rect 5337 4986 5349 4996
rect 5337 4978 5375 4986
rect 5251 4939 5253 4953
rect 4731 4818 4743 4824
rect 4771 4818 4783 4824
rect 4827 4818 4839 4824
rect 4871 4818 4883 4824
rect 4911 4818 4923 4824
rect 4951 4818 4963 4824
rect 4977 4818 4989 4824
rect 5017 4818 5029 4824
rect 5195 4864 5203 4919
rect 5251 4904 5259 4939
rect 5294 4864 5302 4978
rect 5358 4864 5366 4978
rect 5401 4953 5409 4996
rect 5407 4939 5409 4953
rect 5500 4953 5507 4996
rect 5579 4988 5591 4996
rect 5579 4982 5603 4988
rect 5401 4904 5409 4939
rect 5493 4916 5499 4939
rect 5595 4933 5603 4982
rect 5754 4996 5780 5007
rect 5837 4997 5853 5003
rect 5686 4978 5704 4980
rect 5674 4969 5704 4978
rect 5696 4941 5704 4969
rect 5754 4953 5762 4996
rect 5472 4910 5499 4916
rect 5472 4904 5484 4910
rect 5057 4818 5069 4824
rect 5101 4818 5113 4824
rect 5171 4818 5183 4824
rect 5211 4818 5223 4824
rect 5267 4818 5279 4824
rect 5311 4818 5323 4824
rect 5463 4824 5491 4830
rect 5503 4896 5531 4902
rect 5595 4864 5603 4919
rect 5698 4872 5705 4927
rect 5754 4904 5762 4939
rect 5837 4923 5843 4997
rect 5856 4978 5874 4980
rect 5856 4969 5886 4978
rect 6020 5036 6032 5042
rect 6076 5036 6088 5042
rect 6210 5036 6222 5042
rect 6257 5036 6269 5042
rect 6410 5036 6422 5042
rect 6510 5036 6522 5042
rect 6137 4997 6153 5003
rect 5959 4988 5971 4996
rect 5959 4982 5983 4988
rect 5856 4941 5864 4969
rect 5927 4957 5943 4963
rect 5787 4917 5843 4923
rect 5658 4866 5705 4872
rect 5658 4864 5669 4866
rect 5337 4818 5349 4824
rect 5381 4818 5393 4824
rect 5511 4818 5523 4824
rect 5571 4818 5583 4824
rect 5611 4818 5623 4824
rect 5697 4864 5705 4866
rect 5783 4898 5823 4904
rect 5811 4896 5823 4898
rect 5855 4872 5862 4927
rect 5937 4883 5943 4957
rect 5975 4933 5983 4982
rect 6053 4953 6060 4996
rect 5927 4877 5943 4883
rect 5855 4866 5902 4872
rect 5855 4864 5863 4866
rect 5891 4864 5902 4866
rect 5975 4864 5983 4919
rect 6061 4916 6067 4939
rect 6061 4910 6088 4916
rect 6076 4904 6088 4910
rect 6137 4907 6143 4997
rect 6156 4978 6174 4980
rect 6156 4969 6186 4978
rect 6249 4996 6277 5002
rect 6237 4993 6289 4996
rect 6297 4982 6305 4996
rect 6280 4975 6305 4982
rect 6356 4978 6374 4980
rect 6156 4941 6164 4969
rect 6279 4953 6287 4975
rect 6356 4969 6386 4978
rect 6456 4978 6474 4980
rect 6456 4969 6486 4978
rect 6539 5036 6551 5042
rect 6651 5036 6663 5042
rect 6569 4988 6581 4996
rect 6557 4982 6581 4988
rect 6356 4941 6364 4969
rect 6456 4941 6464 4969
rect 5637 4818 5649 4824
rect 5677 4818 5689 4824
rect 5791 4818 5803 4824
rect 5871 4818 5883 4824
rect 5911 4818 5923 4824
rect 6029 4896 6057 4902
rect 6069 4824 6097 4830
rect 6155 4872 6162 4927
rect 6273 4904 6281 4939
rect 6317 4917 6333 4923
rect 6155 4866 6202 4872
rect 6155 4864 6163 4866
rect 6191 4864 6202 4866
rect 5951 4818 5963 4824
rect 5991 4818 6003 4824
rect 6037 4818 6049 4824
rect 6171 4818 6183 4824
rect 6211 4818 6223 4824
rect 6317 4883 6323 4917
rect 6307 4877 6323 4883
rect 6355 4872 6362 4927
rect 6455 4872 6462 4927
rect 6557 4933 6565 4982
rect 6617 4927 6623 4993
rect 6636 4961 6644 5016
rect 6355 4866 6402 4872
rect 6355 4864 6363 4866
rect 6391 4864 6402 4866
rect 6455 4866 6502 4872
rect 6455 4864 6463 4866
rect 6491 4864 6502 4866
rect 6557 4864 6565 4919
rect 6636 4864 6644 4947
rect 6242 4818 6254 4824
rect 6292 4818 6304 4824
rect 6371 4818 6383 4824
rect 6411 4818 6423 4824
rect 6471 4818 6483 4824
rect 6511 4818 6523 4824
rect 6537 4818 6549 4824
rect 6577 4818 6589 4824
rect 6651 4818 6663 4824
rect 4427 4816 6736 4818
rect -62 4804 4 4816
rect -62 4802 1673 4804
rect -62 4338 -2 4802
rect 17 4796 29 4802
rect 57 4796 69 4802
rect 97 4796 109 4802
rect 137 4796 149 4802
rect 177 4796 189 4802
rect 271 4796 283 4802
rect 331 4796 343 4802
rect 411 4796 423 4802
rect 491 4796 503 4802
rect 571 4796 583 4802
rect 627 4796 639 4802
rect 671 4796 683 4802
rect 37 4710 49 4716
rect 77 4710 89 4716
rect 117 4710 129 4716
rect 157 4710 169 4716
rect 37 4702 63 4710
rect 77 4702 102 4710
rect 117 4702 142 4710
rect 157 4702 175 4710
rect 243 4709 260 4716
rect 55 4656 63 4702
rect 94 4656 102 4702
rect 134 4656 142 4702
rect 168 4673 175 4702
rect 168 4659 173 4673
rect 253 4661 260 4709
rect 316 4673 324 4756
rect 431 4722 443 4724
rect 403 4716 443 4722
rect 374 4681 382 4716
rect 55 4644 70 4656
rect 94 4644 110 4656
rect 134 4644 150 4656
rect 55 4638 63 4644
rect 94 4638 102 4644
rect 134 4638 142 4644
rect 168 4638 175 4659
rect 36 4630 63 4638
rect 77 4630 102 4638
rect 116 4630 142 4638
rect 156 4631 175 4638
rect 476 4673 484 4756
rect 697 4796 709 4802
rect 809 4796 821 4802
rect 871 4796 883 4802
rect 911 4796 923 4802
rect 957 4796 969 4802
rect 1015 4796 1027 4802
rect 1061 4796 1073 4802
rect 1127 4796 1139 4802
rect 1196 4796 1208 4802
rect 1246 4796 1258 4802
rect 543 4709 560 4716
rect 156 4630 174 4631
rect 36 4624 48 4630
rect 77 4624 89 4630
rect 116 4624 128 4630
rect 156 4624 168 4630
rect 253 4604 260 4647
rect 316 4604 324 4659
rect 357 4623 363 4653
rect 347 4617 363 4623
rect 374 4624 382 4667
rect 553 4661 560 4709
rect 611 4681 619 4716
rect 611 4667 613 4681
rect 374 4613 400 4624
rect 17 4578 29 4584
rect 57 4578 69 4584
rect 97 4578 109 4584
rect 137 4578 149 4584
rect 177 4578 189 4584
rect 231 4578 243 4584
rect 271 4578 283 4584
rect 331 4578 343 4584
rect 476 4604 484 4659
rect 553 4604 560 4647
rect 611 4624 619 4667
rect 654 4642 662 4756
rect 720 4709 737 4716
rect 720 4661 727 4709
rect 791 4681 799 4716
rect 835 4710 843 4756
rect 817 4704 843 4710
rect 817 4698 820 4704
rect 895 4701 903 4756
rect 987 4742 999 4776
rect 1041 4750 1053 4756
rect 1095 4750 1103 4756
rect 1045 4738 1067 4750
rect 1095 4736 1113 4750
rect 993 4718 999 4736
rect 1017 4726 1047 4732
rect 1095 4730 1103 4736
rect 791 4667 793 4681
rect 645 4634 683 4642
rect 671 4624 683 4634
rect 611 4614 621 4624
rect 378 4578 390 4584
rect 428 4578 440 4584
rect 491 4578 503 4584
rect 720 4604 727 4647
rect 791 4624 799 4667
rect 813 4642 820 4698
rect 817 4636 820 4642
rect 895 4638 903 4687
rect 817 4630 839 4636
rect 831 4604 839 4630
rect 879 4632 903 4638
rect 937 4653 945 4716
rect 959 4704 973 4712
rect 993 4712 1033 4718
rect 953 4653 967 4667
rect 937 4639 953 4653
rect 1027 4640 1033 4712
rect 1041 4712 1047 4726
rect 1065 4722 1103 4730
rect 1291 4796 1303 4802
rect 1331 4796 1343 4802
rect 1357 4796 1369 4802
rect 1397 4796 1409 4802
rect 1456 4796 1468 4802
rect 1506 4796 1518 4802
rect 1041 4706 1085 4712
rect 1097 4708 1159 4716
rect 1087 4667 1114 4674
rect 1134 4656 1140 4661
rect 1106 4648 1140 4656
rect 1094 4640 1101 4648
rect 879 4624 891 4632
rect 937 4624 945 4639
rect 1027 4634 1101 4640
rect 1027 4632 1033 4634
rect 1094 4628 1101 4634
rect 987 4610 998 4618
rect 991 4604 998 4610
rect 1048 4616 1069 4623
rect 1153 4624 1159 4708
rect 1219 4681 1227 4716
rect 1315 4701 1323 4756
rect 1377 4701 1385 4756
rect 1407 4737 1433 4743
rect 1407 4717 1423 4723
rect 1213 4645 1221 4667
rect 1195 4638 1220 4645
rect 1315 4638 1323 4687
rect 1195 4624 1203 4638
rect 1299 4632 1323 4638
rect 1377 4638 1385 4687
rect 1417 4663 1423 4717
rect 1537 4796 1549 4802
rect 1617 4796 1629 4802
rect 1687 4802 1813 4804
rect 1697 4796 1709 4802
rect 1757 4796 1769 4802
rect 1479 4681 1487 4716
rect 1560 4709 1577 4716
rect 1640 4709 1657 4716
rect 1417 4657 1433 4663
rect 1473 4645 1481 4667
rect 1560 4661 1567 4709
rect 1640 4661 1647 4709
rect 1716 4673 1724 4756
rect 1827 4802 3733 4804
rect 1842 4796 1854 4802
rect 1892 4796 1904 4802
rect 1957 4796 1969 4802
rect 2015 4796 2027 4802
rect 2061 4796 2073 4802
rect 2127 4796 2139 4802
rect 2191 4796 2203 4802
rect 2231 4796 2243 4802
rect 2301 4796 2313 4802
rect 2357 4796 2369 4802
rect 2397 4796 2409 4802
rect 1987 4742 1999 4776
rect 2041 4750 2053 4756
rect 2095 4750 2103 4756
rect 2045 4738 2067 4750
rect 2095 4736 2113 4750
rect 1993 4718 1999 4736
rect 2017 4726 2047 4732
rect 2095 4730 2103 4736
rect 1455 4638 1480 4645
rect 1377 4632 1401 4638
rect 1048 4604 1055 4616
rect 1113 4604 1120 4610
rect 1107 4598 1120 4604
rect 1211 4624 1263 4627
rect 1223 4618 1251 4624
rect 1299 4624 1311 4632
rect 1389 4624 1401 4632
rect 1455 4624 1463 4638
rect 531 4578 543 4584
rect 571 4578 583 4584
rect 641 4578 653 4584
rect 697 4578 709 4584
rect 737 4578 749 4584
rect 809 4578 821 4584
rect 909 4578 921 4584
rect 959 4578 971 4584
rect 1017 4578 1029 4584
rect 1065 4578 1077 4584
rect 1127 4578 1139 4584
rect 1231 4578 1243 4584
rect 1329 4578 1341 4584
rect 1471 4624 1523 4627
rect 1483 4618 1511 4624
rect 1560 4604 1567 4647
rect 1640 4604 1647 4647
rect 1716 4604 1724 4659
rect 1737 4643 1743 4713
rect 1780 4709 1797 4716
rect 1780 4661 1787 4709
rect 1737 4637 1753 4643
rect 1780 4604 1787 4647
rect 1817 4627 1823 4693
rect 1873 4681 1881 4716
rect 1879 4645 1887 4667
rect 1937 4653 1945 4716
rect 1959 4704 1973 4712
rect 1993 4712 2033 4718
rect 1953 4653 1967 4667
rect 1880 4638 1905 4645
rect 1837 4624 1889 4627
rect 1359 4578 1371 4584
rect 1491 4578 1503 4584
rect 1537 4578 1549 4584
rect 1577 4578 1589 4584
rect 1617 4578 1629 4584
rect 1657 4578 1669 4584
rect 1849 4618 1877 4624
rect 1897 4624 1905 4638
rect 1937 4639 1953 4653
rect 2027 4640 2033 4712
rect 2041 4712 2047 4726
rect 2065 4722 2103 4730
rect 2041 4706 2085 4712
rect 2097 4708 2159 4716
rect 2087 4667 2114 4674
rect 2134 4656 2140 4661
rect 2106 4648 2140 4656
rect 2094 4640 2101 4648
rect 1937 4624 1945 4639
rect 2027 4634 2101 4640
rect 2027 4632 2033 4634
rect 2094 4628 2101 4634
rect 1987 4610 1998 4618
rect 1991 4604 1998 4610
rect 2048 4616 2069 4623
rect 2153 4624 2159 4708
rect 2215 4701 2223 4756
rect 2277 4717 2281 4726
rect 2215 4638 2223 4687
rect 2277 4673 2286 4717
rect 2437 4796 2449 4802
rect 2537 4796 2549 4802
rect 2651 4796 2663 4802
rect 2697 4796 2709 4802
rect 2755 4796 2767 4802
rect 2801 4796 2813 4802
rect 2867 4796 2879 4802
rect 2922 4796 2934 4802
rect 2972 4796 2984 4802
rect 3037 4796 3049 4802
rect 3095 4796 3107 4802
rect 3141 4796 3153 4802
rect 3207 4796 3219 4802
rect 3277 4796 3289 4802
rect 3335 4796 3347 4802
rect 3381 4796 3393 4802
rect 3447 4796 3459 4802
rect 3516 4796 3528 4802
rect 3566 4796 3578 4802
rect 3631 4796 3643 4802
rect 2335 4708 2343 4716
rect 2307 4700 2343 4708
rect 2377 4701 2385 4756
rect 2517 4722 2529 4724
rect 2517 4716 2557 4722
rect 2460 4709 2477 4716
rect 2048 4604 2055 4616
rect 2113 4604 2120 4610
rect 2107 4598 2120 4604
rect 2199 4632 2223 4638
rect 2199 4624 2211 4632
rect 2273 4624 2280 4659
rect 2296 4644 2302 4699
rect 2377 4638 2385 4687
rect 2460 4661 2467 4709
rect 2507 4697 2553 4703
rect 2578 4681 2586 4716
rect 2636 4673 2644 4756
rect 2727 4742 2739 4776
rect 2781 4750 2793 4756
rect 2835 4750 2843 4756
rect 2785 4738 2807 4750
rect 2835 4736 2853 4750
rect 2733 4718 2739 4736
rect 2757 4726 2787 4732
rect 2835 4730 2843 4736
rect 2307 4632 2317 4638
rect 2377 4632 2401 4638
rect 2311 4604 2317 4632
rect 2389 4624 2401 4632
rect 1697 4578 1709 4584
rect 1757 4578 1769 4584
rect 1797 4578 1809 4584
rect 1857 4578 1869 4584
rect 1959 4578 1971 4584
rect 2017 4578 2029 4584
rect 2065 4578 2077 4584
rect 2127 4578 2139 4584
rect 2229 4578 2241 4584
rect 2291 4578 2303 4584
rect 2335 4578 2343 4584
rect 2460 4604 2467 4647
rect 2578 4624 2586 4667
rect 2359 4578 2371 4584
rect 2437 4578 2449 4584
rect 2477 4578 2489 4584
rect 2560 4613 2586 4624
rect 2636 4604 2644 4659
rect 2677 4653 2685 4716
rect 2699 4704 2713 4712
rect 2733 4712 2773 4718
rect 2693 4653 2707 4667
rect 2677 4639 2693 4653
rect 2767 4640 2773 4712
rect 2781 4712 2787 4726
rect 2805 4722 2843 4730
rect 3067 4742 3079 4776
rect 3121 4750 3133 4756
rect 3175 4750 3183 4756
rect 3125 4738 3147 4750
rect 3175 4736 3193 4750
rect 3073 4718 3079 4736
rect 3097 4726 3127 4732
rect 3175 4730 3183 4736
rect 2781 4706 2825 4712
rect 2837 4708 2899 4716
rect 2827 4667 2854 4674
rect 2874 4656 2880 4661
rect 2846 4648 2880 4656
rect 2834 4640 2841 4648
rect 2677 4624 2685 4639
rect 2767 4634 2841 4640
rect 2767 4632 2773 4634
rect 2834 4628 2841 4634
rect 2727 4610 2738 4618
rect 2731 4604 2738 4610
rect 2788 4616 2809 4623
rect 2893 4624 2899 4708
rect 2953 4681 2961 4716
rect 2959 4645 2967 4667
rect 3017 4653 3025 4716
rect 3039 4704 3053 4712
rect 3073 4712 3113 4718
rect 3033 4653 3047 4667
rect 2960 4638 2985 4645
rect 2788 4604 2795 4616
rect 2853 4604 2860 4610
rect 2847 4598 2860 4604
rect 2917 4624 2969 4627
rect 2929 4618 2957 4624
rect 2977 4624 2985 4638
rect 3017 4639 3033 4653
rect 3107 4640 3113 4712
rect 3121 4712 3127 4726
rect 3145 4722 3183 4730
rect 3121 4706 3165 4712
rect 3177 4708 3239 4716
rect 3167 4667 3194 4674
rect 3214 4656 3220 4661
rect 3186 4648 3220 4656
rect 3174 4640 3181 4648
rect 3017 4624 3025 4639
rect 3107 4634 3181 4640
rect 3107 4632 3113 4634
rect 3174 4628 3181 4634
rect 3067 4610 3078 4618
rect 3071 4604 3078 4610
rect 3128 4616 3149 4623
rect 3233 4624 3239 4708
rect 3128 4604 3135 4616
rect 3193 4604 3200 4610
rect 3187 4598 3200 4604
rect 3307 4742 3319 4776
rect 3361 4750 3373 4756
rect 3415 4750 3423 4756
rect 3365 4738 3387 4750
rect 3415 4736 3433 4750
rect 3313 4718 3319 4736
rect 3337 4726 3367 4732
rect 3415 4730 3423 4736
rect 3257 4653 3265 4716
rect 3279 4704 3293 4712
rect 3313 4712 3353 4718
rect 3273 4653 3287 4667
rect 3257 4639 3273 4653
rect 3347 4640 3353 4712
rect 3361 4712 3367 4726
rect 3385 4722 3423 4730
rect 3671 4796 3683 4802
rect 3711 4796 3723 4802
rect 3747 4802 6736 4804
rect 3756 4796 3768 4802
rect 3806 4796 3818 4802
rect 3861 4796 3873 4802
rect 3927 4796 3939 4802
rect 3973 4796 3985 4802
rect 4031 4796 4043 4802
rect 4111 4796 4123 4802
rect 3361 4706 3405 4712
rect 3417 4708 3479 4716
rect 3407 4667 3434 4674
rect 3454 4656 3460 4661
rect 3426 4648 3460 4656
rect 3414 4640 3421 4648
rect 3257 4624 3265 4639
rect 3347 4634 3421 4640
rect 3347 4632 3353 4634
rect 3414 4628 3421 4634
rect 3307 4610 3318 4618
rect 3311 4604 3318 4610
rect 3368 4616 3389 4623
rect 3473 4624 3479 4708
rect 3539 4681 3547 4716
rect 3616 4681 3624 4716
rect 3695 4701 3703 4756
rect 3727 4717 3743 4723
rect 3533 4645 3541 4667
rect 3515 4638 3540 4645
rect 3515 4624 3523 4638
rect 3368 4604 3375 4616
rect 3433 4604 3440 4610
rect 3427 4598 3440 4604
rect 3531 4624 3583 4627
rect 3616 4624 3624 4667
rect 3695 4638 3703 4687
rect 3679 4632 3703 4638
rect 3737 4643 3743 4717
rect 3897 4750 3905 4756
rect 3947 4750 3959 4756
rect 3887 4736 3905 4750
rect 3933 4738 3955 4750
rect 4001 4742 4013 4776
rect 3897 4730 3905 4736
rect 3897 4722 3935 4730
rect 3953 4726 3983 4732
rect 3779 4681 3787 4716
rect 3841 4708 3903 4716
rect 3773 4645 3781 4667
rect 3727 4637 3743 4643
rect 3755 4638 3780 4645
rect 3679 4624 3691 4632
rect 3755 4624 3763 4638
rect 3543 4618 3571 4624
rect 3771 4624 3823 4627
rect 3783 4618 3811 4624
rect 3841 4624 3847 4708
rect 3953 4712 3959 4726
rect 4001 4718 4007 4736
rect 3915 4706 3959 4712
rect 3967 4712 4007 4718
rect 3886 4667 3913 4674
rect 3860 4656 3866 4661
rect 3860 4648 3894 4656
rect 3899 4640 3906 4648
rect 3967 4640 3973 4712
rect 4151 4796 4163 4802
rect 4191 4796 4203 4802
rect 4237 4796 4249 4802
rect 4295 4796 4307 4802
rect 4341 4796 4353 4802
rect 4407 4796 4419 4802
rect 4491 4796 4503 4802
rect 4531 4796 4543 4802
rect 4027 4704 4041 4712
rect 4033 4653 4047 4667
rect 4055 4653 4063 4716
rect 4096 4681 4104 4716
rect 4175 4701 4183 4756
rect 4267 4742 4279 4776
rect 4321 4750 4333 4756
rect 4375 4750 4383 4756
rect 4325 4738 4347 4750
rect 4375 4736 4393 4750
rect 4273 4718 4279 4736
rect 4297 4726 4327 4732
rect 4375 4730 4383 4736
rect 3899 4634 3973 4640
rect 4047 4639 4063 4653
rect 3899 4628 3906 4634
rect 3967 4632 3973 4634
rect 3931 4616 3952 4623
rect 4055 4624 4063 4639
rect 4096 4624 4104 4667
rect 4175 4638 4183 4687
rect 4159 4632 4183 4638
rect 4217 4653 4225 4716
rect 4239 4704 4253 4712
rect 4273 4712 4313 4718
rect 4233 4653 4247 4667
rect 4217 4639 4233 4653
rect 4307 4640 4313 4712
rect 4321 4712 4327 4726
rect 4345 4722 4383 4730
rect 4321 4706 4365 4712
rect 4377 4708 4439 4716
rect 4367 4667 4394 4674
rect 4414 4656 4420 4661
rect 4386 4648 4420 4656
rect 4374 4640 4381 4648
rect 4159 4624 4171 4632
rect 4217 4624 4225 4639
rect 4307 4634 4381 4640
rect 4307 4632 4313 4634
rect 3880 4604 3887 4610
rect 3945 4604 3952 4616
rect 4002 4610 4013 4618
rect 4002 4604 4009 4610
rect 3880 4598 3893 4604
rect 4374 4628 4381 4634
rect 4267 4610 4278 4618
rect 4271 4604 4278 4610
rect 4328 4616 4349 4623
rect 4433 4624 4439 4708
rect 4475 4754 4483 4756
rect 4557 4796 4569 4802
rect 4617 4796 4629 4802
rect 4711 4796 4723 4802
rect 4511 4754 4522 4756
rect 4475 4748 4522 4754
rect 4475 4693 4482 4748
rect 4476 4651 4484 4679
rect 4576 4673 4584 4756
rect 4742 4796 4754 4802
rect 4792 4796 4804 4802
rect 4636 4681 4644 4716
rect 4476 4642 4506 4651
rect 4696 4673 4704 4756
rect 4837 4796 4849 4802
rect 4917 4796 4929 4802
rect 4957 4796 4969 4802
rect 4997 4796 5009 4802
rect 5037 4796 5049 4802
rect 5091 4796 5103 4802
rect 5131 4796 5143 4802
rect 5162 4796 5174 4802
rect 5212 4796 5224 4802
rect 4773 4681 4781 4716
rect 4860 4709 4877 4716
rect 4476 4640 4494 4642
rect 4328 4604 4335 4616
rect 4393 4604 4400 4610
rect 4387 4598 4400 4604
rect 4576 4604 4584 4659
rect 4636 4624 4644 4667
rect 2520 4578 2532 4584
rect 2570 4578 2582 4584
rect 2651 4578 2663 4584
rect 2699 4578 2711 4584
rect 2757 4578 2769 4584
rect 2805 4578 2817 4584
rect 2867 4578 2879 4584
rect 2937 4578 2949 4584
rect 3039 4578 3051 4584
rect 3097 4578 3109 4584
rect 3145 4578 3157 4584
rect 3207 4578 3219 4584
rect 3279 4578 3291 4584
rect 3337 4578 3349 4584
rect 3385 4578 3397 4584
rect 3447 4578 3459 4584
rect 3551 4578 3563 4584
rect 3631 4578 3643 4584
rect 3709 4578 3721 4584
rect 3791 4578 3803 4584
rect 3861 4578 3873 4584
rect 3923 4578 3935 4584
rect 3971 4578 3983 4584
rect 4029 4578 4041 4584
rect 4111 4578 4123 4584
rect 4189 4578 4201 4584
rect 4239 4578 4251 4584
rect 4297 4578 4309 4584
rect 4345 4578 4357 4584
rect 4407 4578 4419 4584
rect 4530 4578 4542 4584
rect 4696 4604 4704 4659
rect 4779 4645 4787 4667
rect 4860 4661 4867 4709
rect 4937 4701 4945 4756
rect 4967 4717 4983 4723
rect 4780 4638 4805 4645
rect 4737 4624 4789 4627
rect 4749 4618 4777 4624
rect 4797 4624 4805 4638
rect 4860 4604 4867 4647
rect 4937 4638 4945 4687
rect 4977 4687 4983 4717
rect 5017 4701 5025 4756
rect 5047 4737 5073 4743
rect 5077 4717 5093 4723
rect 5017 4638 5025 4687
rect 5077 4683 5083 4717
rect 5115 4701 5123 4756
rect 5281 4796 5293 4802
rect 5351 4796 5363 4802
rect 5377 4796 5389 4802
rect 5417 4796 5429 4802
rect 5471 4796 5483 4802
rect 5511 4796 5523 4802
rect 5537 4796 5549 4802
rect 5577 4796 5589 4802
rect 5651 4796 5663 4802
rect 5691 4796 5703 4802
rect 5067 4677 5083 4683
rect 5115 4638 5123 4687
rect 5193 4681 5201 4716
rect 5315 4681 5323 4716
rect 5397 4701 5405 4756
rect 5427 4737 5473 4743
rect 5457 4717 5473 4723
rect 5199 4645 5207 4667
rect 5200 4638 5225 4645
rect 5316 4641 5324 4667
rect 4937 4632 4961 4638
rect 5017 4632 5041 4638
rect 4949 4624 4961 4632
rect 5029 4624 5041 4632
rect 4557 4578 4569 4584
rect 4617 4578 4629 4584
rect 4711 4578 4723 4584
rect 4757 4578 4769 4584
rect 4837 4578 4849 4584
rect 4877 4578 4889 4584
rect 5099 4632 5123 4638
rect 5099 4624 5111 4632
rect 5157 4624 5209 4627
rect 5169 4618 5197 4624
rect 5217 4624 5225 4638
rect 5295 4634 5324 4641
rect 5397 4638 5405 4687
rect 5295 4624 5301 4634
rect 5397 4632 5421 4638
rect 5457 4643 5463 4717
rect 5495 4701 5503 4756
rect 5558 4754 5569 4756
rect 5717 4796 5729 4802
rect 5757 4796 5769 4802
rect 5851 4796 5863 4802
rect 5597 4754 5605 4756
rect 5558 4748 5605 4754
rect 5447 4637 5463 4643
rect 5495 4638 5503 4687
rect 5598 4693 5605 4748
rect 5675 4701 5683 4756
rect 5738 4754 5749 4756
rect 5877 4796 5889 4802
rect 5917 4796 5929 4802
rect 6007 4796 6019 4802
rect 6051 4796 6063 4802
rect 5777 4754 5785 4756
rect 5738 4748 5785 4754
rect 5596 4651 5604 4679
rect 5311 4624 5363 4626
rect 5409 4624 5421 4632
rect 5283 4584 5311 4590
rect 5323 4620 5351 4624
rect 5479 4632 5503 4638
rect 5479 4624 5491 4632
rect 4919 4578 4931 4584
rect 4999 4578 5011 4584
rect 5129 4578 5141 4584
rect 5177 4578 5189 4584
rect 5331 4578 5343 4584
rect 5379 4578 5391 4584
rect 5509 4578 5521 4584
rect 5574 4642 5604 4651
rect 5586 4640 5604 4642
rect 5675 4638 5683 4687
rect 5778 4693 5785 4748
rect 5776 4651 5784 4679
rect 5836 4673 5844 4756
rect 5898 4754 5909 4756
rect 5937 4754 5945 4756
rect 5898 4748 5945 4754
rect 5938 4693 5945 4748
rect 6082 4796 6094 4802
rect 6132 4796 6144 4802
rect 5991 4681 5999 4716
rect 5659 4632 5683 4638
rect 5659 4624 5671 4632
rect 5538 4578 5550 4584
rect 5689 4578 5701 4584
rect 5754 4642 5784 4651
rect 5766 4640 5784 4642
rect 5836 4604 5844 4659
rect 5936 4651 5944 4679
rect 5718 4578 5730 4584
rect 5851 4578 5863 4584
rect 5914 4642 5944 4651
rect 5926 4640 5944 4642
rect 5991 4667 5993 4681
rect 5991 4624 5999 4667
rect 6034 4642 6042 4756
rect 6191 4796 6203 4802
rect 6231 4796 6243 4802
rect 6277 4796 6289 4802
rect 6357 4796 6369 4802
rect 6397 4796 6409 4802
rect 6487 4796 6499 4802
rect 6531 4796 6543 4802
rect 6591 4796 6603 4802
rect 6631 4796 6643 4802
rect 6147 4737 6163 4743
rect 6113 4681 6121 4716
rect 6157 4667 6163 4737
rect 6215 4701 6223 4756
rect 6257 4722 6269 4724
rect 6257 4716 6297 4722
rect 6378 4754 6389 4756
rect 6417 4754 6425 4756
rect 6378 4748 6425 4754
rect 6119 4645 6127 4667
rect 6025 4634 6063 4642
rect 6120 4638 6145 4645
rect 6215 4638 6223 4687
rect 6318 4681 6326 4716
rect 6418 4693 6425 4748
rect 6471 4681 6479 4716
rect 6051 4624 6063 4634
rect 5991 4614 6001 4624
rect 6077 4624 6129 4627
rect 6089 4618 6117 4624
rect 6137 4624 6145 4638
rect 6199 4632 6223 4638
rect 6199 4624 6211 4632
rect 6318 4624 6326 4667
rect 6416 4651 6424 4679
rect 5878 4578 5890 4584
rect 6021 4578 6033 4584
rect 6097 4578 6109 4584
rect 6229 4578 6241 4584
rect 6300 4613 6326 4624
rect 6260 4578 6272 4584
rect 6310 4578 6322 4584
rect 6394 4642 6424 4651
rect 6406 4640 6424 4642
rect 6471 4667 6473 4681
rect 6471 4624 6479 4667
rect 6514 4642 6522 4756
rect 6575 4754 6583 4756
rect 6611 4754 6622 4756
rect 6575 4748 6622 4754
rect 6557 4647 6563 4733
rect 6575 4693 6582 4748
rect 6647 4737 6663 4743
rect 6657 4703 6663 4737
rect 6657 4697 6673 4703
rect 6576 4651 6584 4679
rect 6505 4634 6543 4642
rect 6531 4624 6543 4634
rect 6576 4642 6606 4651
rect 6576 4640 6594 4642
rect 6471 4614 6481 4624
rect 6358 4578 6370 4584
rect 6501 4578 6513 4584
rect 6630 4578 6642 4584
rect 6742 4578 6802 5042
rect 4 4576 6802 4578
rect 6736 4564 6802 4576
rect 4 4562 6802 4564
rect 51 4556 63 4562
rect 91 4556 103 4562
rect 131 4556 143 4562
rect 191 4556 203 4562
rect 237 4556 249 4562
rect 331 4556 343 4562
rect 371 4556 383 4562
rect 417 4556 429 4562
rect 497 4556 505 4562
rect 537 4556 549 4562
rect 600 4556 612 4562
rect 650 4556 662 4562
rect 731 4556 743 4562
rect 36 4481 44 4536
rect 113 4493 120 4536
rect 176 4481 184 4536
rect 229 4516 257 4522
rect 217 4513 269 4516
rect 277 4502 285 4516
rect 260 4495 285 4502
rect 36 4384 44 4467
rect 113 4431 120 4479
rect 103 4424 120 4431
rect 176 4384 184 4467
rect 259 4473 267 4495
rect 353 4493 360 4536
rect 409 4516 437 4522
rect 397 4513 449 4516
rect 457 4502 465 4516
rect 523 4508 529 4536
rect 757 4556 769 4562
rect 797 4556 809 4562
rect 837 4556 849 4562
rect 897 4556 909 4562
rect 937 4556 949 4562
rect 977 4556 989 4562
rect 1037 4556 1049 4562
rect 1077 4556 1089 4562
rect 1117 4556 1129 4562
rect 1157 4556 1169 4562
rect 1197 4556 1209 4562
rect 1259 4556 1271 4562
rect 1351 4556 1363 4562
rect 640 4516 666 4527
rect 523 4502 533 4508
rect 440 4495 465 4502
rect 253 4424 261 4459
rect 353 4431 360 4479
rect 439 4473 447 4495
rect 343 4424 360 4431
rect 433 4424 441 4459
rect 538 4441 544 4496
rect 560 4481 567 4516
rect 658 4473 666 4516
rect 716 4481 724 4536
rect 780 4493 787 4536
rect 497 4432 533 4440
rect 497 4424 505 4432
rect 51 4338 63 4344
rect 131 4338 143 4344
rect 191 4338 203 4344
rect 222 4338 234 4344
rect 272 4338 284 4344
rect 371 4338 383 4344
rect 554 4423 563 4467
rect 856 4481 864 4536
rect 920 4493 927 4536
rect 658 4424 666 4459
rect 559 4414 563 4423
rect 597 4418 637 4424
rect 597 4416 609 4418
rect 716 4384 724 4467
rect 780 4431 787 4479
rect 996 4481 1004 4536
rect 1056 4510 1068 4516
rect 1097 4510 1109 4516
rect 1136 4510 1148 4516
rect 1176 4510 1188 4516
rect 1241 4510 1249 4536
rect 1391 4556 1403 4562
rect 1431 4556 1443 4562
rect 1509 4556 1521 4562
rect 1056 4502 1083 4510
rect 1097 4502 1122 4510
rect 1136 4502 1162 4510
rect 1176 4509 1194 4510
rect 1176 4502 1195 4509
rect 1241 4504 1263 4510
rect 1075 4496 1083 4502
rect 1114 4496 1122 4502
rect 1154 4496 1162 4502
rect 1075 4484 1090 4496
rect 1114 4484 1130 4496
rect 1154 4484 1170 4496
rect 780 4424 797 4431
rect 402 4338 414 4344
rect 452 4338 464 4344
rect 527 4338 539 4344
rect 617 4338 629 4344
rect 731 4338 743 4344
rect 856 4384 864 4467
rect 920 4431 927 4479
rect 920 4424 937 4431
rect 996 4384 1004 4467
rect 1075 4438 1083 4484
rect 1114 4438 1122 4484
rect 1154 4438 1162 4484
rect 1188 4481 1195 4502
rect 1260 4498 1263 4504
rect 1188 4467 1193 4481
rect 1188 4438 1195 4467
rect 1057 4430 1083 4438
rect 1097 4430 1122 4438
rect 1137 4430 1162 4438
rect 1177 4430 1195 4438
rect 1260 4442 1267 4498
rect 1281 4473 1289 4516
rect 1336 4481 1344 4536
rect 1377 4497 1393 4503
rect 1287 4459 1289 4473
rect 1260 4436 1263 4442
rect 1237 4430 1263 4436
rect 1057 4424 1069 4430
rect 1097 4424 1109 4430
rect 1137 4424 1149 4430
rect 1177 4424 1189 4430
rect 1237 4384 1245 4430
rect 1281 4424 1289 4459
rect 1336 4384 1344 4467
rect 1377 4443 1383 4497
rect 1413 4493 1420 4536
rect 1539 4556 1551 4562
rect 1631 4556 1643 4562
rect 1671 4556 1683 4562
rect 1711 4556 1723 4562
rect 1761 4556 1773 4562
rect 1823 4556 1835 4562
rect 1871 4556 1883 4562
rect 1929 4556 1941 4562
rect 1979 4556 1991 4562
rect 2079 4556 2091 4562
rect 2137 4556 2149 4562
rect 2185 4556 2197 4562
rect 2247 4556 2259 4562
rect 2297 4556 2309 4562
rect 2357 4556 2369 4562
rect 2397 4556 2409 4562
rect 1780 4536 1793 4542
rect 1780 4530 1787 4536
rect 1845 4524 1852 4536
rect 1479 4508 1491 4516
rect 1569 4508 1581 4516
rect 1447 4497 1463 4503
rect 1479 4502 1503 4508
rect 1367 4437 1383 4443
rect 1413 4431 1420 4479
rect 1403 4424 1420 4431
rect 1457 4423 1463 4497
rect 1495 4453 1503 4502
rect 1557 4502 1581 4508
rect 1655 4510 1663 4516
rect 1695 4510 1703 4516
rect 1655 4502 1703 4510
rect 1557 4453 1565 4502
rect 1655 4473 1663 4502
rect 1457 4417 1473 4423
rect 1495 4384 1503 4439
rect 1557 4384 1565 4439
rect 1655 4436 1663 4459
rect 1655 4430 1703 4436
rect 1655 4424 1663 4430
rect 1691 4424 1703 4430
rect 1741 4432 1747 4516
rect 1831 4517 1852 4524
rect 1902 4530 1909 4536
rect 1902 4522 1913 4530
rect 1799 4506 1806 4512
rect 1867 4506 1873 4508
rect 1799 4500 1873 4506
rect 1955 4501 1963 4516
rect 2009 4508 2021 4516
rect 1799 4492 1806 4500
rect 1760 4484 1794 4492
rect 1760 4479 1766 4484
rect 1786 4466 1813 4473
rect 1741 4424 1803 4432
rect 1815 4428 1859 4434
rect 757 4338 769 4344
rect 837 4338 849 4344
rect 897 4338 909 4344
rect 977 4338 989 4344
rect 1037 4338 1049 4344
rect 1077 4338 1089 4344
rect 1117 4338 1129 4344
rect 1157 4338 1169 4344
rect 1197 4338 1209 4344
rect 1259 4338 1271 4344
rect 1351 4338 1363 4344
rect 1431 4338 1443 4344
rect 1471 4338 1483 4344
rect 1511 4338 1523 4344
rect 1537 4338 1549 4344
rect 1577 4338 1589 4344
rect 1797 4410 1835 4418
rect 1853 4414 1859 4428
rect 1867 4428 1873 4500
rect 1947 4487 1963 4501
rect 1933 4473 1947 4487
rect 1867 4422 1907 4428
rect 1927 4428 1941 4436
rect 1955 4424 1963 4487
rect 1997 4502 2021 4508
rect 2227 4536 2240 4542
rect 2111 4530 2118 4536
rect 2107 4522 2118 4530
rect 2168 4524 2175 4536
rect 2233 4530 2240 4536
rect 1997 4453 2005 4502
rect 2057 4501 2065 4516
rect 2168 4517 2189 4524
rect 2437 4556 2449 4562
rect 2477 4556 2489 4562
rect 2517 4556 2529 4562
rect 2599 4556 2611 4562
rect 2657 4556 2669 4562
rect 2705 4556 2717 4562
rect 2767 4556 2779 4562
rect 2837 4556 2849 4562
rect 2919 4556 2931 4562
rect 3031 4556 3043 4562
rect 3077 4556 3089 4562
rect 3179 4556 3191 4562
rect 3237 4556 3249 4562
rect 3285 4556 3297 4562
rect 3347 4556 3359 4562
rect 3417 4556 3429 4562
rect 3551 4556 3563 4562
rect 3621 4556 3633 4562
rect 3683 4556 3695 4562
rect 3731 4556 3743 4562
rect 3789 4556 3801 4562
rect 3857 4556 3869 4562
rect 3961 4556 3973 4562
rect 4023 4556 4035 4562
rect 4071 4556 4083 4562
rect 4129 4556 4141 4562
rect 4250 4556 4262 4562
rect 4297 4556 4309 4562
rect 4391 4556 4403 4562
rect 4431 4556 4443 4562
rect 2147 4506 2153 4508
rect 2214 4506 2221 4512
rect 2057 4487 2073 4501
rect 2147 4500 2221 4506
rect 1797 4404 1805 4410
rect 1853 4408 1883 4414
rect 1901 4404 1907 4422
rect 1787 4390 1805 4404
rect 1833 4390 1855 4402
rect 1797 4384 1805 4390
rect 1847 4384 1859 4390
rect 1901 4364 1913 4398
rect 1997 4384 2005 4439
rect 2057 4424 2065 4487
rect 2073 4473 2087 4487
rect 2079 4428 2093 4436
rect 2147 4428 2153 4500
rect 2214 4492 2221 4500
rect 2226 4484 2260 4492
rect 2254 4479 2260 4484
rect 2207 4466 2234 4473
rect 2113 4422 2153 4428
rect 2161 4428 2205 4434
rect 2113 4404 2119 4422
rect 2161 4414 2167 4428
rect 2273 4432 2279 4516
rect 2316 4481 2324 4536
rect 2380 4493 2387 4536
rect 2460 4493 2467 4536
rect 2536 4481 2544 4536
rect 2747 4536 2760 4542
rect 2631 4530 2638 4536
rect 2627 4522 2638 4530
rect 2688 4524 2695 4536
rect 2753 4530 2760 4536
rect 2577 4501 2585 4516
rect 2688 4517 2709 4524
rect 2667 4506 2673 4508
rect 2734 4506 2741 4512
rect 2577 4487 2593 4501
rect 2667 4500 2741 4506
rect 2217 4424 2279 4432
rect 2137 4408 2167 4414
rect 2185 4410 2223 4418
rect 2215 4404 2223 4410
rect 2107 4364 2119 4398
rect 2165 4390 2187 4402
rect 2215 4390 2233 4404
rect 2161 4384 2173 4390
rect 2215 4384 2223 4390
rect 2316 4384 2324 4467
rect 2380 4431 2387 4479
rect 2460 4431 2467 4479
rect 2380 4424 2397 4431
rect 2460 4424 2477 4431
rect 2536 4384 2544 4467
rect 2577 4424 2585 4487
rect 2593 4473 2607 4487
rect 2599 4428 2613 4436
rect 2667 4428 2673 4500
rect 2734 4492 2741 4500
rect 2746 4484 2780 4492
rect 2774 4479 2780 4484
rect 2727 4466 2754 4473
rect 2633 4422 2673 4428
rect 2681 4428 2725 4434
rect 2633 4404 2639 4422
rect 2681 4414 2687 4428
rect 2793 4432 2799 4516
rect 2829 4516 2857 4522
rect 2817 4513 2869 4516
rect 2877 4502 2885 4516
rect 2949 4508 2961 4516
rect 2860 4495 2885 4502
rect 2937 4502 2961 4508
rect 2859 4473 2867 4495
rect 2737 4424 2799 4432
rect 2853 4424 2861 4459
rect 2937 4453 2945 4502
rect 3016 4481 3024 4536
rect 3069 4516 3097 4522
rect 3057 4513 3109 4516
rect 3327 4536 3340 4542
rect 3211 4530 3218 4536
rect 3207 4522 3218 4530
rect 3268 4524 3275 4536
rect 3333 4530 3340 4536
rect 3117 4502 3125 4516
rect 3100 4495 3125 4502
rect 3157 4501 3165 4516
rect 3268 4517 3289 4524
rect 3247 4506 3253 4508
rect 3314 4506 3321 4512
rect 2657 4408 2687 4414
rect 2705 4410 2743 4418
rect 2735 4404 2743 4410
rect 2627 4364 2639 4398
rect 2685 4390 2707 4402
rect 2735 4390 2753 4404
rect 2681 4384 2693 4390
rect 2735 4384 2743 4390
rect 2937 4384 2945 4439
rect 3016 4384 3024 4467
rect 3099 4473 3107 4495
rect 3157 4487 3173 4501
rect 3247 4500 3321 4506
rect 3093 4424 3101 4459
rect 3157 4424 3165 4487
rect 3173 4473 3187 4487
rect 3179 4428 3193 4436
rect 1631 4338 1643 4344
rect 1671 4338 1683 4344
rect 1711 4338 1723 4344
rect 1761 4338 1773 4344
rect 1827 4338 1839 4344
rect 1873 4338 1885 4344
rect 1931 4338 1943 4344
rect 1977 4338 1989 4344
rect 2017 4338 2029 4344
rect 2077 4338 2089 4344
rect 2135 4338 2147 4344
rect 2181 4338 2193 4344
rect 2247 4338 2259 4344
rect 2297 4338 2309 4344
rect 2357 4338 2369 4344
rect 2437 4338 2449 4344
rect 2517 4338 2529 4344
rect 2597 4338 2609 4344
rect 2655 4338 2667 4344
rect 2701 4338 2713 4344
rect 2767 4338 2779 4344
rect 2822 4338 2834 4344
rect 2872 4338 2884 4344
rect 2917 4338 2929 4344
rect 2957 4338 2969 4344
rect 3031 4338 3043 4344
rect 3247 4428 3253 4500
rect 3314 4492 3321 4500
rect 3326 4484 3360 4492
rect 3354 4479 3360 4484
rect 3307 4466 3334 4473
rect 3213 4422 3253 4428
rect 3261 4428 3305 4434
rect 3213 4404 3219 4422
rect 3261 4414 3267 4428
rect 3373 4432 3379 4516
rect 3409 4516 3437 4522
rect 3397 4513 3449 4516
rect 3457 4502 3465 4516
rect 3440 4495 3465 4502
rect 3515 4502 3523 4516
rect 3543 4516 3571 4522
rect 3531 4513 3583 4516
rect 3640 4536 3653 4542
rect 3640 4530 3647 4536
rect 3705 4524 3712 4536
rect 3515 4495 3540 4502
rect 3439 4473 3447 4495
rect 3497 4477 3513 4483
rect 3317 4424 3379 4432
rect 3433 4424 3441 4459
rect 3237 4408 3267 4414
rect 3285 4410 3323 4418
rect 3315 4404 3323 4410
rect 3207 4364 3219 4398
rect 3265 4390 3287 4402
rect 3315 4390 3333 4404
rect 3261 4384 3273 4390
rect 3315 4384 3323 4390
rect 3497 4403 3503 4477
rect 3533 4473 3541 4495
rect 3539 4424 3547 4459
rect 3601 4432 3607 4516
rect 3691 4517 3712 4524
rect 3762 4530 3769 4536
rect 3762 4522 3773 4530
rect 3659 4506 3666 4512
rect 3727 4506 3733 4508
rect 3659 4500 3733 4506
rect 3815 4501 3823 4516
rect 3849 4516 3877 4522
rect 3837 4513 3889 4516
rect 3980 4536 3993 4542
rect 3980 4530 3987 4536
rect 4045 4524 4052 4536
rect 3897 4502 3905 4516
rect 3659 4492 3666 4500
rect 3620 4484 3654 4492
rect 3620 4479 3626 4484
rect 3646 4466 3673 4473
rect 3601 4424 3663 4432
rect 3675 4428 3719 4434
rect 3497 4397 3513 4403
rect 3062 4338 3074 4344
rect 3112 4338 3124 4344
rect 3177 4338 3189 4344
rect 3235 4338 3247 4344
rect 3281 4338 3293 4344
rect 3347 4338 3359 4344
rect 3402 4338 3414 4344
rect 3452 4338 3464 4344
rect -62 4336 3493 4338
rect 3657 4410 3695 4418
rect 3713 4414 3719 4428
rect 3727 4428 3733 4500
rect 3807 4487 3823 4501
rect 3880 4495 3905 4502
rect 3793 4473 3807 4487
rect 3727 4422 3767 4428
rect 3787 4428 3801 4436
rect 3815 4424 3823 4487
rect 3879 4473 3887 4495
rect 3873 4424 3881 4459
rect 3941 4432 3947 4516
rect 4031 4517 4052 4524
rect 4102 4530 4109 4536
rect 4102 4522 4113 4530
rect 3999 4506 4006 4512
rect 4067 4506 4073 4508
rect 3999 4500 4073 4506
rect 4155 4501 4163 4516
rect 3999 4492 4006 4500
rect 3960 4484 3994 4492
rect 3960 4479 3966 4484
rect 3986 4466 4013 4473
rect 3941 4424 4003 4432
rect 4015 4428 4059 4434
rect 3657 4404 3665 4410
rect 3713 4408 3743 4414
rect 3761 4404 3767 4422
rect 3647 4390 3665 4404
rect 3693 4390 3715 4402
rect 3657 4384 3665 4390
rect 3707 4384 3719 4390
rect 3761 4364 3773 4398
rect 3997 4410 4035 4418
rect 4053 4414 4059 4428
rect 4067 4428 4073 4500
rect 4147 4487 4163 4501
rect 4133 4473 4147 4487
rect 4067 4422 4107 4428
rect 4127 4428 4141 4436
rect 4155 4424 4163 4487
rect 4196 4498 4214 4500
rect 4196 4489 4226 4498
rect 4289 4516 4317 4522
rect 4277 4513 4329 4516
rect 4478 4556 4490 4562
rect 4528 4556 4540 4562
rect 4337 4502 4345 4516
rect 4320 4495 4345 4502
rect 4196 4461 4204 4489
rect 4319 4473 4327 4495
rect 4413 4493 4420 4536
rect 4474 4516 4500 4527
rect 4558 4556 4570 4562
rect 4691 4556 4703 4562
rect 4737 4556 4749 4562
rect 4851 4556 4863 4562
rect 4895 4556 4903 4562
rect 4969 4556 4981 4562
rect 5070 4556 5082 4562
rect 5117 4556 5129 4562
rect 5231 4556 5243 4562
rect 5275 4556 5283 4562
rect 5317 4556 5329 4562
rect 5397 4556 5409 4562
rect 5530 4556 5542 4562
rect 3997 4404 4005 4410
rect 4053 4408 4083 4414
rect 4101 4404 4107 4422
rect 3987 4390 4005 4404
rect 4033 4390 4055 4402
rect 3997 4384 4005 4390
rect 4047 4384 4059 4390
rect 4101 4364 4113 4398
rect 4195 4392 4202 4447
rect 4313 4424 4321 4459
rect 4413 4431 4420 4479
rect 4474 4473 4482 4516
rect 4606 4498 4624 4500
rect 4594 4489 4624 4498
rect 4616 4461 4624 4489
rect 4676 4481 4684 4536
rect 4729 4516 4757 4522
rect 4717 4513 4769 4516
rect 4777 4502 4785 4516
rect 4760 4495 4785 4502
rect 4403 4424 4420 4431
rect 4474 4424 4482 4459
rect 4195 4386 4242 4392
rect 4195 4384 4203 4386
rect 4231 4384 4242 4386
rect 3516 4338 3528 4344
rect 3566 4338 3578 4344
rect 3621 4338 3633 4344
rect 3687 4338 3699 4344
rect 3733 4338 3745 4344
rect 3791 4338 3803 4344
rect 3842 4338 3854 4344
rect 3892 4338 3904 4344
rect 3961 4338 3973 4344
rect 4027 4338 4039 4344
rect 4073 4338 4085 4344
rect 4131 4338 4143 4344
rect 4211 4338 4223 4344
rect 4251 4338 4263 4344
rect 4282 4338 4294 4344
rect 4332 4338 4344 4344
rect 3507 4336 4373 4338
rect 4503 4418 4543 4424
rect 4531 4416 4543 4418
rect 4618 4392 4625 4447
rect 4578 4386 4625 4392
rect 4578 4384 4589 4386
rect 4617 4384 4625 4386
rect 4676 4384 4684 4467
rect 4759 4473 4767 4495
rect 4833 4481 4840 4516
rect 4871 4508 4877 4536
rect 4867 4502 4877 4508
rect 4939 4508 4951 4516
rect 4939 4502 4963 4508
rect 4753 4424 4761 4459
rect 4431 4338 4443 4344
rect 4511 4338 4523 4344
rect 4557 4338 4569 4344
rect 4597 4338 4609 4344
rect 4691 4338 4703 4344
rect 4837 4423 4846 4467
rect 4856 4441 4862 4496
rect 4955 4453 4963 4502
rect 5016 4498 5034 4500
rect 5016 4489 5046 4498
rect 5109 4516 5137 4522
rect 5097 4513 5149 4516
rect 5157 4502 5165 4516
rect 5140 4495 5165 4502
rect 5016 4461 5024 4489
rect 4867 4432 4903 4440
rect 5139 4473 5147 4495
rect 5213 4481 5220 4516
rect 5251 4508 5257 4536
rect 5309 4516 5337 4522
rect 5297 4513 5349 4516
rect 5247 4502 5257 4508
rect 5357 4502 5365 4516
rect 4895 4424 4903 4432
rect 4837 4414 4841 4423
rect 4955 4384 4963 4439
rect 5015 4392 5022 4447
rect 5133 4424 5141 4459
rect 5015 4386 5062 4392
rect 5015 4384 5023 4386
rect 5051 4384 5062 4386
rect 4722 4338 4734 4344
rect 4772 4338 4784 4344
rect 4861 4338 4873 4344
rect 4931 4338 4943 4344
rect 4971 4338 4983 4344
rect 5031 4338 5043 4344
rect 5071 4338 5083 4344
rect 5217 4423 5226 4467
rect 5236 4441 5242 4496
rect 5340 4495 5365 4502
rect 5339 4473 5347 4495
rect 5367 4477 5383 4483
rect 5416 4481 5424 4536
rect 5247 4432 5283 4440
rect 5275 4424 5283 4432
rect 5333 4424 5341 4459
rect 5377 4427 5383 4477
rect 5217 4414 5221 4423
rect 5416 4384 5424 4467
rect 5457 4407 5463 4533
rect 5476 4498 5494 4500
rect 5476 4489 5506 4498
rect 5559 4556 5571 4562
rect 5657 4556 5669 4562
rect 5789 4556 5801 4562
rect 5890 4556 5902 4562
rect 5971 4556 5983 4562
rect 6017 4556 6029 4562
rect 6111 4556 6123 4562
rect 5589 4508 5601 4516
rect 5649 4516 5677 4522
rect 5637 4513 5689 4516
rect 5577 4502 5601 4508
rect 5476 4461 5484 4489
rect 5475 4392 5482 4447
rect 5577 4453 5585 4502
rect 5617 4497 5633 4503
rect 5475 4386 5522 4392
rect 5475 4384 5483 4386
rect 5102 4338 5114 4344
rect 5152 4338 5164 4344
rect 5241 4338 5253 4344
rect 5302 4338 5314 4344
rect 5352 4338 5364 4344
rect 5511 4384 5522 4386
rect 5577 4384 5585 4439
rect 5617 4427 5623 4497
rect 5697 4502 5705 4516
rect 5759 4508 5771 4516
rect 5759 4502 5783 4508
rect 5680 4495 5705 4502
rect 5679 4473 5687 4495
rect 5707 4477 5723 4483
rect 5673 4424 5681 4459
rect 5397 4338 5409 4344
rect 5491 4338 5503 4344
rect 5531 4338 5543 4344
rect 5557 4338 5569 4344
rect 5597 4338 5609 4344
rect 5717 4423 5723 4477
rect 5775 4453 5783 4502
rect 5836 4498 5854 4500
rect 5836 4489 5866 4498
rect 5935 4502 5943 4516
rect 5963 4516 5991 4522
rect 6138 4556 6150 4562
rect 6291 4556 6303 4562
rect 6338 4556 6350 4562
rect 6438 4556 6450 4562
rect 6557 4556 6569 4562
rect 6637 4556 6649 4562
rect 5951 4513 6003 4516
rect 5935 4495 5960 4502
rect 5836 4461 5844 4489
rect 5887 4477 5923 4483
rect 5717 4417 5753 4423
rect 5775 4384 5783 4439
rect 5835 4392 5842 4447
rect 5917 4447 5923 4477
rect 5953 4473 5961 4495
rect 6036 4481 6044 4536
rect 6096 4481 6104 4536
rect 6255 4502 6263 4516
rect 6283 4516 6311 4522
rect 6271 4513 6323 4516
rect 6186 4498 6204 4500
rect 6174 4489 6204 4498
rect 6255 4495 6280 4502
rect 6386 4498 6404 4500
rect 5959 4424 5967 4459
rect 5835 4386 5882 4392
rect 5835 4384 5843 4386
rect 5642 4338 5654 4344
rect 5692 4338 5704 4344
rect 5871 4384 5882 4386
rect 5751 4338 5763 4344
rect 5791 4338 5803 4344
rect 5851 4338 5863 4344
rect 5891 4338 5903 4344
rect 6036 4384 6044 4467
rect 6096 4384 6104 4467
rect 6196 4461 6204 4489
rect 6273 4473 6281 4495
rect 6374 4489 6404 4498
rect 6549 4516 6577 4522
rect 6537 4513 6589 4516
rect 6597 4502 6605 4516
rect 6486 4498 6504 4500
rect 6474 4489 6504 4498
rect 6580 4495 6605 4502
rect 6396 4461 6404 4489
rect 6417 4477 6433 4483
rect 6198 4392 6205 4447
rect 6279 4424 6287 4459
rect 6158 4386 6205 4392
rect 6158 4384 6169 4386
rect 5936 4338 5948 4344
rect 5986 4338 5998 4344
rect 6017 4338 6029 4344
rect 6111 4338 6123 4344
rect 6197 4384 6205 4386
rect 6398 4392 6405 4447
rect 6417 4403 6423 4477
rect 6496 4461 6504 4489
rect 6579 4473 6587 4495
rect 6656 4481 6664 4536
rect 6417 4397 6433 4403
rect 6498 4392 6505 4447
rect 6573 4424 6581 4459
rect 6358 4386 6405 4392
rect 6358 4384 6369 4386
rect 6137 4338 6149 4344
rect 6177 4338 6189 4344
rect 6256 4338 6268 4344
rect 6306 4338 6318 4344
rect 6397 4384 6405 4386
rect 6458 4386 6505 4392
rect 6458 4384 6469 4386
rect 6497 4384 6505 4386
rect 6656 4384 6664 4467
rect 6337 4338 6349 4344
rect 6377 4338 6389 4344
rect 6437 4338 6449 4344
rect 6477 4338 6489 4344
rect 6542 4338 6554 4344
rect 6592 4338 6604 4344
rect 6637 4338 6649 4344
rect 4387 4336 6736 4338
rect -62 4324 4 4336
rect -62 4322 93 4324
rect -62 3858 -2 4322
rect 49 4316 61 4322
rect 107 4322 2733 4324
rect 116 4316 128 4322
rect 166 4316 178 4322
rect 31 4201 39 4236
rect 75 4230 83 4276
rect 202 4316 214 4322
rect 252 4316 264 4322
rect 321 4316 333 4322
rect 387 4316 399 4322
rect 433 4316 445 4322
rect 491 4316 503 4322
rect 537 4316 549 4322
rect 577 4316 589 4322
rect 691 4316 703 4322
rect 771 4316 783 4322
rect 817 4316 829 4322
rect 875 4316 887 4322
rect 921 4316 933 4322
rect 987 4316 999 4322
rect 1037 4316 1049 4322
rect 1077 4316 1089 4322
rect 1137 4316 1149 4322
rect 1195 4316 1207 4322
rect 1241 4316 1253 4322
rect 1307 4316 1319 4322
rect 1357 4316 1369 4322
rect 1397 4316 1409 4322
rect 357 4270 365 4276
rect 407 4270 419 4276
rect 347 4256 365 4270
rect 393 4258 415 4270
rect 461 4262 473 4296
rect 357 4250 365 4256
rect 357 4242 395 4250
rect 413 4246 443 4252
rect 57 4224 83 4230
rect 57 4218 60 4224
rect 31 4187 33 4201
rect 31 4144 39 4187
rect 53 4162 60 4218
rect 139 4201 147 4236
rect 233 4201 241 4236
rect 301 4228 363 4236
rect 133 4165 141 4187
rect 239 4165 247 4187
rect 57 4156 60 4162
rect 115 4158 140 4165
rect 240 4158 265 4165
rect 57 4150 79 4156
rect 71 4124 79 4150
rect 115 4144 123 4158
rect 131 4144 183 4147
rect 143 4138 171 4144
rect 197 4144 249 4147
rect 209 4138 237 4144
rect 257 4144 265 4158
rect 301 4144 307 4228
rect 413 4232 419 4246
rect 461 4238 467 4256
rect 375 4226 419 4232
rect 427 4232 467 4238
rect 346 4187 373 4194
rect 320 4176 326 4181
rect 320 4168 354 4176
rect 359 4160 366 4168
rect 427 4160 433 4232
rect 487 4224 501 4232
rect 493 4173 507 4187
rect 515 4173 523 4236
rect 557 4221 565 4276
rect 597 4223 603 4253
rect 643 4310 671 4316
rect 683 4238 711 4244
rect 652 4230 664 4236
rect 652 4224 679 4230
rect 597 4217 623 4223
rect 359 4154 433 4160
rect 507 4159 523 4173
rect 359 4148 366 4154
rect 427 4152 433 4154
rect 391 4136 412 4143
rect 515 4144 523 4159
rect 557 4158 565 4207
rect 617 4163 623 4217
rect 673 4201 679 4224
rect 557 4152 581 4158
rect 617 4157 633 4163
rect 569 4144 581 4152
rect 680 4144 687 4187
rect 737 4167 743 4213
rect 756 4193 764 4276
rect 847 4262 859 4296
rect 901 4270 913 4276
rect 955 4270 963 4276
rect 905 4258 927 4270
rect 955 4256 973 4270
rect 853 4238 859 4256
rect 877 4246 907 4252
rect 955 4250 963 4256
rect 340 4124 347 4130
rect 405 4124 412 4136
rect 462 4130 473 4138
rect 462 4124 469 4130
rect 340 4118 353 4124
rect 756 4124 764 4179
rect 797 4173 805 4236
rect 819 4224 833 4232
rect 853 4232 893 4238
rect 813 4173 827 4187
rect 797 4159 813 4173
rect 887 4160 893 4232
rect 901 4232 907 4246
rect 925 4242 963 4250
rect 901 4226 945 4232
rect 957 4228 1019 4236
rect 947 4187 974 4194
rect 994 4176 1000 4181
rect 966 4168 1000 4176
rect 954 4160 961 4168
rect 797 4144 805 4159
rect 887 4154 961 4160
rect 887 4152 893 4154
rect 954 4148 961 4154
rect 847 4130 858 4138
rect 851 4124 858 4130
rect 908 4136 929 4143
rect 1013 4144 1019 4228
rect 1057 4221 1065 4276
rect 1167 4262 1179 4296
rect 1221 4270 1233 4276
rect 1275 4270 1283 4276
rect 1225 4258 1247 4270
rect 1275 4256 1293 4270
rect 1173 4238 1179 4256
rect 1197 4246 1227 4252
rect 1275 4250 1283 4256
rect 1057 4158 1065 4207
rect 1117 4173 1125 4236
rect 1139 4224 1153 4232
rect 1173 4232 1213 4238
rect 1133 4173 1147 4187
rect 1117 4159 1133 4173
rect 1207 4160 1213 4232
rect 1221 4232 1227 4246
rect 1245 4242 1283 4250
rect 1437 4316 1449 4322
rect 1516 4316 1528 4322
rect 1566 4316 1578 4322
rect 1651 4316 1663 4322
rect 1711 4316 1723 4322
rect 1751 4316 1763 4322
rect 1221 4226 1265 4232
rect 1277 4228 1339 4236
rect 1267 4187 1294 4194
rect 1314 4176 1320 4181
rect 1286 4168 1320 4176
rect 1274 4160 1281 4168
rect 1057 4152 1081 4158
rect 1069 4144 1081 4152
rect 908 4124 915 4136
rect 973 4124 980 4130
rect 967 4118 980 4124
rect 1117 4144 1125 4159
rect 1207 4154 1281 4160
rect 1207 4152 1213 4154
rect 1274 4148 1281 4154
rect 1167 4130 1178 4138
rect 1171 4124 1178 4130
rect 1228 4136 1249 4143
rect 1333 4144 1339 4228
rect 1377 4221 1385 4276
rect 1377 4158 1385 4207
rect 1456 4193 1464 4276
rect 1777 4316 1789 4322
rect 1817 4316 1829 4322
rect 1877 4316 1889 4322
rect 1935 4316 1947 4322
rect 1981 4316 1993 4322
rect 2047 4316 2059 4322
rect 2097 4316 2109 4322
rect 2137 4316 2149 4322
rect 1671 4242 1683 4244
rect 1643 4236 1683 4242
rect 1539 4201 1547 4236
rect 1614 4201 1622 4236
rect 1735 4221 1743 4276
rect 1797 4221 1805 4276
rect 1907 4262 1919 4296
rect 1961 4270 1973 4276
rect 2015 4270 2023 4276
rect 1965 4258 1987 4270
rect 2015 4256 2033 4270
rect 1913 4238 1919 4256
rect 1937 4246 1967 4252
rect 2015 4250 2023 4256
rect 1377 4152 1401 4158
rect 1389 4144 1401 4152
rect 1228 4124 1235 4136
rect 1293 4124 1300 4130
rect 1287 4118 1300 4124
rect 1456 4124 1464 4179
rect 1533 4165 1541 4187
rect 1515 4158 1540 4165
rect 1515 4144 1523 4158
rect 1531 4144 1583 4147
rect 1543 4138 1571 4144
rect 1614 4144 1622 4187
rect 1735 4158 1743 4207
rect 1719 4152 1743 4158
rect 1797 4158 1805 4207
rect 1857 4173 1865 4236
rect 1879 4224 1893 4232
rect 1913 4232 1953 4238
rect 1873 4173 1887 4187
rect 1857 4159 1873 4173
rect 1947 4160 1953 4232
rect 1961 4232 1967 4246
rect 1985 4242 2023 4250
rect 2196 4316 2208 4322
rect 2246 4316 2258 4322
rect 2301 4316 2313 4322
rect 2367 4316 2379 4322
rect 2413 4316 2425 4322
rect 2471 4316 2483 4322
rect 2571 4316 2583 4322
rect 1961 4226 2005 4232
rect 2017 4228 2079 4236
rect 2007 4187 2034 4194
rect 2054 4176 2060 4181
rect 2026 4168 2060 4176
rect 2014 4160 2021 4168
rect 1797 4152 1821 4158
rect 1719 4144 1731 4152
rect 1809 4144 1821 4152
rect 1614 4133 1640 4144
rect 49 4098 61 4104
rect 151 4098 163 4104
rect 217 4098 229 4104
rect 321 4098 333 4104
rect 383 4098 395 4104
rect 431 4098 443 4104
rect 489 4098 501 4104
rect 539 4098 551 4104
rect 652 4098 664 4104
rect 708 4098 720 4104
rect 771 4098 783 4104
rect 819 4098 831 4104
rect 877 4098 889 4104
rect 925 4098 937 4104
rect 987 4098 999 4104
rect 1039 4098 1051 4104
rect 1139 4098 1151 4104
rect 1197 4098 1209 4104
rect 1245 4098 1257 4104
rect 1307 4098 1319 4104
rect 1359 4098 1371 4104
rect 1437 4098 1449 4104
rect 1551 4098 1563 4104
rect 1618 4098 1630 4104
rect 1668 4098 1680 4104
rect 1749 4098 1761 4104
rect 1857 4144 1865 4159
rect 1947 4154 2021 4160
rect 1947 4152 1953 4154
rect 2014 4148 2021 4154
rect 1907 4130 1918 4138
rect 1911 4124 1918 4130
rect 1968 4136 1989 4143
rect 2073 4144 2079 4228
rect 2117 4221 2125 4276
rect 2337 4270 2345 4276
rect 2387 4270 2399 4276
rect 2327 4256 2345 4270
rect 2373 4258 2395 4270
rect 2441 4262 2453 4296
rect 2337 4250 2345 4256
rect 2337 4242 2375 4250
rect 2393 4246 2423 4252
rect 2117 4158 2125 4207
rect 2219 4201 2227 4236
rect 2281 4228 2343 4236
rect 2213 4165 2221 4187
rect 2195 4158 2220 4165
rect 2117 4152 2141 4158
rect 2129 4144 2141 4152
rect 2195 4144 2203 4158
rect 1968 4124 1975 4136
rect 2033 4124 2040 4130
rect 2027 4118 2040 4124
rect 2211 4144 2263 4147
rect 2223 4138 2251 4144
rect 2281 4144 2287 4228
rect 2393 4232 2399 4246
rect 2441 4238 2447 4256
rect 2355 4226 2399 4232
rect 2407 4232 2447 4238
rect 2326 4187 2353 4194
rect 2300 4176 2306 4181
rect 2300 4168 2334 4176
rect 2339 4160 2346 4168
rect 2407 4160 2413 4232
rect 2467 4224 2481 4232
rect 2473 4173 2487 4187
rect 2495 4173 2503 4236
rect 2597 4316 2609 4322
rect 2662 4316 2674 4322
rect 2712 4316 2724 4322
rect 2543 4229 2560 4236
rect 2339 4154 2413 4160
rect 2487 4159 2503 4173
rect 2339 4148 2346 4154
rect 2407 4152 2413 4154
rect 2371 4136 2392 4143
rect 2495 4144 2503 4159
rect 2320 4124 2327 4130
rect 2385 4124 2392 4136
rect 2442 4130 2453 4138
rect 2442 4124 2449 4130
rect 2320 4118 2333 4124
rect 2553 4181 2560 4229
rect 2616 4193 2624 4276
rect 2747 4322 2833 4324
rect 2757 4316 2769 4322
rect 2797 4316 2809 4322
rect 2847 4322 3053 4324
rect 2856 4316 2868 4322
rect 2906 4316 2918 4322
rect 2693 4201 2701 4236
rect 2777 4221 2785 4276
rect 2937 4316 2949 4322
rect 2997 4316 3009 4322
rect 2553 4124 2560 4167
rect 2616 4124 2624 4179
rect 2699 4165 2707 4187
rect 2700 4158 2725 4165
rect 2657 4144 2709 4147
rect 1779 4098 1791 4104
rect 1879 4098 1891 4104
rect 1937 4098 1949 4104
rect 1985 4098 1997 4104
rect 2047 4098 2059 4104
rect 2099 4098 2111 4104
rect 2231 4098 2243 4104
rect 2301 4098 2313 4104
rect 2363 4098 2375 4104
rect 2411 4098 2423 4104
rect 2469 4098 2481 4104
rect 2531 4098 2543 4104
rect 2571 4098 2583 4104
rect 2669 4138 2697 4144
rect 2717 4144 2725 4158
rect 2777 4158 2785 4207
rect 2879 4201 2887 4236
rect 2873 4165 2881 4187
rect 2956 4193 2964 4276
rect 3067 4322 4073 4324
rect 3111 4316 3123 4322
rect 3157 4316 3169 4322
rect 3215 4316 3227 4322
rect 3261 4316 3273 4322
rect 3327 4316 3339 4322
rect 3377 4316 3389 4322
rect 3447 4316 3459 4322
rect 3020 4229 3037 4236
rect 3020 4181 3027 4229
rect 3096 4193 3104 4276
rect 3187 4262 3199 4296
rect 3241 4270 3253 4276
rect 3295 4270 3303 4276
rect 3245 4258 3267 4270
rect 3295 4256 3313 4270
rect 3193 4238 3199 4256
rect 3217 4246 3247 4252
rect 3295 4250 3303 4256
rect 2855 4158 2880 4165
rect 2777 4152 2801 4158
rect 2789 4144 2801 4152
rect 2855 4144 2863 4158
rect 2871 4144 2923 4147
rect 2883 4138 2911 4144
rect 2956 4124 2964 4179
rect 3020 4124 3027 4167
rect 3096 4124 3104 4179
rect 3137 4173 3145 4236
rect 3159 4224 3173 4232
rect 3193 4232 3233 4238
rect 3153 4173 3167 4187
rect 3137 4159 3153 4173
rect 3227 4160 3233 4232
rect 3241 4232 3247 4246
rect 3265 4242 3303 4250
rect 3497 4316 3509 4322
rect 3537 4316 3549 4322
rect 3577 4316 3589 4322
rect 3617 4316 3629 4322
rect 3657 4316 3669 4322
rect 3697 4316 3709 4322
rect 3737 4316 3749 4322
rect 3241 4226 3285 4232
rect 3297 4228 3359 4236
rect 3287 4187 3314 4194
rect 3334 4176 3340 4181
rect 3306 4168 3340 4176
rect 3294 4160 3301 4168
rect 3137 4144 3145 4159
rect 3227 4154 3301 4160
rect 3227 4152 3233 4154
rect 3294 4148 3301 4154
rect 3187 4130 3198 4138
rect 3191 4124 3198 4130
rect 3248 4136 3269 4143
rect 3353 4144 3359 4228
rect 3417 4201 3425 4236
rect 3517 4221 3525 4276
rect 3777 4316 3789 4322
rect 3817 4316 3829 4322
rect 3857 4316 3869 4322
rect 3897 4316 3909 4322
rect 3951 4316 3963 4322
rect 3991 4316 4003 4322
rect 4017 4316 4029 4322
rect 4087 4322 4513 4324
rect 4096 4316 4108 4322
rect 4146 4316 4158 4322
rect 3597 4230 3609 4236
rect 3637 4230 3649 4236
rect 3677 4230 3689 4236
rect 3717 4230 3729 4236
rect 3597 4222 3623 4230
rect 3637 4222 3662 4230
rect 3677 4222 3702 4230
rect 3717 4222 3735 4230
rect 3416 4161 3424 4187
rect 3416 4154 3445 4161
rect 3248 4124 3255 4136
rect 3313 4124 3320 4130
rect 3307 4118 3320 4124
rect 3377 4144 3429 4146
rect 3439 4144 3445 4154
rect 3517 4158 3525 4207
rect 3615 4176 3623 4222
rect 3654 4176 3662 4222
rect 3694 4176 3702 4222
rect 3728 4193 3735 4222
rect 3797 4221 3805 4276
rect 3877 4221 3885 4276
rect 3975 4221 3983 4276
rect 3728 4179 3733 4193
rect 3615 4164 3630 4176
rect 3654 4164 3670 4176
rect 3694 4164 3710 4176
rect 3615 4158 3623 4164
rect 3654 4158 3662 4164
rect 3694 4158 3702 4164
rect 3728 4158 3735 4179
rect 3517 4152 3541 4158
rect 3529 4144 3541 4152
rect 3596 4150 3623 4158
rect 3637 4150 3662 4158
rect 3676 4150 3702 4158
rect 3716 4151 3735 4158
rect 3797 4158 3805 4207
rect 3877 4158 3885 4207
rect 3975 4158 3983 4207
rect 4036 4193 4044 4276
rect 4182 4316 4194 4322
rect 4232 4316 4244 4322
rect 4301 4316 4313 4322
rect 4367 4316 4379 4322
rect 4413 4316 4425 4322
rect 4471 4316 4483 4322
rect 4337 4270 4345 4276
rect 4387 4270 4399 4276
rect 4327 4256 4345 4270
rect 4373 4258 4395 4270
rect 4441 4262 4453 4296
rect 4337 4250 4345 4256
rect 4337 4242 4375 4250
rect 4393 4246 4423 4252
rect 4119 4201 4127 4236
rect 4213 4201 4221 4236
rect 4281 4228 4343 4236
rect 3797 4152 3821 4158
rect 3877 4152 3901 4158
rect 3716 4150 3734 4151
rect 3596 4144 3608 4150
rect 3637 4144 3649 4150
rect 3676 4144 3688 4150
rect 3716 4144 3728 4150
rect 3809 4144 3821 4152
rect 3889 4144 3901 4152
rect 3389 4140 3417 4144
rect 3429 4104 3457 4110
rect 2597 4098 2609 4104
rect 2677 4098 2689 4104
rect 2759 4098 2771 4104
rect 2891 4098 2903 4104
rect 2937 4098 2949 4104
rect 2997 4098 3009 4104
rect 3037 4098 3049 4104
rect 3111 4098 3123 4104
rect 3159 4098 3171 4104
rect 3217 4098 3229 4104
rect 3265 4098 3277 4104
rect 3327 4098 3339 4104
rect 3397 4098 3409 4104
rect 3499 4098 3511 4104
rect 3577 4098 3589 4104
rect 3617 4098 3629 4104
rect 3657 4098 3669 4104
rect 3697 4098 3709 4104
rect 3737 4098 3749 4104
rect 3959 4152 3983 4158
rect 3959 4144 3971 4152
rect 4036 4124 4044 4179
rect 4113 4165 4121 4187
rect 4219 4165 4227 4187
rect 4095 4158 4120 4165
rect 4220 4158 4245 4165
rect 4095 4144 4103 4158
rect 3779 4098 3791 4104
rect 3859 4098 3871 4104
rect 3989 4098 4001 4104
rect 4111 4144 4163 4147
rect 4123 4138 4151 4144
rect 4177 4144 4229 4147
rect 4189 4138 4217 4144
rect 4237 4144 4245 4158
rect 4281 4144 4287 4228
rect 4393 4232 4399 4246
rect 4441 4238 4447 4256
rect 4355 4226 4399 4232
rect 4407 4232 4447 4238
rect 4326 4187 4353 4194
rect 4300 4176 4306 4181
rect 4300 4168 4334 4176
rect 4339 4160 4346 4168
rect 4407 4160 4413 4232
rect 4527 4322 5253 4324
rect 4536 4316 4548 4322
rect 4586 4316 4598 4322
rect 4641 4316 4653 4322
rect 4707 4316 4719 4322
rect 4753 4316 4765 4322
rect 4811 4316 4823 4322
rect 4891 4316 4903 4322
rect 4971 4316 4983 4322
rect 5017 4316 5029 4322
rect 5057 4316 5069 4322
rect 5151 4316 5163 4322
rect 4677 4270 4685 4276
rect 4727 4270 4739 4276
rect 4667 4256 4685 4270
rect 4713 4258 4735 4270
rect 4781 4262 4793 4296
rect 4677 4250 4685 4256
rect 4677 4242 4715 4250
rect 4733 4246 4763 4252
rect 4467 4224 4481 4232
rect 4473 4173 4487 4187
rect 4495 4173 4503 4236
rect 4559 4201 4567 4236
rect 4621 4228 4683 4236
rect 4339 4154 4413 4160
rect 4487 4159 4503 4173
rect 4553 4165 4561 4187
rect 4339 4148 4346 4154
rect 4407 4152 4413 4154
rect 4371 4136 4392 4143
rect 4495 4144 4503 4159
rect 4535 4158 4560 4165
rect 4535 4144 4543 4158
rect 4320 4124 4327 4130
rect 4385 4124 4392 4136
rect 4442 4130 4453 4138
rect 4442 4124 4449 4130
rect 4320 4118 4333 4124
rect 4551 4144 4603 4147
rect 4563 4138 4591 4144
rect 4621 4144 4627 4228
rect 4733 4232 4739 4246
rect 4781 4238 4787 4256
rect 4695 4226 4739 4232
rect 4747 4232 4787 4238
rect 4666 4187 4693 4194
rect 4640 4176 4646 4181
rect 4640 4168 4674 4176
rect 4679 4160 4686 4168
rect 4747 4160 4753 4232
rect 5038 4274 5049 4276
rect 5182 4316 5194 4322
rect 5232 4316 5244 4322
rect 5077 4274 5085 4276
rect 5038 4268 5085 4274
rect 4991 4242 5003 4244
rect 4963 4236 5003 4242
rect 4807 4224 4821 4232
rect 4813 4173 4827 4187
rect 4835 4173 4843 4236
rect 4876 4201 4884 4236
rect 4934 4201 4942 4236
rect 5078 4213 5085 4268
rect 4679 4154 4753 4160
rect 4827 4159 4843 4173
rect 4679 4148 4686 4154
rect 4747 4152 4753 4154
rect 4711 4136 4732 4143
rect 4835 4144 4843 4159
rect 4876 4144 4884 4187
rect 4934 4144 4942 4187
rect 5076 4171 5084 4199
rect 4660 4124 4667 4130
rect 4725 4124 4732 4136
rect 4782 4130 4793 4138
rect 4782 4124 4789 4130
rect 4660 4118 4673 4124
rect 4934 4133 4960 4144
rect 4017 4098 4029 4104
rect 4131 4098 4143 4104
rect 4197 4098 4209 4104
rect 4301 4098 4313 4104
rect 4363 4098 4375 4104
rect 4411 4098 4423 4104
rect 4469 4098 4481 4104
rect 4571 4098 4583 4104
rect 4641 4098 4653 4104
rect 4703 4098 4715 4104
rect 4751 4098 4763 4104
rect 4809 4098 4821 4104
rect 4891 4098 4903 4104
rect 4938 4098 4950 4104
rect 4988 4098 5000 4104
rect 5054 4162 5084 4171
rect 5066 4160 5084 4162
rect 5097 4143 5103 4233
rect 5136 4193 5144 4276
rect 5267 4322 6736 4324
rect 5301 4316 5313 4322
rect 5367 4316 5379 4322
rect 5413 4316 5425 4322
rect 5471 4316 5483 4322
rect 5517 4316 5529 4322
rect 5557 4316 5569 4322
rect 5337 4270 5345 4276
rect 5387 4270 5399 4276
rect 5327 4256 5345 4270
rect 5373 4258 5395 4270
rect 5441 4262 5453 4296
rect 5337 4250 5345 4256
rect 5337 4242 5375 4250
rect 5393 4246 5423 4252
rect 5213 4201 5221 4236
rect 5281 4228 5343 4236
rect 5087 4137 5103 4143
rect 5136 4124 5144 4179
rect 5219 4165 5227 4187
rect 5220 4158 5245 4165
rect 5177 4144 5229 4147
rect 5189 4138 5217 4144
rect 5237 4144 5245 4158
rect 5281 4144 5287 4228
rect 5393 4232 5399 4246
rect 5441 4238 5447 4256
rect 5355 4226 5399 4232
rect 5407 4232 5447 4238
rect 5326 4187 5353 4194
rect 5300 4176 5306 4181
rect 5300 4168 5334 4176
rect 5339 4160 5346 4168
rect 5407 4160 5413 4232
rect 5597 4316 5609 4322
rect 5662 4316 5674 4322
rect 5712 4316 5724 4322
rect 5787 4316 5799 4322
rect 5831 4316 5843 4322
rect 5467 4224 5481 4232
rect 5473 4173 5487 4187
rect 5495 4173 5503 4236
rect 5537 4221 5545 4276
rect 5339 4154 5413 4160
rect 5487 4159 5503 4173
rect 5339 4148 5346 4154
rect 5407 4152 5413 4154
rect 5371 4136 5392 4143
rect 5495 4144 5503 4159
rect 5537 4158 5545 4207
rect 5616 4193 5624 4276
rect 5857 4316 5869 4322
rect 5897 4316 5909 4322
rect 5991 4316 6003 4322
rect 5693 4201 5701 4236
rect 5771 4201 5779 4236
rect 5537 4152 5561 4158
rect 5549 4144 5561 4152
rect 5320 4124 5327 4130
rect 5385 4124 5392 4136
rect 5442 4130 5453 4138
rect 5442 4124 5449 4130
rect 5320 4118 5333 4124
rect 5616 4124 5624 4179
rect 5699 4165 5707 4187
rect 5771 4187 5773 4201
rect 5700 4158 5725 4165
rect 5657 4144 5709 4147
rect 5669 4138 5697 4144
rect 5717 4144 5725 4158
rect 5771 4144 5779 4187
rect 5814 4162 5822 4276
rect 5878 4274 5889 4276
rect 5917 4274 5925 4276
rect 5878 4268 5925 4274
rect 5918 4213 5925 4268
rect 6022 4316 6034 4322
rect 6072 4316 6084 4322
rect 6139 4316 6151 4322
rect 6197 4316 6209 4322
rect 6237 4316 6249 4322
rect 6307 4316 6319 4322
rect 6351 4316 6363 4322
rect 5916 4171 5924 4199
rect 5976 4201 5984 4236
rect 6053 4201 6061 4236
rect 6117 4230 6125 4276
rect 6117 4224 6143 4230
rect 6140 4218 6143 4224
rect 5805 4154 5843 4162
rect 5831 4144 5843 4154
rect 5771 4134 5781 4144
rect 5894 4162 5924 4171
rect 5957 4163 5963 4193
rect 5906 4160 5924 4162
rect 5937 4157 5963 4163
rect 5937 4143 5943 4157
rect 5976 4144 5984 4187
rect 6059 4165 6067 4187
rect 6060 4158 6085 4165
rect 6017 4144 6069 4147
rect 5927 4137 5943 4143
rect 6029 4138 6057 4144
rect 6077 4144 6085 4158
rect 6140 4162 6147 4218
rect 6161 4201 6169 4236
rect 6217 4221 6225 4276
rect 6377 4316 6389 4322
rect 6417 4316 6429 4322
rect 6457 4316 6469 4322
rect 6571 4316 6583 4322
rect 6617 4316 6629 4322
rect 6657 4316 6669 4322
rect 6167 4187 6169 4201
rect 6140 4156 6143 4162
rect 6121 4150 6143 4156
rect 6121 4124 6129 4150
rect 6161 4144 6169 4187
rect 6217 4158 6225 4207
rect 6291 4201 6299 4236
rect 6291 4187 6293 4201
rect 6217 4152 6241 4158
rect 6229 4144 6241 4152
rect 6291 4144 6299 4187
rect 6334 4162 6342 4276
rect 6397 4221 6405 4276
rect 6437 4217 6453 4223
rect 6325 4154 6363 4162
rect 6351 4144 6363 4154
rect 6397 4158 6405 4207
rect 6437 4187 6443 4217
rect 6476 4193 6484 4276
rect 6638 4274 6649 4276
rect 6677 4274 6685 4276
rect 6638 4268 6685 4274
rect 6591 4242 6603 4244
rect 6563 4236 6603 4242
rect 6534 4201 6542 4236
rect 6678 4213 6685 4268
rect 6397 4152 6421 4158
rect 6409 4144 6421 4152
rect 6291 4134 6301 4144
rect 6476 4124 6484 4179
rect 6534 4144 6542 4187
rect 6676 4171 6684 4199
rect 6534 4133 6560 4144
rect 5018 4098 5030 4104
rect 5151 4098 5163 4104
rect 5197 4098 5209 4104
rect 5301 4098 5313 4104
rect 5363 4098 5375 4104
rect 5411 4098 5423 4104
rect 5469 4098 5481 4104
rect 5519 4098 5531 4104
rect 5597 4098 5609 4104
rect 5677 4098 5689 4104
rect 5801 4098 5813 4104
rect 5858 4098 5870 4104
rect 5991 4098 6003 4104
rect 6037 4098 6049 4104
rect 6139 4098 6151 4104
rect 6199 4098 6211 4104
rect 6321 4098 6333 4104
rect 6379 4098 6391 4104
rect 6457 4098 6469 4104
rect 6538 4098 6550 4104
rect 6588 4098 6600 4104
rect 6654 4162 6684 4171
rect 6666 4160 6684 4162
rect 6618 4098 6630 4104
rect 6742 4098 6802 4562
rect 4 4096 6802 4098
rect 6736 4084 6802 4096
rect 4 4082 6802 4084
rect 49 4076 61 4082
rect 119 4076 131 4082
rect 177 4076 189 4082
rect 225 4076 237 4082
rect 287 4076 299 4082
rect 339 4076 351 4082
rect 438 4076 450 4082
rect 488 4076 500 4082
rect 569 4076 581 4082
rect 649 4076 661 4082
rect 709 4076 721 4082
rect 779 4076 791 4082
rect 837 4076 849 4082
rect 885 4076 897 4082
rect 947 4076 959 4082
rect 1049 4076 1061 4082
rect 31 3993 39 4036
rect 71 4030 79 4056
rect 57 4024 79 4030
rect 267 4056 280 4062
rect 151 4050 158 4056
rect 147 4042 158 4050
rect 208 4044 215 4056
rect 273 4050 280 4056
rect 57 4018 60 4024
rect 31 3979 33 3993
rect 31 3944 39 3979
rect 53 3962 60 4018
rect 97 4021 105 4036
rect 208 4037 229 4044
rect 187 4026 193 4028
rect 254 4026 261 4032
rect 97 4007 113 4021
rect 187 4020 261 4026
rect 57 3956 60 3962
rect 57 3950 83 3956
rect 75 3904 83 3950
rect 97 3944 105 4007
rect 113 3993 127 4007
rect 119 3948 133 3956
rect 187 3948 193 4020
rect 254 4012 261 4020
rect 266 4004 300 4012
rect 294 3999 300 4004
rect 247 3986 274 3993
rect 153 3942 193 3948
rect 201 3948 245 3954
rect 153 3924 159 3942
rect 201 3934 207 3948
rect 313 3952 319 4036
rect 369 4028 381 4036
rect 357 4022 381 4028
rect 434 4036 460 4047
rect 357 3973 365 4022
rect 434 3993 442 4036
rect 539 4028 551 4036
rect 619 4028 631 4036
rect 539 4022 563 4028
rect 619 4022 643 4028
rect 257 3944 319 3952
rect 177 3928 207 3934
rect 225 3930 263 3938
rect 255 3924 263 3930
rect 147 3884 159 3918
rect 205 3910 227 3922
rect 255 3910 273 3924
rect 201 3904 213 3910
rect 255 3904 263 3910
rect 357 3904 365 3959
rect 434 3944 442 3979
rect 555 3973 563 4022
rect 635 3973 643 4022
rect 691 3993 699 4036
rect 731 4030 739 4056
rect 717 4024 739 4030
rect 927 4056 940 4062
rect 811 4050 818 4056
rect 807 4042 818 4050
rect 868 4044 875 4056
rect 933 4050 940 4056
rect 717 4018 720 4024
rect 691 3979 693 3993
rect 463 3938 503 3944
rect 491 3936 503 3938
rect 555 3904 563 3959
rect 587 3937 613 3943
rect 635 3904 643 3959
rect 691 3944 699 3979
rect 713 3962 720 4018
rect 757 4021 765 4036
rect 868 4037 889 4044
rect 847 4026 853 4028
rect 914 4026 921 4032
rect 757 4007 773 4021
rect 847 4020 921 4026
rect 717 3956 720 3962
rect 717 3950 743 3956
rect 49 3858 61 3864
rect 117 3858 129 3864
rect 175 3858 187 3864
rect 221 3858 233 3864
rect 287 3858 299 3864
rect 337 3858 349 3864
rect 377 3858 389 3864
rect 471 3858 483 3864
rect 531 3858 543 3864
rect 571 3858 583 3864
rect 735 3904 743 3950
rect 757 3944 765 4007
rect 773 3993 787 4007
rect 779 3948 793 3956
rect 847 3948 853 4020
rect 914 4012 921 4020
rect 926 4004 960 4012
rect 954 3999 960 4004
rect 907 3986 934 3993
rect 813 3942 853 3948
rect 861 3948 905 3954
rect 813 3924 819 3942
rect 861 3934 867 3948
rect 973 3952 979 4036
rect 1079 4076 1091 4082
rect 1159 4076 1171 4082
rect 1258 4076 1270 4082
rect 1308 4076 1320 4082
rect 1359 4076 1371 4082
rect 1417 4076 1429 4082
rect 1465 4076 1477 4082
rect 1527 4076 1539 4082
rect 1629 4076 1641 4082
rect 1679 4076 1691 4082
rect 1739 4076 1751 4082
rect 1839 4076 1851 4082
rect 1897 4076 1909 4082
rect 1945 4076 1957 4082
rect 2007 4076 2019 4082
rect 2059 4076 2071 4082
rect 2191 4076 2203 4082
rect 2289 4076 2301 4082
rect 1019 4028 1031 4036
rect 1109 4028 1121 4036
rect 1189 4028 1201 4036
rect 1019 4022 1043 4028
rect 1035 3973 1043 4022
rect 1097 4022 1121 4028
rect 1097 3973 1105 4022
rect 1177 4022 1201 4028
rect 1254 4036 1280 4047
rect 1507 4056 1520 4062
rect 1391 4050 1398 4056
rect 1387 4042 1398 4050
rect 1448 4044 1455 4056
rect 1513 4050 1520 4056
rect 917 3944 979 3952
rect 837 3928 867 3934
rect 885 3930 923 3938
rect 915 3924 923 3930
rect 807 3884 819 3918
rect 865 3910 887 3922
rect 915 3910 933 3924
rect 861 3904 873 3910
rect 915 3904 923 3910
rect 1035 3904 1043 3959
rect 1097 3904 1105 3959
rect 1137 3927 1143 4013
rect 1177 3973 1185 4022
rect 1254 3993 1262 4036
rect 1337 4021 1345 4036
rect 1448 4037 1469 4044
rect 1427 4026 1433 4028
rect 1494 4026 1501 4032
rect 1337 4007 1353 4021
rect 1427 4020 1501 4026
rect 1177 3904 1185 3959
rect 1254 3944 1262 3979
rect 1337 3944 1345 4007
rect 1353 3993 1367 4007
rect 1359 3948 1373 3956
rect 611 3858 623 3864
rect 651 3858 663 3864
rect 709 3858 721 3864
rect 777 3858 789 3864
rect 835 3858 847 3864
rect 881 3858 893 3864
rect 947 3858 959 3864
rect 1011 3858 1023 3864
rect 1051 3858 1063 3864
rect 1077 3858 1089 3864
rect 1117 3858 1129 3864
rect 1283 3938 1323 3944
rect 1311 3936 1323 3938
rect 1427 3948 1433 4020
rect 1494 4012 1501 4020
rect 1506 4004 1540 4012
rect 1534 3999 1540 4004
rect 1487 3986 1514 3993
rect 1393 3942 1433 3948
rect 1441 3948 1485 3954
rect 1393 3924 1399 3942
rect 1441 3934 1447 3948
rect 1553 3952 1559 4036
rect 1599 4028 1611 4036
rect 1661 4030 1669 4056
rect 1599 4022 1623 4028
rect 1661 4024 1683 4030
rect 1615 3973 1623 4022
rect 1680 4018 1683 4024
rect 1680 3962 1687 4018
rect 1701 3993 1709 4036
rect 1769 4028 1781 4036
rect 1757 4022 1781 4028
rect 1987 4056 2000 4062
rect 1871 4050 1878 4056
rect 1867 4042 1878 4050
rect 1928 4044 1935 4056
rect 1993 4050 2000 4056
rect 1707 3979 1709 3993
rect 1497 3944 1559 3952
rect 1417 3928 1447 3934
rect 1465 3930 1503 3938
rect 1495 3924 1503 3930
rect 1387 3884 1399 3918
rect 1445 3910 1467 3922
rect 1495 3910 1513 3924
rect 1441 3904 1453 3910
rect 1495 3904 1503 3910
rect 1615 3904 1623 3959
rect 1680 3956 1683 3962
rect 1657 3950 1683 3956
rect 1657 3904 1665 3950
rect 1701 3944 1709 3979
rect 1757 3973 1765 4022
rect 1817 4021 1825 4036
rect 1928 4037 1949 4044
rect 1907 4026 1913 4028
rect 1974 4026 1981 4032
rect 1817 4007 1833 4021
rect 1907 4020 1981 4026
rect 1757 3904 1765 3959
rect 1817 3944 1825 4007
rect 1833 3993 1847 4007
rect 1839 3948 1853 3956
rect 1907 3948 1913 4020
rect 1974 4012 1981 4020
rect 1986 4004 2020 4012
rect 2014 3999 2020 4004
rect 1967 3986 1994 3993
rect 1873 3942 1913 3948
rect 1921 3948 1965 3954
rect 1873 3924 1879 3942
rect 1921 3934 1927 3948
rect 2033 3952 2039 4036
rect 2089 4028 2101 4036
rect 2077 4022 2101 4028
rect 2155 4022 2163 4036
rect 2183 4036 2211 4042
rect 2171 4033 2223 4036
rect 2319 4076 2331 4082
rect 2431 4076 2443 4082
rect 2511 4076 2523 4082
rect 2557 4076 2569 4082
rect 2597 4076 2609 4082
rect 2259 4028 2271 4036
rect 2349 4028 2361 4036
rect 2259 4022 2283 4028
rect 2077 3973 2085 4022
rect 2155 4015 2180 4022
rect 2173 3993 2181 4015
rect 1977 3944 2039 3952
rect 1897 3928 1927 3934
rect 1945 3930 1983 3938
rect 1975 3924 1983 3930
rect 1867 3884 1879 3918
rect 1925 3910 1947 3922
rect 1975 3910 1993 3924
rect 1921 3904 1933 3910
rect 1975 3904 1983 3910
rect 2077 3904 2085 3959
rect 2179 3944 2187 3979
rect 2275 3973 2283 4022
rect 2337 4022 2361 4028
rect 2337 3973 2345 4022
rect 2416 4001 2424 4056
rect 2475 4022 2483 4036
rect 2503 4036 2531 4042
rect 2651 4076 2663 4082
rect 2691 4076 2703 4082
rect 2717 4076 2729 4082
rect 2811 4076 2823 4082
rect 2889 4076 2901 4082
rect 2491 4033 2543 4036
rect 2475 4015 2500 4022
rect 2493 3993 2501 4015
rect 2580 4013 2587 4056
rect 1157 3858 1169 3864
rect 1197 3858 1209 3864
rect 1291 3858 1303 3864
rect 1357 3858 1369 3864
rect 1415 3858 1427 3864
rect 1461 3858 1473 3864
rect 1527 3858 1539 3864
rect 1591 3858 1603 3864
rect 1631 3858 1643 3864
rect 1679 3858 1691 3864
rect 1737 3858 1749 3864
rect 1777 3858 1789 3864
rect 1837 3858 1849 3864
rect 1895 3858 1907 3864
rect 1941 3858 1953 3864
rect 2007 3858 2019 3864
rect 2057 3858 2069 3864
rect 2097 3858 2109 3864
rect 2275 3904 2283 3959
rect 2337 3904 2345 3959
rect 2416 3904 2424 3987
rect 2499 3944 2507 3979
rect 2580 3951 2587 3999
rect 2673 4013 2680 4056
rect 2736 4001 2744 4056
rect 2796 4001 2804 4056
rect 2917 4076 2929 4082
rect 2957 4076 2969 4082
rect 3017 4076 3029 4082
rect 3097 4076 3109 4082
rect 3157 4076 3169 4082
rect 3197 4076 3209 4082
rect 3289 4076 3301 4082
rect 3369 4076 3381 4082
rect 3421 4076 3433 4082
rect 3483 4076 3495 4082
rect 3531 4076 3543 4082
rect 3589 4076 3601 4082
rect 3671 4076 3683 4082
rect 3721 4076 3733 4082
rect 3783 4076 3795 4082
rect 3831 4076 3843 4082
rect 3889 4076 3901 4082
rect 4010 4076 4022 4082
rect 2859 4028 2871 4036
rect 2859 4022 2883 4028
rect 2673 3951 2680 3999
rect 2580 3944 2597 3951
rect 2156 3858 2168 3864
rect 2206 3858 2218 3864
rect 2251 3858 2263 3864
rect 2291 3858 2303 3864
rect 2317 3858 2329 3864
rect 2357 3858 2369 3864
rect 2431 3858 2443 3864
rect 2476 3858 2488 3864
rect 2526 3858 2538 3864
rect 2663 3944 2680 3951
rect 2736 3904 2744 3987
rect 2796 3904 2804 3987
rect 2875 3973 2883 4022
rect 2940 4013 2947 4056
rect 3009 4036 3037 4042
rect 2997 4033 3049 4036
rect 3057 4022 3065 4036
rect 3040 4015 3065 4022
rect 2875 3904 2883 3959
rect 2940 3951 2947 3999
rect 3039 3993 3047 4015
rect 3116 4001 3124 4056
rect 3180 4013 3187 4056
rect 3440 4056 3453 4062
rect 3440 4050 3447 4056
rect 3505 4044 3512 4056
rect 3259 4028 3271 4036
rect 3339 4028 3351 4036
rect 3259 4022 3283 4028
rect 3339 4022 3363 4028
rect 2940 3944 2957 3951
rect 3033 3944 3041 3979
rect 2557 3858 2569 3864
rect 2691 3858 2703 3864
rect 2717 3858 2729 3864
rect 2811 3858 2823 3864
rect 2851 3858 2863 3864
rect 2891 3858 2903 3864
rect 3116 3904 3124 3987
rect 3180 3951 3187 3999
rect 3275 3973 3283 4022
rect 3355 3973 3363 4022
rect 3180 3944 3197 3951
rect 2917 3858 2929 3864
rect 3002 3858 3014 3864
rect 3052 3858 3064 3864
rect 3275 3904 3283 3959
rect 3355 3904 3363 3959
rect 3401 3952 3407 4036
rect 3491 4037 3512 4044
rect 3562 4050 3569 4056
rect 3562 4042 3573 4050
rect 3459 4026 3466 4032
rect 3527 4026 3533 4028
rect 3459 4020 3533 4026
rect 3615 4021 3623 4036
rect 3459 4012 3466 4020
rect 3420 4004 3454 4012
rect 3420 3999 3426 4004
rect 3446 3986 3473 3993
rect 3401 3944 3463 3952
rect 3475 3948 3519 3954
rect 3097 3858 3109 3864
rect 3157 3858 3169 3864
rect 3251 3858 3263 3864
rect 3291 3858 3303 3864
rect 3457 3930 3495 3938
rect 3513 3934 3519 3948
rect 3527 3948 3533 4020
rect 3607 4007 3623 4021
rect 3593 3993 3607 4007
rect 3527 3942 3567 3948
rect 3587 3948 3601 3956
rect 3615 3944 3623 4007
rect 3656 4001 3664 4056
rect 3740 4056 3753 4062
rect 3740 4050 3747 4056
rect 3805 4044 3812 4056
rect 3457 3924 3465 3930
rect 3513 3928 3543 3934
rect 3561 3924 3567 3942
rect 3447 3910 3465 3924
rect 3493 3910 3515 3922
rect 3457 3904 3465 3910
rect 3507 3904 3519 3910
rect 3561 3884 3573 3918
rect 3656 3904 3664 3987
rect 3701 3952 3707 4036
rect 3791 4037 3812 4044
rect 3862 4050 3869 4056
rect 3862 4042 3873 4050
rect 3759 4026 3766 4032
rect 3827 4026 3833 4028
rect 3759 4020 3833 4026
rect 3915 4021 3923 4036
rect 3759 4012 3766 4020
rect 3720 4004 3754 4012
rect 3720 3999 3726 4004
rect 3746 3986 3773 3993
rect 3701 3944 3763 3952
rect 3775 3948 3819 3954
rect 3757 3930 3795 3938
rect 3813 3934 3819 3948
rect 3827 3948 3833 4020
rect 3907 4007 3923 4021
rect 3893 3993 3907 4007
rect 3827 3942 3867 3948
rect 3887 3948 3901 3956
rect 3915 3944 3923 4007
rect 3956 4018 3974 4020
rect 3956 4009 3986 4018
rect 4039 4076 4051 4082
rect 4171 4076 4183 4082
rect 4217 4076 4229 4082
rect 4257 4076 4269 4082
rect 4331 4076 4343 4082
rect 4409 4076 4421 4082
rect 4491 4076 4503 4082
rect 4561 4076 4573 4082
rect 4623 4076 4635 4082
rect 4671 4076 4683 4082
rect 4729 4076 4741 4082
rect 4829 4076 4841 4082
rect 4911 4076 4923 4082
rect 4981 4076 4993 4082
rect 5043 4076 5055 4082
rect 5091 4076 5103 4082
rect 5149 4076 5161 4082
rect 5249 4076 5261 4082
rect 5331 4076 5343 4082
rect 5429 4076 5441 4082
rect 5477 4076 5489 4082
rect 5591 4076 5603 4082
rect 5641 4076 5653 4082
rect 5703 4076 5715 4082
rect 5751 4076 5763 4082
rect 5809 4076 5821 4082
rect 5857 4076 5869 4082
rect 5990 4076 6002 4082
rect 6039 4076 6051 4082
rect 6097 4076 6109 4082
rect 6145 4076 6157 4082
rect 6207 4076 6219 4082
rect 6279 4076 6291 4082
rect 6337 4076 6349 4082
rect 6385 4076 6397 4082
rect 6447 4076 6459 4082
rect 6519 4076 6531 4082
rect 6577 4076 6589 4082
rect 6625 4076 6637 4082
rect 6687 4076 6699 4082
rect 4069 4028 4081 4036
rect 4057 4022 4081 4028
rect 3956 3981 3964 4009
rect 3757 3924 3765 3930
rect 3813 3928 3843 3934
rect 3861 3924 3867 3942
rect 3747 3910 3765 3924
rect 3793 3910 3815 3922
rect 3757 3904 3765 3910
rect 3807 3904 3819 3910
rect 3861 3884 3873 3918
rect 3955 3912 3962 3967
rect 4057 3973 4065 4022
rect 4135 4022 4143 4036
rect 4163 4036 4191 4042
rect 4151 4033 4203 4036
rect 4135 4015 4160 4022
rect 3955 3906 4002 3912
rect 3955 3904 3963 3906
rect 3991 3904 4002 3906
rect 4057 3904 4065 3959
rect 4097 3943 4103 4013
rect 4153 3993 4161 4015
rect 4240 4013 4247 4056
rect 4316 4001 4324 4056
rect 4379 4028 4391 4036
rect 4379 4022 4403 4028
rect 4159 3944 4167 3979
rect 4240 3951 4247 3999
rect 4240 3944 4257 3951
rect 4087 3937 4103 3943
rect 3331 3858 3343 3864
rect 3371 3858 3383 3864
rect 3421 3858 3433 3864
rect 3487 3858 3499 3864
rect 3533 3858 3545 3864
rect 3591 3858 3603 3864
rect 3671 3858 3683 3864
rect 3721 3858 3733 3864
rect 3787 3858 3799 3864
rect 3833 3858 3845 3864
rect 3891 3858 3903 3864
rect 3971 3858 3983 3864
rect 4011 3858 4023 3864
rect 4037 3858 4049 3864
rect 4077 3858 4089 3864
rect -62 3856 4113 3858
rect 4136 3858 4148 3864
rect 4186 3858 4198 3864
rect 4316 3904 4324 3987
rect 4395 3973 4403 4022
rect 4455 4022 4463 4036
rect 4483 4036 4511 4042
rect 4471 4033 4523 4036
rect 4580 4056 4593 4062
rect 4580 4050 4587 4056
rect 4645 4044 4652 4056
rect 4455 4015 4480 4022
rect 4473 3993 4481 4015
rect 4395 3904 4403 3959
rect 4479 3944 4487 3979
rect 4541 3952 4547 4036
rect 4631 4037 4652 4044
rect 4702 4050 4709 4056
rect 4702 4042 4713 4050
rect 4599 4026 4606 4032
rect 4667 4026 4673 4028
rect 4599 4020 4673 4026
rect 4755 4021 4763 4036
rect 4799 4028 4811 4036
rect 4799 4022 4823 4028
rect 4599 4012 4606 4020
rect 4560 4004 4594 4012
rect 4560 3999 4566 4004
rect 4586 3986 4613 3993
rect 4541 3944 4603 3952
rect 4615 3948 4659 3954
rect 4217 3858 4229 3864
rect 4331 3858 4343 3864
rect 4371 3858 4383 3864
rect 4411 3858 4423 3864
rect 4127 3856 4433 3858
rect 4597 3930 4635 3938
rect 4653 3934 4659 3948
rect 4667 3948 4673 4020
rect 4747 4007 4763 4021
rect 4733 3993 4747 4007
rect 4667 3942 4707 3948
rect 4727 3948 4741 3956
rect 4755 3944 4763 4007
rect 4815 3973 4823 4022
rect 4875 4022 4883 4036
rect 4903 4036 4931 4042
rect 4891 4033 4943 4036
rect 5000 4056 5013 4062
rect 5000 4050 5007 4056
rect 5065 4044 5072 4056
rect 4875 4015 4900 4022
rect 4893 3993 4901 4015
rect 4597 3924 4605 3930
rect 4653 3928 4683 3934
rect 4701 3924 4707 3942
rect 4587 3910 4605 3924
rect 4633 3910 4655 3922
rect 4597 3904 4605 3910
rect 4647 3904 4659 3910
rect 4701 3884 4713 3918
rect 4815 3904 4823 3959
rect 4899 3944 4907 3979
rect 4961 3952 4967 4036
rect 5051 4037 5072 4044
rect 5122 4050 5129 4056
rect 5122 4042 5133 4050
rect 5019 4026 5026 4032
rect 5087 4026 5093 4028
rect 5019 4020 5093 4026
rect 5175 4021 5183 4036
rect 5219 4028 5231 4036
rect 5219 4022 5243 4028
rect 5019 4012 5026 4020
rect 4980 4004 5014 4012
rect 4980 3999 4986 4004
rect 5006 3986 5033 3993
rect 4961 3944 5023 3952
rect 5035 3948 5079 3954
rect 4456 3858 4468 3864
rect 4506 3858 4518 3864
rect 4561 3858 4573 3864
rect 4627 3858 4639 3864
rect 4673 3858 4685 3864
rect 4731 3858 4743 3864
rect 4791 3858 4803 3864
rect 4831 3858 4843 3864
rect 4447 3856 4853 3858
rect 5017 3930 5055 3938
rect 5073 3934 5079 3948
rect 5087 3948 5093 4020
rect 5167 4007 5183 4021
rect 5153 3993 5167 4007
rect 5087 3942 5127 3948
rect 5147 3948 5161 3956
rect 5175 3944 5183 4007
rect 5235 3973 5243 4022
rect 5295 4022 5303 4036
rect 5323 4036 5351 4042
rect 5311 4033 5363 4036
rect 5469 4036 5497 4042
rect 5399 4028 5411 4036
rect 5457 4033 5509 4036
rect 5399 4022 5423 4028
rect 5517 4022 5525 4036
rect 5295 4015 5320 4022
rect 5313 3993 5321 4015
rect 5017 3924 5025 3930
rect 5073 3928 5103 3934
rect 5121 3924 5127 3942
rect 5007 3910 5025 3924
rect 5053 3910 5075 3922
rect 5017 3904 5025 3910
rect 5067 3904 5079 3910
rect 5121 3884 5133 3918
rect 5235 3904 5243 3959
rect 5319 3944 5327 3979
rect 5415 3973 5423 4022
rect 5500 4015 5525 4022
rect 5499 3993 5507 4015
rect 4876 3858 4888 3864
rect 4926 3858 4938 3864
rect 4981 3858 4993 3864
rect 5047 3858 5059 3864
rect 5093 3858 5105 3864
rect 5151 3858 5163 3864
rect 5211 3858 5223 3864
rect 5251 3858 5263 3864
rect 4867 3856 5273 3858
rect 5415 3904 5423 3959
rect 5493 3944 5501 3979
rect 5557 3967 5563 4033
rect 5576 4001 5584 4056
rect 5660 4056 5673 4062
rect 5660 4050 5667 4056
rect 5725 4044 5732 4056
rect 5296 3858 5308 3864
rect 5346 3858 5358 3864
rect 5391 3858 5403 3864
rect 5431 3858 5443 3864
rect 5576 3904 5584 3987
rect 5621 3952 5627 4036
rect 5711 4037 5732 4044
rect 5782 4050 5789 4056
rect 5782 4042 5793 4050
rect 5679 4026 5686 4032
rect 5747 4026 5753 4028
rect 5679 4020 5753 4026
rect 5835 4021 5843 4036
rect 5679 4012 5686 4020
rect 5640 4004 5674 4012
rect 5640 3999 5646 4004
rect 5666 3986 5693 3993
rect 5621 3944 5683 3952
rect 5695 3948 5739 3954
rect 5677 3930 5715 3938
rect 5733 3934 5739 3948
rect 5747 3948 5753 4020
rect 5827 4007 5843 4021
rect 5813 3993 5827 4007
rect 5747 3942 5787 3948
rect 5807 3948 5821 3956
rect 5835 3944 5843 4007
rect 5876 4001 5884 4056
rect 5936 4018 5954 4020
rect 5936 4009 5966 4018
rect 6187 4056 6200 4062
rect 6071 4050 6078 4056
rect 6067 4042 6078 4050
rect 6128 4044 6135 4056
rect 6193 4050 6200 4056
rect 6017 4021 6025 4036
rect 6128 4037 6149 4044
rect 6107 4026 6113 4028
rect 6174 4026 6181 4032
rect 5677 3924 5685 3930
rect 5733 3928 5763 3934
rect 5781 3924 5787 3942
rect 5667 3910 5685 3924
rect 5713 3910 5735 3922
rect 5677 3904 5685 3910
rect 5727 3904 5739 3910
rect 5781 3884 5793 3918
rect 5876 3904 5884 3987
rect 5936 3981 5944 4009
rect 6017 4007 6033 4021
rect 6107 4020 6181 4026
rect 5935 3912 5942 3967
rect 6017 3944 6025 4007
rect 6033 3993 6047 4007
rect 6039 3948 6053 3956
rect 5935 3906 5982 3912
rect 5935 3904 5943 3906
rect 5971 3904 5982 3906
rect 6107 3948 6113 4020
rect 6174 4012 6181 4020
rect 6186 4004 6220 4012
rect 6214 3999 6220 4004
rect 6167 3986 6194 3993
rect 6073 3942 6113 3948
rect 6121 3948 6165 3954
rect 6073 3924 6079 3942
rect 6121 3934 6127 3948
rect 6233 3952 6239 4036
rect 6177 3944 6239 3952
rect 6097 3928 6127 3934
rect 6145 3930 6183 3938
rect 6175 3924 6183 3930
rect 6067 3884 6079 3918
rect 6125 3910 6147 3922
rect 6175 3910 6193 3924
rect 6121 3904 6133 3910
rect 6175 3904 6183 3910
rect 6427 4056 6440 4062
rect 6311 4050 6318 4056
rect 6307 4042 6318 4050
rect 6368 4044 6375 4056
rect 6433 4050 6440 4056
rect 6257 4021 6265 4036
rect 6368 4037 6389 4044
rect 6347 4026 6353 4028
rect 6414 4026 6421 4032
rect 6257 4007 6273 4021
rect 6347 4020 6421 4026
rect 6257 3944 6265 4007
rect 6273 3993 6287 4007
rect 6279 3948 6293 3956
rect 6347 3948 6353 4020
rect 6414 4012 6421 4020
rect 6426 4004 6460 4012
rect 6454 3999 6460 4004
rect 6407 3986 6434 3993
rect 6313 3942 6353 3948
rect 6361 3948 6405 3954
rect 6313 3924 6319 3942
rect 6361 3934 6367 3948
rect 6473 3952 6479 4036
rect 6417 3944 6479 3952
rect 6337 3928 6367 3934
rect 6385 3930 6423 3938
rect 6415 3924 6423 3930
rect 6307 3884 6319 3918
rect 6365 3910 6387 3922
rect 6415 3910 6433 3924
rect 6361 3904 6373 3910
rect 6415 3904 6423 3910
rect 6667 4056 6680 4062
rect 6551 4050 6558 4056
rect 6547 4042 6558 4050
rect 6608 4044 6615 4056
rect 6673 4050 6680 4056
rect 6497 4021 6505 4036
rect 6608 4037 6629 4044
rect 6587 4026 6593 4028
rect 6654 4026 6661 4032
rect 6497 4007 6513 4021
rect 6587 4020 6661 4026
rect 6497 3944 6505 4007
rect 6513 3993 6527 4007
rect 6519 3948 6533 3956
rect 6587 3948 6593 4020
rect 6654 4012 6661 4020
rect 6666 4004 6700 4012
rect 6694 3999 6700 4004
rect 6647 3986 6674 3993
rect 6553 3942 6593 3948
rect 6601 3948 6645 3954
rect 6553 3924 6559 3942
rect 6601 3934 6607 3948
rect 6713 3952 6719 4036
rect 6657 3944 6719 3952
rect 6577 3928 6607 3934
rect 6625 3930 6663 3938
rect 6655 3924 6663 3930
rect 6547 3884 6559 3918
rect 6605 3910 6627 3922
rect 6655 3910 6673 3924
rect 6601 3904 6613 3910
rect 6655 3904 6663 3910
rect 5462 3858 5474 3864
rect 5512 3858 5524 3864
rect 5591 3858 5603 3864
rect 5641 3858 5653 3864
rect 5707 3858 5719 3864
rect 5753 3858 5765 3864
rect 5811 3858 5823 3864
rect 5857 3858 5869 3864
rect 5951 3858 5963 3864
rect 5991 3858 6003 3864
rect 6037 3858 6049 3864
rect 6095 3858 6107 3864
rect 6141 3858 6153 3864
rect 6207 3858 6219 3864
rect 6277 3858 6289 3864
rect 6335 3858 6347 3864
rect 6381 3858 6393 3864
rect 6447 3858 6459 3864
rect 6517 3858 6529 3864
rect 6575 3858 6587 3864
rect 6621 3858 6633 3864
rect 6687 3858 6699 3864
rect 5287 3856 6736 3858
rect -62 3844 4 3856
rect -62 3842 2053 3844
rect -62 3378 -2 3842
rect 49 3836 61 3842
rect 129 3836 141 3842
rect 191 3836 203 3842
rect 231 3836 243 3842
rect 277 3836 289 3842
rect 335 3836 347 3842
rect 381 3836 393 3842
rect 447 3836 459 3842
rect 551 3836 563 3842
rect 611 3836 623 3842
rect 651 3836 663 3842
rect 31 3721 39 3756
rect 75 3750 83 3796
rect 57 3744 83 3750
rect 57 3738 60 3744
rect 31 3707 33 3721
rect 31 3664 39 3707
rect 53 3682 60 3738
rect 111 3721 119 3756
rect 155 3750 163 3796
rect 137 3744 163 3750
rect 137 3738 140 3744
rect 215 3741 223 3796
rect 307 3782 319 3816
rect 361 3790 373 3796
rect 415 3790 423 3796
rect 365 3778 387 3790
rect 415 3776 433 3790
rect 313 3758 319 3776
rect 337 3766 367 3772
rect 415 3770 423 3776
rect 111 3707 113 3721
rect 57 3676 60 3682
rect 57 3670 79 3676
rect 71 3644 79 3670
rect 111 3664 119 3707
rect 133 3682 140 3738
rect 137 3676 140 3682
rect 215 3678 223 3727
rect 137 3670 159 3676
rect 151 3644 159 3670
rect 199 3672 223 3678
rect 257 3693 265 3756
rect 279 3744 293 3752
rect 313 3752 353 3758
rect 273 3693 287 3707
rect 257 3679 273 3693
rect 347 3680 353 3752
rect 361 3752 367 3766
rect 385 3762 423 3770
rect 677 3836 689 3842
rect 717 3836 729 3842
rect 771 3836 783 3842
rect 811 3836 823 3842
rect 857 3836 869 3842
rect 915 3836 927 3842
rect 961 3836 973 3842
rect 1027 3836 1039 3842
rect 1097 3836 1109 3842
rect 1191 3836 1203 3842
rect 1231 3836 1243 3842
rect 1279 3836 1291 3842
rect 1391 3836 1403 3842
rect 1451 3836 1463 3842
rect 1491 3836 1503 3842
rect 571 3762 583 3764
rect 543 3756 583 3762
rect 597 3757 613 3763
rect 361 3746 405 3752
rect 417 3748 479 3756
rect 407 3707 434 3714
rect 454 3696 460 3701
rect 426 3688 460 3696
rect 414 3680 421 3688
rect 199 3664 211 3672
rect 257 3664 265 3679
rect 347 3674 421 3680
rect 347 3672 353 3674
rect 414 3668 421 3674
rect 307 3650 318 3658
rect 311 3644 318 3650
rect 368 3656 389 3663
rect 473 3664 479 3748
rect 514 3721 522 3756
rect 597 3743 603 3757
rect 587 3737 603 3743
rect 635 3741 643 3796
rect 697 3741 705 3796
rect 795 3741 803 3796
rect 887 3782 899 3816
rect 941 3790 953 3796
rect 995 3790 1003 3796
rect 945 3778 967 3790
rect 995 3776 1013 3790
rect 893 3758 899 3776
rect 917 3766 947 3772
rect 995 3770 1003 3776
rect 368 3644 375 3656
rect 433 3644 440 3650
rect 427 3638 440 3644
rect 514 3664 522 3707
rect 635 3678 643 3727
rect 619 3672 643 3678
rect 697 3678 705 3727
rect 795 3678 803 3727
rect 697 3672 721 3678
rect 619 3664 631 3672
rect 709 3664 721 3672
rect 514 3653 540 3664
rect 49 3618 61 3624
rect 129 3618 141 3624
rect 229 3618 241 3624
rect 279 3618 291 3624
rect 337 3618 349 3624
rect 385 3618 397 3624
rect 447 3618 459 3624
rect 518 3618 530 3624
rect 568 3618 580 3624
rect 649 3618 661 3624
rect 779 3672 803 3678
rect 837 3693 845 3756
rect 859 3744 873 3752
rect 893 3752 933 3758
rect 853 3693 867 3707
rect 837 3679 853 3693
rect 927 3680 933 3752
rect 941 3752 947 3766
rect 965 3762 1003 3770
rect 1077 3762 1089 3764
rect 1077 3756 1117 3762
rect 941 3746 985 3752
rect 997 3748 1059 3756
rect 987 3707 1014 3714
rect 1034 3696 1040 3701
rect 1006 3688 1040 3696
rect 994 3680 1001 3688
rect 779 3664 791 3672
rect 837 3664 845 3679
rect 927 3674 1001 3680
rect 927 3672 933 3674
rect 994 3668 1001 3674
rect 887 3650 898 3658
rect 891 3644 898 3650
rect 948 3656 969 3663
rect 1053 3664 1059 3748
rect 1138 3721 1146 3756
rect 1215 3741 1223 3796
rect 1257 3750 1265 3796
rect 1517 3836 1529 3842
rect 1557 3836 1569 3842
rect 1597 3836 1609 3842
rect 1697 3836 1709 3842
rect 1755 3836 1767 3842
rect 1801 3836 1813 3842
rect 1867 3836 1879 3842
rect 1931 3836 1943 3842
rect 1971 3836 1983 3842
rect 1411 3762 1423 3764
rect 1383 3756 1423 3762
rect 1257 3744 1283 3750
rect 1280 3738 1283 3744
rect 1138 3664 1146 3707
rect 1215 3678 1223 3727
rect 948 3644 955 3656
rect 1013 3644 1020 3650
rect 1007 3638 1020 3644
rect 1120 3653 1146 3664
rect 1199 3672 1223 3678
rect 1280 3682 1287 3738
rect 1301 3721 1309 3756
rect 1354 3721 1362 3756
rect 1475 3741 1483 3796
rect 1537 3741 1545 3796
rect 1620 3749 1637 3756
rect 1727 3782 1739 3816
rect 1781 3790 1793 3796
rect 1835 3790 1843 3796
rect 1785 3778 1807 3790
rect 1835 3776 1853 3790
rect 1733 3758 1739 3776
rect 1757 3766 1787 3772
rect 1835 3770 1843 3776
rect 1307 3707 1309 3721
rect 1280 3676 1283 3682
rect 1199 3664 1211 3672
rect 1261 3670 1283 3676
rect 1261 3644 1269 3670
rect 1301 3664 1309 3707
rect 1337 3667 1343 3693
rect 1354 3664 1362 3707
rect 1475 3678 1483 3727
rect 1459 3672 1483 3678
rect 1537 3678 1545 3727
rect 1620 3701 1627 3749
rect 1537 3672 1561 3678
rect 1459 3664 1471 3672
rect 1549 3664 1561 3672
rect 1354 3653 1380 3664
rect 679 3618 691 3624
rect 809 3618 821 3624
rect 859 3618 871 3624
rect 917 3618 929 3624
rect 965 3618 977 3624
rect 1027 3618 1039 3624
rect 1080 3618 1092 3624
rect 1130 3618 1142 3624
rect 1229 3618 1241 3624
rect 1279 3618 1291 3624
rect 1358 3618 1370 3624
rect 1408 3618 1420 3624
rect 1489 3618 1501 3624
rect 1620 3644 1627 3687
rect 1677 3693 1685 3756
rect 1699 3744 1713 3752
rect 1733 3752 1773 3758
rect 1693 3693 1707 3707
rect 1677 3679 1693 3693
rect 1767 3680 1773 3752
rect 1781 3752 1787 3766
rect 1805 3762 1843 3770
rect 1997 3836 2009 3842
rect 1781 3746 1825 3752
rect 1837 3748 1899 3756
rect 1827 3707 1854 3714
rect 1874 3696 1880 3701
rect 1846 3688 1880 3696
rect 1834 3680 1841 3688
rect 1677 3664 1685 3679
rect 1767 3674 1841 3680
rect 1767 3672 1773 3674
rect 1834 3668 1841 3674
rect 1727 3650 1738 3658
rect 1731 3644 1738 3650
rect 1788 3656 1809 3663
rect 1893 3664 1899 3748
rect 1955 3741 1963 3796
rect 2067 3842 2233 3844
rect 2077 3836 2089 3842
rect 2142 3836 2154 3842
rect 2192 3836 2204 3842
rect 2020 3749 2037 3756
rect 1955 3678 1963 3727
rect 2020 3701 2027 3749
rect 2096 3713 2104 3796
rect 2247 3842 6736 3844
rect 2256 3836 2268 3842
rect 2306 3836 2318 3842
rect 2391 3836 2403 3842
rect 2437 3836 2449 3842
rect 2531 3836 2543 3842
rect 2562 3836 2574 3842
rect 2612 3836 2624 3842
rect 2411 3762 2423 3764
rect 2383 3756 2423 3762
rect 2173 3721 2181 3756
rect 2279 3721 2287 3756
rect 2354 3721 2362 3756
rect 1788 3644 1795 3656
rect 1853 3644 1860 3650
rect 1847 3638 1860 3644
rect 1939 3672 1963 3678
rect 1939 3664 1951 3672
rect 2020 3644 2027 3687
rect 2096 3644 2104 3699
rect 2179 3685 2187 3707
rect 2273 3685 2281 3707
rect 2456 3713 2464 3796
rect 2516 3713 2524 3796
rect 2657 3836 2669 3842
rect 2697 3836 2709 3842
rect 2791 3836 2803 3842
rect 2678 3794 2689 3796
rect 2831 3836 2843 3842
rect 2871 3836 2883 3842
rect 2902 3836 2914 3842
rect 2952 3836 2964 3842
rect 2717 3794 2725 3796
rect 2678 3788 2725 3794
rect 2593 3721 2601 3756
rect 2718 3733 2725 3788
rect 2180 3678 2205 3685
rect 2137 3664 2189 3667
rect 1519 3618 1531 3624
rect 1597 3618 1609 3624
rect 1637 3618 1649 3624
rect 1699 3618 1711 3624
rect 1757 3618 1769 3624
rect 1805 3618 1817 3624
rect 1867 3618 1879 3624
rect 1969 3618 1981 3624
rect 1997 3618 2009 3624
rect 2037 3618 2049 3624
rect 2149 3658 2177 3664
rect 2197 3664 2205 3678
rect 2255 3678 2280 3685
rect 2255 3664 2263 3678
rect 2271 3664 2323 3667
rect 2283 3658 2311 3664
rect 2354 3664 2362 3707
rect 2354 3653 2380 3664
rect 2456 3644 2464 3699
rect 2487 3677 2503 3683
rect 2497 3667 2503 3677
rect 2516 3644 2524 3699
rect 2599 3685 2607 3707
rect 2716 3691 2724 3719
rect 2776 3713 2784 3796
rect 2807 3737 2823 3743
rect 2855 3741 2863 3796
rect 3002 3836 3014 3842
rect 3052 3836 3064 3842
rect 3117 3836 3129 3842
rect 3271 3836 3283 3842
rect 3331 3836 3343 3842
rect 3371 3836 3383 3842
rect 3097 3762 3109 3764
rect 3097 3756 3137 3762
rect 3223 3830 3251 3836
rect 3263 3758 3291 3764
rect 3411 3836 3423 3842
rect 3451 3836 3463 3842
rect 3501 3836 3513 3842
rect 3567 3836 3579 3842
rect 3613 3836 3625 3842
rect 3671 3836 3683 3842
rect 3731 3836 3743 3842
rect 3771 3836 3783 3842
rect 3871 3836 3883 3842
rect 3917 3836 3929 3842
rect 3977 3836 3989 3842
rect 4017 3836 4029 3842
rect 2817 3707 2823 3737
rect 2600 3678 2625 3685
rect 2557 3664 2609 3667
rect 2077 3618 2089 3624
rect 2157 3618 2169 3624
rect 2291 3618 2303 3624
rect 2358 3618 2370 3624
rect 2408 3618 2420 3624
rect 2569 3658 2597 3664
rect 2617 3664 2625 3678
rect 2694 3682 2724 3691
rect 2706 3680 2724 3682
rect 2776 3644 2784 3699
rect 2855 3678 2863 3727
rect 2933 3721 2941 3756
rect 3033 3721 3041 3756
rect 3158 3721 3166 3756
rect 3232 3750 3244 3756
rect 3232 3744 3259 3750
rect 3253 3721 3259 3744
rect 3355 3741 3363 3796
rect 3435 3741 3443 3796
rect 3537 3790 3545 3796
rect 3587 3790 3599 3796
rect 3527 3776 3545 3790
rect 3573 3778 3595 3790
rect 3641 3782 3653 3816
rect 3537 3770 3545 3776
rect 3537 3762 3575 3770
rect 3593 3766 3623 3772
rect 3481 3748 3543 3756
rect 2939 3685 2947 3707
rect 3039 3685 3047 3707
rect 2940 3678 2965 3685
rect 3040 3678 3065 3685
rect 2839 3672 2863 3678
rect 2839 3664 2851 3672
rect 2897 3664 2949 3667
rect 2909 3658 2937 3664
rect 2957 3664 2965 3678
rect 2997 3664 3049 3667
rect 3009 3658 3037 3664
rect 3057 3664 3065 3678
rect 3158 3664 3166 3707
rect 3260 3664 3267 3707
rect 3355 3678 3363 3727
rect 3435 3678 3443 3727
rect 3339 3672 3363 3678
rect 3419 3672 3443 3678
rect 3339 3664 3351 3672
rect 3419 3664 3431 3672
rect 3481 3664 3487 3748
rect 3593 3752 3599 3766
rect 3641 3758 3647 3776
rect 3555 3746 3599 3752
rect 3607 3752 3647 3758
rect 3526 3707 3553 3714
rect 3500 3696 3506 3701
rect 3500 3688 3534 3696
rect 3539 3680 3546 3688
rect 3607 3680 3613 3752
rect 3667 3744 3681 3752
rect 3673 3693 3687 3707
rect 3695 3693 3703 3756
rect 3755 3741 3763 3796
rect 3823 3830 3851 3836
rect 3863 3758 3891 3764
rect 4062 3836 4074 3842
rect 4112 3836 4124 3842
rect 4181 3836 4193 3842
rect 4247 3836 4259 3842
rect 4293 3836 4305 3842
rect 4351 3836 4363 3842
rect 4397 3836 4409 3842
rect 4437 3836 4449 3842
rect 3832 3750 3844 3756
rect 3832 3744 3859 3750
rect 3539 3674 3613 3680
rect 3687 3679 3703 3693
rect 3539 3668 3546 3674
rect 3607 3672 3613 3674
rect 3140 3653 3166 3664
rect 2437 3618 2449 3624
rect 2531 3618 2543 3624
rect 2577 3618 2589 3624
rect 2658 3618 2670 3624
rect 2791 3618 2803 3624
rect 2869 3618 2881 3624
rect 2917 3618 2929 3624
rect 3017 3618 3029 3624
rect 3100 3618 3112 3624
rect 3150 3618 3162 3624
rect 3571 3656 3592 3663
rect 3695 3664 3703 3679
rect 3755 3678 3763 3727
rect 3853 3721 3859 3744
rect 3520 3644 3527 3650
rect 3585 3644 3592 3656
rect 3642 3650 3653 3658
rect 3642 3644 3649 3650
rect 3520 3638 3533 3644
rect 3739 3672 3763 3678
rect 3739 3664 3751 3672
rect 3860 3664 3867 3707
rect 3936 3713 3944 3796
rect 3997 3741 4005 3796
rect 4217 3790 4225 3796
rect 4267 3790 4279 3796
rect 4207 3776 4225 3790
rect 4253 3778 4275 3790
rect 4321 3782 4333 3816
rect 4217 3770 4225 3776
rect 4217 3762 4255 3770
rect 4273 3766 4303 3772
rect 3232 3618 3244 3624
rect 3288 3618 3300 3624
rect 3369 3618 3381 3624
rect 3449 3618 3461 3624
rect 3501 3618 3513 3624
rect 3563 3618 3575 3624
rect 3611 3618 3623 3624
rect 3669 3618 3681 3624
rect 3769 3618 3781 3624
rect 3936 3644 3944 3699
rect 3997 3678 4005 3727
rect 4093 3721 4101 3756
rect 4161 3748 4223 3756
rect 4099 3685 4107 3707
rect 4100 3678 4125 3685
rect 3997 3672 4021 3678
rect 4009 3664 4021 3672
rect 3832 3618 3844 3624
rect 3888 3618 3900 3624
rect 4057 3664 4109 3667
rect 4069 3658 4097 3664
rect 4117 3664 4125 3678
rect 4161 3664 4167 3748
rect 4273 3752 4279 3766
rect 4321 3758 4327 3776
rect 4235 3746 4279 3752
rect 4287 3752 4327 3758
rect 4206 3707 4233 3714
rect 4180 3696 4186 3701
rect 4180 3688 4214 3696
rect 4219 3680 4226 3688
rect 4287 3680 4293 3752
rect 4491 3836 4503 3842
rect 4531 3836 4543 3842
rect 4571 3836 4583 3842
rect 4611 3836 4623 3842
rect 4651 3836 4663 3842
rect 4691 3836 4703 3842
rect 4731 3836 4743 3842
rect 4781 3836 4793 3842
rect 4847 3836 4859 3842
rect 4893 3836 4905 3842
rect 4951 3836 4963 3842
rect 5002 3836 5014 3842
rect 5052 3836 5064 3842
rect 4347 3744 4361 3752
rect 4353 3693 4367 3707
rect 4375 3693 4383 3756
rect 4417 3741 4425 3796
rect 4515 3741 4523 3796
rect 4817 3790 4825 3796
rect 4867 3790 4879 3796
rect 4807 3776 4825 3790
rect 4853 3778 4875 3790
rect 4921 3782 4933 3816
rect 4817 3770 4825 3776
rect 4817 3762 4855 3770
rect 4873 3766 4903 3772
rect 4591 3750 4603 3756
rect 4631 3750 4643 3756
rect 4671 3750 4683 3756
rect 4711 3750 4723 3756
rect 4585 3742 4603 3750
rect 4618 3742 4643 3750
rect 4658 3742 4683 3750
rect 4697 3742 4723 3750
rect 4761 3748 4823 3756
rect 4219 3674 4293 3680
rect 4367 3679 4383 3693
rect 4219 3668 4226 3674
rect 4287 3672 4293 3674
rect 4251 3656 4272 3663
rect 4375 3664 4383 3679
rect 4417 3678 4425 3727
rect 4515 3678 4523 3727
rect 4585 3713 4592 3742
rect 4587 3699 4592 3713
rect 4417 3672 4441 3678
rect 4429 3664 4441 3672
rect 4200 3644 4207 3650
rect 4265 3644 4272 3656
rect 4322 3650 4333 3658
rect 4322 3644 4329 3650
rect 4200 3638 4213 3644
rect 4499 3672 4523 3678
rect 4585 3678 4592 3699
rect 4618 3696 4626 3742
rect 4658 3696 4666 3742
rect 4697 3696 4705 3742
rect 4610 3684 4626 3696
rect 4650 3684 4666 3696
rect 4690 3684 4705 3696
rect 4618 3678 4626 3684
rect 4658 3678 4666 3684
rect 4697 3678 4705 3684
rect 4499 3664 4511 3672
rect 4585 3671 4604 3678
rect 4586 3670 4604 3671
rect 4618 3670 4644 3678
rect 4658 3670 4683 3678
rect 4697 3670 4724 3678
rect 4592 3664 4604 3670
rect 4632 3664 4644 3670
rect 4671 3664 4683 3670
rect 4712 3664 4724 3670
rect 4761 3664 4767 3748
rect 4873 3752 4879 3766
rect 4921 3758 4927 3776
rect 4835 3746 4879 3752
rect 4887 3752 4927 3758
rect 4806 3707 4833 3714
rect 4780 3696 4786 3701
rect 4780 3688 4814 3696
rect 4819 3680 4826 3688
rect 4887 3680 4893 3752
rect 5111 3836 5123 3842
rect 5151 3836 5163 3842
rect 5191 3836 5203 3842
rect 5231 3836 5243 3842
rect 5291 3836 5303 3842
rect 5317 3836 5329 3842
rect 5357 3836 5369 3842
rect 5397 3836 5409 3842
rect 5437 3836 5449 3842
rect 5477 3836 5489 3842
rect 5537 3836 5549 3842
rect 5595 3836 5607 3842
rect 5641 3836 5653 3842
rect 5707 3836 5719 3842
rect 5791 3836 5803 3842
rect 4947 3744 4961 3752
rect 4953 3693 4967 3707
rect 4975 3693 4983 3756
rect 5033 3721 5041 3756
rect 5135 3741 5143 3796
rect 5177 3757 5193 3763
rect 4819 3674 4893 3680
rect 4967 3679 4983 3693
rect 5039 3685 5047 3707
rect 4819 3668 4826 3674
rect 4887 3672 4893 3674
rect 3917 3618 3929 3624
rect 3979 3618 3991 3624
rect 4077 3618 4089 3624
rect 4181 3618 4193 3624
rect 4243 3618 4255 3624
rect 4291 3618 4303 3624
rect 4349 3618 4361 3624
rect 4399 3618 4411 3624
rect 4529 3618 4541 3624
rect 4851 3656 4872 3663
rect 4975 3664 4983 3679
rect 5040 3678 5065 3685
rect 5135 3678 5143 3727
rect 4800 3644 4807 3650
rect 4865 3644 4872 3656
rect 4922 3650 4933 3658
rect 4922 3644 4929 3650
rect 4800 3638 4813 3644
rect 4997 3664 5049 3667
rect 5009 3658 5037 3664
rect 5057 3664 5065 3678
rect 5119 3672 5143 3678
rect 5177 3683 5183 3757
rect 5215 3741 5223 3796
rect 5167 3677 5183 3683
rect 5215 3678 5223 3727
rect 5199 3672 5223 3678
rect 5257 3683 5263 3753
rect 5276 3713 5284 3796
rect 5567 3782 5579 3816
rect 5621 3790 5633 3796
rect 5675 3790 5683 3796
rect 5625 3778 5647 3790
rect 5675 3776 5693 3790
rect 5573 3758 5579 3776
rect 5597 3766 5627 3772
rect 5675 3770 5683 3776
rect 5337 3750 5349 3756
rect 5377 3750 5389 3756
rect 5417 3750 5429 3756
rect 5457 3750 5469 3756
rect 5337 3742 5363 3750
rect 5377 3742 5402 3750
rect 5417 3742 5442 3750
rect 5457 3742 5475 3750
rect 5247 3677 5263 3683
rect 5119 3664 5131 3672
rect 5199 3664 5211 3672
rect 5276 3644 5284 3699
rect 5355 3696 5363 3742
rect 5394 3696 5402 3742
rect 5434 3696 5442 3742
rect 5468 3713 5475 3742
rect 5468 3699 5473 3713
rect 5355 3684 5370 3696
rect 5394 3684 5410 3696
rect 5434 3684 5450 3696
rect 5355 3678 5363 3684
rect 5394 3678 5402 3684
rect 5434 3678 5442 3684
rect 5468 3678 5475 3699
rect 5336 3670 5363 3678
rect 5377 3670 5402 3678
rect 5416 3670 5442 3678
rect 5456 3671 5475 3678
rect 5517 3693 5525 3756
rect 5539 3744 5553 3752
rect 5573 3752 5613 3758
rect 5533 3693 5547 3707
rect 5517 3679 5533 3693
rect 5607 3680 5613 3752
rect 5621 3752 5627 3766
rect 5645 3762 5683 3770
rect 5817 3836 5829 3842
rect 5857 3836 5869 3842
rect 5897 3836 5909 3842
rect 5937 3836 5949 3842
rect 6011 3836 6023 3842
rect 6037 3836 6049 3842
rect 6171 3836 6183 3842
rect 6217 3836 6229 3842
rect 6317 3836 6329 3842
rect 6375 3836 6387 3842
rect 6421 3836 6433 3842
rect 6487 3836 6499 3842
rect 6542 3836 6554 3842
rect 6592 3836 6604 3842
rect 5621 3746 5665 3752
rect 5677 3748 5739 3756
rect 5667 3707 5694 3714
rect 5714 3696 5720 3701
rect 5686 3688 5720 3696
rect 5674 3680 5681 3688
rect 5456 3670 5474 3671
rect 5336 3664 5348 3670
rect 5377 3664 5389 3670
rect 5416 3664 5428 3670
rect 5456 3664 5468 3670
rect 5517 3664 5525 3679
rect 5607 3674 5681 3680
rect 5607 3672 5613 3674
rect 4571 3618 4583 3624
rect 4611 3618 4623 3624
rect 4651 3618 4663 3624
rect 4691 3618 4703 3624
rect 4731 3618 4743 3624
rect 4781 3618 4793 3624
rect 4843 3618 4855 3624
rect 4891 3618 4903 3624
rect 4949 3618 4961 3624
rect 5017 3618 5029 3624
rect 5149 3618 5161 3624
rect 5229 3618 5241 3624
rect 5291 3618 5303 3624
rect 5674 3668 5681 3674
rect 5567 3650 5578 3658
rect 5571 3644 5578 3650
rect 5628 3656 5649 3663
rect 5733 3664 5739 3748
rect 5776 3713 5784 3796
rect 5837 3741 5845 3796
rect 5917 3741 5925 3796
rect 5628 3644 5635 3656
rect 5693 3644 5700 3650
rect 5687 3638 5700 3644
rect 5776 3644 5784 3699
rect 5837 3678 5845 3727
rect 5917 3678 5925 3727
rect 5996 3713 6004 3796
rect 6060 3749 6077 3756
rect 6197 3762 6209 3764
rect 6197 3756 6237 3762
rect 6347 3782 6359 3816
rect 6401 3790 6413 3796
rect 6455 3790 6463 3796
rect 6405 3778 6427 3790
rect 6455 3776 6473 3790
rect 6353 3758 6359 3776
rect 6377 3766 6407 3772
rect 6455 3770 6463 3776
rect 6143 3749 6160 3756
rect 6060 3701 6067 3749
rect 5837 3672 5861 3678
rect 5917 3672 5941 3678
rect 5849 3664 5861 3672
rect 5929 3664 5941 3672
rect 5317 3618 5329 3624
rect 5357 3618 5369 3624
rect 5397 3618 5409 3624
rect 5437 3618 5449 3624
rect 5477 3618 5489 3624
rect 5539 3618 5551 3624
rect 5597 3618 5609 3624
rect 5645 3618 5657 3624
rect 5707 3618 5719 3624
rect 5791 3618 5803 3624
rect 5996 3644 6004 3699
rect 6060 3644 6067 3687
rect 6153 3701 6160 3749
rect 6258 3721 6266 3756
rect 6153 3644 6160 3687
rect 6258 3664 6266 3707
rect 5819 3618 5831 3624
rect 5899 3618 5911 3624
rect 6011 3618 6023 3624
rect 6037 3618 6049 3624
rect 6077 3618 6089 3624
rect 6131 3618 6143 3624
rect 6171 3618 6183 3624
rect 6240 3653 6266 3664
rect 6297 3693 6305 3756
rect 6319 3744 6333 3752
rect 6353 3752 6393 3758
rect 6313 3693 6327 3707
rect 6297 3679 6313 3693
rect 6387 3680 6393 3752
rect 6401 3752 6407 3766
rect 6425 3762 6463 3770
rect 6637 3836 6649 3842
rect 6677 3836 6689 3842
rect 6401 3746 6445 3752
rect 6457 3748 6519 3756
rect 6447 3707 6474 3714
rect 6494 3696 6500 3701
rect 6466 3688 6500 3696
rect 6454 3680 6461 3688
rect 6297 3664 6305 3679
rect 6387 3674 6461 3680
rect 6387 3672 6393 3674
rect 6454 3668 6461 3674
rect 6347 3650 6358 3658
rect 6351 3644 6358 3650
rect 6408 3656 6429 3663
rect 6513 3664 6519 3748
rect 6573 3721 6581 3756
rect 6657 3741 6665 3796
rect 6579 3685 6587 3707
rect 6580 3678 6605 3685
rect 6408 3644 6415 3656
rect 6473 3644 6480 3650
rect 6467 3638 6480 3644
rect 6537 3664 6589 3667
rect 6549 3658 6577 3664
rect 6597 3664 6605 3678
rect 6657 3678 6665 3727
rect 6657 3672 6681 3678
rect 6669 3664 6681 3672
rect 6200 3618 6212 3624
rect 6250 3618 6262 3624
rect 6319 3618 6331 3624
rect 6377 3618 6389 3624
rect 6425 3618 6437 3624
rect 6487 3618 6499 3624
rect 6557 3618 6569 3624
rect 6639 3618 6651 3624
rect 6742 3618 6802 4082
rect 4 3616 6802 3618
rect 6736 3604 6802 3616
rect 4 3602 6802 3604
rect 49 3596 61 3602
rect 119 3596 131 3602
rect 177 3596 189 3602
rect 225 3596 237 3602
rect 287 3596 299 3602
rect 339 3596 351 3602
rect 439 3596 451 3602
rect 518 3596 530 3602
rect 568 3596 580 3602
rect 649 3596 661 3602
rect 709 3596 721 3602
rect 779 3596 791 3602
rect 839 3596 851 3602
rect 949 3596 961 3602
rect 1031 3596 1043 3602
rect 1089 3596 1101 3602
rect 1169 3596 1181 3602
rect 1239 3596 1251 3602
rect 1297 3596 1309 3602
rect 1345 3596 1357 3602
rect 1407 3596 1419 3602
rect 1471 3596 1483 3602
rect 1511 3596 1523 3602
rect 1559 3596 1571 3602
rect 1617 3596 1629 3602
rect 1665 3596 1677 3602
rect 1727 3596 1739 3602
rect 1821 3596 1833 3602
rect 1911 3596 1923 3602
rect 1991 3596 2003 3602
rect 2037 3596 2049 3602
rect 2077 3596 2089 3602
rect 2151 3596 2163 3602
rect 2221 3596 2233 3602
rect 2291 3596 2303 3602
rect 2331 3596 2343 3602
rect 2379 3596 2391 3602
rect 2437 3596 2449 3602
rect 2485 3596 2497 3602
rect 2547 3596 2559 3602
rect 2597 3596 2609 3602
rect 2637 3596 2649 3602
rect 2697 3596 2709 3602
rect 2811 3596 2823 3602
rect 2889 3596 2901 3602
rect 2937 3596 2949 3602
rect 3020 3596 3032 3602
rect 3070 3596 3082 3602
rect 31 3513 39 3556
rect 71 3550 79 3576
rect 57 3544 79 3550
rect 267 3576 280 3582
rect 151 3570 158 3576
rect 147 3562 158 3570
rect 208 3564 215 3576
rect 273 3570 280 3576
rect 57 3538 60 3544
rect 31 3499 33 3513
rect 31 3464 39 3499
rect 53 3482 60 3538
rect 97 3541 105 3556
rect 208 3557 229 3564
rect 187 3546 193 3548
rect 254 3546 261 3552
rect 97 3527 113 3541
rect 187 3540 261 3546
rect 57 3476 60 3482
rect 57 3470 83 3476
rect 75 3424 83 3470
rect 97 3464 105 3527
rect 113 3513 127 3527
rect 119 3468 133 3476
rect 187 3468 193 3540
rect 254 3532 261 3540
rect 266 3524 300 3532
rect 294 3519 300 3524
rect 247 3506 274 3513
rect 153 3462 193 3468
rect 201 3468 245 3474
rect 153 3444 159 3462
rect 201 3454 207 3468
rect 313 3472 319 3556
rect 369 3548 381 3556
rect 357 3542 381 3548
rect 421 3550 429 3576
rect 514 3556 540 3567
rect 421 3544 443 3550
rect 357 3493 365 3542
rect 440 3538 443 3544
rect 440 3482 447 3538
rect 461 3513 469 3556
rect 514 3513 522 3556
rect 619 3548 631 3556
rect 619 3542 643 3548
rect 467 3499 469 3513
rect 257 3464 319 3472
rect 177 3448 207 3454
rect 225 3450 263 3458
rect 255 3444 263 3450
rect 147 3404 159 3438
rect 205 3430 227 3442
rect 255 3430 273 3444
rect 201 3424 213 3430
rect 255 3424 263 3430
rect 357 3424 365 3479
rect 440 3476 443 3482
rect 417 3470 443 3476
rect 417 3424 425 3470
rect 461 3464 469 3499
rect 514 3464 522 3499
rect 635 3493 643 3542
rect 691 3513 699 3556
rect 731 3550 739 3576
rect 717 3544 739 3550
rect 761 3550 769 3576
rect 761 3544 783 3550
rect 717 3538 720 3544
rect 691 3499 693 3513
rect 543 3458 583 3464
rect 571 3456 583 3458
rect 635 3424 643 3479
rect 691 3464 699 3499
rect 713 3482 720 3538
rect 780 3538 783 3544
rect 717 3476 720 3482
rect 780 3482 787 3538
rect 801 3513 809 3556
rect 869 3548 881 3556
rect 857 3542 881 3548
rect 807 3499 809 3513
rect 780 3476 783 3482
rect 717 3470 743 3476
rect 735 3424 743 3470
rect 757 3470 783 3476
rect 757 3424 765 3470
rect 801 3464 809 3499
rect 857 3493 865 3542
rect 931 3513 939 3556
rect 971 3550 979 3576
rect 957 3544 979 3550
rect 957 3538 960 3544
rect 931 3499 933 3513
rect 857 3424 865 3479
rect 931 3464 939 3499
rect 953 3482 960 3538
rect 1016 3521 1024 3576
rect 1071 3513 1079 3556
rect 1111 3550 1119 3576
rect 1097 3544 1119 3550
rect 1097 3538 1100 3544
rect 957 3476 960 3482
rect 957 3470 983 3476
rect 975 3424 983 3470
rect 1016 3424 1024 3507
rect 1071 3499 1073 3513
rect 1071 3464 1079 3499
rect 1093 3482 1100 3538
rect 1151 3513 1159 3556
rect 1191 3550 1199 3576
rect 1177 3544 1199 3550
rect 1387 3576 1400 3582
rect 1271 3570 1278 3576
rect 1267 3562 1278 3570
rect 1328 3564 1335 3576
rect 1393 3570 1400 3576
rect 1177 3538 1180 3544
rect 1151 3499 1153 3513
rect 1097 3476 1100 3482
rect 1097 3470 1123 3476
rect 1115 3424 1123 3470
rect 1151 3464 1159 3499
rect 1173 3482 1180 3538
rect 1217 3541 1225 3556
rect 1328 3557 1349 3564
rect 1307 3546 1313 3548
rect 1374 3546 1381 3552
rect 1217 3527 1233 3541
rect 1307 3540 1381 3546
rect 1177 3476 1180 3482
rect 1177 3470 1203 3476
rect 1195 3424 1203 3470
rect 1217 3464 1225 3527
rect 1233 3513 1247 3527
rect 1239 3468 1253 3476
rect 1307 3468 1313 3540
rect 1374 3532 1381 3540
rect 1386 3524 1420 3532
rect 1414 3519 1420 3524
rect 1367 3506 1394 3513
rect 1273 3462 1313 3468
rect 1321 3468 1365 3474
rect 1273 3444 1279 3462
rect 1321 3454 1327 3468
rect 1433 3472 1439 3556
rect 1493 3533 1500 3576
rect 1707 3576 1720 3582
rect 1591 3570 1598 3576
rect 1587 3562 1598 3570
rect 1648 3564 1655 3576
rect 1713 3570 1720 3576
rect 1537 3541 1545 3556
rect 1648 3557 1669 3564
rect 1627 3546 1633 3548
rect 1694 3546 1701 3552
rect 1537 3527 1553 3541
rect 1627 3540 1701 3546
rect 1377 3464 1439 3472
rect 1493 3471 1500 3519
rect 1297 3448 1327 3454
rect 1345 3450 1383 3458
rect 1375 3444 1383 3450
rect 1267 3404 1279 3438
rect 1325 3430 1347 3442
rect 1375 3430 1393 3444
rect 1321 3424 1333 3430
rect 1375 3424 1383 3430
rect 1483 3464 1500 3471
rect 1537 3464 1545 3527
rect 1553 3513 1567 3527
rect 1559 3468 1573 3476
rect 49 3378 61 3384
rect 117 3378 129 3384
rect 175 3378 187 3384
rect 221 3378 233 3384
rect 287 3378 299 3384
rect 337 3378 349 3384
rect 377 3378 389 3384
rect 439 3378 451 3384
rect 551 3378 563 3384
rect 611 3378 623 3384
rect 651 3378 663 3384
rect 709 3378 721 3384
rect 779 3378 791 3384
rect 837 3378 849 3384
rect 877 3378 889 3384
rect 949 3378 961 3384
rect 1031 3378 1043 3384
rect 1089 3378 1101 3384
rect 1169 3378 1181 3384
rect 1237 3378 1249 3384
rect 1295 3378 1307 3384
rect 1341 3378 1353 3384
rect 1407 3378 1419 3384
rect -62 3376 1453 3378
rect 1627 3468 1633 3540
rect 1694 3532 1701 3540
rect 1706 3524 1740 3532
rect 1734 3519 1740 3524
rect 1687 3506 1714 3513
rect 1593 3462 1633 3468
rect 1641 3468 1685 3474
rect 1593 3444 1599 3462
rect 1641 3454 1647 3468
rect 1753 3472 1759 3556
rect 1697 3464 1759 3472
rect 1791 3556 1801 3566
rect 1791 3513 1799 3556
rect 1851 3546 1863 3556
rect 1825 3538 1863 3546
rect 1791 3499 1793 3513
rect 1791 3464 1799 3499
rect 1617 3448 1647 3454
rect 1665 3450 1703 3458
rect 1695 3444 1703 3450
rect 1587 3404 1599 3438
rect 1645 3430 1667 3442
rect 1695 3430 1713 3444
rect 1641 3424 1653 3430
rect 1695 3424 1703 3430
rect 1834 3424 1842 3538
rect 1896 3521 1904 3576
rect 1955 3542 1963 3556
rect 1983 3556 2011 3562
rect 1971 3553 2023 3556
rect 1955 3535 1980 3542
rect 1973 3513 1981 3535
rect 2060 3533 2067 3576
rect 1896 3424 1904 3507
rect 2136 3521 2144 3576
rect 2191 3556 2201 3566
rect 1979 3464 1987 3499
rect 2060 3471 2067 3519
rect 2191 3513 2199 3556
rect 2251 3546 2263 3556
rect 2225 3538 2263 3546
rect 2060 3464 2077 3471
rect 1511 3378 1523 3384
rect 1557 3378 1569 3384
rect 1615 3378 1627 3384
rect 1661 3378 1673 3384
rect 1727 3378 1739 3384
rect 1807 3378 1819 3384
rect 1851 3378 1863 3384
rect 1911 3378 1923 3384
rect 1956 3378 1968 3384
rect 2006 3378 2018 3384
rect 2136 3424 2144 3507
rect 2191 3499 2193 3513
rect 2191 3464 2199 3499
rect 2234 3424 2242 3538
rect 2313 3533 2320 3576
rect 2527 3576 2540 3582
rect 2411 3570 2418 3576
rect 2407 3562 2418 3570
rect 2468 3564 2475 3576
rect 2533 3570 2540 3576
rect 2357 3541 2365 3556
rect 2468 3557 2489 3564
rect 2447 3546 2453 3548
rect 2514 3546 2521 3552
rect 2357 3527 2373 3541
rect 2447 3540 2521 3546
rect 2313 3471 2320 3519
rect 2303 3464 2320 3471
rect 2357 3464 2365 3527
rect 2373 3513 2387 3527
rect 2379 3468 2393 3476
rect 2447 3468 2453 3540
rect 2514 3532 2521 3540
rect 2526 3524 2560 3532
rect 2554 3519 2560 3524
rect 2507 3506 2534 3513
rect 2413 3462 2453 3468
rect 2461 3468 2505 3474
rect 2413 3444 2419 3462
rect 2461 3454 2467 3468
rect 2573 3472 2579 3556
rect 2620 3533 2627 3576
rect 2689 3556 2717 3562
rect 2677 3553 2729 3556
rect 2737 3542 2745 3556
rect 2720 3535 2745 3542
rect 2517 3464 2579 3472
rect 2620 3471 2627 3519
rect 2719 3513 2727 3535
rect 2796 3521 2804 3576
rect 2929 3556 2957 3562
rect 2859 3548 2871 3556
rect 2917 3553 2969 3556
rect 3117 3596 3129 3602
rect 3212 3596 3224 3602
rect 3268 3596 3280 3602
rect 3331 3596 3343 3602
rect 3379 3596 3391 3602
rect 3437 3596 3449 3602
rect 3485 3596 3497 3602
rect 3547 3596 3559 3602
rect 3632 3596 3644 3602
rect 3688 3596 3700 3602
rect 3739 3596 3751 3602
rect 3797 3596 3809 3602
rect 3845 3596 3857 3602
rect 3907 3596 3919 3602
rect 3991 3596 4003 3602
rect 4039 3596 4051 3602
rect 4097 3596 4109 3602
rect 4145 3596 4157 3602
rect 4207 3596 4219 3602
rect 4291 3596 4303 3602
rect 4351 3596 4363 3602
rect 3060 3556 3086 3567
rect 2859 3542 2883 3548
rect 2977 3542 2985 3556
rect 2620 3464 2637 3471
rect 2713 3464 2721 3499
rect 2437 3448 2467 3454
rect 2485 3450 2523 3458
rect 2515 3444 2523 3450
rect 2407 3404 2419 3438
rect 2465 3430 2487 3442
rect 2515 3430 2533 3444
rect 2461 3424 2473 3430
rect 2515 3424 2523 3430
rect 2796 3424 2804 3507
rect 2875 3493 2883 3542
rect 2960 3535 2985 3542
rect 2959 3513 2967 3535
rect 3078 3513 3086 3556
rect 3136 3513 3144 3556
rect 3240 3513 3247 3556
rect 3316 3521 3324 3576
rect 3527 3576 3540 3582
rect 3411 3570 3418 3576
rect 3407 3562 3418 3570
rect 3468 3564 3475 3576
rect 3533 3570 3540 3576
rect 3357 3541 3365 3556
rect 3468 3557 3489 3564
rect 3887 3576 3900 3582
rect 3771 3570 3778 3576
rect 3767 3562 3778 3570
rect 3828 3564 3835 3576
rect 3893 3570 3900 3576
rect 3447 3546 3453 3548
rect 3514 3546 3521 3552
rect 3357 3527 3373 3541
rect 3447 3540 3521 3546
rect 2875 3424 2883 3479
rect 2953 3464 2961 3499
rect 3078 3464 3086 3499
rect 3136 3464 3144 3499
rect 3233 3476 3239 3499
rect 3212 3470 3239 3476
rect 3212 3464 3224 3470
rect 2037 3378 2049 3384
rect 2151 3378 2163 3384
rect 2207 3378 2219 3384
rect 2251 3378 2263 3384
rect 2331 3378 2343 3384
rect 2377 3378 2389 3384
rect 2435 3378 2447 3384
rect 2481 3378 2493 3384
rect 2547 3378 2559 3384
rect 2597 3378 2609 3384
rect 2682 3378 2694 3384
rect 2732 3378 2744 3384
rect 2811 3378 2823 3384
rect 2851 3378 2863 3384
rect 2891 3378 2903 3384
rect 3017 3458 3057 3464
rect 3017 3456 3029 3458
rect 3203 3384 3231 3390
rect 3243 3456 3271 3462
rect 3316 3424 3324 3507
rect 3357 3464 3365 3527
rect 3373 3513 3387 3527
rect 3379 3468 3393 3476
rect 3447 3468 3453 3540
rect 3514 3532 3521 3540
rect 3526 3524 3560 3532
rect 3554 3519 3560 3524
rect 3507 3506 3534 3513
rect 3413 3462 3453 3468
rect 3461 3468 3505 3474
rect 3413 3444 3419 3462
rect 3461 3454 3467 3468
rect 3573 3472 3579 3556
rect 3660 3513 3667 3556
rect 3717 3541 3725 3556
rect 3828 3557 3849 3564
rect 3807 3546 3813 3548
rect 3874 3546 3881 3552
rect 3717 3527 3733 3541
rect 3807 3540 3881 3546
rect 3653 3476 3659 3499
rect 3517 3464 3579 3472
rect 3632 3470 3659 3476
rect 3632 3464 3644 3470
rect 3717 3464 3725 3527
rect 3733 3513 3747 3527
rect 3739 3468 3753 3476
rect 3437 3448 3467 3454
rect 3485 3450 3523 3458
rect 3515 3444 3523 3450
rect 3407 3404 3419 3438
rect 3465 3430 3487 3442
rect 3515 3430 3533 3444
rect 3461 3424 3473 3430
rect 3515 3424 3523 3430
rect 3623 3384 3651 3390
rect 3663 3456 3691 3462
rect 3807 3468 3813 3540
rect 3874 3532 3881 3540
rect 3886 3524 3920 3532
rect 3914 3519 3920 3524
rect 3867 3506 3894 3513
rect 3773 3462 3813 3468
rect 3821 3468 3865 3474
rect 3773 3444 3779 3462
rect 3821 3454 3827 3468
rect 3933 3472 3939 3556
rect 3976 3521 3984 3576
rect 4187 3576 4200 3582
rect 4071 3570 4078 3576
rect 4067 3562 4078 3570
rect 4128 3564 4135 3576
rect 4193 3570 4200 3576
rect 4017 3541 4025 3556
rect 4128 3557 4149 3564
rect 4379 3596 4391 3602
rect 4481 3596 4493 3602
rect 4543 3596 4555 3602
rect 4591 3596 4603 3602
rect 4649 3596 4661 3602
rect 4731 3596 4743 3602
rect 4779 3596 4791 3602
rect 4837 3596 4849 3602
rect 4885 3596 4897 3602
rect 4947 3596 4959 3602
rect 5032 3596 5044 3602
rect 5088 3596 5100 3602
rect 5151 3596 5163 3602
rect 5199 3596 5211 3602
rect 5257 3596 5269 3602
rect 5305 3596 5317 3602
rect 5367 3596 5379 3602
rect 5439 3596 5451 3602
rect 5497 3596 5509 3602
rect 5545 3596 5557 3602
rect 5607 3596 5619 3602
rect 5677 3596 5689 3602
rect 5777 3596 5789 3602
rect 5891 3596 5903 3602
rect 4107 3546 4113 3548
rect 4174 3546 4181 3552
rect 4017 3527 4033 3541
rect 4107 3540 4181 3546
rect 3877 3464 3939 3472
rect 3797 3448 3827 3454
rect 3845 3450 3883 3458
rect 3875 3444 3883 3450
rect 3767 3404 3779 3438
rect 3825 3430 3847 3442
rect 3875 3430 3893 3444
rect 3821 3424 3833 3430
rect 3875 3424 3883 3430
rect 3976 3424 3984 3507
rect 4017 3464 4025 3527
rect 4033 3513 4047 3527
rect 4039 3468 4053 3476
rect 4107 3468 4113 3540
rect 4174 3532 4181 3540
rect 4186 3524 4220 3532
rect 4214 3519 4220 3524
rect 4167 3506 4194 3513
rect 4073 3462 4113 3468
rect 4121 3468 4165 3474
rect 4073 3444 4079 3462
rect 4121 3454 4127 3468
rect 4233 3472 4239 3556
rect 4276 3521 4284 3576
rect 4336 3521 4344 3576
rect 4409 3548 4421 3556
rect 4397 3542 4421 3548
rect 4500 3576 4513 3582
rect 4500 3570 4507 3576
rect 4565 3564 4572 3576
rect 4177 3464 4239 3472
rect 4097 3448 4127 3454
rect 4145 3450 4183 3458
rect 4175 3444 4183 3450
rect 4067 3404 4079 3438
rect 4125 3430 4147 3442
rect 4175 3430 4193 3444
rect 4121 3424 4133 3430
rect 4175 3424 4183 3430
rect 4276 3424 4284 3507
rect 4336 3424 4344 3507
rect 4397 3493 4405 3542
rect 4397 3424 4405 3479
rect 4461 3472 4467 3556
rect 4551 3557 4572 3564
rect 4622 3570 4629 3576
rect 4622 3562 4633 3570
rect 4519 3546 4526 3552
rect 4587 3546 4593 3548
rect 4519 3540 4593 3546
rect 4675 3541 4683 3556
rect 4519 3532 4526 3540
rect 4480 3524 4514 3532
rect 4480 3519 4486 3524
rect 4506 3506 4533 3513
rect 4461 3464 4523 3472
rect 4535 3468 4579 3474
rect 2922 3378 2934 3384
rect 2972 3378 2984 3384
rect 3037 3378 3049 3384
rect 3117 3378 3129 3384
rect 3251 3378 3263 3384
rect 3331 3378 3343 3384
rect 3377 3378 3389 3384
rect 3435 3378 3447 3384
rect 3481 3378 3493 3384
rect 3547 3378 3559 3384
rect 3671 3378 3683 3384
rect 3737 3378 3749 3384
rect 3795 3378 3807 3384
rect 3841 3378 3853 3384
rect 3907 3378 3919 3384
rect 3991 3378 4003 3384
rect 4037 3378 4049 3384
rect 4095 3378 4107 3384
rect 4141 3378 4153 3384
rect 4207 3378 4219 3384
rect 4291 3378 4303 3384
rect 4351 3378 4363 3384
rect 4517 3450 4555 3458
rect 4573 3454 4579 3468
rect 4587 3468 4593 3540
rect 4667 3527 4683 3541
rect 4653 3513 4667 3527
rect 4587 3462 4627 3468
rect 4647 3468 4661 3476
rect 4675 3464 4683 3527
rect 4716 3521 4724 3576
rect 4927 3576 4940 3582
rect 4811 3570 4818 3576
rect 4807 3562 4818 3570
rect 4868 3564 4875 3576
rect 4933 3570 4940 3576
rect 4757 3541 4765 3556
rect 4868 3557 4889 3564
rect 4847 3546 4853 3548
rect 4914 3546 4921 3552
rect 4757 3527 4773 3541
rect 4847 3540 4921 3546
rect 4517 3444 4525 3450
rect 4573 3448 4603 3454
rect 4621 3444 4627 3462
rect 4507 3430 4525 3444
rect 4553 3430 4575 3442
rect 4517 3424 4525 3430
rect 4567 3424 4579 3430
rect 4621 3404 4633 3438
rect 4716 3424 4724 3507
rect 4757 3464 4765 3527
rect 4773 3513 4787 3527
rect 4779 3468 4793 3476
rect 4847 3468 4853 3540
rect 4914 3532 4921 3540
rect 4926 3524 4960 3532
rect 4954 3519 4960 3524
rect 4907 3506 4934 3513
rect 4813 3462 4853 3468
rect 4861 3468 4905 3474
rect 4813 3444 4819 3462
rect 4861 3454 4867 3468
rect 4973 3472 4979 3556
rect 5060 3513 5067 3556
rect 5136 3521 5144 3576
rect 5347 3576 5360 3582
rect 5231 3570 5238 3576
rect 5227 3562 5238 3570
rect 5288 3564 5295 3576
rect 5353 3570 5360 3576
rect 5177 3541 5185 3556
rect 5288 3557 5309 3564
rect 5267 3546 5273 3548
rect 5334 3546 5341 3552
rect 5177 3527 5193 3541
rect 5267 3540 5341 3546
rect 5053 3476 5059 3499
rect 4917 3464 4979 3472
rect 5032 3470 5059 3476
rect 5032 3464 5044 3470
rect 4837 3448 4867 3454
rect 4885 3450 4923 3458
rect 4915 3444 4923 3450
rect 4807 3404 4819 3438
rect 4865 3430 4887 3442
rect 4915 3430 4933 3444
rect 4861 3424 4873 3430
rect 4915 3424 4923 3430
rect 5023 3384 5051 3390
rect 5063 3456 5091 3462
rect 5136 3424 5144 3507
rect 5177 3464 5185 3527
rect 5193 3513 5207 3527
rect 5199 3468 5213 3476
rect 5267 3468 5273 3540
rect 5334 3532 5341 3540
rect 5346 3524 5380 3532
rect 5374 3519 5380 3524
rect 5327 3506 5354 3513
rect 5233 3462 5273 3468
rect 5281 3468 5325 3474
rect 5233 3444 5239 3462
rect 5281 3454 5287 3468
rect 5393 3472 5399 3556
rect 5337 3464 5399 3472
rect 5257 3448 5287 3454
rect 5305 3450 5343 3458
rect 5335 3444 5343 3450
rect 5227 3404 5239 3438
rect 5285 3430 5307 3442
rect 5335 3430 5353 3444
rect 5281 3424 5293 3430
rect 5335 3424 5343 3430
rect 5587 3576 5600 3582
rect 5471 3570 5478 3576
rect 5467 3562 5478 3570
rect 5528 3564 5535 3576
rect 5593 3570 5600 3576
rect 5417 3541 5425 3556
rect 5528 3557 5549 3564
rect 5507 3546 5513 3548
rect 5574 3546 5581 3552
rect 5417 3527 5433 3541
rect 5507 3540 5581 3546
rect 5417 3464 5425 3527
rect 5433 3513 5447 3527
rect 5439 3468 5453 3476
rect 5507 3468 5513 3540
rect 5574 3532 5581 3540
rect 5586 3524 5620 3532
rect 5614 3519 5620 3524
rect 5567 3506 5594 3513
rect 5473 3462 5513 3468
rect 5521 3468 5565 3474
rect 5473 3444 5479 3462
rect 5521 3454 5527 3468
rect 5633 3472 5639 3556
rect 5669 3556 5697 3562
rect 5657 3553 5709 3556
rect 5769 3556 5797 3562
rect 5717 3542 5725 3556
rect 5757 3553 5809 3556
rect 5952 3596 5964 3602
rect 6008 3596 6020 3602
rect 5817 3542 5825 3556
rect 5700 3535 5725 3542
rect 5800 3535 5825 3542
rect 5699 3513 5707 3535
rect 5799 3513 5807 3535
rect 5876 3521 5884 3576
rect 5907 3557 5923 3563
rect 5577 3464 5639 3472
rect 5693 3464 5701 3499
rect 5793 3464 5801 3499
rect 5497 3448 5527 3454
rect 5545 3450 5583 3458
rect 5575 3444 5583 3450
rect 5467 3404 5479 3438
rect 5525 3430 5547 3442
rect 5575 3430 5593 3444
rect 5521 3424 5533 3430
rect 5575 3424 5583 3430
rect 4377 3378 4389 3384
rect 4417 3378 4429 3384
rect 4481 3378 4493 3384
rect 4547 3378 4559 3384
rect 4593 3378 4605 3384
rect 4651 3378 4663 3384
rect 4731 3378 4743 3384
rect 4777 3378 4789 3384
rect 4835 3378 4847 3384
rect 4881 3378 4893 3384
rect 4947 3378 4959 3384
rect 5071 3378 5083 3384
rect 5151 3378 5163 3384
rect 5197 3378 5209 3384
rect 5255 3378 5267 3384
rect 5301 3378 5313 3384
rect 5367 3378 5379 3384
rect 5437 3378 5449 3384
rect 5495 3378 5507 3384
rect 5541 3378 5553 3384
rect 5607 3378 5619 3384
rect 5662 3378 5674 3384
rect 5712 3378 5724 3384
rect 5876 3424 5884 3507
rect 5917 3483 5923 3557
rect 6039 3596 6051 3602
rect 6151 3596 6163 3602
rect 6195 3596 6209 3602
rect 6237 3596 6249 3602
rect 6391 3596 6403 3602
rect 6439 3596 6451 3602
rect 6497 3596 6509 3602
rect 6545 3596 6557 3602
rect 6607 3596 6619 3602
rect 5980 3513 5987 3556
rect 6069 3548 6081 3556
rect 6057 3542 6081 3548
rect 5907 3477 5923 3483
rect 5973 3476 5979 3499
rect 6057 3493 6065 3542
rect 6136 3521 6144 3576
rect 6222 3570 6229 3576
rect 6262 3570 6269 3576
rect 6222 3564 6294 3570
rect 6286 3521 6294 3564
rect 6376 3521 6384 3576
rect 6587 3576 6600 3582
rect 6471 3570 6478 3576
rect 6467 3562 6478 3570
rect 6528 3564 6535 3576
rect 6593 3570 6600 3576
rect 6417 3541 6425 3556
rect 6528 3557 6549 3564
rect 6507 3546 6513 3548
rect 6574 3546 6581 3552
rect 5952 3470 5979 3476
rect 5952 3464 5964 3470
rect 5943 3384 5971 3390
rect 5983 3456 6011 3462
rect 6057 3424 6065 3479
rect 6136 3424 6144 3507
rect 6286 3507 6293 3521
rect 6417 3527 6433 3541
rect 6507 3540 6581 3546
rect 6286 3472 6294 3507
rect 6286 3464 6309 3472
rect 6177 3450 6229 3456
rect 6177 3444 6189 3450
rect 6217 3444 6229 3450
rect 6237 3452 6293 3454
rect 6237 3448 6281 3452
rect 6237 3444 6249 3448
rect 6229 3384 6257 3390
rect 6301 3448 6309 3464
rect 6281 3390 6293 3392
rect 6376 3424 6384 3507
rect 6417 3464 6425 3527
rect 6433 3513 6447 3527
rect 6439 3468 6453 3476
rect 6321 3390 6333 3392
rect 6281 3384 6333 3390
rect 6507 3468 6513 3540
rect 6574 3532 6581 3540
rect 6586 3524 6620 3532
rect 6614 3519 6620 3524
rect 6567 3506 6594 3513
rect 6473 3462 6513 3468
rect 6521 3468 6565 3474
rect 6473 3444 6479 3462
rect 6521 3454 6527 3468
rect 6633 3472 6639 3556
rect 6577 3464 6639 3472
rect 6497 3448 6527 3454
rect 6545 3450 6583 3458
rect 6575 3444 6583 3450
rect 6467 3404 6479 3438
rect 6525 3430 6547 3442
rect 6575 3430 6593 3444
rect 6521 3424 6533 3430
rect 6575 3424 6583 3430
rect 5762 3378 5774 3384
rect 5812 3378 5824 3384
rect 5891 3378 5903 3384
rect 5991 3378 6003 3384
rect 6037 3378 6049 3384
rect 6077 3378 6089 3384
rect 6151 3378 6163 3384
rect 6197 3378 6209 3384
rect 6391 3378 6403 3384
rect 6437 3378 6449 3384
rect 6495 3378 6507 3384
rect 6541 3378 6553 3384
rect 6607 3378 6619 3384
rect 1467 3376 6736 3378
rect -62 3364 4 3376
rect -62 3362 1153 3364
rect -62 2898 -2 3362
rect 49 3356 61 3362
rect 117 3356 129 3362
rect 175 3356 187 3362
rect 221 3356 233 3362
rect 287 3356 299 3362
rect 337 3356 349 3362
rect 377 3356 389 3362
rect 471 3356 483 3362
rect 531 3356 543 3362
rect 571 3356 583 3362
rect 31 3241 39 3276
rect 75 3270 83 3316
rect 57 3264 83 3270
rect 147 3302 159 3336
rect 201 3310 213 3316
rect 255 3310 263 3316
rect 205 3298 227 3310
rect 255 3296 273 3310
rect 153 3278 159 3296
rect 177 3286 207 3292
rect 255 3290 263 3296
rect 57 3258 60 3264
rect 31 3227 33 3241
rect 31 3184 39 3227
rect 53 3202 60 3258
rect 57 3196 60 3202
rect 97 3213 105 3276
rect 119 3264 133 3272
rect 153 3272 193 3278
rect 113 3213 127 3227
rect 97 3199 113 3213
rect 187 3200 193 3272
rect 201 3272 207 3286
rect 225 3282 263 3290
rect 201 3266 245 3272
rect 257 3268 319 3276
rect 247 3227 274 3234
rect 294 3216 300 3221
rect 266 3208 300 3216
rect 254 3200 261 3208
rect 57 3190 79 3196
rect 71 3164 79 3190
rect 97 3184 105 3199
rect 187 3194 261 3200
rect 187 3192 193 3194
rect 254 3188 261 3194
rect 147 3170 158 3178
rect 151 3164 158 3170
rect 208 3176 229 3183
rect 313 3184 319 3268
rect 357 3261 365 3316
rect 597 3356 609 3362
rect 657 3356 669 3362
rect 697 3356 709 3362
rect 757 3356 769 3362
rect 797 3356 809 3362
rect 491 3282 503 3284
rect 463 3276 503 3282
rect 517 3277 533 3283
rect 357 3198 365 3247
rect 434 3241 442 3276
rect 517 3263 523 3277
rect 507 3257 523 3263
rect 555 3261 563 3316
rect 357 3192 381 3198
rect 369 3184 381 3192
rect 208 3164 215 3176
rect 273 3164 280 3170
rect 267 3158 280 3164
rect 434 3184 442 3227
rect 555 3198 563 3247
rect 616 3233 624 3316
rect 678 3314 689 3316
rect 856 3356 868 3362
rect 906 3356 918 3362
rect 717 3314 725 3316
rect 678 3308 725 3314
rect 539 3192 563 3198
rect 539 3184 551 3192
rect 434 3173 460 3184
rect 616 3164 624 3219
rect 637 3207 643 3273
rect 718 3253 725 3308
rect 777 3261 785 3316
rect 937 3356 949 3362
rect 997 3356 1009 3362
rect 1082 3356 1094 3362
rect 1132 3356 1144 3362
rect 716 3211 724 3239
rect 49 3138 61 3144
rect 119 3138 131 3144
rect 177 3138 189 3144
rect 225 3138 237 3144
rect 287 3138 299 3144
rect 339 3138 351 3144
rect 438 3138 450 3144
rect 488 3138 500 3144
rect 569 3138 581 3144
rect 694 3202 724 3211
rect 706 3200 724 3202
rect 777 3198 785 3247
rect 879 3241 887 3276
rect 873 3205 881 3227
rect 956 3233 964 3316
rect 1167 3362 2373 3364
rect 1182 3356 1194 3362
rect 1232 3356 1244 3362
rect 1277 3356 1289 3362
rect 1317 3356 1329 3362
rect 1377 3356 1389 3362
rect 1435 3356 1447 3362
rect 1481 3356 1493 3362
rect 1547 3356 1559 3362
rect 1627 3356 1639 3362
rect 1671 3356 1683 3362
rect 1751 3356 1763 3362
rect 1831 3356 1843 3362
rect 1871 3356 1883 3362
rect 1917 3356 1929 3362
rect 2021 3356 2033 3362
rect 2087 3356 2099 3362
rect 2133 3356 2145 3362
rect 2191 3356 2203 3362
rect 2237 3356 2249 3362
rect 2277 3356 2289 3362
rect 1020 3269 1037 3276
rect 1020 3221 1027 3269
rect 1113 3241 1121 3276
rect 1213 3241 1221 3276
rect 1297 3261 1305 3316
rect 1407 3302 1419 3336
rect 1461 3310 1473 3316
rect 1515 3310 1523 3316
rect 1465 3298 1487 3310
rect 1515 3296 1533 3310
rect 1413 3278 1419 3296
rect 1437 3286 1467 3292
rect 1515 3290 1523 3296
rect 855 3198 880 3205
rect 777 3192 801 3198
rect 789 3184 801 3192
rect 855 3184 863 3198
rect 871 3184 923 3187
rect 883 3178 911 3184
rect 956 3164 964 3219
rect 1020 3164 1027 3207
rect 1119 3205 1127 3227
rect 1219 3205 1227 3227
rect 1120 3198 1145 3205
rect 1220 3198 1245 3205
rect 1077 3184 1129 3187
rect 1089 3178 1117 3184
rect 1137 3184 1145 3198
rect 1177 3184 1229 3187
rect 1189 3178 1217 3184
rect 1237 3184 1245 3198
rect 1297 3198 1305 3247
rect 1357 3213 1365 3276
rect 1379 3264 1393 3272
rect 1413 3272 1453 3278
rect 1373 3213 1387 3227
rect 1357 3199 1373 3213
rect 1447 3200 1453 3272
rect 1461 3272 1467 3286
rect 1485 3282 1523 3290
rect 1461 3266 1505 3272
rect 1517 3268 1579 3276
rect 1507 3227 1534 3234
rect 1554 3216 1560 3221
rect 1526 3208 1560 3216
rect 1514 3200 1521 3208
rect 1297 3192 1321 3198
rect 1309 3184 1321 3192
rect 1357 3184 1365 3199
rect 1447 3194 1521 3200
rect 1447 3192 1453 3194
rect 1514 3188 1521 3194
rect 1407 3170 1418 3178
rect 1411 3164 1418 3170
rect 1468 3176 1489 3183
rect 1573 3184 1579 3268
rect 1468 3164 1475 3176
rect 1533 3164 1540 3170
rect 1527 3158 1540 3164
rect 1611 3241 1619 3276
rect 1611 3227 1613 3241
rect 1611 3184 1619 3227
rect 1654 3202 1662 3316
rect 1771 3282 1783 3284
rect 1743 3276 1783 3282
rect 1815 3314 1823 3316
rect 1851 3314 1862 3316
rect 1815 3308 1862 3314
rect 1714 3241 1722 3276
rect 1815 3253 1822 3308
rect 1897 3282 1909 3284
rect 1897 3276 1937 3282
rect 2057 3310 2065 3316
rect 2107 3310 2119 3316
rect 2047 3296 2065 3310
rect 2093 3298 2115 3310
rect 2161 3302 2173 3336
rect 2057 3290 2065 3296
rect 2057 3282 2095 3290
rect 2113 3286 2143 3292
rect 1958 3241 1966 3276
rect 2001 3268 2063 3276
rect 1645 3194 1683 3202
rect 1671 3184 1683 3194
rect 1611 3174 1621 3184
rect 1714 3184 1722 3227
rect 1816 3211 1824 3239
rect 1816 3202 1846 3211
rect 1816 3200 1834 3202
rect 1714 3173 1740 3184
rect 1958 3184 1966 3227
rect 597 3138 609 3144
rect 658 3138 670 3144
rect 759 3138 771 3144
rect 891 3138 903 3144
rect 937 3138 949 3144
rect 997 3138 1009 3144
rect 1037 3138 1049 3144
rect 1097 3138 1109 3144
rect 1197 3138 1209 3144
rect 1279 3138 1291 3144
rect 1379 3138 1391 3144
rect 1437 3138 1449 3144
rect 1485 3138 1497 3144
rect 1547 3138 1559 3144
rect 1641 3138 1653 3144
rect 1718 3138 1730 3144
rect 1768 3138 1780 3144
rect 1870 3138 1882 3144
rect 1940 3173 1966 3184
rect 2001 3184 2007 3268
rect 2113 3272 2119 3286
rect 2161 3278 2167 3296
rect 2075 3266 2119 3272
rect 2127 3272 2167 3278
rect 2046 3227 2073 3234
rect 2020 3216 2026 3221
rect 2020 3208 2054 3216
rect 2059 3200 2066 3208
rect 2127 3200 2133 3272
rect 2317 3356 2329 3362
rect 2187 3264 2201 3272
rect 2193 3213 2207 3227
rect 2215 3213 2223 3276
rect 2257 3261 2265 3316
rect 2387 3362 3433 3364
rect 2451 3356 2463 3362
rect 2340 3269 2357 3276
rect 2496 3356 2508 3362
rect 2546 3356 2558 3362
rect 2577 3356 2589 3362
rect 2661 3356 2673 3362
rect 2727 3356 2739 3362
rect 2773 3356 2785 3362
rect 2831 3356 2843 3362
rect 2877 3356 2889 3362
rect 2917 3356 2929 3362
rect 2423 3269 2440 3276
rect 2059 3194 2133 3200
rect 2207 3199 2223 3213
rect 2059 3188 2066 3194
rect 2127 3192 2133 3194
rect 2091 3176 2112 3183
rect 2215 3184 2223 3199
rect 2257 3198 2265 3247
rect 2340 3221 2347 3269
rect 2257 3192 2281 3198
rect 2269 3184 2281 3192
rect 2040 3164 2047 3170
rect 2105 3164 2112 3176
rect 2162 3170 2173 3178
rect 2162 3164 2169 3170
rect 2040 3158 2053 3164
rect 2340 3164 2347 3207
rect 2433 3221 2440 3269
rect 2519 3241 2527 3276
rect 2433 3164 2440 3207
rect 2513 3205 2521 3227
rect 2596 3233 2604 3316
rect 2697 3310 2705 3316
rect 2747 3310 2759 3316
rect 2687 3296 2705 3310
rect 2733 3298 2755 3310
rect 2801 3302 2813 3336
rect 2697 3290 2705 3296
rect 2697 3282 2735 3290
rect 2753 3286 2783 3292
rect 2641 3268 2703 3276
rect 2495 3198 2520 3205
rect 2495 3184 2503 3198
rect 1900 3138 1912 3144
rect 1950 3138 1962 3144
rect 2021 3138 2033 3144
rect 2083 3138 2095 3144
rect 2131 3138 2143 3144
rect 2189 3138 2201 3144
rect 2239 3138 2251 3144
rect 2317 3138 2329 3144
rect 2357 3138 2369 3144
rect 2511 3184 2563 3187
rect 2523 3178 2551 3184
rect 2596 3164 2604 3219
rect 2641 3184 2647 3268
rect 2753 3272 2759 3286
rect 2801 3278 2807 3296
rect 2715 3266 2759 3272
rect 2767 3272 2807 3278
rect 2686 3227 2713 3234
rect 2660 3216 2666 3221
rect 2660 3208 2694 3216
rect 2699 3200 2706 3208
rect 2767 3200 2773 3272
rect 2971 3356 2983 3362
rect 3011 3356 3023 3362
rect 3056 3356 3068 3362
rect 3106 3356 3118 3362
rect 2827 3264 2841 3272
rect 2833 3213 2847 3227
rect 2855 3213 2863 3276
rect 2897 3261 2905 3316
rect 2995 3261 3003 3316
rect 3037 3297 3053 3303
rect 2699 3194 2773 3200
rect 2847 3199 2863 3213
rect 2699 3188 2706 3194
rect 2767 3192 2773 3194
rect 2731 3176 2752 3183
rect 2855 3184 2863 3199
rect 2897 3198 2905 3247
rect 2995 3198 3003 3247
rect 3037 3247 3043 3297
rect 3151 3356 3163 3362
rect 3191 3356 3203 3362
rect 3251 3356 3263 3362
rect 3296 3356 3308 3362
rect 3346 3356 3358 3362
rect 3079 3241 3087 3276
rect 3175 3261 3183 3316
rect 3073 3205 3081 3227
rect 2897 3192 2921 3198
rect 2909 3184 2921 3192
rect 2680 3164 2687 3170
rect 2745 3164 2752 3176
rect 2802 3170 2813 3178
rect 2802 3164 2809 3170
rect 2680 3158 2693 3164
rect 2979 3192 3003 3198
rect 3055 3198 3080 3205
rect 3175 3198 3183 3247
rect 3236 3233 3244 3316
rect 3377 3356 3389 3362
rect 3447 3362 4473 3364
rect 3491 3356 3503 3362
rect 3571 3356 3583 3362
rect 3671 3356 3683 3362
rect 3717 3356 3729 3362
rect 3775 3356 3787 3362
rect 3821 3356 3833 3362
rect 3887 3356 3899 3362
rect 3957 3356 3969 3362
rect 4131 3356 4143 3362
rect 4201 3356 4213 3362
rect 4267 3356 4279 3362
rect 4313 3356 4325 3362
rect 4371 3356 4383 3362
rect 4417 3356 4429 3362
rect 3267 3257 3283 3263
rect 3277 3223 3283 3257
rect 3319 3241 3327 3276
rect 2979 3184 2991 3192
rect 3055 3184 3063 3198
rect 3159 3192 3183 3198
rect 3071 3184 3123 3187
rect 3083 3178 3111 3184
rect 3159 3184 3171 3192
rect 3236 3164 3244 3219
rect 3277 3217 3293 3223
rect 3313 3205 3321 3227
rect 3396 3233 3404 3316
rect 3591 3282 3603 3284
rect 3563 3276 3603 3282
rect 3747 3302 3759 3336
rect 3801 3310 3813 3316
rect 3855 3310 3863 3316
rect 3805 3298 3827 3310
rect 3855 3296 3873 3310
rect 3753 3278 3759 3296
rect 3777 3286 3807 3292
rect 3855 3290 3863 3296
rect 3463 3269 3480 3276
rect 3473 3221 3480 3269
rect 3534 3241 3542 3276
rect 3643 3269 3660 3276
rect 3587 3257 3623 3263
rect 3295 3198 3320 3205
rect 3295 3184 3303 3198
rect 3311 3184 3363 3187
rect 3323 3178 3351 3184
rect 3396 3164 3404 3219
rect 3473 3164 3480 3207
rect 3534 3184 3542 3227
rect 3617 3203 3623 3257
rect 3653 3221 3660 3269
rect 3697 3213 3705 3276
rect 3719 3264 3733 3272
rect 3753 3272 3793 3278
rect 3713 3213 3727 3227
rect 3617 3197 3633 3203
rect 3534 3173 3560 3184
rect 2411 3138 2423 3144
rect 2451 3138 2463 3144
rect 2531 3138 2543 3144
rect 2577 3138 2589 3144
rect 2661 3138 2673 3144
rect 2723 3138 2735 3144
rect 2771 3138 2783 3144
rect 2829 3138 2841 3144
rect 2879 3138 2891 3144
rect 3009 3138 3021 3144
rect 3091 3138 3103 3144
rect 3189 3138 3201 3144
rect 3251 3138 3263 3144
rect 3331 3138 3343 3144
rect 3377 3138 3389 3144
rect 3451 3138 3463 3144
rect 3491 3138 3503 3144
rect 3653 3164 3660 3207
rect 3697 3199 3713 3213
rect 3787 3200 3793 3272
rect 3801 3272 3807 3286
rect 3825 3282 3863 3290
rect 3949 3278 3977 3284
rect 3989 3350 4017 3356
rect 4083 3350 4111 3356
rect 4123 3278 4151 3284
rect 4237 3310 4245 3316
rect 4287 3310 4299 3316
rect 4227 3296 4245 3310
rect 4273 3298 4295 3310
rect 4341 3302 4353 3336
rect 4237 3290 4245 3296
rect 4237 3282 4275 3290
rect 4293 3286 4323 3292
rect 3801 3266 3845 3272
rect 3857 3268 3919 3276
rect 3996 3270 4008 3276
rect 3847 3227 3874 3234
rect 3894 3216 3900 3221
rect 3866 3208 3900 3216
rect 3854 3200 3861 3208
rect 3697 3184 3705 3199
rect 3787 3194 3861 3200
rect 3787 3192 3793 3194
rect 3538 3138 3550 3144
rect 3588 3138 3600 3144
rect 3854 3188 3861 3194
rect 3747 3170 3758 3178
rect 3751 3164 3758 3170
rect 3808 3176 3829 3183
rect 3913 3184 3919 3268
rect 3981 3264 4008 3270
rect 4092 3270 4104 3276
rect 4092 3264 4119 3270
rect 3981 3241 3987 3264
rect 4113 3241 4119 3264
rect 4181 3268 4243 3276
rect 3973 3184 3980 3227
rect 4120 3184 4127 3227
rect 4181 3184 4187 3268
rect 4293 3272 4299 3286
rect 4341 3278 4347 3296
rect 4255 3266 4299 3272
rect 4307 3272 4347 3278
rect 4226 3227 4253 3234
rect 4200 3216 4206 3221
rect 4200 3208 4234 3216
rect 4239 3200 4246 3208
rect 4307 3200 4313 3272
rect 4487 3362 6736 3364
rect 4517 3356 4529 3362
rect 4617 3356 4629 3362
rect 4697 3356 4709 3362
rect 4777 3356 4789 3362
rect 4857 3356 4869 3362
rect 4977 3356 4989 3362
rect 5077 3356 5089 3362
rect 5135 3356 5147 3362
rect 5181 3356 5193 3362
rect 5247 3356 5259 3362
rect 5331 3356 5343 3362
rect 4509 3278 4537 3284
rect 4549 3350 4577 3356
rect 4367 3264 4381 3272
rect 4373 3213 4387 3227
rect 4395 3213 4403 3276
rect 4440 3269 4457 3276
rect 4556 3270 4568 3276
rect 4440 3221 4447 3269
rect 4541 3264 4568 3270
rect 4640 3269 4657 3276
rect 4720 3269 4737 3276
rect 4239 3194 4313 3200
rect 4387 3199 4403 3213
rect 4477 3207 4483 3253
rect 4541 3241 4547 3264
rect 4239 3188 4246 3194
rect 4307 3192 4313 3194
rect 3808 3164 3815 3176
rect 3873 3164 3880 3170
rect 3867 3158 3880 3164
rect 3631 3138 3643 3144
rect 3671 3138 3683 3144
rect 3719 3138 3731 3144
rect 3777 3138 3789 3144
rect 3825 3138 3837 3144
rect 3887 3138 3899 3144
rect 3940 3138 3952 3144
rect 3996 3138 4008 3144
rect 4271 3176 4292 3183
rect 4395 3184 4403 3199
rect 4220 3164 4227 3170
rect 4285 3164 4292 3176
rect 4342 3170 4353 3178
rect 4342 3164 4349 3170
rect 4220 3158 4233 3164
rect 4440 3164 4447 3207
rect 4533 3184 4540 3227
rect 4640 3221 4647 3269
rect 4720 3221 4727 3269
rect 4796 3233 4804 3316
rect 4849 3278 4877 3284
rect 4889 3350 4917 3356
rect 4957 3282 4969 3284
rect 4957 3276 4997 3282
rect 5107 3302 5119 3336
rect 5161 3310 5173 3316
rect 5215 3310 5223 3316
rect 5165 3298 5187 3310
rect 5215 3296 5233 3310
rect 5113 3278 5119 3296
rect 5137 3286 5167 3292
rect 5215 3290 5223 3296
rect 4896 3270 4908 3276
rect 4881 3264 4908 3270
rect 4881 3241 4887 3264
rect 5018 3241 5026 3276
rect 4092 3138 4104 3144
rect 4148 3138 4160 3144
rect 4201 3138 4213 3144
rect 4263 3138 4275 3144
rect 4311 3138 4323 3144
rect 4369 3138 4381 3144
rect 4417 3138 4429 3144
rect 4457 3138 4469 3144
rect 4640 3164 4647 3207
rect 4667 3197 4693 3203
rect 4720 3164 4727 3207
rect 4796 3164 4804 3219
rect 4873 3184 4880 3227
rect 5018 3184 5026 3227
rect 4500 3138 4512 3144
rect 4556 3138 4568 3144
rect 4617 3138 4629 3144
rect 4657 3138 4669 3144
rect 4697 3138 4709 3144
rect 4737 3138 4749 3144
rect 4777 3138 4789 3144
rect 4840 3138 4852 3144
rect 4896 3138 4908 3144
rect 5000 3173 5026 3184
rect 5057 3213 5065 3276
rect 5079 3264 5093 3272
rect 5113 3272 5153 3278
rect 5073 3213 5087 3227
rect 5057 3199 5073 3213
rect 5147 3200 5153 3272
rect 5161 3272 5167 3286
rect 5185 3282 5223 3290
rect 5377 3348 5389 3362
rect 5437 3356 5449 3362
rect 5511 3356 5523 3362
rect 5561 3356 5573 3362
rect 5627 3356 5639 3362
rect 5673 3356 5685 3362
rect 5731 3356 5743 3362
rect 5796 3356 5808 3362
rect 5846 3356 5858 3362
rect 5911 3356 5923 3362
rect 5991 3356 6003 3362
rect 6042 3356 6054 3362
rect 6092 3356 6104 3362
rect 5161 3266 5205 3272
rect 5217 3268 5279 3276
rect 5207 3227 5234 3234
rect 5254 3216 5260 3221
rect 5226 3208 5260 3216
rect 5214 3200 5221 3208
rect 5057 3184 5065 3199
rect 5147 3194 5221 3200
rect 5147 3192 5153 3194
rect 5214 3188 5221 3194
rect 5107 3170 5118 3178
rect 5111 3164 5118 3170
rect 5168 3176 5189 3183
rect 5273 3184 5279 3268
rect 5316 3233 5324 3316
rect 5363 3274 5369 3308
rect 5419 3284 5421 3286
rect 5407 3280 5421 3284
rect 5363 3268 5404 3274
rect 5168 3164 5175 3176
rect 5233 3164 5240 3170
rect 5227 3158 5240 3164
rect 5316 3164 5324 3219
rect 5395 3250 5404 3268
rect 5395 3200 5404 3238
rect 5415 3233 5421 3280
rect 5496 3233 5504 3316
rect 5597 3310 5605 3316
rect 5647 3310 5659 3316
rect 5587 3296 5605 3310
rect 5633 3298 5655 3310
rect 5701 3302 5713 3336
rect 5597 3290 5605 3296
rect 5597 3282 5635 3290
rect 5653 3286 5683 3292
rect 5541 3268 5603 3276
rect 5362 3194 5404 3200
rect 5362 3172 5369 3194
rect 5415 3188 5421 3219
rect 5407 3184 5421 3188
rect 5419 3182 5421 3184
rect 5496 3164 5504 3219
rect 5541 3184 5547 3268
rect 5653 3272 5659 3286
rect 5701 3278 5707 3296
rect 5615 3266 5659 3272
rect 5667 3272 5707 3278
rect 5586 3227 5613 3234
rect 5560 3216 5566 3221
rect 5560 3208 5594 3216
rect 5599 3200 5606 3208
rect 5667 3200 5673 3272
rect 5727 3264 5741 3272
rect 5733 3213 5747 3227
rect 5755 3213 5763 3276
rect 5819 3241 5827 3276
rect 5599 3194 5673 3200
rect 5747 3199 5763 3213
rect 5813 3205 5821 3227
rect 5896 3233 5904 3316
rect 6011 3282 6023 3284
rect 5983 3276 6023 3282
rect 6151 3356 6163 3362
rect 6191 3356 6203 3362
rect 6271 3356 6283 3362
rect 6331 3356 6343 3362
rect 6371 3356 6383 3362
rect 6117 3277 6133 3283
rect 5954 3241 5962 3276
rect 6073 3241 6081 3276
rect 5599 3188 5606 3194
rect 5667 3192 5673 3194
rect 4960 3138 4972 3144
rect 5010 3138 5022 3144
rect 5079 3138 5091 3144
rect 5137 3138 5149 3144
rect 5185 3138 5197 3144
rect 5247 3138 5259 3144
rect 5331 3138 5343 3144
rect 5377 3138 5389 3152
rect 5437 3138 5449 3152
rect 5631 3176 5652 3183
rect 5755 3184 5763 3199
rect 5795 3198 5820 3205
rect 5795 3184 5803 3198
rect 5580 3164 5587 3170
rect 5645 3164 5652 3176
rect 5702 3170 5713 3178
rect 5702 3164 5709 3170
rect 5580 3158 5593 3164
rect 5811 3184 5863 3187
rect 5823 3178 5851 3184
rect 5896 3164 5904 3219
rect 5954 3184 5962 3227
rect 6079 3205 6087 3227
rect 6117 3207 6123 3277
rect 6175 3261 6183 3316
rect 6402 3356 6414 3362
rect 6452 3356 6464 3362
rect 6517 3356 6529 3362
rect 6575 3356 6587 3362
rect 6621 3356 6633 3362
rect 6687 3356 6699 3362
rect 6291 3282 6303 3284
rect 6263 3276 6303 3282
rect 6080 3198 6105 3205
rect 6037 3184 6089 3187
rect 5954 3173 5980 3184
rect 5511 3138 5523 3144
rect 5561 3138 5573 3144
rect 5623 3138 5635 3144
rect 5671 3138 5683 3144
rect 5729 3138 5741 3144
rect 5831 3138 5843 3144
rect 5911 3138 5923 3144
rect 6049 3178 6077 3184
rect 6097 3184 6105 3198
rect 6175 3198 6183 3247
rect 6234 3241 6242 3276
rect 6355 3261 6363 3316
rect 6547 3302 6559 3336
rect 6601 3310 6613 3316
rect 6655 3310 6663 3316
rect 6605 3298 6627 3310
rect 6655 3296 6673 3310
rect 6553 3278 6559 3296
rect 6577 3286 6607 3292
rect 6655 3290 6663 3296
rect 6159 3192 6183 3198
rect 6159 3184 6171 3192
rect 6234 3184 6242 3227
rect 6355 3198 6363 3247
rect 6433 3241 6441 3276
rect 6439 3205 6447 3227
rect 6497 3213 6505 3276
rect 6519 3264 6533 3272
rect 6553 3272 6593 3278
rect 6513 3213 6527 3227
rect 6440 3198 6465 3205
rect 6339 3192 6363 3198
rect 6339 3184 6351 3192
rect 6397 3184 6449 3187
rect 6234 3173 6260 3184
rect 5958 3138 5970 3144
rect 6008 3138 6020 3144
rect 6057 3138 6069 3144
rect 6189 3138 6201 3144
rect 6409 3178 6437 3184
rect 6457 3184 6465 3198
rect 6497 3199 6513 3213
rect 6587 3200 6593 3272
rect 6601 3272 6607 3286
rect 6625 3282 6663 3290
rect 6601 3266 6645 3272
rect 6657 3268 6719 3276
rect 6647 3227 6674 3234
rect 6694 3216 6700 3221
rect 6666 3208 6700 3216
rect 6654 3200 6661 3208
rect 6497 3184 6505 3199
rect 6587 3194 6661 3200
rect 6587 3192 6593 3194
rect 6654 3188 6661 3194
rect 6547 3170 6558 3178
rect 6551 3164 6558 3170
rect 6608 3176 6629 3183
rect 6713 3184 6719 3268
rect 6608 3164 6615 3176
rect 6673 3164 6680 3170
rect 6667 3158 6680 3164
rect 6238 3138 6250 3144
rect 6288 3138 6300 3144
rect 6369 3138 6381 3144
rect 6417 3138 6429 3144
rect 6519 3138 6531 3144
rect 6577 3138 6589 3144
rect 6625 3138 6637 3144
rect 6687 3138 6699 3144
rect 6742 3138 6802 3602
rect 4 3136 6802 3138
rect 6736 3124 6802 3136
rect 4 3122 6802 3124
rect 17 3116 29 3122
rect 57 3116 69 3122
rect 97 3116 109 3122
rect 137 3116 149 3122
rect 177 3116 189 3122
rect 249 3116 261 3122
rect 321 3116 333 3122
rect 383 3116 395 3122
rect 431 3116 443 3122
rect 489 3116 501 3122
rect 589 3116 601 3122
rect 36 3070 48 3076
rect 77 3070 89 3076
rect 116 3070 128 3076
rect 156 3070 168 3076
rect 36 3062 63 3070
rect 77 3062 102 3070
rect 116 3062 142 3070
rect 156 3069 174 3070
rect 156 3062 175 3069
rect 55 3056 63 3062
rect 94 3056 102 3062
rect 134 3056 142 3062
rect 55 3044 70 3056
rect 94 3044 110 3056
rect 134 3044 150 3056
rect 55 2998 63 3044
rect 94 2998 102 3044
rect 134 2998 142 3044
rect 168 3041 175 3062
rect 168 3027 173 3041
rect 231 3033 239 3076
rect 271 3070 279 3096
rect 257 3064 279 3070
rect 340 3096 353 3102
rect 340 3090 347 3096
rect 405 3084 412 3096
rect 257 3058 260 3064
rect 168 2998 175 3027
rect 37 2990 63 2998
rect 77 2990 102 2998
rect 117 2990 142 2998
rect 157 2990 175 2998
rect 231 3019 233 3033
rect 37 2984 49 2990
rect 77 2984 89 2990
rect 117 2984 129 2990
rect 157 2984 169 2990
rect 231 2984 239 3019
rect 253 3002 260 3058
rect 257 2996 260 3002
rect 257 2990 283 2996
rect 275 2944 283 2990
rect 301 2992 307 3076
rect 391 3077 412 3084
rect 462 3090 469 3096
rect 462 3082 473 3090
rect 359 3066 366 3072
rect 427 3066 433 3068
rect 359 3060 433 3066
rect 515 3061 523 3076
rect 619 3116 631 3122
rect 751 3116 763 3122
rect 849 3116 861 3122
rect 929 3116 941 3122
rect 559 3068 571 3076
rect 649 3068 661 3076
rect 559 3062 583 3068
rect 359 3052 366 3060
rect 320 3044 354 3052
rect 320 3039 326 3044
rect 346 3026 373 3033
rect 301 2984 363 2992
rect 375 2988 419 2994
rect 357 2970 395 2978
rect 413 2974 419 2988
rect 427 2988 433 3060
rect 507 3047 523 3061
rect 493 3033 507 3047
rect 427 2982 467 2988
rect 487 2988 501 2996
rect 515 2984 523 3047
rect 575 3013 583 3062
rect 637 3062 661 3068
rect 677 3063 683 3073
rect 637 3013 645 3062
rect 677 3057 703 3063
rect 357 2964 365 2970
rect 413 2968 443 2974
rect 461 2964 467 2982
rect 347 2950 365 2964
rect 393 2950 415 2962
rect 357 2944 365 2950
rect 407 2944 419 2950
rect 461 2924 473 2958
rect 575 2944 583 2999
rect 637 2944 645 2999
rect 677 2983 683 3033
rect 697 3007 703 3057
rect 715 3062 723 3076
rect 743 3076 771 3082
rect 731 3073 783 3076
rect 960 3116 972 3122
rect 1010 3116 1022 3122
rect 1079 3116 1091 3122
rect 1137 3116 1149 3122
rect 1185 3116 1197 3122
rect 1247 3116 1259 3122
rect 1349 3116 1361 3122
rect 1399 3116 1411 3122
rect 1457 3116 1469 3122
rect 1505 3116 1517 3122
rect 1567 3116 1579 3122
rect 1651 3116 1663 3122
rect 1731 3116 1743 3122
rect 1791 3116 1803 3122
rect 1831 3116 1843 3122
rect 1901 3116 1913 3122
rect 1977 3116 1989 3122
rect 2078 3116 2090 3122
rect 2128 3116 2140 3122
rect 1000 3076 1026 3087
rect 819 3068 831 3076
rect 899 3068 911 3076
rect 715 3055 740 3062
rect 733 3033 741 3055
rect 819 3062 843 3068
rect 739 2984 747 3019
rect 797 2987 803 3053
rect 835 3013 843 3062
rect 867 3057 883 3063
rect 899 3062 923 3068
rect 667 2977 683 2983
rect 17 2898 29 2904
rect 57 2898 69 2904
rect 97 2898 109 2904
rect 137 2898 149 2904
rect 177 2898 189 2904
rect 249 2898 261 2904
rect 321 2898 333 2904
rect 387 2898 399 2904
rect 433 2898 445 2904
rect 491 2898 503 2904
rect 551 2898 563 2904
rect 591 2898 603 2904
rect 617 2898 629 2904
rect 657 2898 669 2904
rect 835 2944 843 2999
rect 877 2967 883 3057
rect 915 3013 923 3062
rect 1018 3033 1026 3076
rect 1227 3096 1240 3102
rect 1111 3090 1118 3096
rect 1107 3082 1118 3090
rect 1168 3084 1175 3096
rect 1233 3090 1240 3096
rect 1057 3061 1065 3076
rect 1168 3077 1189 3084
rect 1147 3066 1153 3068
rect 1214 3066 1221 3072
rect 1057 3047 1073 3061
rect 1147 3060 1221 3066
rect 915 2944 923 2999
rect 1018 2984 1026 3019
rect 1057 2984 1065 3047
rect 1073 3033 1087 3047
rect 1079 2988 1093 2996
rect 957 2978 997 2984
rect 957 2976 969 2978
rect 716 2898 728 2904
rect 766 2898 778 2904
rect 811 2898 823 2904
rect 851 2898 863 2904
rect 1147 2988 1153 3060
rect 1214 3052 1221 3060
rect 1226 3044 1260 3052
rect 1254 3039 1260 3044
rect 1207 3026 1234 3033
rect 1113 2982 1153 2988
rect 1161 2988 1205 2994
rect 1113 2964 1119 2982
rect 1161 2974 1167 2988
rect 1273 2992 1279 3076
rect 1547 3096 1560 3102
rect 1431 3090 1438 3096
rect 1427 3082 1438 3090
rect 1488 3084 1495 3096
rect 1553 3090 1560 3096
rect 1319 3068 1331 3076
rect 1319 3062 1343 3068
rect 1335 3013 1343 3062
rect 1377 3061 1385 3076
rect 1488 3077 1509 3084
rect 1467 3066 1473 3068
rect 1534 3066 1541 3072
rect 1377 3047 1393 3061
rect 1467 3060 1541 3066
rect 1217 2984 1279 2992
rect 1137 2968 1167 2974
rect 1185 2970 1223 2978
rect 1215 2964 1223 2970
rect 1107 2924 1119 2958
rect 1165 2950 1187 2962
rect 1215 2950 1233 2964
rect 1161 2944 1173 2950
rect 1215 2944 1223 2950
rect 1335 2944 1343 2999
rect 1377 2984 1385 3047
rect 1393 3033 1407 3047
rect 1399 2988 1413 2996
rect 1467 2988 1473 3060
rect 1534 3052 1541 3060
rect 1546 3044 1580 3052
rect 1574 3039 1580 3044
rect 1527 3026 1554 3033
rect 1433 2982 1473 2988
rect 1481 2988 1525 2994
rect 1433 2964 1439 2982
rect 1481 2974 1487 2988
rect 1593 2992 1599 3076
rect 1636 3041 1644 3096
rect 1695 3062 1703 3076
rect 1723 3076 1751 3082
rect 1711 3073 1763 3076
rect 1695 3055 1720 3062
rect 1713 3033 1721 3055
rect 1813 3053 1820 3096
rect 1871 3076 1881 3086
rect 1537 2984 1599 2992
rect 1457 2968 1487 2974
rect 1505 2970 1543 2978
rect 1535 2964 1543 2970
rect 1427 2924 1439 2958
rect 1485 2950 1507 2962
rect 1535 2950 1553 2964
rect 1481 2944 1493 2950
rect 1535 2944 1543 2950
rect 1636 2944 1644 3027
rect 1719 2984 1727 3019
rect 1813 2991 1820 3039
rect 1871 3033 1879 3076
rect 1931 3066 1943 3076
rect 1969 3076 1997 3082
rect 1957 3073 2009 3076
rect 2074 3076 2100 3087
rect 2159 3116 2171 3122
rect 2271 3116 2283 3122
rect 2327 3116 2339 3122
rect 2421 3116 2433 3122
rect 2483 3116 2495 3122
rect 2531 3116 2543 3122
rect 2589 3116 2601 3122
rect 2637 3116 2649 3122
rect 2697 3116 2709 3122
rect 2737 3116 2749 3122
rect 2811 3116 2823 3122
rect 2891 3116 2903 3122
rect 2937 3116 2949 3122
rect 3070 3116 3082 3122
rect 3149 3116 3161 3122
rect 3231 3116 3243 3122
rect 3279 3116 3291 3122
rect 3359 3116 3371 3122
rect 3457 3116 3469 3122
rect 3567 3116 3579 3122
rect 3672 3116 3684 3122
rect 3728 3116 3740 3122
rect 1905 3058 1943 3066
rect 2017 3062 2025 3076
rect 1871 3019 1873 3033
rect 1803 2984 1820 2991
rect 1871 2984 1879 3019
rect 891 2898 903 2904
rect 931 2898 943 2904
rect 977 2898 989 2904
rect 1077 2898 1089 2904
rect 1135 2898 1147 2904
rect 1181 2898 1193 2904
rect 1247 2898 1259 2904
rect 1311 2898 1323 2904
rect 1351 2898 1363 2904
rect 1397 2898 1409 2904
rect 1455 2898 1467 2904
rect 1501 2898 1513 2904
rect 1567 2898 1579 2904
rect 1651 2898 1663 2904
rect 1914 2944 1922 3058
rect 2000 3055 2025 3062
rect 1999 3033 2007 3055
rect 2074 3033 2082 3076
rect 2189 3068 2201 3076
rect 2177 3062 2201 3068
rect 1993 2984 2001 3019
rect 2074 2984 2082 3019
rect 2177 3013 2185 3062
rect 2256 3041 2264 3096
rect 2359 3076 2369 3086
rect 2297 3066 2309 3076
rect 2297 3058 2335 3066
rect 1696 2898 1708 2904
rect 1746 2898 1758 2904
rect 1831 2898 1843 2904
rect 1887 2898 1899 2904
rect 1931 2898 1943 2904
rect 2103 2978 2143 2984
rect 2131 2976 2143 2978
rect 2177 2944 2185 2999
rect 2207 2977 2233 2983
rect 2256 2944 2264 3027
rect 2318 2944 2326 3058
rect 2361 3033 2369 3076
rect 2367 3019 2369 3033
rect 2361 2984 2369 3019
rect 2440 3096 2453 3102
rect 2440 3090 2447 3096
rect 2505 3084 2512 3096
rect 2401 2992 2407 3076
rect 2491 3077 2512 3084
rect 2562 3090 2569 3096
rect 2562 3082 2573 3090
rect 2459 3066 2466 3072
rect 2527 3066 2533 3068
rect 2459 3060 2533 3066
rect 2615 3061 2623 3076
rect 2459 3052 2466 3060
rect 2420 3044 2454 3052
rect 2420 3039 2426 3044
rect 2446 3026 2473 3033
rect 2401 2984 2463 2992
rect 2475 2988 2519 2994
rect 1962 2898 1974 2904
rect 2012 2898 2024 2904
rect 2111 2898 2123 2904
rect 2157 2898 2169 2904
rect 2197 2898 2209 2904
rect 2271 2898 2283 2904
rect 2457 2970 2495 2978
rect 2513 2974 2519 2988
rect 2527 2988 2533 3060
rect 2607 3047 2623 3061
rect 2593 3033 2607 3047
rect 2527 2982 2567 2988
rect 2587 2988 2601 2996
rect 2615 2984 2623 3047
rect 2656 3041 2664 3096
rect 2720 3053 2727 3096
rect 2796 3041 2804 3096
rect 2855 3062 2863 3076
rect 2883 3076 2911 3082
rect 2871 3073 2923 3076
rect 2855 3055 2880 3062
rect 2457 2964 2465 2970
rect 2513 2968 2543 2974
rect 2561 2964 2567 2982
rect 2447 2950 2465 2964
rect 2493 2950 2515 2962
rect 2457 2944 2465 2950
rect 2507 2944 2519 2950
rect 2561 2924 2573 2958
rect 2656 2944 2664 3027
rect 2720 2991 2727 3039
rect 2873 3033 2881 3055
rect 2720 2984 2737 2991
rect 2796 2944 2804 3027
rect 2956 3033 2964 3076
rect 3016 3058 3034 3060
rect 3016 3049 3046 3058
rect 3119 3068 3131 3076
rect 3119 3062 3143 3068
rect 3016 3021 3024 3049
rect 2879 2984 2887 3019
rect 2956 2984 2964 3019
rect 2297 2898 2309 2904
rect 2341 2898 2353 2904
rect 2421 2898 2433 2904
rect 2487 2898 2499 2904
rect 2533 2898 2545 2904
rect 2591 2898 2603 2904
rect 2637 2898 2649 2904
rect 2697 2898 2709 2904
rect 2811 2898 2823 2904
rect 2856 2898 2868 2904
rect 2906 2898 2918 2904
rect 3015 2952 3022 3007
rect 3135 3013 3143 3062
rect 3195 3062 3203 3076
rect 3223 3076 3251 3082
rect 3211 3073 3263 3076
rect 3309 3068 3321 3076
rect 3389 3068 3401 3076
rect 3449 3076 3477 3082
rect 3437 3073 3489 3076
rect 3599 3076 3609 3086
rect 3771 3116 3783 3122
rect 3811 3116 3823 3122
rect 3861 3116 3873 3122
rect 3923 3116 3935 3122
rect 3971 3116 3983 3122
rect 4029 3116 4041 3122
rect 4097 3116 4109 3122
rect 4250 3116 4262 3122
rect 4301 3116 4313 3122
rect 4363 3116 4375 3122
rect 4411 3116 4423 3122
rect 4469 3116 4481 3122
rect 4591 3116 4603 3122
rect 4671 3116 4683 3122
rect 3880 3096 3893 3102
rect 3880 3090 3887 3096
rect 3945 3084 3952 3096
rect 3297 3062 3321 3068
rect 3195 3055 3220 3062
rect 3177 3037 3193 3043
rect 3015 2946 3062 2952
rect 3015 2944 3023 2946
rect 3051 2944 3062 2946
rect 3135 2944 3143 2999
rect 3177 2963 3183 3037
rect 3213 3033 3221 3055
rect 3219 2984 3227 3019
rect 3297 3013 3305 3062
rect 3377 3062 3401 3068
rect 3177 2957 3193 2963
rect 2937 2898 2949 2904
rect 3031 2898 3043 2904
rect 3071 2898 3083 2904
rect 3111 2898 3123 2904
rect 3151 2898 3163 2904
rect 3297 2944 3305 2999
rect 3337 2983 3343 3053
rect 3377 3013 3385 3062
rect 3417 3007 3423 3073
rect 3497 3062 3505 3076
rect 3480 3055 3505 3062
rect 3479 3033 3487 3055
rect 3537 3066 3549 3076
rect 3537 3058 3575 3066
rect 3337 2977 3353 2983
rect 3327 2957 3353 2963
rect 3377 2944 3385 2999
rect 3473 2984 3481 3019
rect 3196 2898 3208 2904
rect 3246 2898 3258 2904
rect 3277 2898 3289 2904
rect 3317 2898 3329 2904
rect 3357 2898 3369 2904
rect 3397 2898 3409 2904
rect 3517 2983 3523 3053
rect 3517 2977 3533 2983
rect 3558 2944 3566 3058
rect 3601 3033 3609 3076
rect 3607 3019 3609 3033
rect 3700 3033 3707 3076
rect 3747 3057 3763 3063
rect 3601 2984 3609 3019
rect 3693 2996 3699 3019
rect 3757 3007 3763 3057
rect 3792 3041 3801 3076
rect 3787 3027 3801 3041
rect 3672 2990 3699 2996
rect 3672 2984 3684 2990
rect 3792 2984 3801 3027
rect 3841 2992 3847 3076
rect 3931 3077 3952 3084
rect 4002 3090 4009 3096
rect 4002 3082 4013 3090
rect 3899 3066 3906 3072
rect 3967 3066 3973 3068
rect 3899 3060 3973 3066
rect 4055 3061 4063 3076
rect 4089 3076 4117 3082
rect 4077 3073 4129 3076
rect 4137 3062 4145 3076
rect 3899 3052 3906 3060
rect 3860 3044 3894 3052
rect 3860 3039 3866 3044
rect 3886 3026 3913 3033
rect 3841 2984 3903 2992
rect 3915 2988 3959 2994
rect 3442 2898 3454 2904
rect 3492 2898 3504 2904
rect 3663 2904 3691 2910
rect 3703 2976 3731 2982
rect 3537 2898 3549 2904
rect 3581 2898 3593 2904
rect 3711 2898 3723 2904
rect 3771 2898 3783 2904
rect 3811 2898 3823 2906
rect 3897 2970 3935 2978
rect 3953 2974 3959 2988
rect 3967 2988 3973 3060
rect 4047 3047 4063 3061
rect 4120 3055 4145 3062
rect 4196 3058 4214 3060
rect 4033 3033 4047 3047
rect 3967 2982 4007 2988
rect 4027 2988 4041 2996
rect 4055 2984 4063 3047
rect 4119 3033 4127 3055
rect 4196 3049 4226 3058
rect 4320 3096 4333 3102
rect 4320 3090 4327 3096
rect 4385 3084 4392 3096
rect 4196 3021 4204 3049
rect 4113 2984 4121 3019
rect 3897 2964 3905 2970
rect 3953 2968 3983 2974
rect 4001 2964 4007 2982
rect 3887 2950 3905 2964
rect 3933 2950 3955 2962
rect 3897 2944 3905 2950
rect 3947 2944 3959 2950
rect 4001 2924 4013 2958
rect 4195 2952 4202 3007
rect 4281 2992 4287 3076
rect 4371 3077 4392 3084
rect 4442 3090 4449 3096
rect 4442 3082 4453 3090
rect 4339 3066 4346 3072
rect 4543 3110 4571 3116
rect 4583 3076 4611 3080
rect 4711 3108 4723 3122
rect 4771 3108 4783 3122
rect 4820 3116 4832 3122
rect 4876 3116 4888 3122
rect 4971 3116 4983 3122
rect 4407 3066 4413 3068
rect 4339 3060 4413 3066
rect 4495 3061 4503 3076
rect 4339 3052 4346 3060
rect 4300 3044 4334 3052
rect 4300 3039 4306 3044
rect 4326 3026 4353 3033
rect 4281 2984 4343 2992
rect 4355 2988 4399 2994
rect 4195 2946 4242 2952
rect 4195 2944 4203 2946
rect 4231 2944 4242 2946
rect 4337 2970 4375 2978
rect 4393 2974 4399 2988
rect 4407 2988 4413 3060
rect 4487 3047 4503 3061
rect 4555 3066 4561 3076
rect 4571 3074 4623 3076
rect 4555 3059 4584 3066
rect 4473 3033 4487 3047
rect 4407 2982 4447 2988
rect 4467 2988 4481 2996
rect 4495 2984 4503 3047
rect 4576 3033 4584 3059
rect 4656 3041 4664 3096
rect 4739 3076 4741 3078
rect 4739 3072 4753 3076
rect 4739 3041 4745 3072
rect 4791 3066 4798 3088
rect 5000 3116 5012 3122
rect 5056 3116 5068 3122
rect 4756 3060 4798 3066
rect 4575 2984 4583 3019
rect 4337 2964 4345 2970
rect 4393 2968 4423 2974
rect 4441 2964 4447 2982
rect 4327 2950 4345 2964
rect 4373 2950 4395 2962
rect 4337 2944 4345 2950
rect 4387 2944 4399 2950
rect 4441 2924 4453 2958
rect 4656 2944 4664 3027
rect 3861 2898 3873 2904
rect 3927 2898 3939 2904
rect 3973 2898 3985 2904
rect 4031 2898 4043 2904
rect 4082 2898 4094 2904
rect 4132 2898 4144 2904
rect 4211 2898 4223 2904
rect 4251 2898 4263 2904
rect 4301 2898 4313 2904
rect 4367 2898 4379 2904
rect 4413 2898 4425 2904
rect 4471 2898 4483 2904
rect 4541 2898 4553 2904
rect 4611 2898 4623 2904
rect 4671 2898 4683 2904
rect 4739 2980 4745 3027
rect 4756 3022 4765 3060
rect 4756 2992 4765 3010
rect 4853 3033 4860 3076
rect 4956 3041 4964 3096
rect 5117 3116 5129 3122
rect 5177 3116 5189 3122
rect 5217 3116 5229 3122
rect 5281 3116 5293 3122
rect 5343 3116 5355 3122
rect 5391 3116 5403 3122
rect 5449 3116 5461 3122
rect 5511 3116 5523 3122
rect 5551 3116 5563 3122
rect 5597 3116 5609 3122
rect 5750 3116 5762 3122
rect 5851 3116 5863 3122
rect 5897 3116 5909 3122
rect 4861 2996 4867 3019
rect 4756 2986 4797 2992
rect 4861 2990 4888 2996
rect 4739 2976 4753 2980
rect 4739 2974 4741 2976
rect 4791 2952 4797 2986
rect 4876 2984 4888 2990
rect 4711 2898 4723 2904
rect 4771 2898 4783 2912
rect 4829 2976 4857 2982
rect 4869 2904 4897 2910
rect 4956 2944 4964 3027
rect 5033 3033 5040 3076
rect 5136 3041 5144 3096
rect 5200 3053 5207 3096
rect 5041 2996 5047 3019
rect 5041 2990 5068 2996
rect 5056 2984 5068 2990
rect 5009 2976 5037 2982
rect 5049 2904 5077 2910
rect 5136 2944 5144 3027
rect 5200 2991 5207 3039
rect 5300 3096 5313 3102
rect 5300 3090 5307 3096
rect 5365 3084 5372 3096
rect 5261 2992 5267 3076
rect 5351 3077 5372 3084
rect 5422 3090 5429 3096
rect 5422 3082 5433 3090
rect 5319 3066 5326 3072
rect 5387 3066 5393 3068
rect 5319 3060 5393 3066
rect 5475 3061 5483 3076
rect 5319 3052 5326 3060
rect 5280 3044 5314 3052
rect 5280 3039 5286 3044
rect 5306 3026 5333 3033
rect 5200 2984 5217 2991
rect 5261 2984 5323 2992
rect 5335 2988 5379 2994
rect 5317 2970 5355 2978
rect 5373 2974 5379 2988
rect 5387 2988 5393 3060
rect 5467 3047 5483 3061
rect 5453 3033 5467 3047
rect 5387 2982 5427 2988
rect 5447 2988 5461 2996
rect 5475 2984 5483 3047
rect 5533 3053 5540 3096
rect 5589 3076 5617 3082
rect 5577 3073 5629 3076
rect 5637 3062 5645 3076
rect 5620 3055 5645 3062
rect 5696 3058 5714 3060
rect 5533 2991 5540 3039
rect 5619 3033 5627 3055
rect 5696 3049 5726 3058
rect 5803 3110 5831 3116
rect 5843 3076 5871 3080
rect 5977 3108 5989 3122
rect 6037 3108 6049 3122
rect 5815 3066 5821 3076
rect 5831 3074 5883 3076
rect 5815 3059 5844 3066
rect 5317 2964 5325 2970
rect 5373 2968 5403 2974
rect 5421 2964 5427 2982
rect 5307 2950 5325 2964
rect 5353 2950 5375 2962
rect 5317 2944 5325 2950
rect 5367 2944 5379 2950
rect 5421 2924 5433 2958
rect 5523 2984 5540 2991
rect 5613 2984 5621 3019
rect 5696 3021 5704 3049
rect 4837 2898 4849 2904
rect 4971 2898 4983 2904
rect 5017 2898 5029 2904
rect 5117 2898 5129 2904
rect 5177 2898 5189 2904
rect 5281 2898 5293 2904
rect 5347 2898 5359 2904
rect 5393 2898 5405 2904
rect 5451 2898 5463 2904
rect 5551 2898 5563 2904
rect 5657 2963 5663 3013
rect 5836 3033 5844 3059
rect 5916 3041 5924 3096
rect 5962 3066 5969 3088
rect 6019 3076 6021 3078
rect 6007 3072 6021 3076
rect 5962 3060 6004 3066
rect 5647 2957 5663 2963
rect 5695 2952 5702 3007
rect 5835 2984 5843 3019
rect 5695 2946 5742 2952
rect 5695 2944 5703 2946
rect 5731 2944 5742 2946
rect 5582 2898 5594 2904
rect 5632 2898 5644 2904
rect 5711 2898 5723 2904
rect 5751 2898 5763 2904
rect 5916 2944 5924 3027
rect 5995 3022 6004 3060
rect 6015 3041 6021 3072
rect 6098 3116 6110 3122
rect 6148 3116 6160 3122
rect 6094 3076 6120 3087
rect 6191 3116 6203 3122
rect 6231 3116 6243 3122
rect 6257 3116 6269 3122
rect 6352 3116 6364 3122
rect 6408 3116 6420 3122
rect 6471 3116 6483 3122
rect 6094 3033 6102 3076
rect 6213 3053 6220 3096
rect 5995 2992 6004 3010
rect 5963 2986 6004 2992
rect 5963 2952 5969 2986
rect 6015 2980 6021 3027
rect 6276 3041 6284 3096
rect 6497 3116 6509 3122
rect 6577 3116 6589 3122
rect 6094 2984 6102 3019
rect 6213 2991 6220 3039
rect 6203 2984 6220 2991
rect 6007 2976 6021 2980
rect 5801 2898 5813 2904
rect 5871 2898 5883 2904
rect 6019 2974 6021 2976
rect 5897 2898 5909 2904
rect 5977 2898 5989 2912
rect 6123 2978 6163 2984
rect 6151 2976 6163 2978
rect 6276 2944 6284 3027
rect 6380 3033 6387 3076
rect 6456 3041 6464 3096
rect 6516 3041 6524 3096
rect 6569 3076 6597 3082
rect 6557 3073 6609 3076
rect 6617 3062 6625 3076
rect 6600 3055 6625 3062
rect 6373 2996 6379 3019
rect 6352 2990 6379 2996
rect 6352 2984 6364 2990
rect 6037 2898 6049 2904
rect 6131 2898 6143 2904
rect 6231 2898 6243 2904
rect 6343 2904 6371 2910
rect 6383 2976 6411 2982
rect 6456 2944 6464 3027
rect 6516 2944 6524 3027
rect 6599 3033 6607 3055
rect 6593 2984 6601 3019
rect 6257 2898 6269 2904
rect 6391 2898 6403 2904
rect 6471 2898 6483 2904
rect 6497 2898 6509 2904
rect 6562 2898 6574 2904
rect 6612 2898 6624 2904
rect -62 2896 6736 2898
rect -62 2884 4 2896
rect -62 2882 2053 2884
rect -62 2418 -2 2882
rect 17 2876 29 2882
rect 131 2876 143 2882
rect 181 2876 193 2882
rect 247 2876 259 2882
rect 293 2876 305 2882
rect 351 2876 363 2882
rect 397 2876 409 2882
rect 511 2876 523 2882
rect 561 2876 573 2882
rect 627 2876 639 2882
rect 673 2876 685 2882
rect 731 2876 743 2882
rect 809 2876 821 2882
rect 36 2753 44 2836
rect 217 2830 225 2836
rect 267 2830 279 2836
rect 207 2816 225 2830
rect 253 2818 275 2830
rect 321 2822 333 2856
rect 217 2810 225 2816
rect 217 2802 255 2810
rect 273 2806 303 2812
rect 103 2789 120 2796
rect 113 2741 120 2789
rect 161 2788 223 2796
rect 36 2684 44 2739
rect 113 2684 120 2727
rect 161 2704 167 2788
rect 273 2792 279 2806
rect 321 2798 327 2816
rect 235 2786 279 2792
rect 287 2792 327 2798
rect 206 2747 233 2754
rect 180 2736 186 2741
rect 180 2728 214 2736
rect 219 2720 226 2728
rect 287 2720 293 2792
rect 347 2784 361 2792
rect 353 2733 367 2747
rect 375 2733 383 2796
rect 416 2753 424 2836
rect 597 2830 605 2836
rect 647 2830 659 2836
rect 587 2816 605 2830
rect 633 2818 655 2830
rect 701 2822 713 2856
rect 597 2810 605 2816
rect 597 2802 635 2810
rect 653 2806 683 2812
rect 483 2789 500 2796
rect 219 2714 293 2720
rect 367 2719 383 2733
rect 493 2741 500 2789
rect 541 2788 603 2796
rect 219 2708 226 2714
rect 287 2712 293 2714
rect 251 2696 272 2703
rect 375 2704 383 2719
rect 200 2684 207 2690
rect 265 2684 272 2696
rect 322 2690 333 2698
rect 322 2684 329 2690
rect 200 2678 213 2684
rect 416 2684 424 2739
rect 447 2717 473 2723
rect 493 2684 500 2727
rect 541 2704 547 2788
rect 653 2792 659 2806
rect 701 2798 707 2816
rect 615 2786 659 2792
rect 667 2792 707 2798
rect 586 2747 613 2754
rect 560 2736 566 2741
rect 560 2728 594 2736
rect 599 2720 606 2728
rect 667 2720 673 2792
rect 727 2784 741 2792
rect 733 2733 747 2747
rect 755 2733 763 2796
rect 599 2714 673 2720
rect 747 2719 763 2733
rect 599 2708 606 2714
rect 667 2712 673 2714
rect 631 2696 652 2703
rect 755 2704 763 2719
rect 791 2761 799 2796
rect 835 2790 843 2836
rect 857 2874 869 2882
rect 897 2876 909 2882
rect 937 2876 949 2882
rect 977 2876 989 2882
rect 1017 2876 1029 2882
rect 1057 2876 1069 2882
rect 1097 2876 1109 2882
rect 1177 2876 1189 2882
rect 1331 2876 1343 2882
rect 1411 2876 1423 2882
rect 817 2784 843 2790
rect 817 2778 820 2784
rect 791 2747 793 2761
rect 791 2704 799 2747
rect 813 2722 820 2778
rect 879 2753 888 2796
rect 957 2781 965 2836
rect 1037 2781 1045 2836
rect 879 2739 893 2753
rect 817 2716 820 2722
rect 817 2710 839 2716
rect 580 2684 587 2690
rect 645 2684 652 2696
rect 702 2690 713 2698
rect 702 2684 709 2690
rect 580 2678 593 2684
rect 831 2684 839 2710
rect 879 2704 888 2739
rect 957 2718 965 2767
rect 1037 2718 1045 2767
rect 1116 2753 1124 2836
rect 1169 2798 1197 2804
rect 1209 2870 1237 2876
rect 1456 2876 1468 2882
rect 1506 2876 1518 2882
rect 1351 2802 1363 2804
rect 1323 2796 1363 2802
rect 1216 2790 1228 2796
rect 1201 2784 1228 2790
rect 1201 2761 1207 2784
rect 1294 2761 1302 2796
rect 957 2712 981 2718
rect 1037 2712 1061 2718
rect 969 2704 981 2712
rect 1049 2704 1061 2712
rect 17 2658 29 2664
rect 91 2658 103 2664
rect 131 2658 143 2664
rect 181 2658 193 2664
rect 243 2658 255 2664
rect 291 2658 303 2664
rect 349 2658 361 2664
rect 397 2658 409 2664
rect 471 2658 483 2664
rect 511 2658 523 2664
rect 561 2658 573 2664
rect 623 2658 635 2664
rect 671 2658 683 2664
rect 729 2658 741 2664
rect 809 2658 821 2664
rect 857 2658 869 2664
rect 897 2658 909 2664
rect 1116 2684 1124 2739
rect 1193 2704 1200 2747
rect 1396 2753 1404 2836
rect 1537 2876 1549 2882
rect 1617 2876 1629 2882
rect 1657 2876 1669 2882
rect 1697 2876 1709 2882
rect 1796 2876 1808 2882
rect 1846 2876 1858 2882
rect 1907 2876 1919 2882
rect 1982 2876 1994 2882
rect 2032 2876 2044 2882
rect 1479 2761 1487 2796
rect 1560 2789 1577 2796
rect 1294 2704 1302 2747
rect 1294 2693 1320 2704
rect 939 2658 951 2664
rect 1019 2658 1031 2664
rect 1097 2658 1109 2664
rect 1160 2658 1172 2664
rect 1216 2658 1228 2664
rect 1396 2684 1404 2739
rect 1473 2725 1481 2747
rect 1560 2741 1567 2789
rect 1455 2718 1480 2725
rect 1455 2704 1463 2718
rect 1471 2704 1523 2707
rect 1483 2698 1511 2704
rect 1560 2684 1567 2727
rect 1597 2723 1603 2793
rect 1637 2781 1645 2836
rect 1939 2797 1943 2806
rect 1720 2789 1737 2796
rect 1597 2717 1613 2723
rect 1637 2718 1645 2767
rect 1720 2741 1727 2789
rect 1819 2761 1827 2796
rect 1877 2788 1885 2796
rect 1877 2780 1913 2788
rect 1637 2712 1661 2718
rect 1649 2704 1661 2712
rect 1298 2658 1310 2664
rect 1348 2658 1360 2664
rect 1411 2658 1423 2664
rect 1491 2658 1503 2664
rect 1537 2658 1549 2664
rect 1577 2658 1589 2664
rect 1720 2684 1727 2727
rect 1813 2725 1821 2747
rect 1795 2718 1820 2725
rect 1918 2724 1924 2779
rect 1934 2753 1943 2797
rect 2067 2882 3793 2884
rect 2131 2876 2143 2882
rect 2201 2876 2213 2882
rect 2267 2876 2279 2882
rect 2313 2876 2325 2882
rect 2371 2876 2383 2882
rect 2417 2876 2429 2882
rect 2457 2876 2469 2882
rect 2151 2802 2163 2804
rect 2123 2796 2163 2802
rect 2237 2830 2245 2836
rect 2287 2830 2299 2836
rect 2227 2816 2245 2830
rect 2273 2818 2295 2830
rect 2341 2822 2353 2856
rect 2237 2810 2245 2816
rect 2237 2802 2275 2810
rect 2293 2806 2323 2812
rect 2013 2761 2021 2796
rect 2094 2761 2102 2796
rect 2181 2788 2243 2796
rect 1795 2704 1803 2718
rect 1903 2712 1913 2718
rect 1811 2704 1863 2707
rect 1823 2698 1851 2704
rect 1903 2684 1909 2712
rect 1940 2704 1947 2739
rect 2019 2725 2027 2747
rect 2020 2718 2045 2725
rect 1977 2704 2029 2707
rect 1989 2698 2017 2704
rect 2037 2704 2045 2718
rect 2094 2704 2102 2747
rect 2181 2704 2187 2788
rect 2293 2792 2299 2806
rect 2341 2798 2347 2816
rect 2255 2786 2299 2792
rect 2307 2792 2347 2798
rect 2226 2747 2253 2754
rect 2200 2736 2206 2741
rect 2200 2728 2234 2736
rect 2239 2720 2246 2728
rect 2307 2720 2313 2792
rect 2497 2876 2509 2882
rect 2591 2876 2603 2882
rect 2641 2876 2653 2882
rect 2707 2876 2719 2882
rect 2753 2876 2765 2882
rect 2811 2876 2823 2882
rect 2862 2876 2874 2882
rect 2912 2876 2924 2882
rect 3011 2876 3023 2882
rect 3077 2876 3089 2882
rect 3135 2876 3147 2882
rect 3181 2876 3193 2882
rect 3247 2876 3259 2882
rect 3297 2876 3309 2882
rect 3357 2876 3369 2882
rect 3427 2876 3439 2882
rect 2367 2784 2381 2792
rect 2373 2733 2387 2747
rect 2395 2733 2403 2796
rect 2437 2781 2445 2836
rect 2239 2714 2313 2720
rect 2387 2719 2403 2733
rect 2239 2708 2246 2714
rect 2307 2712 2313 2714
rect 2094 2693 2120 2704
rect 2271 2696 2292 2703
rect 2395 2704 2403 2719
rect 2437 2718 2445 2767
rect 2516 2753 2524 2836
rect 2576 2753 2584 2836
rect 2677 2830 2685 2836
rect 2727 2830 2739 2836
rect 2667 2816 2685 2830
rect 2713 2818 2735 2830
rect 2781 2822 2793 2856
rect 2677 2810 2685 2816
rect 2677 2802 2715 2810
rect 2733 2806 2763 2812
rect 2621 2788 2683 2796
rect 2437 2712 2461 2718
rect 2449 2704 2461 2712
rect 2220 2684 2227 2690
rect 2285 2684 2292 2696
rect 2342 2690 2353 2698
rect 2342 2684 2349 2690
rect 2220 2678 2233 2684
rect 2516 2684 2524 2739
rect 2576 2684 2584 2739
rect 2621 2704 2627 2788
rect 2733 2792 2739 2806
rect 2781 2798 2787 2816
rect 2695 2786 2739 2792
rect 2747 2792 2787 2798
rect 2666 2747 2693 2754
rect 2640 2736 2646 2741
rect 2640 2728 2674 2736
rect 2679 2720 2686 2728
rect 2747 2720 2753 2792
rect 3031 2802 3043 2804
rect 3003 2796 3043 2802
rect 3107 2822 3119 2856
rect 3161 2830 3173 2836
rect 3215 2830 3223 2836
rect 3165 2818 3187 2830
rect 3215 2816 3233 2830
rect 3113 2798 3119 2816
rect 3137 2806 3167 2812
rect 3215 2810 3223 2816
rect 2807 2784 2821 2792
rect 2813 2733 2827 2747
rect 2835 2733 2843 2796
rect 2893 2761 2901 2796
rect 2974 2761 2982 2796
rect 2679 2714 2753 2720
rect 2827 2719 2843 2733
rect 2899 2725 2907 2747
rect 2679 2708 2686 2714
rect 2747 2712 2753 2714
rect 2711 2696 2732 2703
rect 2835 2704 2843 2719
rect 2900 2718 2925 2725
rect 2660 2684 2667 2690
rect 2725 2684 2732 2696
rect 2782 2690 2793 2698
rect 2782 2684 2789 2690
rect 2660 2678 2673 2684
rect 2857 2704 2909 2707
rect 2869 2698 2897 2704
rect 2917 2704 2925 2718
rect 2974 2704 2982 2747
rect 3057 2733 3065 2796
rect 3079 2784 3093 2792
rect 3113 2792 3153 2798
rect 3073 2733 3087 2747
rect 3057 2719 3073 2733
rect 3147 2720 3153 2792
rect 3161 2792 3167 2806
rect 3185 2802 3223 2810
rect 3161 2786 3205 2792
rect 3217 2788 3279 2796
rect 3207 2747 3234 2754
rect 3254 2736 3260 2741
rect 3226 2728 3260 2736
rect 3214 2720 3221 2728
rect 3057 2704 3065 2719
rect 3147 2714 3221 2720
rect 3147 2712 3153 2714
rect 2974 2693 3000 2704
rect 3214 2708 3221 2714
rect 3107 2690 3118 2698
rect 3111 2684 3118 2690
rect 3168 2696 3189 2703
rect 3273 2704 3279 2788
rect 3316 2753 3324 2836
rect 3482 2876 3494 2882
rect 3532 2876 3544 2882
rect 3601 2876 3613 2882
rect 3671 2876 3683 2882
rect 3702 2876 3714 2882
rect 3752 2876 3764 2882
rect 3807 2882 6736 2884
rect 3821 2876 3833 2882
rect 3891 2876 3903 2882
rect 3951 2876 3963 2882
rect 3397 2761 3405 2796
rect 3513 2761 3521 2796
rect 3635 2761 3643 2796
rect 3733 2761 3741 2796
rect 3977 2876 3989 2882
rect 4057 2876 4069 2882
rect 4191 2876 4203 2882
rect 4242 2876 4254 2882
rect 4292 2876 4304 2882
rect 4371 2876 4383 2882
rect 4411 2876 4423 2882
rect 4461 2876 4473 2882
rect 4527 2876 4539 2882
rect 4573 2876 4585 2882
rect 4631 2876 4643 2882
rect 4677 2876 4689 2882
rect 4737 2876 4749 2882
rect 4822 2876 4834 2882
rect 4872 2876 4884 2882
rect 4971 2876 4983 2882
rect 3168 2684 3175 2696
rect 3233 2684 3240 2690
rect 3227 2678 3240 2684
rect 3316 2684 3324 2739
rect 3396 2721 3404 2747
rect 3519 2725 3527 2747
rect 3396 2714 3425 2721
rect 3520 2718 3545 2725
rect 3636 2721 3644 2747
rect 3739 2725 3747 2747
rect 3357 2704 3409 2706
rect 3419 2704 3425 2714
rect 3477 2704 3529 2707
rect 3369 2700 3397 2704
rect 3409 2664 3437 2670
rect 3489 2698 3517 2704
rect 3537 2704 3545 2718
rect 3615 2714 3644 2721
rect 3740 2718 3765 2725
rect 3615 2704 3621 2714
rect 3631 2704 3683 2706
rect 3603 2664 3631 2670
rect 3643 2700 3671 2704
rect 3697 2704 3749 2707
rect 3709 2698 3737 2704
rect 3757 2704 3765 2718
rect 3797 2723 3803 2793
rect 3855 2761 3863 2796
rect 3797 2717 3813 2723
rect 3856 2721 3864 2747
rect 3835 2714 3864 2721
rect 3835 2704 3841 2714
rect 3917 2723 3923 2773
rect 3936 2753 3944 2836
rect 4000 2789 4017 2796
rect 4000 2741 4007 2789
rect 3907 2717 3923 2723
rect 3851 2704 3903 2706
rect 3823 2664 3851 2670
rect 3863 2700 3891 2704
rect 3936 2684 3944 2739
rect 4000 2684 4007 2727
rect 4037 2723 4043 2853
rect 4211 2802 4223 2804
rect 4183 2796 4223 2802
rect 4355 2834 4363 2836
rect 4391 2834 4402 2836
rect 4355 2828 4402 2834
rect 4307 2817 4343 2823
rect 4080 2789 4097 2796
rect 4080 2741 4087 2789
rect 4154 2761 4162 2796
rect 4273 2761 4281 2796
rect 4027 2717 4043 2723
rect 4080 2684 4087 2727
rect 4154 2704 4162 2747
rect 4337 2747 4343 2817
rect 4355 2773 4362 2828
rect 4497 2830 4505 2836
rect 4547 2830 4559 2836
rect 4487 2816 4505 2830
rect 4533 2818 4555 2830
rect 4601 2822 4613 2856
rect 4497 2810 4505 2816
rect 4497 2802 4535 2810
rect 4553 2806 4583 2812
rect 4441 2788 4503 2796
rect 4279 2725 4287 2747
rect 4356 2731 4364 2759
rect 4280 2718 4305 2725
rect 4356 2722 4386 2731
rect 4356 2720 4374 2722
rect 4237 2704 4289 2707
rect 4154 2693 4180 2704
rect 1619 2658 1631 2664
rect 1697 2658 1709 2664
rect 1737 2658 1749 2664
rect 1831 2658 1843 2664
rect 1877 2658 1885 2664
rect 1917 2658 1929 2664
rect 1997 2658 2009 2664
rect 2098 2658 2110 2664
rect 2148 2658 2160 2664
rect 2201 2658 2213 2664
rect 2263 2658 2275 2664
rect 2311 2658 2323 2664
rect 2369 2658 2381 2664
rect 2419 2658 2431 2664
rect 2497 2658 2509 2664
rect 2591 2658 2603 2664
rect 2641 2658 2653 2664
rect 2703 2658 2715 2664
rect 2751 2658 2763 2664
rect 2809 2658 2821 2664
rect 2877 2658 2889 2664
rect 2978 2658 2990 2664
rect 3028 2658 3040 2664
rect 3079 2658 3091 2664
rect 3137 2658 3149 2664
rect 3185 2658 3197 2664
rect 3247 2658 3259 2664
rect 3297 2658 3309 2664
rect 3377 2658 3389 2664
rect 3497 2658 3509 2664
rect 3651 2658 3663 2664
rect 3717 2658 3729 2664
rect 3871 2658 3883 2664
rect 3951 2658 3963 2664
rect 3977 2658 3989 2664
rect 4017 2658 4029 2664
rect 4057 2658 4069 2664
rect 4097 2658 4109 2664
rect 4249 2698 4277 2704
rect 4297 2704 4305 2718
rect 4441 2704 4447 2788
rect 4553 2792 4559 2806
rect 4601 2798 4607 2816
rect 4515 2786 4559 2792
rect 4567 2792 4607 2798
rect 4486 2747 4513 2754
rect 4460 2736 4466 2741
rect 4460 2728 4494 2736
rect 4499 2720 4506 2728
rect 4567 2720 4573 2792
rect 4627 2784 4641 2792
rect 4633 2733 4647 2747
rect 4655 2733 4663 2796
rect 4696 2753 4704 2836
rect 5021 2876 5033 2882
rect 5091 2876 5103 2882
rect 5137 2876 5149 2882
rect 5239 2876 5251 2882
rect 5302 2876 5314 2882
rect 5352 2876 5364 2882
rect 5117 2802 5129 2804
rect 5117 2796 5157 2802
rect 4760 2789 4777 2796
rect 4499 2714 4573 2720
rect 4647 2719 4663 2733
rect 4760 2741 4767 2789
rect 4853 2761 4861 2796
rect 4943 2789 4960 2796
rect 4499 2708 4506 2714
rect 4567 2712 4573 2714
rect 4531 2696 4552 2703
rect 4655 2704 4663 2719
rect 4480 2684 4487 2690
rect 4545 2684 4552 2696
rect 4602 2690 4613 2698
rect 4602 2684 4609 2690
rect 4480 2678 4493 2684
rect 4696 2684 4704 2739
rect 4760 2684 4767 2727
rect 4787 2717 4813 2723
rect 4859 2725 4867 2747
rect 4953 2741 4960 2789
rect 5055 2761 5063 2796
rect 5178 2761 5186 2796
rect 5217 2790 5225 2836
rect 5421 2876 5433 2882
rect 5491 2876 5503 2882
rect 5551 2876 5563 2882
rect 5601 2876 5613 2882
rect 5667 2876 5679 2882
rect 5713 2876 5725 2882
rect 5771 2876 5783 2882
rect 5217 2784 5243 2790
rect 5240 2778 5243 2784
rect 5197 2767 5203 2773
rect 4860 2718 4885 2725
rect 4817 2704 4869 2707
rect 4829 2698 4857 2704
rect 4877 2704 4885 2718
rect 4953 2684 4960 2727
rect 5056 2721 5064 2747
rect 5035 2714 5064 2721
rect 5035 2704 5041 2714
rect 5051 2704 5103 2706
rect 5178 2704 5186 2747
rect 5240 2722 5247 2778
rect 5261 2761 5269 2796
rect 5333 2761 5341 2796
rect 5267 2747 5269 2761
rect 5240 2716 5243 2722
rect 5023 2664 5051 2670
rect 5063 2700 5091 2704
rect 5160 2693 5186 2704
rect 5221 2710 5243 2716
rect 5221 2684 5229 2710
rect 5261 2704 5269 2747
rect 5455 2761 5463 2796
rect 5339 2725 5347 2747
rect 5397 2743 5403 2753
rect 5367 2737 5403 2743
rect 5340 2718 5365 2725
rect 5456 2721 5464 2747
rect 5536 2753 5544 2836
rect 5637 2830 5645 2836
rect 5687 2830 5699 2836
rect 5627 2816 5645 2830
rect 5673 2818 5695 2830
rect 5741 2822 5753 2856
rect 5637 2810 5645 2816
rect 5637 2802 5675 2810
rect 5693 2806 5723 2812
rect 5581 2788 5643 2796
rect 5297 2704 5349 2707
rect 5309 2698 5337 2704
rect 5357 2704 5365 2718
rect 5435 2714 5464 2721
rect 5435 2704 5441 2714
rect 5451 2704 5503 2706
rect 5423 2664 5451 2670
rect 5463 2700 5491 2704
rect 5536 2684 5544 2739
rect 5581 2704 5587 2788
rect 5693 2792 5699 2806
rect 5741 2798 5747 2816
rect 5655 2786 5699 2792
rect 5707 2792 5747 2798
rect 5626 2747 5653 2754
rect 5600 2736 5606 2741
rect 5600 2728 5634 2736
rect 5639 2720 5646 2728
rect 5707 2720 5713 2792
rect 5837 2868 5849 2882
rect 5897 2876 5909 2882
rect 5767 2784 5781 2792
rect 5773 2733 5787 2747
rect 5795 2733 5803 2796
rect 5823 2794 5829 2828
rect 5879 2804 5881 2806
rect 5867 2800 5881 2804
rect 5823 2788 5864 2794
rect 5855 2770 5864 2788
rect 5639 2714 5713 2720
rect 5787 2719 5803 2733
rect 5855 2720 5864 2758
rect 5875 2753 5881 2800
rect 5957 2868 5969 2882
rect 6017 2876 6029 2882
rect 5943 2794 5949 2828
rect 5999 2804 6001 2806
rect 5987 2800 6001 2804
rect 5943 2788 5984 2794
rect 5975 2770 5984 2788
rect 5639 2708 5646 2714
rect 5707 2712 5713 2714
rect 5671 2696 5692 2703
rect 5795 2704 5803 2719
rect 5620 2684 5627 2690
rect 5685 2684 5692 2696
rect 5742 2690 5753 2698
rect 5742 2684 5749 2690
rect 5620 2678 5633 2684
rect 5822 2714 5864 2720
rect 5822 2692 5829 2714
rect 5875 2708 5881 2739
rect 5975 2720 5984 2758
rect 5995 2753 6001 2800
rect 6077 2868 6089 2882
rect 6137 2876 6149 2882
rect 6207 2876 6219 2882
rect 6251 2876 6263 2882
rect 6063 2794 6069 2828
rect 6119 2804 6121 2806
rect 6107 2800 6121 2804
rect 6063 2788 6104 2794
rect 6095 2770 6104 2788
rect 5942 2714 5984 2720
rect 5867 2704 5881 2708
rect 5879 2702 5881 2704
rect 5942 2692 5949 2714
rect 5995 2708 6001 2739
rect 6095 2720 6104 2758
rect 6115 2753 6121 2800
rect 6291 2876 6303 2882
rect 6191 2761 6199 2796
rect 6191 2747 6193 2761
rect 6062 2714 6104 2720
rect 5987 2704 6001 2708
rect 5999 2702 6001 2704
rect 6062 2692 6069 2714
rect 6115 2708 6121 2739
rect 6107 2704 6121 2708
rect 6119 2702 6121 2704
rect 6191 2704 6199 2747
rect 6234 2722 6242 2836
rect 6331 2874 6343 2882
rect 6357 2876 6369 2882
rect 6401 2876 6413 2882
rect 6477 2876 6489 2882
rect 6535 2876 6547 2882
rect 6581 2876 6593 2882
rect 6647 2876 6659 2882
rect 6312 2753 6321 2796
rect 6307 2739 6321 2753
rect 6225 2714 6263 2722
rect 6251 2704 6263 2714
rect 6312 2704 6321 2739
rect 6378 2722 6386 2836
rect 6507 2822 6519 2856
rect 6561 2830 6573 2836
rect 6615 2830 6623 2836
rect 6565 2818 6587 2830
rect 6615 2816 6633 2830
rect 6513 2798 6519 2816
rect 6537 2806 6567 2812
rect 6615 2810 6623 2816
rect 6421 2761 6429 2796
rect 6427 2747 6429 2761
rect 6357 2714 6395 2722
rect 6357 2704 6369 2714
rect 6421 2704 6429 2747
rect 6191 2694 6201 2704
rect 4158 2658 4170 2664
rect 4208 2658 4220 2664
rect 4257 2658 4269 2664
rect 4410 2658 4422 2664
rect 4461 2658 4473 2664
rect 4523 2658 4535 2664
rect 4571 2658 4583 2664
rect 4629 2658 4641 2664
rect 4677 2658 4689 2664
rect 4737 2658 4749 2664
rect 4777 2658 4789 2664
rect 4837 2658 4849 2664
rect 4931 2658 4943 2664
rect 4971 2658 4983 2664
rect 5071 2658 5083 2664
rect 5120 2658 5132 2664
rect 5170 2658 5182 2664
rect 5239 2658 5251 2664
rect 5317 2658 5329 2664
rect 5471 2658 5483 2664
rect 5551 2658 5563 2664
rect 5601 2658 5613 2664
rect 5663 2658 5675 2664
rect 5711 2658 5723 2664
rect 5769 2658 5781 2664
rect 5837 2658 5849 2672
rect 5897 2658 5909 2672
rect 5957 2658 5969 2672
rect 6017 2658 6029 2672
rect 6077 2658 6089 2672
rect 6137 2658 6149 2672
rect 6419 2694 6429 2704
rect 6457 2733 6465 2796
rect 6479 2784 6493 2792
rect 6513 2792 6553 2798
rect 6473 2733 6487 2747
rect 6457 2719 6473 2733
rect 6547 2720 6553 2792
rect 6561 2792 6567 2806
rect 6585 2802 6623 2810
rect 6561 2786 6605 2792
rect 6617 2788 6679 2796
rect 6607 2747 6634 2754
rect 6654 2736 6660 2741
rect 6626 2728 6660 2736
rect 6614 2720 6621 2728
rect 6457 2704 6465 2719
rect 6547 2714 6621 2720
rect 6547 2712 6553 2714
rect 6614 2708 6621 2714
rect 6507 2690 6518 2698
rect 6511 2684 6518 2690
rect 6568 2696 6589 2703
rect 6673 2704 6679 2788
rect 6568 2684 6575 2696
rect 6633 2684 6640 2690
rect 6627 2678 6640 2684
rect 6221 2658 6233 2664
rect 6291 2658 6303 2664
rect 6331 2658 6343 2664
rect 6387 2658 6399 2664
rect 6479 2658 6491 2664
rect 6537 2658 6549 2664
rect 6585 2658 6597 2664
rect 6647 2658 6659 2664
rect 6742 2658 6802 3122
rect 4 2656 6802 2658
rect 6736 2644 6802 2656
rect 4 2642 6802 2644
rect 39 2636 51 2642
rect 97 2636 109 2642
rect 145 2636 157 2642
rect 207 2636 219 2642
rect 289 2636 301 2642
rect 359 2636 371 2642
rect 417 2636 429 2642
rect 465 2636 477 2642
rect 527 2636 539 2642
rect 598 2636 610 2642
rect 648 2636 660 2642
rect 187 2616 200 2622
rect 71 2610 78 2616
rect 67 2602 78 2610
rect 128 2604 135 2616
rect 193 2610 200 2616
rect 17 2581 25 2596
rect 128 2597 149 2604
rect 107 2586 113 2588
rect 174 2586 181 2592
rect 17 2567 33 2581
rect 107 2580 181 2586
rect 17 2504 25 2567
rect 33 2553 47 2567
rect 39 2508 53 2516
rect 107 2508 113 2580
rect 174 2572 181 2580
rect 186 2564 220 2572
rect 214 2559 220 2564
rect 167 2546 194 2553
rect 73 2502 113 2508
rect 121 2508 165 2514
rect 73 2484 79 2502
rect 121 2494 127 2508
rect 233 2512 239 2596
rect 177 2504 239 2512
rect 271 2553 279 2596
rect 311 2590 319 2616
rect 297 2584 319 2590
rect 507 2616 520 2622
rect 391 2610 398 2616
rect 387 2602 398 2610
rect 448 2604 455 2616
rect 513 2610 520 2616
rect 297 2578 300 2584
rect 271 2539 273 2553
rect 271 2504 279 2539
rect 293 2522 300 2578
rect 337 2581 345 2596
rect 448 2597 469 2604
rect 427 2586 433 2588
rect 494 2586 501 2592
rect 337 2567 353 2581
rect 427 2580 501 2586
rect 297 2516 300 2522
rect 297 2510 323 2516
rect 97 2488 127 2494
rect 145 2490 183 2498
rect 175 2484 183 2490
rect 67 2444 79 2478
rect 125 2470 147 2482
rect 175 2470 193 2484
rect 121 2464 133 2470
rect 175 2464 183 2470
rect 315 2464 323 2510
rect 337 2504 345 2567
rect 353 2553 367 2567
rect 359 2508 373 2516
rect 427 2508 433 2580
rect 494 2572 501 2580
rect 506 2564 540 2572
rect 534 2559 540 2564
rect 487 2546 514 2553
rect 393 2502 433 2508
rect 441 2508 485 2514
rect 393 2484 399 2502
rect 441 2494 447 2508
rect 553 2512 559 2596
rect 594 2596 620 2607
rect 679 2636 691 2642
rect 809 2636 821 2642
rect 594 2553 602 2596
rect 709 2588 721 2596
rect 697 2582 721 2588
rect 851 2636 863 2642
rect 891 2636 903 2642
rect 931 2636 943 2642
rect 971 2636 983 2642
rect 1011 2636 1023 2642
rect 1059 2636 1071 2642
rect 1117 2636 1129 2642
rect 1165 2636 1177 2642
rect 1227 2636 1239 2642
rect 1329 2636 1341 2642
rect 1207 2616 1220 2622
rect 1091 2610 1098 2616
rect 1087 2602 1098 2610
rect 1148 2604 1155 2616
rect 1213 2610 1220 2616
rect 779 2588 791 2596
rect 872 2590 884 2596
rect 912 2590 924 2596
rect 951 2590 963 2596
rect 992 2590 1004 2596
rect 866 2589 884 2590
rect 779 2582 803 2588
rect 497 2504 559 2512
rect 594 2504 602 2539
rect 697 2533 705 2582
rect 795 2533 803 2582
rect 865 2582 884 2589
rect 898 2582 924 2590
rect 938 2582 963 2590
rect 977 2582 1004 2590
rect 865 2561 872 2582
rect 898 2576 906 2582
rect 938 2576 946 2582
rect 977 2576 985 2582
rect 890 2564 906 2576
rect 930 2564 946 2576
rect 970 2564 985 2576
rect 1037 2581 1045 2596
rect 1148 2597 1169 2604
rect 1127 2586 1133 2588
rect 1194 2586 1201 2592
rect 867 2547 872 2561
rect 417 2488 447 2494
rect 465 2490 503 2498
rect 495 2484 503 2490
rect 387 2444 399 2478
rect 445 2470 467 2482
rect 495 2470 513 2484
rect 441 2464 453 2470
rect 495 2464 503 2470
rect 623 2498 663 2504
rect 651 2496 663 2498
rect 697 2464 705 2519
rect 795 2464 803 2519
rect 865 2518 872 2547
rect 898 2518 906 2564
rect 938 2518 946 2564
rect 977 2518 985 2564
rect 1037 2567 1053 2581
rect 1127 2580 1201 2586
rect 865 2510 883 2518
rect 898 2510 923 2518
rect 938 2510 963 2518
rect 977 2510 1003 2518
rect 871 2504 883 2510
rect 911 2504 923 2510
rect 951 2504 963 2510
rect 991 2504 1003 2510
rect 1037 2504 1045 2567
rect 1053 2553 1067 2567
rect 1059 2508 1073 2516
rect 37 2418 49 2424
rect 95 2418 107 2424
rect 141 2418 153 2424
rect 207 2418 219 2424
rect 289 2418 301 2424
rect 357 2418 369 2424
rect 415 2418 427 2424
rect 461 2418 473 2424
rect 527 2418 539 2424
rect 631 2418 643 2424
rect 677 2418 689 2424
rect 717 2418 729 2424
rect 771 2418 783 2424
rect 811 2418 823 2424
rect 1127 2508 1133 2580
rect 1194 2572 1201 2580
rect 1206 2564 1240 2572
rect 1234 2559 1240 2564
rect 1187 2546 1214 2553
rect 1093 2502 1133 2508
rect 1141 2508 1185 2514
rect 1093 2484 1099 2502
rect 1141 2494 1147 2508
rect 1253 2512 1259 2596
rect 1357 2636 1369 2642
rect 1397 2636 1409 2642
rect 1437 2636 1449 2642
rect 1551 2636 1563 2642
rect 1621 2636 1633 2642
rect 1683 2636 1695 2642
rect 1731 2636 1743 2642
rect 1789 2636 1801 2642
rect 1837 2636 1849 2642
rect 1897 2636 1909 2642
rect 1977 2636 1989 2642
rect 2077 2636 2089 2642
rect 2117 2636 2129 2642
rect 1299 2588 1311 2596
rect 1299 2582 1323 2588
rect 1315 2533 1323 2582
rect 1380 2573 1387 2616
rect 1456 2561 1464 2616
rect 1515 2582 1523 2596
rect 1543 2596 1571 2602
rect 1531 2593 1583 2596
rect 1640 2616 1653 2622
rect 1640 2610 1647 2616
rect 1705 2604 1712 2616
rect 1515 2575 1540 2582
rect 1197 2504 1259 2512
rect 1117 2488 1147 2494
rect 1165 2490 1203 2498
rect 1195 2484 1203 2490
rect 1087 2444 1099 2478
rect 1145 2470 1167 2482
rect 1195 2470 1213 2484
rect 1141 2464 1153 2470
rect 1195 2464 1203 2470
rect 1315 2464 1323 2519
rect 1380 2511 1387 2559
rect 1533 2553 1541 2575
rect 1380 2504 1397 2511
rect 851 2418 863 2424
rect 891 2418 903 2424
rect 931 2418 943 2424
rect 971 2418 983 2424
rect 1011 2418 1023 2424
rect 1057 2418 1069 2424
rect 1115 2418 1127 2424
rect 1161 2418 1173 2424
rect 1227 2418 1239 2424
rect 1291 2418 1303 2424
rect 1331 2418 1343 2424
rect 1456 2464 1464 2547
rect 1539 2504 1547 2539
rect 1601 2512 1607 2596
rect 1691 2597 1712 2604
rect 1762 2610 1769 2616
rect 1762 2602 1773 2610
rect 1659 2586 1666 2592
rect 1727 2586 1733 2588
rect 1659 2580 1733 2586
rect 1815 2581 1823 2596
rect 1659 2572 1666 2580
rect 1620 2564 1654 2572
rect 1620 2559 1626 2564
rect 1646 2546 1673 2553
rect 1601 2504 1663 2512
rect 1675 2508 1719 2514
rect 1657 2490 1695 2498
rect 1713 2494 1719 2508
rect 1727 2508 1733 2580
rect 1807 2567 1823 2581
rect 1793 2553 1807 2567
rect 1727 2502 1767 2508
rect 1787 2508 1801 2516
rect 1815 2504 1823 2567
rect 1856 2561 1864 2616
rect 1916 2561 1924 2616
rect 1969 2596 1997 2600
rect 2009 2630 2037 2636
rect 2177 2628 2189 2642
rect 2237 2628 2249 2642
rect 2297 2628 2309 2642
rect 2357 2628 2369 2642
rect 2421 2636 2433 2642
rect 2483 2636 2495 2642
rect 2531 2636 2543 2642
rect 2589 2636 2601 2642
rect 1957 2594 2009 2596
rect 2019 2586 2025 2596
rect 1996 2579 2025 2586
rect 1657 2484 1665 2490
rect 1713 2488 1743 2494
rect 1761 2484 1767 2502
rect 1647 2470 1665 2484
rect 1693 2470 1715 2482
rect 1657 2464 1665 2470
rect 1707 2464 1719 2470
rect 1761 2444 1773 2478
rect 1856 2464 1864 2547
rect 1916 2464 1924 2547
rect 1996 2553 2004 2579
rect 2077 2583 2083 2593
rect 2047 2577 2083 2583
rect 2100 2573 2107 2616
rect 2162 2586 2169 2608
rect 2219 2596 2221 2598
rect 2207 2592 2221 2596
rect 2162 2580 2204 2586
rect 1997 2504 2005 2539
rect 2100 2511 2107 2559
rect 2195 2542 2204 2580
rect 2215 2561 2221 2592
rect 2282 2586 2289 2608
rect 2339 2596 2341 2598
rect 2327 2592 2341 2596
rect 2282 2580 2324 2586
rect 2195 2512 2204 2530
rect 2100 2504 2117 2511
rect 1357 2418 1369 2424
rect 1437 2418 1449 2424
rect 1516 2418 1528 2424
rect 1566 2418 1578 2424
rect 1621 2418 1633 2424
rect 1687 2418 1699 2424
rect 1733 2418 1745 2424
rect 1791 2418 1803 2424
rect 1837 2418 1849 2424
rect 1897 2418 1909 2424
rect 1957 2418 1969 2424
rect 2027 2418 2039 2424
rect 2163 2506 2204 2512
rect 2163 2472 2169 2506
rect 2215 2500 2221 2547
rect 2315 2542 2324 2580
rect 2335 2561 2341 2592
rect 2440 2616 2453 2622
rect 2440 2610 2447 2616
rect 2505 2604 2512 2616
rect 2315 2512 2324 2530
rect 2283 2506 2324 2512
rect 2207 2496 2221 2500
rect 2219 2494 2221 2496
rect 2077 2418 2089 2424
rect 2177 2418 2189 2432
rect 2283 2472 2289 2506
rect 2335 2500 2341 2547
rect 2401 2512 2407 2596
rect 2491 2597 2512 2604
rect 2562 2610 2569 2616
rect 2562 2602 2573 2610
rect 2459 2586 2466 2592
rect 2657 2628 2669 2642
rect 2717 2628 2729 2642
rect 2527 2586 2533 2588
rect 2459 2580 2533 2586
rect 2615 2581 2623 2596
rect 2459 2572 2466 2580
rect 2420 2564 2454 2572
rect 2420 2559 2426 2564
rect 2446 2546 2473 2553
rect 2401 2504 2463 2512
rect 2475 2508 2519 2514
rect 2327 2496 2341 2500
rect 2339 2494 2341 2496
rect 2237 2418 2249 2424
rect 2297 2418 2309 2432
rect 2457 2490 2495 2498
rect 2513 2494 2519 2508
rect 2527 2508 2533 2580
rect 2607 2567 2623 2581
rect 2642 2586 2649 2608
rect 2699 2596 2701 2598
rect 2687 2592 2701 2596
rect 2642 2580 2684 2586
rect 2593 2553 2607 2567
rect 2527 2502 2567 2508
rect 2587 2508 2601 2516
rect 2615 2504 2623 2567
rect 2675 2542 2684 2580
rect 2695 2561 2701 2592
rect 2771 2636 2783 2642
rect 2811 2636 2823 2642
rect 2851 2628 2863 2642
rect 2911 2628 2923 2642
rect 3031 2636 3043 2642
rect 3111 2636 3123 2642
rect 3161 2636 3173 2642
rect 3223 2636 3235 2642
rect 3271 2636 3283 2642
rect 3329 2636 3341 2642
rect 3377 2636 3389 2642
rect 3417 2636 3429 2642
rect 3509 2636 3521 2642
rect 2793 2573 2800 2616
rect 2879 2596 2881 2598
rect 2879 2592 2893 2596
rect 2879 2561 2885 2592
rect 2931 2586 2938 2608
rect 2983 2630 3011 2636
rect 3023 2596 3051 2600
rect 2896 2580 2938 2586
rect 2995 2586 3001 2596
rect 3011 2594 3063 2596
rect 2675 2512 2684 2530
rect 2457 2484 2465 2490
rect 2513 2488 2543 2494
rect 2561 2484 2567 2502
rect 2447 2470 2465 2484
rect 2493 2470 2515 2482
rect 2457 2464 2465 2470
rect 2507 2464 2519 2470
rect 2561 2444 2573 2478
rect 2643 2506 2684 2512
rect 2643 2472 2649 2506
rect 2695 2500 2701 2547
rect 2793 2511 2800 2559
rect 2783 2504 2800 2511
rect 2687 2496 2701 2500
rect 2699 2494 2701 2496
rect 2357 2418 2369 2424
rect 2421 2418 2433 2424
rect 2487 2418 2499 2424
rect 2533 2418 2545 2424
rect 2591 2418 2603 2424
rect 2657 2418 2669 2432
rect 2717 2418 2729 2424
rect 2811 2418 2823 2424
rect 2879 2500 2885 2547
rect 2896 2542 2905 2580
rect 2995 2579 3024 2586
rect 2896 2512 2905 2530
rect 3016 2553 3024 2579
rect 3096 2561 3104 2616
rect 3180 2616 3193 2622
rect 3180 2610 3187 2616
rect 3245 2604 3252 2616
rect 2896 2506 2937 2512
rect 2879 2496 2893 2500
rect 2879 2494 2881 2496
rect 2931 2472 2937 2506
rect 3015 2504 3023 2539
rect 2851 2418 2863 2424
rect 2911 2418 2923 2432
rect 3096 2464 3104 2547
rect 3141 2512 3147 2596
rect 3231 2597 3252 2604
rect 3302 2610 3309 2616
rect 3302 2602 3313 2610
rect 3199 2586 3206 2592
rect 3267 2586 3273 2588
rect 3199 2580 3273 2586
rect 3355 2581 3363 2596
rect 3199 2572 3206 2580
rect 3160 2564 3194 2572
rect 3160 2559 3166 2564
rect 3186 2546 3213 2553
rect 3141 2504 3203 2512
rect 3215 2508 3259 2514
rect 3197 2490 3235 2498
rect 3253 2494 3259 2508
rect 3267 2508 3273 2580
rect 3347 2567 3363 2581
rect 3400 2573 3407 2616
rect 3537 2636 3549 2642
rect 3598 2636 3610 2642
rect 3698 2636 3710 2642
rect 3870 2636 3882 2642
rect 3917 2636 3929 2642
rect 4000 2636 4012 2642
rect 4050 2636 4062 2642
rect 3479 2588 3491 2596
rect 3479 2582 3503 2588
rect 3333 2553 3347 2567
rect 3267 2502 3307 2508
rect 3327 2508 3341 2516
rect 3355 2504 3363 2567
rect 3400 2511 3407 2559
rect 3495 2533 3503 2582
rect 3556 2561 3564 2616
rect 3646 2578 3664 2580
rect 3634 2569 3664 2578
rect 3746 2578 3764 2580
rect 3734 2569 3764 2578
rect 3577 2557 3623 2563
rect 3400 2504 3417 2511
rect 3197 2484 3205 2490
rect 3253 2488 3283 2494
rect 3301 2484 3307 2502
rect 3187 2470 3205 2484
rect 3233 2470 3255 2482
rect 3197 2464 3205 2470
rect 3247 2464 3259 2470
rect 3301 2444 3313 2478
rect 3495 2464 3503 2519
rect 3556 2464 3564 2547
rect 3577 2483 3583 2557
rect 3617 2547 3623 2557
rect 3656 2541 3664 2569
rect 3756 2541 3764 2569
rect 3816 2578 3834 2580
rect 3816 2569 3846 2578
rect 3909 2596 3937 2602
rect 3897 2593 3949 2596
rect 4111 2636 4123 2642
rect 4151 2636 4163 2642
rect 4251 2636 4263 2642
rect 4321 2636 4333 2642
rect 4383 2636 4395 2642
rect 4431 2636 4443 2642
rect 4489 2636 4501 2642
rect 4571 2636 4583 2642
rect 4671 2636 4683 2642
rect 4040 2596 4066 2607
rect 3957 2582 3965 2596
rect 3940 2575 3965 2582
rect 3816 2541 3824 2569
rect 3577 2477 3593 2483
rect 3658 2472 3665 2527
rect 3677 2483 3683 2533
rect 3939 2553 3947 2575
rect 3967 2557 3983 2563
rect 3677 2477 3693 2483
rect 3758 2472 3765 2527
rect 3618 2466 3665 2472
rect 3618 2464 3629 2466
rect 2981 2418 2993 2424
rect 3051 2418 3063 2424
rect 3111 2418 3123 2424
rect 3161 2418 3173 2424
rect 3227 2418 3239 2424
rect 3273 2418 3285 2424
rect 3331 2418 3343 2424
rect 3377 2418 3389 2424
rect 3471 2418 3483 2424
rect 3511 2418 3523 2424
rect 3657 2464 3665 2466
rect 3718 2466 3765 2472
rect 3718 2464 3729 2466
rect 3757 2464 3765 2466
rect 3815 2472 3822 2527
rect 3933 2504 3941 2539
rect 3977 2523 3983 2557
rect 4058 2553 4066 2596
rect 4133 2573 4140 2616
rect 4203 2630 4231 2636
rect 4243 2596 4271 2600
rect 4215 2586 4221 2596
rect 4231 2594 4283 2596
rect 4340 2616 4353 2622
rect 4340 2610 4347 2616
rect 4405 2604 4412 2616
rect 4215 2579 4244 2586
rect 3977 2517 4033 2523
rect 4058 2504 4066 2539
rect 4133 2511 4140 2559
rect 4236 2553 4244 2579
rect 4123 2504 4140 2511
rect 4235 2504 4243 2539
rect 4301 2512 4307 2596
rect 4391 2597 4412 2604
rect 4462 2610 4469 2616
rect 4462 2602 4473 2610
rect 4359 2586 4366 2592
rect 4427 2586 4433 2588
rect 4359 2580 4433 2586
rect 4515 2581 4523 2596
rect 4359 2572 4366 2580
rect 4320 2564 4354 2572
rect 4320 2559 4326 2564
rect 4346 2546 4373 2553
rect 4301 2504 4363 2512
rect 4375 2508 4419 2514
rect 3815 2466 3862 2472
rect 3815 2464 3823 2466
rect 3851 2464 3862 2466
rect 3537 2418 3549 2424
rect 3597 2418 3609 2424
rect 3637 2418 3649 2424
rect 3697 2418 3709 2424
rect 3737 2418 3749 2424
rect 3831 2418 3843 2424
rect 3871 2418 3883 2424
rect 3997 2498 4037 2504
rect 3997 2496 4009 2498
rect 3902 2418 3914 2424
rect 3952 2418 3964 2424
rect 4017 2418 4029 2424
rect 4151 2418 4163 2424
rect 4357 2490 4395 2498
rect 4413 2494 4419 2508
rect 4427 2508 4433 2580
rect 4507 2567 4523 2581
rect 4493 2553 4507 2567
rect 4427 2502 4467 2508
rect 4487 2508 4501 2516
rect 4515 2504 4523 2567
rect 4556 2561 4564 2616
rect 4623 2630 4651 2636
rect 4663 2596 4691 2600
rect 4737 2628 4749 2642
rect 4797 2628 4809 2642
rect 4859 2636 4871 2642
rect 4917 2636 4929 2642
rect 4965 2636 4977 2642
rect 5027 2636 5039 2642
rect 5077 2636 5089 2642
rect 5157 2636 5169 2642
rect 5277 2636 5289 2642
rect 5357 2636 5369 2642
rect 5397 2636 5409 2642
rect 4635 2586 4641 2596
rect 4651 2594 4703 2596
rect 4722 2586 4729 2608
rect 4779 2596 4781 2598
rect 4767 2592 4781 2596
rect 4635 2579 4664 2586
rect 4722 2580 4764 2586
rect 4357 2484 4365 2490
rect 4413 2488 4443 2494
rect 4461 2484 4467 2502
rect 4347 2470 4365 2484
rect 4393 2470 4415 2482
rect 4357 2464 4365 2470
rect 4407 2464 4419 2470
rect 4461 2444 4473 2478
rect 4556 2464 4564 2547
rect 4656 2553 4664 2579
rect 4655 2504 4663 2539
rect 4755 2542 4764 2580
rect 4775 2561 4781 2592
rect 5007 2616 5020 2622
rect 4891 2610 4898 2616
rect 4887 2602 4898 2610
rect 4948 2604 4955 2616
rect 5013 2610 5020 2616
rect 4837 2581 4845 2596
rect 4948 2597 4969 2604
rect 4927 2586 4933 2588
rect 4994 2586 5001 2592
rect 4837 2567 4853 2581
rect 4927 2580 5001 2586
rect 4755 2512 4764 2530
rect 4723 2506 4764 2512
rect 4201 2418 4213 2424
rect 4271 2418 4283 2424
rect 4321 2418 4333 2424
rect 4387 2418 4399 2424
rect 4433 2418 4445 2424
rect 4491 2418 4503 2424
rect 4571 2418 4583 2424
rect 4723 2472 4729 2506
rect 4775 2500 4781 2547
rect 4837 2504 4845 2567
rect 4853 2553 4867 2567
rect 4859 2508 4873 2516
rect 4767 2496 4781 2500
rect 4779 2494 4781 2496
rect 4621 2418 4633 2424
rect 4691 2418 4703 2424
rect 4737 2418 4749 2432
rect 4927 2508 4933 2580
rect 4994 2572 5001 2580
rect 5006 2564 5040 2572
rect 5034 2559 5040 2564
rect 4987 2546 5014 2553
rect 4893 2502 4933 2508
rect 4941 2508 4985 2514
rect 4893 2484 4899 2502
rect 4941 2494 4947 2508
rect 5053 2512 5059 2596
rect 5096 2561 5104 2616
rect 5149 2596 5177 2600
rect 5189 2630 5217 2636
rect 5269 2596 5297 2602
rect 5137 2594 5189 2596
rect 5199 2586 5205 2596
rect 5257 2593 5309 2596
rect 5451 2636 5463 2642
rect 5491 2636 5503 2642
rect 5517 2636 5529 2642
rect 5557 2636 5569 2642
rect 5597 2636 5609 2642
rect 5637 2636 5649 2642
rect 5677 2636 5689 2642
rect 5176 2579 5205 2586
rect 5317 2582 5325 2596
rect 4997 2504 5059 2512
rect 4917 2488 4947 2494
rect 4965 2490 5003 2498
rect 4995 2484 5003 2490
rect 4887 2444 4899 2478
rect 4945 2470 4967 2482
rect 4995 2470 5013 2484
rect 4941 2464 4953 2470
rect 4995 2464 5003 2470
rect 5096 2464 5104 2547
rect 5176 2553 5184 2579
rect 5300 2575 5325 2582
rect 5299 2553 5307 2575
rect 5380 2573 5387 2616
rect 5177 2504 5185 2539
rect 5293 2504 5301 2539
rect 5380 2511 5387 2559
rect 5473 2573 5480 2616
rect 5731 2636 5743 2642
rect 5771 2636 5783 2642
rect 5817 2636 5829 2642
rect 5971 2636 5983 2642
rect 6051 2636 6063 2642
rect 6099 2636 6111 2642
rect 6157 2636 6169 2642
rect 6205 2636 6217 2642
rect 6267 2636 6279 2642
rect 6352 2636 6364 2642
rect 6408 2636 6420 2642
rect 5536 2590 5548 2596
rect 5577 2590 5589 2596
rect 5616 2590 5628 2596
rect 5656 2590 5668 2596
rect 5536 2582 5563 2590
rect 5577 2582 5602 2590
rect 5616 2582 5642 2590
rect 5656 2589 5674 2590
rect 5656 2582 5675 2589
rect 5555 2576 5563 2582
rect 5594 2576 5602 2582
rect 5634 2576 5642 2582
rect 5555 2564 5570 2576
rect 5594 2564 5610 2576
rect 5634 2564 5650 2576
rect 5473 2511 5480 2559
rect 5555 2518 5563 2564
rect 5594 2518 5602 2564
rect 5634 2518 5642 2564
rect 5668 2561 5675 2582
rect 5753 2573 5760 2616
rect 5809 2596 5837 2602
rect 5797 2593 5849 2596
rect 5923 2630 5951 2636
rect 5963 2596 5991 2600
rect 5857 2582 5865 2596
rect 5840 2575 5865 2582
rect 5935 2586 5941 2596
rect 5951 2594 6003 2596
rect 5935 2579 5964 2586
rect 5668 2547 5673 2561
rect 5668 2518 5675 2547
rect 5380 2504 5397 2511
rect 4797 2418 4809 2424
rect 4857 2418 4869 2424
rect 4915 2418 4927 2424
rect 4961 2418 4973 2424
rect 5027 2418 5039 2424
rect 5077 2418 5089 2424
rect 5137 2418 5149 2424
rect 5207 2418 5219 2424
rect 5262 2418 5274 2424
rect 5312 2418 5324 2424
rect 5463 2504 5480 2511
rect 5537 2510 5563 2518
rect 5577 2510 5602 2518
rect 5617 2510 5642 2518
rect 5657 2510 5675 2518
rect 5753 2511 5760 2559
rect 5839 2553 5847 2575
rect 5956 2553 5964 2579
rect 6036 2561 6044 2616
rect 6247 2616 6260 2622
rect 6131 2610 6138 2616
rect 6127 2602 6138 2610
rect 6188 2604 6195 2616
rect 6253 2610 6260 2616
rect 6077 2581 6085 2596
rect 6188 2597 6209 2604
rect 6437 2636 6449 2642
rect 6477 2636 6489 2642
rect 6517 2636 6529 2642
rect 6580 2636 6592 2642
rect 6636 2636 6648 2642
rect 6167 2586 6173 2588
rect 6234 2586 6241 2592
rect 6077 2567 6093 2581
rect 6167 2580 6241 2586
rect 5537 2504 5549 2510
rect 5577 2504 5589 2510
rect 5617 2504 5629 2510
rect 5657 2504 5669 2510
rect 5743 2504 5760 2511
rect 5833 2504 5841 2539
rect 5955 2504 5963 2539
rect 5357 2418 5369 2424
rect 5491 2418 5503 2424
rect 5517 2418 5529 2424
rect 5557 2418 5569 2424
rect 5597 2418 5609 2424
rect 5637 2418 5649 2424
rect 5677 2418 5689 2424
rect 5771 2418 5783 2424
rect 5802 2418 5814 2424
rect 5852 2418 5864 2424
rect 6036 2464 6044 2547
rect 6077 2504 6085 2567
rect 6093 2553 6107 2567
rect 6099 2508 6113 2516
rect 6167 2508 6173 2580
rect 6234 2572 6241 2580
rect 6246 2564 6280 2572
rect 6274 2559 6280 2564
rect 6227 2546 6254 2553
rect 6133 2502 6173 2508
rect 6181 2508 6225 2514
rect 6133 2484 6139 2502
rect 6181 2494 6187 2508
rect 6293 2512 6299 2596
rect 6380 2553 6387 2596
rect 6459 2561 6468 2596
rect 6459 2547 6473 2561
rect 6536 2561 6544 2616
rect 6373 2516 6379 2539
rect 6237 2504 6299 2512
rect 6352 2510 6379 2516
rect 6352 2504 6364 2510
rect 6459 2504 6468 2547
rect 6157 2488 6187 2494
rect 6205 2490 6243 2498
rect 6235 2484 6243 2490
rect 6127 2444 6139 2478
rect 6185 2470 6207 2482
rect 6235 2470 6253 2484
rect 6181 2464 6193 2470
rect 6235 2464 6243 2470
rect 6343 2424 6371 2430
rect 6383 2496 6411 2502
rect 5921 2418 5933 2424
rect 5991 2418 6003 2424
rect 6051 2418 6063 2424
rect 6097 2418 6109 2424
rect 6155 2418 6167 2424
rect 6201 2418 6213 2424
rect 6267 2418 6279 2424
rect 6391 2418 6403 2424
rect 6437 2418 6449 2426
rect 6536 2464 6544 2547
rect 6613 2553 6620 2596
rect 6621 2516 6627 2539
rect 6621 2510 6648 2516
rect 6636 2504 6648 2510
rect 6477 2418 6489 2424
rect 6589 2496 6617 2502
rect 6629 2424 6657 2430
rect 6517 2418 6529 2424
rect 6597 2418 6609 2424
rect -62 2416 6736 2418
rect -62 2404 4 2416
rect -62 2402 6736 2404
rect -62 1938 -2 2402
rect 41 2396 53 2402
rect 107 2396 119 2402
rect 153 2396 165 2402
rect 211 2396 223 2402
rect 289 2396 301 2402
rect 371 2396 383 2402
rect 431 2396 443 2402
rect 511 2396 523 2402
rect 77 2350 85 2356
rect 127 2350 139 2356
rect 67 2336 85 2350
rect 113 2338 135 2350
rect 181 2342 193 2376
rect 77 2330 85 2336
rect 77 2322 115 2330
rect 133 2326 163 2332
rect 21 2308 83 2316
rect 21 2224 27 2308
rect 133 2312 139 2326
rect 181 2318 187 2336
rect 95 2306 139 2312
rect 147 2312 187 2318
rect 66 2267 93 2274
rect 40 2256 46 2261
rect 40 2248 74 2256
rect 79 2240 86 2248
rect 147 2240 153 2312
rect 207 2304 221 2312
rect 213 2253 227 2267
rect 235 2253 243 2316
rect 79 2234 153 2240
rect 227 2239 243 2253
rect 79 2228 86 2234
rect 147 2232 153 2234
rect 111 2216 132 2223
rect 235 2224 243 2239
rect 271 2281 279 2316
rect 315 2310 323 2356
rect 297 2304 323 2310
rect 297 2298 300 2304
rect 271 2267 273 2281
rect 271 2224 279 2267
rect 293 2242 300 2298
rect 356 2281 364 2316
rect 416 2273 424 2356
rect 542 2396 554 2402
rect 592 2396 604 2402
rect 667 2396 679 2402
rect 711 2396 723 2402
rect 737 2396 749 2402
rect 777 2396 789 2402
rect 837 2396 849 2402
rect 877 2396 889 2402
rect 937 2396 949 2402
rect 995 2396 1007 2402
rect 1041 2396 1053 2402
rect 1107 2396 1119 2402
rect 1157 2396 1169 2402
rect 1241 2396 1253 2402
rect 1307 2396 1319 2402
rect 1353 2396 1365 2402
rect 1411 2396 1423 2402
rect 1491 2396 1503 2402
rect 483 2309 500 2316
rect 297 2236 300 2242
rect 297 2230 319 2236
rect 60 2204 67 2210
rect 125 2204 132 2216
rect 182 2210 193 2218
rect 182 2204 189 2210
rect 60 2198 73 2204
rect 311 2204 319 2230
rect 356 2224 364 2267
rect 493 2261 500 2309
rect 573 2281 581 2316
rect 651 2281 659 2316
rect 416 2204 424 2259
rect 493 2204 500 2247
rect 579 2245 587 2267
rect 651 2267 653 2281
rect 580 2238 605 2245
rect 537 2224 589 2227
rect 41 2178 53 2184
rect 103 2178 115 2184
rect 151 2178 163 2184
rect 209 2178 221 2184
rect 289 2178 301 2184
rect 371 2178 383 2184
rect 431 2178 443 2184
rect 549 2218 577 2224
rect 597 2224 605 2238
rect 651 2224 659 2267
rect 694 2242 702 2356
rect 758 2354 769 2356
rect 797 2354 805 2356
rect 758 2348 805 2354
rect 798 2293 805 2348
rect 857 2301 865 2356
rect 967 2342 979 2376
rect 1021 2350 1033 2356
rect 1075 2350 1083 2356
rect 1025 2338 1047 2350
rect 1075 2336 1093 2350
rect 973 2318 979 2336
rect 997 2326 1027 2332
rect 1075 2330 1083 2336
rect 796 2251 804 2279
rect 685 2234 723 2242
rect 711 2224 723 2234
rect 651 2214 661 2224
rect 774 2242 804 2251
rect 786 2240 804 2242
rect 857 2238 865 2287
rect 917 2253 925 2316
rect 939 2304 953 2312
rect 973 2312 1013 2318
rect 933 2253 947 2267
rect 917 2239 933 2253
rect 1007 2240 1013 2312
rect 1021 2312 1027 2326
rect 1045 2322 1083 2330
rect 1021 2306 1065 2312
rect 1077 2308 1139 2316
rect 1067 2267 1094 2274
rect 1114 2256 1120 2261
rect 1086 2248 1120 2256
rect 1074 2240 1081 2248
rect 857 2232 881 2238
rect 869 2224 881 2232
rect 917 2224 925 2239
rect 1007 2234 1081 2240
rect 1007 2232 1013 2234
rect 1074 2228 1081 2234
rect 967 2210 978 2218
rect 971 2204 978 2210
rect 1028 2216 1049 2223
rect 1133 2224 1139 2308
rect 1176 2273 1184 2356
rect 1277 2350 1285 2356
rect 1327 2350 1339 2356
rect 1267 2336 1285 2350
rect 1313 2338 1335 2350
rect 1381 2342 1393 2376
rect 1277 2330 1285 2336
rect 1277 2322 1315 2330
rect 1333 2326 1363 2332
rect 1221 2308 1283 2316
rect 1028 2204 1035 2216
rect 1093 2204 1100 2210
rect 1087 2198 1100 2204
rect 1176 2204 1184 2259
rect 1221 2224 1227 2308
rect 1333 2312 1339 2326
rect 1381 2318 1387 2336
rect 1295 2306 1339 2312
rect 1347 2312 1387 2318
rect 1266 2267 1293 2274
rect 1240 2256 1246 2261
rect 1240 2248 1274 2256
rect 1279 2240 1286 2248
rect 1347 2240 1353 2312
rect 1517 2396 1529 2402
rect 1587 2396 1599 2402
rect 1407 2304 1421 2312
rect 1413 2253 1427 2267
rect 1435 2253 1443 2316
rect 1476 2273 1484 2356
rect 1642 2396 1654 2402
rect 1692 2396 1704 2402
rect 1791 2396 1803 2402
rect 1871 2396 1883 2402
rect 1921 2396 1933 2402
rect 1991 2396 2003 2402
rect 2051 2396 2063 2402
rect 2101 2396 2113 2402
rect 2167 2396 2179 2402
rect 2213 2396 2225 2402
rect 2271 2396 2283 2402
rect 2371 2396 2383 2402
rect 1557 2281 1565 2316
rect 1673 2281 1681 2316
rect 1763 2309 1780 2316
rect 1843 2309 1860 2316
rect 1279 2234 1353 2240
rect 1427 2239 1443 2253
rect 1279 2228 1286 2234
rect 1347 2232 1353 2234
rect 1311 2216 1332 2223
rect 1435 2224 1443 2239
rect 1260 2204 1267 2210
rect 1325 2204 1332 2216
rect 1382 2210 1393 2218
rect 1382 2204 1389 2210
rect 1260 2198 1273 2204
rect 1476 2204 1484 2259
rect 1556 2241 1564 2267
rect 1679 2245 1687 2267
rect 1773 2261 1780 2309
rect 1853 2261 1860 2309
rect 1955 2281 1963 2316
rect 1556 2234 1585 2241
rect 1680 2238 1705 2245
rect 1517 2224 1569 2226
rect 1579 2224 1585 2234
rect 1637 2224 1689 2227
rect 1529 2220 1557 2224
rect 1569 2184 1597 2190
rect 1649 2218 1677 2224
rect 1697 2224 1705 2238
rect 1773 2204 1780 2247
rect 1853 2204 1860 2247
rect 1956 2241 1964 2267
rect 2036 2273 2044 2356
rect 2137 2350 2145 2356
rect 2187 2350 2199 2356
rect 2127 2336 2145 2350
rect 2173 2338 2195 2350
rect 2241 2342 2253 2376
rect 2137 2330 2145 2336
rect 2137 2322 2175 2330
rect 2193 2326 2223 2332
rect 2081 2308 2143 2316
rect 1935 2234 1964 2241
rect 1935 2224 1941 2234
rect 1951 2224 2003 2226
rect 471 2178 483 2184
rect 511 2178 523 2184
rect 557 2178 569 2184
rect 681 2178 693 2184
rect 738 2178 750 2184
rect 839 2178 851 2184
rect 939 2178 951 2184
rect 997 2178 1009 2184
rect 1045 2178 1057 2184
rect 1107 2178 1119 2184
rect 1157 2178 1169 2184
rect 1241 2178 1253 2184
rect 1303 2178 1315 2184
rect 1351 2178 1363 2184
rect 1409 2178 1421 2184
rect 1491 2178 1503 2184
rect 1537 2178 1549 2184
rect 1657 2178 1669 2184
rect 1751 2178 1763 2184
rect 1791 2178 1803 2184
rect 1923 2184 1951 2190
rect 1963 2220 1991 2224
rect 2036 2204 2044 2259
rect 2081 2224 2087 2308
rect 2193 2312 2199 2326
rect 2241 2318 2247 2336
rect 2155 2306 2199 2312
rect 2207 2312 2247 2318
rect 2126 2267 2153 2274
rect 2100 2256 2106 2261
rect 2100 2248 2134 2256
rect 2139 2240 2146 2248
rect 2207 2240 2213 2312
rect 2267 2304 2281 2312
rect 2273 2253 2287 2267
rect 2295 2253 2303 2316
rect 2402 2396 2414 2402
rect 2452 2396 2464 2402
rect 2531 2396 2543 2402
rect 2571 2396 2583 2402
rect 2651 2396 2663 2402
rect 2702 2396 2714 2402
rect 2752 2396 2764 2402
rect 2851 2396 2863 2402
rect 2897 2396 2909 2402
rect 2955 2396 2967 2402
rect 3001 2396 3013 2402
rect 3067 2396 3079 2402
rect 3122 2396 3134 2402
rect 3172 2396 3184 2402
rect 2515 2354 2523 2356
rect 2551 2354 2562 2356
rect 2515 2348 2562 2354
rect 2467 2337 2483 2343
rect 2343 2309 2360 2316
rect 2139 2234 2213 2240
rect 2287 2239 2303 2253
rect 2139 2228 2146 2234
rect 2207 2232 2213 2234
rect 2171 2216 2192 2223
rect 2295 2224 2303 2239
rect 2120 2204 2127 2210
rect 2185 2204 2192 2216
rect 2242 2210 2253 2218
rect 2242 2204 2249 2210
rect 2120 2198 2133 2204
rect 2353 2261 2360 2309
rect 2433 2281 2441 2316
rect 2477 2303 2483 2337
rect 2477 2297 2503 2303
rect 2353 2204 2360 2247
rect 2439 2245 2447 2267
rect 2440 2238 2465 2245
rect 2397 2224 2449 2227
rect 2409 2218 2437 2224
rect 2457 2224 2465 2238
rect 2497 2223 2503 2297
rect 2515 2293 2522 2348
rect 2671 2322 2683 2324
rect 2643 2316 2683 2322
rect 2927 2342 2939 2376
rect 2981 2350 2993 2356
rect 3035 2350 3043 2356
rect 2985 2338 3007 2350
rect 3035 2336 3053 2350
rect 2933 2318 2939 2336
rect 2957 2326 2987 2332
rect 3035 2330 3043 2336
rect 2597 2287 2603 2293
rect 2516 2251 2524 2279
rect 2614 2281 2622 2316
rect 2733 2281 2741 2316
rect 2823 2309 2840 2316
rect 2557 2263 2563 2273
rect 2557 2257 2593 2263
rect 2516 2242 2546 2251
rect 2516 2240 2534 2242
rect 2497 2217 2513 2223
rect 2614 2224 2622 2267
rect 2739 2245 2747 2267
rect 2833 2261 2840 2309
rect 2877 2253 2885 2316
rect 2899 2304 2913 2312
rect 2933 2312 2973 2318
rect 2893 2253 2907 2267
rect 2740 2238 2765 2245
rect 2697 2224 2749 2227
rect 2614 2213 2640 2224
rect 1831 2178 1843 2184
rect 1871 2178 1883 2184
rect 1971 2178 1983 2184
rect 2051 2178 2063 2184
rect 2101 2178 2113 2184
rect 2163 2178 2175 2184
rect 2211 2178 2223 2184
rect 2269 2178 2281 2184
rect 2331 2178 2343 2184
rect 2371 2178 2383 2184
rect 2417 2178 2429 2184
rect 2570 2178 2582 2184
rect 2709 2218 2737 2224
rect 2757 2224 2765 2238
rect 2833 2204 2840 2247
rect 2877 2239 2893 2253
rect 2967 2240 2973 2312
rect 2981 2312 2987 2326
rect 3005 2322 3043 2330
rect 3241 2396 3253 2402
rect 3311 2396 3323 2402
rect 3391 2396 3403 2402
rect 3451 2396 3463 2402
rect 3531 2396 3543 2402
rect 3581 2396 3593 2402
rect 3647 2396 3659 2402
rect 3693 2396 3705 2402
rect 3751 2396 3763 2402
rect 3797 2396 3809 2402
rect 3837 2396 3849 2402
rect 2981 2306 3025 2312
rect 3037 2308 3099 2316
rect 3027 2267 3054 2274
rect 3074 2256 3080 2261
rect 3046 2248 3080 2256
rect 3034 2240 3041 2248
rect 2877 2224 2885 2239
rect 2967 2234 3041 2240
rect 2967 2232 2973 2234
rect 3034 2228 3041 2234
rect 2927 2210 2938 2218
rect 2931 2204 2938 2210
rect 2988 2216 3009 2223
rect 3093 2224 3099 2308
rect 3153 2281 3161 2316
rect 3275 2281 3283 2316
rect 3363 2309 3380 2316
rect 3159 2245 3167 2267
rect 3160 2238 3185 2245
rect 3276 2241 3284 2267
rect 3373 2261 3380 2309
rect 3436 2273 3444 2356
rect 3617 2350 3625 2356
rect 3667 2350 3679 2356
rect 3607 2336 3625 2350
rect 3653 2338 3675 2350
rect 3721 2342 3733 2376
rect 3617 2330 3625 2336
rect 3617 2322 3655 2330
rect 3673 2326 3703 2332
rect 3503 2309 3520 2316
rect 3467 2297 3483 2303
rect 2988 2204 2995 2216
rect 3053 2204 3060 2210
rect 3047 2198 3060 2204
rect 3117 2224 3169 2227
rect 3129 2218 3157 2224
rect 3177 2224 3185 2238
rect 3255 2234 3284 2241
rect 3255 2224 3261 2234
rect 3271 2224 3323 2226
rect 3243 2184 3271 2190
rect 3283 2220 3311 2224
rect 3373 2204 3380 2247
rect 3436 2204 3444 2259
rect 3477 2243 3483 2297
rect 3513 2261 3520 2309
rect 3561 2308 3623 2316
rect 3477 2237 3493 2243
rect 3513 2204 3520 2247
rect 3561 2224 3567 2308
rect 3673 2312 3679 2326
rect 3721 2318 3727 2336
rect 3635 2306 3679 2312
rect 3687 2312 3727 2318
rect 3606 2267 3633 2274
rect 3580 2256 3586 2261
rect 3580 2248 3614 2256
rect 3619 2240 3626 2248
rect 3687 2240 3693 2312
rect 3877 2396 3889 2402
rect 3917 2396 3929 2402
rect 3747 2304 3761 2312
rect 3753 2253 3767 2267
rect 3775 2253 3783 2316
rect 3817 2301 3825 2356
rect 3898 2354 3909 2356
rect 3997 2388 4009 2402
rect 4057 2396 4069 2402
rect 3937 2354 3945 2356
rect 3898 2348 3945 2354
rect 3619 2234 3693 2240
rect 3767 2239 3783 2253
rect 3619 2228 3626 2234
rect 3687 2232 3693 2234
rect 2618 2178 2630 2184
rect 2668 2178 2680 2184
rect 2717 2178 2729 2184
rect 2811 2178 2823 2184
rect 2851 2178 2863 2184
rect 2899 2178 2911 2184
rect 2957 2178 2969 2184
rect 3005 2178 3017 2184
rect 3067 2178 3079 2184
rect 3137 2178 3149 2184
rect 3291 2178 3303 2184
rect 3351 2178 3363 2184
rect 3391 2178 3403 2184
rect 3451 2178 3463 2184
rect 3651 2216 3672 2223
rect 3775 2224 3783 2239
rect 3817 2238 3825 2287
rect 3938 2293 3945 2348
rect 3983 2314 3989 2348
rect 4039 2324 4041 2326
rect 4027 2320 4041 2324
rect 3983 2308 4024 2314
rect 3936 2251 3944 2279
rect 4015 2290 4024 2308
rect 3817 2232 3841 2238
rect 3829 2224 3841 2232
rect 3600 2204 3607 2210
rect 3665 2204 3672 2216
rect 3722 2210 3733 2218
rect 3722 2204 3729 2210
rect 3600 2198 3613 2204
rect 3914 2242 3944 2251
rect 3926 2240 3944 2242
rect 4015 2240 4024 2278
rect 4035 2273 4041 2320
rect 4117 2388 4129 2402
rect 4177 2396 4189 2402
rect 4103 2314 4109 2348
rect 4159 2324 4161 2326
rect 4147 2320 4161 2324
rect 4103 2308 4144 2314
rect 4135 2290 4144 2308
rect 3982 2234 4024 2240
rect 3982 2212 3989 2234
rect 4035 2228 4041 2259
rect 4135 2240 4144 2278
rect 4155 2273 4161 2320
rect 4237 2388 4249 2402
rect 4297 2396 4309 2402
rect 4359 2396 4371 2402
rect 4471 2396 4483 2402
rect 4223 2314 4229 2348
rect 4279 2324 4281 2326
rect 4267 2320 4281 2324
rect 4223 2308 4264 2314
rect 4255 2290 4264 2308
rect 4102 2234 4144 2240
rect 4027 2224 4041 2228
rect 4039 2222 4041 2224
rect 4102 2212 4109 2234
rect 4155 2228 4161 2259
rect 4255 2240 4264 2278
rect 4275 2273 4281 2320
rect 4337 2310 4345 2356
rect 4517 2388 4529 2402
rect 4577 2396 4589 2402
rect 4337 2304 4363 2310
rect 4360 2298 4363 2304
rect 4222 2234 4264 2240
rect 4147 2224 4161 2228
rect 4159 2222 4161 2224
rect 4222 2212 4229 2234
rect 4275 2228 4281 2259
rect 4360 2242 4367 2298
rect 4381 2281 4389 2316
rect 4443 2309 4460 2316
rect 4387 2267 4389 2281
rect 4360 2236 4363 2242
rect 4267 2224 4281 2228
rect 4279 2222 4281 2224
rect 4341 2230 4363 2236
rect 4341 2204 4349 2230
rect 4381 2224 4389 2267
rect 4453 2261 4460 2309
rect 4503 2314 4509 2348
rect 4559 2324 4561 2326
rect 4547 2320 4561 2324
rect 4503 2308 4544 2314
rect 4535 2290 4544 2308
rect 3491 2178 3503 2184
rect 3531 2178 3543 2184
rect 3581 2178 3593 2184
rect 3643 2178 3655 2184
rect 3691 2178 3703 2184
rect 3749 2178 3761 2184
rect 3799 2178 3811 2184
rect 3878 2178 3890 2184
rect 3997 2178 4009 2192
rect 4057 2178 4069 2192
rect 4117 2178 4129 2192
rect 4177 2178 4189 2192
rect 4237 2178 4249 2192
rect 4297 2178 4309 2192
rect 4453 2204 4460 2247
rect 4535 2240 4544 2278
rect 4555 2273 4561 2320
rect 4631 2396 4643 2402
rect 4691 2388 4703 2402
rect 4757 2388 4769 2402
rect 4817 2396 4829 2402
rect 4659 2324 4661 2326
rect 4659 2320 4673 2324
rect 4659 2273 4665 2320
rect 4711 2314 4717 2348
rect 4676 2308 4717 2314
rect 4743 2314 4749 2348
rect 4799 2324 4801 2326
rect 4787 2320 4801 2324
rect 4743 2308 4784 2314
rect 4676 2290 4685 2308
rect 4502 2234 4544 2240
rect 4502 2212 4509 2234
rect 4555 2228 4561 2259
rect 4547 2224 4561 2228
rect 4559 2222 4561 2224
rect 4359 2178 4371 2184
rect 4431 2178 4443 2184
rect 4471 2178 4483 2184
rect 4517 2178 4529 2192
rect 4577 2178 4589 2192
rect 4659 2228 4665 2259
rect 4676 2240 4685 2278
rect 4775 2290 4784 2308
rect 4775 2240 4784 2278
rect 4795 2273 4801 2320
rect 4857 2396 4869 2402
rect 4957 2388 4969 2402
rect 5017 2396 5029 2402
rect 5111 2396 5123 2402
rect 5157 2396 5169 2402
rect 5217 2396 5229 2402
rect 5287 2396 5299 2402
rect 4880 2309 4897 2316
rect 4943 2314 4949 2348
rect 4999 2324 5001 2326
rect 4987 2320 5001 2324
rect 4880 2261 4887 2309
rect 4943 2308 4984 2314
rect 4676 2234 4718 2240
rect 4659 2224 4673 2228
rect 4659 2222 4661 2224
rect 4711 2212 4718 2234
rect 4742 2234 4784 2240
rect 4742 2212 4749 2234
rect 4795 2228 4801 2259
rect 4975 2290 4984 2308
rect 4787 2224 4801 2228
rect 4799 2222 4801 2224
rect 4880 2204 4887 2247
rect 4975 2240 4984 2278
rect 4995 2273 5001 2320
rect 5131 2322 5143 2324
rect 5103 2316 5143 2322
rect 5074 2281 5082 2316
rect 5176 2273 5184 2356
rect 5351 2396 5363 2402
rect 5411 2388 5423 2402
rect 5477 2388 5489 2402
rect 5537 2396 5549 2402
rect 5379 2324 5381 2326
rect 5379 2320 5393 2324
rect 5257 2281 5265 2316
rect 4942 2234 4984 2240
rect 4942 2212 4949 2234
rect 4995 2228 5001 2259
rect 4987 2224 5001 2228
rect 4631 2178 4643 2192
rect 4691 2178 4703 2192
rect 4757 2178 4769 2192
rect 4817 2178 4829 2192
rect 4999 2222 5001 2224
rect 5074 2224 5082 2267
rect 5074 2213 5100 2224
rect 4857 2178 4869 2184
rect 4897 2178 4909 2184
rect 4957 2178 4969 2192
rect 5017 2178 5029 2192
rect 5176 2204 5184 2259
rect 5256 2241 5264 2267
rect 5379 2273 5385 2320
rect 5431 2314 5437 2348
rect 5396 2308 5437 2314
rect 5463 2314 5469 2348
rect 5519 2324 5521 2326
rect 5507 2320 5521 2324
rect 5463 2308 5504 2314
rect 5396 2290 5405 2308
rect 5256 2234 5285 2241
rect 5217 2224 5269 2226
rect 5279 2224 5285 2234
rect 5078 2178 5090 2184
rect 5128 2178 5140 2184
rect 5229 2220 5257 2224
rect 5269 2184 5297 2190
rect 5379 2228 5385 2259
rect 5396 2240 5405 2278
rect 5495 2290 5504 2308
rect 5495 2240 5504 2278
rect 5515 2273 5521 2320
rect 5597 2388 5609 2402
rect 5657 2396 5669 2402
rect 5731 2396 5743 2402
rect 5771 2396 5783 2402
rect 5831 2396 5843 2402
rect 5871 2396 5883 2402
rect 5931 2396 5943 2402
rect 6031 2396 6043 2402
rect 6091 2396 6103 2402
rect 5583 2314 5589 2348
rect 5639 2324 5641 2326
rect 5627 2320 5641 2324
rect 5583 2308 5624 2314
rect 5615 2290 5624 2308
rect 5396 2234 5438 2240
rect 5379 2224 5393 2228
rect 5379 2222 5381 2224
rect 5431 2212 5438 2234
rect 5462 2234 5504 2240
rect 5462 2212 5469 2234
rect 5515 2228 5521 2259
rect 5615 2240 5624 2278
rect 5635 2273 5641 2320
rect 5715 2354 5723 2356
rect 5751 2354 5762 2356
rect 5715 2348 5762 2354
rect 5815 2354 5823 2356
rect 5851 2354 5862 2356
rect 5815 2348 5862 2354
rect 5715 2293 5722 2348
rect 5797 2287 5803 2333
rect 5815 2293 5822 2348
rect 5582 2234 5624 2240
rect 5507 2224 5521 2228
rect 5519 2222 5521 2224
rect 5582 2212 5589 2234
rect 5635 2228 5641 2259
rect 5716 2251 5724 2279
rect 5816 2251 5824 2279
rect 5916 2273 5924 2356
rect 5983 2390 6011 2396
rect 6023 2318 6051 2324
rect 6151 2388 6163 2402
rect 6211 2396 6223 2402
rect 6119 2324 6121 2326
rect 6119 2320 6133 2324
rect 5992 2310 6004 2316
rect 5992 2304 6019 2310
rect 6013 2281 6019 2304
rect 5716 2242 5746 2251
rect 5716 2240 5734 2242
rect 5627 2224 5641 2228
rect 5639 2222 5641 2224
rect 5157 2178 5169 2184
rect 5237 2178 5249 2184
rect 5351 2178 5363 2192
rect 5411 2178 5423 2192
rect 5477 2178 5489 2192
rect 5537 2178 5549 2192
rect 5597 2178 5609 2192
rect 5657 2178 5669 2192
rect 5816 2242 5846 2251
rect 5816 2240 5834 2242
rect 5916 2204 5924 2259
rect 6020 2224 6027 2267
rect 6119 2273 6125 2320
rect 6171 2314 6177 2348
rect 6271 2388 6283 2402
rect 6317 2396 6329 2402
rect 6382 2396 6394 2402
rect 6432 2396 6444 2402
rect 6239 2324 6241 2326
rect 6239 2320 6253 2324
rect 6136 2308 6177 2314
rect 6136 2290 6145 2308
rect 5770 2178 5782 2184
rect 5870 2178 5882 2184
rect 5931 2178 5943 2184
rect 5992 2178 6004 2184
rect 6048 2178 6060 2184
rect 6119 2228 6125 2259
rect 6136 2240 6145 2278
rect 6239 2273 6245 2320
rect 6291 2314 6297 2348
rect 6256 2308 6297 2314
rect 6256 2290 6265 2308
rect 6136 2234 6178 2240
rect 6119 2224 6133 2228
rect 6119 2222 6121 2224
rect 6171 2212 6178 2234
rect 6239 2228 6245 2259
rect 6256 2240 6265 2278
rect 6336 2273 6344 2356
rect 6477 2396 6489 2402
rect 6517 2396 6529 2402
rect 6577 2396 6589 2402
rect 6657 2396 6669 2402
rect 6447 2337 6463 2343
rect 6413 2281 6421 2316
rect 6256 2234 6298 2240
rect 6239 2224 6253 2228
rect 6239 2222 6241 2224
rect 6291 2212 6298 2234
rect 6336 2204 6344 2259
rect 6419 2245 6427 2267
rect 6420 2238 6445 2245
rect 6377 2224 6429 2227
rect 6091 2178 6103 2192
rect 6151 2178 6163 2192
rect 6211 2178 6223 2192
rect 6271 2178 6283 2192
rect 6389 2218 6417 2224
rect 6437 2224 6445 2238
rect 6457 2243 6463 2337
rect 6497 2301 6505 2356
rect 6557 2322 6569 2324
rect 6557 2316 6597 2322
rect 6457 2237 6473 2243
rect 6497 2238 6505 2287
rect 6618 2281 6626 2316
rect 6676 2273 6684 2356
rect 6497 2232 6521 2238
rect 6509 2224 6521 2232
rect 6618 2224 6626 2267
rect 6600 2213 6626 2224
rect 6676 2204 6684 2259
rect 6317 2178 6329 2184
rect 6397 2178 6409 2184
rect 6479 2178 6491 2184
rect 6560 2178 6572 2184
rect 6610 2178 6622 2184
rect 6657 2178 6669 2184
rect 6742 2178 6802 2642
rect 4 2176 6802 2178
rect 6736 2164 6802 2176
rect 4 2162 6802 2164
rect 31 2156 43 2162
rect 71 2156 83 2162
rect 149 2156 161 2162
rect 250 2156 262 2162
rect 350 2156 362 2162
rect 429 2156 441 2162
rect 53 2093 60 2136
rect 119 2108 131 2116
rect 87 2097 103 2103
rect 119 2102 143 2108
rect 53 2031 60 2079
rect 43 2024 60 2031
rect 97 2007 103 2097
rect 135 2053 143 2102
rect 196 2098 214 2100
rect 135 1984 143 2039
rect 177 2023 183 2093
rect 196 2089 226 2098
rect 296 2098 314 2100
rect 196 2061 204 2089
rect 167 2017 183 2023
rect 195 1992 202 2047
rect 277 2003 283 2093
rect 296 2089 326 2098
rect 458 2156 470 2162
rect 571 2156 583 2162
rect 611 2156 623 2162
rect 657 2156 669 2162
rect 738 2156 750 2162
rect 837 2156 849 2162
rect 877 2156 889 2162
rect 969 2156 981 2162
rect 296 2061 304 2089
rect 267 1997 283 2003
rect 295 1992 302 2047
rect 377 2003 383 2113
rect 399 2108 411 2116
rect 399 2102 423 2108
rect 415 2053 423 2102
rect 527 2117 573 2123
rect 506 2098 524 2100
rect 494 2089 524 2098
rect 516 2061 524 2089
rect 557 2097 573 2103
rect 367 1997 383 2003
rect 195 1986 242 1992
rect 195 1984 203 1986
rect 71 1938 83 1944
rect 231 1984 242 1986
rect 295 1986 342 1992
rect 295 1984 303 1986
rect 331 1984 342 1986
rect 415 1984 423 2039
rect 518 1992 525 2047
rect 557 2043 563 2097
rect 593 2093 600 2136
rect 649 2116 677 2122
rect 637 2113 689 2116
rect 697 2102 705 2116
rect 680 2095 705 2102
rect 786 2098 804 2100
rect 547 2037 563 2043
rect 593 2031 600 2079
rect 679 2073 687 2095
rect 774 2089 804 2098
rect 860 2093 867 2136
rect 1017 2148 1029 2162
rect 1077 2148 1089 2162
rect 1141 2156 1153 2162
rect 1203 2156 1215 2162
rect 1251 2156 1263 2162
rect 1309 2156 1321 2162
rect 1357 2156 1369 2162
rect 1437 2156 1449 2162
rect 1591 2156 1603 2162
rect 1691 2156 1703 2162
rect 1751 2156 1763 2162
rect 1791 2156 1803 2162
rect 1871 2156 1883 2162
rect 939 2108 951 2116
rect 939 2102 963 2108
rect 796 2061 804 2089
rect 478 1986 525 1992
rect 478 1984 489 1986
rect 111 1938 123 1944
rect 151 1938 163 1944
rect 211 1938 223 1944
rect 251 1938 263 1944
rect 311 1938 323 1944
rect 351 1938 363 1944
rect 391 1938 403 1944
rect 431 1938 443 1944
rect 517 1984 525 1986
rect 583 2024 600 2031
rect 673 2024 681 2059
rect 457 1938 469 1944
rect 497 1938 509 1944
rect 611 1938 623 1944
rect 798 1992 805 2047
rect 860 2031 867 2079
rect 955 2053 963 2102
rect 1002 2106 1009 2128
rect 1059 2116 1061 2118
rect 1047 2112 1061 2116
rect 1002 2100 1044 2106
rect 1035 2062 1044 2100
rect 1055 2081 1061 2112
rect 1160 2136 1173 2142
rect 1160 2130 1167 2136
rect 1225 2124 1232 2136
rect 860 2024 877 2031
rect 758 1986 805 1992
rect 758 1984 769 1986
rect 642 1938 654 1944
rect 692 1938 704 1944
rect 797 1984 805 1986
rect 955 1984 963 2039
rect 1035 2032 1044 2050
rect 1003 2026 1044 2032
rect 1003 1992 1009 2026
rect 1055 2020 1061 2067
rect 1121 2032 1127 2116
rect 1211 2117 1232 2124
rect 1282 2130 1289 2136
rect 1282 2122 1293 2130
rect 1179 2106 1186 2112
rect 1247 2106 1253 2108
rect 1179 2100 1253 2106
rect 1335 2101 1343 2116
rect 1179 2092 1186 2100
rect 1140 2084 1174 2092
rect 1140 2079 1146 2084
rect 1166 2066 1193 2073
rect 1121 2024 1183 2032
rect 1195 2028 1239 2034
rect 1047 2016 1061 2020
rect 1059 2014 1061 2016
rect 737 1938 749 1944
rect 777 1938 789 1944
rect 837 1938 849 1944
rect 931 1938 943 1944
rect 971 1938 983 1944
rect 1017 1938 1029 1952
rect 1177 2010 1215 2018
rect 1233 2014 1239 2028
rect 1247 2028 1253 2100
rect 1327 2087 1343 2101
rect 1313 2073 1327 2087
rect 1247 2022 1287 2028
rect 1307 2028 1321 2036
rect 1335 2024 1343 2087
rect 1376 2081 1384 2136
rect 1429 2116 1457 2120
rect 1469 2150 1497 2156
rect 1417 2114 1469 2116
rect 1479 2106 1485 2116
rect 1456 2099 1485 2106
rect 1177 2004 1185 2010
rect 1233 2008 1263 2014
rect 1281 2004 1287 2022
rect 1167 1990 1185 2004
rect 1213 1990 1235 2002
rect 1177 1984 1185 1990
rect 1227 1984 1239 1990
rect 1281 1964 1293 1998
rect 1376 1984 1384 2067
rect 1456 2073 1464 2099
rect 1507 2097 1523 2103
rect 1457 2024 1465 2059
rect 1517 2047 1523 2097
rect 1555 2102 1563 2116
rect 1583 2116 1611 2122
rect 1571 2113 1623 2116
rect 1655 2102 1663 2116
rect 1683 2116 1711 2122
rect 1671 2113 1723 2116
rect 1555 2095 1580 2102
rect 1655 2095 1680 2102
rect 1573 2073 1581 2095
rect 1673 2073 1681 2095
rect 1773 2093 1780 2136
rect 1835 2102 1843 2116
rect 1863 2116 1891 2122
rect 1851 2113 1903 2116
rect 1931 2148 1943 2162
rect 1991 2148 2003 2162
rect 2051 2148 2063 2162
rect 2111 2148 2123 2162
rect 2181 2156 2193 2162
rect 2243 2156 2255 2162
rect 2291 2156 2303 2162
rect 2349 2156 2361 2162
rect 2451 2156 2463 2162
rect 2497 2156 2509 2162
rect 2537 2156 2549 2162
rect 2650 2156 2662 2162
rect 1959 2116 1961 2118
rect 1959 2112 1973 2116
rect 1835 2095 1860 2102
rect 1579 2024 1587 2059
rect 1679 2024 1687 2059
rect 1773 2031 1780 2079
rect 1853 2073 1861 2095
rect 1959 2081 1965 2112
rect 2011 2106 2018 2128
rect 2079 2116 2081 2118
rect 2079 2112 2093 2116
rect 1976 2100 2018 2106
rect 1763 2024 1780 2031
rect 1859 2024 1867 2059
rect 1077 1938 1089 1944
rect 1141 1938 1153 1944
rect 1207 1938 1219 1944
rect 1253 1938 1265 1944
rect 1311 1938 1323 1944
rect 1357 1938 1369 1944
rect 1417 1938 1429 1944
rect 1487 1938 1499 1944
rect 1556 1938 1568 1944
rect 1606 1938 1618 1944
rect 1656 1938 1668 1944
rect 1706 1938 1718 1944
rect 1791 1938 1803 1944
rect 1836 1938 1848 1944
rect 1886 1938 1898 1944
rect 1959 2020 1965 2067
rect 1976 2062 1985 2100
rect 2079 2081 2085 2112
rect 2131 2106 2138 2128
rect 2096 2100 2138 2106
rect 2200 2136 2213 2142
rect 2200 2130 2207 2136
rect 2265 2124 2272 2136
rect 1976 2032 1985 2050
rect 1976 2026 2017 2032
rect 1959 2016 1973 2020
rect 1959 2014 1961 2016
rect 2011 1992 2017 2026
rect 1931 1938 1943 1944
rect 1991 1938 2003 1952
rect 2079 2020 2085 2067
rect 2096 2062 2105 2100
rect 2096 2032 2105 2050
rect 2161 2032 2167 2116
rect 2251 2117 2272 2124
rect 2322 2130 2329 2136
rect 2322 2122 2333 2130
rect 2219 2106 2226 2112
rect 2287 2106 2293 2108
rect 2219 2100 2293 2106
rect 2375 2101 2383 2116
rect 2219 2092 2226 2100
rect 2180 2084 2214 2092
rect 2180 2079 2186 2084
rect 2206 2066 2233 2073
rect 2096 2026 2137 2032
rect 2079 2016 2093 2020
rect 2079 2014 2081 2016
rect 2131 1992 2137 2026
rect 2161 2024 2223 2032
rect 2235 2028 2279 2034
rect 2051 1938 2063 1944
rect 2111 1938 2123 1952
rect 2217 2010 2255 2018
rect 2273 2014 2279 2028
rect 2287 2028 2293 2100
rect 2367 2087 2383 2101
rect 2415 2102 2423 2116
rect 2443 2116 2471 2122
rect 2431 2113 2483 2116
rect 2415 2095 2440 2102
rect 2353 2073 2367 2087
rect 2287 2022 2327 2028
rect 2347 2028 2361 2036
rect 2375 2024 2383 2087
rect 2433 2073 2441 2095
rect 2520 2093 2527 2136
rect 2439 2024 2447 2059
rect 2520 2031 2527 2079
rect 2596 2098 2614 2100
rect 2596 2089 2626 2098
rect 2697 2148 2709 2162
rect 2757 2148 2769 2162
rect 2682 2106 2689 2128
rect 2739 2116 2741 2118
rect 2727 2112 2741 2116
rect 2682 2100 2724 2106
rect 2596 2061 2604 2089
rect 2520 2024 2537 2031
rect 2217 2004 2225 2010
rect 2273 2008 2303 2014
rect 2321 2004 2327 2022
rect 2207 1990 2225 2004
rect 2253 1990 2275 2002
rect 2217 1984 2225 1990
rect 2267 1984 2279 1990
rect 2321 1964 2333 1998
rect 2181 1938 2193 1944
rect 2247 1938 2259 1944
rect 2293 1938 2305 1944
rect 2351 1938 2363 1944
rect 2416 1938 2428 1944
rect 2466 1938 2478 1944
rect 2595 1992 2602 2047
rect 2715 2062 2724 2100
rect 2735 2081 2741 2112
rect 2811 2148 2823 2162
rect 2871 2148 2883 2162
rect 2917 2156 2929 2162
rect 2997 2156 3009 2162
rect 3118 2156 3130 2162
rect 3168 2156 3180 2162
rect 2839 2116 2841 2118
rect 2839 2112 2853 2116
rect 2839 2081 2845 2112
rect 2891 2106 2898 2128
rect 2856 2100 2898 2106
rect 2715 2032 2724 2050
rect 2683 2026 2724 2032
rect 2683 1992 2689 2026
rect 2735 2020 2741 2067
rect 2727 2016 2741 2020
rect 2595 1986 2642 1992
rect 2595 1984 2603 1986
rect 2631 1984 2642 1986
rect 2739 2014 2741 2016
rect 2497 1938 2509 1944
rect 2611 1938 2623 1944
rect 2651 1938 2663 1944
rect 2697 1938 2709 1952
rect 2757 1938 2769 1944
rect 2839 2020 2845 2067
rect 2856 2062 2865 2100
rect 2856 2032 2865 2050
rect 2936 2081 2944 2136
rect 2989 2116 3017 2120
rect 3029 2150 3057 2156
rect 3114 2116 3140 2127
rect 3197 2156 3209 2162
rect 3277 2156 3289 2162
rect 3377 2156 3389 2162
rect 3417 2156 3429 2162
rect 3481 2156 3493 2162
rect 3543 2156 3555 2162
rect 3591 2156 3603 2162
rect 3649 2156 3661 2162
rect 3711 2156 3723 2162
rect 3751 2156 3763 2162
rect 3851 2156 3863 2162
rect 3931 2156 3943 2162
rect 3977 2156 3989 2162
rect 4059 2156 4071 2162
rect 4151 2156 4163 2162
rect 4191 2156 4203 2162
rect 4241 2156 4253 2162
rect 4303 2156 4315 2162
rect 4351 2156 4363 2162
rect 4409 2156 4421 2162
rect 4457 2156 4469 2162
rect 4537 2156 4549 2162
rect 4637 2156 4649 2162
rect 4677 2156 4689 2162
rect 4771 2156 4783 2162
rect 4831 2156 4843 2162
rect 4871 2156 4883 2162
rect 4917 2156 4929 2162
rect 5069 2156 5081 2162
rect 2977 2114 3029 2116
rect 2957 2097 2973 2103
rect 2957 2067 2963 2097
rect 3039 2106 3045 2116
rect 3016 2099 3045 2106
rect 2856 2026 2897 2032
rect 2839 2016 2853 2020
rect 2839 2014 2841 2016
rect 2891 1992 2897 2026
rect 2936 1984 2944 2067
rect 3016 2073 3024 2099
rect 3114 2073 3122 2116
rect 3216 2081 3224 2136
rect 3269 2116 3297 2120
rect 3309 2150 3337 2156
rect 3257 2114 3309 2116
rect 3319 2106 3325 2116
rect 3296 2099 3325 2106
rect 3017 2024 3025 2059
rect 3114 2024 3122 2059
rect 2811 1938 2823 1944
rect 2871 1938 2883 1952
rect 3143 2018 3183 2024
rect 3171 2016 3183 2018
rect 3216 1984 3224 2067
rect 3296 2073 3304 2099
rect 3400 2093 3407 2136
rect 3297 2024 3305 2059
rect 3400 2031 3407 2079
rect 3500 2136 3513 2142
rect 3500 2130 3507 2136
rect 3565 2124 3572 2136
rect 3461 2032 3467 2116
rect 3551 2117 3572 2124
rect 3622 2130 3629 2136
rect 3622 2122 3633 2130
rect 3519 2106 3526 2112
rect 3587 2106 3593 2108
rect 3519 2100 3593 2106
rect 3675 2101 3683 2116
rect 3519 2092 3526 2100
rect 3480 2084 3514 2092
rect 3480 2079 3486 2084
rect 3506 2066 3533 2073
rect 3400 2024 3417 2031
rect 2917 1938 2929 1944
rect 2977 1938 2989 1944
rect 3047 1938 3059 1944
rect 3151 1938 3163 1944
rect 3197 1938 3209 1944
rect 3257 1938 3269 1944
rect 3327 1938 3339 1944
rect 3461 2024 3523 2032
rect 3535 2028 3579 2034
rect 3517 2010 3555 2018
rect 3573 2014 3579 2028
rect 3587 2028 3593 2100
rect 3667 2087 3683 2101
rect 3653 2073 3667 2087
rect 3587 2022 3627 2028
rect 3647 2028 3661 2036
rect 3675 2024 3683 2087
rect 3517 2004 3525 2010
rect 3573 2008 3603 2014
rect 3621 2004 3627 2022
rect 3507 1990 3525 2004
rect 3553 1990 3575 2002
rect 3517 1984 3525 1990
rect 3567 1984 3579 1990
rect 3621 1964 3633 1998
rect 3697 2097 3713 2103
rect 3697 2007 3703 2097
rect 3733 2093 3740 2136
rect 3803 2150 3831 2156
rect 3843 2116 3871 2120
rect 3767 2097 3793 2103
rect 3815 2106 3821 2116
rect 3831 2114 3883 2116
rect 3815 2099 3844 2106
rect 3733 2031 3740 2079
rect 3836 2073 3844 2099
rect 3887 2097 3903 2103
rect 3723 2024 3740 2031
rect 3835 2024 3843 2059
rect 3897 2027 3903 2097
rect 3916 2081 3924 2136
rect 3969 2116 3997 2122
rect 3957 2113 4009 2116
rect 4017 2102 4025 2116
rect 4089 2108 4101 2116
rect 4000 2095 4025 2102
rect 4077 2102 4101 2108
rect 3377 1938 3389 1944
rect 3481 1938 3493 1944
rect 3547 1938 3559 1944
rect 3593 1938 3605 1944
rect 3651 1938 3663 1944
rect 3751 1938 3763 1944
rect 3916 1984 3924 2067
rect 3999 2073 4007 2095
rect 3993 2024 4001 2059
rect 3801 1938 3813 1944
rect 3871 1938 3883 1944
rect 3931 1938 3943 1944
rect 4037 2023 4043 2053
rect 4077 2053 4085 2102
rect 4173 2093 4180 2136
rect 4260 2136 4273 2142
rect 4260 2130 4267 2136
rect 4325 2124 4332 2136
rect 4037 2017 4053 2023
rect 4077 1984 4085 2039
rect 4173 2031 4180 2079
rect 4163 2024 4180 2031
rect 4221 2032 4227 2116
rect 4311 2117 4332 2124
rect 4382 2130 4389 2136
rect 4382 2122 4393 2130
rect 4279 2106 4286 2112
rect 4347 2106 4353 2108
rect 4279 2100 4353 2106
rect 4435 2101 4443 2116
rect 4279 2092 4286 2100
rect 4240 2084 4274 2092
rect 4240 2079 4246 2084
rect 4266 2066 4293 2073
rect 4221 2024 4283 2032
rect 4295 2028 4339 2034
rect 3962 1938 3974 1944
rect 4012 1938 4024 1944
rect 4277 2010 4315 2018
rect 4333 2014 4339 2028
rect 4347 2028 4353 2100
rect 4427 2087 4443 2101
rect 4413 2073 4427 2087
rect 4347 2022 4387 2028
rect 4407 2028 4421 2036
rect 4435 2024 4443 2087
rect 4476 2081 4484 2136
rect 4529 2116 4557 2120
rect 4569 2150 4597 2156
rect 4517 2114 4569 2116
rect 4579 2106 4585 2116
rect 4556 2099 4585 2106
rect 4277 2004 4285 2010
rect 4333 2008 4363 2014
rect 4381 2004 4387 2022
rect 4267 1990 4285 2004
rect 4313 1990 4335 2002
rect 4277 1984 4285 1990
rect 4327 1984 4339 1990
rect 4381 1964 4393 1998
rect 4476 1984 4484 2067
rect 4497 2047 4503 2093
rect 4556 2073 4564 2099
rect 4660 2093 4667 2136
rect 4735 2102 4743 2116
rect 4763 2116 4791 2122
rect 4751 2113 4803 2116
rect 4735 2095 4760 2102
rect 4557 2024 4565 2059
rect 4660 2031 4667 2079
rect 4753 2073 4761 2095
rect 4853 2093 4860 2136
rect 4909 2116 4937 2120
rect 4949 2150 4977 2156
rect 5111 2156 5123 2162
rect 5151 2156 5163 2162
rect 5177 2156 5185 2162
rect 5217 2156 5229 2162
rect 5351 2156 5363 2162
rect 5417 2156 5429 2162
rect 5531 2156 5543 2162
rect 5571 2156 5583 2162
rect 5671 2156 5683 2162
rect 5751 2156 5763 2162
rect 4897 2114 4949 2116
rect 4959 2106 4965 2116
rect 4936 2099 4965 2106
rect 5039 2108 5051 2116
rect 5039 2102 5063 2108
rect 4660 2024 4677 2031
rect 4759 2024 4767 2059
rect 4853 2031 4860 2079
rect 4936 2073 4944 2099
rect 4843 2024 4860 2031
rect 4937 2024 4945 2059
rect 5055 2053 5063 2102
rect 5133 2093 5140 2136
rect 5203 2108 5209 2136
rect 5303 2150 5331 2156
rect 5343 2116 5371 2120
rect 5203 2102 5213 2108
rect 4057 1938 4069 1944
rect 4097 1938 4109 1944
rect 4191 1938 4203 1944
rect 4241 1938 4253 1944
rect 4307 1938 4319 1944
rect 4353 1938 4365 1944
rect 4411 1938 4423 1944
rect 4457 1938 4469 1944
rect 4517 1938 4529 1944
rect 4587 1938 4599 1944
rect 4637 1938 4649 1944
rect 4736 1938 4748 1944
rect 4786 1938 4798 1944
rect 4871 1938 4883 1944
rect 5055 1984 5063 2039
rect 5133 2031 5140 2079
rect 5218 2041 5224 2096
rect 5240 2081 5247 2116
rect 5315 2106 5321 2116
rect 5331 2114 5383 2116
rect 5409 2116 5437 2120
rect 5449 2150 5477 2156
rect 5397 2114 5449 2116
rect 5459 2106 5465 2116
rect 5315 2099 5344 2106
rect 5123 2024 5140 2031
rect 5177 2032 5213 2040
rect 5177 2024 5185 2032
rect 4897 1938 4909 1944
rect 4967 1938 4979 1944
rect 5234 2023 5243 2067
rect 5336 2073 5344 2099
rect 5436 2099 5465 2106
rect 5436 2073 5444 2099
rect 5553 2093 5560 2136
rect 5623 2150 5651 2156
rect 5663 2116 5691 2120
rect 5779 2156 5791 2162
rect 5879 2156 5891 2162
rect 5937 2156 5949 2162
rect 5985 2156 5997 2162
rect 6047 2156 6059 2162
rect 6121 2156 6133 2162
rect 6183 2156 6195 2162
rect 6231 2156 6243 2162
rect 6289 2156 6301 2162
rect 5635 2106 5641 2116
rect 5651 2114 5703 2116
rect 5587 2097 5603 2103
rect 5635 2099 5664 2106
rect 5335 2024 5343 2059
rect 5437 2024 5445 2059
rect 5553 2031 5560 2079
rect 5597 2047 5603 2097
rect 5656 2073 5664 2099
rect 5543 2024 5560 2031
rect 5655 2024 5663 2059
rect 5717 2047 5723 2093
rect 5736 2081 5744 2136
rect 5809 2108 5821 2116
rect 5797 2102 5821 2108
rect 6027 2136 6040 2142
rect 5911 2130 5918 2136
rect 5907 2122 5918 2130
rect 5968 2124 5975 2136
rect 6033 2130 6040 2136
rect 5239 2014 5243 2023
rect 5031 1938 5043 1944
rect 5071 1938 5083 1944
rect 5151 1938 5163 1944
rect 5207 1938 5219 1944
rect 5301 1938 5313 1944
rect 5371 1938 5383 1944
rect 5397 1938 5409 1944
rect 5467 1938 5479 1944
rect 5571 1938 5583 1944
rect 5736 1984 5744 2067
rect 5797 2053 5805 2102
rect 5857 2101 5865 2116
rect 5968 2117 5989 2124
rect 5947 2106 5953 2108
rect 6014 2106 6021 2112
rect 5857 2087 5873 2101
rect 5947 2100 6021 2106
rect 5797 1984 5805 2039
rect 5857 2024 5865 2087
rect 5873 2073 5887 2087
rect 5879 2028 5893 2036
rect 5621 1938 5633 1944
rect 5691 1938 5703 1944
rect 5751 1938 5763 1944
rect 5947 2028 5953 2100
rect 6014 2092 6021 2100
rect 6026 2084 6060 2092
rect 6054 2079 6060 2084
rect 6007 2066 6034 2073
rect 5913 2022 5953 2028
rect 5961 2028 6005 2034
rect 5913 2004 5919 2022
rect 5961 2014 5967 2028
rect 6073 2032 6079 2116
rect 6017 2024 6079 2032
rect 5937 2008 5967 2014
rect 5985 2010 6023 2018
rect 6015 2004 6023 2010
rect 5907 1964 5919 1998
rect 5965 1990 5987 2002
rect 6015 1990 6033 2004
rect 5961 1984 5973 1990
rect 6015 1984 6023 1990
rect 6140 2136 6153 2142
rect 6140 2130 6147 2136
rect 6205 2124 6212 2136
rect 6101 2032 6107 2116
rect 6191 2117 6212 2124
rect 6262 2130 6269 2136
rect 6262 2122 6273 2130
rect 6159 2106 6166 2112
rect 6357 2148 6369 2162
rect 6417 2148 6429 2162
rect 6227 2106 6233 2108
rect 6159 2100 6233 2106
rect 6315 2101 6323 2116
rect 6159 2092 6166 2100
rect 6120 2084 6154 2092
rect 6120 2079 6126 2084
rect 6146 2066 6173 2073
rect 6101 2024 6163 2032
rect 6175 2028 6219 2034
rect 6157 2010 6195 2018
rect 6213 2014 6219 2028
rect 6227 2028 6233 2100
rect 6307 2087 6323 2101
rect 6342 2106 6349 2128
rect 6399 2116 6401 2118
rect 6387 2112 6401 2116
rect 6342 2100 6384 2106
rect 6293 2073 6307 2087
rect 6227 2022 6267 2028
rect 6287 2028 6301 2036
rect 6315 2024 6323 2087
rect 6375 2062 6384 2100
rect 6395 2081 6401 2112
rect 6460 2156 6472 2162
rect 6510 2156 6522 2162
rect 6577 2156 6589 2162
rect 6500 2116 6526 2127
rect 6375 2032 6384 2050
rect 6157 2004 6165 2010
rect 6213 2008 6243 2014
rect 6261 2004 6267 2022
rect 6147 1990 6165 2004
rect 6193 1990 6215 2002
rect 6157 1984 6165 1990
rect 6207 1984 6219 1990
rect 6261 1964 6273 1998
rect 6343 2026 6384 2032
rect 6343 1992 6349 2026
rect 6395 2020 6401 2067
rect 6518 2073 6526 2116
rect 6569 2116 6597 2122
rect 6557 2113 6609 2116
rect 6617 2102 6625 2116
rect 6600 2095 6625 2102
rect 6599 2073 6607 2095
rect 6518 2024 6526 2059
rect 6593 2024 6601 2059
rect 6387 2016 6401 2020
rect 6399 2014 6401 2016
rect 5777 1938 5789 1944
rect 5817 1938 5829 1944
rect 5877 1938 5889 1944
rect 5935 1938 5947 1944
rect 5981 1938 5993 1944
rect 6047 1938 6059 1944
rect 6121 1938 6133 1944
rect 6187 1938 6199 1944
rect 6233 1938 6245 1944
rect 6291 1938 6303 1944
rect 6357 1938 6369 1952
rect 6457 2018 6497 2024
rect 6457 2016 6469 2018
rect 6417 1938 6429 1944
rect 6477 1938 6489 1944
rect 6562 1938 6574 1944
rect 6612 1938 6624 1944
rect -62 1936 6736 1938
rect -62 1924 4 1936
rect -62 1922 6736 1924
rect -62 1458 -2 1922
rect 51 1916 63 1922
rect 97 1916 109 1922
rect 155 1916 167 1922
rect 201 1916 213 1922
rect 267 1916 279 1922
rect 317 1916 329 1922
rect 451 1916 463 1922
rect 511 1916 523 1922
rect 36 1793 44 1876
rect 127 1862 139 1896
rect 181 1870 193 1876
rect 235 1870 243 1876
rect 185 1858 207 1870
rect 235 1856 253 1870
rect 133 1838 139 1856
rect 157 1846 187 1852
rect 235 1850 243 1856
rect 36 1724 44 1779
rect 77 1773 85 1836
rect 99 1824 113 1832
rect 133 1832 173 1838
rect 93 1773 107 1787
rect 77 1759 93 1773
rect 167 1760 173 1832
rect 181 1832 187 1846
rect 205 1842 243 1850
rect 181 1826 225 1832
rect 237 1828 299 1836
rect 227 1787 254 1794
rect 274 1776 280 1781
rect 246 1768 280 1776
rect 234 1760 241 1768
rect 77 1744 85 1759
rect 167 1754 241 1760
rect 167 1752 173 1754
rect 234 1748 241 1754
rect 127 1730 138 1738
rect 131 1724 138 1730
rect 188 1736 209 1743
rect 293 1744 299 1828
rect 340 1829 357 1836
rect 556 1916 568 1922
rect 606 1916 618 1922
rect 657 1916 669 1922
rect 715 1916 727 1922
rect 761 1916 773 1922
rect 827 1916 839 1922
rect 911 1916 923 1922
rect 951 1916 963 1922
rect 423 1829 440 1836
rect 340 1781 347 1829
rect 188 1724 195 1736
rect 253 1724 260 1730
rect 247 1718 260 1724
rect 340 1724 347 1767
rect 433 1781 440 1829
rect 496 1793 504 1876
rect 687 1862 699 1896
rect 741 1870 753 1876
rect 795 1870 803 1876
rect 745 1858 767 1870
rect 795 1856 813 1870
rect 693 1838 699 1856
rect 717 1846 747 1852
rect 795 1850 803 1856
rect 579 1801 587 1836
rect 433 1724 440 1767
rect 496 1724 504 1779
rect 573 1765 581 1787
rect 637 1773 645 1836
rect 659 1824 673 1832
rect 693 1832 733 1838
rect 653 1773 667 1787
rect 555 1758 580 1765
rect 637 1759 653 1773
rect 727 1760 733 1832
rect 741 1832 747 1846
rect 765 1842 803 1850
rect 741 1826 785 1832
rect 797 1828 859 1836
rect 787 1787 814 1794
rect 834 1776 840 1781
rect 806 1768 840 1776
rect 794 1760 801 1768
rect 555 1744 563 1758
rect 51 1698 63 1704
rect 99 1698 111 1704
rect 157 1698 169 1704
rect 205 1698 217 1704
rect 267 1698 279 1704
rect 317 1698 329 1704
rect 357 1698 369 1704
rect 571 1744 623 1747
rect 583 1738 611 1744
rect 637 1744 645 1759
rect 727 1754 801 1760
rect 727 1752 733 1754
rect 794 1748 801 1754
rect 687 1730 698 1738
rect 691 1724 698 1730
rect 748 1736 769 1743
rect 853 1744 859 1828
rect 895 1874 903 1876
rect 977 1916 989 1922
rect 1021 1916 1033 1922
rect 1077 1916 1089 1922
rect 1142 1916 1154 1922
rect 1192 1916 1204 1922
rect 931 1874 942 1876
rect 895 1868 942 1874
rect 895 1813 902 1868
rect 896 1771 904 1799
rect 896 1762 926 1771
rect 896 1760 914 1762
rect 748 1724 755 1736
rect 813 1724 820 1730
rect 807 1718 820 1724
rect 998 1762 1006 1876
rect 1041 1801 1049 1836
rect 1047 1787 1049 1801
rect 1096 1793 1104 1876
rect 1251 1916 1263 1922
rect 1291 1916 1303 1922
rect 1351 1916 1363 1922
rect 1391 1916 1403 1922
rect 1173 1801 1181 1836
rect 977 1754 1015 1762
rect 977 1744 989 1754
rect 1041 1744 1049 1787
rect 1039 1734 1049 1744
rect 1096 1724 1104 1779
rect 1179 1765 1187 1787
rect 1237 1783 1243 1853
rect 1275 1821 1283 1876
rect 1335 1874 1343 1876
rect 1417 1916 1429 1922
rect 1501 1916 1513 1922
rect 1567 1916 1579 1922
rect 1613 1916 1625 1922
rect 1671 1916 1683 1922
rect 1717 1916 1729 1922
rect 1777 1916 1789 1922
rect 1847 1916 1859 1922
rect 1371 1874 1382 1876
rect 1335 1868 1382 1874
rect 1335 1813 1342 1868
rect 1207 1777 1243 1783
rect 1180 1758 1205 1765
rect 1275 1758 1283 1807
rect 1336 1771 1344 1799
rect 1436 1793 1444 1876
rect 1537 1870 1545 1876
rect 1587 1870 1599 1876
rect 1527 1856 1545 1870
rect 1573 1858 1595 1870
rect 1641 1862 1653 1896
rect 1537 1850 1545 1856
rect 1537 1842 1575 1850
rect 1593 1846 1623 1852
rect 1481 1828 1543 1836
rect 1336 1762 1366 1771
rect 1336 1760 1354 1762
rect 1137 1744 1189 1747
rect 1149 1738 1177 1744
rect 1197 1744 1205 1758
rect 1259 1752 1283 1758
rect 1259 1744 1271 1752
rect 1436 1724 1444 1779
rect 1481 1744 1487 1828
rect 1593 1832 1599 1846
rect 1641 1838 1647 1856
rect 1555 1826 1599 1832
rect 1607 1832 1647 1838
rect 1526 1787 1553 1794
rect 1500 1776 1506 1781
rect 1500 1768 1534 1776
rect 1539 1760 1546 1768
rect 1607 1760 1613 1832
rect 1667 1824 1681 1832
rect 1673 1773 1687 1787
rect 1695 1773 1703 1836
rect 1736 1793 1744 1876
rect 1897 1916 1909 1922
rect 1982 1916 1994 1922
rect 2032 1916 2044 1922
rect 2097 1916 2109 1922
rect 2155 1916 2167 1922
rect 2201 1916 2213 1922
rect 2267 1916 2279 1922
rect 2341 1916 2353 1922
rect 2411 1916 2423 1922
rect 2127 1862 2139 1896
rect 2181 1870 2193 1876
rect 2235 1870 2243 1876
rect 2185 1858 2207 1870
rect 2235 1856 2253 1870
rect 2133 1838 2139 1856
rect 2157 1846 2187 1852
rect 2235 1850 2243 1856
rect 1817 1801 1825 1836
rect 1920 1829 1937 1836
rect 1539 1754 1613 1760
rect 1687 1759 1703 1773
rect 1539 1748 1546 1754
rect 1607 1752 1613 1754
rect 411 1698 423 1704
rect 451 1698 463 1704
rect 511 1698 523 1704
rect 591 1698 603 1704
rect 659 1698 671 1704
rect 717 1698 729 1704
rect 765 1698 777 1704
rect 827 1698 839 1704
rect 950 1698 962 1704
rect 1007 1698 1019 1704
rect 1077 1698 1089 1704
rect 1157 1698 1169 1704
rect 1289 1698 1301 1704
rect 1390 1698 1402 1704
rect 1571 1736 1592 1743
rect 1695 1744 1703 1759
rect 1520 1724 1527 1730
rect 1585 1724 1592 1736
rect 1642 1730 1653 1738
rect 1642 1724 1649 1730
rect 1520 1718 1533 1724
rect 1736 1724 1744 1779
rect 1816 1761 1824 1787
rect 1920 1781 1927 1829
rect 2013 1801 2021 1836
rect 1816 1754 1845 1761
rect 1777 1744 1829 1746
rect 1839 1744 1845 1754
rect 1789 1740 1817 1744
rect 1829 1704 1857 1710
rect 1920 1724 1927 1767
rect 2019 1765 2027 1787
rect 2077 1773 2085 1836
rect 2099 1824 2113 1832
rect 2133 1832 2173 1838
rect 2093 1773 2107 1787
rect 2020 1758 2045 1765
rect 1977 1744 2029 1747
rect 1989 1738 2017 1744
rect 2037 1744 2045 1758
rect 2077 1759 2093 1773
rect 2167 1760 2173 1832
rect 2181 1832 2187 1846
rect 2205 1842 2243 1850
rect 2437 1916 2449 1922
rect 2497 1916 2509 1922
rect 2597 1916 2609 1922
rect 2655 1916 2667 1922
rect 2701 1916 2713 1922
rect 2767 1916 2779 1922
rect 2817 1916 2829 1922
rect 2857 1916 2869 1922
rect 2936 1916 2948 1922
rect 2986 1916 2998 1922
rect 2181 1826 2225 1832
rect 2237 1828 2299 1836
rect 2227 1787 2254 1794
rect 2274 1776 2280 1781
rect 2246 1768 2280 1776
rect 2234 1760 2241 1768
rect 2077 1744 2085 1759
rect 2167 1754 2241 1760
rect 2167 1752 2173 1754
rect 2234 1748 2241 1754
rect 2127 1730 2138 1738
rect 2131 1724 2138 1730
rect 2188 1736 2209 1743
rect 2293 1744 2299 1828
rect 2375 1801 2383 1836
rect 2376 1761 2384 1787
rect 2456 1793 2464 1876
rect 2520 1829 2537 1836
rect 2627 1862 2639 1896
rect 2681 1870 2693 1876
rect 2735 1870 2743 1876
rect 2685 1858 2707 1870
rect 2735 1856 2753 1870
rect 2633 1838 2639 1856
rect 2657 1846 2687 1852
rect 2735 1850 2743 1856
rect 2520 1781 2527 1829
rect 2355 1754 2384 1761
rect 2355 1744 2361 1754
rect 2371 1744 2423 1746
rect 2188 1724 2195 1736
rect 2253 1724 2260 1730
rect 2247 1718 2260 1724
rect 2343 1704 2371 1710
rect 2383 1740 2411 1744
rect 2456 1724 2464 1779
rect 2520 1724 2527 1767
rect 2577 1773 2585 1836
rect 2599 1824 2613 1832
rect 2633 1832 2673 1838
rect 2593 1773 2607 1787
rect 2577 1759 2593 1773
rect 2667 1760 2673 1832
rect 2681 1832 2687 1846
rect 2705 1842 2743 1850
rect 2838 1874 2849 1876
rect 2877 1874 2885 1876
rect 2838 1868 2885 1874
rect 2681 1826 2725 1832
rect 2737 1828 2799 1836
rect 2727 1787 2754 1794
rect 2774 1776 2780 1781
rect 2746 1768 2780 1776
rect 2734 1760 2741 1768
rect 2577 1744 2585 1759
rect 2667 1754 2741 1760
rect 2667 1752 2673 1754
rect 2734 1748 2741 1754
rect 2627 1730 2638 1738
rect 2631 1724 2638 1730
rect 2688 1736 2709 1743
rect 2793 1744 2799 1828
rect 2878 1813 2885 1868
rect 3017 1916 3029 1922
rect 3151 1916 3163 1922
rect 3251 1916 3263 1922
rect 3329 1916 3341 1922
rect 3391 1916 3403 1922
rect 3431 1916 3443 1922
rect 3171 1842 3183 1844
rect 3143 1836 3183 1842
rect 3271 1842 3283 1844
rect 3243 1836 3283 1842
rect 3457 1916 3469 1922
rect 3537 1916 3549 1922
rect 3577 1916 3589 1922
rect 2959 1801 2967 1836
rect 3040 1829 3057 1836
rect 2876 1771 2884 1799
rect 2688 1724 2695 1736
rect 2753 1724 2760 1730
rect 2747 1718 2760 1724
rect 2854 1762 2884 1771
rect 2953 1765 2961 1787
rect 3040 1781 3047 1829
rect 3114 1801 3122 1836
rect 3214 1801 3222 1836
rect 3311 1801 3319 1836
rect 3355 1830 3363 1876
rect 3337 1824 3363 1830
rect 3337 1818 3340 1824
rect 2866 1760 2884 1762
rect 2935 1758 2960 1765
rect 2935 1744 2943 1758
rect 2951 1744 3003 1747
rect 2963 1738 2991 1744
rect 3040 1724 3047 1767
rect 3114 1744 3122 1787
rect 3214 1744 3222 1787
rect 3311 1787 3313 1801
rect 3311 1744 3319 1787
rect 3333 1762 3340 1818
rect 3377 1767 3383 1833
rect 3415 1821 3423 1876
rect 3622 1916 3634 1922
rect 3672 1916 3684 1922
rect 3480 1829 3497 1836
rect 3337 1756 3340 1762
rect 3337 1750 3359 1756
rect 3415 1758 3423 1807
rect 3480 1781 3487 1829
rect 3557 1821 3565 1876
rect 3731 1916 3743 1922
rect 3771 1916 3783 1922
rect 3831 1916 3843 1922
rect 3857 1916 3869 1922
rect 3897 1916 3909 1922
rect 3937 1916 3949 1922
rect 4017 1916 4029 1922
rect 4087 1916 4099 1922
rect 4191 1916 4203 1922
rect 3114 1733 3140 1744
rect 1417 1698 1429 1704
rect 1501 1698 1513 1704
rect 1563 1698 1575 1704
rect 1611 1698 1623 1704
rect 1669 1698 1681 1704
rect 1717 1698 1729 1704
rect 1797 1698 1809 1704
rect 1897 1698 1909 1704
rect 1937 1698 1949 1704
rect 1997 1698 2009 1704
rect 2099 1698 2111 1704
rect 2157 1698 2169 1704
rect 2205 1698 2217 1704
rect 2267 1698 2279 1704
rect 2391 1698 2403 1704
rect 2437 1698 2449 1704
rect 2497 1698 2509 1704
rect 2537 1698 2549 1704
rect 2599 1698 2611 1704
rect 2657 1698 2669 1704
rect 2705 1698 2717 1704
rect 2767 1698 2779 1704
rect 2818 1698 2830 1704
rect 2971 1698 2983 1704
rect 3017 1698 3029 1704
rect 3057 1698 3069 1704
rect 3214 1733 3240 1744
rect 3118 1698 3130 1704
rect 3168 1698 3180 1704
rect 3351 1724 3359 1750
rect 3399 1752 3423 1758
rect 3399 1744 3411 1752
rect 3480 1724 3487 1767
rect 3557 1758 3565 1807
rect 3653 1801 3661 1836
rect 3755 1821 3763 1876
rect 3659 1765 3667 1787
rect 3717 1783 3723 1813
rect 3687 1777 3723 1783
rect 3660 1758 3685 1765
rect 3755 1758 3763 1807
rect 3816 1793 3824 1876
rect 3877 1821 3885 1876
rect 4222 1916 4234 1922
rect 4272 1916 4284 1922
rect 4317 1914 4329 1922
rect 4357 1916 4369 1922
rect 4287 1857 4303 1863
rect 3960 1829 3977 1836
rect 3557 1752 3581 1758
rect 3569 1744 3581 1752
rect 3218 1698 3230 1704
rect 3268 1698 3280 1704
rect 3329 1698 3341 1704
rect 3429 1698 3441 1704
rect 3457 1698 3469 1704
rect 3497 1698 3509 1704
rect 3617 1744 3669 1747
rect 3629 1738 3657 1744
rect 3677 1744 3685 1758
rect 3739 1752 3763 1758
rect 3739 1744 3751 1752
rect 3816 1724 3824 1779
rect 3877 1758 3885 1807
rect 3960 1781 3967 1829
rect 4057 1801 4065 1836
rect 4163 1829 4180 1836
rect 3877 1752 3901 1758
rect 3889 1744 3901 1752
rect 3539 1698 3551 1704
rect 3637 1698 3649 1704
rect 3769 1698 3781 1704
rect 3831 1698 3843 1704
rect 3960 1724 3967 1767
rect 4056 1761 4064 1787
rect 4173 1781 4180 1829
rect 4253 1801 4261 1836
rect 4297 1807 4303 1857
rect 4402 1916 4414 1922
rect 4452 1916 4464 1922
rect 4551 1916 4563 1922
rect 4487 1877 4503 1883
rect 4467 1857 4483 1863
rect 4339 1793 4348 1836
rect 4056 1754 4085 1761
rect 4017 1744 4069 1746
rect 4079 1744 4085 1754
rect 4029 1740 4057 1744
rect 4069 1704 4097 1710
rect 4173 1724 4180 1767
rect 4259 1765 4267 1787
rect 4339 1779 4353 1793
rect 4260 1758 4285 1765
rect 4217 1744 4269 1747
rect 4229 1738 4257 1744
rect 4277 1744 4285 1758
rect 4339 1744 4348 1779
rect 4377 1763 4383 1813
rect 4433 1801 4441 1836
rect 4377 1757 4393 1763
rect 4439 1765 4447 1787
rect 4477 1767 4483 1857
rect 4440 1758 4465 1765
rect 4397 1744 4449 1747
rect 4409 1738 4437 1744
rect 4457 1744 4465 1758
rect 4497 1763 4503 1877
rect 4601 1916 4613 1922
rect 4671 1916 4683 1922
rect 4731 1916 4743 1922
rect 4777 1916 4789 1922
rect 4835 1916 4847 1922
rect 4881 1916 4893 1922
rect 4947 1916 4959 1922
rect 5017 1916 5029 1922
rect 5097 1916 5109 1922
rect 5182 1916 5194 1922
rect 5232 1916 5244 1922
rect 4523 1829 4540 1836
rect 4533 1781 4540 1829
rect 4635 1801 4643 1836
rect 4497 1757 4513 1763
rect 4533 1724 4540 1767
rect 4636 1761 4644 1787
rect 4716 1793 4724 1876
rect 4807 1862 4819 1896
rect 4861 1870 4873 1876
rect 4915 1870 4923 1876
rect 4865 1858 4887 1870
rect 4915 1856 4933 1870
rect 4813 1838 4819 1856
rect 4837 1846 4867 1852
rect 4915 1850 4923 1856
rect 4615 1754 4644 1761
rect 4615 1744 4621 1754
rect 4631 1744 4683 1746
rect 4603 1704 4631 1710
rect 4643 1740 4671 1744
rect 4716 1724 4724 1779
rect 4757 1773 4765 1836
rect 4779 1824 4793 1832
rect 4813 1832 4853 1838
rect 4773 1773 4787 1787
rect 4757 1759 4773 1773
rect 4847 1760 4853 1832
rect 4861 1832 4867 1846
rect 4885 1842 4923 1850
rect 4997 1842 5009 1844
rect 4997 1836 5037 1842
rect 5277 1916 5289 1922
rect 5317 1916 5329 1922
rect 5399 1916 5411 1922
rect 5491 1916 5503 1922
rect 5551 1916 5563 1922
rect 5298 1874 5309 1876
rect 5337 1874 5345 1876
rect 5298 1868 5345 1874
rect 4861 1826 4905 1832
rect 4917 1828 4979 1836
rect 4907 1787 4934 1794
rect 4954 1776 4960 1781
rect 4926 1768 4960 1776
rect 4914 1760 4921 1768
rect 4757 1744 4765 1759
rect 4847 1754 4921 1760
rect 4847 1752 4853 1754
rect 4914 1748 4921 1754
rect 4807 1730 4818 1738
rect 4811 1724 4818 1730
rect 4868 1736 4889 1743
rect 4973 1744 4979 1828
rect 5058 1801 5066 1836
rect 5120 1829 5137 1836
rect 5058 1744 5066 1787
rect 5120 1781 5127 1829
rect 5213 1801 5221 1836
rect 5338 1813 5345 1868
rect 5377 1830 5385 1876
rect 5377 1824 5403 1830
rect 5400 1818 5403 1824
rect 4868 1724 4875 1736
rect 4933 1724 4940 1730
rect 4927 1718 4940 1724
rect 5040 1733 5066 1744
rect 5120 1724 5127 1767
rect 5219 1765 5227 1787
rect 5336 1771 5344 1799
rect 5220 1758 5245 1765
rect 5177 1744 5229 1747
rect 3859 1698 3871 1704
rect 3937 1698 3949 1704
rect 3977 1698 3989 1704
rect 4037 1698 4049 1704
rect 4151 1698 4163 1704
rect 4191 1698 4203 1704
rect 4237 1698 4249 1704
rect 4317 1698 4329 1704
rect 4357 1698 4369 1704
rect 4417 1698 4429 1704
rect 4511 1698 4523 1704
rect 4551 1698 4563 1704
rect 4651 1698 4663 1704
rect 4731 1698 4743 1704
rect 4779 1698 4791 1704
rect 4837 1698 4849 1704
rect 4885 1698 4897 1704
rect 4947 1698 4959 1704
rect 5000 1698 5012 1704
rect 5050 1698 5062 1704
rect 5189 1738 5217 1744
rect 5237 1744 5245 1758
rect 5314 1762 5344 1771
rect 5326 1760 5344 1762
rect 5400 1762 5407 1818
rect 5421 1801 5429 1836
rect 5427 1787 5429 1801
rect 5476 1793 5484 1876
rect 5596 1916 5608 1922
rect 5646 1916 5658 1922
rect 5677 1916 5689 1922
rect 5717 1916 5729 1922
rect 5831 1916 5843 1922
rect 5899 1916 5911 1922
rect 5976 1916 5988 1922
rect 6026 1916 6038 1922
rect 5536 1801 5544 1836
rect 5619 1801 5627 1836
rect 5697 1821 5705 1876
rect 5783 1910 5811 1916
rect 5823 1838 5851 1844
rect 5792 1830 5804 1836
rect 5877 1830 5885 1876
rect 6081 1916 6093 1922
rect 6151 1916 6163 1922
rect 6197 1908 6209 1922
rect 6257 1916 6269 1922
rect 5400 1756 5403 1762
rect 5381 1750 5403 1756
rect 5381 1724 5389 1750
rect 5421 1744 5429 1787
rect 5476 1724 5484 1779
rect 5536 1744 5544 1787
rect 5613 1765 5621 1787
rect 5792 1824 5819 1830
rect 5877 1824 5903 1830
rect 5747 1817 5763 1823
rect 5595 1758 5620 1765
rect 5697 1758 5705 1807
rect 5757 1763 5763 1817
rect 5813 1801 5819 1824
rect 5900 1818 5903 1824
rect 5595 1744 5603 1758
rect 5697 1752 5721 1758
rect 5757 1757 5773 1763
rect 5611 1744 5663 1747
rect 5709 1744 5721 1752
rect 5820 1744 5827 1787
rect 5900 1762 5907 1818
rect 5921 1801 5929 1836
rect 5999 1801 6007 1836
rect 6115 1801 6123 1836
rect 6183 1834 6189 1868
rect 6239 1844 6241 1846
rect 6227 1840 6241 1844
rect 6183 1828 6224 1834
rect 5927 1787 5929 1801
rect 5900 1756 5903 1762
rect 5881 1750 5903 1756
rect 5623 1738 5651 1744
rect 5881 1724 5889 1750
rect 5921 1744 5929 1787
rect 5993 1765 6001 1787
rect 5975 1758 6000 1765
rect 6116 1761 6124 1787
rect 6215 1810 6224 1828
rect 5975 1744 5983 1758
rect 6095 1754 6124 1761
rect 6215 1760 6224 1798
rect 6235 1793 6241 1840
rect 6317 1908 6329 1922
rect 6377 1916 6389 1922
rect 6303 1834 6309 1868
rect 6359 1844 6361 1846
rect 6347 1840 6361 1844
rect 6303 1828 6344 1834
rect 6335 1810 6344 1828
rect 6182 1754 6224 1760
rect 5991 1744 6043 1747
rect 6095 1744 6101 1754
rect 6111 1744 6163 1746
rect 6003 1738 6031 1744
rect 6083 1704 6111 1710
rect 6123 1740 6151 1744
rect 6182 1732 6189 1754
rect 6235 1748 6241 1779
rect 6335 1760 6344 1798
rect 6355 1793 6361 1840
rect 6417 1916 6429 1922
rect 6482 1916 6494 1922
rect 6532 1916 6544 1922
rect 6436 1793 6444 1876
rect 6591 1916 6603 1922
rect 6631 1916 6643 1922
rect 6513 1801 6521 1836
rect 6615 1821 6623 1876
rect 6302 1754 6344 1760
rect 6227 1744 6241 1748
rect 6239 1742 6241 1744
rect 6302 1732 6309 1754
rect 6355 1748 6361 1779
rect 6347 1744 6361 1748
rect 6359 1742 6361 1744
rect 6436 1724 6444 1779
rect 6519 1765 6527 1787
rect 6520 1758 6545 1765
rect 6615 1758 6623 1807
rect 6477 1744 6529 1747
rect 5097 1698 5109 1704
rect 5137 1698 5149 1704
rect 5197 1698 5209 1704
rect 5278 1698 5290 1704
rect 5399 1698 5411 1704
rect 5491 1698 5503 1704
rect 5551 1698 5563 1704
rect 5631 1698 5643 1704
rect 5679 1698 5691 1704
rect 5792 1698 5804 1704
rect 5848 1698 5860 1704
rect 5899 1698 5911 1704
rect 6011 1698 6023 1704
rect 6131 1698 6143 1704
rect 6197 1698 6209 1712
rect 6257 1698 6269 1712
rect 6317 1698 6329 1712
rect 6377 1698 6389 1712
rect 6489 1738 6517 1744
rect 6537 1744 6545 1758
rect 6599 1752 6623 1758
rect 6599 1744 6611 1752
rect 6417 1698 6429 1704
rect 6497 1698 6509 1704
rect 6629 1698 6641 1704
rect 6742 1698 6802 2162
rect 4 1696 6802 1698
rect 6736 1684 6802 1696
rect 4 1682 6802 1684
rect 31 1676 43 1682
rect 71 1676 83 1682
rect 111 1676 123 1682
rect 151 1676 163 1682
rect 191 1676 203 1682
rect 231 1676 243 1682
rect 271 1676 283 1682
rect 321 1676 333 1682
rect 383 1676 395 1682
rect 431 1676 443 1682
rect 489 1676 501 1682
rect 571 1676 583 1682
rect 53 1613 60 1656
rect 340 1656 353 1662
rect 340 1650 347 1656
rect 405 1644 412 1656
rect 132 1630 144 1636
rect 172 1630 184 1636
rect 211 1630 223 1636
rect 252 1630 264 1636
rect 126 1629 144 1630
rect 125 1622 144 1629
rect 158 1622 184 1630
rect 198 1622 223 1630
rect 237 1622 264 1630
rect 125 1601 132 1622
rect 158 1616 166 1622
rect 198 1616 206 1622
rect 237 1616 245 1622
rect 150 1604 166 1616
rect 190 1604 206 1616
rect 230 1604 245 1616
rect 53 1551 60 1599
rect 127 1587 132 1601
rect 43 1544 60 1551
rect 125 1558 132 1587
rect 158 1558 166 1604
rect 198 1558 206 1604
rect 237 1558 245 1604
rect 125 1550 143 1558
rect 158 1550 183 1558
rect 198 1550 223 1558
rect 237 1550 263 1558
rect 131 1544 143 1550
rect 171 1544 183 1550
rect 211 1544 223 1550
rect 251 1544 263 1550
rect 301 1552 307 1636
rect 391 1637 412 1644
rect 462 1650 469 1656
rect 462 1642 473 1650
rect 359 1626 366 1632
rect 598 1676 610 1682
rect 700 1676 712 1682
rect 750 1676 762 1682
rect 821 1676 833 1682
rect 883 1676 895 1682
rect 931 1676 943 1682
rect 989 1676 1001 1682
rect 1071 1676 1083 1682
rect 1117 1676 1129 1682
rect 1271 1676 1283 1682
rect 1331 1676 1343 1682
rect 1371 1676 1383 1682
rect 427 1626 433 1628
rect 359 1620 433 1626
rect 515 1621 523 1636
rect 359 1612 366 1620
rect 320 1604 354 1612
rect 320 1599 326 1604
rect 346 1586 373 1593
rect 301 1544 363 1552
rect 375 1548 419 1554
rect 71 1458 83 1464
rect 357 1530 395 1538
rect 413 1534 419 1548
rect 427 1548 433 1620
rect 507 1607 523 1621
rect 493 1593 507 1607
rect 427 1542 467 1548
rect 487 1548 501 1556
rect 515 1544 523 1607
rect 556 1601 564 1656
rect 740 1636 766 1647
rect 646 1618 664 1620
rect 634 1609 664 1618
rect 357 1524 365 1530
rect 413 1528 443 1534
rect 461 1524 467 1542
rect 347 1510 365 1524
rect 393 1510 415 1522
rect 357 1504 365 1510
rect 407 1504 419 1510
rect 461 1484 473 1518
rect 556 1504 564 1587
rect 656 1581 664 1609
rect 758 1593 766 1636
rect 840 1656 853 1662
rect 840 1650 847 1656
rect 905 1644 912 1656
rect 658 1512 665 1567
rect 758 1544 766 1579
rect 801 1552 807 1636
rect 891 1637 912 1644
rect 962 1650 969 1656
rect 962 1642 973 1650
rect 859 1626 866 1632
rect 927 1626 933 1628
rect 859 1620 933 1626
rect 1015 1621 1023 1636
rect 859 1612 866 1620
rect 820 1604 854 1612
rect 820 1599 826 1604
rect 846 1586 873 1593
rect 801 1544 863 1552
rect 875 1548 919 1554
rect 618 1506 665 1512
rect 618 1504 629 1506
rect 111 1458 123 1464
rect 151 1458 163 1464
rect 191 1458 203 1464
rect 231 1458 243 1464
rect 271 1458 283 1464
rect 321 1458 333 1464
rect 387 1458 399 1464
rect 433 1458 445 1464
rect 491 1458 503 1464
rect 571 1458 583 1464
rect 657 1504 665 1506
rect 697 1538 737 1544
rect 697 1536 709 1538
rect 857 1530 895 1538
rect 913 1534 919 1548
rect 927 1548 933 1620
rect 1007 1607 1023 1621
rect 993 1593 1007 1607
rect 927 1542 967 1548
rect 987 1548 1001 1556
rect 1015 1544 1023 1607
rect 1056 1601 1064 1656
rect 1109 1636 1137 1640
rect 1149 1670 1177 1676
rect 1097 1634 1149 1636
rect 1159 1626 1165 1636
rect 1136 1619 1165 1626
rect 1235 1622 1243 1636
rect 1263 1636 1291 1642
rect 1411 1668 1423 1682
rect 1471 1668 1483 1682
rect 1531 1668 1543 1682
rect 1591 1668 1603 1682
rect 1651 1668 1663 1682
rect 1711 1668 1723 1682
rect 1779 1676 1791 1682
rect 1837 1676 1849 1682
rect 1885 1676 1897 1682
rect 1947 1676 1959 1682
rect 1251 1633 1303 1636
rect 857 1524 865 1530
rect 913 1528 943 1534
rect 961 1524 967 1542
rect 847 1510 865 1524
rect 893 1510 915 1522
rect 857 1504 865 1510
rect 907 1504 919 1510
rect 961 1484 973 1518
rect 1056 1504 1064 1587
rect 1136 1593 1144 1619
rect 1235 1615 1260 1622
rect 1253 1593 1261 1615
rect 1353 1613 1360 1656
rect 1439 1636 1441 1638
rect 1439 1632 1453 1636
rect 1439 1601 1445 1632
rect 1491 1626 1498 1648
rect 1559 1636 1561 1638
rect 1559 1632 1573 1636
rect 1456 1620 1498 1626
rect 1137 1544 1145 1579
rect 1259 1544 1267 1579
rect 1353 1551 1360 1599
rect 1343 1544 1360 1551
rect 597 1458 609 1464
rect 637 1458 649 1464
rect 717 1458 729 1464
rect 821 1458 833 1464
rect 887 1458 899 1464
rect 933 1458 945 1464
rect 991 1458 1003 1464
rect 1071 1458 1083 1464
rect 1097 1458 1109 1464
rect 1167 1458 1179 1464
rect 1236 1458 1248 1464
rect 1286 1458 1298 1464
rect 1371 1458 1383 1464
rect 1439 1540 1445 1587
rect 1456 1582 1465 1620
rect 1559 1601 1565 1632
rect 1611 1626 1618 1648
rect 1679 1636 1681 1638
rect 1679 1632 1693 1636
rect 1576 1620 1618 1626
rect 1456 1552 1465 1570
rect 1456 1546 1497 1552
rect 1439 1536 1453 1540
rect 1439 1534 1441 1536
rect 1491 1512 1497 1546
rect 1411 1458 1423 1464
rect 1471 1458 1483 1472
rect 1559 1540 1565 1587
rect 1576 1582 1585 1620
rect 1679 1601 1685 1632
rect 1731 1626 1738 1648
rect 1696 1620 1738 1626
rect 1927 1656 1940 1662
rect 1811 1650 1818 1656
rect 1807 1642 1818 1650
rect 1868 1644 1875 1656
rect 1933 1650 1940 1656
rect 1757 1621 1765 1636
rect 1868 1637 1889 1644
rect 2017 1668 2029 1682
rect 2077 1668 2089 1682
rect 1847 1626 1853 1628
rect 1914 1626 1921 1632
rect 1576 1552 1585 1570
rect 1576 1546 1617 1552
rect 1559 1536 1573 1540
rect 1559 1534 1561 1536
rect 1611 1512 1617 1546
rect 1531 1458 1543 1464
rect 1591 1458 1603 1472
rect 1679 1540 1685 1587
rect 1696 1582 1705 1620
rect 1757 1607 1773 1621
rect 1847 1620 1921 1626
rect 1696 1552 1705 1570
rect 1696 1546 1737 1552
rect 1679 1536 1693 1540
rect 1679 1534 1681 1536
rect 1731 1512 1737 1546
rect 1757 1544 1765 1607
rect 1773 1593 1787 1607
rect 1779 1548 1793 1556
rect 1651 1458 1663 1464
rect 1711 1458 1723 1472
rect 1847 1548 1853 1620
rect 1914 1612 1921 1620
rect 1926 1604 1960 1612
rect 1954 1599 1960 1604
rect 1907 1586 1934 1593
rect 1813 1542 1853 1548
rect 1861 1548 1905 1554
rect 1813 1524 1819 1542
rect 1861 1534 1867 1548
rect 1973 1552 1979 1636
rect 2002 1626 2009 1648
rect 2059 1636 2061 1638
rect 2047 1632 2061 1636
rect 2002 1620 2044 1626
rect 2035 1582 2044 1620
rect 2055 1601 2061 1632
rect 2117 1676 2129 1682
rect 2197 1676 2209 1682
rect 2297 1676 2309 1682
rect 2337 1676 2349 1682
rect 2431 1676 2443 1682
rect 2509 1676 2521 1682
rect 2557 1676 2569 1682
rect 2597 1676 2609 1682
rect 2689 1676 2701 1682
rect 2136 1601 2144 1656
rect 2189 1636 2217 1640
rect 2229 1670 2257 1676
rect 2177 1634 2229 1636
rect 2239 1626 2245 1636
rect 2216 1619 2245 1626
rect 2035 1552 2044 1570
rect 1917 1544 1979 1552
rect 1837 1528 1867 1534
rect 1885 1530 1923 1538
rect 1915 1524 1923 1530
rect 1807 1484 1819 1518
rect 1865 1510 1887 1522
rect 1915 1510 1933 1524
rect 1861 1504 1873 1510
rect 1915 1504 1923 1510
rect 2003 1546 2044 1552
rect 2003 1512 2009 1546
rect 2055 1540 2061 1587
rect 2047 1536 2061 1540
rect 2059 1534 2061 1536
rect 1777 1458 1789 1464
rect 1835 1458 1847 1464
rect 1881 1458 1893 1464
rect 1947 1458 1959 1464
rect 2017 1458 2029 1472
rect 2136 1504 2144 1587
rect 2216 1593 2224 1619
rect 2267 1617 2293 1623
rect 2320 1613 2327 1656
rect 2395 1622 2403 1636
rect 2423 1636 2451 1642
rect 2411 1633 2463 1636
rect 2395 1615 2420 1622
rect 2217 1544 2225 1579
rect 2320 1551 2327 1599
rect 2413 1593 2421 1615
rect 2491 1593 2499 1636
rect 2531 1630 2539 1656
rect 2517 1624 2539 1630
rect 2517 1618 2520 1624
rect 2491 1579 2493 1593
rect 2320 1544 2337 1551
rect 2419 1544 2427 1579
rect 2491 1544 2499 1579
rect 2513 1562 2520 1618
rect 2580 1613 2587 1656
rect 2719 1676 2731 1682
rect 2659 1628 2671 1636
rect 2749 1628 2761 1636
rect 2811 1668 2823 1682
rect 2871 1668 2883 1682
rect 2990 1676 3002 1682
rect 3051 1676 3063 1682
rect 3101 1676 3113 1682
rect 3163 1676 3175 1682
rect 3211 1676 3223 1682
rect 3269 1676 3281 1682
rect 3369 1676 3381 1682
rect 3451 1676 3463 1682
rect 3500 1676 3512 1682
rect 3556 1676 3568 1682
rect 3671 1676 3683 1682
rect 3751 1676 3763 1682
rect 2839 1636 2841 1638
rect 2839 1632 2853 1636
rect 2659 1622 2683 1628
rect 2517 1556 2520 1562
rect 2517 1550 2543 1556
rect 2077 1458 2089 1464
rect 2117 1458 2129 1464
rect 2177 1458 2189 1464
rect 2247 1458 2259 1464
rect 2535 1504 2543 1550
rect 2580 1551 2587 1599
rect 2675 1573 2683 1622
rect 2737 1622 2761 1628
rect 2737 1573 2745 1622
rect 2839 1601 2845 1632
rect 2891 1626 2898 1648
rect 2856 1620 2898 1626
rect 2580 1544 2597 1551
rect 2675 1504 2683 1559
rect 2737 1504 2745 1559
rect 2297 1458 2309 1464
rect 2396 1458 2408 1464
rect 2446 1458 2458 1464
rect 2509 1458 2521 1464
rect 2557 1458 2569 1464
rect 2651 1458 2663 1464
rect 2691 1458 2703 1464
rect 2717 1458 2729 1464
rect 2757 1458 2769 1464
rect 2839 1540 2845 1587
rect 2856 1582 2865 1620
rect 2936 1618 2954 1620
rect 2936 1609 2966 1618
rect 3120 1656 3133 1662
rect 3120 1650 3127 1656
rect 3185 1644 3192 1656
rect 2856 1552 2865 1570
rect 2936 1581 2944 1609
rect 3036 1593 3044 1636
rect 2856 1546 2897 1552
rect 2839 1536 2853 1540
rect 2839 1534 2841 1536
rect 2891 1512 2897 1546
rect 2935 1512 2942 1567
rect 3036 1544 3044 1579
rect 3081 1552 3087 1636
rect 3171 1637 3192 1644
rect 3242 1650 3249 1656
rect 3242 1642 3253 1650
rect 3139 1626 3146 1632
rect 3207 1626 3213 1628
rect 3139 1620 3213 1626
rect 3295 1621 3303 1636
rect 3339 1628 3351 1636
rect 3339 1622 3363 1628
rect 3139 1612 3146 1620
rect 3100 1604 3134 1612
rect 3100 1599 3106 1604
rect 3126 1586 3153 1593
rect 3081 1544 3143 1552
rect 3155 1548 3199 1554
rect 2935 1506 2982 1512
rect 2935 1504 2943 1506
rect 2811 1458 2823 1464
rect 2871 1458 2883 1472
rect 2971 1504 2982 1506
rect 3137 1530 3175 1538
rect 3193 1534 3199 1548
rect 3207 1548 3213 1620
rect 3287 1607 3303 1621
rect 3273 1593 3287 1607
rect 3207 1542 3247 1548
rect 3267 1548 3281 1556
rect 3295 1544 3303 1607
rect 3355 1573 3363 1622
rect 3415 1622 3423 1636
rect 3443 1636 3471 1642
rect 3431 1633 3483 1636
rect 3415 1615 3440 1622
rect 3397 1597 3413 1603
rect 3137 1524 3145 1530
rect 3193 1528 3223 1534
rect 3241 1524 3247 1542
rect 3127 1510 3145 1524
rect 3173 1510 3195 1522
rect 3137 1504 3145 1510
rect 3187 1504 3199 1510
rect 3241 1484 3253 1518
rect 3355 1504 3363 1559
rect 3397 1543 3403 1597
rect 3433 1593 3441 1615
rect 3533 1593 3540 1636
rect 3587 1617 3603 1623
rect 3439 1544 3447 1579
rect 3541 1556 3547 1579
rect 3597 1567 3603 1617
rect 3635 1622 3643 1636
rect 3663 1636 3691 1642
rect 3791 1676 3803 1682
rect 3831 1676 3843 1682
rect 3931 1676 3943 1682
rect 4011 1676 4023 1682
rect 4061 1676 4073 1682
rect 4123 1676 4135 1682
rect 4171 1676 4183 1682
rect 4229 1676 4241 1682
rect 3651 1633 3703 1636
rect 3635 1615 3660 1622
rect 3653 1593 3661 1615
rect 3736 1601 3744 1656
rect 3777 1617 3793 1623
rect 3541 1550 3568 1556
rect 3556 1544 3568 1550
rect 3659 1544 3667 1579
rect 3377 1537 3403 1543
rect 3377 1527 3383 1537
rect 2951 1458 2963 1464
rect 2991 1458 3003 1464
rect 3051 1458 3063 1464
rect 3101 1458 3113 1464
rect 3167 1458 3179 1464
rect 3213 1458 3225 1464
rect 3271 1458 3283 1464
rect 3331 1458 3343 1464
rect 3371 1458 3383 1464
rect 3509 1536 3537 1542
rect 3549 1464 3577 1470
rect 3736 1504 3744 1587
rect 3777 1563 3783 1617
rect 3813 1613 3820 1656
rect 3883 1670 3911 1676
rect 3923 1636 3951 1640
rect 3895 1626 3901 1636
rect 3911 1634 3963 1636
rect 3895 1619 3924 1626
rect 3767 1557 3783 1563
rect 3813 1551 3820 1599
rect 3916 1593 3924 1619
rect 3996 1601 4004 1656
rect 4080 1656 4093 1662
rect 4080 1650 4087 1656
rect 4145 1644 4152 1656
rect 3803 1544 3820 1551
rect 3915 1544 3923 1579
rect 3416 1458 3428 1464
rect 3466 1458 3478 1464
rect 3517 1458 3529 1464
rect 3636 1458 3648 1464
rect 3686 1458 3698 1464
rect 3751 1458 3763 1464
rect 3831 1458 3843 1464
rect 3996 1504 4004 1587
rect 4041 1552 4047 1636
rect 4131 1637 4152 1644
rect 4202 1650 4209 1656
rect 4202 1642 4213 1650
rect 4099 1626 4106 1632
rect 4167 1626 4173 1628
rect 4099 1620 4173 1626
rect 4255 1621 4263 1636
rect 4291 1668 4303 1682
rect 4351 1668 4363 1682
rect 4411 1668 4423 1682
rect 4471 1668 4483 1682
rect 4537 1668 4549 1682
rect 4597 1668 4609 1682
rect 4657 1668 4669 1682
rect 4717 1668 4729 1682
rect 4777 1668 4789 1682
rect 4837 1668 4849 1682
rect 4897 1668 4909 1682
rect 4957 1668 4969 1682
rect 5019 1676 5031 1682
rect 5077 1676 5089 1682
rect 5125 1676 5137 1682
rect 5187 1676 5199 1682
rect 5259 1676 5271 1682
rect 5317 1676 5329 1682
rect 5365 1676 5377 1682
rect 5427 1676 5439 1682
rect 5480 1676 5492 1682
rect 5536 1676 5548 1682
rect 4319 1636 4321 1638
rect 4319 1632 4333 1636
rect 4099 1612 4106 1620
rect 4060 1604 4094 1612
rect 4060 1599 4066 1604
rect 4086 1586 4113 1593
rect 4041 1544 4103 1552
rect 4115 1548 4159 1554
rect 4097 1530 4135 1538
rect 4153 1534 4159 1548
rect 4167 1548 4173 1620
rect 4247 1607 4263 1621
rect 4233 1593 4247 1607
rect 4167 1542 4207 1548
rect 4227 1548 4241 1556
rect 4255 1544 4263 1607
rect 4319 1601 4325 1632
rect 4371 1626 4378 1648
rect 4439 1636 4441 1638
rect 4439 1632 4453 1636
rect 4336 1620 4378 1626
rect 4097 1524 4105 1530
rect 4153 1528 4183 1534
rect 4201 1524 4207 1542
rect 4087 1510 4105 1524
rect 4133 1510 4155 1522
rect 4097 1504 4105 1510
rect 4147 1504 4159 1510
rect 4201 1484 4213 1518
rect 4319 1540 4325 1587
rect 4336 1582 4345 1620
rect 4439 1601 4445 1632
rect 4491 1626 4498 1648
rect 4456 1620 4498 1626
rect 4522 1626 4529 1648
rect 4579 1636 4581 1638
rect 4567 1632 4581 1636
rect 4522 1620 4564 1626
rect 4336 1552 4345 1570
rect 4336 1546 4377 1552
rect 4319 1536 4333 1540
rect 4319 1534 4321 1536
rect 4371 1512 4377 1546
rect 3881 1458 3893 1464
rect 3951 1458 3963 1464
rect 4011 1458 4023 1464
rect 4061 1458 4073 1464
rect 4127 1458 4139 1464
rect 4173 1458 4185 1464
rect 4231 1458 4243 1464
rect 4291 1458 4303 1464
rect 4351 1458 4363 1472
rect 4439 1540 4445 1587
rect 4456 1582 4465 1620
rect 4456 1552 4465 1570
rect 4555 1582 4564 1620
rect 4575 1601 4581 1632
rect 4642 1626 4649 1648
rect 4699 1636 4701 1638
rect 4687 1632 4701 1636
rect 4642 1620 4684 1626
rect 4555 1552 4564 1570
rect 4456 1546 4497 1552
rect 4439 1536 4453 1540
rect 4439 1534 4441 1536
rect 4491 1512 4497 1546
rect 4523 1546 4564 1552
rect 4523 1512 4529 1546
rect 4575 1540 4581 1587
rect 4675 1582 4684 1620
rect 4695 1601 4701 1632
rect 4762 1626 4769 1648
rect 4819 1636 4821 1638
rect 4807 1632 4821 1636
rect 4762 1620 4804 1626
rect 4675 1552 4684 1570
rect 4643 1546 4684 1552
rect 4567 1536 4581 1540
rect 4579 1534 4581 1536
rect 4411 1458 4423 1464
rect 4471 1458 4483 1472
rect 4537 1458 4549 1472
rect 4643 1512 4649 1546
rect 4695 1540 4701 1587
rect 4795 1582 4804 1620
rect 4815 1601 4821 1632
rect 4882 1626 4889 1648
rect 4939 1636 4941 1638
rect 4927 1632 4941 1636
rect 4882 1620 4924 1626
rect 4795 1552 4804 1570
rect 4763 1546 4804 1552
rect 4687 1536 4701 1540
rect 4699 1534 4701 1536
rect 4597 1458 4609 1464
rect 4657 1458 4669 1472
rect 4763 1512 4769 1546
rect 4815 1540 4821 1587
rect 4915 1582 4924 1620
rect 4935 1601 4941 1632
rect 5167 1656 5180 1662
rect 5051 1650 5058 1656
rect 5047 1642 5058 1650
rect 5108 1644 5115 1656
rect 5173 1650 5180 1656
rect 4997 1621 5005 1636
rect 5108 1637 5129 1644
rect 5087 1626 5093 1628
rect 5154 1626 5161 1632
rect 4997 1607 5013 1621
rect 5087 1620 5161 1626
rect 4915 1552 4924 1570
rect 4883 1546 4924 1552
rect 4807 1536 4821 1540
rect 4819 1534 4821 1536
rect 4717 1458 4729 1464
rect 4777 1458 4789 1472
rect 4883 1512 4889 1546
rect 4935 1540 4941 1587
rect 4997 1544 5005 1607
rect 5013 1593 5027 1607
rect 5019 1548 5033 1556
rect 4927 1536 4941 1540
rect 4939 1534 4941 1536
rect 4837 1458 4849 1464
rect 4897 1458 4909 1472
rect 5087 1548 5093 1620
rect 5154 1612 5161 1620
rect 5166 1604 5200 1612
rect 5194 1599 5200 1604
rect 5147 1586 5174 1593
rect 5053 1542 5093 1548
rect 5101 1548 5145 1554
rect 5053 1524 5059 1542
rect 5101 1534 5107 1548
rect 5213 1552 5219 1636
rect 5157 1544 5219 1552
rect 5077 1528 5107 1534
rect 5125 1530 5163 1538
rect 5155 1524 5163 1530
rect 5047 1484 5059 1518
rect 5105 1510 5127 1522
rect 5155 1510 5173 1524
rect 5101 1504 5113 1510
rect 5155 1504 5163 1510
rect 5407 1656 5420 1662
rect 5291 1650 5298 1656
rect 5287 1642 5298 1650
rect 5348 1644 5355 1656
rect 5413 1650 5420 1656
rect 5237 1621 5245 1636
rect 5348 1637 5369 1644
rect 5617 1668 5629 1682
rect 5677 1668 5689 1682
rect 5771 1676 5783 1682
rect 5831 1676 5843 1682
rect 5871 1676 5883 1682
rect 5949 1676 5961 1682
rect 6031 1676 6043 1682
rect 6091 1676 6103 1682
rect 6131 1676 6143 1682
rect 6231 1676 6243 1682
rect 5327 1626 5333 1628
rect 5394 1626 5401 1632
rect 5237 1607 5253 1621
rect 5327 1620 5401 1626
rect 5237 1544 5245 1607
rect 5253 1593 5267 1607
rect 5259 1548 5273 1556
rect 5327 1548 5333 1620
rect 5394 1612 5401 1620
rect 5406 1604 5440 1612
rect 5434 1599 5440 1604
rect 5387 1586 5414 1593
rect 5293 1542 5333 1548
rect 5341 1548 5385 1554
rect 5293 1524 5299 1542
rect 5341 1534 5347 1548
rect 5453 1552 5459 1636
rect 5513 1593 5520 1636
rect 5602 1626 5609 1648
rect 5659 1636 5661 1638
rect 5647 1632 5661 1636
rect 5602 1620 5644 1626
rect 5397 1544 5459 1552
rect 5521 1556 5527 1579
rect 5635 1582 5644 1620
rect 5655 1601 5661 1632
rect 5735 1622 5743 1636
rect 5763 1636 5791 1642
rect 5751 1633 5803 1636
rect 5735 1615 5760 1622
rect 5717 1597 5733 1603
rect 5521 1550 5548 1556
rect 5635 1552 5644 1570
rect 5536 1544 5548 1550
rect 5603 1546 5644 1552
rect 5317 1528 5347 1534
rect 5365 1530 5403 1538
rect 5395 1524 5403 1530
rect 5287 1484 5299 1518
rect 5345 1510 5367 1522
rect 5395 1510 5413 1524
rect 5341 1504 5353 1510
rect 5395 1504 5403 1510
rect 5489 1536 5517 1542
rect 5529 1464 5557 1470
rect 5603 1512 5609 1546
rect 5655 1540 5661 1587
rect 5647 1536 5661 1540
rect 5659 1534 5661 1536
rect 4957 1458 4969 1464
rect 5017 1458 5029 1464
rect 5075 1458 5087 1464
rect 5121 1458 5133 1464
rect 5187 1458 5199 1464
rect 5257 1458 5269 1464
rect 5315 1458 5327 1464
rect 5361 1458 5373 1464
rect 5427 1458 5439 1464
rect 5497 1458 5509 1464
rect 5617 1458 5629 1472
rect 5717 1523 5723 1597
rect 5753 1593 5761 1615
rect 5853 1613 5860 1656
rect 5919 1628 5931 1636
rect 5887 1617 5903 1623
rect 5919 1622 5943 1628
rect 5759 1544 5767 1579
rect 5853 1551 5860 1599
rect 5843 1544 5860 1551
rect 5717 1517 5733 1523
rect 5677 1458 5689 1464
rect 5897 1523 5903 1617
rect 5935 1573 5943 1622
rect 5995 1622 6003 1636
rect 6023 1636 6051 1642
rect 6011 1633 6063 1636
rect 5995 1615 6020 1622
rect 6013 1593 6021 1615
rect 6113 1613 6120 1656
rect 6183 1670 6211 1676
rect 6223 1636 6251 1640
rect 6195 1626 6201 1636
rect 6211 1634 6263 1636
rect 6291 1668 6303 1682
rect 6351 1668 6363 1682
rect 6397 1676 6409 1682
rect 6479 1676 6491 1682
rect 6537 1676 6549 1682
rect 6585 1676 6597 1682
rect 6647 1676 6659 1682
rect 6319 1636 6321 1638
rect 6319 1632 6333 1636
rect 6195 1619 6224 1626
rect 5897 1517 5913 1523
rect 5935 1504 5943 1559
rect 6019 1544 6027 1579
rect 6113 1551 6120 1599
rect 6216 1593 6224 1619
rect 6319 1601 6325 1632
rect 6371 1626 6378 1648
rect 6336 1620 6378 1626
rect 6103 1544 6120 1551
rect 6215 1544 6223 1579
rect 5967 1517 5993 1523
rect 5736 1458 5748 1464
rect 5786 1458 5798 1464
rect 5871 1458 5883 1464
rect 5911 1458 5923 1464
rect 5951 1458 5963 1464
rect 5996 1458 6008 1464
rect 6046 1458 6058 1464
rect 6131 1458 6143 1464
rect 6181 1458 6193 1464
rect 6251 1458 6263 1464
rect 6319 1540 6325 1587
rect 6336 1582 6345 1620
rect 6336 1552 6345 1570
rect 6416 1601 6424 1656
rect 6627 1656 6640 1662
rect 6511 1650 6518 1656
rect 6507 1642 6518 1650
rect 6568 1644 6575 1656
rect 6633 1650 6640 1656
rect 6457 1621 6465 1636
rect 6568 1637 6589 1644
rect 6547 1626 6553 1628
rect 6614 1626 6621 1632
rect 6457 1607 6473 1621
rect 6547 1620 6621 1626
rect 6336 1546 6377 1552
rect 6319 1536 6333 1540
rect 6319 1534 6321 1536
rect 6371 1512 6377 1546
rect 6416 1504 6424 1587
rect 6457 1544 6465 1607
rect 6473 1593 6487 1607
rect 6479 1548 6493 1556
rect 6291 1458 6303 1464
rect 6351 1458 6363 1472
rect 6547 1548 6553 1620
rect 6614 1612 6621 1620
rect 6626 1604 6660 1612
rect 6654 1599 6660 1604
rect 6607 1586 6634 1593
rect 6513 1542 6553 1548
rect 6561 1548 6605 1554
rect 6513 1524 6519 1542
rect 6561 1534 6567 1548
rect 6673 1552 6679 1636
rect 6617 1544 6679 1552
rect 6537 1528 6567 1534
rect 6585 1530 6623 1538
rect 6615 1524 6623 1530
rect 6507 1484 6519 1518
rect 6565 1510 6587 1522
rect 6615 1510 6633 1524
rect 6561 1504 6573 1510
rect 6615 1504 6623 1510
rect 6397 1458 6409 1464
rect 6477 1458 6489 1464
rect 6535 1458 6547 1464
rect 6581 1458 6593 1464
rect 6647 1458 6659 1464
rect -62 1456 6736 1458
rect -62 1444 4 1456
rect -62 1442 173 1444
rect -62 978 -2 1442
rect 17 1436 29 1442
rect 61 1436 73 1442
rect 117 1436 129 1442
rect 38 1282 46 1396
rect 187 1442 6736 1444
rect 216 1436 228 1442
rect 266 1436 278 1442
rect 351 1436 363 1442
rect 377 1436 389 1442
rect 437 1436 449 1442
rect 511 1436 523 1442
rect 551 1436 563 1442
rect 597 1436 609 1442
rect 701 1436 713 1442
rect 767 1436 779 1442
rect 813 1436 825 1442
rect 871 1436 883 1442
rect 931 1436 943 1442
rect 971 1436 983 1442
rect 81 1321 89 1356
rect 140 1349 157 1356
rect 87 1307 89 1321
rect 17 1274 55 1282
rect 17 1264 29 1274
rect 81 1264 89 1307
rect 140 1301 147 1349
rect 239 1321 247 1356
rect 323 1349 340 1356
rect 79 1254 89 1264
rect 140 1244 147 1287
rect 233 1285 241 1307
rect 333 1301 340 1349
rect 396 1313 404 1396
rect 456 1313 464 1396
rect 535 1341 543 1396
rect 577 1362 589 1364
rect 577 1356 617 1362
rect 737 1390 745 1396
rect 787 1390 799 1396
rect 727 1376 745 1390
rect 773 1378 795 1390
rect 841 1382 853 1416
rect 737 1370 745 1376
rect 737 1362 775 1370
rect 793 1366 823 1372
rect 215 1278 240 1285
rect 215 1264 223 1278
rect 231 1264 283 1267
rect 243 1258 271 1264
rect 333 1244 340 1287
rect 396 1244 404 1299
rect 456 1244 464 1299
rect 535 1278 543 1327
rect 638 1321 646 1356
rect 681 1348 743 1356
rect 519 1272 543 1278
rect 519 1264 531 1272
rect 638 1264 646 1307
rect 47 1218 59 1224
rect 117 1218 129 1224
rect 157 1218 169 1224
rect 251 1218 263 1224
rect 311 1218 323 1224
rect 351 1218 363 1224
rect 377 1218 389 1224
rect 437 1218 449 1224
rect 549 1218 561 1224
rect 620 1253 646 1264
rect 681 1264 687 1348
rect 793 1352 799 1366
rect 841 1358 847 1376
rect 755 1346 799 1352
rect 807 1352 847 1358
rect 726 1307 753 1314
rect 700 1296 706 1301
rect 700 1288 734 1296
rect 739 1280 746 1288
rect 807 1280 813 1352
rect 997 1436 1009 1442
rect 1037 1436 1049 1442
rect 1097 1436 1109 1442
rect 1201 1436 1213 1442
rect 1267 1436 1279 1442
rect 1313 1436 1325 1442
rect 1371 1436 1383 1442
rect 1431 1436 1443 1442
rect 1471 1436 1483 1442
rect 1511 1436 1523 1442
rect 1551 1436 1563 1442
rect 1591 1436 1603 1442
rect 867 1344 881 1352
rect 873 1293 887 1307
rect 895 1293 903 1356
rect 955 1341 963 1396
rect 1018 1394 1029 1396
rect 1057 1394 1065 1396
rect 1018 1388 1065 1394
rect 739 1274 813 1280
rect 887 1279 903 1293
rect 739 1268 746 1274
rect 807 1272 813 1274
rect 771 1256 792 1263
rect 895 1264 903 1279
rect 955 1278 963 1327
rect 1058 1333 1065 1388
rect 1120 1349 1137 1356
rect 1237 1390 1245 1396
rect 1287 1390 1299 1396
rect 1227 1376 1245 1390
rect 1273 1378 1295 1390
rect 1341 1382 1353 1416
rect 1237 1370 1245 1376
rect 1237 1362 1275 1370
rect 1293 1366 1323 1372
rect 1056 1291 1064 1319
rect 1120 1301 1127 1349
rect 1181 1348 1243 1356
rect 720 1244 727 1250
rect 785 1244 792 1256
rect 842 1250 853 1258
rect 842 1244 849 1250
rect 720 1238 733 1244
rect 939 1272 963 1278
rect 939 1264 951 1272
rect 580 1218 592 1224
rect 630 1218 642 1224
rect 701 1218 713 1224
rect 763 1218 775 1224
rect 811 1218 823 1224
rect 869 1218 881 1224
rect 969 1218 981 1224
rect 1034 1282 1064 1291
rect 1046 1280 1064 1282
rect 1120 1244 1127 1287
rect 1181 1264 1187 1348
rect 1293 1352 1299 1366
rect 1341 1358 1347 1376
rect 1255 1346 1299 1352
rect 1307 1352 1347 1358
rect 1226 1307 1253 1314
rect 1200 1296 1206 1301
rect 1200 1288 1234 1296
rect 1239 1280 1246 1288
rect 1307 1280 1313 1352
rect 1631 1436 1643 1442
rect 1691 1428 1703 1442
rect 1791 1436 1803 1442
rect 1659 1364 1661 1366
rect 1659 1360 1673 1364
rect 1367 1344 1381 1352
rect 1373 1293 1387 1307
rect 1395 1293 1403 1356
rect 1451 1350 1463 1356
rect 1491 1350 1503 1356
rect 1531 1350 1543 1356
rect 1571 1350 1583 1356
rect 1445 1342 1463 1350
rect 1478 1342 1503 1350
rect 1518 1342 1543 1350
rect 1557 1342 1583 1350
rect 1445 1313 1452 1342
rect 1447 1299 1452 1313
rect 1239 1274 1313 1280
rect 1387 1279 1403 1293
rect 1239 1268 1246 1274
rect 1307 1272 1313 1274
rect 1271 1256 1292 1263
rect 1395 1264 1403 1279
rect 1445 1278 1452 1299
rect 1478 1296 1486 1342
rect 1518 1296 1526 1342
rect 1557 1296 1565 1342
rect 1659 1313 1665 1360
rect 1711 1354 1717 1388
rect 1676 1348 1717 1354
rect 1841 1436 1853 1442
rect 1911 1436 1923 1442
rect 1956 1436 1968 1442
rect 2006 1436 2018 1442
rect 2037 1436 2049 1442
rect 2102 1436 2114 1442
rect 2152 1436 2164 1442
rect 1763 1349 1780 1356
rect 1676 1330 1685 1348
rect 1470 1284 1486 1296
rect 1510 1284 1526 1296
rect 1550 1284 1565 1296
rect 1478 1278 1486 1284
rect 1518 1278 1526 1284
rect 1557 1278 1565 1284
rect 1445 1271 1464 1278
rect 1446 1270 1464 1271
rect 1478 1270 1504 1278
rect 1518 1270 1543 1278
rect 1557 1270 1584 1278
rect 1452 1264 1464 1270
rect 1492 1264 1504 1270
rect 1531 1264 1543 1270
rect 1572 1264 1584 1270
rect 1220 1244 1227 1250
rect 1285 1244 1292 1256
rect 1342 1250 1353 1258
rect 1342 1244 1349 1250
rect 1220 1238 1233 1244
rect 998 1218 1010 1224
rect 1097 1218 1109 1224
rect 1137 1218 1149 1224
rect 1201 1218 1213 1224
rect 1263 1218 1275 1224
rect 1311 1218 1323 1224
rect 1369 1218 1381 1224
rect 1431 1218 1443 1224
rect 1471 1218 1483 1224
rect 1511 1218 1523 1224
rect 1551 1218 1563 1224
rect 1591 1218 1603 1224
rect 1659 1268 1665 1299
rect 1676 1280 1685 1318
rect 1773 1301 1780 1349
rect 1875 1321 1883 1356
rect 1979 1321 1987 1356
rect 1676 1274 1718 1280
rect 1659 1264 1673 1268
rect 1659 1262 1661 1264
rect 1711 1252 1718 1274
rect 1773 1244 1780 1287
rect 1876 1281 1884 1307
rect 1973 1285 1981 1307
rect 2056 1313 2064 1396
rect 2197 1436 2209 1442
rect 2237 1436 2249 1442
rect 2297 1428 2309 1442
rect 2357 1436 2369 1442
rect 2133 1321 2141 1356
rect 1855 1274 1884 1281
rect 1955 1278 1980 1285
rect 1855 1264 1861 1274
rect 1871 1264 1923 1266
rect 1955 1264 1963 1278
rect 1631 1218 1643 1232
rect 1691 1218 1703 1232
rect 1843 1224 1871 1230
rect 1883 1260 1911 1264
rect 1971 1264 2023 1267
rect 1983 1258 2011 1264
rect 2056 1244 2064 1299
rect 2139 1285 2147 1307
rect 2177 1303 2183 1353
rect 2217 1341 2225 1396
rect 2283 1354 2289 1388
rect 2339 1364 2341 1366
rect 2327 1360 2341 1364
rect 2283 1348 2324 1354
rect 2167 1297 2183 1303
rect 2140 1278 2165 1285
rect 2097 1264 2149 1267
rect 2109 1258 2137 1264
rect 2157 1264 2165 1278
rect 2217 1278 2225 1327
rect 2315 1330 2324 1348
rect 2315 1280 2324 1318
rect 2335 1313 2341 1360
rect 2411 1436 2423 1442
rect 2471 1428 2483 1442
rect 2591 1436 2603 1442
rect 2657 1436 2669 1442
rect 2831 1436 2843 1442
rect 2899 1436 2911 1442
rect 3031 1436 3043 1442
rect 3111 1436 3123 1442
rect 2439 1364 2441 1366
rect 2439 1360 2453 1364
rect 2439 1313 2445 1360
rect 2491 1354 2497 1388
rect 2543 1430 2571 1436
rect 2583 1358 2611 1364
rect 2649 1358 2677 1364
rect 2689 1430 2717 1436
rect 2783 1430 2811 1436
rect 2823 1358 2851 1364
rect 2456 1348 2497 1354
rect 2552 1350 2564 1356
rect 2696 1350 2708 1356
rect 2456 1330 2465 1348
rect 2552 1344 2579 1350
rect 2217 1272 2241 1278
rect 2229 1264 2241 1272
rect 2282 1274 2324 1280
rect 2282 1252 2289 1274
rect 2335 1268 2341 1299
rect 2327 1264 2341 1268
rect 2339 1262 2341 1264
rect 1751 1218 1763 1224
rect 1791 1218 1803 1224
rect 1891 1218 1903 1224
rect 1991 1218 2003 1224
rect 2037 1218 2049 1224
rect 2117 1218 2129 1224
rect 2199 1218 2211 1224
rect 2297 1218 2309 1232
rect 2357 1218 2369 1232
rect 2439 1268 2445 1299
rect 2456 1280 2465 1318
rect 2573 1321 2579 1344
rect 2681 1344 2708 1350
rect 2792 1350 2804 1356
rect 2877 1350 2885 1396
rect 2983 1430 3011 1436
rect 3023 1358 3051 1364
rect 3151 1436 3163 1442
rect 2792 1344 2819 1350
rect 2877 1344 2903 1350
rect 2681 1321 2687 1344
rect 2813 1321 2819 1344
rect 2900 1338 2903 1344
rect 2456 1274 2498 1280
rect 2439 1264 2453 1268
rect 2439 1262 2441 1264
rect 2491 1252 2498 1274
rect 2580 1264 2587 1307
rect 2673 1264 2680 1307
rect 2820 1264 2827 1307
rect 2900 1282 2907 1338
rect 2921 1321 2929 1356
rect 2992 1350 3004 1356
rect 2992 1344 3019 1350
rect 3013 1321 3019 1344
rect 2927 1307 2929 1321
rect 2900 1276 2903 1282
rect 2881 1270 2903 1276
rect 2411 1218 2423 1232
rect 2471 1218 2483 1232
rect 2552 1218 2564 1224
rect 2608 1218 2620 1224
rect 2640 1218 2652 1224
rect 2696 1218 2708 1224
rect 2881 1244 2889 1270
rect 2921 1264 2929 1307
rect 3020 1264 3027 1307
rect 3096 1313 3104 1396
rect 3211 1428 3223 1442
rect 3281 1436 3293 1442
rect 3347 1436 3359 1442
rect 3393 1436 3405 1442
rect 3451 1436 3463 1442
rect 3551 1436 3563 1442
rect 3179 1364 3181 1366
rect 3179 1360 3193 1364
rect 3179 1313 3185 1360
rect 3231 1354 3237 1388
rect 3196 1348 3237 1354
rect 3317 1390 3325 1396
rect 3367 1390 3379 1396
rect 3307 1376 3325 1390
rect 3353 1378 3375 1390
rect 3421 1382 3433 1416
rect 3317 1370 3325 1376
rect 3317 1362 3355 1370
rect 3373 1366 3403 1372
rect 3261 1348 3323 1356
rect 3196 1330 3205 1348
rect 3096 1244 3104 1299
rect 2792 1218 2804 1224
rect 2848 1218 2860 1224
rect 2899 1218 2911 1224
rect 2992 1218 3004 1224
rect 3048 1218 3060 1224
rect 3111 1218 3123 1224
rect 3179 1268 3185 1299
rect 3196 1280 3205 1318
rect 3196 1274 3238 1280
rect 3179 1264 3193 1268
rect 3179 1262 3181 1264
rect 3231 1252 3238 1274
rect 3261 1264 3267 1348
rect 3373 1352 3379 1366
rect 3421 1358 3427 1376
rect 3335 1346 3379 1352
rect 3387 1352 3427 1358
rect 3306 1307 3333 1314
rect 3280 1296 3286 1301
rect 3280 1288 3314 1296
rect 3319 1280 3326 1288
rect 3387 1280 3393 1352
rect 3447 1344 3461 1352
rect 3453 1293 3467 1307
rect 3475 1293 3483 1356
rect 3601 1436 3613 1442
rect 3671 1436 3683 1442
rect 3716 1436 3728 1442
rect 3766 1436 3778 1442
rect 3831 1436 3843 1442
rect 3877 1436 3889 1442
rect 3935 1436 3947 1442
rect 3981 1436 3993 1442
rect 4047 1436 4059 1442
rect 4117 1436 4129 1442
rect 4175 1436 4187 1442
rect 4221 1436 4233 1442
rect 4287 1436 4299 1442
rect 4371 1436 4383 1442
rect 4417 1436 4429 1442
rect 3523 1349 3540 1356
rect 3319 1274 3393 1280
rect 3467 1279 3483 1293
rect 3319 1268 3326 1274
rect 3387 1272 3393 1274
rect 3151 1218 3163 1232
rect 3211 1218 3223 1232
rect 3351 1256 3372 1263
rect 3475 1264 3483 1279
rect 3300 1244 3307 1250
rect 3365 1244 3372 1256
rect 3422 1250 3433 1258
rect 3422 1244 3429 1250
rect 3300 1238 3313 1244
rect 3533 1301 3540 1349
rect 3635 1321 3643 1356
rect 3739 1321 3747 1356
rect 3533 1244 3540 1287
rect 3577 1283 3583 1313
rect 3577 1277 3593 1283
rect 3636 1281 3644 1307
rect 3697 1297 3713 1303
rect 3615 1274 3644 1281
rect 3615 1264 3621 1274
rect 3697 1283 3703 1297
rect 3733 1285 3741 1307
rect 3816 1313 3824 1396
rect 3907 1382 3919 1416
rect 3961 1390 3973 1396
rect 4015 1390 4023 1396
rect 3965 1378 3987 1390
rect 4015 1376 4033 1390
rect 3913 1358 3919 1376
rect 3937 1366 3967 1372
rect 4015 1370 4023 1376
rect 3687 1277 3703 1283
rect 3715 1278 3740 1285
rect 3631 1264 3683 1266
rect 3715 1264 3723 1278
rect 3603 1224 3631 1230
rect 3643 1260 3671 1264
rect 3731 1264 3783 1267
rect 3743 1258 3771 1264
rect 3816 1244 3824 1299
rect 3857 1293 3865 1356
rect 3879 1344 3893 1352
rect 3913 1352 3953 1358
rect 3873 1293 3887 1307
rect 3857 1279 3873 1293
rect 3947 1280 3953 1352
rect 3961 1352 3967 1366
rect 3985 1362 4023 1370
rect 3961 1346 4005 1352
rect 4017 1348 4079 1356
rect 4007 1307 4034 1314
rect 4054 1296 4060 1301
rect 4026 1288 4060 1296
rect 4014 1280 4021 1288
rect 3857 1264 3865 1279
rect 3947 1274 4021 1280
rect 3947 1272 3953 1274
rect 4014 1268 4021 1274
rect 3907 1250 3918 1258
rect 3911 1244 3918 1250
rect 3968 1256 3989 1263
rect 4073 1264 4079 1348
rect 3968 1244 3975 1256
rect 4033 1244 4040 1250
rect 4027 1238 4040 1244
rect 4147 1382 4159 1416
rect 4201 1390 4213 1396
rect 4255 1390 4263 1396
rect 4205 1378 4227 1390
rect 4255 1376 4273 1390
rect 4153 1358 4159 1376
rect 4177 1366 4207 1372
rect 4255 1370 4263 1376
rect 4097 1293 4105 1356
rect 4119 1344 4133 1352
rect 4153 1352 4193 1358
rect 4113 1293 4127 1307
rect 4097 1279 4113 1293
rect 4187 1280 4193 1352
rect 4201 1352 4207 1366
rect 4225 1362 4263 1370
rect 4201 1346 4245 1352
rect 4257 1348 4319 1356
rect 4247 1307 4274 1314
rect 4294 1296 4300 1301
rect 4266 1288 4300 1296
rect 4254 1280 4261 1288
rect 4097 1264 4105 1279
rect 4187 1274 4261 1280
rect 4187 1272 4193 1274
rect 4254 1268 4261 1274
rect 4147 1250 4158 1258
rect 4151 1244 4158 1250
rect 4208 1256 4229 1263
rect 4313 1264 4319 1348
rect 4337 1287 4343 1353
rect 4356 1313 4364 1396
rect 4409 1358 4437 1364
rect 4449 1430 4477 1436
rect 4537 1428 4549 1442
rect 4597 1436 4609 1442
rect 4711 1436 4723 1442
rect 4789 1436 4801 1442
rect 4851 1436 4863 1442
rect 4891 1436 4903 1442
rect 4456 1350 4468 1356
rect 4441 1344 4468 1350
rect 4523 1354 4529 1388
rect 4579 1364 4581 1366
rect 4567 1360 4581 1364
rect 4523 1348 4564 1354
rect 4441 1321 4447 1344
rect 4208 1244 4215 1256
rect 4273 1244 4280 1250
rect 4267 1238 4280 1244
rect 4356 1244 4364 1299
rect 4433 1264 4440 1307
rect 4555 1330 4564 1348
rect 4555 1280 4564 1318
rect 4575 1313 4581 1360
rect 4663 1430 4691 1436
rect 4703 1358 4731 1364
rect 4931 1436 4943 1442
rect 4971 1436 4983 1442
rect 5021 1436 5033 1442
rect 5091 1436 5103 1442
rect 4672 1350 4684 1356
rect 4672 1344 4699 1350
rect 4627 1337 4643 1343
rect 4522 1274 4564 1280
rect 3281 1218 3293 1224
rect 3343 1218 3355 1224
rect 3391 1218 3403 1224
rect 3449 1218 3461 1224
rect 3511 1218 3523 1224
rect 3551 1218 3563 1224
rect 3651 1218 3663 1224
rect 3751 1218 3763 1224
rect 3831 1218 3843 1224
rect 3879 1218 3891 1224
rect 3937 1218 3949 1224
rect 3985 1218 3997 1224
rect 4047 1218 4059 1224
rect 4119 1218 4131 1224
rect 4177 1218 4189 1224
rect 4225 1218 4237 1224
rect 4287 1218 4299 1224
rect 4371 1218 4383 1224
rect 4522 1252 4529 1274
rect 4575 1268 4581 1299
rect 4637 1283 4643 1337
rect 4693 1321 4699 1344
rect 4771 1321 4779 1356
rect 4815 1350 4823 1396
rect 4797 1344 4823 1350
rect 4797 1338 4800 1344
rect 4875 1341 4883 1396
rect 4937 1363 4943 1373
rect 4917 1357 4943 1363
rect 4637 1277 4653 1283
rect 4567 1264 4581 1268
rect 4579 1262 4581 1264
rect 4700 1264 4707 1307
rect 4771 1307 4773 1321
rect 4771 1264 4779 1307
rect 4793 1282 4800 1338
rect 4797 1276 4800 1282
rect 4875 1278 4883 1327
rect 4797 1270 4819 1276
rect 4400 1218 4412 1224
rect 4456 1218 4468 1224
rect 4537 1218 4549 1232
rect 4597 1218 4609 1232
rect 4811 1244 4819 1270
rect 4859 1272 4883 1278
rect 4917 1283 4923 1357
rect 4955 1341 4963 1396
rect 5141 1436 5153 1442
rect 5211 1436 5223 1442
rect 4907 1277 4923 1283
rect 4955 1278 4963 1327
rect 5055 1321 5063 1356
rect 5237 1436 5249 1442
rect 5311 1436 5323 1442
rect 5351 1436 5363 1442
rect 5377 1436 5389 1442
rect 5447 1436 5459 1442
rect 5551 1436 5563 1442
rect 5597 1436 5609 1442
rect 5056 1281 5064 1307
rect 4939 1272 4963 1278
rect 5035 1274 5064 1281
rect 5117 1283 5123 1353
rect 5175 1321 5183 1356
rect 5256 1321 5264 1356
rect 5335 1341 5343 1396
rect 5571 1362 5583 1364
rect 5543 1356 5583 1362
rect 5677 1428 5689 1442
rect 5737 1436 5749 1442
rect 5117 1277 5133 1283
rect 4859 1264 4871 1272
rect 4939 1264 4951 1272
rect 5035 1264 5041 1274
rect 5176 1281 5184 1307
rect 5155 1274 5184 1281
rect 5051 1264 5103 1266
rect 5155 1264 5161 1274
rect 5171 1264 5223 1266
rect 5256 1264 5264 1307
rect 5335 1278 5343 1327
rect 5417 1321 5425 1356
rect 5319 1272 5343 1278
rect 5416 1281 5424 1307
rect 5416 1274 5445 1281
rect 5319 1264 5331 1272
rect 5377 1264 5429 1266
rect 5439 1264 5445 1274
rect 5497 1283 5503 1333
rect 5514 1321 5522 1356
rect 5616 1321 5624 1356
rect 5663 1354 5669 1388
rect 5719 1364 5721 1366
rect 5707 1360 5721 1364
rect 5663 1348 5704 1354
rect 5467 1277 5503 1283
rect 5514 1264 5522 1307
rect 5616 1264 5624 1307
rect 5695 1330 5704 1348
rect 5695 1280 5704 1318
rect 5715 1313 5721 1360
rect 5791 1436 5803 1442
rect 5831 1436 5843 1442
rect 5876 1436 5888 1442
rect 5926 1436 5938 1442
rect 5991 1436 6003 1442
rect 5815 1341 5823 1396
rect 6022 1436 6034 1442
rect 6072 1436 6084 1442
rect 5662 1274 5704 1280
rect 5023 1224 5051 1230
rect 5063 1260 5091 1264
rect 5143 1224 5171 1230
rect 5183 1260 5211 1264
rect 5389 1260 5417 1264
rect 5429 1224 5457 1230
rect 5514 1253 5540 1264
rect 4672 1218 4684 1224
rect 4728 1218 4740 1224
rect 4789 1218 4801 1224
rect 4889 1218 4901 1224
rect 4969 1218 4981 1224
rect 5071 1218 5083 1224
rect 5191 1218 5203 1224
rect 5237 1218 5249 1224
rect 5349 1218 5361 1224
rect 5397 1218 5409 1224
rect 5518 1218 5530 1224
rect 5568 1218 5580 1224
rect 5662 1252 5669 1274
rect 5715 1268 5721 1299
rect 5815 1278 5823 1327
rect 5899 1321 5907 1356
rect 5893 1285 5901 1307
rect 5976 1313 5984 1396
rect 6117 1436 6129 1442
rect 6187 1436 6199 1442
rect 6257 1436 6269 1442
rect 6315 1436 6327 1442
rect 6361 1436 6373 1442
rect 6427 1436 6439 1442
rect 6497 1436 6509 1442
rect 6555 1436 6567 1442
rect 6601 1436 6613 1442
rect 6667 1436 6679 1442
rect 6087 1377 6103 1383
rect 6053 1321 6061 1356
rect 5799 1272 5823 1278
rect 5875 1278 5900 1285
rect 5707 1264 5721 1268
rect 5719 1262 5721 1264
rect 5597 1218 5609 1224
rect 5677 1218 5689 1232
rect 5737 1218 5749 1232
rect 5799 1264 5811 1272
rect 5875 1264 5883 1278
rect 5891 1264 5943 1267
rect 5903 1258 5931 1264
rect 5976 1244 5984 1299
rect 6059 1285 6067 1307
rect 6060 1278 6085 1285
rect 6017 1264 6069 1267
rect 6029 1258 6057 1264
rect 6077 1264 6085 1278
rect 6097 1283 6103 1377
rect 6287 1382 6299 1416
rect 6341 1390 6353 1396
rect 6395 1390 6403 1396
rect 6345 1378 6367 1390
rect 6395 1376 6413 1390
rect 6293 1358 6299 1376
rect 6317 1366 6347 1372
rect 6395 1370 6403 1376
rect 6157 1321 6165 1356
rect 6097 1277 6113 1283
rect 6156 1281 6164 1307
rect 6237 1293 6245 1356
rect 6259 1344 6273 1352
rect 6293 1352 6333 1358
rect 6253 1293 6267 1307
rect 6156 1274 6185 1281
rect 6117 1264 6169 1266
rect 6179 1264 6185 1274
rect 6237 1279 6253 1293
rect 6327 1280 6333 1352
rect 6341 1352 6347 1366
rect 6365 1362 6403 1370
rect 6341 1346 6385 1352
rect 6397 1348 6459 1356
rect 6387 1307 6414 1314
rect 6434 1296 6440 1301
rect 6406 1288 6440 1296
rect 6394 1280 6401 1288
rect 6237 1264 6245 1279
rect 6327 1274 6401 1280
rect 6327 1272 6333 1274
rect 6129 1260 6157 1264
rect 6169 1224 6197 1230
rect 6394 1268 6401 1274
rect 6287 1250 6298 1258
rect 6291 1244 6298 1250
rect 6348 1256 6369 1263
rect 6453 1264 6459 1348
rect 6348 1244 6355 1256
rect 6413 1244 6420 1250
rect 6407 1238 6420 1244
rect 6527 1382 6539 1416
rect 6581 1390 6593 1396
rect 6635 1390 6643 1396
rect 6585 1378 6607 1390
rect 6635 1376 6653 1390
rect 6533 1358 6539 1376
rect 6557 1366 6587 1372
rect 6635 1370 6643 1376
rect 6477 1293 6485 1356
rect 6499 1344 6513 1352
rect 6533 1352 6573 1358
rect 6493 1293 6507 1307
rect 6477 1279 6493 1293
rect 6567 1280 6573 1352
rect 6581 1352 6587 1366
rect 6605 1362 6643 1370
rect 6581 1346 6625 1352
rect 6637 1348 6699 1356
rect 6627 1307 6654 1314
rect 6674 1296 6680 1301
rect 6646 1288 6680 1296
rect 6634 1280 6641 1288
rect 6477 1264 6485 1279
rect 6567 1274 6641 1280
rect 6567 1272 6573 1274
rect 6634 1268 6641 1274
rect 6527 1250 6538 1258
rect 6531 1244 6538 1250
rect 6588 1256 6609 1263
rect 6693 1264 6699 1348
rect 6588 1244 6595 1256
rect 6653 1244 6660 1250
rect 6647 1238 6660 1244
rect 5829 1218 5841 1224
rect 5911 1218 5923 1224
rect 5991 1218 6003 1224
rect 6037 1218 6049 1224
rect 6137 1218 6149 1224
rect 6259 1218 6271 1224
rect 6317 1218 6329 1224
rect 6365 1218 6377 1224
rect 6427 1218 6439 1224
rect 6499 1218 6511 1224
rect 6557 1218 6569 1224
rect 6605 1218 6617 1224
rect 6667 1218 6679 1224
rect 6742 1218 6802 1682
rect 4 1216 6802 1218
rect 6736 1204 6802 1216
rect 4 1202 6802 1204
rect 39 1196 51 1202
rect 97 1196 109 1202
rect 145 1196 157 1202
rect 207 1196 219 1202
rect 291 1196 303 1202
rect 339 1196 351 1202
rect 397 1196 409 1202
rect 445 1196 457 1202
rect 507 1196 519 1202
rect 557 1196 569 1202
rect 618 1196 630 1202
rect 717 1196 729 1202
rect 757 1196 769 1202
rect 187 1176 200 1182
rect 71 1170 78 1176
rect 67 1162 78 1170
rect 128 1164 135 1176
rect 193 1170 200 1176
rect 17 1141 25 1156
rect 128 1157 149 1164
rect 107 1146 113 1148
rect 174 1146 181 1152
rect 17 1127 33 1141
rect 107 1140 181 1146
rect 17 1064 25 1127
rect 33 1113 47 1127
rect 39 1068 53 1076
rect 107 1068 113 1140
rect 174 1132 181 1140
rect 186 1124 220 1132
rect 214 1119 220 1124
rect 167 1106 194 1113
rect 73 1062 113 1068
rect 121 1068 165 1074
rect 73 1044 79 1062
rect 121 1054 127 1068
rect 233 1072 239 1156
rect 276 1121 284 1176
rect 487 1176 500 1182
rect 371 1170 378 1176
rect 367 1162 378 1170
rect 428 1164 435 1176
rect 493 1170 500 1176
rect 317 1141 325 1156
rect 428 1157 449 1164
rect 407 1146 413 1148
rect 474 1146 481 1152
rect 317 1127 333 1141
rect 407 1140 481 1146
rect 177 1064 239 1072
rect 97 1048 127 1054
rect 145 1050 183 1058
rect 175 1044 183 1050
rect 67 1004 79 1038
rect 125 1030 147 1042
rect 175 1030 193 1044
rect 121 1024 133 1030
rect 175 1024 183 1030
rect 276 1024 284 1107
rect 317 1064 325 1127
rect 333 1113 347 1127
rect 339 1068 353 1076
rect 407 1068 413 1140
rect 474 1132 481 1140
rect 486 1124 520 1132
rect 514 1119 520 1124
rect 467 1106 494 1113
rect 373 1062 413 1068
rect 421 1068 465 1074
rect 373 1044 379 1062
rect 421 1054 427 1068
rect 533 1072 539 1156
rect 576 1121 584 1176
rect 798 1196 810 1202
rect 899 1196 911 1202
rect 977 1196 989 1202
rect 1061 1196 1073 1202
rect 1123 1196 1135 1202
rect 1171 1196 1183 1202
rect 1229 1196 1241 1202
rect 1277 1196 1289 1202
rect 1317 1196 1329 1202
rect 1357 1196 1369 1202
rect 1397 1196 1409 1202
rect 1437 1196 1449 1202
rect 1501 1196 1513 1202
rect 1563 1196 1575 1202
rect 1611 1196 1623 1202
rect 1669 1196 1681 1202
rect 1731 1196 1743 1202
rect 1771 1196 1783 1202
rect 1871 1196 1883 1202
rect 1971 1196 1983 1202
rect 2071 1196 2083 1202
rect 2131 1196 2143 1202
rect 2171 1196 2183 1202
rect 2271 1196 2283 1202
rect 2341 1196 2353 1202
rect 2403 1196 2415 1202
rect 2451 1196 2463 1202
rect 2509 1196 2521 1202
rect 2591 1196 2603 1202
rect 2637 1196 2649 1202
rect 2749 1196 2761 1202
rect 2797 1196 2809 1202
rect 2892 1196 2904 1202
rect 2948 1196 2960 1202
rect 3001 1196 3013 1202
rect 3063 1196 3075 1202
rect 3111 1196 3123 1202
rect 3169 1196 3181 1202
rect 3219 1196 3231 1202
rect 666 1138 684 1140
rect 654 1129 684 1138
rect 740 1133 747 1176
rect 929 1148 941 1156
rect 917 1142 941 1148
rect 846 1138 864 1140
rect 597 1117 633 1123
rect 477 1064 539 1072
rect 397 1048 427 1054
rect 445 1050 483 1058
rect 475 1044 483 1050
rect 367 1004 379 1038
rect 425 1030 447 1042
rect 475 1030 493 1044
rect 421 1024 433 1030
rect 475 1024 483 1030
rect 576 1024 584 1107
rect 597 1043 603 1117
rect 676 1101 684 1129
rect 834 1129 864 1138
rect 597 1037 613 1043
rect 678 1032 685 1087
rect 740 1071 747 1119
rect 787 1117 813 1123
rect 856 1101 864 1129
rect 917 1093 925 1142
rect 996 1121 1004 1176
rect 1080 1176 1093 1182
rect 1080 1170 1087 1176
rect 1145 1164 1152 1176
rect 740 1064 757 1071
rect 638 1026 685 1032
rect 638 1024 649 1026
rect 677 1024 685 1026
rect 858 1032 865 1087
rect 818 1026 865 1032
rect 818 1024 829 1026
rect 857 1024 865 1026
rect 917 1024 925 1079
rect 996 1024 1004 1107
rect 1041 1072 1047 1156
rect 1131 1157 1152 1164
rect 1202 1170 1209 1176
rect 1202 1162 1213 1170
rect 1099 1146 1106 1152
rect 1520 1176 1533 1182
rect 1520 1170 1527 1176
rect 1585 1164 1592 1176
rect 1167 1146 1173 1148
rect 1099 1140 1173 1146
rect 1255 1141 1263 1156
rect 1296 1150 1308 1156
rect 1337 1150 1349 1156
rect 1376 1150 1388 1156
rect 1416 1150 1428 1156
rect 1296 1142 1323 1150
rect 1337 1142 1362 1150
rect 1376 1142 1402 1150
rect 1416 1149 1434 1150
rect 1416 1142 1435 1149
rect 1099 1132 1106 1140
rect 1060 1124 1094 1132
rect 1060 1119 1066 1124
rect 1086 1106 1113 1113
rect 1041 1064 1103 1072
rect 1115 1068 1159 1074
rect 37 978 49 984
rect 95 978 107 984
rect 141 978 153 984
rect 207 978 219 984
rect 291 978 303 984
rect 337 978 349 984
rect 395 978 407 984
rect 441 978 453 984
rect 507 978 519 984
rect 557 978 569 984
rect 617 978 629 984
rect 657 978 669 984
rect 717 978 729 984
rect 797 978 809 984
rect 837 978 849 984
rect 897 978 909 984
rect 937 978 949 984
rect 1097 1050 1135 1058
rect 1153 1054 1159 1068
rect 1167 1068 1173 1140
rect 1247 1127 1263 1141
rect 1315 1136 1323 1142
rect 1354 1136 1362 1142
rect 1394 1136 1402 1142
rect 1233 1113 1247 1127
rect 1167 1062 1207 1068
rect 1227 1068 1241 1076
rect 1255 1064 1263 1127
rect 1315 1124 1330 1136
rect 1354 1124 1370 1136
rect 1394 1124 1410 1136
rect 1315 1078 1323 1124
rect 1354 1078 1362 1124
rect 1394 1078 1402 1124
rect 1428 1121 1435 1142
rect 1428 1107 1433 1121
rect 1428 1078 1435 1107
rect 1297 1070 1323 1078
rect 1337 1070 1362 1078
rect 1377 1070 1402 1078
rect 1417 1070 1435 1078
rect 1481 1072 1487 1156
rect 1571 1157 1592 1164
rect 1642 1170 1649 1176
rect 1642 1162 1653 1170
rect 1539 1146 1546 1152
rect 1607 1146 1613 1148
rect 1539 1140 1613 1146
rect 1695 1141 1703 1156
rect 1539 1132 1546 1140
rect 1500 1124 1534 1132
rect 1500 1119 1506 1124
rect 1526 1106 1553 1113
rect 1297 1064 1309 1070
rect 1337 1064 1349 1070
rect 1377 1064 1389 1070
rect 1417 1064 1429 1070
rect 1481 1064 1543 1072
rect 1555 1068 1599 1074
rect 1097 1044 1105 1050
rect 1153 1048 1183 1054
rect 1201 1044 1207 1062
rect 1087 1030 1105 1044
rect 1133 1030 1155 1042
rect 1097 1024 1105 1030
rect 1147 1024 1159 1030
rect 1201 1004 1213 1038
rect 1537 1050 1575 1058
rect 1593 1054 1599 1068
rect 1607 1068 1613 1140
rect 1687 1127 1703 1141
rect 1673 1113 1687 1127
rect 1607 1062 1647 1068
rect 1667 1068 1681 1076
rect 1695 1064 1703 1127
rect 1753 1133 1760 1176
rect 1823 1190 1851 1196
rect 1863 1156 1891 1160
rect 1835 1146 1841 1156
rect 1851 1154 1903 1156
rect 1835 1139 1864 1146
rect 1753 1071 1760 1119
rect 1856 1113 1864 1139
rect 1935 1142 1943 1156
rect 1963 1156 1991 1162
rect 1951 1153 2003 1156
rect 1935 1135 1960 1142
rect 1953 1113 1961 1135
rect 2007 1137 2023 1143
rect 1537 1044 1545 1050
rect 1593 1048 1623 1054
rect 1641 1044 1647 1062
rect 1527 1030 1545 1044
rect 1573 1030 1595 1042
rect 1537 1024 1545 1030
rect 1587 1024 1599 1030
rect 1641 1004 1653 1038
rect 1743 1064 1760 1071
rect 1855 1064 1863 1099
rect 1959 1064 1967 1099
rect 977 978 989 984
rect 1061 978 1073 984
rect 1127 978 1139 984
rect 1173 978 1185 984
rect 1231 978 1243 984
rect 1277 978 1289 984
rect 1317 978 1329 984
rect 1357 978 1369 984
rect 1397 978 1409 984
rect 1437 978 1449 984
rect 1501 978 1513 984
rect 1567 978 1579 984
rect 1613 978 1625 984
rect 1671 978 1683 984
rect 1771 978 1783 984
rect 1821 978 1833 984
rect 1891 978 1903 984
rect 2017 1043 2023 1137
rect 2035 1142 2043 1156
rect 2063 1156 2091 1162
rect 2051 1153 2103 1156
rect 2035 1135 2060 1142
rect 2053 1113 2061 1135
rect 2153 1133 2160 1176
rect 2223 1190 2251 1196
rect 2263 1156 2291 1160
rect 2235 1146 2241 1156
rect 2251 1154 2303 1156
rect 2360 1176 2373 1182
rect 2360 1170 2367 1176
rect 2425 1164 2432 1176
rect 2235 1139 2264 1146
rect 2059 1064 2067 1099
rect 2153 1071 2160 1119
rect 2256 1113 2264 1139
rect 2143 1064 2160 1071
rect 2255 1064 2263 1099
rect 2321 1072 2327 1156
rect 2411 1157 2432 1164
rect 2482 1170 2489 1176
rect 2482 1162 2493 1170
rect 2379 1146 2386 1152
rect 2447 1146 2453 1148
rect 2379 1140 2453 1146
rect 2535 1141 2543 1156
rect 2379 1132 2386 1140
rect 2340 1124 2374 1132
rect 2340 1119 2346 1124
rect 2366 1106 2393 1113
rect 2321 1064 2383 1072
rect 2395 1068 2439 1074
rect 2017 1037 2033 1043
rect 1936 978 1948 984
rect 1986 978 1998 984
rect 2036 978 2048 984
rect 2086 978 2098 984
rect 2171 978 2183 984
rect 2377 1050 2415 1058
rect 2433 1054 2439 1068
rect 2447 1068 2453 1140
rect 2527 1127 2543 1141
rect 2513 1113 2527 1127
rect 2447 1062 2487 1068
rect 2507 1068 2521 1076
rect 2535 1064 2543 1127
rect 2576 1121 2584 1176
rect 2629 1156 2657 1162
rect 2617 1153 2669 1156
rect 2677 1142 2685 1156
rect 2660 1135 2685 1142
rect 2377 1044 2385 1050
rect 2433 1048 2463 1054
rect 2481 1044 2487 1062
rect 2367 1030 2385 1044
rect 2413 1030 2435 1042
rect 2377 1024 2385 1030
rect 2427 1024 2439 1030
rect 2481 1004 2493 1038
rect 2576 1024 2584 1107
rect 2659 1113 2667 1135
rect 2731 1113 2739 1156
rect 2771 1150 2779 1176
rect 2757 1144 2779 1150
rect 2757 1138 2760 1144
rect 2731 1099 2733 1113
rect 2653 1064 2661 1099
rect 2731 1064 2739 1099
rect 2753 1082 2760 1138
rect 2816 1121 2824 1176
rect 3020 1176 3033 1182
rect 3020 1170 3027 1176
rect 3085 1164 3092 1176
rect 2757 1076 2760 1082
rect 2757 1070 2783 1076
rect 2221 978 2233 984
rect 2291 978 2303 984
rect 2341 978 2353 984
rect 2407 978 2419 984
rect 2453 978 2465 984
rect 2511 978 2523 984
rect 2591 978 2603 984
rect 2775 1024 2783 1070
rect 2816 1024 2824 1107
rect 2920 1113 2927 1156
rect 2913 1076 2919 1099
rect 2892 1070 2919 1076
rect 2981 1072 2987 1156
rect 3071 1157 3092 1164
rect 3142 1170 3149 1176
rect 3142 1162 3153 1170
rect 3039 1146 3046 1152
rect 3107 1146 3113 1148
rect 3039 1140 3113 1146
rect 3195 1141 3203 1156
rect 3249 1148 3261 1156
rect 3311 1188 3323 1202
rect 3371 1188 3383 1202
rect 3437 1188 3449 1202
rect 3497 1188 3509 1202
rect 3569 1196 3581 1202
rect 3641 1196 3653 1202
rect 3703 1196 3715 1202
rect 3751 1196 3763 1202
rect 3809 1196 3821 1202
rect 3339 1156 3341 1158
rect 3339 1152 3353 1156
rect 3039 1132 3046 1140
rect 3000 1124 3034 1132
rect 3000 1119 3006 1124
rect 3026 1106 3053 1113
rect 2892 1064 2904 1070
rect 2981 1064 3043 1072
rect 3055 1068 3099 1074
rect 2883 984 2911 990
rect 2923 1056 2951 1062
rect 3037 1050 3075 1058
rect 3093 1054 3099 1068
rect 3107 1068 3113 1140
rect 3187 1127 3203 1141
rect 3173 1113 3187 1127
rect 3107 1062 3147 1068
rect 3167 1068 3181 1076
rect 3195 1064 3203 1127
rect 3237 1142 3261 1148
rect 3237 1093 3245 1142
rect 3339 1121 3345 1152
rect 3391 1146 3398 1168
rect 3356 1140 3398 1146
rect 3422 1146 3429 1168
rect 3479 1156 3481 1158
rect 3467 1152 3481 1156
rect 3422 1140 3464 1146
rect 3037 1044 3045 1050
rect 3093 1048 3123 1054
rect 3141 1044 3147 1062
rect 3027 1030 3045 1044
rect 3073 1030 3095 1042
rect 3037 1024 3045 1030
rect 3087 1024 3099 1030
rect 3141 1004 3153 1038
rect 3237 1024 3245 1079
rect 2622 978 2634 984
rect 2672 978 2684 984
rect 2749 978 2761 984
rect 2797 978 2809 984
rect 2931 978 2943 984
rect 3001 978 3013 984
rect 3067 978 3079 984
rect 3113 978 3125 984
rect 3171 978 3183 984
rect 3217 978 3229 984
rect 3257 978 3269 984
rect 3339 1060 3345 1107
rect 3356 1102 3365 1140
rect 3356 1072 3365 1090
rect 3455 1102 3464 1140
rect 3475 1121 3481 1152
rect 3551 1113 3559 1156
rect 3591 1150 3599 1176
rect 3577 1144 3599 1150
rect 3660 1176 3673 1182
rect 3660 1170 3667 1176
rect 3725 1164 3732 1176
rect 3577 1138 3580 1144
rect 3455 1072 3464 1090
rect 3356 1066 3397 1072
rect 3339 1056 3353 1060
rect 3339 1054 3341 1056
rect 3391 1032 3397 1066
rect 3423 1066 3464 1072
rect 3423 1032 3429 1066
rect 3475 1060 3481 1107
rect 3551 1099 3553 1113
rect 3551 1064 3559 1099
rect 3573 1082 3580 1138
rect 3577 1076 3580 1082
rect 3577 1070 3603 1076
rect 3467 1056 3481 1060
rect 3479 1054 3481 1056
rect 3311 978 3323 984
rect 3371 978 3383 992
rect 3437 978 3449 992
rect 3595 1024 3603 1070
rect 3621 1072 3627 1156
rect 3711 1157 3732 1164
rect 3782 1170 3789 1176
rect 3782 1162 3793 1170
rect 3679 1146 3686 1152
rect 3877 1188 3889 1202
rect 3937 1188 3949 1202
rect 3747 1146 3753 1148
rect 3679 1140 3753 1146
rect 3835 1141 3843 1156
rect 3679 1132 3686 1140
rect 3640 1124 3674 1132
rect 3640 1119 3646 1124
rect 3666 1106 3693 1113
rect 3621 1064 3683 1072
rect 3695 1068 3739 1074
rect 3677 1050 3715 1058
rect 3733 1054 3739 1068
rect 3747 1068 3753 1140
rect 3827 1127 3843 1141
rect 3862 1146 3869 1168
rect 3919 1156 3921 1158
rect 3907 1152 3921 1156
rect 3862 1140 3904 1146
rect 3813 1113 3827 1127
rect 3747 1062 3787 1068
rect 3807 1068 3821 1076
rect 3835 1064 3843 1127
rect 3895 1102 3904 1140
rect 3915 1121 3921 1152
rect 3991 1188 4003 1202
rect 4051 1188 4063 1202
rect 4097 1196 4109 1202
rect 4177 1196 4189 1202
rect 4277 1196 4289 1202
rect 4317 1196 4329 1202
rect 4411 1196 4423 1202
rect 4478 1196 4490 1202
rect 4528 1196 4540 1202
rect 4581 1196 4593 1202
rect 4643 1196 4655 1202
rect 4691 1196 4703 1202
rect 4749 1196 4761 1202
rect 4817 1196 4829 1202
rect 4931 1196 4943 1202
rect 4971 1196 4983 1202
rect 5051 1196 5063 1202
rect 5111 1196 5123 1202
rect 5151 1196 5163 1202
rect 4019 1156 4021 1158
rect 4019 1152 4033 1156
rect 4019 1121 4025 1152
rect 4071 1146 4078 1168
rect 4036 1140 4078 1146
rect 3895 1072 3904 1090
rect 3677 1044 3685 1050
rect 3733 1048 3763 1054
rect 3781 1044 3787 1062
rect 3667 1030 3685 1044
rect 3713 1030 3735 1042
rect 3677 1024 3685 1030
rect 3727 1024 3739 1030
rect 3781 1004 3793 1038
rect 3863 1066 3904 1072
rect 3863 1032 3869 1066
rect 3915 1060 3921 1107
rect 3907 1056 3921 1060
rect 3919 1054 3921 1056
rect 3497 978 3509 984
rect 3569 978 3581 984
rect 3641 978 3653 984
rect 3707 978 3719 984
rect 3753 978 3765 984
rect 3811 978 3823 984
rect 3877 978 3889 992
rect 3937 978 3949 984
rect 4019 1060 4025 1107
rect 4036 1102 4045 1140
rect 4036 1072 4045 1090
rect 4116 1121 4124 1176
rect 4169 1156 4197 1160
rect 4209 1190 4237 1196
rect 4157 1154 4209 1156
rect 4137 1137 4153 1143
rect 4036 1066 4077 1072
rect 4019 1056 4033 1060
rect 4019 1054 4021 1056
rect 4071 1032 4077 1066
rect 4116 1024 4124 1107
rect 4137 1067 4143 1137
rect 4219 1146 4225 1156
rect 4196 1139 4225 1146
rect 4196 1113 4204 1139
rect 4300 1133 4307 1176
rect 4375 1142 4383 1156
rect 4403 1156 4431 1162
rect 4391 1153 4443 1156
rect 4474 1156 4500 1167
rect 4600 1176 4613 1182
rect 4600 1170 4607 1176
rect 4665 1164 4672 1176
rect 4375 1135 4400 1142
rect 4197 1064 4205 1099
rect 4300 1071 4307 1119
rect 4393 1113 4401 1135
rect 4474 1113 4482 1156
rect 4300 1064 4317 1071
rect 4399 1064 4407 1099
rect 4474 1064 4482 1099
rect 4561 1072 4567 1156
rect 4651 1157 4672 1164
rect 4722 1170 4729 1176
rect 4722 1162 4733 1170
rect 4619 1146 4626 1152
rect 4687 1146 4693 1148
rect 4619 1140 4693 1146
rect 4775 1141 4783 1156
rect 4809 1156 4837 1160
rect 4849 1190 4877 1196
rect 4797 1154 4849 1156
rect 4859 1146 4865 1156
rect 4619 1132 4626 1140
rect 4580 1124 4614 1132
rect 4580 1119 4586 1124
rect 4606 1106 4633 1113
rect 4561 1064 4623 1072
rect 4635 1068 4679 1074
rect 3991 978 4003 984
rect 4051 978 4063 992
rect 4097 978 4109 984
rect 4157 978 4169 984
rect 4227 978 4239 984
rect 4503 1058 4543 1064
rect 4531 1056 4543 1058
rect 4617 1050 4655 1058
rect 4673 1054 4679 1068
rect 4687 1068 4693 1140
rect 4767 1127 4783 1141
rect 4836 1139 4865 1146
rect 4753 1113 4767 1127
rect 4687 1062 4727 1068
rect 4747 1068 4761 1076
rect 4775 1064 4783 1127
rect 4836 1113 4844 1139
rect 4953 1133 4960 1176
rect 5015 1142 5023 1156
rect 5043 1156 5071 1162
rect 5177 1196 5189 1202
rect 5217 1196 5229 1202
rect 5257 1196 5269 1202
rect 5297 1196 5309 1202
rect 5369 1196 5381 1202
rect 5417 1196 5429 1202
rect 5457 1196 5469 1202
rect 5031 1153 5083 1156
rect 5015 1135 5040 1142
rect 4837 1064 4845 1099
rect 4953 1071 4960 1119
rect 5033 1113 5041 1135
rect 5133 1133 5140 1176
rect 5200 1133 5207 1176
rect 5280 1133 5287 1176
rect 5497 1196 5509 1202
rect 5537 1196 5549 1202
rect 5580 1196 5592 1202
rect 5630 1196 5642 1202
rect 4943 1064 4960 1071
rect 5039 1064 5047 1099
rect 5097 1067 5103 1133
rect 5133 1071 5140 1119
rect 4617 1044 4625 1050
rect 4673 1048 4703 1054
rect 4721 1044 4727 1062
rect 4607 1030 4625 1044
rect 4653 1030 4675 1042
rect 4617 1024 4625 1030
rect 4667 1024 4679 1030
rect 4721 1004 4733 1038
rect 4277 978 4289 984
rect 4376 978 4388 984
rect 4426 978 4438 984
rect 4511 978 4523 984
rect 4581 978 4593 984
rect 4647 978 4659 984
rect 4693 978 4705 984
rect 4751 978 4763 984
rect 4797 978 4809 984
rect 4867 978 4879 984
rect 4971 978 4983 984
rect 5123 1064 5140 1071
rect 5200 1071 5207 1119
rect 5280 1071 5287 1119
rect 5351 1113 5359 1156
rect 5391 1150 5399 1176
rect 5377 1144 5399 1150
rect 5377 1138 5380 1144
rect 5351 1099 5353 1113
rect 5200 1064 5217 1071
rect 5280 1064 5297 1071
rect 5351 1064 5359 1099
rect 5373 1082 5380 1138
rect 5440 1133 5447 1176
rect 5520 1133 5527 1176
rect 5677 1196 5685 1202
rect 5717 1196 5729 1202
rect 5791 1196 5803 1202
rect 5831 1196 5843 1202
rect 5877 1196 5889 1202
rect 6030 1196 6042 1202
rect 6077 1196 6089 1202
rect 6171 1196 6183 1202
rect 6211 1196 6223 1202
rect 5620 1156 5646 1167
rect 5547 1137 5563 1143
rect 5377 1076 5380 1082
rect 5377 1070 5403 1076
rect 5016 978 5028 984
rect 5066 978 5078 984
rect 5151 978 5163 984
rect 5395 1024 5403 1070
rect 5440 1071 5447 1119
rect 5520 1071 5527 1119
rect 5557 1083 5563 1137
rect 5638 1113 5646 1156
rect 5703 1148 5709 1176
rect 5703 1142 5713 1148
rect 5557 1077 5573 1083
rect 5440 1064 5457 1071
rect 5520 1064 5537 1071
rect 5638 1064 5646 1099
rect 5718 1081 5724 1136
rect 5740 1121 5747 1156
rect 5813 1133 5820 1176
rect 5869 1156 5897 1162
rect 5857 1153 5909 1156
rect 5917 1142 5925 1156
rect 5900 1135 5925 1142
rect 5976 1138 5994 1140
rect 5677 1072 5713 1080
rect 5677 1064 5685 1072
rect 5577 1058 5617 1064
rect 5577 1056 5589 1058
rect 5734 1063 5743 1107
rect 5813 1071 5820 1119
rect 5899 1113 5907 1135
rect 5976 1129 6006 1138
rect 6069 1156 6097 1162
rect 6057 1153 6109 1156
rect 6237 1196 6249 1202
rect 6277 1196 6289 1202
rect 6339 1196 6351 1202
rect 6397 1196 6409 1202
rect 6445 1196 6457 1202
rect 6507 1196 6519 1202
rect 6577 1196 6589 1202
rect 6117 1142 6125 1156
rect 6100 1135 6125 1142
rect 5927 1117 5943 1123
rect 5739 1054 5743 1063
rect 5803 1064 5820 1071
rect 5893 1064 5901 1099
rect 5937 1067 5943 1117
rect 5976 1101 5984 1129
rect 6099 1113 6107 1135
rect 6193 1133 6200 1176
rect 6260 1133 6267 1176
rect 6127 1117 6143 1123
rect 5177 978 5189 984
rect 5257 978 5269 984
rect 5369 978 5381 984
rect 5417 978 5429 984
rect 5497 978 5509 984
rect 5597 978 5609 984
rect 5707 978 5719 984
rect 5831 978 5843 984
rect 5975 1032 5982 1087
rect 6093 1064 6101 1099
rect 5975 1026 6022 1032
rect 5975 1024 5983 1026
rect 6011 1024 6022 1026
rect 5862 978 5874 984
rect 5912 978 5924 984
rect 5991 978 6003 984
rect 6031 978 6043 984
rect 6137 1043 6143 1117
rect 6193 1071 6200 1119
rect 6127 1037 6143 1043
rect 6183 1064 6200 1071
rect 6260 1071 6267 1119
rect 6487 1176 6500 1182
rect 6371 1170 6378 1176
rect 6367 1162 6378 1170
rect 6428 1164 6435 1176
rect 6493 1170 6500 1176
rect 6317 1141 6325 1156
rect 6428 1157 6449 1164
rect 6407 1146 6413 1148
rect 6474 1146 6481 1152
rect 6317 1127 6333 1141
rect 6407 1140 6481 1146
rect 6260 1064 6277 1071
rect 6062 978 6074 984
rect 6112 978 6124 984
rect 6211 978 6223 984
rect 6317 1064 6325 1127
rect 6333 1113 6347 1127
rect 6339 1068 6353 1076
rect 6407 1068 6413 1140
rect 6474 1132 6481 1140
rect 6486 1124 6520 1132
rect 6514 1119 6520 1124
rect 6467 1106 6494 1113
rect 6373 1062 6413 1068
rect 6421 1068 6465 1074
rect 6373 1044 6379 1062
rect 6421 1054 6427 1068
rect 6533 1072 6539 1156
rect 6569 1156 6597 1160
rect 6609 1190 6637 1196
rect 6557 1154 6609 1156
rect 6619 1146 6625 1156
rect 6596 1139 6625 1146
rect 6596 1113 6604 1139
rect 6477 1064 6539 1072
rect 6597 1064 6605 1099
rect 6397 1048 6427 1054
rect 6445 1050 6483 1058
rect 6475 1044 6483 1050
rect 6367 1004 6379 1038
rect 6425 1030 6447 1042
rect 6475 1030 6493 1044
rect 6421 1024 6433 1030
rect 6475 1024 6483 1030
rect 6237 978 6249 984
rect 6337 978 6349 984
rect 6395 978 6407 984
rect 6441 978 6453 984
rect 6507 978 6519 984
rect 6557 978 6569 984
rect 6627 978 6639 984
rect -62 976 6736 978
rect -62 964 4 976
rect -62 962 6736 964
rect -62 498 -2 962
rect 47 956 59 962
rect 131 956 143 962
rect 171 956 183 962
rect 217 956 229 962
rect 275 956 287 962
rect 321 956 333 962
rect 387 956 399 962
rect 471 956 483 962
rect 551 956 563 962
rect 79 877 83 886
rect 17 868 25 876
rect 17 860 53 868
rect 58 804 64 859
rect 74 833 83 877
rect 155 861 163 916
rect 247 902 259 936
rect 301 910 313 916
rect 355 910 363 916
rect 305 898 327 910
rect 355 896 373 910
rect 253 878 259 896
rect 277 886 307 892
rect 355 890 363 896
rect 43 792 53 798
rect 43 764 49 792
rect 80 784 87 819
rect 155 798 163 847
rect 139 792 163 798
rect 197 813 205 876
rect 219 864 233 872
rect 253 872 293 878
rect 213 813 227 827
rect 197 799 213 813
rect 287 800 293 872
rect 301 872 307 886
rect 325 882 363 890
rect 301 866 345 872
rect 357 868 419 876
rect 347 827 374 834
rect 394 816 400 821
rect 366 808 400 816
rect 354 800 361 808
rect 139 784 151 792
rect 197 784 205 799
rect 287 794 361 800
rect 287 792 293 794
rect 354 788 361 794
rect 247 770 258 778
rect 251 764 258 770
rect 308 776 329 783
rect 413 784 419 868
rect 456 833 464 916
rect 577 956 589 962
rect 657 956 669 962
rect 697 956 709 962
rect 737 956 749 962
rect 777 956 789 962
rect 837 956 849 962
rect 907 956 919 962
rect 523 869 540 876
rect 308 764 315 776
rect 373 764 380 770
rect 367 758 380 764
rect 456 764 464 819
rect 497 783 503 833
rect 487 777 503 783
rect 533 821 540 869
rect 600 869 617 876
rect 600 821 607 869
rect 677 861 685 916
rect 758 914 769 916
rect 797 914 805 916
rect 758 908 805 914
rect 707 877 723 883
rect 533 764 540 807
rect 600 764 607 807
rect 677 798 685 847
rect 717 823 723 877
rect 798 853 805 908
rect 962 956 974 962
rect 1012 956 1024 962
rect 877 841 885 876
rect 1062 956 1074 962
rect 1112 956 1124 962
rect 1291 956 1303 962
rect 1342 956 1354 962
rect 1392 956 1404 962
rect 1471 956 1483 962
rect 1521 956 1533 962
rect 1587 956 1599 962
rect 1633 956 1645 962
rect 1691 956 1703 962
rect 1737 956 1749 962
rect 1167 950 1219 956
rect 1167 948 1179 950
rect 1207 948 1219 950
rect 1191 876 1199 892
rect 1243 950 1271 956
rect 1251 892 1263 896
rect 1219 888 1263 892
rect 1207 886 1263 888
rect 1271 890 1283 896
rect 1311 890 1323 896
rect 1271 884 1323 890
rect 717 817 733 823
rect 796 811 804 839
rect 677 792 701 798
rect 689 784 701 792
rect 17 738 25 744
rect 57 738 69 744
rect 169 738 181 744
rect 219 738 231 744
rect 277 738 289 744
rect 325 738 337 744
rect 387 738 399 744
rect 471 738 483 744
rect 511 738 523 744
rect 551 738 563 744
rect 577 738 589 744
rect 617 738 629 744
rect 774 802 804 811
rect 786 800 804 802
rect 876 801 884 827
rect 937 803 943 873
rect 993 841 1001 876
rect 1093 841 1101 876
rect 1191 868 1214 876
rect 876 794 905 801
rect 937 797 953 803
rect 837 784 889 786
rect 899 784 905 794
rect 999 805 1007 827
rect 1027 817 1043 823
rect 1206 833 1214 868
rect 1373 841 1381 876
rect 1000 798 1025 805
rect 957 784 1009 787
rect 849 780 877 784
rect 889 744 917 750
rect 969 778 997 784
rect 1017 784 1025 798
rect 1037 803 1043 817
rect 1037 797 1053 803
rect 1099 805 1107 827
rect 1127 817 1153 823
rect 1207 819 1214 833
rect 1456 833 1464 916
rect 1557 910 1565 916
rect 1607 910 1619 916
rect 1547 896 1565 910
rect 1593 898 1615 910
rect 1661 902 1673 936
rect 1557 890 1565 896
rect 1557 882 1595 890
rect 1613 886 1643 892
rect 1501 868 1563 876
rect 1100 798 1125 805
rect 1057 784 1109 787
rect 1069 778 1097 784
rect 1117 784 1125 798
rect 1206 776 1214 819
rect 1379 805 1387 827
rect 1380 798 1405 805
rect 1337 784 1389 787
rect 1206 770 1278 776
rect 1231 764 1238 770
rect 1271 764 1278 770
rect 1349 778 1377 784
rect 1397 784 1405 798
rect 1456 764 1464 819
rect 1501 784 1507 868
rect 1613 872 1619 886
rect 1661 878 1667 896
rect 1575 866 1619 872
rect 1627 872 1667 878
rect 1546 827 1573 834
rect 1520 816 1526 821
rect 1520 808 1554 816
rect 1559 800 1566 808
rect 1627 800 1633 872
rect 1817 948 1829 962
rect 1877 956 1889 962
rect 1687 864 1701 872
rect 1693 813 1707 827
rect 1715 813 1723 876
rect 1756 833 1764 916
rect 1803 874 1809 908
rect 1859 884 1861 886
rect 1847 880 1861 884
rect 1803 868 1844 874
rect 1559 794 1633 800
rect 1707 799 1723 813
rect 1835 850 1844 868
rect 1559 788 1566 794
rect 1627 792 1633 794
rect 1591 776 1612 783
rect 1715 784 1723 799
rect 1540 764 1547 770
rect 1605 764 1612 776
rect 1662 770 1673 778
rect 1662 764 1669 770
rect 1540 758 1553 764
rect 1756 764 1764 819
rect 1835 800 1844 838
rect 1855 833 1861 880
rect 1922 956 1934 962
rect 1972 956 1984 962
rect 2017 956 2029 962
rect 2057 956 2069 962
rect 2117 956 2129 962
rect 2175 956 2187 962
rect 2221 956 2233 962
rect 2287 956 2299 962
rect 2337 956 2349 962
rect 2397 956 2409 962
rect 2467 956 2479 962
rect 1953 841 1961 876
rect 2037 861 2045 916
rect 2147 902 2159 936
rect 2201 910 2213 916
rect 2255 910 2263 916
rect 2205 898 2227 910
rect 2255 896 2273 910
rect 2153 878 2159 896
rect 2177 886 2207 892
rect 2255 890 2263 896
rect 1802 794 1844 800
rect 1802 772 1809 794
rect 1855 788 1861 819
rect 1959 805 1967 827
rect 1960 798 1985 805
rect 1847 784 1861 788
rect 1859 782 1861 784
rect 659 738 671 744
rect 738 738 750 744
rect 857 738 869 744
rect 977 738 989 744
rect 1077 738 1089 744
rect 1251 738 1263 744
rect 1291 738 1305 744
rect 1357 738 1369 744
rect 1471 738 1483 744
rect 1521 738 1533 744
rect 1583 738 1595 744
rect 1631 738 1643 744
rect 1689 738 1701 744
rect 1737 738 1749 744
rect 1817 738 1829 752
rect 1877 738 1889 752
rect 1917 784 1969 787
rect 1929 778 1957 784
rect 1977 784 1985 798
rect 2037 798 2045 847
rect 2097 813 2105 876
rect 2119 864 2133 872
rect 2153 872 2193 878
rect 2113 813 2127 827
rect 2097 799 2113 813
rect 2187 800 2193 872
rect 2201 872 2207 886
rect 2225 882 2263 890
rect 2201 866 2245 872
rect 2257 868 2319 876
rect 2247 827 2274 834
rect 2294 816 2300 821
rect 2266 808 2300 816
rect 2254 800 2261 808
rect 2037 792 2061 798
rect 2049 784 2061 792
rect 2097 784 2105 799
rect 2187 794 2261 800
rect 2187 792 2193 794
rect 2254 788 2261 794
rect 2147 770 2158 778
rect 2151 764 2158 770
rect 2208 776 2229 783
rect 2313 784 2319 868
rect 2356 833 2364 916
rect 2517 956 2529 962
rect 2616 956 2628 962
rect 2666 956 2678 962
rect 2711 956 2723 962
rect 2751 956 2763 962
rect 2791 956 2803 962
rect 2831 956 2843 962
rect 2871 956 2883 962
rect 2917 956 2929 962
rect 3051 956 3063 962
rect 3111 956 3123 962
rect 2897 882 2909 884
rect 2897 876 2937 882
rect 3071 882 3083 884
rect 3043 876 3083 882
rect 3171 948 3183 962
rect 3231 956 3243 962
rect 3139 884 3141 886
rect 3139 880 3153 884
rect 2208 764 2215 776
rect 2273 764 2280 770
rect 2267 758 2280 764
rect 2356 764 2364 819
rect 2377 803 2383 853
rect 2437 841 2445 876
rect 2540 869 2557 876
rect 2377 797 2393 803
rect 2436 801 2444 827
rect 2540 821 2547 869
rect 2639 841 2647 876
rect 2731 870 2743 876
rect 2771 870 2783 876
rect 2811 870 2823 876
rect 2851 870 2863 876
rect 2725 862 2743 870
rect 2758 862 2783 870
rect 2798 862 2823 870
rect 2837 862 2863 870
rect 2436 794 2465 801
rect 2397 784 2449 786
rect 2459 784 2465 794
rect 2409 780 2437 784
rect 2449 744 2477 750
rect 2540 764 2547 807
rect 2633 805 2641 827
rect 2725 833 2732 862
rect 2727 819 2732 833
rect 2615 798 2640 805
rect 2725 798 2732 819
rect 2758 816 2766 862
rect 2798 816 2806 862
rect 2837 816 2845 862
rect 2887 857 2933 863
rect 2958 841 2966 876
rect 3014 841 3022 876
rect 2750 804 2766 816
rect 2790 804 2806 816
rect 2830 804 2845 816
rect 2758 798 2766 804
rect 2798 798 2806 804
rect 2837 798 2845 804
rect 2615 784 2623 798
rect 2725 791 2744 798
rect 2726 790 2744 791
rect 2758 790 2784 798
rect 2798 790 2823 798
rect 2837 790 2864 798
rect 2631 784 2683 787
rect 2732 784 2744 790
rect 2772 784 2784 790
rect 2811 784 2823 790
rect 2852 784 2864 790
rect 2958 784 2966 827
rect 2643 778 2671 784
rect 1937 738 1949 744
rect 2019 738 2031 744
rect 2119 738 2131 744
rect 2177 738 2189 744
rect 2225 738 2237 744
rect 2287 738 2299 744
rect 2337 738 2349 744
rect 2417 738 2429 744
rect 2517 738 2529 744
rect 2557 738 2569 744
rect 2651 738 2663 744
rect 2711 738 2723 744
rect 2751 738 2763 744
rect 2791 738 2803 744
rect 2831 738 2843 744
rect 2871 738 2883 744
rect 2940 773 2966 784
rect 3014 784 3022 827
rect 3139 833 3145 880
rect 3191 874 3197 908
rect 3291 948 3303 962
rect 3356 956 3368 962
rect 3406 956 3418 962
rect 3259 884 3261 886
rect 3259 880 3273 884
rect 3156 868 3197 874
rect 3156 850 3165 868
rect 3014 773 3040 784
rect 2900 738 2912 744
rect 2950 738 2962 744
rect 3018 738 3030 744
rect 3068 738 3080 744
rect 3139 788 3145 819
rect 3156 800 3165 838
rect 3259 833 3265 880
rect 3311 874 3317 908
rect 3437 956 3449 962
rect 3477 956 3489 962
rect 3537 948 3549 962
rect 3597 956 3609 962
rect 3671 956 3683 962
rect 3276 868 3317 874
rect 3276 850 3285 868
rect 3156 794 3198 800
rect 3139 784 3153 788
rect 3139 782 3141 784
rect 3191 772 3198 794
rect 3259 788 3265 819
rect 3276 800 3285 838
rect 3379 841 3387 876
rect 3457 861 3465 916
rect 3523 874 3529 908
rect 3579 884 3581 886
rect 3567 880 3581 884
rect 3523 868 3564 874
rect 3373 805 3381 827
rect 3276 794 3318 800
rect 3259 784 3273 788
rect 3259 782 3261 784
rect 3311 772 3318 794
rect 3355 798 3380 805
rect 3457 798 3465 847
rect 3555 850 3564 868
rect 3555 800 3564 838
rect 3575 833 3581 880
rect 3711 956 3723 962
rect 3656 833 3664 916
rect 3771 948 3783 962
rect 3841 956 3853 962
rect 3907 956 3919 962
rect 3953 956 3965 962
rect 4011 956 4023 962
rect 3739 884 3741 886
rect 3739 880 3753 884
rect 3739 833 3745 880
rect 3791 874 3797 908
rect 3756 868 3797 874
rect 3877 910 3885 916
rect 3927 910 3939 916
rect 3867 896 3885 910
rect 3913 898 3935 910
rect 3981 902 3993 936
rect 3877 890 3885 896
rect 3877 882 3915 890
rect 3933 886 3963 892
rect 3821 868 3883 876
rect 3756 850 3765 868
rect 3355 784 3363 798
rect 3457 792 3481 798
rect 3111 738 3123 752
rect 3171 738 3183 752
rect 3231 738 3243 752
rect 3291 738 3303 752
rect 3371 784 3423 787
rect 3469 784 3481 792
rect 3383 778 3411 784
rect 3522 794 3564 800
rect 3522 772 3529 794
rect 3575 788 3581 819
rect 3567 784 3581 788
rect 3579 782 3581 784
rect 3656 764 3664 819
rect 3391 738 3403 744
rect 3439 738 3451 744
rect 3537 738 3549 752
rect 3597 738 3609 752
rect 3671 738 3683 744
rect 3739 788 3745 819
rect 3756 800 3765 838
rect 3756 794 3798 800
rect 3739 784 3753 788
rect 3739 782 3741 784
rect 3791 772 3798 794
rect 3821 784 3827 868
rect 3933 872 3939 886
rect 3981 878 3987 896
rect 3895 866 3939 872
rect 3947 872 3987 878
rect 3866 827 3893 834
rect 3840 816 3846 821
rect 3840 808 3874 816
rect 3879 800 3886 808
rect 3947 800 3953 872
rect 4077 948 4089 962
rect 4137 956 4149 962
rect 4197 956 4209 962
rect 4282 956 4294 962
rect 4332 956 4344 962
rect 4411 956 4423 962
rect 4451 956 4463 962
rect 4007 864 4021 872
rect 4013 813 4027 827
rect 4035 813 4043 876
rect 4063 874 4069 908
rect 4119 884 4121 886
rect 4107 880 4121 884
rect 4063 868 4104 874
rect 4095 850 4104 868
rect 3879 794 3953 800
rect 4027 799 4043 813
rect 4095 800 4104 838
rect 4115 833 4121 880
rect 4177 882 4189 884
rect 4177 876 4217 882
rect 4395 914 4403 916
rect 4477 956 4489 962
rect 4542 956 4554 962
rect 4592 956 4604 962
rect 4431 914 4442 916
rect 4395 908 4442 914
rect 4167 857 4213 863
rect 4238 841 4246 876
rect 3879 788 3886 794
rect 3947 792 3953 794
rect 3711 738 3723 752
rect 3771 738 3783 752
rect 3911 776 3932 783
rect 4035 784 4043 799
rect 3860 764 3867 770
rect 3925 764 3932 776
rect 3982 770 3993 778
rect 3982 764 3989 770
rect 3860 758 3873 764
rect 4062 794 4104 800
rect 4062 772 4069 794
rect 4115 788 4121 819
rect 4107 784 4121 788
rect 4119 782 4121 784
rect 4238 784 4246 827
rect 4257 803 4263 853
rect 4313 841 4321 876
rect 4395 853 4402 908
rect 4257 797 4273 803
rect 4319 805 4327 827
rect 4396 811 4404 839
rect 4496 833 4504 916
rect 4637 956 4649 962
rect 4677 956 4689 962
rect 4751 956 4763 962
rect 4782 956 4794 962
rect 4832 956 4844 962
rect 4573 841 4581 876
rect 4320 798 4345 805
rect 4396 802 4426 811
rect 4396 800 4414 802
rect 3841 738 3853 744
rect 3903 738 3915 744
rect 3951 738 3963 744
rect 4009 738 4021 744
rect 4077 738 4089 752
rect 4137 738 4149 752
rect 4220 773 4246 784
rect 4277 784 4329 787
rect 4289 778 4317 784
rect 4337 784 4345 798
rect 4496 764 4504 819
rect 4579 805 4587 827
rect 4617 823 4623 873
rect 4657 861 4665 916
rect 4607 817 4623 823
rect 4580 798 4605 805
rect 4537 784 4589 787
rect 4180 738 4192 744
rect 4230 738 4242 744
rect 4297 738 4309 744
rect 4450 738 4462 744
rect 4549 778 4577 784
rect 4597 784 4605 798
rect 4657 798 4665 847
rect 4736 833 4744 916
rect 4877 956 4889 962
rect 4917 956 4929 962
rect 4977 948 4989 962
rect 5037 956 5049 962
rect 4857 877 4873 883
rect 4813 841 4821 876
rect 4657 792 4681 798
rect 4669 784 4681 792
rect 4736 764 4744 819
rect 4819 805 4827 827
rect 4857 823 4863 877
rect 4897 861 4905 916
rect 4963 874 4969 908
rect 5019 884 5021 886
rect 5007 880 5021 884
rect 4963 868 5004 874
rect 4847 817 4863 823
rect 4820 798 4845 805
rect 4777 784 4829 787
rect 4789 778 4817 784
rect 4837 784 4845 798
rect 4897 798 4905 847
rect 4995 850 5004 868
rect 4995 800 5004 838
rect 5015 833 5021 880
rect 5091 956 5103 962
rect 5151 948 5163 962
rect 5197 956 5209 962
rect 5237 956 5249 962
rect 5277 956 5289 962
rect 5317 956 5329 962
rect 5357 956 5369 962
rect 5417 956 5429 962
rect 5531 956 5543 962
rect 5119 884 5121 886
rect 5119 880 5133 884
rect 5119 833 5125 880
rect 5171 874 5177 908
rect 5397 882 5409 884
rect 5397 876 5437 882
rect 5562 956 5574 962
rect 5612 956 5624 962
rect 5136 868 5177 874
rect 5217 870 5229 876
rect 5257 870 5269 876
rect 5297 870 5309 876
rect 5337 870 5349 876
rect 5136 850 5145 868
rect 5217 862 5243 870
rect 5257 862 5282 870
rect 5297 862 5322 870
rect 5337 862 5355 870
rect 4897 792 4921 798
rect 4909 784 4921 792
rect 4962 794 5004 800
rect 4962 772 4969 794
rect 5015 788 5021 819
rect 5007 784 5021 788
rect 5019 782 5021 784
rect 4477 738 4489 744
rect 4557 738 4569 744
rect 4639 738 4651 744
rect 4751 738 4763 744
rect 4797 738 4809 744
rect 4879 738 4891 744
rect 4977 738 4989 752
rect 5037 738 5049 752
rect 5119 788 5125 819
rect 5136 800 5145 838
rect 5235 816 5243 862
rect 5274 816 5282 862
rect 5314 816 5322 862
rect 5348 833 5355 862
rect 5458 841 5466 876
rect 5348 819 5353 833
rect 5235 804 5250 816
rect 5274 804 5290 816
rect 5314 804 5330 816
rect 5136 794 5178 800
rect 5235 798 5243 804
rect 5274 798 5282 804
rect 5314 798 5322 804
rect 5348 798 5355 819
rect 5516 833 5524 916
rect 5657 956 5669 962
rect 5697 956 5709 962
rect 5742 956 5754 962
rect 5792 956 5804 962
rect 5871 956 5883 962
rect 5911 956 5923 962
rect 5961 956 5973 962
rect 6027 956 6039 962
rect 6073 956 6085 962
rect 6131 956 6143 962
rect 6182 956 6194 962
rect 6232 956 6244 962
rect 5593 841 5601 876
rect 5677 861 5685 916
rect 5855 914 5863 916
rect 5891 914 5902 916
rect 5855 908 5902 914
rect 5119 784 5133 788
rect 5119 782 5121 784
rect 5171 772 5178 794
rect 5216 790 5243 798
rect 5257 790 5282 798
rect 5296 790 5322 798
rect 5336 791 5355 798
rect 5336 790 5354 791
rect 5216 784 5228 790
rect 5257 784 5269 790
rect 5296 784 5308 790
rect 5336 784 5348 790
rect 5458 784 5466 827
rect 5091 738 5103 752
rect 5151 738 5163 752
rect 5197 738 5209 744
rect 5237 738 5249 744
rect 5277 738 5289 744
rect 5317 738 5329 744
rect 5357 738 5369 744
rect 5440 773 5466 784
rect 5516 764 5524 819
rect 5599 805 5607 827
rect 5600 798 5625 805
rect 5557 784 5609 787
rect 5569 778 5597 784
rect 5617 784 5625 798
rect 5677 798 5685 847
rect 5773 841 5781 876
rect 5855 853 5862 908
rect 5997 910 6005 916
rect 6047 910 6059 916
rect 5987 896 6005 910
rect 6033 898 6055 910
rect 6101 902 6113 936
rect 5997 890 6005 896
rect 5997 882 6035 890
rect 6053 886 6083 892
rect 5941 868 6003 876
rect 5779 805 5787 827
rect 5856 811 5864 839
rect 5780 798 5805 805
rect 5856 802 5886 811
rect 5856 800 5874 802
rect 5677 792 5701 798
rect 5689 784 5701 792
rect 5737 784 5789 787
rect 5749 778 5777 784
rect 5797 784 5805 798
rect 5941 784 5947 868
rect 6053 872 6059 886
rect 6101 878 6107 896
rect 6015 866 6059 872
rect 6067 872 6107 878
rect 5986 827 6013 834
rect 5960 816 5966 821
rect 5960 808 5994 816
rect 5999 800 6006 808
rect 6067 800 6073 872
rect 6282 956 6294 962
rect 6332 956 6344 962
rect 6391 956 6403 962
rect 6431 956 6443 962
rect 6481 956 6493 962
rect 6547 956 6559 962
rect 6593 956 6605 962
rect 6651 956 6663 962
rect 6127 864 6141 872
rect 6133 813 6147 827
rect 6155 813 6163 876
rect 6213 841 6221 876
rect 6313 841 6321 876
rect 6415 861 6423 916
rect 6517 910 6525 916
rect 6567 910 6579 916
rect 6507 896 6525 910
rect 6553 898 6575 910
rect 6621 902 6633 936
rect 6517 890 6525 896
rect 6517 882 6555 890
rect 6573 886 6603 892
rect 6461 868 6523 876
rect 5999 794 6073 800
rect 6147 799 6163 813
rect 6219 805 6227 827
rect 6319 805 6327 827
rect 5999 788 6006 794
rect 6067 792 6073 794
rect 6031 776 6052 783
rect 6155 784 6163 799
rect 6220 798 6245 805
rect 6320 798 6345 805
rect 6415 798 6423 847
rect 5980 764 5987 770
rect 6045 764 6052 776
rect 6102 770 6113 778
rect 6102 764 6109 770
rect 5980 758 5993 764
rect 6177 784 6229 787
rect 6189 778 6217 784
rect 6237 784 6245 798
rect 6277 784 6329 787
rect 6289 778 6317 784
rect 6337 784 6345 798
rect 6399 792 6423 798
rect 6399 784 6411 792
rect 6461 784 6467 868
rect 6573 872 6579 886
rect 6621 878 6627 896
rect 6535 866 6579 872
rect 6587 872 6627 878
rect 6506 827 6533 834
rect 6480 816 6486 821
rect 6480 808 6514 816
rect 6519 800 6526 808
rect 6587 800 6593 872
rect 6647 864 6661 872
rect 6653 813 6667 827
rect 6675 813 6683 876
rect 6519 794 6593 800
rect 6667 799 6683 813
rect 6519 788 6526 794
rect 6587 792 6593 794
rect 6551 776 6572 783
rect 6675 784 6683 799
rect 6500 764 6507 770
rect 6565 764 6572 776
rect 6622 770 6633 778
rect 6622 764 6629 770
rect 6500 758 6513 764
rect 5400 738 5412 744
rect 5450 738 5462 744
rect 5531 738 5543 744
rect 5577 738 5589 744
rect 5659 738 5671 744
rect 5757 738 5769 744
rect 5910 738 5922 744
rect 5961 738 5973 744
rect 6023 738 6035 744
rect 6071 738 6083 744
rect 6129 738 6141 744
rect 6197 738 6209 744
rect 6297 738 6309 744
rect 6429 738 6441 744
rect 6481 738 6493 744
rect 6543 738 6555 744
rect 6591 738 6603 744
rect 6649 738 6661 744
rect 6742 738 6802 1202
rect 4 736 6802 738
rect 6736 724 6802 736
rect 4 722 6802 724
rect 17 716 29 722
rect 79 716 91 722
rect 160 716 172 722
rect 210 716 222 722
rect 36 641 44 696
rect 257 716 269 722
rect 338 716 350 722
rect 388 716 400 722
rect 200 676 226 687
rect 109 668 121 676
rect 97 662 121 668
rect 36 544 44 627
rect 97 613 105 662
rect 218 633 226 676
rect 276 641 284 696
rect 334 676 360 687
rect 418 716 430 722
rect 569 716 581 722
rect 670 716 682 722
rect 334 633 342 676
rect 539 668 551 676
rect 539 662 563 668
rect 466 658 484 660
rect 97 544 105 599
rect 218 584 226 619
rect 157 578 197 584
rect 157 576 169 578
rect 276 544 284 627
rect 454 649 484 658
rect 476 621 484 649
rect 334 584 342 619
rect 555 613 563 662
rect 616 658 634 660
rect 616 649 646 658
rect 697 716 709 722
rect 757 716 769 722
rect 831 716 843 722
rect 871 716 883 722
rect 991 716 1003 722
rect 1031 716 1045 722
rect 1101 716 1113 722
rect 1163 716 1175 722
rect 1211 716 1223 722
rect 1269 716 1281 722
rect 1339 716 1351 722
rect 1399 716 1411 722
rect 1501 716 1513 722
rect 1563 716 1575 722
rect 1611 716 1623 722
rect 1669 716 1681 722
rect 1741 716 1753 722
rect 1803 716 1815 722
rect 1851 716 1863 722
rect 1909 716 1921 722
rect 1981 716 1993 722
rect 2043 716 2055 722
rect 2091 716 2103 722
rect 2149 716 2161 722
rect 2221 716 2233 722
rect 2283 716 2295 722
rect 2331 716 2343 722
rect 2389 716 2401 722
rect 2459 716 2471 722
rect 2517 716 2529 722
rect 2565 716 2577 722
rect 2627 716 2639 722
rect 2712 716 2724 722
rect 2768 716 2780 722
rect 2831 716 2843 722
rect 616 621 624 649
rect 716 641 724 696
rect 776 641 784 696
rect 853 653 860 696
rect 971 690 978 696
rect 1011 690 1018 696
rect 946 684 1018 690
rect 946 641 954 684
rect 1120 696 1133 702
rect 1120 690 1127 696
rect 1185 684 1192 696
rect 363 578 403 584
rect 391 576 403 578
rect 478 552 485 607
rect 438 546 485 552
rect 438 544 449 546
rect 477 544 485 546
rect 555 544 563 599
rect 615 552 622 607
rect 615 546 662 552
rect 615 544 623 546
rect 651 544 662 546
rect 716 544 724 627
rect 776 544 784 627
rect 853 591 860 639
rect 947 627 954 641
rect 946 592 954 627
rect 843 584 860 591
rect 931 584 954 592
rect 1081 592 1087 676
rect 1171 677 1192 684
rect 1242 690 1249 696
rect 1242 682 1253 690
rect 1139 666 1146 672
rect 1207 666 1213 668
rect 1139 660 1213 666
rect 1295 661 1303 676
rect 1321 670 1329 696
rect 1321 664 1343 670
rect 1139 652 1146 660
rect 1100 644 1134 652
rect 1100 639 1106 644
rect 1126 626 1153 633
rect 1081 584 1143 592
rect 1155 588 1199 594
rect 17 498 29 504
rect 77 498 89 504
rect 117 498 129 504
rect 177 498 189 504
rect 257 498 269 504
rect 371 498 383 504
rect 417 498 429 504
rect 457 498 469 504
rect 531 498 543 504
rect 571 498 583 504
rect 631 498 643 504
rect 671 498 683 504
rect 931 568 939 584
rect 947 572 1003 574
rect 907 510 919 512
rect 959 568 1003 572
rect 991 564 1003 568
rect 947 510 959 512
rect 907 504 959 510
rect 1011 570 1063 576
rect 1011 564 1023 570
rect 1051 564 1063 570
rect 983 504 1011 510
rect 1137 570 1175 578
rect 1193 574 1199 588
rect 1207 588 1213 660
rect 1287 647 1303 661
rect 1273 633 1287 647
rect 1207 582 1247 588
rect 1267 588 1281 596
rect 1295 584 1303 647
rect 1340 658 1343 664
rect 1340 602 1347 658
rect 1361 633 1369 676
rect 1429 668 1441 676
rect 1417 662 1441 668
rect 1520 696 1533 702
rect 1520 690 1527 696
rect 1585 684 1592 696
rect 1367 619 1369 633
rect 1340 596 1343 602
rect 1137 564 1145 570
rect 1193 568 1223 574
rect 1241 564 1247 582
rect 1127 550 1145 564
rect 1173 550 1195 562
rect 1137 544 1145 550
rect 1187 544 1199 550
rect 1241 524 1253 558
rect 1317 590 1343 596
rect 1317 544 1325 590
rect 1361 584 1369 619
rect 1417 613 1425 662
rect 1417 544 1425 599
rect 1481 592 1487 676
rect 1571 677 1592 684
rect 1642 690 1649 696
rect 1642 682 1653 690
rect 1539 666 1546 672
rect 1607 666 1613 668
rect 1539 660 1613 666
rect 1695 661 1703 676
rect 1539 652 1546 660
rect 1500 644 1534 652
rect 1500 639 1506 644
rect 1526 626 1553 633
rect 1481 584 1543 592
rect 1555 588 1599 594
rect 1537 570 1575 578
rect 1593 574 1599 588
rect 1607 588 1613 660
rect 1687 647 1703 661
rect 1673 633 1687 647
rect 1607 582 1647 588
rect 1667 588 1681 596
rect 1695 584 1703 647
rect 1537 564 1545 570
rect 1593 568 1623 574
rect 1641 564 1647 582
rect 1527 550 1545 564
rect 1573 550 1595 562
rect 1537 544 1545 550
rect 1587 544 1599 550
rect 1641 524 1653 558
rect 1760 696 1773 702
rect 1760 690 1767 696
rect 1825 684 1832 696
rect 1721 592 1727 676
rect 1811 677 1832 684
rect 1882 690 1889 696
rect 1882 682 1893 690
rect 1779 666 1786 672
rect 1847 666 1853 668
rect 1779 660 1853 666
rect 1935 661 1943 676
rect 1779 652 1786 660
rect 1740 644 1774 652
rect 1740 639 1746 644
rect 1766 626 1793 633
rect 1721 584 1783 592
rect 1795 588 1839 594
rect 1777 570 1815 578
rect 1833 574 1839 588
rect 1847 588 1853 660
rect 1927 647 1943 661
rect 1913 633 1927 647
rect 1847 582 1887 588
rect 1907 588 1921 596
rect 1935 584 1943 647
rect 1777 564 1785 570
rect 1833 568 1863 574
rect 1881 564 1887 582
rect 1767 550 1785 564
rect 1813 550 1835 562
rect 1777 544 1785 550
rect 1827 544 1839 550
rect 1881 524 1893 558
rect 2000 696 2013 702
rect 2000 690 2007 696
rect 2065 684 2072 696
rect 1961 592 1967 676
rect 2051 677 2072 684
rect 2122 690 2129 696
rect 2122 682 2133 690
rect 2019 666 2026 672
rect 2087 666 2093 668
rect 2019 660 2093 666
rect 2175 661 2183 676
rect 2019 652 2026 660
rect 1980 644 2014 652
rect 1980 639 1986 644
rect 2006 626 2033 633
rect 1961 584 2023 592
rect 2035 588 2079 594
rect 2017 570 2055 578
rect 2073 574 2079 588
rect 2087 588 2093 660
rect 2167 647 2183 661
rect 2153 633 2167 647
rect 2087 582 2127 588
rect 2147 588 2161 596
rect 2175 584 2183 647
rect 2017 564 2025 570
rect 2073 568 2103 574
rect 2121 564 2127 582
rect 2007 550 2025 564
rect 2053 550 2075 562
rect 2017 544 2025 550
rect 2067 544 2079 550
rect 2121 524 2133 558
rect 2240 696 2253 702
rect 2240 690 2247 696
rect 2305 684 2312 696
rect 2201 592 2207 676
rect 2291 677 2312 684
rect 2362 690 2369 696
rect 2362 682 2373 690
rect 2259 666 2266 672
rect 2327 666 2333 668
rect 2259 660 2333 666
rect 2415 661 2423 676
rect 2259 652 2266 660
rect 2220 644 2254 652
rect 2220 639 2226 644
rect 2246 626 2273 633
rect 2201 584 2263 592
rect 2275 588 2319 594
rect 2257 570 2295 578
rect 2313 574 2319 588
rect 2327 588 2333 660
rect 2407 647 2423 661
rect 2393 633 2407 647
rect 2327 582 2367 588
rect 2387 588 2401 596
rect 2415 584 2423 647
rect 2257 564 2265 570
rect 2313 568 2343 574
rect 2361 564 2367 582
rect 2247 550 2265 564
rect 2293 550 2315 562
rect 2257 544 2265 550
rect 2307 544 2319 550
rect 2361 524 2373 558
rect 2607 696 2620 702
rect 2491 690 2498 696
rect 2487 682 2498 690
rect 2548 684 2555 696
rect 2613 690 2620 696
rect 2437 661 2445 676
rect 2548 677 2569 684
rect 2878 716 2890 722
rect 2928 716 2940 722
rect 2527 666 2533 668
rect 2594 666 2601 672
rect 2437 647 2453 661
rect 2527 660 2601 666
rect 2437 584 2445 647
rect 2453 633 2467 647
rect 2459 588 2473 596
rect 2527 588 2533 660
rect 2594 652 2601 660
rect 2606 644 2640 652
rect 2634 639 2640 644
rect 2587 626 2614 633
rect 2493 582 2533 588
rect 2541 588 2585 594
rect 2493 564 2499 582
rect 2541 574 2547 588
rect 2653 592 2659 676
rect 2740 633 2747 676
rect 2816 641 2824 696
rect 2874 676 2900 687
rect 2957 716 2969 722
rect 3037 716 3049 722
rect 3119 716 3131 722
rect 3198 716 3210 722
rect 3297 716 3309 722
rect 3377 716 3389 722
rect 3459 716 3471 722
rect 3540 716 3552 722
rect 3590 716 3602 722
rect 2874 633 2882 676
rect 2733 596 2739 619
rect 2597 584 2659 592
rect 2712 590 2739 596
rect 2712 584 2724 590
rect 2517 568 2547 574
rect 2565 570 2603 578
rect 2595 564 2603 570
rect 2487 524 2499 558
rect 2545 550 2567 562
rect 2595 550 2613 564
rect 2541 544 2553 550
rect 2595 544 2603 550
rect 2703 504 2731 510
rect 2743 576 2771 582
rect 2816 544 2824 627
rect 2976 641 2984 696
rect 3029 676 3057 682
rect 3017 673 3069 676
rect 2874 584 2882 619
rect 2903 578 2943 584
rect 2931 576 2943 578
rect 2976 544 2984 627
rect 2997 587 3003 673
rect 3077 662 3085 676
rect 3149 668 3161 676
rect 3060 655 3085 662
rect 3097 657 3113 663
rect 3059 633 3067 655
rect 3097 643 3103 657
rect 3137 662 3161 668
rect 3087 637 3103 643
rect 3053 584 3061 619
rect 3137 613 3145 662
rect 3246 658 3264 660
rect 3234 649 3264 658
rect 3177 637 3193 643
rect 3137 544 3145 599
rect 3177 587 3183 637
rect 3256 621 3264 649
rect 3316 641 3324 696
rect 3369 676 3397 682
rect 3357 673 3409 676
rect 3637 716 3649 722
rect 3677 716 3689 722
rect 3737 716 3749 722
rect 3890 716 3902 722
rect 3939 716 3951 722
rect 3997 716 4009 722
rect 4045 716 4057 722
rect 4107 716 4119 722
rect 4171 716 4183 722
rect 4211 716 4223 722
rect 4259 716 4271 722
rect 4317 716 4329 722
rect 4365 716 4377 722
rect 4427 716 4439 722
rect 4477 716 4489 722
rect 4540 716 4552 722
rect 4596 716 4608 722
rect 3580 676 3606 687
rect 3417 662 3425 676
rect 3489 668 3501 676
rect 3400 655 3425 662
rect 3477 662 3501 668
rect 3258 552 3265 607
rect 3218 546 3265 552
rect 3218 544 3229 546
rect 697 498 709 504
rect 757 498 769 504
rect 871 498 883 504
rect 1031 498 1043 504
rect 1101 498 1113 504
rect 1167 498 1179 504
rect 1213 498 1225 504
rect 1271 498 1283 504
rect 1339 498 1351 504
rect 1397 498 1409 504
rect 1437 498 1449 504
rect 1501 498 1513 504
rect 1567 498 1579 504
rect 1613 498 1625 504
rect 1671 498 1683 504
rect 1741 498 1753 504
rect 1807 498 1819 504
rect 1853 498 1865 504
rect 1911 498 1923 504
rect 1981 498 1993 504
rect 2047 498 2059 504
rect 2093 498 2105 504
rect 2151 498 2163 504
rect 2221 498 2233 504
rect 2287 498 2299 504
rect 2333 498 2345 504
rect 2391 498 2403 504
rect 2457 498 2469 504
rect 2515 498 2527 504
rect 2561 498 2573 504
rect 2627 498 2639 504
rect 2751 498 2763 504
rect 2831 498 2843 504
rect 2911 498 2923 504
rect 2957 498 2969 504
rect 3022 498 3034 504
rect 3072 498 3084 504
rect 3117 498 3129 504
rect 3157 498 3169 504
rect 3257 544 3265 546
rect 3316 544 3324 627
rect 3399 633 3407 655
rect 3393 584 3401 619
rect 3477 613 3485 662
rect 3598 633 3606 676
rect 3660 653 3667 696
rect 3729 676 3757 682
rect 3717 673 3769 676
rect 3777 662 3785 676
rect 3760 655 3785 662
rect 3477 544 3485 599
rect 3598 584 3606 619
rect 3660 591 3667 639
rect 3759 633 3767 655
rect 3817 643 3823 693
rect 3787 637 3823 643
rect 3836 658 3854 660
rect 3836 649 3866 658
rect 4087 696 4100 702
rect 3971 690 3978 696
rect 3967 682 3978 690
rect 4028 684 4035 696
rect 4093 690 4100 696
rect 3917 661 3925 676
rect 4028 677 4049 684
rect 4007 666 4013 668
rect 4074 666 4081 672
rect 3836 621 3844 649
rect 3917 647 3933 661
rect 4007 660 4081 666
rect 3660 584 3677 591
rect 3753 584 3761 619
rect 3537 578 3577 584
rect 3537 576 3549 578
rect 3197 498 3209 504
rect 3237 498 3249 504
rect 3297 498 3309 504
rect 3362 498 3374 504
rect 3412 498 3424 504
rect 3835 552 3842 607
rect 3917 584 3925 647
rect 3933 633 3947 647
rect 3939 588 3953 596
rect 3835 546 3882 552
rect 3835 544 3843 546
rect 3871 544 3882 546
rect 4007 588 4013 660
rect 4074 652 4081 660
rect 4086 644 4120 652
rect 4114 639 4120 644
rect 4067 626 4094 633
rect 3973 582 4013 588
rect 4021 588 4065 594
rect 3973 564 3979 582
rect 4021 574 4027 588
rect 4133 592 4139 676
rect 4193 653 4200 696
rect 4407 696 4420 702
rect 4291 690 4298 696
rect 4287 682 4298 690
rect 4348 684 4355 696
rect 4413 690 4420 696
rect 4237 661 4245 676
rect 4348 677 4369 684
rect 4327 666 4333 668
rect 4394 666 4401 672
rect 4237 647 4253 661
rect 4327 660 4401 666
rect 4077 584 4139 592
rect 4193 591 4200 639
rect 3997 568 4027 574
rect 4045 570 4083 578
rect 4075 564 4083 570
rect 3967 524 3979 558
rect 4025 550 4047 562
rect 4075 550 4093 564
rect 4021 544 4033 550
rect 4075 544 4083 550
rect 4183 584 4200 591
rect 4237 584 4245 647
rect 4253 633 4267 647
rect 4259 588 4273 596
rect 4327 588 4333 660
rect 4394 652 4401 660
rect 4406 644 4440 652
rect 4434 639 4440 644
rect 4387 626 4414 633
rect 4293 582 4333 588
rect 4341 588 4385 594
rect 4293 564 4299 582
rect 4341 574 4347 588
rect 4453 592 4459 676
rect 4496 641 4504 696
rect 4678 716 4690 722
rect 4728 716 4740 722
rect 4811 716 4823 722
rect 4859 716 4871 722
rect 4971 716 4983 722
rect 4674 676 4700 687
rect 4397 584 4459 592
rect 4317 568 4347 574
rect 4365 570 4403 578
rect 4395 564 4403 570
rect 4287 524 4299 558
rect 4345 550 4367 562
rect 4395 550 4413 564
rect 4341 544 4353 550
rect 4395 544 4403 550
rect 4496 544 4504 627
rect 4573 633 4580 676
rect 4674 633 4682 676
rect 4775 662 4783 676
rect 4803 676 4831 682
rect 5011 708 5023 722
rect 5071 708 5083 722
rect 5118 716 5130 722
rect 5239 716 5251 722
rect 5297 716 5309 722
rect 5345 716 5357 722
rect 5407 716 5419 722
rect 5457 716 5469 722
rect 4791 673 4843 676
rect 4889 668 4901 676
rect 4877 662 4901 668
rect 4775 655 4800 662
rect 4757 637 4773 643
rect 4581 596 4587 619
rect 4581 590 4608 596
rect 4596 584 4608 590
rect 4674 584 4682 619
rect 4757 587 4763 637
rect 4793 633 4801 655
rect 4549 576 4577 582
rect 4589 504 4617 510
rect 4703 578 4743 584
rect 4731 576 4743 578
rect 4799 584 4807 619
rect 4877 613 4885 662
rect 4956 641 4964 696
rect 5039 676 5041 678
rect 5039 672 5053 676
rect 5039 641 5045 672
rect 5091 666 5098 688
rect 5056 660 5098 666
rect 4877 544 4885 599
rect 4956 544 4964 627
rect 3457 498 3469 504
rect 3497 498 3509 504
rect 3557 498 3569 504
rect 3637 498 3649 504
rect 3722 498 3734 504
rect 3772 498 3784 504
rect 3851 498 3863 504
rect 3891 498 3903 504
rect 3937 498 3949 504
rect 3995 498 4007 504
rect 4041 498 4053 504
rect 4107 498 4119 504
rect 4211 498 4223 504
rect 4257 498 4269 504
rect 4315 498 4327 504
rect 4361 498 4373 504
rect 4427 498 4439 504
rect 4477 498 4489 504
rect 4557 498 4569 504
rect 4711 498 4723 504
rect 4776 498 4788 504
rect 4826 498 4838 504
rect 4857 498 4869 504
rect 4897 498 4909 504
rect 4971 498 4983 504
rect 5039 580 5045 627
rect 5056 622 5065 660
rect 5387 696 5400 702
rect 5271 690 5278 696
rect 5267 682 5278 690
rect 5328 684 5335 696
rect 5393 690 5400 696
rect 5217 661 5225 676
rect 5328 677 5349 684
rect 5537 708 5549 722
rect 5597 708 5609 722
rect 5307 666 5313 668
rect 5374 666 5381 672
rect 5166 658 5184 660
rect 5154 649 5184 658
rect 5056 592 5065 610
rect 5176 621 5184 649
rect 5217 647 5233 661
rect 5307 660 5381 666
rect 5056 586 5097 592
rect 5039 576 5053 580
rect 5039 574 5041 576
rect 5091 552 5097 586
rect 5178 552 5185 607
rect 5138 546 5185 552
rect 5138 544 5149 546
rect 5011 498 5023 504
rect 5071 498 5083 512
rect 5177 544 5185 546
rect 5217 584 5225 647
rect 5233 633 5247 647
rect 5239 588 5253 596
rect 5307 588 5313 660
rect 5374 652 5381 660
rect 5386 644 5420 652
rect 5414 639 5420 644
rect 5367 626 5394 633
rect 5273 582 5313 588
rect 5321 588 5365 594
rect 5273 564 5279 582
rect 5321 574 5327 588
rect 5433 592 5439 676
rect 5476 633 5484 676
rect 5522 666 5529 688
rect 5579 676 5581 678
rect 5567 672 5581 676
rect 5522 660 5564 666
rect 5377 584 5439 592
rect 5476 584 5484 619
rect 5555 622 5564 660
rect 5575 641 5581 672
rect 5651 716 5663 722
rect 5691 716 5703 722
rect 5731 716 5743 722
rect 5771 716 5783 722
rect 5811 716 5823 722
rect 5851 716 5863 722
rect 5877 716 5889 722
rect 5917 716 5929 722
rect 5971 716 5983 722
rect 6011 716 6023 722
rect 6057 716 6069 722
rect 6157 716 6169 722
rect 6289 716 6301 722
rect 6341 716 6353 722
rect 6403 716 6415 722
rect 6451 716 6463 722
rect 6509 716 6521 722
rect 6557 716 6569 722
rect 6617 716 6629 722
rect 5673 653 5680 696
rect 5707 657 5723 663
rect 5555 592 5564 610
rect 5523 586 5564 592
rect 5297 568 5327 574
rect 5345 570 5383 578
rect 5375 564 5383 570
rect 5267 524 5279 558
rect 5325 550 5347 562
rect 5375 550 5393 564
rect 5321 544 5333 550
rect 5375 544 5383 550
rect 5523 552 5529 586
rect 5575 580 5581 627
rect 5673 591 5680 639
rect 5717 607 5723 657
rect 5753 653 5760 696
rect 5833 653 5840 696
rect 5900 653 5907 696
rect 5927 657 5943 663
rect 5753 591 5760 639
rect 5833 591 5840 639
rect 5663 584 5680 591
rect 5743 584 5760 591
rect 5823 584 5840 591
rect 5900 591 5907 639
rect 5937 603 5943 657
rect 5993 653 6000 696
rect 6049 676 6077 682
rect 6037 673 6089 676
rect 6149 676 6177 682
rect 6097 662 6105 676
rect 6137 673 6189 676
rect 6360 696 6373 702
rect 6360 690 6367 696
rect 6425 684 6432 696
rect 6197 662 6205 676
rect 6259 668 6271 676
rect 6259 662 6283 668
rect 6080 655 6105 662
rect 6180 655 6205 662
rect 5937 597 5953 603
rect 5993 591 6000 639
rect 6079 633 6087 655
rect 6179 633 6187 655
rect 5900 584 5917 591
rect 5567 576 5581 580
rect 5579 574 5581 576
rect 5117 498 5129 504
rect 5157 498 5169 504
rect 5237 498 5249 504
rect 5295 498 5307 504
rect 5341 498 5353 504
rect 5407 498 5419 504
rect 5457 498 5469 504
rect 5537 498 5549 512
rect 5597 498 5609 504
rect 5691 498 5703 504
rect 5771 498 5783 504
rect 5851 498 5863 504
rect 5983 584 6000 591
rect 6073 584 6081 619
rect 6173 584 6181 619
rect 6275 613 6283 662
rect 5877 498 5889 504
rect 6011 498 6023 504
rect 6042 498 6054 504
rect 6092 498 6104 504
rect 6275 544 6283 599
rect 6321 592 6327 676
rect 6411 677 6432 684
rect 6482 690 6489 696
rect 6482 682 6493 690
rect 6379 666 6386 672
rect 6447 666 6453 668
rect 6379 660 6453 666
rect 6535 661 6543 676
rect 6379 652 6386 660
rect 6340 644 6374 652
rect 6340 639 6346 644
rect 6366 626 6393 633
rect 6321 584 6383 592
rect 6395 588 6439 594
rect 6142 498 6154 504
rect 6192 498 6204 504
rect 6377 570 6415 578
rect 6433 574 6439 588
rect 6447 588 6453 660
rect 6527 647 6543 661
rect 6513 633 6527 647
rect 6447 582 6487 588
rect 6507 588 6521 596
rect 6535 584 6543 647
rect 6576 641 6584 696
rect 6636 641 6644 696
rect 6377 564 6385 570
rect 6433 568 6463 574
rect 6481 564 6487 582
rect 6367 550 6385 564
rect 6413 550 6435 562
rect 6377 544 6385 550
rect 6427 544 6439 550
rect 6481 524 6493 558
rect 6576 544 6584 627
rect 6636 544 6644 627
rect 6251 498 6263 504
rect 6291 498 6303 504
rect 6341 498 6353 504
rect 6407 498 6419 504
rect 6453 498 6465 504
rect 6511 498 6523 504
rect 6557 498 6569 504
rect 6617 498 6629 504
rect -62 496 6736 498
rect -62 484 4 496
rect -62 482 6736 484
rect -62 18 -2 482
rect 37 476 49 482
rect 95 476 107 482
rect 141 476 153 482
rect 207 476 219 482
rect 281 476 293 482
rect 347 476 359 482
rect 393 476 405 482
rect 451 476 463 482
rect 497 476 509 482
rect 537 476 549 482
rect 597 476 609 482
rect 731 476 743 482
rect 67 422 79 456
rect 121 430 133 436
rect 175 430 183 436
rect 125 418 147 430
rect 175 416 193 430
rect 73 398 79 416
rect 97 406 127 412
rect 175 410 183 416
rect 17 333 25 396
rect 39 384 53 392
rect 73 392 113 398
rect 33 333 47 347
rect 17 319 33 333
rect 107 320 113 392
rect 121 392 127 406
rect 145 402 183 410
rect 121 386 165 392
rect 177 388 239 396
rect 167 347 194 354
rect 214 336 220 341
rect 186 328 220 336
rect 174 320 181 328
rect 17 304 25 319
rect 107 314 181 320
rect 107 312 113 314
rect 174 308 181 314
rect 67 290 78 298
rect 71 284 78 290
rect 128 296 149 303
rect 233 304 239 388
rect 128 284 135 296
rect 193 284 200 290
rect 187 278 200 284
rect 317 430 325 436
rect 367 430 379 436
rect 307 416 325 430
rect 353 418 375 430
rect 421 422 433 456
rect 317 410 325 416
rect 317 402 355 410
rect 373 406 403 412
rect 261 388 323 396
rect 261 304 267 388
rect 373 392 379 406
rect 421 398 427 416
rect 335 386 379 392
rect 387 392 427 398
rect 306 347 333 354
rect 280 336 286 341
rect 280 328 314 336
rect 319 320 326 328
rect 387 320 393 392
rect 518 434 529 436
rect 557 434 565 436
rect 518 428 565 434
rect 447 384 461 392
rect 453 333 467 347
rect 475 333 483 396
rect 558 373 565 428
rect 319 314 393 320
rect 467 319 483 333
rect 556 331 564 359
rect 319 308 326 314
rect 387 312 393 314
rect 351 296 372 303
rect 475 304 483 319
rect 300 284 307 290
rect 365 284 372 296
rect 422 290 433 298
rect 422 284 429 290
rect 300 278 313 284
rect 534 322 564 331
rect 546 320 564 322
rect 577 323 583 393
rect 620 389 637 396
rect 757 476 769 482
rect 797 476 809 482
rect 871 476 883 482
rect 921 476 933 482
rect 987 476 999 482
rect 1033 476 1045 482
rect 1091 476 1103 482
rect 1169 476 1181 482
rect 1239 476 1251 482
rect 1319 476 1331 482
rect 1411 476 1423 482
rect 703 389 720 396
rect 620 341 627 389
rect 577 317 593 323
rect 620 284 627 327
rect 713 341 720 389
rect 777 381 785 436
rect 713 284 720 327
rect 777 318 785 367
rect 856 353 864 436
rect 957 430 965 436
rect 1007 430 1019 436
rect 947 416 965 430
rect 993 418 1015 430
rect 1061 422 1073 456
rect 957 410 965 416
rect 957 402 995 410
rect 1013 406 1043 412
rect 901 388 963 396
rect 777 312 801 318
rect 789 304 801 312
rect 39 258 51 264
rect 97 258 109 264
rect 145 258 157 264
rect 207 258 219 264
rect 281 258 293 264
rect 343 258 355 264
rect 391 258 403 264
rect 449 258 461 264
rect 498 258 510 264
rect 597 258 609 264
rect 637 258 649 264
rect 691 258 703 264
rect 731 258 743 264
rect 856 284 864 339
rect 901 304 907 388
rect 1013 392 1019 406
rect 1061 398 1067 416
rect 975 386 1019 392
rect 1027 392 1067 398
rect 946 347 973 354
rect 920 336 926 341
rect 920 328 954 336
rect 959 320 966 328
rect 1027 320 1033 392
rect 1087 384 1101 392
rect 1093 333 1107 347
rect 1115 333 1123 396
rect 959 314 1033 320
rect 1107 319 1123 333
rect 959 308 966 314
rect 1027 312 1033 314
rect 991 296 1012 303
rect 1115 304 1123 319
rect 1151 361 1159 396
rect 1195 390 1203 436
rect 1177 384 1203 390
rect 1217 390 1225 436
rect 1217 384 1243 390
rect 1177 378 1180 384
rect 1151 347 1153 361
rect 1151 304 1159 347
rect 1173 322 1180 378
rect 1240 378 1243 384
rect 1177 316 1180 322
rect 1240 322 1247 378
rect 1261 361 1269 396
rect 1297 390 1305 436
rect 1442 476 1454 482
rect 1492 476 1504 482
rect 1571 476 1583 482
rect 1297 384 1323 390
rect 1320 378 1323 384
rect 1267 347 1269 361
rect 1240 316 1243 322
rect 1177 310 1199 316
rect 940 284 947 290
rect 1005 284 1012 296
rect 1062 290 1073 298
rect 1062 284 1069 290
rect 940 278 953 284
rect 1191 284 1199 310
rect 1221 310 1243 316
rect 1221 284 1229 310
rect 1261 304 1269 347
rect 1320 322 1327 378
rect 1341 361 1349 396
rect 1347 347 1349 361
rect 1396 353 1404 436
rect 1602 476 1614 482
rect 1652 476 1664 482
rect 1721 476 1733 482
rect 1787 476 1799 482
rect 1833 476 1845 482
rect 1891 476 1903 482
rect 1971 476 1983 482
rect 2031 476 2043 482
rect 1473 361 1481 396
rect 1320 316 1323 322
rect 1301 310 1323 316
rect 1301 284 1309 310
rect 1341 304 1349 347
rect 1396 284 1404 339
rect 1556 353 1564 436
rect 1757 430 1765 436
rect 1807 430 1819 436
rect 1747 416 1765 430
rect 1793 418 1815 430
rect 1861 422 1873 456
rect 1757 410 1765 416
rect 1757 402 1795 410
rect 1813 406 1843 412
rect 1633 361 1641 396
rect 1701 388 1763 396
rect 1479 325 1487 347
rect 1480 318 1505 325
rect 1437 304 1489 307
rect 1449 298 1477 304
rect 1497 304 1505 318
rect 1556 284 1564 339
rect 1639 325 1647 347
rect 1640 318 1665 325
rect 1597 304 1649 307
rect 1609 298 1637 304
rect 1657 304 1665 318
rect 1701 304 1707 388
rect 1813 392 1819 406
rect 1861 398 1867 416
rect 1775 386 1819 392
rect 1827 392 1867 398
rect 1746 347 1773 354
rect 1720 336 1726 341
rect 1720 328 1754 336
rect 1759 320 1766 328
rect 1827 320 1833 392
rect 2062 476 2074 482
rect 2112 476 2124 482
rect 1887 384 1901 392
rect 1893 333 1907 347
rect 1915 333 1923 396
rect 1956 353 1964 436
rect 2016 353 2024 436
rect 2157 476 2169 482
rect 2217 476 2229 482
rect 2287 476 2299 482
rect 2093 361 2101 396
rect 1759 314 1833 320
rect 1907 319 1923 333
rect 1759 308 1766 314
rect 1827 312 1833 314
rect 1791 296 1812 303
rect 1915 304 1923 319
rect 1740 284 1747 290
rect 1805 284 1812 296
rect 1862 290 1873 298
rect 1862 284 1869 290
rect 1740 278 1753 284
rect 1956 284 1964 339
rect 2016 284 2024 339
rect 2176 353 2184 436
rect 2356 476 2368 482
rect 2406 476 2418 482
rect 2437 476 2449 482
rect 2541 476 2553 482
rect 2607 476 2619 482
rect 2653 476 2665 482
rect 2711 476 2723 482
rect 2776 476 2788 482
rect 2826 476 2838 482
rect 2099 325 2107 347
rect 2100 318 2125 325
rect 2057 304 2109 307
rect 2069 298 2097 304
rect 2117 304 2125 318
rect 2176 284 2184 339
rect 2197 307 2203 373
rect 2257 361 2265 396
rect 2256 321 2264 347
rect 2379 361 2387 396
rect 2460 389 2477 396
rect 2577 430 2585 436
rect 2627 430 2639 436
rect 2567 416 2585 430
rect 2613 418 2635 430
rect 2681 422 2693 456
rect 2577 410 2585 416
rect 2577 402 2615 410
rect 2633 406 2663 412
rect 2256 314 2285 321
rect 2217 304 2269 306
rect 2279 304 2285 314
rect 2337 323 2343 353
rect 2373 325 2381 347
rect 2460 341 2467 389
rect 2521 388 2583 396
rect 2307 317 2343 323
rect 2355 318 2380 325
rect 2355 304 2363 318
rect 2229 300 2257 304
rect 2269 264 2297 270
rect 2371 304 2423 307
rect 2383 298 2411 304
rect 2460 284 2467 327
rect 2521 304 2527 388
rect 2633 392 2639 406
rect 2681 398 2687 416
rect 2595 386 2639 392
rect 2647 392 2687 398
rect 2566 347 2593 354
rect 2540 336 2546 341
rect 2540 328 2574 336
rect 2579 320 2586 328
rect 2647 320 2653 392
rect 2857 476 2869 482
rect 2961 476 2973 482
rect 3027 476 3039 482
rect 3073 476 3085 482
rect 3131 476 3143 482
rect 3177 476 3189 482
rect 3217 476 3229 482
rect 2707 384 2721 392
rect 2713 333 2727 347
rect 2735 333 2743 396
rect 2799 361 2807 396
rect 2880 389 2897 396
rect 2997 430 3005 436
rect 3047 430 3059 436
rect 2987 416 3005 430
rect 3033 418 3055 430
rect 3101 422 3113 456
rect 2997 410 3005 416
rect 2997 402 3035 410
rect 3053 406 3083 412
rect 2579 314 2653 320
rect 2727 319 2743 333
rect 2793 325 2801 347
rect 2880 341 2887 389
rect 2941 388 3003 396
rect 2579 308 2586 314
rect 2647 312 2653 314
rect 2611 296 2632 303
rect 2735 304 2743 319
rect 2775 318 2800 325
rect 2775 304 2783 318
rect 2560 284 2567 290
rect 2625 284 2632 296
rect 2682 290 2693 298
rect 2682 284 2689 290
rect 2560 278 2573 284
rect 2791 304 2843 307
rect 2803 298 2831 304
rect 2880 284 2887 327
rect 2941 304 2947 388
rect 3053 392 3059 406
rect 3101 398 3107 416
rect 3015 386 3059 392
rect 3067 392 3107 398
rect 2986 347 3013 354
rect 2960 336 2966 341
rect 2960 328 2994 336
rect 2999 320 3006 328
rect 3067 320 3073 392
rect 3276 476 3288 482
rect 3326 476 3338 482
rect 3127 384 3141 392
rect 3133 333 3147 347
rect 3155 333 3163 396
rect 3197 381 3205 436
rect 3357 476 3369 482
rect 3491 476 3503 482
rect 3542 476 3554 482
rect 3592 476 3604 482
rect 3511 402 3523 404
rect 3483 396 3523 402
rect 3637 476 3649 482
rect 3737 476 3749 482
rect 3871 476 3883 482
rect 3717 402 3729 404
rect 3717 396 3757 402
rect 3902 476 3914 482
rect 3952 476 3964 482
rect 4031 476 4043 482
rect 4071 476 4083 482
rect 4015 434 4023 436
rect 4097 476 4109 482
rect 4197 476 4209 482
rect 4255 476 4267 482
rect 4301 476 4313 482
rect 4367 476 4379 482
rect 4417 476 4429 482
rect 4516 476 4528 482
rect 4566 476 4578 482
rect 4051 434 4062 436
rect 4015 428 4062 434
rect 2999 314 3073 320
rect 3147 319 3163 333
rect 2999 308 3006 314
rect 3067 312 3073 314
rect 3031 296 3052 303
rect 3155 304 3163 319
rect 3197 318 3205 367
rect 3299 361 3307 396
rect 3380 389 3397 396
rect 3293 325 3301 347
rect 3380 341 3387 389
rect 3454 361 3462 396
rect 3573 361 3581 396
rect 3660 389 3677 396
rect 3275 318 3300 325
rect 3197 312 3221 318
rect 3209 304 3221 312
rect 3275 304 3283 318
rect 2980 284 2987 290
rect 3045 284 3052 296
rect 3102 290 3113 298
rect 3102 284 3109 290
rect 2980 278 2993 284
rect 3291 304 3343 307
rect 3303 298 3331 304
rect 3380 284 3387 327
rect 3454 304 3462 347
rect 3579 325 3587 347
rect 3660 341 3667 389
rect 3697 377 3713 383
rect 3580 318 3605 325
rect 3537 304 3589 307
rect 3454 293 3480 304
rect 759 258 771 264
rect 871 258 883 264
rect 921 258 933 264
rect 983 258 995 264
rect 1031 258 1043 264
rect 1089 258 1101 264
rect 1169 258 1181 264
rect 1239 258 1251 264
rect 1319 258 1331 264
rect 1411 258 1423 264
rect 1457 258 1469 264
rect 1571 258 1583 264
rect 1617 258 1629 264
rect 1721 258 1733 264
rect 1783 258 1795 264
rect 1831 258 1843 264
rect 1889 258 1901 264
rect 1971 258 1983 264
rect 2031 258 2043 264
rect 2077 258 2089 264
rect 2157 258 2169 264
rect 2237 258 2249 264
rect 2391 258 2403 264
rect 2437 258 2449 264
rect 2477 258 2489 264
rect 2541 258 2553 264
rect 2603 258 2615 264
rect 2651 258 2663 264
rect 2709 258 2721 264
rect 2811 258 2823 264
rect 2857 258 2869 264
rect 2897 258 2909 264
rect 2961 258 2973 264
rect 3023 258 3035 264
rect 3071 258 3083 264
rect 3129 258 3141 264
rect 3179 258 3191 264
rect 3311 258 3323 264
rect 3357 258 3369 264
rect 3397 258 3409 264
rect 3549 298 3577 304
rect 3597 304 3605 318
rect 3660 284 3667 327
rect 3697 323 3703 377
rect 3778 361 3786 396
rect 3843 389 3860 396
rect 3687 317 3703 323
rect 3778 304 3786 347
rect 3458 258 3470 264
rect 3508 258 3520 264
rect 3557 258 3569 264
rect 3637 258 3649 264
rect 3677 258 3689 264
rect 3760 293 3786 304
rect 3853 341 3860 389
rect 3933 361 3941 396
rect 4015 373 4022 428
rect 4120 389 4137 396
rect 4227 422 4239 456
rect 4281 430 4293 436
rect 4335 430 4343 436
rect 4285 418 4307 430
rect 4335 416 4353 430
rect 4233 398 4239 416
rect 4257 406 4287 412
rect 4335 410 4343 416
rect 3853 284 3860 327
rect 3939 325 3947 347
rect 4016 331 4024 359
rect 4120 341 4127 389
rect 3940 318 3965 325
rect 4016 322 4046 331
rect 4016 320 4034 322
rect 3897 304 3949 307
rect 3720 258 3732 264
rect 3770 258 3782 264
rect 3909 298 3937 304
rect 3957 304 3965 318
rect 4120 284 4127 327
rect 4157 323 4163 393
rect 4147 317 4163 323
rect 4177 333 4185 396
rect 4199 384 4213 392
rect 4233 392 4273 398
rect 4193 333 4207 347
rect 4177 319 4193 333
rect 4267 320 4273 392
rect 4281 392 4287 406
rect 4305 402 4343 410
rect 4597 476 4609 482
rect 4701 476 4713 482
rect 4771 476 4783 482
rect 4831 476 4843 482
rect 4881 476 4893 482
rect 4947 476 4959 482
rect 4993 476 5005 482
rect 5051 476 5063 482
rect 5151 476 5163 482
rect 5197 476 5209 482
rect 5296 476 5308 482
rect 5346 476 5358 482
rect 4281 386 4325 392
rect 4337 388 4399 396
rect 4327 347 4354 354
rect 4374 336 4380 341
rect 4346 328 4380 336
rect 4334 320 4341 328
rect 4177 304 4185 319
rect 4267 314 4341 320
rect 4267 312 4273 314
rect 3831 258 3843 264
rect 3871 258 3883 264
rect 3917 258 3929 264
rect 4070 258 4082 264
rect 4334 308 4341 314
rect 4227 290 4238 298
rect 4231 284 4238 290
rect 4288 296 4309 303
rect 4393 304 4399 388
rect 4440 389 4457 396
rect 4440 341 4447 389
rect 4539 361 4547 396
rect 4620 389 4637 396
rect 4288 284 4295 296
rect 4353 284 4360 290
rect 4347 278 4360 284
rect 4440 284 4447 327
rect 4533 325 4541 347
rect 4620 341 4627 389
rect 4735 361 4743 396
rect 4515 318 4540 325
rect 4515 304 4523 318
rect 4531 304 4583 307
rect 4543 298 4571 304
rect 4620 284 4627 327
rect 4736 321 4744 347
rect 4816 353 4824 436
rect 4917 430 4925 436
rect 4967 430 4979 436
rect 4907 416 4925 430
rect 4953 418 4975 430
rect 5021 422 5033 456
rect 4917 410 4925 416
rect 4917 402 4955 410
rect 4973 406 5003 412
rect 4861 388 4923 396
rect 4715 314 4744 321
rect 4715 304 4721 314
rect 4731 304 4783 306
rect 4703 264 4731 270
rect 4743 300 4771 304
rect 4816 284 4824 339
rect 4861 304 4867 388
rect 4973 392 4979 406
rect 5021 398 5027 416
rect 4935 386 4979 392
rect 4987 392 5027 398
rect 4906 347 4933 354
rect 4880 336 4886 341
rect 4880 328 4914 336
rect 4919 320 4926 328
rect 4987 320 4993 392
rect 5171 402 5183 404
rect 5143 396 5183 402
rect 5377 476 5389 482
rect 5477 476 5489 482
rect 5557 476 5569 482
rect 5597 476 5609 482
rect 5662 476 5674 482
rect 5712 476 5724 482
rect 5457 402 5469 404
rect 5457 396 5497 402
rect 5578 434 5589 436
rect 5617 434 5625 436
rect 5578 428 5625 434
rect 5047 384 5061 392
rect 5053 333 5067 347
rect 5075 333 5083 396
rect 5114 361 5122 396
rect 5220 389 5237 396
rect 4919 314 4993 320
rect 5067 319 5083 333
rect 4919 308 4926 314
rect 4987 312 4993 314
rect 4951 296 4972 303
rect 5075 304 5083 319
rect 4900 284 4907 290
rect 4965 284 4972 296
rect 5022 290 5033 298
rect 5022 284 5029 290
rect 4900 278 4913 284
rect 5114 304 5122 347
rect 5220 341 5227 389
rect 5114 293 5140 304
rect 5220 284 5227 327
rect 5257 323 5263 373
rect 5319 361 5327 396
rect 5400 389 5417 396
rect 5313 325 5321 347
rect 5400 341 5407 389
rect 5518 361 5526 396
rect 5618 373 5625 428
rect 5771 476 5783 482
rect 5811 476 5823 482
rect 5856 476 5868 482
rect 5906 476 5918 482
rect 5693 361 5701 396
rect 5795 381 5803 436
rect 5942 476 5954 482
rect 5992 476 6004 482
rect 6042 476 6054 482
rect 6092 476 6104 482
rect 6191 476 6203 482
rect 6271 476 6283 482
rect 5247 317 5263 323
rect 5295 318 5320 325
rect 5295 304 5303 318
rect 4097 258 4109 264
rect 4137 258 4149 264
rect 4199 258 4211 264
rect 4257 258 4269 264
rect 4305 258 4317 264
rect 4367 258 4379 264
rect 4417 258 4429 264
rect 4457 258 4469 264
rect 4551 258 4563 264
rect 4597 258 4609 264
rect 4637 258 4649 264
rect 4751 258 4763 264
rect 4831 258 4843 264
rect 4881 258 4893 264
rect 4943 258 4955 264
rect 4991 258 5003 264
rect 5049 258 5061 264
rect 5118 258 5130 264
rect 5168 258 5180 264
rect 5311 304 5363 307
rect 5323 298 5351 304
rect 5400 284 5407 327
rect 5518 304 5526 347
rect 5616 331 5624 359
rect 5197 258 5209 264
rect 5237 258 5249 264
rect 5331 258 5343 264
rect 5377 258 5389 264
rect 5417 258 5429 264
rect 5500 293 5526 304
rect 5460 258 5472 264
rect 5510 258 5522 264
rect 5594 322 5624 331
rect 5699 325 5707 347
rect 5606 320 5624 322
rect 5700 318 5725 325
rect 5795 318 5803 367
rect 5879 361 5887 396
rect 5973 361 5981 396
rect 6073 361 6081 396
rect 6321 476 6333 482
rect 6391 476 6403 482
rect 6441 476 6453 482
rect 6507 476 6519 482
rect 6553 476 6565 482
rect 6611 476 6623 482
rect 5873 325 5881 347
rect 5979 325 5987 347
rect 6079 325 6087 347
rect 5657 304 5709 307
rect 5669 298 5697 304
rect 5717 304 5725 318
rect 5779 312 5803 318
rect 5855 318 5880 325
rect 5980 318 6005 325
rect 6080 318 6105 325
rect 5779 304 5791 312
rect 5855 304 5863 318
rect 5871 304 5923 307
rect 5883 298 5911 304
rect 5937 304 5989 307
rect 5949 298 5977 304
rect 5997 304 6005 318
rect 6037 304 6089 307
rect 6049 298 6077 304
rect 6097 304 6105 318
rect 6137 323 6143 393
rect 6163 389 6180 396
rect 6243 389 6260 396
rect 6477 430 6485 436
rect 6527 430 6539 436
rect 6467 416 6485 430
rect 6513 418 6535 430
rect 6581 422 6593 456
rect 6477 410 6485 416
rect 6477 402 6515 410
rect 6533 406 6563 412
rect 6173 341 6180 389
rect 6253 341 6260 389
rect 6297 327 6303 393
rect 6355 361 6363 396
rect 6421 388 6483 396
rect 6137 317 6153 323
rect 6173 284 6180 327
rect 6253 284 6260 327
rect 6356 321 6364 347
rect 6335 314 6364 321
rect 6335 304 6341 314
rect 6351 304 6403 306
rect 5558 258 5570 264
rect 5677 258 5689 264
rect 5809 258 5821 264
rect 5891 258 5903 264
rect 5957 258 5969 264
rect 6057 258 6069 264
rect 6151 258 6163 264
rect 6191 258 6203 264
rect 6323 264 6351 270
rect 6363 300 6391 304
rect 6421 304 6427 388
rect 6533 392 6539 406
rect 6581 398 6587 416
rect 6495 386 6539 392
rect 6547 392 6587 398
rect 6466 347 6493 354
rect 6440 336 6446 341
rect 6440 328 6474 336
rect 6479 320 6486 328
rect 6547 320 6553 392
rect 6607 384 6621 392
rect 6613 333 6627 347
rect 6635 333 6643 396
rect 6479 314 6553 320
rect 6627 319 6643 333
rect 6479 308 6486 314
rect 6547 312 6553 314
rect 6511 296 6532 303
rect 6635 304 6643 319
rect 6460 284 6467 290
rect 6525 284 6532 296
rect 6582 290 6593 298
rect 6582 284 6589 290
rect 6460 278 6473 284
rect 6231 258 6243 264
rect 6271 258 6283 264
rect 6371 258 6383 264
rect 6441 258 6453 264
rect 6503 258 6515 264
rect 6551 258 6563 264
rect 6609 258 6621 264
rect 6742 258 6802 722
rect 4 256 6802 258
rect 6736 244 6802 256
rect 4 242 6802 244
rect 39 236 51 242
rect 97 236 109 242
rect 145 236 157 242
rect 207 236 219 242
rect 279 236 291 242
rect 337 236 349 242
rect 385 236 397 242
rect 447 236 459 242
rect 529 236 541 242
rect 599 236 611 242
rect 689 236 701 242
rect 759 236 771 242
rect 817 236 829 242
rect 865 236 877 242
rect 927 236 939 242
rect 999 236 1011 242
rect 1109 236 1121 242
rect 1191 236 1203 242
rect 1261 236 1273 242
rect 1323 236 1335 242
rect 1371 236 1383 242
rect 1429 236 1441 242
rect 1511 236 1523 242
rect 187 216 200 222
rect 71 210 78 216
rect 67 202 78 210
rect 128 204 135 216
rect 193 210 200 216
rect 17 181 25 196
rect 128 197 149 204
rect 107 186 113 188
rect 174 186 181 192
rect 17 167 33 181
rect 107 180 181 186
rect 17 104 25 167
rect 33 153 47 167
rect 39 108 53 116
rect 107 108 113 180
rect 174 172 181 180
rect 186 164 220 172
rect 214 159 220 164
rect 167 146 194 153
rect 73 102 113 108
rect 121 108 165 114
rect 73 84 79 102
rect 121 94 127 108
rect 233 112 239 196
rect 177 104 239 112
rect 97 88 127 94
rect 145 90 183 98
rect 175 84 183 90
rect 67 44 79 78
rect 125 70 147 82
rect 175 70 193 84
rect 121 64 133 70
rect 175 64 183 70
rect 427 216 440 222
rect 311 210 318 216
rect 307 202 318 210
rect 368 204 375 216
rect 433 210 440 216
rect 257 181 265 196
rect 368 197 389 204
rect 347 186 353 188
rect 414 186 421 192
rect 257 167 273 181
rect 347 180 421 186
rect 257 104 265 167
rect 273 153 287 167
rect 279 108 293 116
rect 347 108 353 180
rect 414 172 421 180
rect 426 164 460 172
rect 454 159 460 164
rect 407 146 434 153
rect 313 102 353 108
rect 361 108 405 114
rect 313 84 319 102
rect 361 94 367 108
rect 473 112 479 196
rect 417 104 479 112
rect 511 153 519 196
rect 551 190 559 216
rect 537 184 559 190
rect 581 190 589 216
rect 581 184 603 190
rect 537 178 540 184
rect 511 139 513 153
rect 511 104 519 139
rect 533 122 540 178
rect 600 178 603 184
rect 537 116 540 122
rect 600 122 607 178
rect 621 153 629 196
rect 627 139 629 153
rect 600 116 603 122
rect 537 110 563 116
rect 337 88 367 94
rect 385 90 423 98
rect 415 84 423 90
rect 307 44 319 78
rect 365 70 387 82
rect 415 70 433 84
rect 361 64 373 70
rect 415 64 423 70
rect 555 64 563 110
rect 577 110 603 116
rect 577 64 585 110
rect 621 104 629 139
rect 671 153 679 196
rect 711 190 719 216
rect 697 184 719 190
rect 907 216 920 222
rect 791 210 798 216
rect 787 202 798 210
rect 848 204 855 216
rect 913 210 920 216
rect 697 178 700 184
rect 671 139 673 153
rect 671 104 679 139
rect 693 122 700 178
rect 737 181 745 196
rect 848 197 869 204
rect 827 186 833 188
rect 894 186 901 192
rect 737 167 753 181
rect 827 180 901 186
rect 697 116 700 122
rect 697 110 723 116
rect 715 64 723 110
rect 737 104 745 167
rect 753 153 767 167
rect 759 108 773 116
rect 827 108 833 180
rect 894 172 901 180
rect 906 164 940 172
rect 934 159 940 164
rect 887 146 914 153
rect 793 102 833 108
rect 841 108 885 114
rect 793 84 799 102
rect 841 94 847 108
rect 953 112 959 196
rect 981 190 989 216
rect 981 184 1003 190
rect 1000 178 1003 184
rect 1000 122 1007 178
rect 1021 153 1029 196
rect 1079 188 1091 196
rect 1079 182 1103 188
rect 1027 139 1029 153
rect 1000 116 1003 122
rect 897 104 959 112
rect 817 88 847 94
rect 865 90 903 98
rect 895 84 903 90
rect 787 44 799 78
rect 845 70 867 82
rect 895 70 913 84
rect 841 64 853 70
rect 895 64 903 70
rect 977 110 1003 116
rect 977 64 985 110
rect 1021 104 1029 139
rect 1095 133 1103 182
rect 1155 182 1163 196
rect 1183 196 1211 202
rect 1171 193 1223 196
rect 1280 216 1293 222
rect 1280 210 1287 216
rect 1345 204 1352 216
rect 1155 175 1180 182
rect 1173 153 1181 175
rect 1095 64 1103 119
rect 1179 104 1187 139
rect 1241 112 1247 196
rect 1331 197 1352 204
rect 1402 210 1409 216
rect 1402 202 1413 210
rect 1299 186 1306 192
rect 1539 236 1551 242
rect 1671 236 1683 242
rect 1717 236 1729 242
rect 1779 236 1791 242
rect 1859 236 1871 242
rect 1939 236 1951 242
rect 2071 236 2083 242
rect 2141 236 2153 242
rect 2203 236 2215 242
rect 2251 236 2263 242
rect 2309 236 2321 242
rect 2359 236 2371 242
rect 2489 236 2501 242
rect 2571 236 2583 242
rect 2651 236 2663 242
rect 2701 236 2713 242
rect 2763 236 2775 242
rect 2811 236 2823 242
rect 2869 236 2881 242
rect 2971 236 2983 242
rect 3031 236 3043 242
rect 3071 236 3083 242
rect 3171 236 3183 242
rect 3251 236 3263 242
rect 3299 236 3311 242
rect 3357 236 3369 242
rect 3405 236 3417 242
rect 3467 236 3479 242
rect 3569 236 3581 242
rect 3651 236 3663 242
rect 3717 236 3729 242
rect 3819 236 3831 242
rect 3877 236 3889 242
rect 3925 236 3937 242
rect 3987 236 3999 242
rect 4057 236 4069 242
rect 4157 236 4169 242
rect 4239 236 4251 242
rect 4339 236 4351 242
rect 4397 236 4409 242
rect 4445 236 4457 242
rect 4507 236 4519 242
rect 4577 236 4589 242
rect 4677 236 4689 242
rect 4759 236 4771 242
rect 4859 236 4871 242
rect 4917 236 4929 242
rect 4965 236 4977 242
rect 5027 236 5039 242
rect 5131 236 5143 242
rect 5197 236 5209 242
rect 5279 236 5291 242
rect 5379 236 5391 242
rect 5437 236 5449 242
rect 5485 236 5497 242
rect 5547 236 5559 242
rect 5619 236 5631 242
rect 5677 236 5689 242
rect 5725 236 5737 242
rect 5787 236 5799 242
rect 5859 236 5871 242
rect 5917 236 5929 242
rect 5965 236 5977 242
rect 6027 236 6039 242
rect 6111 236 6123 242
rect 6157 236 6169 242
rect 6311 236 6323 242
rect 6391 236 6403 242
rect 6439 236 6451 242
rect 6497 236 6509 242
rect 6545 236 6557 242
rect 6607 236 6619 242
rect 1367 186 1373 188
rect 1299 180 1373 186
rect 1455 181 1463 196
rect 1299 172 1306 180
rect 1260 164 1294 172
rect 1260 159 1266 164
rect 1286 146 1313 153
rect 1241 104 1303 112
rect 1315 108 1359 114
rect 37 18 49 24
rect 95 18 107 24
rect 141 18 153 24
rect 207 18 219 24
rect 277 18 289 24
rect 335 18 347 24
rect 381 18 393 24
rect 447 18 459 24
rect 529 18 541 24
rect 599 18 611 24
rect 689 18 701 24
rect 757 18 769 24
rect 815 18 827 24
rect 861 18 873 24
rect 927 18 939 24
rect 999 18 1011 24
rect 1071 18 1083 24
rect 1111 18 1123 24
rect 1297 90 1335 98
rect 1353 94 1359 108
rect 1367 108 1373 180
rect 1447 167 1463 181
rect 1433 153 1447 167
rect 1367 102 1407 108
rect 1427 108 1441 116
rect 1455 104 1463 167
rect 1496 161 1504 216
rect 1569 188 1581 196
rect 1557 182 1581 188
rect 1635 182 1643 196
rect 1663 196 1691 202
rect 1651 193 1703 196
rect 1297 84 1305 90
rect 1353 88 1383 94
rect 1401 84 1407 102
rect 1287 70 1305 84
rect 1333 70 1355 82
rect 1297 64 1305 70
rect 1347 64 1359 70
rect 1401 44 1413 78
rect 1496 64 1504 147
rect 1557 133 1565 182
rect 1635 175 1660 182
rect 1653 153 1661 175
rect 1736 161 1744 216
rect 1809 188 1821 196
rect 1889 188 1901 196
rect 1969 188 1981 196
rect 1797 182 1821 188
rect 1877 182 1901 188
rect 1957 182 1981 188
rect 2035 182 2043 196
rect 2063 196 2091 202
rect 2051 193 2103 196
rect 2160 216 2173 222
rect 2160 210 2167 216
rect 2225 204 2232 216
rect 1557 64 1565 119
rect 1659 104 1667 139
rect 1156 18 1168 24
rect 1206 18 1218 24
rect 1261 18 1273 24
rect 1327 18 1339 24
rect 1373 18 1385 24
rect 1431 18 1443 24
rect 1511 18 1523 24
rect 1537 18 1549 24
rect 1577 18 1589 24
rect 1736 64 1744 147
rect 1797 133 1805 182
rect 1877 133 1885 182
rect 1957 133 1965 182
rect 2035 175 2060 182
rect 2053 153 2061 175
rect 1797 64 1805 119
rect 1877 64 1885 119
rect 1957 64 1965 119
rect 2059 104 2067 139
rect 2121 112 2127 196
rect 2211 197 2232 204
rect 2282 210 2289 216
rect 2282 202 2293 210
rect 2179 186 2186 192
rect 2247 186 2253 188
rect 2179 180 2253 186
rect 2335 181 2343 196
rect 2389 188 2401 196
rect 2179 172 2186 180
rect 2140 164 2174 172
rect 2140 159 2146 164
rect 2166 146 2193 153
rect 2121 104 2183 112
rect 2195 108 2239 114
rect 1636 18 1648 24
rect 1686 18 1698 24
rect 1717 18 1729 24
rect 1777 18 1789 24
rect 1817 18 1829 24
rect 1857 18 1869 24
rect 1897 18 1909 24
rect 1937 18 1949 24
rect 1977 18 1989 24
rect 2177 90 2215 98
rect 2233 94 2239 108
rect 2247 108 2253 180
rect 2327 167 2343 181
rect 2313 153 2327 167
rect 2247 102 2287 108
rect 2307 108 2321 116
rect 2335 104 2343 167
rect 2377 182 2401 188
rect 2459 188 2471 196
rect 2459 182 2483 188
rect 2377 133 2385 182
rect 2475 133 2483 182
rect 2535 182 2543 196
rect 2563 196 2591 202
rect 2551 193 2603 196
rect 2535 175 2560 182
rect 2553 153 2561 175
rect 2636 161 2644 216
rect 2720 216 2733 222
rect 2720 210 2727 216
rect 2785 204 2792 216
rect 2177 84 2185 90
rect 2233 88 2263 94
rect 2281 84 2287 102
rect 2167 70 2185 84
rect 2213 70 2235 82
rect 2177 64 2185 70
rect 2227 64 2239 70
rect 2281 44 2293 78
rect 2377 64 2385 119
rect 2475 64 2483 119
rect 2559 104 2567 139
rect 2036 18 2048 24
rect 2086 18 2098 24
rect 2141 18 2153 24
rect 2207 18 2219 24
rect 2253 18 2265 24
rect 2311 18 2323 24
rect 2357 18 2369 24
rect 2397 18 2409 24
rect 2451 18 2463 24
rect 2491 18 2503 24
rect 2636 64 2644 147
rect 2681 112 2687 196
rect 2771 197 2792 204
rect 2842 210 2849 216
rect 2842 202 2853 210
rect 2739 186 2746 192
rect 2807 186 2813 188
rect 2739 180 2813 186
rect 2895 181 2903 196
rect 2739 172 2746 180
rect 2700 164 2734 172
rect 2700 159 2706 164
rect 2726 146 2753 153
rect 2681 104 2743 112
rect 2755 108 2799 114
rect 2737 90 2775 98
rect 2793 94 2799 108
rect 2807 108 2813 180
rect 2887 167 2903 181
rect 2935 182 2943 196
rect 2963 196 2991 202
rect 2951 193 3003 196
rect 2935 175 2960 182
rect 2873 153 2887 167
rect 2807 102 2847 108
rect 2867 108 2881 116
rect 2895 104 2903 167
rect 2953 153 2961 175
rect 3053 173 3060 216
rect 3123 230 3151 236
rect 3163 196 3191 200
rect 3135 186 3141 196
rect 3151 194 3203 196
rect 3135 179 3164 186
rect 2959 104 2967 139
rect 3053 111 3060 159
rect 3156 153 3164 179
rect 3236 161 3244 216
rect 3447 216 3460 222
rect 3331 210 3338 216
rect 3327 202 3338 210
rect 3388 204 3395 216
rect 3453 210 3460 216
rect 3277 181 3285 196
rect 3388 197 3409 204
rect 3367 186 3373 188
rect 3434 186 3441 192
rect 3277 167 3293 181
rect 3367 180 3441 186
rect 3043 104 3060 111
rect 3155 104 3163 139
rect 2737 84 2745 90
rect 2793 88 2823 94
rect 2841 84 2847 102
rect 2727 70 2745 84
rect 2773 70 2795 82
rect 2737 64 2745 70
rect 2787 64 2799 70
rect 2841 44 2853 78
rect 2536 18 2548 24
rect 2586 18 2598 24
rect 2651 18 2663 24
rect 2701 18 2713 24
rect 2767 18 2779 24
rect 2813 18 2825 24
rect 2871 18 2883 24
rect 2936 18 2948 24
rect 2986 18 2998 24
rect 3071 18 3083 24
rect 3236 64 3244 147
rect 3277 104 3285 167
rect 3293 153 3307 167
rect 3299 108 3313 116
rect 3367 108 3373 180
rect 3434 172 3441 180
rect 3446 164 3480 172
rect 3474 159 3480 164
rect 3427 146 3454 153
rect 3333 102 3373 108
rect 3381 108 3425 114
rect 3333 84 3339 102
rect 3381 94 3387 108
rect 3493 112 3499 196
rect 3539 188 3551 196
rect 3539 182 3563 188
rect 3555 133 3563 182
rect 3615 182 3623 196
rect 3643 196 3671 202
rect 3631 193 3683 196
rect 3709 196 3737 202
rect 3697 193 3749 196
rect 3967 216 3980 222
rect 3851 210 3858 216
rect 3847 202 3858 210
rect 3908 204 3915 216
rect 3973 210 3980 216
rect 3757 182 3765 196
rect 3615 175 3640 182
rect 3740 175 3765 182
rect 3797 181 3805 196
rect 3908 197 3929 204
rect 3887 186 3893 188
rect 3954 186 3961 192
rect 3633 153 3641 175
rect 3739 153 3747 175
rect 3797 167 3813 181
rect 3887 180 3961 186
rect 3437 104 3499 112
rect 3357 88 3387 94
rect 3405 90 3443 98
rect 3435 84 3443 90
rect 3327 44 3339 78
rect 3385 70 3407 82
rect 3435 70 3453 84
rect 3381 64 3393 70
rect 3435 64 3443 70
rect 3555 64 3563 119
rect 3639 104 3647 139
rect 3733 104 3741 139
rect 3797 104 3805 167
rect 3813 153 3827 167
rect 3819 108 3833 116
rect 3121 18 3133 24
rect 3191 18 3203 24
rect 3251 18 3263 24
rect 3297 18 3309 24
rect 3355 18 3367 24
rect 3401 18 3413 24
rect 3467 18 3479 24
rect 3531 18 3543 24
rect 3571 18 3583 24
rect 3616 18 3628 24
rect 3666 18 3678 24
rect 3887 108 3893 180
rect 3954 172 3961 180
rect 3966 164 4000 172
rect 3994 159 4000 164
rect 3947 146 3974 153
rect 3853 102 3893 108
rect 3901 108 3945 114
rect 3853 84 3859 102
rect 3901 94 3907 108
rect 4013 112 4019 196
rect 4049 196 4077 202
rect 4037 193 4089 196
rect 4149 196 4177 202
rect 4097 182 4105 196
rect 4137 193 4189 196
rect 4197 182 4205 196
rect 4269 188 4281 196
rect 4080 175 4105 182
rect 4180 175 4205 182
rect 4257 182 4281 188
rect 4487 216 4500 222
rect 4371 210 4378 216
rect 4367 202 4378 210
rect 4428 204 4435 216
rect 4493 210 4500 216
rect 4079 153 4087 175
rect 4179 153 4187 175
rect 3957 104 4019 112
rect 4073 104 4081 139
rect 4173 104 4181 139
rect 4257 133 4265 182
rect 4317 181 4325 196
rect 4428 197 4449 204
rect 4407 186 4413 188
rect 4474 186 4481 192
rect 4317 167 4333 181
rect 4407 180 4481 186
rect 3877 88 3907 94
rect 3925 90 3963 98
rect 3955 84 3963 90
rect 3847 44 3859 78
rect 3905 70 3927 82
rect 3955 70 3973 84
rect 3901 64 3913 70
rect 3955 64 3963 70
rect 3702 18 3714 24
rect 3752 18 3764 24
rect 3817 18 3829 24
rect 3875 18 3887 24
rect 3921 18 3933 24
rect 3987 18 3999 24
rect 4042 18 4054 24
rect 4092 18 4104 24
rect 4257 64 4265 119
rect 4317 104 4325 167
rect 4333 153 4347 167
rect 4339 108 4353 116
rect 4142 18 4154 24
rect 4192 18 4204 24
rect 4407 108 4413 180
rect 4474 172 4481 180
rect 4486 164 4520 172
rect 4514 159 4520 164
rect 4467 146 4494 153
rect 4373 102 4413 108
rect 4421 108 4465 114
rect 4373 84 4379 102
rect 4421 94 4427 108
rect 4533 112 4539 196
rect 4569 196 4597 202
rect 4557 193 4609 196
rect 4669 196 4697 202
rect 4617 182 4625 196
rect 4657 193 4709 196
rect 4717 182 4725 196
rect 4789 188 4801 196
rect 4600 175 4625 182
rect 4700 175 4725 182
rect 4777 182 4801 188
rect 5007 216 5020 222
rect 4891 210 4898 216
rect 4887 202 4898 210
rect 4948 204 4955 216
rect 5013 210 5020 216
rect 4599 153 4607 175
rect 4699 153 4707 175
rect 4477 104 4539 112
rect 4593 104 4601 139
rect 4693 104 4701 139
rect 4777 133 4785 182
rect 4837 181 4845 196
rect 4948 197 4969 204
rect 4927 186 4933 188
rect 4994 186 5001 192
rect 4837 167 4853 181
rect 4927 180 5001 186
rect 4397 88 4427 94
rect 4445 90 4483 98
rect 4475 84 4483 90
rect 4367 44 4379 78
rect 4425 70 4447 82
rect 4475 70 4493 84
rect 4421 64 4433 70
rect 4475 64 4483 70
rect 4237 18 4249 24
rect 4277 18 4289 24
rect 4337 18 4349 24
rect 4395 18 4407 24
rect 4441 18 4453 24
rect 4507 18 4519 24
rect 4562 18 4574 24
rect 4612 18 4624 24
rect 4777 64 4785 119
rect 4837 104 4845 167
rect 4853 153 4867 167
rect 4859 108 4873 116
rect 4662 18 4674 24
rect 4712 18 4724 24
rect 4927 108 4933 180
rect 4994 172 5001 180
rect 5006 164 5040 172
rect 5034 159 5040 164
rect 4987 146 5014 153
rect 4893 102 4933 108
rect 4941 108 4985 114
rect 4893 84 4899 102
rect 4941 94 4947 108
rect 5053 112 5059 196
rect 5095 182 5103 196
rect 5123 196 5151 202
rect 5111 193 5163 196
rect 5189 196 5217 202
rect 5177 193 5229 196
rect 5237 182 5245 196
rect 5309 188 5321 196
rect 5095 175 5120 182
rect 5220 175 5245 182
rect 5297 182 5321 188
rect 5527 216 5540 222
rect 5411 210 5418 216
rect 5407 202 5418 210
rect 5468 204 5475 216
rect 5533 210 5540 216
rect 5113 153 5121 175
rect 5219 153 5227 175
rect 4997 104 5059 112
rect 5119 104 5127 139
rect 5213 104 5221 139
rect 5297 133 5305 182
rect 5357 181 5365 196
rect 5468 197 5489 204
rect 5447 186 5453 188
rect 5514 186 5521 192
rect 5357 167 5373 181
rect 5447 180 5521 186
rect 4917 88 4947 94
rect 4965 90 5003 98
rect 4995 84 5003 90
rect 4887 44 4899 78
rect 4945 70 4967 82
rect 4995 70 5013 84
rect 4941 64 4953 70
rect 4995 64 5003 70
rect 4757 18 4769 24
rect 4797 18 4809 24
rect 4857 18 4869 24
rect 4915 18 4927 24
rect 4961 18 4973 24
rect 5027 18 5039 24
rect 5096 18 5108 24
rect 5146 18 5158 24
rect 5297 64 5305 119
rect 5357 104 5365 167
rect 5373 153 5387 167
rect 5379 108 5393 116
rect 5182 18 5194 24
rect 5232 18 5244 24
rect 5447 108 5453 180
rect 5514 172 5521 180
rect 5526 164 5560 172
rect 5554 159 5560 164
rect 5507 146 5534 153
rect 5413 102 5453 108
rect 5461 108 5505 114
rect 5413 84 5419 102
rect 5461 94 5467 108
rect 5573 112 5579 196
rect 5517 104 5579 112
rect 5437 88 5467 94
rect 5485 90 5523 98
rect 5515 84 5523 90
rect 5407 44 5419 78
rect 5465 70 5487 82
rect 5515 70 5533 84
rect 5461 64 5473 70
rect 5515 64 5523 70
rect 5767 216 5780 222
rect 5651 210 5658 216
rect 5647 202 5658 210
rect 5708 204 5715 216
rect 5773 210 5780 216
rect 5597 181 5605 196
rect 5708 197 5729 204
rect 5687 186 5693 188
rect 5754 186 5761 192
rect 5597 167 5613 181
rect 5687 180 5761 186
rect 5597 104 5605 167
rect 5613 153 5627 167
rect 5619 108 5633 116
rect 5687 108 5693 180
rect 5754 172 5761 180
rect 5766 164 5800 172
rect 5794 159 5800 164
rect 5747 146 5774 153
rect 5653 102 5693 108
rect 5701 108 5745 114
rect 5653 84 5659 102
rect 5701 94 5707 108
rect 5813 112 5819 196
rect 5757 104 5819 112
rect 5677 88 5707 94
rect 5725 90 5763 98
rect 5755 84 5763 90
rect 5647 44 5659 78
rect 5705 70 5727 82
rect 5755 70 5773 84
rect 5701 64 5713 70
rect 5755 64 5763 70
rect 6007 216 6020 222
rect 5891 210 5898 216
rect 5887 202 5898 210
rect 5948 204 5955 216
rect 6013 210 6020 216
rect 5837 181 5845 196
rect 5948 197 5969 204
rect 6149 196 6177 202
rect 5927 186 5933 188
rect 5994 186 6001 192
rect 5837 167 5853 181
rect 5927 180 6001 186
rect 5837 104 5845 167
rect 5853 153 5867 167
rect 5859 108 5873 116
rect 5927 108 5933 180
rect 5994 172 6001 180
rect 6006 164 6040 172
rect 6034 159 6040 164
rect 5987 146 6014 153
rect 5893 102 5933 108
rect 5941 108 5985 114
rect 5893 84 5899 102
rect 5941 94 5947 108
rect 6053 112 6059 196
rect 6096 153 6104 196
rect 6137 193 6189 196
rect 6263 230 6291 236
rect 6303 196 6331 200
rect 6197 182 6205 196
rect 6180 175 6205 182
rect 6275 186 6281 196
rect 6291 194 6343 196
rect 6275 179 6304 186
rect 6179 153 6187 175
rect 6296 153 6304 179
rect 6376 161 6384 216
rect 6587 216 6600 222
rect 6471 210 6478 216
rect 6467 202 6478 210
rect 6528 204 6535 216
rect 6593 210 6600 216
rect 6417 181 6425 196
rect 6528 197 6549 204
rect 6507 186 6513 188
rect 6574 186 6581 192
rect 6417 167 6433 181
rect 6507 180 6581 186
rect 5997 104 6059 112
rect 6096 104 6104 139
rect 6173 104 6181 139
rect 6295 104 6303 139
rect 5917 88 5947 94
rect 5965 90 6003 98
rect 5995 84 6003 90
rect 5887 44 5899 78
rect 5945 70 5967 82
rect 5995 70 6013 84
rect 5941 64 5953 70
rect 5995 64 6003 70
rect 5277 18 5289 24
rect 5317 18 5329 24
rect 5377 18 5389 24
rect 5435 18 5447 24
rect 5481 18 5493 24
rect 5547 18 5559 24
rect 5617 18 5629 24
rect 5675 18 5687 24
rect 5721 18 5733 24
rect 5787 18 5799 24
rect 5857 18 5869 24
rect 5915 18 5927 24
rect 5961 18 5973 24
rect 6027 18 6039 24
rect 6111 18 6123 24
rect 6142 18 6154 24
rect 6192 18 6204 24
rect 6376 64 6384 147
rect 6417 104 6425 167
rect 6433 153 6447 167
rect 6439 108 6453 116
rect 6507 108 6513 180
rect 6574 172 6581 180
rect 6586 164 6620 172
rect 6614 159 6620 164
rect 6567 146 6594 153
rect 6473 102 6513 108
rect 6521 108 6565 114
rect 6473 84 6479 102
rect 6521 94 6527 108
rect 6633 112 6639 196
rect 6577 104 6639 112
rect 6497 88 6527 94
rect 6545 90 6583 98
rect 6575 84 6583 90
rect 6467 44 6479 78
rect 6525 70 6547 82
rect 6575 70 6593 84
rect 6521 64 6533 70
rect 6575 64 6583 70
rect 6261 18 6273 24
rect 6331 18 6343 24
rect 6391 18 6403 24
rect 6437 18 6449 24
rect 6495 18 6507 24
rect 6541 18 6553 24
rect 6607 18 6619 24
rect -62 16 6736 18
rect -62 4 4 16
rect -62 2 6736 4
rect 6742 2 6802 242
<< m2contact >>
rect 53 6436 67 6450
rect 193 6436 207 6450
rect 93 6379 107 6393
rect 133 6379 147 6393
rect 213 6407 227 6421
rect 193 6342 207 6356
rect 293 6379 307 6393
rect 313 6387 327 6401
rect 333 6379 347 6393
rect 273 6359 287 6373
rect 353 6367 367 6381
rect 373 6359 387 6373
rect 393 6367 407 6381
rect 53 6310 67 6324
rect 193 6304 207 6318
rect 433 6413 447 6427
rect 453 6367 467 6381
rect 633 6436 647 6450
rect 473 6359 487 6373
rect 493 6367 507 6381
rect 513 6367 527 6381
rect 773 6436 787 6450
rect 613 6407 627 6421
rect 533 6359 547 6373
rect 553 6367 567 6381
rect 393 6313 407 6327
rect 633 6342 647 6356
rect 693 6379 707 6393
rect 733 6379 747 6393
rect 833 6399 847 6413
rect 853 6387 867 6401
rect 633 6304 647 6318
rect 773 6310 787 6324
rect 893 6379 907 6393
rect 913 6387 927 6401
rect 1113 6436 1127 6450
rect 1253 6436 1267 6450
rect 933 6379 947 6393
rect 953 6387 967 6401
rect 973 6379 987 6393
rect 1033 6387 1047 6401
rect 1053 6399 1067 6413
rect 1093 6407 1107 6421
rect 1113 6342 1127 6356
rect 1173 6379 1187 6393
rect 1213 6379 1227 6393
rect 1313 6379 1327 6393
rect 1333 6387 1347 6401
rect 1353 6379 1367 6393
rect 1373 6387 1387 6401
rect 1413 6393 1427 6407
rect 1453 6393 1467 6407
rect 1393 6379 1407 6393
rect 1473 6379 1487 6393
rect 1493 6387 1507 6401
rect 1513 6379 1527 6393
rect 1553 6379 1567 6393
rect 1453 6359 1467 6373
rect 1573 6367 1587 6381
rect 1113 6304 1127 6318
rect 1253 6310 1267 6324
rect 1433 6256 1447 6267
rect 1733 6436 1747 6450
rect 1873 6436 1887 6450
rect 1613 6379 1627 6393
rect 1653 6387 1667 6401
rect 1673 6399 1687 6413
rect 1713 6407 1727 6421
rect 1733 6342 1747 6356
rect 1793 6379 1807 6393
rect 1833 6379 1847 6393
rect 1933 6379 1947 6393
rect 1953 6387 1967 6401
rect 1973 6379 1987 6393
rect 1993 6359 2007 6373
rect 2033 6367 2047 6381
rect 2053 6359 2067 6373
rect 2073 6367 2087 6381
rect 2153 6379 2167 6393
rect 2173 6387 2187 6401
rect 2193 6379 2207 6393
rect 2233 6379 2247 6393
rect 2253 6387 2267 6401
rect 2273 6399 2287 6413
rect 2293 6387 2307 6401
rect 2133 6359 2147 6373
rect 1733 6304 1747 6318
rect 1873 6310 1887 6324
rect 2333 6367 2347 6381
rect 2433 6399 2447 6413
rect 2493 6399 2507 6413
rect 2353 6359 2367 6373
rect 2373 6367 2387 6381
rect 2413 6379 2427 6393
rect 2113 6256 2127 6267
rect 2453 6379 2467 6393
rect 2473 6379 2487 6393
rect 2513 6379 2527 6393
rect 2553 6367 2567 6381
rect 2573 6359 2587 6373
rect 2593 6367 2607 6381
rect 2653 6367 2667 6381
rect 2673 6359 2687 6373
rect 2713 6359 2727 6373
rect 2733 6367 2747 6381
rect 2753 6359 2767 6373
rect 2773 6367 2787 6381
rect 2833 6367 2847 6381
rect 2953 6379 2967 6393
rect 2973 6387 2987 6401
rect 2993 6379 3007 6393
rect 3053 6379 3067 6393
rect 3073 6387 3087 6401
rect 3093 6379 3107 6393
rect 3133 6387 3147 6401
rect 3153 6399 3167 6413
rect 3193 6387 3207 6401
rect 3213 6399 3227 6413
rect 3233 6387 3247 6401
rect 3253 6399 3267 6413
rect 3273 6387 3287 6401
rect 2693 6339 2707 6353
rect 2853 6359 2867 6373
rect 2893 6359 2907 6373
rect 2933 6359 2947 6373
rect 2873 6339 2887 6353
rect 3033 6359 3047 6373
rect 3293 6379 3307 6393
rect 3333 6379 3347 6393
rect 3353 6387 3367 6401
rect 3373 6379 3387 6393
rect 3453 6379 3467 6393
rect 3473 6387 3487 6401
rect 3493 6399 3507 6413
rect 3513 6387 3527 6401
rect 3553 6379 3567 6393
rect 3573 6387 3587 6401
rect 3593 6399 3607 6413
rect 3613 6387 3627 6401
rect 3393 6359 3407 6373
rect 3633 6359 3647 6373
rect 3673 6359 3687 6373
rect 3693 6367 3707 6381
rect 3773 6379 3787 6393
rect 3793 6387 3807 6401
rect 3813 6379 3827 6393
rect 3833 6379 3847 6393
rect 3853 6387 3867 6401
rect 3933 6399 3947 6413
rect 3873 6379 3887 6393
rect 3953 6387 3967 6401
rect 3653 6339 3667 6353
rect 3753 6359 3767 6373
rect 3893 6359 3907 6373
rect 3993 6367 4007 6381
rect 4013 6359 4027 6373
rect 4033 6367 4047 6381
rect 4093 6379 4107 6393
rect 4113 6367 4127 6381
rect 4153 6379 4167 6393
rect 4173 6367 4187 6381
rect 4553 6399 4567 6413
rect 4573 6387 4587 6401
rect 4613 6387 4627 6401
rect 4633 6399 4647 6413
rect 4653 6387 4667 6401
rect 4693 6413 4707 6427
rect 4193 6359 4207 6373
rect 4213 6367 4227 6381
rect 4273 6367 4287 6381
rect 4293 6359 4307 6373
rect 4333 6359 4347 6373
rect 4373 6367 4387 6381
rect 4313 6339 4327 6353
rect 4393 6359 4407 6373
rect 4433 6359 4447 6373
rect 4473 6367 4487 6381
rect 4413 6339 4427 6353
rect 4493 6359 4507 6373
rect 4533 6359 4547 6373
rect 4513 6339 4527 6353
rect 4673 6379 4687 6393
rect 4593 6353 4607 6367
rect 4633 6353 4647 6367
rect 4713 6387 4727 6401
rect 4733 6399 4747 6413
rect 4753 6387 4767 6401
rect 4773 6379 4787 6393
rect 4813 6379 4827 6393
rect 4833 6387 4847 6401
rect 4873 6393 4887 6407
rect 4893 6393 4907 6407
rect 4853 6379 4867 6393
rect 4953 6379 4967 6393
rect 4973 6387 4987 6401
rect 4993 6379 5007 6393
rect 5013 6379 5027 6393
rect 5033 6387 5047 6401
rect 5053 6379 5067 6393
rect 5213 6433 5227 6447
rect 4713 6353 4727 6367
rect 4873 6359 4887 6373
rect 4933 6359 4947 6373
rect 5073 6359 5087 6373
rect 5133 6367 5147 6381
rect 4873 6313 4887 6327
rect 4913 6313 4927 6327
rect 5153 6359 5167 6373
rect 5193 6359 5207 6373
rect 5173 6339 5187 6353
rect 5193 6313 5207 6327
rect 5273 6393 5287 6407
rect 5313 6393 5327 6407
rect 5413 6387 5427 6401
rect 5433 6399 5447 6413
rect 5453 6387 5467 6401
rect 5233 6367 5247 6381
rect 5253 6359 5267 6373
rect 5293 6359 5307 6373
rect 5333 6367 5347 6381
rect 5473 6379 5487 6393
rect 5533 6379 5547 6393
rect 5553 6387 5567 6401
rect 5573 6399 5587 6413
rect 5593 6387 5607 6401
rect 5633 6387 5647 6401
rect 5653 6399 5667 6413
rect 5673 6387 5687 6401
rect 5693 6399 5707 6413
rect 5713 6387 5727 6401
rect 5273 6339 5287 6353
rect 5353 6359 5367 6373
rect 5393 6359 5407 6373
rect 5373 6339 5387 6353
rect 5733 6379 5747 6393
rect 5773 6359 5787 6373
rect 5813 6359 5827 6373
rect 5833 6367 5847 6381
rect 5893 6379 5907 6393
rect 5913 6387 5927 6401
rect 5933 6399 5947 6413
rect 6013 6433 6027 6447
rect 5953 6387 5967 6401
rect 5993 6387 6007 6401
rect 6013 6399 6027 6413
rect 5793 6339 5807 6353
rect 6013 6353 6027 6367
rect 6053 6379 6067 6393
rect 6073 6387 6087 6401
rect 6093 6399 6107 6413
rect 6113 6387 6127 6401
rect 6153 6393 6167 6407
rect 6173 6379 6187 6393
rect 6193 6387 6207 6401
rect 6213 6379 6227 6393
rect 6253 6379 6267 6393
rect 6273 6387 6287 6401
rect 6293 6399 6307 6413
rect 6313 6387 6327 6401
rect 6533 6399 6547 6413
rect 6553 6387 6567 6401
rect 6153 6359 6167 6373
rect 6333 6359 6347 6373
rect 6373 6359 6387 6373
rect 6393 6367 6407 6381
rect 6453 6367 6467 6381
rect 6153 6313 6167 6327
rect 6353 6339 6367 6353
rect 6473 6359 6487 6373
rect 6513 6359 6527 6373
rect 6493 6339 6507 6353
rect 6593 6379 6607 6393
rect 6613 6387 6627 6401
rect 6633 6379 6647 6393
rect 6653 6387 6667 6401
rect 6673 6379 6687 6393
rect 1433 6253 1447 6256
rect 2113 6253 2127 6256
rect 1893 6244 1907 6247
rect 53 6182 67 6196
rect 193 6176 207 6190
rect 53 6144 67 6158
rect 33 6079 47 6093
rect 113 6107 127 6121
rect 153 6107 167 6121
rect 53 6050 67 6064
rect 273 6107 287 6121
rect 373 6119 387 6133
rect 393 6127 407 6141
rect 193 6050 207 6064
rect 293 6099 307 6113
rect 313 6087 327 6101
rect 333 6099 347 6113
rect 413 6119 427 6133
rect 433 6107 447 6121
rect 473 6107 487 6121
rect 533 6119 547 6133
rect 553 6127 567 6141
rect 453 6087 467 6101
rect 573 6119 587 6133
rect 653 6127 667 6141
rect 713 6127 727 6141
rect 593 6107 607 6121
rect 613 6099 627 6113
rect 633 6107 647 6121
rect 733 6107 747 6121
rect 753 6099 767 6113
rect 773 6107 787 6121
rect 793 6107 807 6121
rect 833 6107 847 6121
rect 893 6107 907 6121
rect 813 6087 827 6101
rect 913 6099 927 6113
rect 933 6087 947 6101
rect 953 6099 967 6113
rect 993 6107 1007 6121
rect 973 6087 987 6101
rect 1033 6099 1047 6113
rect 1093 6099 1107 6113
rect 1133 6107 1147 6121
rect 1233 6127 1247 6141
rect 1173 6107 1187 6121
rect 1253 6107 1267 6121
rect 1113 6087 1127 6101
rect 1153 6087 1167 6101
rect 1273 6099 1287 6113
rect 1293 6107 1307 6121
rect 1333 6099 1347 6113
rect 1353 6087 1367 6101
rect 1393 6099 1407 6113
rect 1433 6107 1447 6121
rect 1473 6107 1487 6121
rect 1513 6107 1527 6121
rect 1553 6107 1567 6121
rect 1893 6233 1907 6244
rect 1413 6087 1427 6101
rect 1453 6087 1467 6101
rect 1533 6087 1547 6101
rect 1593 6087 1607 6101
rect 1613 6099 1627 6113
rect 1653 6107 1667 6121
rect 1693 6107 1707 6121
rect 1713 6113 1727 6127
rect 1673 6087 1687 6101
rect 1693 6073 1707 6087
rect 1733 6107 1747 6121
rect 1793 6133 1807 6147
rect 1773 6107 1787 6121
rect 1753 6087 1767 6101
rect 1873 6127 1887 6141
rect 1813 6107 1827 6121
rect 1833 6099 1847 6113
rect 1853 6107 1867 6121
rect 1913 6087 1927 6101
rect 1933 6099 1947 6113
rect 1993 6107 2007 6121
rect 2133 6153 2147 6167
rect 1773 6053 1787 6067
rect 2013 6099 2027 6113
rect 2033 6087 2047 6101
rect 2053 6099 2067 6113
rect 2073 6087 2087 6101
rect 2093 6099 2107 6113
rect 2153 6127 2167 6141
rect 2173 6107 2187 6121
rect 2133 6073 2147 6087
rect 2193 6099 2207 6113
rect 2213 6107 2227 6121
rect 2233 6087 2247 6101
rect 2253 6099 2267 6113
rect 2313 6173 2327 6187
rect 2313 6127 2327 6141
rect 2453 6147 2467 6161
rect 2333 6107 2347 6121
rect 2313 6093 2327 6107
rect 2353 6099 2367 6113
rect 2373 6107 2387 6121
rect 2413 6119 2427 6133
rect 2433 6127 2447 6141
rect 2473 6127 2487 6141
rect 2513 6107 2527 6121
rect 2533 6099 2547 6113
rect 2553 6087 2567 6101
rect 2573 6099 2587 6113
rect 2613 6107 2627 6121
rect 2733 6147 2747 6161
rect 2653 6107 2667 6121
rect 2693 6119 2707 6133
rect 2713 6127 2727 6141
rect 2753 6127 2767 6141
rect 2633 6087 2647 6101
rect 2793 6107 2807 6121
rect 2813 6099 2827 6113
rect 2833 6107 2847 6121
rect 2853 6099 2867 6113
rect 2873 6107 2887 6121
rect 2973 6147 2987 6161
rect 2953 6127 2967 6141
rect 2993 6127 3007 6141
rect 3013 6119 3027 6133
rect 3213 6147 3227 6161
rect 2913 6099 2927 6113
rect 2933 6087 2947 6101
rect 3073 6107 3087 6121
rect 3173 6119 3187 6133
rect 3193 6127 3207 6141
rect 3233 6127 3247 6141
rect 3093 6099 3107 6113
rect 3113 6087 3127 6101
rect 3133 6099 3147 6113
rect 3273 6107 3287 6121
rect 3473 6147 3487 6161
rect 3533 6147 3547 6161
rect 3433 6119 3447 6133
rect 3453 6127 3467 6141
rect 3493 6127 3507 6141
rect 3513 6127 3527 6141
rect 3553 6127 3567 6141
rect 3593 6153 3607 6167
rect 3573 6119 3587 6133
rect 3293 6099 3307 6113
rect 3313 6087 3327 6101
rect 3333 6099 3347 6113
rect 3373 6099 3387 6113
rect 3393 6087 3407 6101
rect 3613 6087 3627 6101
rect 3633 6099 3647 6113
rect 3673 6099 3687 6113
rect 3593 6073 3607 6087
rect 3693 6087 3707 6101
rect 3713 6099 3727 6113
rect 3733 6107 3747 6121
rect 3793 6119 3807 6133
rect 3813 6127 3827 6141
rect 3833 6119 3847 6133
rect 3853 6119 3867 6133
rect 3873 6127 3887 6141
rect 3893 6119 3907 6133
rect 3953 6127 3967 6141
rect 4093 6127 4107 6141
rect 3973 6107 3987 6121
rect 3993 6099 4007 6113
rect 4013 6107 4027 6121
rect 4033 6107 4047 6121
rect 4053 6099 4067 6113
rect 4073 6107 4087 6121
rect 4153 6107 4167 6121
rect 4193 6107 4207 6121
rect 4293 6119 4307 6133
rect 4313 6127 4327 6141
rect 4173 6087 4187 6101
rect 4213 6087 4227 6101
rect 4233 6099 4247 6113
rect 4333 6119 4347 6133
rect 4353 6107 4367 6121
rect 4393 6119 4407 6133
rect 4473 6127 4487 6141
rect 4673 6147 4687 6161
rect 4653 6127 4667 6141
rect 4693 6127 4707 6141
rect 4413 6107 4427 6121
rect 4493 6107 4507 6121
rect 4513 6099 4527 6113
rect 4533 6107 4547 6121
rect 4573 6107 4587 6121
rect 4713 6119 4727 6133
rect 4913 6147 4927 6161
rect 4973 6147 4987 6161
rect 4593 6099 4607 6113
rect 4613 6087 4627 6101
rect 4633 6099 4647 6113
rect 4773 6107 4787 6121
rect 4873 6119 4887 6133
rect 4893 6127 4907 6141
rect 4933 6127 4947 6141
rect 4953 6127 4967 6141
rect 4993 6127 5007 6141
rect 5013 6119 5027 6133
rect 5073 6127 5087 6141
rect 4793 6099 4807 6113
rect 4813 6087 4827 6101
rect 4833 6099 4847 6113
rect 5093 6107 5107 6121
rect 5113 6099 5127 6113
rect 5133 6107 5147 6121
rect 5173 6119 5187 6133
rect 5193 6127 5207 6141
rect 5213 6119 5227 6133
rect 5233 6107 5247 6121
rect 5273 6119 5287 6133
rect 5393 6127 5407 6141
rect 5593 6147 5607 6161
rect 5653 6147 5667 6161
rect 5293 6107 5307 6121
rect 5333 6107 5347 6121
rect 5353 6099 5367 6113
rect 5373 6107 5387 6121
rect 5453 6107 5467 6121
rect 5553 6119 5567 6133
rect 5573 6127 5587 6141
rect 5613 6127 5627 6141
rect 5633 6127 5647 6141
rect 5673 6127 5687 6141
rect 5693 6119 5707 6133
rect 5853 6147 5867 6161
rect 5833 6127 5847 6141
rect 5873 6127 5887 6141
rect 5473 6099 5487 6113
rect 5493 6087 5507 6101
rect 5513 6099 5527 6113
rect 5753 6107 5767 6121
rect 5893 6119 5907 6133
rect 5993 6127 6007 6141
rect 6153 6147 6167 6161
rect 6093 6127 6107 6141
rect 6133 6127 6147 6141
rect 6173 6127 6187 6141
rect 5773 6099 5787 6113
rect 5793 6087 5807 6101
rect 5813 6099 5827 6113
rect 5933 6107 5947 6121
rect 5953 6099 5967 6113
rect 5973 6107 5987 6121
rect 6033 6107 6047 6121
rect 6053 6099 6067 6113
rect 6073 6107 6087 6121
rect 6193 6119 6207 6133
rect 6233 6173 6247 6187
rect 6253 6147 6267 6161
rect 6233 6127 6247 6141
rect 6273 6127 6287 6141
rect 6393 6147 6407 6161
rect 6293 6119 6307 6133
rect 6353 6119 6367 6133
rect 6373 6127 6387 6141
rect 6413 6127 6427 6141
rect 6233 6093 6247 6107
rect 6453 6107 6467 6121
rect 6473 6099 6487 6113
rect 6493 6087 6507 6101
rect 6513 6099 6527 6113
rect 6533 6087 6547 6101
rect 6553 6099 6567 6113
rect 6593 6087 6607 6101
rect 6613 6099 6627 6113
rect 33 5899 47 5913
rect 73 5899 87 5913
rect 93 5887 107 5901
rect 113 5879 127 5893
rect 133 5887 147 5901
rect 173 5887 187 5901
rect 193 5879 207 5893
rect 213 5887 227 5901
rect 273 5899 287 5913
rect 293 5907 307 5921
rect 313 5919 327 5933
rect 333 5907 347 5921
rect 373 5887 387 5901
rect 433 5919 447 5933
rect 453 5907 467 5921
rect 533 5919 547 5933
rect 593 5919 607 5933
rect 393 5879 407 5893
rect 413 5887 427 5901
rect 513 5899 527 5913
rect 553 5899 567 5913
rect 573 5899 587 5913
rect 613 5899 627 5913
rect 653 5933 667 5947
rect 653 5899 667 5913
rect 673 5907 687 5921
rect 693 5899 707 5913
rect 773 5907 787 5921
rect 793 5919 807 5933
rect 833 5919 847 5933
rect 633 5853 647 5867
rect 713 5879 727 5893
rect 813 5899 827 5913
rect 853 5899 867 5913
rect 913 5887 927 5901
rect 933 5879 947 5893
rect 953 5887 967 5901
rect 1013 5899 1027 5913
rect 1033 5907 1047 5921
rect 1093 5919 1107 5933
rect 1253 5956 1267 5970
rect 1393 5956 1407 5970
rect 1053 5899 1067 5913
rect 1073 5899 1087 5913
rect 993 5879 1007 5893
rect 1113 5899 1127 5913
rect 1173 5907 1187 5921
rect 1193 5919 1207 5933
rect 1233 5927 1247 5941
rect 1253 5862 1267 5876
rect 1313 5899 1327 5913
rect 1353 5899 1367 5913
rect 1453 5887 1467 5901
rect 1633 5913 1647 5927
rect 1473 5879 1487 5893
rect 1493 5887 1507 5901
rect 1553 5887 1567 5901
rect 1253 5824 1267 5838
rect 1393 5830 1407 5844
rect 1573 5879 1587 5893
rect 1613 5879 1627 5893
rect 1593 5859 1607 5873
rect 1613 5833 1627 5847
rect 1673 5899 1687 5913
rect 1693 5907 1707 5921
rect 1773 5919 1787 5933
rect 1713 5899 1727 5913
rect 1753 5899 1767 5913
rect 1653 5879 1667 5893
rect 1793 5899 1807 5913
rect 1913 5919 1927 5933
rect 1933 5907 1947 5921
rect 1953 5913 1967 5927
rect 1833 5887 1847 5901
rect 1633 5776 1647 5787
rect 1733 5776 1747 5787
rect 1853 5879 1867 5893
rect 1893 5879 1907 5893
rect 1873 5859 1887 5873
rect 1953 5833 1967 5847
rect 1993 5913 2007 5927
rect 2013 5899 2027 5913
rect 2033 5907 2047 5921
rect 2053 5899 2067 5913
rect 1993 5879 2007 5893
rect 2073 5879 2087 5893
rect 2113 5879 2127 5893
rect 2133 5887 2147 5901
rect 2193 5899 2207 5913
rect 2213 5907 2227 5921
rect 2233 5919 2247 5933
rect 2253 5907 2267 5921
rect 2273 5899 2287 5913
rect 2293 5907 2307 5921
rect 2313 5899 2327 5913
rect 1993 5833 2007 5847
rect 2093 5859 2107 5873
rect 2333 5879 2347 5893
rect 2393 5887 2407 5901
rect 2413 5879 2427 5893
rect 2433 5887 2447 5901
rect 2473 5887 2487 5901
rect 2573 5899 2587 5913
rect 2593 5907 2607 5921
rect 2613 5919 2627 5933
rect 2633 5907 2647 5921
rect 2493 5879 2507 5893
rect 2533 5879 2547 5893
rect 2513 5859 2527 5873
rect 2653 5887 2667 5901
rect 2953 5953 2967 5967
rect 2673 5879 2687 5893
rect 2693 5887 2707 5901
rect 2753 5887 2767 5901
rect 2773 5879 2787 5893
rect 2813 5879 2827 5893
rect 2853 5887 2867 5901
rect 2893 5893 2907 5907
rect 3093 5913 3107 5927
rect 3133 5913 3147 5927
rect 2793 5859 2807 5873
rect 2873 5879 2887 5893
rect 2913 5879 2927 5893
rect 2953 5887 2967 5901
rect 2893 5859 2907 5873
rect 2973 5879 2987 5893
rect 3013 5879 3027 5893
rect 3053 5887 3067 5901
rect 2993 5859 3007 5873
rect 3073 5879 3087 5893
rect 3113 5879 3127 5893
rect 3133 5879 3147 5893
rect 3173 5879 3187 5893
rect 3193 5887 3207 5901
rect 3273 5899 3287 5913
rect 3293 5907 3307 5921
rect 3313 5899 3327 5913
rect 3333 5899 3347 5913
rect 3353 5907 3367 5921
rect 3373 5899 3387 5913
rect 3453 5899 3467 5913
rect 3473 5907 3487 5921
rect 3493 5919 3507 5933
rect 3513 5907 3527 5921
rect 3573 5899 3587 5913
rect 3593 5907 3607 5921
rect 3613 5899 3627 5913
rect 3733 5907 3747 5921
rect 3753 5919 3767 5933
rect 3773 5907 3787 5921
rect 3093 5859 3107 5873
rect 3153 5859 3167 5873
rect 3253 5879 3267 5893
rect 3393 5879 3407 5893
rect 3553 5879 3567 5893
rect 3653 5887 3667 5901
rect 3793 5899 3807 5913
rect 3673 5879 3687 5893
rect 3713 5879 3727 5893
rect 3693 5859 3707 5873
rect 3853 5887 3867 5901
rect 3953 5899 3967 5913
rect 3973 5907 3987 5921
rect 3993 5919 4007 5933
rect 4013 5907 4027 5921
rect 4093 5913 4107 5927
rect 3873 5879 3887 5893
rect 3913 5879 3927 5893
rect 3893 5859 3907 5873
rect 4053 5887 4067 5901
rect 4093 5893 4107 5907
rect 4153 5899 4167 5913
rect 4173 5907 4187 5921
rect 4193 5919 4207 5933
rect 4213 5907 4227 5921
rect 3973 5873 3987 5887
rect 4013 5873 4027 5887
rect 4073 5879 4087 5893
rect 4113 5879 4127 5893
rect 4093 5859 4107 5873
rect 4233 5879 4247 5893
rect 4273 5879 4287 5893
rect 4293 5887 4307 5901
rect 4333 5887 4347 5901
rect 4253 5859 4267 5873
rect 4353 5879 4367 5893
rect 4373 5887 4387 5901
rect 4453 5899 4467 5913
rect 4473 5907 4487 5921
rect 4553 5919 4567 5933
rect 4493 5899 4507 5913
rect 4533 5899 4547 5913
rect 4433 5879 4447 5893
rect 4573 5899 4587 5913
rect 4593 5899 4607 5913
rect 4633 5887 4647 5901
rect 4653 5899 4667 5913
rect 4713 5899 4727 5913
rect 4733 5907 4747 5921
rect 4753 5919 4767 5933
rect 4773 5907 4787 5921
rect 4793 5887 4807 5901
rect 4893 5907 4907 5921
rect 4913 5919 4927 5933
rect 4813 5879 4827 5893
rect 4833 5887 4847 5901
rect 5033 5907 5047 5921
rect 5053 5919 5067 5933
rect 5073 5907 5087 5921
rect 4953 5887 4967 5901
rect 5093 5899 5107 5913
rect 5133 5899 5147 5913
rect 5153 5907 5167 5921
rect 5173 5899 5187 5913
rect 5233 5899 5247 5913
rect 5253 5907 5267 5921
rect 5273 5899 5287 5913
rect 5333 5899 5347 5913
rect 5353 5907 5367 5921
rect 5373 5899 5387 5913
rect 5393 5907 5407 5921
rect 5413 5899 5427 5913
rect 4973 5879 4987 5893
rect 5013 5879 5027 5893
rect 4993 5859 5007 5873
rect 5193 5879 5207 5893
rect 5293 5879 5307 5893
rect 5473 5887 5487 5901
rect 5533 5919 5547 5933
rect 5573 5933 5587 5947
rect 5553 5907 5567 5921
rect 5493 5879 5507 5893
rect 5513 5887 5527 5901
rect 5613 5953 5627 5967
rect 5693 5907 5707 5921
rect 5713 5919 5727 5933
rect 5733 5907 5747 5921
rect 5613 5887 5627 5901
rect 5753 5899 5767 5913
rect 5833 5899 5847 5913
rect 5853 5907 5867 5921
rect 5873 5899 5887 5913
rect 5893 5899 5907 5913
rect 5913 5907 5927 5921
rect 5933 5899 5947 5913
rect 6033 5899 6047 5913
rect 6053 5907 6067 5921
rect 6073 5899 6087 5913
rect 6093 5899 6107 5913
rect 6113 5907 6127 5921
rect 6133 5899 6147 5913
rect 6153 5907 6167 5921
rect 6173 5899 6187 5913
rect 5593 5853 5607 5867
rect 5573 5833 5587 5847
rect 5633 5879 5647 5893
rect 5673 5879 5687 5893
rect 5653 5859 5667 5873
rect 5693 5873 5707 5887
rect 5733 5873 5747 5887
rect 5813 5879 5827 5893
rect 5953 5879 5967 5893
rect 6013 5879 6027 5893
rect 6233 5887 6247 5901
rect 6253 5879 6267 5893
rect 6273 5887 6287 5901
rect 6293 5899 6307 5913
rect 6333 5887 6347 5901
rect 6353 5899 6367 5913
rect 6393 5899 6407 5913
rect 6413 5907 6427 5921
rect 6473 5913 6487 5927
rect 6433 5899 6447 5913
rect 6453 5879 6467 5893
rect 6493 5879 6507 5893
rect 6533 5879 6547 5893
rect 6553 5887 6567 5901
rect 6573 5893 6587 5907
rect 6513 5859 6527 5873
rect 6493 5833 6507 5847
rect 6593 5887 6607 5901
rect 6613 5879 6627 5893
rect 6633 5887 6647 5901
rect 6593 5853 6607 5867
rect 1633 5773 1647 5776
rect 1733 5773 1747 5776
rect 33 5627 47 5641
rect 213 5702 227 5716
rect 353 5696 367 5710
rect 73 5627 87 5641
rect 113 5627 127 5641
rect 153 5627 167 5641
rect 213 5664 227 5678
rect 193 5599 207 5613
rect 273 5627 287 5641
rect 313 5627 327 5641
rect 213 5570 227 5584
rect 433 5627 447 5641
rect 353 5570 367 5584
rect 473 5627 487 5641
rect 453 5607 467 5621
rect 493 5619 507 5633
rect 513 5607 527 5621
rect 533 5619 547 5633
rect 553 5627 567 5641
rect 593 5639 607 5653
rect 613 5647 627 5661
rect 633 5639 647 5653
rect 673 5627 687 5641
rect 713 5639 727 5653
rect 733 5627 747 5641
rect 773 5639 787 5653
rect 793 5647 807 5661
rect 813 5639 827 5653
rect 853 5639 867 5653
rect 873 5647 887 5661
rect 893 5639 907 5653
rect 933 5627 947 5641
rect 973 5627 987 5641
rect 953 5607 967 5621
rect 1013 5607 1027 5621
rect 1033 5619 1047 5633
rect 1093 5627 1107 5641
rect 1073 5607 1087 5621
rect 1133 5619 1147 5633
rect 1173 5627 1187 5641
rect 1213 5627 1227 5641
rect 1193 5607 1207 5621
rect 1253 5607 1267 5621
rect 1273 5619 1287 5633
rect 1313 5627 1327 5641
rect 1353 5627 1367 5641
rect 1493 5702 1507 5716
rect 1633 5696 1647 5710
rect 1333 5607 1347 5621
rect 1393 5607 1407 5621
rect 1413 5619 1427 5633
rect 1493 5664 1507 5678
rect 1473 5599 1487 5613
rect 1553 5627 1567 5641
rect 1593 5627 1607 5641
rect 1493 5570 1507 5584
rect 1833 5647 1847 5661
rect 1693 5627 1707 5641
rect 1713 5619 1727 5633
rect 1733 5627 1747 5641
rect 1753 5619 1767 5633
rect 1773 5627 1787 5641
rect 1853 5627 1867 5641
rect 1873 5619 1887 5633
rect 1893 5627 1907 5641
rect 1933 5639 1947 5653
rect 1953 5647 1967 5661
rect 1633 5570 1647 5584
rect 1973 5639 1987 5653
rect 1993 5607 2007 5621
rect 2013 5619 2027 5633
rect 2073 5627 2087 5641
rect 2093 5619 2107 5633
rect 2113 5607 2127 5621
rect 2133 5619 2147 5633
rect 2153 5627 2167 5641
rect 2193 5627 2207 5641
rect 2233 5639 2247 5653
rect 2253 5647 2267 5661
rect 2173 5607 2187 5621
rect 2273 5639 2287 5653
rect 2573 5673 2587 5687
rect 2353 5619 2367 5633
rect 2393 5627 2407 5641
rect 2413 5619 2427 5633
rect 2453 5627 2467 5641
rect 2513 5639 2527 5653
rect 2533 5647 2547 5661
rect 2553 5639 2567 5653
rect 2553 5593 2567 5607
rect 2633 5667 2647 5681
rect 2673 5673 2687 5687
rect 2593 5639 2607 5653
rect 2613 5647 2627 5661
rect 2653 5647 2667 5661
rect 2733 5667 2747 5681
rect 2693 5639 2707 5653
rect 2713 5647 2727 5661
rect 2753 5647 2767 5661
rect 2773 5639 2787 5653
rect 2793 5647 2807 5661
rect 2673 5613 2687 5627
rect 2813 5639 2827 5653
rect 2913 5647 2927 5661
rect 3013 5667 3027 5681
rect 2853 5627 2867 5641
rect 2873 5619 2887 5633
rect 2893 5627 2907 5641
rect 2973 5639 2987 5653
rect 2993 5647 3007 5661
rect 3033 5647 3047 5661
rect 3173 5647 3187 5661
rect 3053 5619 3067 5633
rect 3073 5607 3087 5621
rect 3093 5619 3107 5633
rect 3113 5627 3127 5641
rect 3193 5627 3207 5641
rect 3213 5619 3227 5633
rect 3233 5627 3247 5641
rect 3333 5667 3347 5681
rect 3313 5647 3327 5661
rect 3353 5647 3367 5661
rect 3473 5667 3487 5681
rect 3373 5639 3387 5653
rect 3433 5639 3447 5653
rect 3453 5647 3467 5661
rect 3493 5647 3507 5661
rect 3573 5667 3587 5681
rect 3533 5639 3547 5653
rect 3553 5647 3567 5661
rect 3593 5647 3607 5661
rect 3273 5619 3287 5633
rect 3293 5607 3307 5621
rect 3473 5613 3487 5627
rect 3513 5613 3527 5627
rect 3693 5647 3707 5661
rect 3633 5619 3647 5633
rect 3713 5627 3727 5641
rect 3653 5607 3667 5621
rect 3733 5619 3747 5633
rect 3753 5627 3767 5641
rect 3793 5627 3807 5641
rect 3913 5647 3927 5661
rect 3833 5627 3847 5641
rect 3853 5627 3867 5641
rect 3813 5607 3827 5621
rect 3873 5619 3887 5633
rect 3893 5627 3907 5641
rect 3973 5619 3987 5633
rect 4033 5627 4047 5641
rect 3993 5607 4007 5621
rect 4053 5619 4067 5633
rect 4073 5627 4087 5641
rect 4093 5619 4107 5633
rect 4113 5627 4127 5641
rect 4153 5693 4167 5707
rect 4153 5647 4167 5661
rect 4293 5667 4307 5681
rect 4173 5627 4187 5641
rect 4153 5613 4167 5627
rect 4193 5619 4207 5633
rect 4213 5627 4227 5641
rect 4253 5639 4267 5653
rect 4273 5647 4287 5661
rect 4313 5647 4327 5661
rect 4413 5647 4427 5661
rect 4333 5607 4347 5621
rect 4353 5619 4367 5633
rect 4433 5627 4447 5641
rect 4453 5619 4467 5633
rect 4473 5627 4487 5641
rect 4513 5627 4527 5641
rect 4533 5639 4547 5653
rect 4853 5713 4867 5727
rect 4573 5627 4587 5641
rect 4593 5639 4607 5653
rect 4613 5647 4627 5661
rect 4633 5639 4647 5653
rect 4693 5647 4707 5661
rect 4833 5647 4847 5661
rect 4713 5627 4727 5641
rect 4733 5619 4747 5633
rect 4753 5627 4767 5641
rect 4773 5627 4787 5641
rect 4793 5619 4807 5633
rect 4813 5627 4827 5641
rect 4833 5613 4847 5627
rect 4933 5667 4947 5681
rect 4893 5639 4907 5653
rect 4913 5647 4927 5661
rect 4953 5647 4967 5661
rect 5053 5653 5067 5667
rect 4973 5619 4987 5633
rect 4993 5607 5007 5621
rect 5013 5619 5027 5633
rect 5033 5627 5047 5641
rect 4893 5573 4907 5587
rect 5133 5647 5147 5661
rect 5073 5627 5087 5641
rect 5093 5619 5107 5633
rect 5113 5627 5127 5641
rect 5173 5693 5187 5707
rect 5193 5667 5207 5681
rect 5173 5647 5187 5661
rect 5213 5647 5227 5661
rect 5253 5673 5267 5687
rect 5233 5639 5247 5653
rect 5193 5613 5207 5627
rect 5053 5573 5067 5587
rect 5233 5573 5247 5587
rect 5373 5667 5387 5681
rect 5273 5639 5287 5653
rect 5293 5647 5307 5661
rect 5313 5639 5327 5653
rect 5353 5647 5367 5661
rect 5393 5647 5407 5661
rect 5413 5639 5427 5653
rect 5453 5619 5467 5633
rect 5473 5607 5487 5621
rect 5493 5619 5507 5633
rect 5513 5627 5527 5641
rect 5553 5639 5567 5653
rect 5573 5647 5587 5661
rect 5593 5639 5607 5653
rect 5653 5673 5667 5687
rect 5653 5639 5667 5653
rect 5673 5647 5687 5661
rect 5693 5639 5707 5653
rect 5853 5647 5867 5661
rect 5713 5627 5727 5641
rect 5733 5619 5747 5633
rect 5753 5627 5767 5641
rect 5773 5619 5787 5633
rect 5793 5627 5807 5641
rect 5873 5627 5887 5641
rect 5893 5619 5907 5633
rect 5913 5627 5927 5641
rect 6133 5667 6147 5681
rect 6113 5647 6127 5661
rect 6153 5647 6167 5661
rect 5933 5607 5947 5621
rect 5953 5619 5967 5633
rect 5993 5627 6007 5641
rect 6013 5619 6027 5633
rect 5633 5553 5647 5567
rect 6033 5627 6047 5641
rect 6053 5619 6067 5633
rect 6073 5627 6087 5641
rect 6173 5639 6187 5653
rect 6353 5653 6367 5667
rect 6393 5667 6407 5681
rect 6233 5619 6247 5633
rect 6253 5607 6267 5621
rect 6273 5619 6287 5633
rect 6293 5607 6307 5621
rect 6313 5619 6327 5633
rect 6333 5627 6347 5641
rect 6373 5647 6387 5661
rect 6413 5647 6427 5661
rect 6453 5693 6467 5707
rect 6433 5639 6447 5653
rect 6493 5667 6507 5681
rect 6473 5647 6487 5661
rect 6513 5647 6527 5661
rect 6593 5667 6607 5681
rect 6533 5639 6547 5653
rect 6573 5647 6587 5661
rect 6613 5647 6627 5661
rect 6633 5639 6647 5653
rect 6453 5613 6467 5627
rect 6353 5593 6367 5607
rect 53 5476 67 5490
rect 193 5476 207 5490
rect 33 5447 47 5461
rect 53 5382 67 5396
rect 113 5419 127 5433
rect 153 5419 167 5433
rect 253 5407 267 5421
rect 273 5399 287 5413
rect 293 5407 307 5421
rect 353 5419 367 5433
rect 373 5427 387 5441
rect 393 5439 407 5453
rect 413 5427 427 5441
rect 53 5344 67 5358
rect 193 5350 207 5364
rect 453 5407 467 5421
rect 473 5399 487 5413
rect 493 5407 507 5421
rect 533 5419 547 5433
rect 553 5407 567 5421
rect 913 5473 927 5487
rect 633 5439 647 5453
rect 713 5439 727 5453
rect 593 5419 607 5433
rect 613 5419 627 5433
rect 653 5419 667 5433
rect 693 5419 707 5433
rect 733 5419 747 5433
rect 773 5407 787 5421
rect 793 5399 807 5413
rect 813 5407 827 5421
rect 853 5407 867 5421
rect 873 5399 887 5413
rect 893 5407 907 5421
rect 933 5439 947 5453
rect 1253 5476 1267 5490
rect 953 5427 967 5441
rect 993 5427 1007 5441
rect 1013 5439 1027 5453
rect 1033 5427 1047 5441
rect 933 5393 947 5407
rect 1053 5419 1067 5433
rect 1113 5419 1127 5433
rect 1133 5427 1147 5441
rect 1393 5476 1407 5490
rect 1153 5419 1167 5433
rect 1233 5447 1247 5461
rect 1173 5427 1187 5441
rect 1193 5419 1207 5433
rect 973 5393 987 5407
rect 1013 5393 1027 5407
rect 1253 5382 1267 5396
rect 1313 5419 1327 5433
rect 1353 5419 1367 5433
rect 1613 5433 1627 5447
rect 1653 5433 1667 5447
rect 1673 5427 1687 5441
rect 1693 5439 1707 5453
rect 1473 5407 1487 5421
rect 1253 5344 1267 5358
rect 1393 5350 1407 5364
rect 1493 5399 1507 5413
rect 1533 5399 1547 5413
rect 1573 5407 1587 5421
rect 1513 5379 1527 5393
rect 1593 5399 1607 5413
rect 1633 5399 1647 5413
rect 1613 5379 1627 5393
rect 1693 5393 1707 5407
rect 1733 5433 1747 5447
rect 1753 5419 1767 5433
rect 1773 5427 1787 5441
rect 1793 5419 1807 5433
rect 1833 5419 1847 5433
rect 1733 5399 1747 5413
rect 1853 5407 1867 5421
rect 1713 5296 1727 5307
rect 1893 5419 1907 5433
rect 1933 5407 1947 5421
rect 1953 5399 1967 5413
rect 1973 5407 1987 5421
rect 2033 5419 2047 5433
rect 2053 5427 2067 5441
rect 2073 5419 2087 5433
rect 2013 5399 2027 5413
rect 2093 5407 2107 5421
rect 2193 5427 2207 5441
rect 2213 5439 2227 5453
rect 2113 5399 2127 5413
rect 2133 5407 2147 5421
rect 2273 5419 2287 5433
rect 2293 5427 2307 5441
rect 2353 5439 2367 5453
rect 2313 5419 2327 5433
rect 2333 5419 2347 5433
rect 2253 5399 2267 5413
rect 2373 5419 2387 5433
rect 2433 5427 2447 5441
rect 2453 5439 2467 5453
rect 2493 5419 2507 5433
rect 2513 5427 2527 5441
rect 2533 5439 2547 5453
rect 2553 5427 2567 5441
rect 2573 5419 2587 5433
rect 2593 5427 2607 5441
rect 2613 5419 2627 5433
rect 2633 5399 2647 5413
rect 2673 5407 2687 5421
rect 2693 5399 2707 5413
rect 2713 5407 2727 5421
rect 2773 5407 2787 5421
rect 2793 5399 2807 5413
rect 2833 5399 2847 5413
rect 2873 5407 2887 5421
rect 2973 5439 2987 5453
rect 2893 5399 2907 5413
rect 2913 5407 2927 5421
rect 2953 5419 2967 5433
rect 2813 5379 2827 5393
rect 2993 5419 3007 5433
rect 3013 5419 3027 5433
rect 3033 5427 3047 5441
rect 3053 5419 3067 5433
rect 3073 5399 3087 5413
rect 3133 5407 3147 5421
rect 3153 5399 3167 5413
rect 3173 5407 3187 5421
rect 3193 5419 3207 5433
rect 3213 5427 3227 5441
rect 3233 5419 3247 5433
rect 3313 5419 3327 5433
rect 2933 5296 2947 5307
rect 3253 5399 3267 5413
rect 3333 5407 3347 5421
rect 3413 5439 3427 5453
rect 3473 5439 3487 5453
rect 3373 5419 3387 5433
rect 3393 5419 3407 5433
rect 3433 5419 3447 5433
rect 3493 5419 3507 5433
rect 3533 5427 3547 5441
rect 3573 5419 3587 5433
rect 3593 5427 3607 5441
rect 3713 5439 3727 5453
rect 3613 5419 3627 5433
rect 3693 5419 3707 5433
rect 3633 5399 3647 5413
rect 3733 5419 3747 5433
rect 3753 5419 3767 5433
rect 3773 5427 3787 5441
rect 3793 5419 3807 5433
rect 3813 5427 3827 5441
rect 3913 5439 3927 5453
rect 3833 5419 3847 5433
rect 3893 5419 3907 5433
rect 3933 5419 3947 5433
rect 3953 5419 3967 5433
rect 3973 5427 3987 5441
rect 3993 5419 4007 5433
rect 4013 5399 4027 5413
rect 4073 5407 4087 5421
rect 4093 5399 4107 5413
rect 4133 5399 4147 5413
rect 4173 5407 4187 5421
rect 4233 5439 4247 5453
rect 4253 5427 4267 5441
rect 4193 5399 4207 5413
rect 4213 5407 4227 5421
rect 4113 5379 4127 5393
rect 4333 5419 4347 5433
rect 4353 5427 4367 5441
rect 4373 5419 4387 5433
rect 4313 5399 4327 5413
rect 4413 5407 4427 5421
rect 4433 5399 4447 5413
rect 4453 5407 4467 5421
rect 4473 5407 4487 5421
rect 4493 5399 4507 5413
rect 4513 5407 4527 5421
rect 4573 5433 4587 5447
rect 4593 5419 4607 5433
rect 4613 5427 4627 5441
rect 4653 5433 4667 5447
rect 4633 5419 4647 5433
rect 4573 5399 4587 5413
rect 4693 5419 4707 5433
rect 4713 5427 4727 5441
rect 4733 5419 4747 5433
rect 4773 5419 4787 5433
rect 4673 5399 4687 5413
rect 4573 5353 4587 5367
rect 4653 5373 4667 5387
rect 4793 5407 4807 5421
rect 4833 5419 4847 5433
rect 4893 5419 4907 5433
rect 4913 5427 4927 5441
rect 4933 5419 4947 5433
rect 4873 5399 4887 5413
rect 4973 5407 4987 5421
rect 4993 5399 5007 5413
rect 5013 5407 5027 5421
rect 5053 5419 5067 5433
rect 5073 5407 5087 5421
rect 5113 5419 5127 5433
rect 5133 5407 5147 5421
rect 5153 5399 5167 5413
rect 5173 5407 5187 5421
rect 5213 5419 5227 5433
rect 5233 5427 5247 5441
rect 5253 5419 5267 5433
rect 5333 5419 5347 5433
rect 5273 5399 5287 5413
rect 5353 5407 5367 5421
rect 5393 5419 5407 5433
rect 5413 5419 5427 5433
rect 5433 5427 5447 5441
rect 5473 5433 5487 5447
rect 5453 5419 5467 5433
rect 5473 5399 5487 5413
rect 5473 5353 5487 5367
rect 5513 5407 5527 5421
rect 5533 5399 5547 5413
rect 5553 5407 5567 5421
rect 5613 5433 5627 5447
rect 5593 5399 5607 5413
rect 5633 5399 5647 5413
rect 5653 5407 5667 5421
rect 5713 5419 5727 5433
rect 5613 5379 5627 5393
rect 5573 5353 5587 5367
rect 5733 5407 5747 5421
rect 5773 5419 5787 5433
rect 5813 5419 5827 5433
rect 5833 5427 5847 5441
rect 5853 5419 5867 5433
rect 5873 5427 5887 5441
rect 5893 5419 5907 5433
rect 5913 5407 5927 5421
rect 6093 5427 6107 5441
rect 6113 5439 6127 5453
rect 6133 5427 6147 5441
rect 5933 5399 5947 5413
rect 5953 5407 5967 5421
rect 5993 5399 6007 5413
rect 6033 5399 6047 5413
rect 6053 5407 6067 5421
rect 6153 5419 6167 5433
rect 6233 5419 6247 5433
rect 6253 5427 6267 5441
rect 6273 5419 6287 5433
rect 6293 5419 6307 5433
rect 6313 5427 6327 5441
rect 6333 5419 6347 5433
rect 6013 5379 6027 5393
rect 6213 5399 6227 5413
rect 6353 5399 6367 5413
rect 6353 5353 6367 5367
rect 6413 5433 6427 5447
rect 6393 5413 6407 5427
rect 6433 5419 6447 5433
rect 6453 5427 6467 5441
rect 6473 5419 6487 5433
rect 6553 5433 6567 5447
rect 6573 5433 6587 5447
rect 6413 5399 6427 5413
rect 6513 5407 6527 5421
rect 6613 5419 6627 5433
rect 6633 5427 6647 5441
rect 6653 5439 6667 5453
rect 6673 5427 6687 5441
rect 6413 5353 6427 5367
rect 6533 5399 6547 5413
rect 6573 5399 6587 5413
rect 6553 5379 6567 5393
rect 1713 5293 1727 5296
rect 2933 5293 2947 5296
rect 1013 5284 1027 5287
rect 3673 5284 3687 5287
rect 4113 5284 4127 5287
rect 133 5222 147 5236
rect 273 5216 287 5230
rect 33 5147 47 5161
rect 73 5147 87 5161
rect 133 5184 147 5198
rect 113 5119 127 5133
rect 193 5147 207 5161
rect 233 5147 247 5161
rect 133 5090 147 5104
rect 333 5159 347 5173
rect 353 5167 367 5181
rect 373 5159 387 5173
rect 633 5216 647 5230
rect 773 5222 787 5236
rect 433 5147 447 5161
rect 533 5159 547 5173
rect 553 5167 567 5181
rect 273 5090 287 5104
rect 453 5139 467 5153
rect 473 5127 487 5141
rect 493 5139 507 5153
rect 573 5159 587 5173
rect 673 5147 687 5161
rect 713 5147 727 5161
rect 773 5184 787 5198
rect 1013 5273 1027 5284
rect 833 5159 847 5173
rect 853 5167 867 5181
rect 793 5119 807 5133
rect 633 5090 647 5104
rect 873 5159 887 5173
rect 933 5167 947 5181
rect 1033 5167 1047 5181
rect 953 5147 967 5161
rect 973 5139 987 5153
rect 993 5147 1007 5161
rect 1053 5147 1067 5161
rect 1073 5139 1087 5153
rect 1093 5147 1107 5161
rect 1133 5147 1147 5161
rect 1153 5159 1167 5173
rect 773 5090 787 5104
rect 1253 5222 1267 5236
rect 1393 5216 1407 5230
rect 1193 5147 1207 5161
rect 1253 5184 1267 5198
rect 1233 5119 1247 5133
rect 1313 5147 1327 5161
rect 1353 5147 1367 5161
rect 1253 5090 1267 5104
rect 1653 5222 1667 5236
rect 1793 5216 1807 5230
rect 1473 5159 1487 5173
rect 1493 5167 1507 5181
rect 1513 5159 1527 5173
rect 1533 5159 1547 5173
rect 1553 5167 1567 5181
rect 1393 5090 1407 5104
rect 1573 5159 1587 5173
rect 1653 5184 1667 5198
rect 1633 5119 1647 5133
rect 1713 5147 1727 5161
rect 1753 5147 1767 5161
rect 1653 5090 1667 5104
rect 1873 5147 1887 5161
rect 1893 5139 1907 5153
rect 1913 5147 1927 5161
rect 1933 5139 1947 5153
rect 1953 5147 1967 5161
rect 1973 5127 1987 5141
rect 1993 5139 2007 5153
rect 2053 5147 2067 5161
rect 2073 5159 2087 5173
rect 1793 5090 1807 5104
rect 2113 5147 2127 5161
rect 2133 5159 2147 5173
rect 2153 5167 2167 5181
rect 2173 5159 2187 5173
rect 2233 5139 2247 5153
rect 2273 5147 2287 5161
rect 2333 5159 2347 5173
rect 2353 5167 2367 5181
rect 2453 5187 2467 5201
rect 2293 5127 2307 5141
rect 2373 5159 2387 5173
rect 2413 5159 2427 5173
rect 2433 5167 2447 5181
rect 2473 5167 2487 5181
rect 2513 5147 2527 5161
rect 2553 5147 2567 5161
rect 2533 5127 2547 5141
rect 2573 5127 2587 5141
rect 2593 5139 2607 5153
rect 2653 5147 2667 5161
rect 2673 5159 2687 5173
rect 2713 5147 2727 5161
rect 2733 5147 2747 5161
rect 2773 5147 2787 5161
rect 2833 5159 2847 5173
rect 2853 5167 2867 5181
rect 2753 5127 2767 5141
rect 2873 5159 2887 5173
rect 2913 5159 2927 5173
rect 2933 5167 2947 5181
rect 2953 5159 2967 5173
rect 2993 5147 3007 5161
rect 2973 5127 2987 5141
rect 3033 5139 3047 5153
rect 3093 5147 3107 5161
rect 3113 5159 3127 5173
rect 3153 5147 3167 5161
rect 3173 5159 3187 5173
rect 3193 5167 3207 5181
rect 3313 5187 3327 5201
rect 3213 5159 3227 5173
rect 3273 5159 3287 5173
rect 3293 5167 3307 5181
rect 3333 5167 3347 5181
rect 3673 5273 3687 5284
rect 3653 5213 3667 5227
rect 3373 5139 3387 5153
rect 3433 5147 3447 5161
rect 3393 5127 3407 5141
rect 3453 5139 3467 5153
rect 3473 5127 3487 5141
rect 3493 5139 3507 5153
rect 3533 5147 3547 5161
rect 3653 5167 3667 5181
rect 3573 5147 3587 5161
rect 3593 5147 3607 5161
rect 3553 5127 3567 5141
rect 3613 5139 3627 5153
rect 3633 5147 3647 5161
rect 3653 5133 3667 5147
rect 3713 5167 3727 5181
rect 3733 5147 3747 5161
rect 3753 5139 3767 5153
rect 3773 5147 3787 5161
rect 3793 5147 3807 5161
rect 3833 5147 3847 5161
rect 3813 5127 3827 5141
rect 3873 5193 3887 5207
rect 3913 5193 3927 5207
rect 3873 5159 3887 5173
rect 3893 5167 3907 5181
rect 3873 5113 3887 5127
rect 3913 5159 3927 5173
rect 4113 5273 4127 5284
rect 4093 5213 4107 5227
rect 4153 5213 4167 5227
rect 3973 5159 3987 5173
rect 3993 5167 4007 5181
rect 4013 5159 4027 5173
rect 4093 5167 4107 5181
rect 4033 5147 4047 5161
rect 4053 5139 4067 5153
rect 4073 5147 4087 5161
rect 4153 5159 4167 5173
rect 4173 5167 4187 5181
rect 4193 5159 4207 5173
rect 4233 5147 4247 5161
rect 4253 5159 4267 5173
rect 3953 5073 3967 5087
rect 4293 5193 4307 5207
rect 4333 5193 4347 5207
rect 4293 5147 4307 5161
rect 4333 5159 4347 5173
rect 4353 5167 4367 5181
rect 4373 5159 4387 5173
rect 4413 5167 4427 5181
rect 4433 5147 4447 5161
rect 4453 5139 4467 5153
rect 4473 5147 4487 5161
rect 4513 5213 4527 5227
rect 4513 5167 4527 5181
rect 4633 5193 4647 5207
rect 4533 5147 4547 5161
rect 4513 5133 4527 5147
rect 4553 5139 4567 5153
rect 4573 5147 4587 5161
rect 4593 5159 4607 5173
rect 4613 5167 4627 5181
rect 4633 5159 4647 5173
rect 4713 5193 4727 5207
rect 4753 5193 4767 5207
rect 4673 5159 4687 5173
rect 4693 5167 4707 5181
rect 4653 5113 4667 5127
rect 4713 5159 4727 5173
rect 4753 5173 4767 5187
rect 4793 5193 4807 5207
rect 4733 5133 4747 5147
rect 4753 5127 4767 5141
rect 4773 5139 4787 5153
rect 4873 5187 4887 5201
rect 4973 5213 4987 5227
rect 4813 5153 4827 5167
rect 4833 5159 4847 5173
rect 4853 5167 4867 5181
rect 4893 5167 4907 5181
rect 4973 5167 4987 5181
rect 4913 5147 4927 5161
rect 4933 5139 4947 5153
rect 4953 5147 4967 5161
rect 4793 5113 4807 5127
rect 4813 5113 4827 5127
rect 4973 5133 4987 5147
rect 5013 5139 5027 5153
rect 5033 5147 5047 5161
rect 5073 5159 5087 5173
rect 5093 5167 5107 5181
rect 5113 5159 5127 5173
rect 5273 5213 5287 5227
rect 5233 5159 5247 5173
rect 5253 5167 5267 5181
rect 5153 5139 5167 5153
rect 5193 5139 5207 5153
rect 5273 5159 5287 5173
rect 5433 5187 5447 5201
rect 5373 5167 5387 5181
rect 5413 5167 5427 5181
rect 5453 5167 5467 5181
rect 5493 5193 5507 5207
rect 5313 5147 5327 5161
rect 5333 5139 5347 5153
rect 5353 5147 5367 5161
rect 5473 5159 5487 5173
rect 5313 5113 5327 5127
rect 5373 5133 5387 5147
rect 5413 5133 5427 5147
rect 5533 5187 5547 5201
rect 5513 5167 5527 5181
rect 5553 5167 5567 5181
rect 5573 5159 5587 5173
rect 5533 5133 5547 5147
rect 5573 5093 5587 5107
rect 5613 5173 5627 5187
rect 5693 5187 5707 5201
rect 5673 5167 5687 5181
rect 5713 5167 5727 5181
rect 5733 5159 5747 5173
rect 5833 5167 5847 5181
rect 5853 5173 5867 5187
rect 5973 5187 5987 5201
rect 5613 5127 5627 5141
rect 5633 5139 5647 5153
rect 5773 5147 5787 5161
rect 5793 5139 5807 5153
rect 5813 5147 5827 5161
rect 5833 5133 5847 5147
rect 5893 5159 5907 5173
rect 5913 5167 5927 5181
rect 5933 5159 5947 5173
rect 5953 5167 5967 5181
rect 5993 5167 6007 5181
rect 6093 5193 6107 5207
rect 6013 5159 6027 5173
rect 6053 5159 6067 5173
rect 6073 5167 6087 5181
rect 6093 5159 6107 5173
rect 6193 5173 6207 5187
rect 6153 5147 6167 5161
rect 6113 5093 6127 5107
rect 6173 5139 6187 5153
rect 6193 5127 6207 5141
rect 6213 5139 6227 5153
rect 6273 5173 6287 5187
rect 6253 5139 6267 5153
rect 6233 5113 6247 5127
rect 6273 5127 6287 5141
rect 6273 5093 6287 5107
rect 6373 5213 6387 5227
rect 6353 5187 6367 5201
rect 6313 5159 6327 5173
rect 6333 5167 6347 5181
rect 6373 5167 6387 5181
rect 6453 5187 6467 5201
rect 6393 5153 6407 5167
rect 6413 5159 6427 5173
rect 6433 5167 6447 5181
rect 6473 5167 6487 5181
rect 6553 5213 6567 5227
rect 6493 5127 6507 5141
rect 6513 5139 6527 5153
rect 6613 5187 6627 5201
rect 6713 5193 6727 5207
rect 6573 5159 6587 5173
rect 6593 5167 6607 5181
rect 6633 5167 6647 5181
rect 6653 5159 6667 5173
rect 6673 5167 6687 5181
rect 6573 5093 6587 5107
rect 6693 5159 6707 5173
rect 6713 5113 6727 5127
rect 33 4939 47 4953
rect 293 4996 307 5010
rect 73 4939 87 4953
rect 113 4939 127 4953
rect 153 4939 167 4953
rect 193 4927 207 4941
rect 433 4996 447 5010
rect 273 4967 287 4981
rect 213 4919 227 4933
rect 233 4927 247 4941
rect 293 4902 307 4916
rect 353 4939 367 4953
rect 393 4939 407 4953
rect 513 4939 527 4953
rect 533 4947 547 4961
rect 553 4959 567 4973
rect 573 4947 587 4961
rect 613 4927 627 4941
rect 873 4996 887 5010
rect 553 4913 567 4927
rect 633 4919 647 4933
rect 653 4927 667 4941
rect 673 4927 687 4941
rect 733 4953 747 4967
rect 693 4919 707 4933
rect 713 4927 727 4941
rect 293 4864 307 4878
rect 433 4870 447 4884
rect 613 4893 627 4907
rect 773 4927 787 4941
rect 1013 4996 1027 5010
rect 853 4967 867 4981
rect 793 4919 807 4933
rect 813 4927 827 4941
rect 733 4873 747 4887
rect 873 4902 887 4916
rect 933 4939 947 4953
rect 973 4939 987 4953
rect 1093 4939 1107 4953
rect 1253 4993 1267 5007
rect 1133 4939 1147 4953
rect 1173 4939 1187 4953
rect 1193 4947 1207 4961
rect 1213 4959 1227 4973
rect 1233 4947 1247 4961
rect 873 4864 887 4878
rect 1013 4870 1027 4884
rect 1213 4913 1227 4927
rect 1273 4927 1287 4941
rect 1293 4919 1307 4933
rect 1313 4927 1327 4941
rect 1353 4939 1367 4953
rect 1393 4939 1407 4953
rect 1413 4927 1427 4941
rect 1433 4919 1447 4933
rect 1453 4927 1467 4941
rect 1513 4927 1527 4941
rect 1673 4993 1687 5007
rect 1533 4919 1547 4933
rect 1553 4927 1567 4941
rect 1613 4939 1627 4953
rect 1633 4947 1647 4961
rect 1653 4939 1667 4953
rect 1593 4919 1607 4933
rect 1693 4927 1707 4941
rect 1713 4919 1727 4933
rect 1733 4927 1747 4941
rect 1793 4939 1807 4953
rect 1813 4947 1827 4961
rect 1833 4939 1847 4953
rect 1773 4919 1787 4933
rect 1673 4893 1687 4907
rect 1853 4927 1867 4941
rect 1873 4919 1887 4933
rect 1893 4927 1907 4941
rect 1973 4939 1987 4953
rect 1993 4947 2007 4961
rect 2033 4953 2047 4967
rect 2013 4939 2027 4953
rect 1913 4913 1927 4927
rect 1953 4919 1967 4933
rect 1893 4893 1907 4907
rect 2073 4939 2087 4953
rect 2093 4947 2107 4961
rect 2113 4939 2127 4953
rect 2153 4939 2167 4953
rect 2053 4919 2067 4933
rect 2173 4927 2187 4941
rect 2053 4873 2067 4887
rect 2033 4816 2047 4827
rect 2233 4959 2247 4973
rect 2213 4939 2227 4953
rect 2253 4947 2267 4961
rect 2333 4959 2347 4973
rect 2313 4939 2327 4953
rect 2353 4939 2367 4953
rect 2393 4947 2407 4961
rect 2453 4959 2467 4973
rect 2433 4939 2447 4953
rect 2493 4927 2507 4941
rect 2513 4919 2527 4933
rect 2533 4927 2547 4941
rect 2593 4939 2607 4953
rect 2613 4947 2627 4961
rect 2633 4939 2647 4953
rect 2693 4939 2707 4953
rect 2713 4947 2727 4961
rect 2733 4939 2747 4953
rect 2773 4947 2787 4961
rect 2793 4959 2807 4973
rect 2573 4919 2587 4933
rect 2673 4919 2687 4933
rect 2553 4816 2567 4827
rect 2813 4939 2827 4953
rect 2833 4947 2847 4961
rect 2853 4939 2867 4953
rect 2953 4939 2967 4953
rect 2973 4947 2987 4961
rect 2993 4939 3007 4953
rect 3053 4939 3067 4953
rect 3073 4947 3087 4961
rect 3153 4959 3167 4973
rect 3093 4939 3107 4953
rect 3133 4939 3147 4953
rect 2873 4919 2887 4933
rect 2933 4919 2947 4933
rect 3033 4919 3047 4933
rect 3173 4939 3187 4953
rect 3213 4939 3227 4953
rect 3233 4947 3247 4961
rect 3273 4927 3287 4941
rect 3473 4996 3487 5010
rect 3293 4919 3307 4933
rect 3313 4927 3327 4941
rect 3373 4939 3387 4953
rect 3393 4947 3407 4961
rect 3413 4939 3427 4953
rect 3353 4919 3367 4933
rect 2913 4816 2927 4827
rect 3613 4996 3627 5010
rect 3513 4939 3527 4953
rect 3553 4939 3567 4953
rect 3633 4967 3647 4981
rect 3613 4902 3627 4916
rect 3673 4939 3687 4953
rect 3693 4947 3707 4961
rect 3713 4939 3727 4953
rect 3793 4939 3807 4953
rect 3813 4947 3827 4961
rect 3833 4959 3847 4973
rect 3853 4947 3867 4961
rect 3733 4919 3747 4933
rect 3833 4913 3847 4927
rect 3893 4993 3907 5007
rect 3893 4927 3907 4941
rect 3993 4939 4007 4953
rect 4013 4947 4027 4961
rect 4033 4959 4047 4973
rect 4053 4947 4067 4961
rect 4093 4939 4107 4953
rect 4113 4947 4127 4961
rect 4153 4939 4167 4953
rect 3473 4870 3487 4884
rect 3613 4864 3627 4878
rect 3913 4919 3927 4933
rect 3953 4919 3967 4933
rect 3933 4899 3947 4913
rect 4013 4913 4027 4927
rect 4073 4913 4087 4927
rect 4173 4927 4187 4941
rect 4213 4939 4227 4953
rect 4253 4927 4267 4941
rect 4273 4919 4287 4933
rect 4293 4927 4307 4941
rect 4313 4939 4327 4953
rect 4353 4927 4367 4941
rect 4373 4939 4387 4953
rect 4453 4939 4467 4953
rect 4473 4947 4487 4961
rect 4493 4939 4507 4953
rect 4433 4919 4447 4933
rect 4513 4919 4527 4933
rect 4553 4919 4567 4933
rect 4573 4927 4587 4941
rect 4613 4939 4627 4953
rect 4633 4947 4647 4961
rect 4673 4953 4687 4967
rect 4653 4939 4667 4953
rect 4413 4816 4427 4827
rect 4533 4899 4547 4913
rect 4673 4919 4687 4933
rect 4673 4873 4687 4887
rect 4733 4927 4747 4941
rect 4713 4913 4727 4927
rect 4753 4919 4767 4933
rect 4773 4927 4787 4941
rect 4813 4939 4827 4953
rect 4733 4893 4747 4907
rect 4833 4927 4847 4941
rect 4893 4973 4907 4987
rect 4873 4939 4887 4953
rect 4913 4927 4927 4941
rect 4933 4919 4947 4933
rect 4953 4927 4967 4941
rect 4973 4927 4987 4941
rect 4993 4919 5007 4933
rect 5013 4927 5027 4941
rect 5053 4939 5067 4953
rect 4913 4893 4927 4907
rect 5093 4927 5107 4941
rect 5113 4939 5127 4953
rect 5173 4927 5187 4941
rect 5193 4919 5207 4933
rect 5213 4927 5227 4941
rect 5253 4939 5267 4953
rect 5273 4927 5287 4941
rect 5313 4939 5327 4953
rect 5333 4939 5347 4953
rect 5373 4927 5387 4941
rect 5393 4939 5407 4953
rect 5453 4939 5467 4953
rect 5473 4947 5487 4961
rect 5493 4939 5507 4953
rect 5513 4947 5527 4961
rect 5533 4939 5547 4953
rect 5573 4927 5587 4941
rect 5593 4919 5607 4933
rect 5613 4927 5627 4941
rect 5633 4919 5647 4933
rect 5673 4919 5687 4933
rect 5693 4927 5707 4941
rect 5753 4939 5767 4953
rect 5773 4947 5787 4961
rect 5793 4959 5807 4973
rect 5813 4947 5827 4961
rect 5653 4899 5667 4913
rect 5773 4913 5787 4927
rect 5853 4993 5867 5007
rect 5913 4953 5927 4967
rect 5853 4927 5867 4941
rect 5873 4919 5887 4933
rect 5913 4919 5927 4933
rect 5893 4899 5907 4913
rect 5913 4873 5927 4887
rect 5953 4927 5967 4941
rect 5973 4919 5987 4933
rect 5993 4927 6007 4941
rect 6013 4939 6027 4953
rect 6033 4947 6047 4961
rect 6053 4939 6067 4953
rect 6073 4947 6087 4961
rect 6093 4939 6107 4953
rect 6153 4993 6167 5007
rect 6153 4927 6167 4941
rect 6233 4939 6247 4953
rect 6253 4947 6267 4961
rect 6273 4939 6287 4953
rect 6613 4993 6627 5007
rect 6133 4893 6147 4907
rect 6173 4919 6187 4933
rect 6213 4919 6227 4933
rect 6193 4899 6207 4913
rect 6293 4919 6307 4933
rect 6353 4927 6367 4941
rect 6293 4873 6307 4887
rect 6333 4913 6347 4927
rect 6373 4919 6387 4933
rect 6413 4919 6427 4933
rect 6453 4927 6467 4941
rect 6393 4899 6407 4913
rect 6473 4919 6487 4933
rect 6513 4919 6527 4933
rect 6533 4927 6547 4941
rect 6553 4919 6567 4933
rect 6573 4927 6587 4941
rect 6633 4947 6647 4961
rect 6653 4959 6667 4973
rect 6493 4899 6507 4913
rect 6613 4913 6627 4927
rect 2033 4813 2047 4816
rect 2553 4813 2567 4816
rect 2913 4813 2927 4816
rect 4413 4813 4427 4816
rect 1673 4804 1687 4807
rect 1813 4804 1827 4807
rect 3733 4804 3747 4807
rect 33 4659 47 4673
rect 173 4659 187 4673
rect 233 4667 247 4681
rect 273 4667 287 4681
rect 253 4647 267 4661
rect 313 4659 327 4673
rect 373 4667 387 4681
rect 333 4647 347 4661
rect 353 4653 367 4667
rect 333 4613 347 4627
rect 393 4659 407 4673
rect 413 4647 427 4661
rect 433 4659 447 4673
rect 473 4659 487 4673
rect 533 4667 547 4681
rect 573 4667 587 4681
rect 613 4667 627 4681
rect 633 4679 647 4693
rect 493 4647 507 4661
rect 553 4647 567 4661
rect 673 4667 687 4681
rect 693 4667 707 4681
rect 973 4742 987 4756
rect 1113 4736 1127 4750
rect 733 4667 747 4681
rect 793 4667 807 4681
rect 713 4647 727 4661
rect 833 4667 847 4681
rect 873 4679 887 4693
rect 893 4687 907 4701
rect 913 4679 927 4693
rect 973 4704 987 4718
rect 953 4639 967 4653
rect 1033 4667 1047 4681
rect 1073 4667 1087 4681
rect 973 4610 987 4624
rect 1193 4687 1207 4701
rect 1393 4733 1407 4747
rect 1433 4733 1447 4747
rect 1393 4713 1407 4727
rect 1213 4667 1227 4681
rect 1233 4659 1247 4673
rect 1253 4667 1267 4681
rect 1293 4679 1307 4693
rect 1313 4687 1327 4701
rect 1333 4679 1347 4693
rect 1353 4679 1367 4693
rect 1373 4687 1387 4701
rect 1393 4679 1407 4693
rect 1673 4793 1687 4804
rect 1453 4687 1467 4701
rect 1473 4667 1487 4681
rect 1433 4653 1447 4667
rect 1493 4659 1507 4673
rect 1513 4667 1527 4681
rect 1533 4667 1547 4681
rect 1573 4667 1587 4681
rect 1613 4667 1627 4681
rect 1653 4667 1667 4681
rect 1733 4713 1747 4727
rect 1813 4793 1827 4804
rect 1973 4742 1987 4756
rect 2113 4736 2127 4750
rect 1553 4647 1567 4661
rect 1633 4647 1647 4661
rect 1693 4647 1707 4661
rect 1713 4659 1727 4673
rect 1113 4610 1127 4624
rect 1753 4667 1767 4681
rect 1813 4693 1827 4707
rect 1793 4667 1807 4681
rect 1773 4647 1787 4661
rect 1753 4633 1767 4647
rect 1893 4687 1907 4701
rect 1833 4667 1847 4681
rect 1853 4659 1867 4673
rect 1873 4667 1887 4681
rect 1973 4704 1987 4718
rect 1813 4613 1827 4627
rect 1953 4639 1967 4653
rect 2033 4667 2047 4681
rect 2073 4667 2087 4681
rect 1973 4610 1987 4624
rect 2193 4679 2207 4693
rect 2213 4687 2227 4701
rect 2233 4679 2247 4693
rect 2113 4610 2127 4624
rect 2273 4659 2287 4673
rect 2313 4667 2327 4681
rect 2353 4679 2367 4693
rect 2373 4687 2387 4701
rect 2333 4647 2347 4661
rect 2393 4679 2407 4693
rect 2433 4667 2447 4681
rect 2493 4693 2507 4707
rect 2553 4693 2567 4707
rect 2473 4667 2487 4681
rect 2453 4647 2467 4661
rect 2513 4659 2527 4673
rect 2533 4647 2547 4661
rect 2553 4659 2567 4673
rect 2573 4667 2587 4681
rect 2713 4742 2727 4756
rect 2853 4736 2867 4750
rect 2633 4659 2647 4673
rect 2653 4647 2667 4661
rect 2713 4704 2727 4718
rect 2693 4639 2707 4653
rect 3053 4742 3067 4756
rect 3193 4736 3207 4750
rect 2773 4667 2787 4681
rect 2813 4667 2827 4681
rect 2713 4610 2727 4624
rect 2973 4687 2987 4701
rect 2913 4667 2927 4681
rect 2933 4659 2947 4673
rect 2953 4667 2967 4681
rect 3053 4704 3067 4718
rect 2853 4610 2867 4624
rect 3033 4639 3047 4653
rect 3113 4667 3127 4681
rect 3153 4667 3167 4681
rect 3053 4610 3067 4624
rect 3193 4610 3207 4624
rect 3293 4742 3307 4756
rect 3433 4736 3447 4750
rect 3293 4704 3307 4718
rect 3273 4639 3287 4653
rect 3733 4793 3747 4804
rect 3353 4667 3367 4681
rect 3393 4667 3407 4681
rect 3293 4610 3307 4624
rect 3513 4687 3527 4701
rect 3713 4713 3727 4727
rect 3533 4667 3547 4681
rect 3553 4659 3567 4673
rect 3573 4667 3587 4681
rect 3613 4667 3627 4681
rect 3673 4679 3687 4693
rect 3693 4687 3707 4701
rect 3433 4610 3447 4624
rect 3633 4659 3647 4673
rect 3713 4679 3727 4693
rect 3713 4633 3727 4647
rect 3873 4736 3887 4750
rect 4013 4742 4027 4756
rect 3753 4687 3767 4701
rect 3773 4667 3787 4681
rect 3793 4659 3807 4673
rect 3813 4667 3827 4681
rect 3913 4667 3927 4681
rect 3953 4667 3967 4681
rect 4013 4704 4027 4718
rect 4253 4742 4267 4756
rect 4393 4736 4407 4750
rect 4093 4667 4107 4681
rect 4153 4679 4167 4693
rect 4173 4687 4187 4701
rect 4033 4639 4047 4653
rect 3873 4610 3887 4624
rect 4113 4659 4127 4673
rect 4193 4679 4207 4693
rect 4253 4704 4267 4718
rect 4233 4639 4247 4653
rect 4313 4667 4327 4681
rect 4353 4667 4367 4681
rect 4013 4610 4027 4624
rect 4253 4610 4267 4624
rect 4513 4707 4527 4721
rect 4473 4679 4487 4693
rect 4493 4687 4507 4701
rect 4533 4687 4547 4701
rect 4553 4647 4567 4661
rect 4573 4659 4587 4673
rect 4613 4659 4627 4673
rect 4633 4667 4647 4681
rect 4793 4687 4807 4701
rect 4393 4610 4407 4624
rect 4693 4659 4707 4673
rect 4733 4667 4747 4681
rect 4713 4647 4727 4661
rect 4753 4659 4767 4673
rect 4773 4667 4787 4681
rect 4833 4667 4847 4681
rect 4953 4713 4967 4727
rect 4873 4667 4887 4681
rect 4913 4679 4927 4693
rect 4933 4687 4947 4701
rect 4853 4647 4867 4661
rect 4953 4679 4967 4693
rect 5033 4733 5047 4747
rect 5073 4733 5087 4747
rect 4973 4673 4987 4687
rect 4993 4679 5007 4693
rect 5013 4687 5027 4701
rect 5033 4679 5047 4693
rect 5053 4673 5067 4687
rect 5093 4713 5107 4727
rect 5093 4679 5107 4693
rect 5113 4687 5127 4701
rect 5133 4679 5147 4693
rect 5213 4687 5227 4701
rect 5413 4733 5427 4747
rect 5473 4733 5487 4747
rect 5153 4667 5167 4681
rect 5173 4659 5187 4673
rect 5193 4667 5207 4681
rect 5273 4667 5287 4681
rect 5293 4659 5307 4673
rect 5313 4667 5327 4681
rect 5333 4659 5347 4673
rect 5353 4667 5367 4681
rect 5373 4679 5387 4693
rect 5393 4687 5407 4701
rect 5413 4679 5427 4693
rect 5433 4633 5447 4647
rect 5473 4713 5487 4727
rect 5553 4707 5567 4721
rect 5473 4679 5487 4693
rect 5493 4687 5507 4701
rect 5513 4679 5527 4693
rect 5533 4687 5547 4701
rect 5573 4687 5587 4701
rect 5733 4707 5747 4721
rect 5593 4679 5607 4693
rect 5653 4679 5667 4693
rect 5673 4687 5687 4701
rect 5693 4679 5707 4693
rect 5713 4687 5727 4701
rect 5753 4687 5767 4701
rect 5773 4679 5787 4693
rect 5893 4707 5907 4721
rect 5873 4687 5887 4701
rect 5913 4687 5927 4701
rect 5933 4679 5947 4693
rect 5833 4659 5847 4673
rect 5853 4647 5867 4661
rect 5993 4667 6007 4681
rect 6013 4679 6027 4693
rect 6133 4733 6147 4747
rect 6133 4687 6147 4701
rect 6053 4667 6067 4681
rect 6073 4667 6087 4681
rect 6093 4659 6107 4673
rect 6113 4667 6127 4681
rect 6193 4679 6207 4693
rect 6213 4687 6227 4701
rect 6153 4653 6167 4667
rect 6233 4679 6247 4693
rect 6373 4707 6387 4721
rect 6353 4687 6367 4701
rect 6393 4687 6407 4701
rect 6253 4659 6267 4673
rect 6273 4647 6287 4661
rect 6293 4659 6307 4673
rect 6313 4667 6327 4681
rect 6413 4679 6427 4693
rect 6473 4667 6487 4681
rect 6493 4679 6507 4693
rect 6553 4733 6567 4747
rect 6533 4667 6547 4681
rect 6633 4733 6647 4747
rect 6613 4707 6627 4721
rect 6573 4679 6587 4693
rect 6593 4687 6607 4701
rect 6633 4687 6647 4701
rect 6673 4693 6687 4707
rect 6553 4633 6567 4647
rect 33 4467 47 4481
rect 53 4479 67 4493
rect 113 4479 127 4493
rect 93 4459 107 4473
rect 133 4459 147 4473
rect 173 4467 187 4481
rect 193 4479 207 4493
rect 213 4459 227 4473
rect 233 4467 247 4481
rect 353 4479 367 4493
rect 253 4459 267 4473
rect 333 4459 347 4473
rect 273 4439 287 4453
rect 373 4459 387 4473
rect 393 4459 407 4473
rect 413 4467 427 4481
rect 493 4479 507 4493
rect 433 4459 447 4473
rect 513 4459 527 4473
rect 453 4439 467 4453
rect 553 4467 567 4481
rect 593 4467 607 4481
rect 613 4479 627 4493
rect 633 4467 647 4481
rect 653 4459 667 4473
rect 713 4467 727 4481
rect 733 4479 747 4493
rect 773 4479 787 4493
rect 833 4479 847 4493
rect 753 4459 767 4473
rect 793 4459 807 4473
rect 853 4467 867 4481
rect 913 4479 927 4493
rect 973 4479 987 4493
rect 893 4459 907 4473
rect 933 4459 947 4473
rect 993 4467 1007 4481
rect 1053 4467 1067 4481
rect 1193 4467 1207 4481
rect 1233 4459 1247 4473
rect 1273 4459 1287 4473
rect 1333 4467 1347 4481
rect 1353 4479 1367 4493
rect 1353 4433 1367 4447
rect 1393 4493 1407 4507
rect 1773 4516 1787 4530
rect 1433 4493 1447 4507
rect 1413 4479 1427 4493
rect 1393 4459 1407 4473
rect 1433 4459 1447 4473
rect 1473 4447 1487 4461
rect 1493 4439 1507 4453
rect 1513 4447 1527 4461
rect 1533 4447 1547 4461
rect 1553 4439 1567 4453
rect 1573 4447 1587 4461
rect 1653 4459 1667 4473
rect 1693 4459 1707 4473
rect 1473 4413 1487 4427
rect 1913 4516 1927 4530
rect 1813 4459 1827 4473
rect 1853 4459 1867 4473
rect 1933 4487 1947 4501
rect 1913 4422 1927 4436
rect 2093 4516 2107 4530
rect 1973 4447 1987 4461
rect 2233 4516 2247 4530
rect 2073 4487 2087 4501
rect 1993 4439 2007 4453
rect 2013 4447 2027 4461
rect 1773 4390 1787 4404
rect 1913 4384 1927 4398
rect 2093 4422 2107 4436
rect 2153 4459 2167 4473
rect 2193 4459 2207 4473
rect 2293 4479 2307 4493
rect 2313 4467 2327 4481
rect 2373 4479 2387 4493
rect 2453 4479 2467 4493
rect 2513 4479 2527 4493
rect 2613 4516 2627 4530
rect 2753 4516 2767 4530
rect 2593 4487 2607 4501
rect 2093 4384 2107 4398
rect 2233 4390 2247 4404
rect 2353 4459 2367 4473
rect 2393 4459 2407 4473
rect 2433 4459 2447 4473
rect 2473 4459 2487 4473
rect 2533 4467 2547 4481
rect 2613 4422 2627 4436
rect 2673 4459 2687 4473
rect 2713 4459 2727 4473
rect 2813 4459 2827 4473
rect 2833 4467 2847 4481
rect 2853 4459 2867 4473
rect 2873 4439 2887 4453
rect 2913 4447 2927 4461
rect 3193 4516 3207 4530
rect 3333 4516 3347 4530
rect 3013 4467 3027 4481
rect 3033 4479 3047 4493
rect 2933 4439 2947 4453
rect 2953 4447 2967 4461
rect 2613 4384 2627 4398
rect 2753 4390 2767 4404
rect 3053 4459 3067 4473
rect 3073 4467 3087 4481
rect 3093 4459 3107 4473
rect 3173 4487 3187 4501
rect 3113 4439 3127 4453
rect 3193 4422 3207 4436
rect 3253 4459 3267 4473
rect 3293 4459 3307 4473
rect 3633 4516 3647 4530
rect 3393 4459 3407 4473
rect 3413 4467 3427 4481
rect 3433 4459 3447 4473
rect 3453 4439 3467 4453
rect 3193 4384 3207 4398
rect 3333 4390 3347 4404
rect 3513 4473 3527 4487
rect 3533 4459 3547 4473
rect 3553 4467 3567 4481
rect 3573 4459 3587 4473
rect 3513 4439 3527 4453
rect 3773 4516 3787 4530
rect 3973 4516 3987 4530
rect 3673 4459 3687 4473
rect 3713 4459 3727 4473
rect 3513 4393 3527 4407
rect 3493 4336 3507 4347
rect 3793 4487 3807 4501
rect 3773 4422 3787 4436
rect 3833 4459 3847 4473
rect 3853 4467 3867 4481
rect 3873 4459 3887 4473
rect 3893 4439 3907 4453
rect 4113 4516 4127 4530
rect 4013 4459 4027 4473
rect 4053 4459 4067 4473
rect 3633 4390 3647 4404
rect 3773 4384 3787 4398
rect 4133 4487 4147 4501
rect 4113 4422 4127 4436
rect 4193 4447 4207 4461
rect 4273 4459 4287 4473
rect 4293 4467 4307 4481
rect 4413 4479 4427 4493
rect 4313 4459 4327 4473
rect 4393 4459 4407 4473
rect 3973 4390 3987 4404
rect 4113 4384 4127 4398
rect 4213 4439 4227 4453
rect 4253 4439 4267 4453
rect 4233 4419 4247 4433
rect 4333 4439 4347 4453
rect 4433 4459 4447 4473
rect 4473 4459 4487 4473
rect 4493 4467 4507 4481
rect 4513 4479 4527 4493
rect 4533 4467 4547 4481
rect 4673 4467 4687 4481
rect 4693 4479 4707 4493
rect 4553 4439 4567 4453
rect 4593 4439 4607 4453
rect 4613 4447 4627 4461
rect 4373 4336 4387 4347
rect 4573 4419 4587 4433
rect 4713 4459 4727 4473
rect 4733 4467 4747 4481
rect 4753 4459 4767 4473
rect 4833 4467 4847 4481
rect 4773 4439 4787 4453
rect 4893 4479 4907 4493
rect 4873 4459 4887 4473
rect 4933 4447 4947 4461
rect 4953 4439 4967 4453
rect 4973 4447 4987 4461
rect 5013 4447 5027 4461
rect 5093 4459 5107 4473
rect 5113 4467 5127 4481
rect 5133 4459 5147 4473
rect 5213 4467 5227 4481
rect 5033 4439 5047 4453
rect 5073 4439 5087 4453
rect 5053 4419 5067 4433
rect 5153 4439 5167 4453
rect 5273 4479 5287 4493
rect 5253 4459 5267 4473
rect 5293 4459 5307 4473
rect 5313 4467 5327 4481
rect 5353 4473 5367 4487
rect 5393 4479 5407 4493
rect 5453 4533 5467 4547
rect 5333 4459 5347 4473
rect 5353 4439 5367 4453
rect 5413 4467 5427 4481
rect 5373 4413 5387 4427
rect 5473 4447 5487 4461
rect 5453 4393 5467 4407
rect 5493 4439 5507 4453
rect 5533 4439 5547 4453
rect 5553 4447 5567 4461
rect 5573 4439 5587 4453
rect 5593 4447 5607 4461
rect 5513 4419 5527 4433
rect 5633 4493 5647 4507
rect 5633 4459 5647 4473
rect 5653 4467 5667 4481
rect 5693 4473 5707 4487
rect 5673 4459 5687 4473
rect 5613 4413 5627 4427
rect 5693 4439 5707 4453
rect 5753 4447 5767 4461
rect 5873 4473 5887 4487
rect 5773 4439 5787 4453
rect 5793 4447 5807 4461
rect 5833 4447 5847 4461
rect 5753 4413 5767 4427
rect 5853 4439 5867 4453
rect 5893 4439 5907 4453
rect 5953 4459 5967 4473
rect 5973 4467 5987 4481
rect 6013 4479 6027 4493
rect 5993 4459 6007 4473
rect 6033 4467 6047 4481
rect 6093 4467 6107 4481
rect 6113 4479 6127 4493
rect 5873 4419 5887 4433
rect 5913 4433 5927 4447
rect 5933 4439 5947 4453
rect 6133 4439 6147 4453
rect 6173 4439 6187 4453
rect 6193 4447 6207 4461
rect 6273 4459 6287 4473
rect 6293 4467 6307 4481
rect 6313 4459 6327 4473
rect 6153 4419 6167 4433
rect 6253 4439 6267 4453
rect 6333 4439 6347 4453
rect 6373 4439 6387 4453
rect 6393 4447 6407 4461
rect 6353 4419 6367 4433
rect 6433 4473 6447 4487
rect 6433 4439 6447 4453
rect 6473 4439 6487 4453
rect 6493 4447 6507 4461
rect 6533 4459 6547 4473
rect 6553 4467 6567 4481
rect 6633 4479 6647 4493
rect 6573 4459 6587 4473
rect 6653 4467 6667 4481
rect 6453 4419 6467 4433
rect 6433 4393 6447 4407
rect 6593 4439 6607 4453
rect 3493 4333 3507 4336
rect 4373 4333 4387 4336
rect 93 4324 107 4327
rect 2733 4324 2747 4327
rect 2833 4324 2847 4327
rect 3053 4324 3067 4327
rect 4073 4324 4087 4327
rect 4513 4324 4527 4327
rect 5253 4324 5267 4327
rect 93 4313 107 4324
rect 333 4256 347 4270
rect 473 4262 487 4276
rect 33 4187 47 4201
rect 113 4207 127 4221
rect 253 4207 267 4221
rect 73 4187 87 4201
rect 133 4187 147 4201
rect 153 4179 167 4193
rect 173 4187 187 4201
rect 193 4187 207 4201
rect 213 4179 227 4193
rect 233 4187 247 4201
rect 373 4187 387 4201
rect 413 4187 427 4201
rect 473 4224 487 4238
rect 593 4253 607 4267
rect 533 4199 547 4213
rect 553 4207 567 4221
rect 493 4159 507 4173
rect 333 4130 347 4144
rect 573 4199 587 4213
rect 733 4213 747 4227
rect 633 4187 647 4201
rect 653 4179 667 4193
rect 673 4187 687 4201
rect 633 4153 647 4167
rect 693 4179 707 4193
rect 713 4187 727 4201
rect 833 4262 847 4276
rect 973 4256 987 4270
rect 753 4179 767 4193
rect 733 4153 747 4167
rect 473 4130 487 4144
rect 773 4167 787 4181
rect 833 4224 847 4238
rect 813 4159 827 4173
rect 893 4187 907 4201
rect 933 4187 947 4201
rect 833 4130 847 4144
rect 1153 4262 1167 4276
rect 1293 4256 1307 4270
rect 1033 4199 1047 4213
rect 1053 4207 1067 4221
rect 1073 4199 1087 4213
rect 1153 4224 1167 4238
rect 1133 4159 1147 4173
rect 1213 4187 1227 4201
rect 1253 4187 1267 4201
rect 973 4130 987 4144
rect 1153 4130 1167 4144
rect 1353 4199 1367 4213
rect 1373 4207 1387 4221
rect 1393 4199 1407 4213
rect 1513 4207 1527 4221
rect 1893 4262 1907 4276
rect 2033 4256 2047 4270
rect 1433 4167 1447 4181
rect 1453 4179 1467 4193
rect 1533 4187 1547 4201
rect 1293 4130 1307 4144
rect 1553 4179 1567 4193
rect 1573 4187 1587 4201
rect 1613 4187 1627 4201
rect 1713 4199 1727 4213
rect 1733 4207 1747 4221
rect 1633 4179 1647 4193
rect 1653 4167 1667 4181
rect 1673 4179 1687 4193
rect 1753 4199 1767 4213
rect 1773 4199 1787 4213
rect 1793 4207 1807 4221
rect 1813 4199 1827 4213
rect 1893 4224 1907 4238
rect 1873 4159 1887 4173
rect 1953 4187 1967 4201
rect 1993 4187 2007 4201
rect 1893 4130 1907 4144
rect 2313 4256 2327 4270
rect 2453 4262 2467 4276
rect 2093 4199 2107 4213
rect 2113 4207 2127 4221
rect 2133 4199 2147 4213
rect 2193 4207 2207 4221
rect 2213 4187 2227 4201
rect 2233 4179 2247 4193
rect 2253 4187 2267 4201
rect 2033 4130 2047 4144
rect 2353 4187 2367 4201
rect 2393 4187 2407 4201
rect 2453 4224 2467 4238
rect 2533 4187 2547 4201
rect 2473 4159 2487 4173
rect 2313 4130 2327 4144
rect 2453 4130 2467 4144
rect 2573 4187 2587 4201
rect 2733 4313 2747 4324
rect 2833 4313 2847 4324
rect 2713 4207 2727 4221
rect 2553 4167 2567 4181
rect 2593 4167 2607 4181
rect 2613 4179 2627 4193
rect 2653 4187 2667 4201
rect 2673 4179 2687 4193
rect 2693 4187 2707 4201
rect 2753 4199 2767 4213
rect 2773 4207 2787 4221
rect 2793 4199 2807 4213
rect 2853 4207 2867 4221
rect 2873 4187 2887 4201
rect 2893 4179 2907 4193
rect 2913 4187 2927 4201
rect 3053 4313 3067 4324
rect 2933 4167 2947 4181
rect 2953 4179 2967 4193
rect 2993 4187 3007 4201
rect 3033 4187 3047 4201
rect 3173 4262 3187 4276
rect 3313 4256 3327 4270
rect 3013 4167 3027 4181
rect 3093 4179 3107 4193
rect 3113 4167 3127 4181
rect 3173 4224 3187 4238
rect 3153 4159 3167 4173
rect 3233 4187 3247 4201
rect 3273 4187 3287 4201
rect 3173 4130 3187 4144
rect 4073 4313 4087 4324
rect 3373 4187 3387 4201
rect 3393 4179 3407 4193
rect 3413 4187 3427 4201
rect 3433 4179 3447 4193
rect 3453 4187 3467 4201
rect 3493 4199 3507 4213
rect 3513 4207 3527 4221
rect 3313 4130 3327 4144
rect 3533 4199 3547 4213
rect 3593 4179 3607 4193
rect 3773 4199 3787 4213
rect 3793 4207 3807 4221
rect 3733 4179 3747 4193
rect 3813 4199 3827 4213
rect 3853 4199 3867 4213
rect 3873 4207 3887 4221
rect 3893 4199 3907 4213
rect 3953 4199 3967 4213
rect 3973 4207 3987 4221
rect 3993 4199 4007 4213
rect 4313 4256 4327 4270
rect 4453 4262 4467 4276
rect 4093 4207 4107 4221
rect 4233 4207 4247 4221
rect 4013 4167 4027 4181
rect 4033 4179 4047 4193
rect 4113 4187 4127 4201
rect 4133 4179 4147 4193
rect 4153 4187 4167 4201
rect 4173 4187 4187 4201
rect 4193 4179 4207 4193
rect 4213 4187 4227 4201
rect 4353 4187 4367 4201
rect 4393 4187 4407 4201
rect 4453 4224 4467 4238
rect 4513 4313 4527 4324
rect 4653 4256 4667 4270
rect 4793 4262 4807 4276
rect 4533 4207 4547 4221
rect 4473 4159 4487 4173
rect 4553 4187 4567 4201
rect 4573 4179 4587 4193
rect 4593 4187 4607 4201
rect 4313 4130 4327 4144
rect 4453 4130 4467 4144
rect 4693 4187 4707 4201
rect 4733 4187 4747 4201
rect 4793 4224 4807 4238
rect 5033 4227 5047 4241
rect 5013 4207 5027 4221
rect 5053 4207 5067 4221
rect 5093 4233 5107 4247
rect 4873 4187 4887 4201
rect 4813 4159 4827 4173
rect 4653 4130 4667 4144
rect 4893 4179 4907 4193
rect 4933 4187 4947 4201
rect 5073 4199 5087 4213
rect 4953 4179 4967 4193
rect 4973 4167 4987 4181
rect 4993 4179 5007 4193
rect 4793 4130 4807 4144
rect 5073 4133 5087 4147
rect 5253 4313 5267 4324
rect 5313 4256 5327 4270
rect 5453 4262 5467 4276
rect 5233 4207 5247 4221
rect 5133 4179 5147 4193
rect 5173 4187 5187 4201
rect 5153 4167 5167 4181
rect 5193 4179 5207 4193
rect 5213 4187 5227 4201
rect 5353 4187 5367 4201
rect 5393 4187 5407 4201
rect 5453 4224 5467 4238
rect 5513 4199 5527 4213
rect 5533 4207 5547 4221
rect 5473 4159 5487 4173
rect 5313 4130 5327 4144
rect 5553 4199 5567 4213
rect 5713 4207 5727 4221
rect 5593 4167 5607 4181
rect 5613 4179 5627 4193
rect 5653 4187 5667 4201
rect 5673 4179 5687 4193
rect 5693 4187 5707 4201
rect 5453 4130 5467 4144
rect 5773 4187 5787 4201
rect 5793 4199 5807 4213
rect 5873 4227 5887 4241
rect 5853 4207 5867 4221
rect 5893 4207 5907 4221
rect 5833 4187 5847 4201
rect 5913 4199 5927 4213
rect 5953 4193 5967 4207
rect 6073 4207 6087 4221
rect 5973 4187 5987 4201
rect 5913 4133 5927 4147
rect 5993 4179 6007 4193
rect 6013 4187 6027 4201
rect 6033 4179 6047 4193
rect 6053 4187 6067 4201
rect 6113 4187 6127 4201
rect 6153 4187 6167 4201
rect 6193 4199 6207 4213
rect 6213 4207 6227 4221
rect 6233 4199 6247 4213
rect 6293 4187 6307 4201
rect 6313 4199 6327 4213
rect 6353 4187 6367 4201
rect 6373 4199 6387 4213
rect 6393 4207 6407 4221
rect 6413 4199 6427 4213
rect 6453 4213 6467 4227
rect 6633 4227 6647 4241
rect 6613 4207 6627 4221
rect 6653 4207 6667 4221
rect 6433 4173 6447 4187
rect 6453 4167 6467 4181
rect 6473 4179 6487 4193
rect 6533 4187 6547 4201
rect 6673 4199 6687 4213
rect 6553 4179 6567 4193
rect 6573 4167 6587 4181
rect 6593 4179 6607 4193
rect 133 4036 147 4050
rect 33 3979 47 3993
rect 273 4036 287 4050
rect 113 4007 127 4021
rect 73 3979 87 3993
rect 133 3942 147 3956
rect 193 3979 207 3993
rect 233 3979 247 3993
rect 333 3967 347 3981
rect 353 3959 367 3973
rect 373 3967 387 3981
rect 433 3979 447 3993
rect 453 3987 467 4001
rect 473 3999 487 4013
rect 493 3987 507 4001
rect 133 3904 147 3918
rect 273 3910 287 3924
rect 533 3967 547 3981
rect 553 3959 567 3973
rect 573 3967 587 3981
rect 613 3967 627 3981
rect 793 4036 807 4050
rect 633 3959 647 3973
rect 653 3967 667 3981
rect 693 3979 707 3993
rect 573 3933 587 3947
rect 613 3933 627 3947
rect 933 4036 947 4050
rect 773 4007 787 4021
rect 733 3979 747 3993
rect 793 3942 807 3956
rect 853 3979 867 3993
rect 893 3979 907 3993
rect 1013 3967 1027 3981
rect 1033 3959 1047 3973
rect 1053 3967 1067 3981
rect 1073 3967 1087 3981
rect 1133 4013 1147 4027
rect 1373 4036 1387 4050
rect 1093 3959 1107 3973
rect 1113 3967 1127 3981
rect 793 3904 807 3918
rect 933 3910 947 3924
rect 1153 3967 1167 3981
rect 1513 4036 1527 4050
rect 1173 3959 1187 3973
rect 1193 3967 1207 3981
rect 1253 3979 1267 3993
rect 1273 3987 1287 4001
rect 1293 3999 1307 4013
rect 1353 4007 1367 4021
rect 1313 3987 1327 4001
rect 1133 3913 1147 3927
rect 1373 3942 1387 3956
rect 1433 3979 1447 3993
rect 1473 3979 1487 3993
rect 1593 3967 1607 3981
rect 1613 3959 1627 3973
rect 1633 3967 1647 3981
rect 1653 3979 1667 3993
rect 1853 4036 1867 4050
rect 1693 3979 1707 3993
rect 1373 3904 1387 3918
rect 1513 3910 1527 3924
rect 1733 3967 1747 3981
rect 1993 4036 2007 4050
rect 1833 4007 1847 4021
rect 1753 3959 1767 3973
rect 1773 3967 1787 3981
rect 1853 3942 1867 3956
rect 1913 3979 1927 3993
rect 1953 3979 1967 3993
rect 2053 3967 2067 3981
rect 2073 3959 2087 3973
rect 2093 3967 2107 3981
rect 2173 3979 2187 3993
rect 2193 3987 2207 4001
rect 2213 3979 2227 3993
rect 2153 3959 2167 3973
rect 1853 3904 1867 3918
rect 1993 3910 2007 3924
rect 2253 3967 2267 3981
rect 2273 3959 2287 3973
rect 2293 3967 2307 3981
rect 2313 3967 2327 3981
rect 2413 3987 2427 4001
rect 2433 3999 2447 4013
rect 2333 3959 2347 3973
rect 2353 3967 2367 3981
rect 2493 3979 2507 3993
rect 2513 3987 2527 4001
rect 2573 3999 2587 4013
rect 2533 3979 2547 3993
rect 2553 3979 2567 3993
rect 2473 3959 2487 3973
rect 2673 3999 2687 4013
rect 2713 3999 2727 4013
rect 2593 3979 2607 3993
rect 2653 3979 2667 3993
rect 2693 3979 2707 3993
rect 2733 3987 2747 4001
rect 2793 3987 2807 4001
rect 2813 3999 2827 4013
rect 2853 3967 2867 3981
rect 2933 3999 2947 4013
rect 2873 3959 2887 3973
rect 2893 3967 2907 3981
rect 2913 3979 2927 3993
rect 2953 3979 2967 3993
rect 2993 3979 3007 3993
rect 3013 3987 3027 4001
rect 3093 3999 3107 4013
rect 3433 4036 3447 4050
rect 3033 3979 3047 3993
rect 3113 3987 3127 4001
rect 3173 3999 3187 4013
rect 3053 3959 3067 3973
rect 3153 3979 3167 3993
rect 3193 3979 3207 3993
rect 3253 3967 3267 3981
rect 3273 3959 3287 3973
rect 3293 3967 3307 3981
rect 3333 3967 3347 3981
rect 3353 3959 3367 3973
rect 3373 3967 3387 3981
rect 3573 4036 3587 4050
rect 3473 3979 3487 3993
rect 3513 3979 3527 3993
rect 3593 4007 3607 4021
rect 3573 3942 3587 3956
rect 3733 4036 3747 4050
rect 3653 3987 3667 4001
rect 3673 3999 3687 4013
rect 3433 3910 3447 3924
rect 3573 3904 3587 3918
rect 3873 4036 3887 4050
rect 3773 3979 3787 3993
rect 3813 3979 3827 3993
rect 3893 4007 3907 4021
rect 3873 3942 3887 3956
rect 3953 3967 3967 3981
rect 3733 3910 3747 3924
rect 3873 3904 3887 3918
rect 3973 3959 3987 3973
rect 4013 3959 4027 3973
rect 4033 3967 4047 3981
rect 4093 4013 4107 4027
rect 4053 3959 4067 3973
rect 4073 3967 4087 3981
rect 3993 3939 4007 3953
rect 4073 3933 4087 3947
rect 4153 3979 4167 3993
rect 4173 3987 4187 4001
rect 4233 3999 4247 4013
rect 4193 3979 4207 3993
rect 4213 3979 4227 3993
rect 4133 3959 4147 3973
rect 4253 3979 4267 3993
rect 4313 3987 4327 4001
rect 4333 3999 4347 4013
rect 4113 3856 4127 3867
rect 4373 3967 4387 3981
rect 4573 4036 4587 4050
rect 4393 3959 4407 3973
rect 4413 3967 4427 3981
rect 4473 3979 4487 3993
rect 4493 3987 4507 4001
rect 4513 3979 4527 3993
rect 4453 3959 4467 3973
rect 4713 4036 4727 4050
rect 4613 3979 4627 3993
rect 4653 3979 4667 3993
rect 4433 3856 4447 3867
rect 4733 4007 4747 4021
rect 4713 3942 4727 3956
rect 4793 3967 4807 3981
rect 4993 4036 5007 4050
rect 4813 3959 4827 3973
rect 4833 3967 4847 3981
rect 4893 3979 4907 3993
rect 4913 3987 4927 4001
rect 4933 3979 4947 3993
rect 4873 3959 4887 3973
rect 4573 3910 4587 3924
rect 4713 3904 4727 3918
rect 5133 4036 5147 4050
rect 5033 3979 5047 3993
rect 5073 3979 5087 3993
rect 4853 3856 4867 3867
rect 5153 4007 5167 4021
rect 5133 3942 5147 3956
rect 5213 3967 5227 3981
rect 5553 4033 5567 4047
rect 5233 3959 5247 3973
rect 5253 3967 5267 3981
rect 5313 3979 5327 3993
rect 5333 3987 5347 4001
rect 5353 3979 5367 3993
rect 5293 3959 5307 3973
rect 4993 3910 5007 3924
rect 5133 3904 5147 3918
rect 5393 3967 5407 3981
rect 5413 3959 5427 3973
rect 5433 3967 5447 3981
rect 5453 3979 5467 3993
rect 5473 3987 5487 4001
rect 5493 3979 5507 3993
rect 5273 3856 5287 3867
rect 5513 3959 5527 3973
rect 5653 4036 5667 4050
rect 5573 3987 5587 4001
rect 5593 3999 5607 4013
rect 5553 3953 5567 3967
rect 5793 4036 5807 4050
rect 5693 3979 5707 3993
rect 5733 3979 5747 3993
rect 5813 4007 5827 4021
rect 5793 3942 5807 3956
rect 5853 3999 5867 4013
rect 6053 4036 6067 4050
rect 6193 4036 6207 4050
rect 5873 3987 5887 4001
rect 5653 3910 5667 3924
rect 5793 3904 5807 3918
rect 6033 4007 6047 4021
rect 5933 3967 5947 3981
rect 5953 3959 5967 3973
rect 5993 3959 6007 3973
rect 5973 3939 5987 3953
rect 6053 3942 6067 3956
rect 6113 3979 6127 3993
rect 6153 3979 6167 3993
rect 6053 3904 6067 3918
rect 6193 3910 6207 3924
rect 6293 4036 6307 4050
rect 6433 4036 6447 4050
rect 6273 4007 6287 4021
rect 6293 3942 6307 3956
rect 6353 3979 6367 3993
rect 6393 3979 6407 3993
rect 6293 3904 6307 3918
rect 6433 3910 6447 3924
rect 6533 4036 6547 4050
rect 6673 4036 6687 4050
rect 6513 4007 6527 4021
rect 6533 3942 6547 3956
rect 6593 3979 6607 3993
rect 6633 3979 6647 3993
rect 6533 3904 6547 3918
rect 6673 3910 6687 3924
rect 4113 3853 4127 3856
rect 4433 3853 4447 3856
rect 4853 3853 4867 3856
rect 5273 3853 5287 3856
rect 2053 3844 2067 3847
rect 2233 3844 2247 3847
rect 33 3707 47 3721
rect 293 3782 307 3796
rect 433 3776 447 3790
rect 73 3707 87 3721
rect 113 3707 127 3721
rect 153 3707 167 3721
rect 193 3719 207 3733
rect 213 3727 227 3741
rect 233 3719 247 3733
rect 293 3744 307 3758
rect 273 3679 287 3693
rect 353 3707 367 3721
rect 393 3707 407 3721
rect 293 3650 307 3664
rect 573 3733 587 3747
rect 613 3753 627 3767
rect 873 3782 887 3796
rect 1013 3776 1027 3790
rect 513 3707 527 3721
rect 613 3719 627 3733
rect 633 3727 647 3741
rect 433 3650 447 3664
rect 533 3699 547 3713
rect 553 3687 567 3701
rect 573 3699 587 3713
rect 653 3719 667 3733
rect 673 3719 687 3733
rect 693 3727 707 3741
rect 713 3719 727 3733
rect 773 3719 787 3733
rect 793 3727 807 3741
rect 813 3719 827 3733
rect 873 3744 887 3758
rect 853 3679 867 3693
rect 933 3707 947 3721
rect 973 3707 987 3721
rect 873 3650 887 3664
rect 1073 3699 1087 3713
rect 1093 3687 1107 3701
rect 1113 3699 1127 3713
rect 1133 3707 1147 3721
rect 1193 3719 1207 3733
rect 1213 3727 1227 3741
rect 1233 3719 1247 3733
rect 1253 3707 1267 3721
rect 1013 3650 1027 3664
rect 1713 3782 1727 3796
rect 1853 3776 1867 3790
rect 1293 3707 1307 3721
rect 1353 3707 1367 3721
rect 1453 3719 1467 3733
rect 1473 3727 1487 3741
rect 1333 3693 1347 3707
rect 1333 3653 1347 3667
rect 1373 3699 1387 3713
rect 1393 3687 1407 3701
rect 1413 3699 1427 3713
rect 1493 3719 1507 3733
rect 1513 3719 1527 3733
rect 1533 3727 1547 3741
rect 1553 3719 1567 3733
rect 1593 3707 1607 3721
rect 1633 3707 1647 3721
rect 1613 3687 1627 3701
rect 1713 3744 1727 3758
rect 1693 3679 1707 3693
rect 1773 3707 1787 3721
rect 1813 3707 1827 3721
rect 1713 3650 1727 3664
rect 2053 3833 2067 3844
rect 1933 3719 1947 3733
rect 1953 3727 1967 3741
rect 1973 3719 1987 3733
rect 1993 3707 2007 3721
rect 2033 3707 2047 3721
rect 2233 3833 2247 3844
rect 2193 3727 2207 3741
rect 2253 3727 2267 3741
rect 2013 3687 2027 3701
rect 2073 3687 2087 3701
rect 2093 3699 2107 3713
rect 2133 3707 2147 3721
rect 2153 3699 2167 3713
rect 2173 3707 2187 3721
rect 1853 3650 1867 3664
rect 2273 3707 2287 3721
rect 2293 3699 2307 3713
rect 2313 3707 2327 3721
rect 2353 3707 2367 3721
rect 2673 3747 2687 3761
rect 2613 3727 2627 3741
rect 2653 3727 2667 3741
rect 2693 3727 2707 3741
rect 2373 3699 2387 3713
rect 2393 3687 2407 3701
rect 2413 3699 2427 3713
rect 2433 3687 2447 3701
rect 2453 3699 2467 3713
rect 2513 3699 2527 3713
rect 2553 3707 2567 3721
rect 2473 3673 2487 3687
rect 2493 3653 2507 3667
rect 2533 3687 2547 3701
rect 2573 3699 2587 3713
rect 2593 3707 2607 3721
rect 2713 3719 2727 3733
rect 2793 3733 2807 3747
rect 2773 3699 2787 3713
rect 2833 3719 2847 3733
rect 2853 3727 2867 3741
rect 2793 3687 2807 3701
rect 2813 3693 2827 3707
rect 2873 3719 2887 3733
rect 2953 3727 2967 3741
rect 3053 3727 3067 3741
rect 3513 3776 3527 3790
rect 3653 3782 3667 3796
rect 2893 3707 2907 3721
rect 2913 3699 2927 3713
rect 2933 3707 2947 3721
rect 2993 3707 3007 3721
rect 3013 3699 3027 3713
rect 3033 3707 3047 3721
rect 3093 3699 3107 3713
rect 3113 3687 3127 3701
rect 3133 3699 3147 3713
rect 3153 3707 3167 3721
rect 3213 3707 3227 3721
rect 3233 3699 3247 3713
rect 3253 3707 3267 3721
rect 3273 3699 3287 3713
rect 3293 3707 3307 3721
rect 3333 3719 3347 3733
rect 3353 3727 3367 3741
rect 3373 3719 3387 3733
rect 3413 3719 3427 3733
rect 3433 3727 3447 3741
rect 3453 3719 3467 3733
rect 3553 3707 3567 3721
rect 3593 3707 3607 3721
rect 3653 3744 3667 3758
rect 3733 3719 3747 3733
rect 3753 3727 3767 3741
rect 3673 3679 3687 3693
rect 3513 3650 3527 3664
rect 3773 3719 3787 3733
rect 3813 3707 3827 3721
rect 3833 3699 3847 3713
rect 3853 3707 3867 3721
rect 3653 3650 3667 3664
rect 3873 3699 3887 3713
rect 3893 3707 3907 3721
rect 4193 3776 4207 3790
rect 4333 3782 4347 3796
rect 3973 3719 3987 3733
rect 3993 3727 4007 3741
rect 3913 3687 3927 3701
rect 3933 3699 3947 3713
rect 4013 3719 4027 3733
rect 4113 3727 4127 3741
rect 4053 3707 4067 3721
rect 4073 3699 4087 3713
rect 4093 3707 4107 3721
rect 4233 3707 4247 3721
rect 4273 3707 4287 3721
rect 4333 3744 4347 3758
rect 4793 3776 4807 3790
rect 4933 3782 4947 3796
rect 4393 3719 4407 3733
rect 4413 3727 4427 3741
rect 4353 3679 4367 3693
rect 4193 3650 4207 3664
rect 4433 3719 4447 3733
rect 4493 3719 4507 3733
rect 4513 3727 4527 3741
rect 4533 3719 4547 3733
rect 4573 3699 4587 3713
rect 4333 3650 4347 3664
rect 4713 3699 4727 3713
rect 4833 3707 4847 3721
rect 4873 3707 4887 3721
rect 4933 3744 4947 3758
rect 5053 3727 5067 3741
rect 4993 3707 5007 3721
rect 5013 3699 5027 3713
rect 5033 3707 5047 3721
rect 5113 3719 5127 3733
rect 5133 3727 5147 3741
rect 4953 3679 4967 3693
rect 4793 3650 4807 3664
rect 5153 3719 5167 3733
rect 4933 3650 4947 3664
rect 5153 3673 5167 3687
rect 5193 3753 5207 3767
rect 5253 3753 5267 3767
rect 5193 3719 5207 3733
rect 5213 3727 5227 3741
rect 5233 3719 5247 3733
rect 5233 3673 5247 3687
rect 5553 3782 5567 3796
rect 5693 3776 5707 3790
rect 5273 3699 5287 3713
rect 5293 3687 5307 3701
rect 5333 3699 5347 3713
rect 5473 3699 5487 3713
rect 5553 3744 5567 3758
rect 5533 3679 5547 3693
rect 5613 3707 5627 3721
rect 5653 3707 5667 3721
rect 5553 3650 5567 3664
rect 5813 3719 5827 3733
rect 5833 3727 5847 3741
rect 5773 3699 5787 3713
rect 5693 3650 5707 3664
rect 5793 3687 5807 3701
rect 5853 3719 5867 3733
rect 5893 3719 5907 3733
rect 5913 3727 5927 3741
rect 5933 3719 5947 3733
rect 6333 3782 6347 3796
rect 6473 3776 6487 3790
rect 5993 3699 6007 3713
rect 6033 3707 6047 3721
rect 6073 3707 6087 3721
rect 6133 3707 6147 3721
rect 6013 3687 6027 3701
rect 6053 3687 6067 3701
rect 6173 3707 6187 3721
rect 6153 3687 6167 3701
rect 6193 3699 6207 3713
rect 6213 3687 6227 3701
rect 6233 3699 6247 3713
rect 6253 3707 6267 3721
rect 6333 3744 6347 3758
rect 6313 3679 6327 3693
rect 6393 3707 6407 3721
rect 6433 3707 6447 3721
rect 6333 3650 6347 3664
rect 6593 3727 6607 3741
rect 6533 3707 6547 3721
rect 6553 3699 6567 3713
rect 6573 3707 6587 3721
rect 6633 3719 6647 3733
rect 6653 3727 6667 3741
rect 6473 3650 6487 3664
rect 6673 3719 6687 3733
rect 133 3556 147 3570
rect 33 3499 47 3513
rect 273 3556 287 3570
rect 113 3527 127 3541
rect 73 3499 87 3513
rect 133 3462 147 3476
rect 193 3499 207 3513
rect 233 3499 247 3513
rect 333 3487 347 3501
rect 353 3479 367 3493
rect 373 3487 387 3501
rect 413 3499 427 3513
rect 453 3499 467 3513
rect 513 3499 527 3513
rect 533 3507 547 3521
rect 553 3519 567 3533
rect 573 3507 587 3521
rect 133 3424 147 3438
rect 273 3430 287 3444
rect 613 3487 627 3501
rect 633 3479 647 3493
rect 653 3487 667 3501
rect 693 3499 707 3513
rect 733 3499 747 3513
rect 753 3499 767 3513
rect 793 3499 807 3513
rect 833 3487 847 3501
rect 853 3479 867 3493
rect 873 3487 887 3501
rect 933 3499 947 3513
rect 973 3499 987 3513
rect 1013 3507 1027 3521
rect 1033 3519 1047 3533
rect 1073 3499 1087 3513
rect 1253 3556 1267 3570
rect 1113 3499 1127 3513
rect 1153 3499 1167 3513
rect 1393 3556 1407 3570
rect 1233 3527 1247 3541
rect 1193 3499 1207 3513
rect 1253 3462 1267 3476
rect 1313 3499 1327 3513
rect 1353 3499 1367 3513
rect 1573 3556 1587 3570
rect 1713 3556 1727 3570
rect 1493 3519 1507 3533
rect 1553 3527 1567 3541
rect 1473 3499 1487 3513
rect 1513 3499 1527 3513
rect 1253 3424 1267 3438
rect 1393 3430 1407 3444
rect 1453 3376 1467 3387
rect 1573 3462 1587 3476
rect 1633 3499 1647 3513
rect 1673 3499 1687 3513
rect 1793 3499 1807 3513
rect 1813 3487 1827 3501
rect 1573 3424 1587 3438
rect 1713 3430 1727 3444
rect 1853 3499 1867 3513
rect 1893 3507 1907 3521
rect 1913 3519 1927 3533
rect 1973 3499 1987 3513
rect 1993 3507 2007 3521
rect 2053 3519 2067 3533
rect 2013 3499 2027 3513
rect 2033 3499 2047 3513
rect 1953 3479 1967 3493
rect 2073 3499 2087 3513
rect 2133 3507 2147 3521
rect 2153 3519 2167 3533
rect 2193 3499 2207 3513
rect 2213 3487 2227 3501
rect 2393 3556 2407 3570
rect 2533 3556 2547 3570
rect 2313 3519 2327 3533
rect 2373 3527 2387 3541
rect 2253 3499 2267 3513
rect 2293 3499 2307 3513
rect 2333 3499 2347 3513
rect 2393 3462 2407 3476
rect 2453 3499 2467 3513
rect 2493 3499 2507 3513
rect 2613 3519 2627 3533
rect 2593 3499 2607 3513
rect 2633 3499 2647 3513
rect 2673 3499 2687 3513
rect 2693 3507 2707 3521
rect 2713 3499 2727 3513
rect 2793 3507 2807 3521
rect 2813 3519 2827 3533
rect 2733 3479 2747 3493
rect 2393 3424 2407 3438
rect 2533 3430 2547 3444
rect 2853 3487 2867 3501
rect 2873 3479 2887 3493
rect 2893 3487 2907 3501
rect 2913 3499 2927 3513
rect 2933 3507 2947 3521
rect 2953 3499 2967 3513
rect 3013 3507 3027 3521
rect 3033 3519 3047 3533
rect 3053 3507 3067 3521
rect 3073 3499 3087 3513
rect 3113 3507 3127 3521
rect 3133 3499 3147 3513
rect 3193 3499 3207 3513
rect 3213 3507 3227 3521
rect 3233 3499 3247 3513
rect 3393 3556 3407 3570
rect 3533 3556 3547 3570
rect 3753 3556 3767 3570
rect 3253 3507 3267 3521
rect 3273 3499 3287 3513
rect 3313 3507 3327 3521
rect 3333 3519 3347 3533
rect 3373 3527 3387 3541
rect 2973 3479 2987 3493
rect 3393 3462 3407 3476
rect 3453 3499 3467 3513
rect 3493 3499 3507 3513
rect 3613 3499 3627 3513
rect 3633 3507 3647 3521
rect 3893 3556 3907 3570
rect 3653 3499 3667 3513
rect 3733 3527 3747 3541
rect 3673 3507 3687 3521
rect 3693 3499 3707 3513
rect 3393 3424 3407 3438
rect 3533 3430 3547 3444
rect 3753 3462 3767 3476
rect 3813 3499 3827 3513
rect 3853 3499 3867 3513
rect 4053 3556 4067 3570
rect 4193 3556 4207 3570
rect 3973 3507 3987 3521
rect 3993 3519 4007 3533
rect 4033 3527 4047 3541
rect 3753 3424 3767 3438
rect 3893 3430 3907 3444
rect 4053 3462 4067 3476
rect 4113 3499 4127 3513
rect 4153 3499 4167 3513
rect 4273 3507 4287 3521
rect 4293 3519 4307 3533
rect 4493 3556 4507 3570
rect 4333 3507 4347 3521
rect 4353 3519 4367 3533
rect 4053 3424 4067 3438
rect 4193 3430 4207 3444
rect 4373 3487 4387 3501
rect 4393 3479 4407 3493
rect 4413 3487 4427 3501
rect 4633 3556 4647 3570
rect 4533 3499 4547 3513
rect 4573 3499 4587 3513
rect 4653 3527 4667 3541
rect 4633 3462 4647 3476
rect 4793 3556 4807 3570
rect 4933 3556 4947 3570
rect 4713 3507 4727 3521
rect 4733 3519 4747 3533
rect 4773 3527 4787 3541
rect 4493 3430 4507 3444
rect 4633 3424 4647 3438
rect 4793 3462 4807 3476
rect 4853 3499 4867 3513
rect 4893 3499 4907 3513
rect 5013 3499 5027 3513
rect 5033 3507 5047 3521
rect 5053 3499 5067 3513
rect 5213 3556 5227 3570
rect 5353 3556 5367 3570
rect 5073 3507 5087 3521
rect 5093 3499 5107 3513
rect 5133 3507 5147 3521
rect 5153 3519 5167 3533
rect 5193 3527 5207 3541
rect 4793 3424 4807 3438
rect 4933 3430 4947 3444
rect 5213 3462 5227 3476
rect 5273 3499 5287 3513
rect 5313 3499 5327 3513
rect 5213 3424 5227 3438
rect 5353 3430 5367 3444
rect 5453 3556 5467 3570
rect 5593 3556 5607 3570
rect 5433 3527 5447 3541
rect 5453 3462 5467 3476
rect 5513 3499 5527 3513
rect 5553 3499 5567 3513
rect 5653 3499 5667 3513
rect 5673 3507 5687 3521
rect 5693 3499 5707 3513
rect 5753 3499 5767 3513
rect 5773 3507 5787 3521
rect 5893 3553 5907 3567
rect 5793 3499 5807 3513
rect 5873 3507 5887 3521
rect 5893 3519 5907 3533
rect 5713 3479 5727 3493
rect 5813 3479 5827 3493
rect 5453 3424 5467 3438
rect 5593 3430 5607 3444
rect 5893 3473 5907 3487
rect 5933 3499 5947 3513
rect 5953 3507 5967 3521
rect 5973 3499 5987 3513
rect 5993 3507 6007 3521
rect 6013 3499 6027 3513
rect 6033 3487 6047 3501
rect 6133 3507 6147 3521
rect 6153 3519 6167 3533
rect 6453 3556 6467 3570
rect 6593 3556 6607 3570
rect 6053 3479 6067 3493
rect 6073 3487 6087 3501
rect 6193 3499 6207 3513
rect 6233 3507 6247 3521
rect 6253 3499 6267 3513
rect 6293 3507 6307 3521
rect 6373 3507 6387 3521
rect 6393 3519 6407 3533
rect 6433 3527 6447 3541
rect 6453 3462 6467 3476
rect 6513 3499 6527 3513
rect 6553 3499 6567 3513
rect 6453 3424 6467 3438
rect 6593 3430 6607 3444
rect 1453 3373 1467 3376
rect 1153 3364 1167 3367
rect 2373 3364 2387 3367
rect 3433 3364 3447 3367
rect 4473 3364 4487 3367
rect 133 3302 147 3316
rect 273 3296 287 3310
rect 33 3227 47 3241
rect 73 3227 87 3241
rect 133 3264 147 3278
rect 113 3199 127 3213
rect 193 3227 207 3241
rect 233 3227 247 3241
rect 133 3170 147 3184
rect 333 3239 347 3253
rect 353 3247 367 3261
rect 373 3239 387 3253
rect 493 3253 507 3267
rect 533 3273 547 3287
rect 433 3227 447 3241
rect 533 3239 547 3253
rect 553 3247 567 3261
rect 273 3170 287 3184
rect 453 3219 467 3233
rect 473 3207 487 3221
rect 493 3219 507 3233
rect 573 3239 587 3253
rect 633 3273 647 3287
rect 593 3207 607 3221
rect 613 3219 627 3233
rect 673 3267 687 3281
rect 653 3247 667 3261
rect 693 3247 707 3261
rect 713 3239 727 3253
rect 753 3239 767 3253
rect 773 3247 787 3261
rect 633 3193 647 3207
rect 793 3239 807 3253
rect 853 3247 867 3261
rect 873 3227 887 3241
rect 893 3219 907 3233
rect 913 3227 927 3241
rect 1153 3353 1167 3364
rect 933 3207 947 3221
rect 953 3219 967 3233
rect 993 3227 1007 3241
rect 1133 3247 1147 3261
rect 1393 3302 1407 3316
rect 1533 3296 1547 3310
rect 1233 3247 1247 3261
rect 1033 3227 1047 3241
rect 1073 3227 1087 3241
rect 1013 3207 1027 3221
rect 1093 3219 1107 3233
rect 1113 3227 1127 3241
rect 1173 3227 1187 3241
rect 1193 3219 1207 3233
rect 1213 3227 1227 3241
rect 1273 3239 1287 3253
rect 1293 3247 1307 3261
rect 1313 3239 1327 3253
rect 1393 3264 1407 3278
rect 1373 3199 1387 3213
rect 1453 3227 1467 3241
rect 1493 3227 1507 3241
rect 1393 3170 1407 3184
rect 1533 3170 1547 3184
rect 1613 3227 1627 3241
rect 1633 3239 1647 3253
rect 1853 3267 1867 3281
rect 2033 3296 2047 3310
rect 2173 3302 2187 3316
rect 1673 3227 1687 3241
rect 1713 3227 1727 3241
rect 1813 3239 1827 3253
rect 1833 3247 1847 3261
rect 1873 3247 1887 3261
rect 1733 3219 1747 3233
rect 1753 3207 1767 3221
rect 1773 3219 1787 3233
rect 1893 3219 1907 3233
rect 1913 3207 1927 3221
rect 1933 3219 1947 3233
rect 1953 3227 1967 3241
rect 2073 3227 2087 3241
rect 2113 3227 2127 3241
rect 2173 3264 2187 3278
rect 2373 3353 2387 3364
rect 2233 3239 2247 3253
rect 2253 3247 2267 3261
rect 2193 3199 2207 3213
rect 2033 3170 2047 3184
rect 2273 3239 2287 3253
rect 2313 3227 2327 3241
rect 2353 3227 2367 3241
rect 2413 3227 2427 3241
rect 2333 3207 2347 3221
rect 2173 3170 2187 3184
rect 2493 3247 2507 3261
rect 2453 3227 2467 3241
rect 2513 3227 2527 3241
rect 2433 3207 2447 3221
rect 2533 3219 2547 3233
rect 2553 3227 2567 3241
rect 2673 3296 2687 3310
rect 2813 3302 2827 3316
rect 2573 3207 2587 3221
rect 2593 3219 2607 3233
rect 2713 3227 2727 3241
rect 2753 3227 2767 3241
rect 2813 3264 2827 3278
rect 2873 3239 2887 3253
rect 2893 3247 2907 3261
rect 2833 3199 2847 3213
rect 2673 3170 2687 3184
rect 2913 3239 2927 3253
rect 2973 3239 2987 3253
rect 2993 3247 3007 3261
rect 3013 3239 3027 3253
rect 3053 3293 3067 3307
rect 3053 3247 3067 3261
rect 3033 3233 3047 3247
rect 3073 3227 3087 3241
rect 3093 3219 3107 3233
rect 3113 3227 3127 3241
rect 3153 3239 3167 3253
rect 3173 3247 3187 3261
rect 2813 3170 2827 3184
rect 3193 3239 3207 3253
rect 3433 3353 3447 3364
rect 3253 3253 3267 3267
rect 3233 3219 3247 3233
rect 3293 3247 3307 3261
rect 3313 3227 3327 3241
rect 3253 3207 3267 3221
rect 3293 3213 3307 3227
rect 3333 3219 3347 3233
rect 3353 3227 3367 3241
rect 3733 3302 3747 3316
rect 3873 3296 3887 3310
rect 3373 3207 3387 3221
rect 3393 3219 3407 3233
rect 3453 3227 3467 3241
rect 3573 3253 3587 3267
rect 3493 3227 3507 3241
rect 3533 3227 3547 3241
rect 3473 3207 3487 3221
rect 3553 3219 3567 3233
rect 3573 3207 3587 3221
rect 3593 3219 3607 3233
rect 3633 3227 3647 3241
rect 3673 3227 3687 3241
rect 3653 3207 3667 3221
rect 3733 3264 3747 3278
rect 3633 3193 3647 3207
rect 3713 3199 3727 3213
rect 4213 3296 4227 3310
rect 4353 3302 4367 3316
rect 3793 3227 3807 3241
rect 3833 3227 3847 3241
rect 3733 3170 3747 3184
rect 3933 3227 3947 3241
rect 3953 3219 3967 3233
rect 3973 3227 3987 3241
rect 3993 3219 4007 3233
rect 4013 3227 4027 3241
rect 4073 3227 4087 3241
rect 4093 3219 4107 3233
rect 4113 3227 4127 3241
rect 4133 3219 4147 3233
rect 4153 3227 4167 3241
rect 4253 3227 4267 3241
rect 4293 3227 4307 3241
rect 4353 3264 4367 3278
rect 4473 3353 4487 3364
rect 4413 3227 4427 3241
rect 4473 3253 4487 3267
rect 4453 3227 4467 3241
rect 4373 3199 4387 3213
rect 4433 3207 4447 3221
rect 4493 3227 4507 3241
rect 4513 3219 4527 3233
rect 4533 3227 4547 3241
rect 3873 3170 3887 3184
rect 4213 3170 4227 3184
rect 4353 3170 4367 3184
rect 4473 3193 4487 3207
rect 4553 3219 4567 3233
rect 4573 3227 4587 3241
rect 4613 3227 4627 3241
rect 4653 3227 4667 3241
rect 4693 3227 4707 3241
rect 4733 3227 4747 3241
rect 5093 3302 5107 3316
rect 5233 3296 5247 3310
rect 4633 3207 4647 3221
rect 4713 3207 4727 3221
rect 4773 3207 4787 3221
rect 4793 3219 4807 3233
rect 4833 3227 4847 3241
rect 4853 3219 4867 3233
rect 4653 3193 4667 3207
rect 4693 3193 4707 3207
rect 4873 3227 4887 3241
rect 4893 3219 4907 3233
rect 4913 3227 4927 3241
rect 4953 3219 4967 3233
rect 4973 3207 4987 3221
rect 4993 3219 5007 3233
rect 5013 3227 5027 3241
rect 5093 3264 5107 3278
rect 5073 3199 5087 3213
rect 5153 3227 5167 3241
rect 5193 3227 5207 3241
rect 5093 3170 5107 3184
rect 5313 3219 5327 3233
rect 5233 3170 5247 3184
rect 5333 3207 5347 3221
rect 5353 3219 5367 3233
rect 5373 3227 5387 3241
rect 5413 3219 5427 3233
rect 5433 3227 5447 3241
rect 5573 3296 5587 3310
rect 5713 3302 5727 3316
rect 5493 3219 5507 3233
rect 5513 3207 5527 3221
rect 5613 3227 5627 3241
rect 5653 3227 5667 3241
rect 5713 3264 5727 3278
rect 5793 3247 5807 3261
rect 5733 3199 5747 3213
rect 5813 3227 5827 3241
rect 5833 3219 5847 3233
rect 5853 3227 5867 3241
rect 6093 3247 6107 3261
rect 5893 3219 5907 3233
rect 5953 3227 5967 3241
rect 5573 3170 5587 3184
rect 5713 3170 5727 3184
rect 5913 3207 5927 3221
rect 5973 3219 5987 3233
rect 5993 3207 6007 3221
rect 6013 3219 6027 3233
rect 6033 3227 6047 3241
rect 6053 3219 6067 3233
rect 6073 3227 6087 3241
rect 6133 3273 6147 3287
rect 6153 3239 6167 3253
rect 6173 3247 6187 3261
rect 6113 3193 6127 3207
rect 6193 3239 6207 3253
rect 6533 3302 6547 3316
rect 6673 3296 6687 3310
rect 6233 3227 6247 3241
rect 6333 3239 6347 3253
rect 6353 3247 6367 3261
rect 6253 3219 6267 3233
rect 6273 3207 6287 3221
rect 6293 3219 6307 3233
rect 6373 3239 6387 3253
rect 6453 3247 6467 3261
rect 6393 3227 6407 3241
rect 6413 3219 6427 3233
rect 6433 3227 6447 3241
rect 6533 3264 6547 3278
rect 6513 3199 6527 3213
rect 6593 3227 6607 3241
rect 6633 3227 6647 3241
rect 6533 3170 6547 3184
rect 6673 3170 6687 3184
rect 33 3027 47 3041
rect 173 3027 187 3041
rect 333 3076 347 3090
rect 233 3019 247 3033
rect 273 3019 287 3033
rect 473 3076 487 3090
rect 673 3073 687 3087
rect 373 3019 387 3033
rect 413 3019 427 3033
rect 493 3047 507 3061
rect 473 2982 487 2996
rect 553 3007 567 3021
rect 573 2999 587 3013
rect 593 3007 607 3021
rect 613 3007 627 3021
rect 673 3033 687 3047
rect 633 2999 647 3013
rect 653 3007 667 3021
rect 333 2950 347 2964
rect 473 2944 487 2958
rect 653 2973 667 2987
rect 793 3053 807 3067
rect 733 3019 747 3033
rect 753 3027 767 3041
rect 773 3019 787 3033
rect 693 2993 707 3007
rect 713 2999 727 3013
rect 813 3007 827 3021
rect 853 3053 867 3067
rect 833 2999 847 3013
rect 853 3007 867 3021
rect 793 2973 807 2987
rect 893 3007 907 3021
rect 953 3027 967 3041
rect 973 3039 987 3053
rect 993 3027 1007 3041
rect 1093 3076 1107 3090
rect 1233 3076 1247 3090
rect 1073 3047 1087 3061
rect 913 2999 927 3013
rect 933 3007 947 3021
rect 1013 3019 1027 3033
rect 873 2953 887 2967
rect 1093 2982 1107 2996
rect 1153 3019 1167 3033
rect 1193 3019 1207 3033
rect 1413 3076 1427 3090
rect 1313 3007 1327 3021
rect 1553 3076 1567 3090
rect 1393 3047 1407 3061
rect 1333 2999 1347 3013
rect 1353 3007 1367 3021
rect 1093 2944 1107 2958
rect 1233 2950 1247 2964
rect 1413 2982 1427 2996
rect 1473 3019 1487 3033
rect 1513 3019 1527 3033
rect 1633 3027 1647 3041
rect 1653 3039 1667 3053
rect 1413 2944 1427 2958
rect 1553 2950 1567 2964
rect 1713 3019 1727 3033
rect 1733 3027 1747 3041
rect 1813 3039 1827 3053
rect 1753 3019 1767 3033
rect 1793 3019 1807 3033
rect 1693 2999 1707 3013
rect 1833 3019 1847 3033
rect 1873 3019 1887 3033
rect 1893 3007 1907 3021
rect 1933 3019 1947 3033
rect 1953 3019 1967 3033
rect 1973 3027 1987 3041
rect 1993 3019 2007 3033
rect 2073 3019 2087 3033
rect 2093 3027 2107 3041
rect 2113 3039 2127 3053
rect 2133 3027 2147 3041
rect 2013 2999 2027 3013
rect 2153 3007 2167 3021
rect 2253 3027 2267 3041
rect 2273 3039 2287 3053
rect 2173 2999 2187 3013
rect 2193 3007 2207 3021
rect 2193 2973 2207 2987
rect 2233 2973 2247 2987
rect 2293 3019 2307 3033
rect 2333 3007 2347 3021
rect 2353 3019 2367 3033
rect 2433 3076 2447 3090
rect 2573 3076 2587 3090
rect 2473 3019 2487 3033
rect 2513 3019 2527 3033
rect 2593 3047 2607 3061
rect 2573 2982 2587 2996
rect 2633 3039 2647 3053
rect 2653 3027 2667 3041
rect 2713 3039 2727 3053
rect 2433 2950 2447 2964
rect 2573 2944 2587 2958
rect 2693 3019 2707 3033
rect 2733 3019 2747 3033
rect 2793 3027 2807 3041
rect 2813 3039 2827 3053
rect 2873 3019 2887 3033
rect 2893 3027 2907 3041
rect 2913 3019 2927 3033
rect 2933 3027 2947 3041
rect 2953 3019 2967 3033
rect 2853 2999 2867 3013
rect 3013 3007 3027 3021
rect 3033 2999 3047 3013
rect 3073 2999 3087 3013
rect 3113 3007 3127 3021
rect 3413 3073 3427 3087
rect 3873 3076 3887 3090
rect 3133 2999 3147 3013
rect 3153 3007 3167 3021
rect 3053 2979 3067 2993
rect 3193 3033 3207 3047
rect 3213 3019 3227 3033
rect 3233 3027 3247 3041
rect 3253 3019 3267 3033
rect 3193 2999 3207 3013
rect 3273 3007 3287 3021
rect 3333 3053 3347 3067
rect 3293 2999 3307 3013
rect 3313 3007 3327 3021
rect 3193 2953 3207 2967
rect 3353 3007 3367 3021
rect 3373 2999 3387 3013
rect 3393 3007 3407 3021
rect 3433 3019 3447 3033
rect 3453 3027 3467 3041
rect 3513 3053 3527 3067
rect 3473 3019 3487 3033
rect 3353 2973 3367 2987
rect 3313 2953 3327 2967
rect 3353 2953 3367 2967
rect 3413 2993 3427 3007
rect 3493 2999 3507 3013
rect 3533 3019 3547 3033
rect 3533 2973 3547 2987
rect 3573 3007 3587 3021
rect 3593 3019 3607 3033
rect 3653 3019 3667 3033
rect 3673 3027 3687 3041
rect 3733 3053 3747 3067
rect 3693 3019 3707 3033
rect 3713 3027 3727 3041
rect 3733 3019 3747 3033
rect 3773 3027 3787 3041
rect 3813 3027 3827 3041
rect 3753 2993 3767 3007
rect 4013 3076 4027 3090
rect 3913 3019 3927 3033
rect 3953 3019 3967 3033
rect 4033 3047 4047 3061
rect 4013 2982 4027 2996
rect 4073 3019 4087 3033
rect 4093 3027 4107 3041
rect 4113 3019 4127 3033
rect 4313 3076 4327 3090
rect 4133 2999 4147 3013
rect 4193 3007 4207 3021
rect 3873 2950 3887 2964
rect 4013 2944 4027 2958
rect 4213 2999 4227 3013
rect 4253 2999 4267 3013
rect 4233 2979 4247 2993
rect 4453 3076 4467 3090
rect 4353 3019 4367 3033
rect 4393 3019 4407 3033
rect 4473 3047 4487 3061
rect 4453 2982 4467 2996
rect 4533 3019 4547 3033
rect 4553 3027 4567 3041
rect 4573 3019 4587 3033
rect 4593 3027 4607 3041
rect 4613 3019 4627 3033
rect 4653 3027 4667 3041
rect 4673 3039 4687 3053
rect 4313 2950 4327 2964
rect 4453 2944 4467 2958
rect 4713 3019 4727 3033
rect 4733 3027 4747 3041
rect 4773 3019 4787 3033
rect 4793 3027 4807 3041
rect 4813 3019 4827 3033
rect 4833 3027 4847 3041
rect 4853 3019 4867 3033
rect 4873 3027 4887 3041
rect 4893 3019 4907 3033
rect 4953 3027 4967 3041
rect 4973 3039 4987 3053
rect 4993 3019 5007 3033
rect 5013 3027 5027 3041
rect 5033 3019 5047 3033
rect 5053 3027 5067 3041
rect 5113 3039 5127 3053
rect 5073 3019 5087 3033
rect 5133 3027 5147 3041
rect 5193 3039 5207 3053
rect 5173 3019 5187 3033
rect 5293 3076 5307 3090
rect 5213 3019 5227 3033
rect 5433 3076 5447 3090
rect 5333 3019 5347 3033
rect 5373 3019 5387 3033
rect 5453 3047 5467 3061
rect 5433 2982 5447 2996
rect 5533 3039 5547 3053
rect 5513 3019 5527 3033
rect 5553 3019 5567 3033
rect 5573 3019 5587 3033
rect 5593 3027 5607 3041
rect 5613 3019 5627 3033
rect 5293 2950 5307 2964
rect 5433 2944 5447 2958
rect 5653 3013 5667 3027
rect 5633 2999 5647 3013
rect 5633 2953 5647 2967
rect 5693 3007 5707 3021
rect 5793 3019 5807 3033
rect 5813 3027 5827 3041
rect 5833 3019 5847 3033
rect 5853 3027 5867 3041
rect 5893 3039 5907 3053
rect 5873 3019 5887 3033
rect 5913 3027 5927 3041
rect 5953 3027 5967 3041
rect 5713 2999 5727 3013
rect 5753 2999 5767 3013
rect 5733 2979 5747 2993
rect 5973 3019 5987 3033
rect 6013 3027 6027 3041
rect 6033 3019 6047 3033
rect 6093 3019 6107 3033
rect 6113 3027 6127 3041
rect 6133 3039 6147 3053
rect 6153 3027 6167 3041
rect 6213 3039 6227 3053
rect 6253 3039 6267 3053
rect 6193 3019 6207 3033
rect 6233 3019 6247 3033
rect 6273 3027 6287 3041
rect 6333 3019 6347 3033
rect 6353 3027 6367 3041
rect 6373 3019 6387 3033
rect 6393 3027 6407 3041
rect 6413 3019 6427 3033
rect 6453 3027 6467 3041
rect 6473 3039 6487 3053
rect 6493 3039 6507 3053
rect 6513 3027 6527 3041
rect 6553 3019 6567 3033
rect 6573 3027 6587 3041
rect 6593 3019 6607 3033
rect 6613 2999 6627 3013
rect 2053 2884 2067 2887
rect 3793 2884 3807 2887
rect 193 2816 207 2830
rect 333 2822 347 2836
rect 13 2727 27 2741
rect 33 2739 47 2753
rect 93 2747 107 2761
rect 133 2747 147 2761
rect 113 2727 127 2741
rect 233 2747 247 2761
rect 273 2747 287 2761
rect 333 2784 347 2798
rect 573 2816 587 2830
rect 713 2822 727 2836
rect 353 2719 367 2733
rect 393 2727 407 2741
rect 413 2739 427 2753
rect 473 2747 487 2761
rect 513 2747 527 2761
rect 193 2690 207 2704
rect 333 2690 347 2704
rect 493 2727 507 2741
rect 433 2713 447 2727
rect 473 2713 487 2727
rect 613 2747 627 2761
rect 653 2747 667 2761
rect 713 2784 727 2798
rect 733 2719 747 2733
rect 573 2690 587 2704
rect 793 2747 807 2761
rect 833 2747 847 2761
rect 933 2759 947 2773
rect 953 2767 967 2781
rect 853 2739 867 2753
rect 893 2739 907 2753
rect 713 2690 727 2704
rect 973 2759 987 2773
rect 1013 2759 1027 2773
rect 1033 2767 1047 2781
rect 1053 2759 1067 2773
rect 1093 2727 1107 2741
rect 1113 2739 1127 2753
rect 1153 2747 1167 2761
rect 1173 2739 1187 2753
rect 1193 2747 1207 2761
rect 1213 2739 1227 2753
rect 1233 2747 1247 2761
rect 1293 2747 1307 2761
rect 1453 2767 1467 2781
rect 1593 2793 1607 2807
rect 1313 2739 1327 2753
rect 1333 2727 1347 2741
rect 1353 2739 1367 2753
rect 1393 2739 1407 2753
rect 1473 2747 1487 2761
rect 1413 2727 1427 2741
rect 1493 2739 1507 2753
rect 1513 2747 1527 2761
rect 1533 2747 1547 2761
rect 1573 2747 1587 2761
rect 1553 2727 1567 2741
rect 1613 2759 1627 2773
rect 1633 2767 1647 2781
rect 1613 2713 1627 2727
rect 1653 2759 1667 2773
rect 1693 2747 1707 2761
rect 1793 2767 1807 2781
rect 1733 2747 1747 2761
rect 1813 2747 1827 2761
rect 1713 2727 1727 2741
rect 1833 2739 1847 2753
rect 1853 2747 1867 2761
rect 1893 2747 1907 2761
rect 1873 2727 1887 2741
rect 2053 2873 2067 2884
rect 2213 2816 2227 2830
rect 2353 2822 2367 2836
rect 2033 2767 2047 2781
rect 1933 2739 1947 2753
rect 1973 2747 1987 2761
rect 1993 2739 2007 2753
rect 2013 2747 2027 2761
rect 2093 2747 2107 2761
rect 2113 2739 2127 2753
rect 2133 2727 2147 2741
rect 2153 2739 2167 2753
rect 2253 2747 2267 2761
rect 2293 2747 2307 2761
rect 2353 2784 2367 2798
rect 2413 2759 2427 2773
rect 2433 2767 2447 2781
rect 2373 2719 2387 2733
rect 2213 2690 2227 2704
rect 2453 2759 2467 2773
rect 2653 2816 2667 2830
rect 2793 2822 2807 2836
rect 2493 2727 2507 2741
rect 2513 2739 2527 2753
rect 2573 2739 2587 2753
rect 2353 2690 2367 2704
rect 2593 2727 2607 2741
rect 2693 2747 2707 2761
rect 2733 2747 2747 2761
rect 2793 2784 2807 2798
rect 3093 2822 3107 2836
rect 3233 2816 3247 2830
rect 2913 2767 2927 2781
rect 2853 2747 2867 2761
rect 2873 2739 2887 2753
rect 2893 2747 2907 2761
rect 2973 2747 2987 2761
rect 2813 2719 2827 2733
rect 2653 2690 2667 2704
rect 2793 2690 2807 2704
rect 2993 2739 3007 2753
rect 3013 2727 3027 2741
rect 3033 2739 3047 2753
rect 3093 2784 3107 2798
rect 3073 2719 3087 2733
rect 3153 2747 3167 2761
rect 3193 2747 3207 2761
rect 3093 2690 3107 2704
rect 3793 2873 3807 2884
rect 3533 2767 3547 2781
rect 3793 2793 3807 2807
rect 3753 2767 3767 2781
rect 3293 2727 3307 2741
rect 3313 2739 3327 2753
rect 3353 2747 3367 2761
rect 3373 2739 3387 2753
rect 3393 2747 3407 2761
rect 3233 2690 3247 2704
rect 3413 2739 3427 2753
rect 3433 2747 3447 2761
rect 3473 2747 3487 2761
rect 3493 2739 3507 2753
rect 3513 2747 3527 2761
rect 3593 2747 3607 2761
rect 3613 2739 3627 2753
rect 3633 2747 3647 2761
rect 3653 2739 3667 2753
rect 3673 2747 3687 2761
rect 3693 2747 3707 2761
rect 3713 2739 3727 2753
rect 3733 2747 3747 2761
rect 3913 2773 3927 2787
rect 3813 2747 3827 2761
rect 3833 2739 3847 2753
rect 3853 2747 3867 2761
rect 3813 2713 3827 2727
rect 3873 2739 3887 2753
rect 3893 2747 3907 2761
rect 3893 2713 3907 2727
rect 4033 2853 4047 2867
rect 3933 2739 3947 2753
rect 3973 2747 3987 2761
rect 4013 2747 4027 2761
rect 3953 2727 3967 2741
rect 3993 2727 4007 2741
rect 4013 2713 4027 2727
rect 4293 2813 4307 2827
rect 4053 2747 4067 2761
rect 4293 2767 4307 2781
rect 4093 2747 4107 2761
rect 4153 2747 4167 2761
rect 4073 2727 4087 2741
rect 4173 2739 4187 2753
rect 4193 2727 4207 2741
rect 4213 2739 4227 2753
rect 4233 2747 4247 2761
rect 4253 2739 4267 2753
rect 4273 2747 4287 2761
rect 4393 2787 4407 2801
rect 4473 2816 4487 2830
rect 4613 2822 4627 2836
rect 4353 2759 4367 2773
rect 4373 2767 4387 2781
rect 4413 2767 4427 2781
rect 4333 2733 4347 2747
rect 4513 2747 4527 2761
rect 4553 2747 4567 2761
rect 4613 2784 4627 2798
rect 4633 2719 4647 2733
rect 4673 2727 4687 2741
rect 4693 2739 4707 2753
rect 4733 2747 4747 2761
rect 4873 2767 4887 2781
rect 4773 2747 4787 2761
rect 4813 2747 4827 2761
rect 4473 2690 4487 2704
rect 4613 2690 4627 2704
rect 4753 2727 4767 2741
rect 4833 2739 4847 2753
rect 4853 2747 4867 2761
rect 4933 2747 4947 2761
rect 4773 2713 4787 2727
rect 4813 2713 4827 2727
rect 5193 2773 5207 2787
rect 4973 2747 4987 2761
rect 5013 2747 5027 2761
rect 4953 2727 4967 2741
rect 5033 2739 5047 2753
rect 5053 2747 5067 2761
rect 5073 2739 5087 2753
rect 5093 2747 5107 2761
rect 5113 2739 5127 2753
rect 5133 2727 5147 2741
rect 5153 2739 5167 2753
rect 5173 2747 5187 2761
rect 5193 2753 5207 2767
rect 5213 2747 5227 2761
rect 5353 2767 5367 2781
rect 5253 2747 5267 2761
rect 5293 2747 5307 2761
rect 5313 2739 5327 2753
rect 5333 2747 5347 2761
rect 5393 2753 5407 2767
rect 5353 2733 5367 2747
rect 5413 2747 5427 2761
rect 5433 2739 5447 2753
rect 5453 2747 5467 2761
rect 5473 2739 5487 2753
rect 5493 2747 5507 2761
rect 5613 2816 5627 2830
rect 5753 2822 5767 2836
rect 5533 2739 5547 2753
rect 5553 2727 5567 2741
rect 5653 2747 5667 2761
rect 5693 2747 5707 2761
rect 5753 2784 5767 2798
rect 5813 2739 5827 2753
rect 5833 2747 5847 2761
rect 5773 2719 5787 2733
rect 5873 2739 5887 2753
rect 5893 2747 5907 2761
rect 5933 2739 5947 2753
rect 5953 2747 5967 2761
rect 5613 2690 5627 2704
rect 5753 2690 5767 2704
rect 5993 2739 6007 2753
rect 6013 2747 6027 2761
rect 6053 2739 6067 2753
rect 6073 2747 6087 2761
rect 6113 2739 6127 2753
rect 6133 2747 6147 2761
rect 6193 2747 6207 2761
rect 6213 2759 6227 2773
rect 6253 2747 6267 2761
rect 6293 2739 6307 2753
rect 6333 2739 6347 2753
rect 6353 2747 6367 2761
rect 6493 2822 6507 2836
rect 6633 2816 6647 2830
rect 6393 2759 6407 2773
rect 6413 2747 6427 2761
rect 6493 2784 6507 2798
rect 6473 2719 6487 2733
rect 6553 2747 6567 2761
rect 6593 2747 6607 2761
rect 6493 2690 6507 2704
rect 6633 2690 6647 2704
rect 53 2596 67 2610
rect 193 2596 207 2610
rect 33 2567 47 2581
rect 53 2502 67 2516
rect 113 2539 127 2553
rect 153 2539 167 2553
rect 373 2596 387 2610
rect 273 2539 287 2553
rect 513 2596 527 2610
rect 353 2567 367 2581
rect 313 2539 327 2553
rect 53 2464 67 2478
rect 193 2470 207 2484
rect 373 2502 387 2516
rect 433 2539 447 2553
rect 473 2539 487 2553
rect 1073 2596 1087 2610
rect 593 2539 607 2553
rect 613 2547 627 2561
rect 633 2559 647 2573
rect 653 2547 667 2561
rect 673 2527 687 2541
rect 693 2519 707 2533
rect 713 2527 727 2541
rect 773 2527 787 2541
rect 1213 2596 1227 2610
rect 853 2547 867 2561
rect 793 2519 807 2533
rect 813 2527 827 2541
rect 373 2464 387 2478
rect 513 2470 527 2484
rect 1053 2567 1067 2581
rect 993 2547 1007 2561
rect 1073 2502 1087 2516
rect 1133 2539 1147 2553
rect 1173 2539 1187 2553
rect 1293 2527 1307 2541
rect 1373 2559 1387 2573
rect 1433 2559 1447 2573
rect 1633 2596 1647 2610
rect 1313 2519 1327 2533
rect 1333 2527 1347 2541
rect 1353 2539 1367 2553
rect 1073 2464 1087 2478
rect 1213 2470 1227 2484
rect 1393 2539 1407 2553
rect 1453 2547 1467 2561
rect 1533 2539 1547 2553
rect 1553 2547 1567 2561
rect 1573 2539 1587 2553
rect 1513 2519 1527 2533
rect 1773 2596 1787 2610
rect 1673 2539 1687 2553
rect 1713 2539 1727 2553
rect 1793 2567 1807 2581
rect 1773 2502 1787 2516
rect 1833 2559 1847 2573
rect 1853 2547 1867 2561
rect 1893 2559 1907 2573
rect 2073 2593 2087 2607
rect 1913 2547 1927 2561
rect 1633 2470 1647 2484
rect 1773 2464 1787 2478
rect 1953 2539 1967 2553
rect 1973 2547 1987 2561
rect 2033 2573 2047 2587
rect 1993 2539 2007 2553
rect 2013 2547 2027 2561
rect 2093 2559 2107 2573
rect 2033 2539 2047 2553
rect 2073 2539 2087 2553
rect 2113 2539 2127 2553
rect 2153 2547 2167 2561
rect 2173 2539 2187 2553
rect 2213 2547 2227 2561
rect 2233 2539 2247 2553
rect 2273 2547 2287 2561
rect 2293 2539 2307 2553
rect 2433 2596 2447 2610
rect 2333 2547 2347 2561
rect 2353 2539 2367 2553
rect 2573 2596 2587 2610
rect 2473 2539 2487 2553
rect 2513 2539 2527 2553
rect 2593 2567 2607 2581
rect 2573 2502 2587 2516
rect 2633 2547 2647 2561
rect 2653 2539 2667 2553
rect 2693 2547 2707 2561
rect 2793 2559 2807 2573
rect 2433 2470 2447 2484
rect 2573 2464 2587 2478
rect 2713 2539 2727 2553
rect 2773 2539 2787 2553
rect 2813 2539 2827 2553
rect 2853 2539 2867 2553
rect 2873 2547 2887 2561
rect 2913 2539 2927 2553
rect 2933 2547 2947 2561
rect 2973 2539 2987 2553
rect 2993 2547 3007 2561
rect 3173 2596 3187 2610
rect 3013 2539 3027 2553
rect 3033 2547 3047 2561
rect 3053 2539 3067 2553
rect 3093 2547 3107 2561
rect 3113 2559 3127 2573
rect 3313 2596 3327 2610
rect 3213 2539 3227 2553
rect 3253 2539 3267 2553
rect 3333 2567 3347 2581
rect 3313 2502 3327 2516
rect 3393 2559 3407 2573
rect 3373 2539 3387 2553
rect 3413 2539 3427 2553
rect 3473 2527 3487 2541
rect 3533 2559 3547 2573
rect 3553 2547 3567 2561
rect 3493 2519 3507 2533
rect 3513 2527 3527 2541
rect 3173 2470 3187 2484
rect 3313 2464 3327 2478
rect 3613 2533 3627 2547
rect 3593 2519 3607 2533
rect 3633 2519 3647 2533
rect 3653 2527 3667 2541
rect 3673 2533 3687 2547
rect 3613 2499 3627 2513
rect 3593 2473 3607 2487
rect 3693 2519 3707 2533
rect 3733 2519 3747 2533
rect 3753 2527 3767 2541
rect 3813 2527 3827 2541
rect 3893 2539 3907 2553
rect 3913 2547 3927 2561
rect 3953 2553 3967 2567
rect 3933 2539 3947 2553
rect 3713 2499 3727 2513
rect 3693 2473 3707 2487
rect 3833 2519 3847 2533
rect 3873 2519 3887 2533
rect 3853 2499 3867 2513
rect 3953 2519 3967 2533
rect 3993 2547 4007 2561
rect 4013 2559 4027 2573
rect 4033 2547 4047 2561
rect 4333 2596 4347 2610
rect 4133 2559 4147 2573
rect 4053 2539 4067 2553
rect 4113 2539 4127 2553
rect 4033 2513 4047 2527
rect 4153 2539 4167 2553
rect 4193 2539 4207 2553
rect 4213 2547 4227 2561
rect 4233 2539 4247 2553
rect 4253 2547 4267 2561
rect 4273 2539 4287 2553
rect 4473 2596 4487 2610
rect 4373 2539 4387 2553
rect 4413 2539 4427 2553
rect 4493 2567 4507 2581
rect 4473 2502 4487 2516
rect 4553 2547 4567 2561
rect 4573 2559 4587 2573
rect 4333 2470 4347 2484
rect 4473 2464 4487 2478
rect 4613 2539 4627 2553
rect 4633 2547 4647 2561
rect 4653 2539 4667 2553
rect 4673 2547 4687 2561
rect 4693 2539 4707 2553
rect 4713 2547 4727 2561
rect 4733 2539 4747 2553
rect 4873 2596 4887 2610
rect 5013 2596 5027 2610
rect 4853 2567 4867 2581
rect 4773 2547 4787 2561
rect 4793 2539 4807 2553
rect 4873 2502 4887 2516
rect 4933 2539 4947 2553
rect 4973 2539 4987 2553
rect 5073 2559 5087 2573
rect 5093 2547 5107 2561
rect 4873 2464 4887 2478
rect 5013 2470 5027 2484
rect 5133 2539 5147 2553
rect 5153 2547 5167 2561
rect 5173 2539 5187 2553
rect 5193 2547 5207 2561
rect 5213 2539 5227 2553
rect 5253 2539 5267 2553
rect 5273 2547 5287 2561
rect 5373 2559 5387 2573
rect 5293 2539 5307 2553
rect 5353 2539 5367 2553
rect 5313 2519 5327 2533
rect 5473 2559 5487 2573
rect 5393 2539 5407 2553
rect 5453 2539 5467 2553
rect 5493 2539 5507 2553
rect 5533 2547 5547 2561
rect 5673 2547 5687 2561
rect 5753 2559 5767 2573
rect 5733 2539 5747 2553
rect 5773 2539 5787 2553
rect 5793 2539 5807 2553
rect 5813 2547 5827 2561
rect 5833 2539 5847 2553
rect 5913 2539 5927 2553
rect 5933 2547 5947 2561
rect 6113 2596 6127 2610
rect 6253 2596 6267 2610
rect 5953 2539 5967 2553
rect 5973 2547 5987 2561
rect 5993 2539 6007 2553
rect 6033 2547 6047 2561
rect 6053 2559 6067 2573
rect 6093 2567 6107 2581
rect 5853 2519 5867 2533
rect 6113 2502 6127 2516
rect 6173 2539 6187 2553
rect 6213 2539 6227 2553
rect 6333 2539 6347 2553
rect 6353 2547 6367 2561
rect 6373 2539 6387 2553
rect 6393 2547 6407 2561
rect 6413 2539 6427 2553
rect 6433 2547 6447 2561
rect 6473 2547 6487 2561
rect 6513 2559 6527 2573
rect 6533 2547 6547 2561
rect 6113 2464 6127 2478
rect 6253 2470 6267 2484
rect 6573 2539 6587 2553
rect 6593 2547 6607 2561
rect 6613 2539 6627 2553
rect 6633 2547 6647 2561
rect 6653 2539 6667 2553
rect 53 2336 67 2350
rect 193 2342 207 2356
rect 93 2267 107 2281
rect 133 2267 147 2281
rect 193 2304 207 2318
rect 213 2239 227 2253
rect 53 2210 67 2224
rect 273 2267 287 2281
rect 313 2267 327 2281
rect 353 2267 367 2281
rect 193 2210 207 2224
rect 373 2259 387 2273
rect 413 2259 427 2273
rect 473 2267 487 2281
rect 593 2287 607 2301
rect 513 2267 527 2281
rect 533 2267 547 2281
rect 433 2247 447 2261
rect 493 2247 507 2261
rect 553 2259 567 2273
rect 573 2267 587 2281
rect 653 2267 667 2281
rect 673 2279 687 2293
rect 753 2307 767 2321
rect 733 2287 747 2301
rect 773 2287 787 2301
rect 953 2342 967 2356
rect 1093 2336 1107 2350
rect 713 2267 727 2281
rect 793 2279 807 2293
rect 833 2279 847 2293
rect 853 2287 867 2301
rect 873 2279 887 2293
rect 953 2304 967 2318
rect 933 2239 947 2253
rect 1013 2267 1027 2281
rect 1053 2267 1067 2281
rect 953 2210 967 2224
rect 1253 2336 1267 2350
rect 1393 2342 1407 2356
rect 1153 2247 1167 2261
rect 1173 2259 1187 2273
rect 1093 2210 1107 2224
rect 1293 2267 1307 2281
rect 1333 2267 1347 2281
rect 1393 2304 1407 2318
rect 1693 2287 1707 2301
rect 1473 2259 1487 2273
rect 1513 2267 1527 2281
rect 1413 2239 1427 2253
rect 1253 2210 1267 2224
rect 1393 2210 1407 2224
rect 1493 2247 1507 2261
rect 1533 2259 1547 2273
rect 1553 2267 1567 2281
rect 1573 2259 1587 2273
rect 1593 2267 1607 2281
rect 1633 2267 1647 2281
rect 1653 2259 1667 2273
rect 1673 2267 1687 2281
rect 1753 2267 1767 2281
rect 1793 2267 1807 2281
rect 1833 2267 1847 2281
rect 1873 2267 1887 2281
rect 1913 2267 1927 2281
rect 1773 2247 1787 2261
rect 1853 2247 1867 2261
rect 1933 2259 1947 2273
rect 1953 2267 1967 2281
rect 1973 2259 1987 2273
rect 1993 2267 2007 2281
rect 2113 2336 2127 2350
rect 2253 2342 2267 2356
rect 2033 2259 2047 2273
rect 2053 2247 2067 2261
rect 2153 2267 2167 2281
rect 2193 2267 2207 2281
rect 2253 2304 2267 2318
rect 2453 2333 2467 2347
rect 2333 2267 2347 2281
rect 2273 2239 2287 2253
rect 2113 2210 2127 2224
rect 2253 2210 2267 2224
rect 2453 2287 2467 2301
rect 2373 2267 2387 2281
rect 2393 2267 2407 2281
rect 2353 2247 2367 2261
rect 2413 2259 2427 2273
rect 2433 2267 2447 2281
rect 2553 2307 2567 2321
rect 2913 2342 2927 2356
rect 3053 2336 3067 2350
rect 2513 2279 2527 2293
rect 2533 2287 2547 2301
rect 2573 2287 2587 2301
rect 2593 2293 2607 2307
rect 2553 2273 2567 2287
rect 2593 2273 2607 2287
rect 2753 2287 2767 2301
rect 2613 2267 2627 2281
rect 2593 2253 2607 2267
rect 2513 2213 2527 2227
rect 2633 2259 2647 2273
rect 2653 2247 2667 2261
rect 2673 2259 2687 2273
rect 2693 2267 2707 2281
rect 2713 2259 2727 2273
rect 2733 2267 2747 2281
rect 2813 2267 2827 2281
rect 2853 2267 2867 2281
rect 2833 2247 2847 2261
rect 2913 2304 2927 2318
rect 2893 2239 2907 2253
rect 2973 2267 2987 2281
rect 3013 2267 3027 2281
rect 2913 2210 2927 2224
rect 3173 2287 3187 2301
rect 3113 2267 3127 2281
rect 3133 2259 3147 2273
rect 3153 2267 3167 2281
rect 3233 2267 3247 2281
rect 3253 2259 3267 2273
rect 3273 2267 3287 2281
rect 3293 2259 3307 2273
rect 3313 2267 3327 2281
rect 3353 2267 3367 2281
rect 3393 2267 3407 2281
rect 3593 2336 3607 2350
rect 3733 2342 3747 2356
rect 3453 2293 3467 2307
rect 3373 2247 3387 2261
rect 3433 2259 3447 2273
rect 3053 2210 3067 2224
rect 3453 2247 3467 2261
rect 3493 2267 3507 2281
rect 3533 2267 3547 2281
rect 3513 2247 3527 2261
rect 3493 2233 3507 2247
rect 3633 2267 3647 2281
rect 3673 2267 3687 2281
rect 3733 2304 3747 2318
rect 3893 2307 3907 2321
rect 3793 2279 3807 2293
rect 3813 2287 3827 2301
rect 3753 2239 3767 2253
rect 3593 2210 3607 2224
rect 3833 2279 3847 2293
rect 3873 2287 3887 2301
rect 3913 2287 3927 2301
rect 3933 2279 3947 2293
rect 3973 2259 3987 2273
rect 3993 2267 4007 2281
rect 3733 2210 3747 2224
rect 4033 2259 4047 2273
rect 4053 2267 4067 2281
rect 4093 2259 4107 2273
rect 4113 2267 4127 2281
rect 4153 2259 4167 2273
rect 4173 2267 4187 2281
rect 4213 2259 4227 2273
rect 4233 2267 4247 2281
rect 4273 2259 4287 2273
rect 4293 2267 4307 2281
rect 4333 2267 4347 2281
rect 4373 2267 4387 2281
rect 4433 2267 4447 2281
rect 4473 2267 4487 2281
rect 4453 2247 4467 2261
rect 4493 2259 4507 2273
rect 4513 2267 4527 2281
rect 4553 2259 4567 2273
rect 4573 2267 4587 2281
rect 4633 2267 4647 2281
rect 4653 2259 4667 2273
rect 4693 2267 4707 2281
rect 4713 2259 4727 2273
rect 4733 2259 4747 2273
rect 4753 2267 4767 2281
rect 4793 2259 4807 2273
rect 4813 2267 4827 2281
rect 4853 2267 4867 2281
rect 4893 2267 4907 2281
rect 4873 2247 4887 2261
rect 4933 2259 4947 2273
rect 4953 2267 4967 2281
rect 4993 2259 5007 2273
rect 5013 2267 5027 2281
rect 5073 2267 5087 2281
rect 5093 2259 5107 2273
rect 5113 2247 5127 2261
rect 5133 2259 5147 2273
rect 5153 2247 5167 2261
rect 5173 2259 5187 2273
rect 5213 2267 5227 2281
rect 5233 2259 5247 2273
rect 5253 2267 5267 2281
rect 5273 2259 5287 2273
rect 5293 2267 5307 2281
rect 5353 2267 5367 2281
rect 5373 2259 5387 2273
rect 5413 2267 5427 2281
rect 5433 2259 5447 2273
rect 5453 2259 5467 2273
rect 5473 2267 5487 2281
rect 5513 2259 5527 2273
rect 5533 2267 5547 2281
rect 5573 2259 5587 2273
rect 5593 2267 5607 2281
rect 5793 2333 5807 2347
rect 5753 2307 5767 2321
rect 5633 2259 5647 2273
rect 5653 2267 5667 2281
rect 5713 2279 5727 2293
rect 5733 2287 5747 2301
rect 5773 2287 5787 2301
rect 5853 2307 5867 2321
rect 5793 2273 5807 2287
rect 5813 2279 5827 2293
rect 5833 2287 5847 2301
rect 5873 2287 5887 2301
rect 5913 2259 5927 2273
rect 5973 2267 5987 2281
rect 5933 2247 5947 2261
rect 5993 2259 6007 2273
rect 6013 2267 6027 2281
rect 6033 2259 6047 2273
rect 6053 2267 6067 2281
rect 6093 2267 6107 2281
rect 6113 2259 6127 2273
rect 6153 2267 6167 2281
rect 6173 2259 6187 2273
rect 6213 2267 6227 2281
rect 6233 2259 6247 2273
rect 6273 2267 6287 2281
rect 6433 2333 6447 2347
rect 6433 2287 6447 2301
rect 6293 2259 6307 2273
rect 6313 2247 6327 2261
rect 6333 2259 6347 2273
rect 6373 2267 6387 2281
rect 6393 2259 6407 2273
rect 6413 2267 6427 2281
rect 6473 2279 6487 2293
rect 6493 2287 6507 2301
rect 6473 2233 6487 2247
rect 6513 2279 6527 2293
rect 6553 2259 6567 2273
rect 6573 2247 6587 2261
rect 6593 2259 6607 2273
rect 6613 2267 6627 2281
rect 6653 2247 6667 2261
rect 6673 2259 6687 2273
rect 73 2093 87 2107
rect 53 2079 67 2093
rect 33 2059 47 2073
rect 73 2059 87 2073
rect 113 2047 127 2061
rect 173 2093 187 2107
rect 133 2039 147 2053
rect 153 2047 167 2061
rect 93 1993 107 2007
rect 153 2013 167 2027
rect 273 2093 287 2107
rect 193 2047 207 2061
rect 213 2039 227 2053
rect 253 2039 267 2053
rect 233 2019 247 2033
rect 253 1993 267 2007
rect 373 2113 387 2127
rect 293 2047 307 2061
rect 313 2039 327 2053
rect 353 2039 367 2053
rect 333 2019 347 2033
rect 353 1993 367 2007
rect 393 2047 407 2061
rect 513 2113 527 2127
rect 573 2113 587 2127
rect 413 2039 427 2053
rect 433 2047 447 2061
rect 453 2039 467 2053
rect 493 2039 507 2053
rect 513 2047 527 2061
rect 473 2019 487 2033
rect 533 2033 547 2047
rect 573 2093 587 2107
rect 593 2079 607 2093
rect 573 2059 587 2073
rect 613 2059 627 2073
rect 633 2059 647 2073
rect 653 2067 667 2081
rect 673 2059 687 2073
rect 853 2079 867 2093
rect 693 2039 707 2053
rect 733 2039 747 2053
rect 773 2039 787 2053
rect 793 2047 807 2061
rect 833 2059 847 2073
rect 753 2019 767 2033
rect 873 2059 887 2073
rect 933 2047 947 2061
rect 993 2067 1007 2081
rect 953 2039 967 2053
rect 973 2047 987 2061
rect 1013 2059 1027 2073
rect 1153 2116 1167 2130
rect 1053 2067 1067 2081
rect 1073 2059 1087 2073
rect 1293 2116 1307 2130
rect 1193 2059 1207 2073
rect 1233 2059 1247 2073
rect 1313 2087 1327 2101
rect 1293 2022 1307 2036
rect 1353 2079 1367 2093
rect 1373 2067 1387 2081
rect 1153 1990 1167 2004
rect 1293 1984 1307 1998
rect 1413 2059 1427 2073
rect 1433 2067 1447 2081
rect 1493 2093 1507 2107
rect 1453 2059 1467 2073
rect 1473 2067 1487 2081
rect 1493 2059 1507 2073
rect 1573 2059 1587 2073
rect 1593 2067 1607 2081
rect 1613 2059 1627 2073
rect 1673 2059 1687 2073
rect 1693 2067 1707 2081
rect 1773 2079 1787 2093
rect 1713 2059 1727 2073
rect 1753 2059 1767 2073
rect 1513 2033 1527 2047
rect 1553 2039 1567 2053
rect 1653 2039 1667 2053
rect 1793 2059 1807 2073
rect 1853 2059 1867 2073
rect 1873 2067 1887 2081
rect 1893 2059 1907 2073
rect 1933 2059 1947 2073
rect 1953 2067 1967 2081
rect 1833 2039 1847 2053
rect 2193 2116 2207 2130
rect 1993 2059 2007 2073
rect 2013 2067 2027 2081
rect 2053 2059 2067 2073
rect 2073 2067 2087 2081
rect 2113 2059 2127 2073
rect 2133 2067 2147 2081
rect 2333 2116 2347 2130
rect 2233 2059 2247 2073
rect 2273 2059 2287 2073
rect 2353 2087 2367 2101
rect 2333 2022 2347 2036
rect 2433 2059 2447 2073
rect 2453 2067 2467 2081
rect 2513 2079 2527 2093
rect 2473 2059 2487 2073
rect 2493 2059 2507 2073
rect 2413 2039 2427 2053
rect 2533 2059 2547 2073
rect 2673 2067 2687 2081
rect 2593 2047 2607 2061
rect 2693 2059 2707 2073
rect 2193 1990 2207 2004
rect 2333 1984 2347 1998
rect 2613 2039 2627 2053
rect 2653 2039 2667 2053
rect 2733 2067 2747 2081
rect 2633 2019 2647 2033
rect 2753 2059 2767 2073
rect 2813 2059 2827 2073
rect 2833 2067 2847 2081
rect 2873 2059 2887 2073
rect 2893 2067 2907 2081
rect 2913 2079 2927 2093
rect 2933 2067 2947 2081
rect 2973 2093 2987 2107
rect 2953 2053 2967 2067
rect 2973 2059 2987 2073
rect 2993 2067 3007 2081
rect 3013 2059 3027 2073
rect 3033 2067 3047 2081
rect 3053 2059 3067 2073
rect 3113 2059 3127 2073
rect 3133 2067 3147 2081
rect 3153 2079 3167 2093
rect 3173 2067 3187 2081
rect 3193 2079 3207 2093
rect 3213 2067 3227 2081
rect 3253 2059 3267 2073
rect 3273 2067 3287 2081
rect 3293 2059 3307 2073
rect 3313 2067 3327 2081
rect 3393 2079 3407 2093
rect 3333 2059 3347 2073
rect 3373 2059 3387 2073
rect 3493 2116 3507 2130
rect 3413 2059 3427 2073
rect 3633 2116 3647 2130
rect 3533 2059 3547 2073
rect 3573 2059 3587 2073
rect 3653 2087 3667 2101
rect 3633 2022 3647 2036
rect 3493 1990 3507 2004
rect 3633 1984 3647 1998
rect 3713 2093 3727 2107
rect 3753 2093 3767 2107
rect 3793 2093 3807 2107
rect 3733 2079 3747 2093
rect 3713 2059 3727 2073
rect 3753 2059 3767 2073
rect 3793 2059 3807 2073
rect 3813 2067 3827 2081
rect 3873 2093 3887 2107
rect 3833 2059 3847 2073
rect 3853 2067 3867 2081
rect 3873 2059 3887 2073
rect 3913 2067 3927 2081
rect 3933 2079 3947 2093
rect 3693 1993 3707 2007
rect 3893 2013 3907 2027
rect 3953 2059 3967 2073
rect 3973 2067 3987 2081
rect 3993 2059 4007 2073
rect 4033 2053 4047 2067
rect 4013 2039 4027 2053
rect 4053 2047 4067 2061
rect 4253 2116 4267 2130
rect 4173 2079 4187 2093
rect 4073 2039 4087 2053
rect 4093 2047 4107 2061
rect 4153 2059 4167 2073
rect 4053 2013 4067 2027
rect 4193 2059 4207 2073
rect 4393 2116 4407 2130
rect 4293 2059 4307 2073
rect 4333 2059 4347 2073
rect 4413 2087 4427 2101
rect 4393 2022 4407 2036
rect 4453 2079 4467 2093
rect 4493 2093 4507 2107
rect 4473 2067 4487 2081
rect 4253 1990 4267 2004
rect 4393 1984 4407 1998
rect 4513 2059 4527 2073
rect 4533 2067 4547 2081
rect 4553 2059 4567 2073
rect 4573 2067 4587 2081
rect 4653 2079 4667 2093
rect 4593 2059 4607 2073
rect 4633 2059 4647 2073
rect 4493 2033 4507 2047
rect 4673 2059 4687 2073
rect 4753 2059 4767 2073
rect 4773 2067 4787 2081
rect 4853 2079 4867 2093
rect 4793 2059 4807 2073
rect 4833 2059 4847 2073
rect 4733 2039 4747 2053
rect 4873 2059 4887 2073
rect 4893 2059 4907 2073
rect 4913 2067 4927 2081
rect 4933 2059 4947 2073
rect 4953 2067 4967 2081
rect 4973 2059 4987 2073
rect 5033 2047 5047 2061
rect 5133 2079 5147 2093
rect 5173 2079 5187 2093
rect 5053 2039 5067 2053
rect 5073 2047 5087 2061
rect 5113 2059 5127 2073
rect 5153 2059 5167 2073
rect 5193 2059 5207 2073
rect 5233 2067 5247 2081
rect 5293 2059 5307 2073
rect 5313 2067 5327 2081
rect 5333 2059 5347 2073
rect 5353 2067 5367 2081
rect 5373 2059 5387 2073
rect 5393 2059 5407 2073
rect 5413 2067 5427 2081
rect 5573 2093 5587 2107
rect 5433 2059 5447 2073
rect 5453 2067 5467 2081
rect 5553 2079 5567 2093
rect 5473 2059 5487 2073
rect 5533 2059 5547 2073
rect 5573 2059 5587 2073
rect 5613 2059 5627 2073
rect 5633 2067 5647 2081
rect 5713 2093 5727 2107
rect 5653 2059 5667 2073
rect 5673 2067 5687 2081
rect 5693 2059 5707 2073
rect 5593 2033 5607 2047
rect 5893 2116 5907 2130
rect 5733 2067 5747 2081
rect 5753 2079 5767 2093
rect 5713 2033 5727 2047
rect 5773 2047 5787 2061
rect 6033 2116 6047 2130
rect 5873 2087 5887 2101
rect 5793 2039 5807 2053
rect 5813 2047 5827 2061
rect 5893 2022 5907 2036
rect 5953 2059 5967 2073
rect 5993 2059 6007 2073
rect 5893 1984 5907 1998
rect 6033 1990 6047 2004
rect 6133 2116 6147 2130
rect 6273 2116 6287 2130
rect 6173 2059 6187 2073
rect 6213 2059 6227 2073
rect 6293 2087 6307 2101
rect 6273 2022 6287 2036
rect 6333 2067 6347 2081
rect 6353 2059 6367 2073
rect 6393 2067 6407 2081
rect 6133 1990 6147 2004
rect 6273 1984 6287 1998
rect 6413 2059 6427 2073
rect 6453 2067 6467 2081
rect 6473 2079 6487 2093
rect 6493 2067 6507 2081
rect 6513 2059 6527 2073
rect 6553 2059 6567 2073
rect 6573 2067 6587 2081
rect 6593 2059 6607 2073
rect 6613 2039 6627 2053
rect 113 1862 127 1876
rect 253 1856 267 1870
rect 33 1779 47 1793
rect 53 1767 67 1781
rect 113 1824 127 1838
rect 93 1759 107 1773
rect 173 1787 187 1801
rect 213 1787 227 1801
rect 113 1730 127 1744
rect 313 1787 327 1801
rect 353 1787 367 1801
rect 413 1787 427 1801
rect 333 1767 347 1781
rect 253 1730 267 1744
rect 453 1787 467 1801
rect 673 1862 687 1876
rect 813 1856 827 1870
rect 553 1807 567 1821
rect 433 1767 447 1781
rect 493 1779 507 1793
rect 573 1787 587 1801
rect 513 1767 527 1781
rect 593 1779 607 1793
rect 613 1787 627 1801
rect 673 1824 687 1838
rect 653 1759 667 1773
rect 733 1787 747 1801
rect 773 1787 787 1801
rect 673 1730 687 1744
rect 933 1827 947 1841
rect 893 1799 907 1813
rect 913 1807 927 1821
rect 953 1807 967 1821
rect 973 1787 987 1801
rect 813 1730 827 1744
rect 1013 1799 1027 1813
rect 1033 1787 1047 1801
rect 1233 1853 1247 1867
rect 1193 1807 1207 1821
rect 1073 1767 1087 1781
rect 1093 1779 1107 1793
rect 1133 1787 1147 1801
rect 1153 1779 1167 1793
rect 1173 1787 1187 1801
rect 1193 1773 1207 1787
rect 1253 1799 1267 1813
rect 1273 1807 1287 1821
rect 1373 1827 1387 1841
rect 1293 1799 1307 1813
rect 1333 1799 1347 1813
rect 1353 1807 1367 1821
rect 1393 1807 1407 1821
rect 1513 1856 1527 1870
rect 1653 1862 1667 1876
rect 1413 1767 1427 1781
rect 1433 1779 1447 1793
rect 1553 1787 1567 1801
rect 1593 1787 1607 1801
rect 1653 1824 1667 1838
rect 2113 1862 2127 1876
rect 2253 1856 2267 1870
rect 1673 1759 1687 1773
rect 1713 1767 1727 1781
rect 1733 1779 1747 1793
rect 1773 1787 1787 1801
rect 1793 1779 1807 1793
rect 1813 1787 1827 1801
rect 1513 1730 1527 1744
rect 1653 1730 1667 1744
rect 1833 1779 1847 1793
rect 1853 1787 1867 1801
rect 1893 1787 1907 1801
rect 2033 1807 2047 1821
rect 1933 1787 1947 1801
rect 1973 1787 1987 1801
rect 1913 1767 1927 1781
rect 1993 1779 2007 1793
rect 2013 1787 2027 1801
rect 2113 1824 2127 1838
rect 2093 1759 2107 1773
rect 2173 1787 2187 1801
rect 2213 1787 2227 1801
rect 2113 1730 2127 1744
rect 2333 1787 2347 1801
rect 2353 1779 2367 1793
rect 2373 1787 2387 1801
rect 2393 1779 2407 1793
rect 2413 1787 2427 1801
rect 2613 1862 2627 1876
rect 2753 1856 2767 1870
rect 2433 1767 2447 1781
rect 2453 1779 2467 1793
rect 2493 1787 2507 1801
rect 2533 1787 2547 1801
rect 2253 1730 2267 1744
rect 2513 1767 2527 1781
rect 2613 1824 2627 1838
rect 2593 1759 2607 1773
rect 2673 1787 2687 1801
rect 2713 1787 2727 1801
rect 2613 1730 2627 1744
rect 2833 1827 2847 1841
rect 2813 1807 2827 1821
rect 2853 1807 2867 1821
rect 2873 1799 2887 1813
rect 2933 1807 2947 1821
rect 2753 1730 2767 1744
rect 2953 1787 2967 1801
rect 2973 1779 2987 1793
rect 2993 1787 3007 1801
rect 3013 1787 3027 1801
rect 3373 1833 3387 1847
rect 3053 1787 3067 1801
rect 3113 1787 3127 1801
rect 3033 1767 3047 1781
rect 3133 1779 3147 1793
rect 3153 1767 3167 1781
rect 3173 1779 3187 1793
rect 3213 1787 3227 1801
rect 3233 1779 3247 1793
rect 3253 1767 3267 1781
rect 3273 1779 3287 1793
rect 3313 1787 3327 1801
rect 3353 1787 3367 1801
rect 3393 1799 3407 1813
rect 3413 1807 3427 1821
rect 3373 1753 3387 1767
rect 3433 1799 3447 1813
rect 3453 1787 3467 1801
rect 3493 1787 3507 1801
rect 3533 1799 3547 1813
rect 3553 1807 3567 1821
rect 3473 1767 3487 1781
rect 3573 1799 3587 1813
rect 3673 1807 3687 1821
rect 3713 1813 3727 1827
rect 3613 1787 3627 1801
rect 3633 1779 3647 1793
rect 3653 1787 3667 1801
rect 3673 1773 3687 1787
rect 3733 1799 3747 1813
rect 3753 1807 3767 1821
rect 3773 1799 3787 1813
rect 4273 1853 4287 1867
rect 3853 1799 3867 1813
rect 3873 1807 3887 1821
rect 3813 1779 3827 1793
rect 3833 1767 3847 1781
rect 3893 1799 3907 1813
rect 3933 1787 3947 1801
rect 3973 1787 3987 1801
rect 4013 1787 4027 1801
rect 3953 1767 3967 1781
rect 4033 1779 4047 1793
rect 4053 1787 4067 1801
rect 4073 1779 4087 1793
rect 4093 1787 4107 1801
rect 4153 1787 4167 1801
rect 4273 1807 4287 1821
rect 4473 1873 4487 1887
rect 4453 1853 4467 1867
rect 4193 1787 4207 1801
rect 4213 1787 4227 1801
rect 4173 1767 4187 1781
rect 4233 1779 4247 1793
rect 4253 1787 4267 1801
rect 4293 1793 4307 1807
rect 4373 1813 4387 1827
rect 4313 1779 4327 1793
rect 4353 1779 4367 1793
rect 4453 1807 4467 1821
rect 4393 1787 4407 1801
rect 4413 1779 4427 1793
rect 4433 1787 4447 1801
rect 4393 1753 4407 1767
rect 4473 1753 4487 1767
rect 4513 1787 4527 1801
rect 4553 1787 4567 1801
rect 4593 1787 4607 1801
rect 4533 1767 4547 1781
rect 4613 1779 4627 1793
rect 4633 1787 4647 1801
rect 4513 1753 4527 1767
rect 4653 1779 4667 1793
rect 4673 1787 4687 1801
rect 4793 1862 4807 1876
rect 4933 1856 4947 1870
rect 4713 1779 4727 1793
rect 4733 1767 4747 1781
rect 4793 1824 4807 1838
rect 4773 1759 4787 1773
rect 4853 1787 4867 1801
rect 4893 1787 4907 1801
rect 4793 1730 4807 1744
rect 4993 1779 5007 1793
rect 5013 1767 5027 1781
rect 5033 1779 5047 1793
rect 5053 1787 5067 1801
rect 5093 1787 5107 1801
rect 5293 1827 5307 1841
rect 5233 1807 5247 1821
rect 5273 1807 5287 1821
rect 5313 1807 5327 1821
rect 5133 1787 5147 1801
rect 5173 1787 5187 1801
rect 5113 1767 5127 1781
rect 5193 1779 5207 1793
rect 5213 1787 5227 1801
rect 5333 1799 5347 1813
rect 4933 1730 4947 1744
rect 5373 1787 5387 1801
rect 5413 1787 5427 1801
rect 5593 1807 5607 1821
rect 5473 1779 5487 1793
rect 5533 1787 5547 1801
rect 5493 1767 5507 1781
rect 5553 1779 5567 1793
rect 5613 1787 5627 1801
rect 5633 1779 5647 1793
rect 5653 1787 5667 1801
rect 5673 1799 5687 1813
rect 5693 1807 5707 1821
rect 5733 1813 5747 1827
rect 5713 1799 5727 1813
rect 5773 1787 5787 1801
rect 5793 1779 5807 1793
rect 5813 1787 5827 1801
rect 5773 1753 5787 1767
rect 5833 1779 5847 1793
rect 5853 1787 5867 1801
rect 5873 1787 5887 1801
rect 5973 1807 5987 1821
rect 5913 1787 5927 1801
rect 5993 1787 6007 1801
rect 6013 1779 6027 1793
rect 6033 1787 6047 1801
rect 6073 1787 6087 1801
rect 6093 1779 6107 1793
rect 6113 1787 6127 1801
rect 6133 1779 6147 1793
rect 6153 1787 6167 1801
rect 6173 1779 6187 1793
rect 6193 1787 6207 1801
rect 6233 1779 6247 1793
rect 6253 1787 6267 1801
rect 6293 1779 6307 1793
rect 6313 1787 6327 1801
rect 6353 1779 6367 1793
rect 6373 1787 6387 1801
rect 6533 1807 6547 1821
rect 6413 1767 6427 1781
rect 6433 1779 6447 1793
rect 6473 1787 6487 1801
rect 6493 1779 6507 1793
rect 6513 1787 6527 1801
rect 6593 1799 6607 1813
rect 6613 1807 6627 1821
rect 6633 1799 6647 1813
rect 333 1636 347 1650
rect 53 1599 67 1613
rect 33 1579 47 1593
rect 73 1579 87 1593
rect 113 1587 127 1601
rect 253 1587 267 1601
rect 473 1636 487 1650
rect 373 1579 387 1593
rect 413 1579 427 1593
rect 493 1607 507 1621
rect 473 1542 487 1556
rect 553 1587 567 1601
rect 573 1599 587 1613
rect 333 1510 347 1524
rect 473 1504 487 1518
rect 693 1587 707 1601
rect 713 1599 727 1613
rect 733 1587 747 1601
rect 833 1636 847 1650
rect 593 1559 607 1573
rect 633 1559 647 1573
rect 653 1567 667 1581
rect 753 1579 767 1593
rect 613 1539 627 1553
rect 973 1636 987 1650
rect 873 1579 887 1593
rect 913 1579 927 1593
rect 993 1607 1007 1621
rect 973 1542 987 1556
rect 1053 1587 1067 1601
rect 1073 1599 1087 1613
rect 833 1510 847 1524
rect 973 1504 987 1518
rect 1093 1579 1107 1593
rect 1113 1587 1127 1601
rect 1133 1579 1147 1593
rect 1153 1587 1167 1601
rect 1173 1579 1187 1593
rect 1253 1579 1267 1593
rect 1273 1587 1287 1601
rect 1353 1599 1367 1613
rect 1293 1579 1307 1593
rect 1333 1579 1347 1593
rect 1233 1559 1247 1573
rect 1373 1579 1387 1593
rect 1413 1579 1427 1593
rect 1433 1587 1447 1601
rect 1473 1579 1487 1593
rect 1493 1587 1507 1601
rect 1533 1579 1547 1593
rect 1553 1587 1567 1601
rect 1793 1636 1807 1650
rect 1933 1636 1947 1650
rect 1593 1579 1607 1593
rect 1613 1587 1627 1601
rect 1653 1579 1667 1593
rect 1673 1587 1687 1601
rect 1773 1607 1787 1621
rect 1713 1579 1727 1593
rect 1733 1587 1747 1601
rect 1793 1542 1807 1556
rect 1853 1579 1867 1593
rect 1893 1579 1907 1593
rect 1993 1587 2007 1601
rect 2013 1579 2027 1593
rect 2053 1587 2067 1601
rect 2113 1599 2127 1613
rect 1793 1504 1807 1518
rect 1933 1510 1947 1524
rect 2073 1579 2087 1593
rect 2133 1587 2147 1601
rect 2173 1579 2187 1593
rect 2193 1587 2207 1601
rect 2253 1613 2267 1627
rect 2293 1613 2307 1627
rect 2213 1579 2227 1593
rect 2233 1587 2247 1601
rect 2313 1599 2327 1613
rect 2253 1579 2267 1593
rect 2293 1579 2307 1593
rect 2333 1579 2347 1593
rect 2413 1579 2427 1593
rect 2433 1587 2447 1601
rect 2453 1579 2467 1593
rect 2493 1579 2507 1593
rect 2393 1559 2407 1573
rect 2573 1599 2587 1613
rect 2533 1579 2547 1593
rect 2553 1579 2567 1593
rect 2593 1579 2607 1593
rect 2653 1567 2667 1581
rect 2673 1559 2687 1573
rect 2693 1567 2707 1581
rect 2713 1567 2727 1581
rect 2733 1559 2747 1573
rect 2753 1567 2767 1581
rect 2813 1579 2827 1593
rect 2833 1587 2847 1601
rect 3113 1636 3127 1650
rect 2873 1579 2887 1593
rect 2893 1587 2907 1601
rect 2933 1567 2947 1581
rect 3033 1579 3047 1593
rect 3053 1587 3067 1601
rect 2953 1559 2967 1573
rect 2993 1559 3007 1573
rect 2973 1539 2987 1553
rect 3253 1636 3267 1650
rect 3153 1579 3167 1593
rect 3193 1579 3207 1593
rect 3273 1607 3287 1621
rect 3253 1542 3267 1556
rect 3333 1567 3347 1581
rect 3353 1559 3367 1573
rect 3373 1567 3387 1581
rect 3113 1510 3127 1524
rect 3253 1504 3267 1518
rect 3413 1593 3427 1607
rect 3433 1579 3447 1593
rect 3453 1587 3467 1601
rect 3473 1579 3487 1593
rect 3493 1579 3507 1593
rect 3513 1587 3527 1601
rect 3573 1613 3587 1627
rect 3533 1579 3547 1593
rect 3553 1587 3567 1601
rect 3573 1579 3587 1593
rect 3413 1559 3427 1573
rect 3653 1579 3667 1593
rect 3673 1587 3687 1601
rect 3693 1579 3707 1593
rect 3733 1587 3747 1601
rect 3753 1599 3767 1613
rect 3593 1553 3607 1567
rect 3633 1559 3647 1573
rect 3373 1513 3387 1527
rect 3753 1553 3767 1567
rect 3793 1613 3807 1627
rect 3813 1599 3827 1613
rect 3793 1579 3807 1593
rect 3833 1579 3847 1593
rect 3873 1579 3887 1593
rect 3893 1587 3907 1601
rect 4073 1636 4087 1650
rect 3913 1579 3927 1593
rect 3933 1587 3947 1601
rect 3953 1579 3967 1593
rect 3993 1587 4007 1601
rect 4013 1599 4027 1613
rect 4213 1636 4227 1650
rect 4113 1579 4127 1593
rect 4153 1579 4167 1593
rect 4233 1607 4247 1621
rect 4213 1542 4227 1556
rect 4293 1579 4307 1593
rect 4313 1587 4327 1601
rect 4073 1510 4087 1524
rect 4213 1504 4227 1518
rect 4353 1579 4367 1593
rect 4373 1587 4387 1601
rect 4413 1579 4427 1593
rect 4433 1587 4447 1601
rect 4473 1579 4487 1593
rect 4493 1587 4507 1601
rect 4513 1587 4527 1601
rect 4533 1579 4547 1593
rect 4573 1587 4587 1601
rect 4593 1579 4607 1593
rect 4633 1587 4647 1601
rect 4653 1579 4667 1593
rect 4693 1587 4707 1601
rect 4713 1579 4727 1593
rect 4753 1587 4767 1601
rect 4773 1579 4787 1593
rect 4813 1587 4827 1601
rect 4833 1579 4847 1593
rect 4873 1587 4887 1601
rect 4893 1579 4907 1593
rect 5033 1636 5047 1650
rect 5173 1636 5187 1650
rect 5013 1607 5027 1621
rect 4933 1587 4947 1601
rect 4953 1579 4967 1593
rect 5033 1542 5047 1556
rect 5093 1579 5107 1593
rect 5133 1579 5147 1593
rect 5033 1504 5047 1518
rect 5173 1510 5187 1524
rect 5273 1636 5287 1650
rect 5413 1636 5427 1650
rect 5253 1607 5267 1621
rect 5273 1542 5287 1556
rect 5333 1579 5347 1593
rect 5373 1579 5387 1593
rect 5473 1579 5487 1593
rect 5493 1587 5507 1601
rect 5513 1579 5527 1593
rect 5533 1587 5547 1601
rect 5553 1579 5567 1593
rect 5593 1587 5607 1601
rect 5613 1579 5627 1593
rect 5653 1587 5667 1601
rect 5273 1504 5287 1518
rect 5413 1510 5427 1524
rect 5673 1579 5687 1593
rect 5733 1593 5747 1607
rect 5873 1613 5887 1627
rect 5753 1579 5767 1593
rect 5773 1587 5787 1601
rect 5853 1599 5867 1613
rect 5793 1579 5807 1593
rect 5833 1579 5847 1593
rect 5733 1559 5747 1573
rect 5873 1579 5887 1593
rect 5733 1513 5747 1527
rect 5913 1567 5927 1581
rect 5933 1559 5947 1573
rect 5953 1567 5967 1581
rect 6013 1579 6027 1593
rect 6033 1587 6047 1601
rect 6113 1599 6127 1613
rect 6053 1579 6067 1593
rect 6093 1579 6107 1593
rect 5993 1559 6007 1573
rect 5913 1513 5927 1527
rect 6133 1579 6147 1593
rect 6173 1579 6187 1593
rect 6193 1587 6207 1601
rect 6213 1579 6227 1593
rect 6233 1587 6247 1601
rect 6253 1579 6267 1593
rect 6293 1579 6307 1593
rect 6313 1587 6327 1601
rect 5953 1513 5967 1527
rect 5993 1513 6007 1527
rect 6353 1579 6367 1593
rect 6373 1587 6387 1601
rect 6393 1599 6407 1613
rect 6493 1636 6507 1650
rect 6633 1636 6647 1650
rect 6473 1607 6487 1621
rect 6413 1587 6427 1601
rect 6493 1542 6507 1556
rect 6553 1579 6567 1593
rect 6593 1579 6607 1593
rect 6493 1504 6507 1518
rect 6633 1510 6647 1524
rect 173 1444 187 1447
rect 13 1307 27 1321
rect 173 1433 187 1444
rect 53 1319 67 1333
rect 73 1307 87 1321
rect 113 1307 127 1321
rect 213 1327 227 1341
rect 153 1307 167 1321
rect 233 1307 247 1321
rect 133 1287 147 1301
rect 253 1299 267 1313
rect 273 1307 287 1321
rect 313 1307 327 1321
rect 353 1307 367 1321
rect 713 1376 727 1390
rect 853 1382 867 1396
rect 513 1319 527 1333
rect 533 1327 547 1341
rect 333 1287 347 1301
rect 373 1287 387 1301
rect 393 1299 407 1313
rect 433 1287 447 1301
rect 453 1299 467 1313
rect 553 1319 567 1333
rect 573 1299 587 1313
rect 593 1287 607 1301
rect 613 1299 627 1313
rect 633 1307 647 1321
rect 753 1307 767 1321
rect 793 1307 807 1321
rect 853 1344 867 1358
rect 1013 1347 1027 1361
rect 933 1319 947 1333
rect 953 1327 967 1341
rect 873 1279 887 1293
rect 713 1250 727 1264
rect 973 1319 987 1333
rect 993 1327 1007 1341
rect 1033 1327 1047 1341
rect 1213 1376 1227 1390
rect 1353 1382 1367 1396
rect 1053 1319 1067 1333
rect 1093 1307 1107 1321
rect 1133 1307 1147 1321
rect 853 1250 867 1264
rect 1113 1287 1127 1301
rect 1253 1307 1267 1321
rect 1293 1307 1307 1321
rect 1353 1344 1367 1358
rect 1433 1299 1447 1313
rect 1373 1279 1387 1293
rect 1213 1250 1227 1264
rect 1573 1299 1587 1313
rect 1633 1307 1647 1321
rect 1653 1299 1667 1313
rect 1353 1250 1367 1264
rect 1693 1307 1707 1321
rect 1713 1299 1727 1313
rect 1753 1307 1767 1321
rect 1953 1327 1967 1341
rect 1793 1307 1807 1321
rect 1833 1307 1847 1321
rect 1773 1287 1787 1301
rect 1853 1299 1867 1313
rect 1873 1307 1887 1321
rect 1893 1299 1907 1313
rect 1913 1307 1927 1321
rect 1973 1307 1987 1321
rect 1993 1299 2007 1313
rect 2013 1307 2027 1321
rect 2173 1353 2187 1367
rect 2153 1327 2167 1341
rect 2033 1287 2047 1301
rect 2053 1299 2067 1313
rect 2093 1307 2107 1321
rect 2113 1299 2127 1313
rect 2133 1307 2147 1321
rect 2153 1293 2167 1307
rect 2193 1319 2207 1333
rect 2213 1327 2227 1341
rect 2233 1319 2247 1333
rect 2273 1299 2287 1313
rect 2293 1307 2307 1321
rect 2333 1299 2347 1313
rect 2353 1307 2367 1321
rect 2413 1307 2427 1321
rect 2433 1299 2447 1313
rect 2473 1307 2487 1321
rect 2493 1299 2507 1313
rect 2533 1307 2547 1321
rect 2553 1299 2567 1313
rect 2573 1307 2587 1321
rect 2593 1299 2607 1313
rect 2613 1307 2627 1321
rect 2633 1307 2647 1321
rect 2653 1299 2667 1313
rect 2673 1307 2687 1321
rect 2693 1299 2707 1313
rect 2713 1307 2727 1321
rect 2773 1307 2787 1321
rect 2793 1299 2807 1313
rect 2813 1307 2827 1321
rect 2833 1299 2847 1313
rect 2853 1307 2867 1321
rect 2873 1307 2887 1321
rect 2913 1307 2927 1321
rect 2973 1307 2987 1321
rect 2993 1299 3007 1313
rect 3013 1307 3027 1321
rect 3033 1299 3047 1313
rect 3053 1307 3067 1321
rect 3093 1299 3107 1313
rect 3153 1307 3167 1321
rect 3293 1376 3307 1390
rect 3433 1382 3447 1396
rect 3113 1287 3127 1301
rect 3173 1299 3187 1313
rect 3213 1307 3227 1321
rect 3233 1299 3247 1313
rect 3333 1307 3347 1321
rect 3373 1307 3387 1321
rect 3433 1344 3447 1358
rect 3513 1307 3527 1321
rect 3453 1279 3467 1293
rect 3293 1250 3307 1264
rect 3433 1250 3447 1264
rect 3553 1307 3567 1321
rect 3573 1313 3587 1327
rect 3713 1327 3727 1341
rect 3533 1287 3547 1301
rect 3593 1307 3607 1321
rect 3613 1299 3627 1313
rect 3633 1307 3647 1321
rect 3593 1273 3607 1287
rect 3653 1299 3667 1313
rect 3673 1307 3687 1321
rect 3733 1307 3747 1321
rect 3673 1273 3687 1287
rect 3713 1293 3727 1307
rect 3753 1299 3767 1313
rect 3773 1307 3787 1321
rect 3893 1382 3907 1396
rect 4033 1376 4047 1390
rect 3813 1299 3827 1313
rect 3833 1287 3847 1301
rect 3893 1344 3907 1358
rect 3873 1279 3887 1293
rect 3953 1307 3967 1321
rect 3993 1307 4007 1321
rect 3893 1250 3907 1264
rect 4033 1250 4047 1264
rect 4133 1382 4147 1396
rect 4273 1376 4287 1390
rect 4133 1344 4147 1358
rect 4113 1279 4127 1293
rect 4333 1353 4347 1367
rect 4193 1307 4207 1321
rect 4233 1307 4247 1321
rect 4133 1250 4147 1264
rect 4353 1299 4367 1313
rect 4393 1307 4407 1321
rect 4333 1273 4347 1287
rect 4273 1250 4287 1264
rect 4373 1287 4387 1301
rect 4413 1299 4427 1313
rect 4433 1307 4447 1321
rect 4453 1299 4467 1313
rect 4473 1307 4487 1321
rect 4513 1299 4527 1313
rect 4533 1307 4547 1321
rect 4613 1333 4627 1347
rect 4573 1299 4587 1313
rect 4593 1307 4607 1321
rect 4933 1373 4947 1387
rect 4653 1307 4667 1321
rect 4673 1299 4687 1313
rect 4693 1307 4707 1321
rect 4653 1273 4667 1287
rect 4713 1299 4727 1313
rect 4733 1307 4747 1321
rect 4773 1307 4787 1321
rect 4813 1307 4827 1321
rect 4853 1319 4867 1333
rect 4873 1327 4887 1341
rect 4893 1319 4907 1333
rect 4893 1273 4907 1287
rect 4933 1319 4947 1333
rect 4953 1327 4967 1341
rect 4973 1319 4987 1333
rect 5113 1353 5127 1367
rect 5013 1307 5027 1321
rect 5033 1299 5047 1313
rect 5053 1307 5067 1321
rect 5073 1299 5087 1313
rect 5093 1307 5107 1321
rect 5133 1307 5147 1321
rect 5153 1299 5167 1313
rect 5173 1307 5187 1321
rect 5133 1273 5147 1287
rect 5193 1299 5207 1313
rect 5213 1307 5227 1321
rect 5233 1299 5247 1313
rect 5253 1307 5267 1321
rect 5313 1319 5327 1333
rect 5333 1327 5347 1341
rect 5353 1319 5367 1333
rect 5493 1333 5507 1347
rect 5373 1307 5387 1321
rect 5393 1299 5407 1313
rect 5413 1307 5427 1321
rect 5433 1299 5447 1313
rect 5453 1307 5467 1321
rect 5453 1273 5467 1287
rect 5513 1307 5527 1321
rect 5533 1299 5547 1313
rect 5553 1287 5567 1301
rect 5573 1299 5587 1313
rect 5593 1299 5607 1313
rect 5613 1307 5627 1321
rect 5653 1299 5667 1313
rect 5673 1307 5687 1321
rect 5713 1299 5727 1313
rect 5733 1307 5747 1321
rect 5793 1319 5807 1333
rect 5813 1327 5827 1341
rect 5833 1319 5847 1333
rect 5873 1327 5887 1341
rect 5893 1307 5907 1321
rect 5913 1299 5927 1313
rect 5933 1307 5947 1321
rect 6073 1373 6087 1387
rect 6073 1327 6087 1341
rect 5973 1299 5987 1313
rect 6013 1307 6027 1321
rect 5993 1287 6007 1301
rect 6033 1299 6047 1313
rect 6053 1307 6067 1321
rect 6273 1382 6287 1396
rect 6413 1376 6427 1390
rect 6113 1307 6127 1321
rect 6133 1299 6147 1313
rect 6153 1307 6167 1321
rect 6113 1273 6127 1287
rect 6173 1299 6187 1313
rect 6193 1307 6207 1321
rect 6273 1344 6287 1358
rect 6253 1279 6267 1293
rect 6333 1307 6347 1321
rect 6373 1307 6387 1321
rect 6273 1250 6287 1264
rect 6413 1250 6427 1264
rect 6513 1382 6527 1396
rect 6653 1376 6667 1390
rect 6513 1344 6527 1358
rect 6493 1279 6507 1293
rect 6573 1307 6587 1321
rect 6613 1307 6627 1321
rect 6513 1250 6527 1264
rect 6653 1250 6667 1264
rect 53 1156 67 1170
rect 193 1156 207 1170
rect 33 1127 47 1141
rect 53 1062 67 1076
rect 113 1099 127 1113
rect 153 1099 167 1113
rect 353 1156 367 1170
rect 493 1156 507 1170
rect 273 1107 287 1121
rect 293 1119 307 1133
rect 333 1127 347 1141
rect 53 1024 67 1038
rect 193 1030 207 1044
rect 353 1062 367 1076
rect 413 1099 427 1113
rect 453 1099 467 1113
rect 553 1119 567 1133
rect 573 1107 587 1121
rect 353 1024 367 1038
rect 493 1030 507 1044
rect 633 1113 647 1127
rect 733 1119 747 1133
rect 613 1079 627 1093
rect 653 1079 667 1093
rect 673 1087 687 1101
rect 713 1099 727 1113
rect 633 1059 647 1073
rect 613 1033 627 1047
rect 773 1113 787 1127
rect 813 1113 827 1127
rect 753 1099 767 1113
rect 793 1079 807 1093
rect 833 1079 847 1093
rect 853 1087 867 1101
rect 893 1087 907 1101
rect 973 1119 987 1133
rect 1073 1156 1087 1170
rect 993 1107 1007 1121
rect 813 1059 827 1073
rect 913 1079 927 1093
rect 933 1087 947 1101
rect 1213 1156 1227 1170
rect 1513 1156 1527 1170
rect 1113 1099 1127 1113
rect 1153 1099 1167 1113
rect 1233 1127 1247 1141
rect 1213 1062 1227 1076
rect 1293 1107 1307 1121
rect 1433 1107 1447 1121
rect 1653 1156 1667 1170
rect 1553 1099 1567 1113
rect 1593 1099 1607 1113
rect 1073 1030 1087 1044
rect 1213 1024 1227 1038
rect 1673 1127 1687 1141
rect 1653 1062 1667 1076
rect 1753 1119 1767 1133
rect 1733 1099 1747 1113
rect 1773 1099 1787 1113
rect 1813 1099 1827 1113
rect 1833 1107 1847 1121
rect 1853 1099 1867 1113
rect 1873 1107 1887 1121
rect 1993 1133 2007 1147
rect 1893 1099 1907 1113
rect 1953 1099 1967 1113
rect 1973 1107 1987 1121
rect 1993 1099 2007 1113
rect 1513 1030 1527 1044
rect 1653 1024 1667 1038
rect 1933 1079 1947 1093
rect 2353 1156 2367 1170
rect 2053 1099 2067 1113
rect 2073 1107 2087 1121
rect 2153 1119 2167 1133
rect 2093 1099 2107 1113
rect 2133 1099 2147 1113
rect 2033 1079 2047 1093
rect 2173 1099 2187 1113
rect 2213 1099 2227 1113
rect 2233 1107 2247 1121
rect 2253 1099 2267 1113
rect 2273 1107 2287 1121
rect 2293 1099 2307 1113
rect 2493 1156 2507 1170
rect 2393 1099 2407 1113
rect 2433 1099 2447 1113
rect 2033 1033 2047 1047
rect 2513 1127 2527 1141
rect 2493 1062 2507 1076
rect 2573 1107 2587 1121
rect 2593 1119 2607 1133
rect 2353 1030 2367 1044
rect 2493 1024 2507 1038
rect 2613 1099 2627 1113
rect 2633 1107 2647 1121
rect 2653 1099 2667 1113
rect 2733 1099 2747 1113
rect 2673 1079 2687 1093
rect 2793 1119 2807 1133
rect 3013 1156 3027 1170
rect 2773 1099 2787 1113
rect 2813 1107 2827 1121
rect 2873 1099 2887 1113
rect 2893 1107 2907 1121
rect 2913 1099 2927 1113
rect 2933 1107 2947 1121
rect 2953 1099 2967 1113
rect 3153 1156 3167 1170
rect 3053 1099 3067 1113
rect 3093 1099 3107 1113
rect 3173 1127 3187 1141
rect 3153 1062 3167 1076
rect 3213 1087 3227 1101
rect 3233 1079 3247 1093
rect 3253 1087 3267 1101
rect 3313 1099 3327 1113
rect 3333 1107 3347 1121
rect 3013 1030 3027 1044
rect 3153 1024 3167 1038
rect 3373 1099 3387 1113
rect 3393 1107 3407 1121
rect 3413 1107 3427 1121
rect 3433 1099 3447 1113
rect 3473 1107 3487 1121
rect 3653 1156 3667 1170
rect 3493 1099 3507 1113
rect 3553 1099 3567 1113
rect 3593 1099 3607 1113
rect 3793 1156 3807 1170
rect 3693 1099 3707 1113
rect 3733 1099 3747 1113
rect 3813 1127 3827 1141
rect 3793 1062 3807 1076
rect 3853 1107 3867 1121
rect 3873 1099 3887 1113
rect 3913 1107 3927 1121
rect 3653 1030 3667 1044
rect 3793 1024 3807 1038
rect 3933 1099 3947 1113
rect 3993 1099 4007 1113
rect 4013 1107 4027 1121
rect 4053 1099 4067 1113
rect 4073 1107 4087 1121
rect 4093 1119 4107 1133
rect 4113 1107 4127 1121
rect 4153 1133 4167 1147
rect 4153 1099 4167 1113
rect 4173 1107 4187 1121
rect 4593 1156 4607 1170
rect 4193 1099 4207 1113
rect 4213 1107 4227 1121
rect 4293 1119 4307 1133
rect 4233 1099 4247 1113
rect 4273 1099 4287 1113
rect 4133 1053 4147 1067
rect 4313 1099 4327 1113
rect 4393 1099 4407 1113
rect 4413 1107 4427 1121
rect 4433 1099 4447 1113
rect 4473 1099 4487 1113
rect 4493 1107 4507 1121
rect 4513 1119 4527 1133
rect 4533 1107 4547 1121
rect 4373 1079 4387 1093
rect 4733 1156 4747 1170
rect 4633 1099 4647 1113
rect 4673 1099 4687 1113
rect 4753 1127 4767 1141
rect 4733 1062 4747 1076
rect 4793 1099 4807 1113
rect 4813 1107 4827 1121
rect 4833 1099 4847 1113
rect 4853 1107 4867 1121
rect 4953 1119 4967 1133
rect 4873 1099 4887 1113
rect 4933 1099 4947 1113
rect 5093 1133 5107 1147
rect 4973 1099 4987 1113
rect 5033 1099 5047 1113
rect 5053 1107 5067 1121
rect 5073 1099 5087 1113
rect 5013 1079 5027 1093
rect 5133 1119 5147 1133
rect 5193 1119 5207 1133
rect 5273 1119 5287 1133
rect 5113 1099 5127 1113
rect 5153 1099 5167 1113
rect 5173 1099 5187 1113
rect 4593 1030 4607 1044
rect 4733 1024 4747 1038
rect 5093 1053 5107 1067
rect 5213 1099 5227 1113
rect 5253 1099 5267 1113
rect 5293 1099 5307 1113
rect 5353 1099 5367 1113
rect 5533 1133 5547 1147
rect 5433 1119 5447 1133
rect 5513 1119 5527 1133
rect 5393 1099 5407 1113
rect 5413 1099 5427 1113
rect 5453 1099 5467 1113
rect 5493 1099 5507 1113
rect 5533 1099 5547 1113
rect 5573 1107 5587 1121
rect 5593 1119 5607 1133
rect 5613 1107 5627 1121
rect 5673 1119 5687 1133
rect 5633 1099 5647 1113
rect 5693 1099 5707 1113
rect 5573 1073 5587 1087
rect 5733 1107 5747 1121
rect 5813 1119 5827 1133
rect 5793 1099 5807 1113
rect 5833 1099 5847 1113
rect 5853 1099 5867 1113
rect 5873 1107 5887 1121
rect 5913 1113 5927 1127
rect 5893 1099 5907 1113
rect 5913 1079 5927 1093
rect 5973 1087 5987 1101
rect 6053 1099 6067 1113
rect 6073 1107 6087 1121
rect 6113 1113 6127 1127
rect 6093 1099 6107 1113
rect 5933 1053 5947 1067
rect 5993 1079 6007 1093
rect 6033 1079 6047 1093
rect 6013 1059 6027 1073
rect 6113 1079 6127 1093
rect 6113 1033 6127 1047
rect 6193 1119 6207 1133
rect 6253 1119 6267 1133
rect 6173 1099 6187 1113
rect 6213 1099 6227 1113
rect 6233 1099 6247 1113
rect 6353 1156 6367 1170
rect 6493 1156 6507 1170
rect 6333 1127 6347 1141
rect 6273 1099 6287 1113
rect 6353 1062 6367 1076
rect 6413 1099 6427 1113
rect 6453 1099 6467 1113
rect 6553 1099 6567 1113
rect 6573 1107 6587 1121
rect 6593 1099 6607 1113
rect 6613 1107 6627 1121
rect 6633 1099 6647 1113
rect 6353 1024 6367 1038
rect 6493 1030 6507 1044
rect 33 827 47 841
rect 13 807 27 821
rect 233 902 247 916
rect 373 896 387 910
rect 133 839 147 853
rect 153 847 167 861
rect 73 819 87 833
rect 173 839 187 853
rect 233 864 247 878
rect 213 799 227 813
rect 293 827 307 841
rect 333 827 347 841
rect 233 770 247 784
rect 493 833 507 847
rect 453 819 467 833
rect 373 770 387 784
rect 473 807 487 821
rect 473 773 487 787
rect 513 827 527 841
rect 553 827 567 841
rect 573 827 587 841
rect 693 873 707 887
rect 613 827 627 841
rect 653 839 667 853
rect 673 847 687 861
rect 533 807 547 821
rect 593 807 607 821
rect 693 839 707 853
rect 753 867 767 881
rect 733 847 747 861
rect 773 847 787 861
rect 793 839 807 853
rect 933 873 947 887
rect 733 813 747 827
rect 833 827 847 841
rect 853 819 867 833
rect 873 827 887 841
rect 893 819 907 833
rect 913 827 927 841
rect 1013 847 1027 861
rect 1113 847 1127 861
rect 953 827 967 841
rect 973 819 987 833
rect 993 827 1007 841
rect 1053 827 1067 841
rect 953 793 967 807
rect 1013 813 1027 827
rect 1073 819 1087 833
rect 1093 827 1107 841
rect 1393 847 1407 861
rect 1053 793 1067 807
rect 1113 813 1127 827
rect 1153 813 1167 827
rect 1193 819 1207 833
rect 1233 827 1247 841
rect 1253 819 1267 833
rect 1293 827 1307 841
rect 1333 827 1347 841
rect 1353 819 1367 833
rect 1373 827 1387 841
rect 1533 896 1547 910
rect 1673 902 1687 916
rect 1453 819 1467 833
rect 1473 807 1487 821
rect 1573 827 1587 841
rect 1613 827 1627 841
rect 1673 864 1687 878
rect 1693 799 1707 813
rect 1733 807 1747 821
rect 1753 819 1767 833
rect 1793 819 1807 833
rect 1813 827 1827 841
rect 1533 770 1547 784
rect 1673 770 1687 784
rect 2133 902 2147 916
rect 2273 896 2287 910
rect 1973 847 1987 861
rect 1853 819 1867 833
rect 1873 827 1887 841
rect 1913 827 1927 841
rect 1933 819 1947 833
rect 1953 827 1967 841
rect 2013 839 2027 853
rect 2033 847 2047 861
rect 2053 839 2067 853
rect 2133 864 2147 878
rect 2113 799 2127 813
rect 2193 827 2207 841
rect 2233 827 2247 841
rect 2133 770 2147 784
rect 2373 853 2387 867
rect 2333 807 2347 821
rect 2353 819 2367 833
rect 2273 770 2287 784
rect 2393 827 2407 841
rect 2413 819 2427 833
rect 2433 827 2447 841
rect 2393 793 2407 807
rect 2453 819 2467 833
rect 2473 827 2487 841
rect 2513 827 2527 841
rect 2613 847 2627 861
rect 2553 827 2567 841
rect 2633 827 2647 841
rect 2533 807 2547 821
rect 2653 819 2667 833
rect 2673 827 2687 841
rect 2713 819 2727 833
rect 2873 853 2887 867
rect 2933 853 2947 867
rect 2853 819 2867 833
rect 2893 819 2907 833
rect 2913 807 2927 821
rect 2933 819 2947 833
rect 2953 827 2967 841
rect 3013 827 3027 841
rect 3033 819 3047 833
rect 3053 807 3067 821
rect 3073 819 3087 833
rect 3113 827 3127 841
rect 3133 819 3147 833
rect 3173 827 3187 841
rect 3193 819 3207 833
rect 3233 827 3247 841
rect 3253 819 3267 833
rect 3353 847 3367 861
rect 3293 827 3307 841
rect 3313 819 3327 833
rect 3373 827 3387 841
rect 3393 819 3407 833
rect 3413 827 3427 841
rect 3433 839 3447 853
rect 3453 847 3467 861
rect 3473 839 3487 853
rect 3513 819 3527 833
rect 3533 827 3547 841
rect 3573 819 3587 833
rect 3593 827 3607 841
rect 3653 819 3667 833
rect 3713 827 3727 841
rect 3853 896 3867 910
rect 3993 902 4007 916
rect 3673 807 3687 821
rect 3733 819 3747 833
rect 3773 827 3787 841
rect 3793 819 3807 833
rect 3893 827 3907 841
rect 3933 827 3947 841
rect 3993 864 4007 878
rect 4053 819 4067 833
rect 4073 827 4087 841
rect 4013 799 4027 813
rect 4153 853 4167 867
rect 4213 853 4227 867
rect 4253 853 4267 867
rect 4113 819 4127 833
rect 4133 827 4147 841
rect 4173 819 4187 833
rect 3853 770 3867 784
rect 3993 770 4007 784
rect 4193 807 4207 821
rect 4213 819 4227 833
rect 4233 827 4247 841
rect 4333 847 4347 861
rect 4433 867 4447 881
rect 4273 827 4287 841
rect 4293 819 4307 833
rect 4313 827 4327 841
rect 4393 839 4407 853
rect 4413 847 4427 861
rect 4453 847 4467 861
rect 4273 793 4287 807
rect 4613 873 4627 887
rect 4593 847 4607 861
rect 4473 807 4487 821
rect 4493 819 4507 833
rect 4533 827 4547 841
rect 4553 819 4567 833
rect 4573 827 4587 841
rect 4593 813 4607 827
rect 4633 839 4647 853
rect 4653 847 4667 861
rect 4673 839 4687 853
rect 4833 847 4847 861
rect 4733 819 4747 833
rect 4773 827 4787 841
rect 4753 807 4767 821
rect 4793 819 4807 833
rect 4813 827 4827 841
rect 4833 813 4847 827
rect 4873 873 4887 887
rect 4873 839 4887 853
rect 4893 847 4907 861
rect 4913 839 4927 853
rect 4953 819 4967 833
rect 4973 827 4987 841
rect 5013 819 5027 833
rect 5033 827 5047 841
rect 5093 827 5107 841
rect 5113 819 5127 833
rect 5153 827 5167 841
rect 5173 819 5187 833
rect 5213 819 5227 833
rect 5353 819 5367 833
rect 5393 819 5407 833
rect 5413 807 5427 821
rect 5433 819 5447 833
rect 5453 827 5467 841
rect 5613 847 5627 861
rect 5513 819 5527 833
rect 5553 827 5567 841
rect 5533 807 5547 821
rect 5573 819 5587 833
rect 5593 827 5607 841
rect 5653 839 5667 853
rect 5673 847 5687 861
rect 5693 839 5707 853
rect 5793 847 5807 861
rect 5893 867 5907 881
rect 5973 896 5987 910
rect 6113 902 6127 916
rect 5733 827 5747 841
rect 5753 819 5767 833
rect 5773 827 5787 841
rect 5853 839 5867 853
rect 5873 847 5887 861
rect 5913 847 5927 861
rect 6013 827 6027 841
rect 6053 827 6067 841
rect 6113 864 6127 878
rect 6233 847 6247 861
rect 6493 896 6507 910
rect 6633 902 6647 916
rect 6333 847 6347 861
rect 6173 827 6187 841
rect 6193 819 6207 833
rect 6213 827 6227 841
rect 6273 827 6287 841
rect 6133 799 6147 813
rect 6293 819 6307 833
rect 6313 827 6327 841
rect 6393 839 6407 853
rect 6413 847 6427 861
rect 5973 770 5987 784
rect 6433 839 6447 853
rect 6113 770 6127 784
rect 6533 827 6547 841
rect 6573 827 6587 841
rect 6633 864 6647 878
rect 6653 799 6667 813
rect 6493 770 6507 784
rect 6633 770 6647 784
rect 13 639 27 653
rect 33 627 47 641
rect 73 607 87 621
rect 153 627 167 641
rect 173 639 187 653
rect 193 627 207 641
rect 253 639 267 653
rect 93 599 107 613
rect 113 607 127 621
rect 213 619 227 633
rect 273 627 287 641
rect 333 619 347 633
rect 353 627 367 641
rect 373 639 387 653
rect 393 627 407 641
rect 413 599 427 613
rect 453 599 467 613
rect 473 607 487 621
rect 533 607 547 621
rect 693 639 707 653
rect 713 627 727 641
rect 753 639 767 653
rect 773 627 787 641
rect 853 639 867 653
rect 1113 676 1127 690
rect 433 579 447 593
rect 553 599 567 613
rect 573 607 587 621
rect 613 607 627 621
rect 633 599 647 613
rect 673 599 687 613
rect 653 579 667 593
rect 833 619 847 633
rect 873 619 887 633
rect 933 627 947 641
rect 973 619 987 633
rect 993 627 1007 641
rect 1033 619 1047 633
rect 1253 676 1267 690
rect 1153 619 1167 633
rect 1193 619 1207 633
rect 1273 647 1287 661
rect 1253 582 1267 596
rect 1313 619 1327 633
rect 1513 676 1527 690
rect 1353 619 1367 633
rect 1113 550 1127 564
rect 1253 544 1267 558
rect 1393 607 1407 621
rect 1413 599 1427 613
rect 1433 607 1447 621
rect 1653 676 1667 690
rect 1553 619 1567 633
rect 1593 619 1607 633
rect 1673 647 1687 661
rect 1653 582 1667 596
rect 1513 550 1527 564
rect 1653 544 1667 558
rect 1753 676 1767 690
rect 1893 676 1907 690
rect 1793 619 1807 633
rect 1833 619 1847 633
rect 1913 647 1927 661
rect 1893 582 1907 596
rect 1753 550 1767 564
rect 1893 544 1907 558
rect 1993 676 2007 690
rect 2133 676 2147 690
rect 2033 619 2047 633
rect 2073 619 2087 633
rect 2153 647 2167 661
rect 2133 582 2147 596
rect 1993 550 2007 564
rect 2133 544 2147 558
rect 2233 676 2247 690
rect 2373 676 2387 690
rect 2273 619 2287 633
rect 2313 619 2327 633
rect 2393 647 2407 661
rect 2373 582 2387 596
rect 2233 550 2247 564
rect 2373 544 2387 558
rect 2473 676 2487 690
rect 2613 676 2627 690
rect 2453 647 2467 661
rect 2473 582 2487 596
rect 2533 619 2547 633
rect 2573 619 2587 633
rect 2693 619 2707 633
rect 2713 627 2727 641
rect 2733 619 2747 633
rect 2753 627 2767 641
rect 2773 619 2787 633
rect 2813 627 2827 641
rect 2833 639 2847 653
rect 2473 544 2487 558
rect 2613 550 2627 564
rect 2873 619 2887 633
rect 2893 627 2907 641
rect 2913 639 2927 653
rect 2933 627 2947 641
rect 2953 639 2967 653
rect 2993 673 3007 687
rect 2973 627 2987 641
rect 3013 619 3027 633
rect 3033 627 3047 641
rect 3073 633 3087 647
rect 3113 653 3127 667
rect 3053 619 3067 633
rect 2993 573 3007 587
rect 3073 599 3087 613
rect 3113 607 3127 621
rect 3133 599 3147 613
rect 3153 607 3167 621
rect 3193 633 3207 647
rect 3293 639 3307 653
rect 3313 627 3327 641
rect 3193 599 3207 613
rect 3233 599 3247 613
rect 3253 607 3267 621
rect 3173 573 3187 587
rect 3213 579 3227 593
rect 3353 619 3367 633
rect 3373 627 3387 641
rect 3393 619 3407 633
rect 3413 599 3427 613
rect 3453 607 3467 621
rect 3533 627 3547 641
rect 3553 639 3567 653
rect 3573 627 3587 641
rect 3813 693 3827 707
rect 3653 639 3667 653
rect 3473 599 3487 613
rect 3493 607 3507 621
rect 3593 619 3607 633
rect 3633 619 3647 633
rect 3673 619 3687 633
rect 3713 619 3727 633
rect 3733 627 3747 641
rect 3773 633 3787 647
rect 3953 676 3967 690
rect 4093 676 4107 690
rect 3753 619 3767 633
rect 3933 647 3947 661
rect 3773 599 3787 613
rect 3833 607 3847 621
rect 3853 599 3867 613
rect 3893 599 3907 613
rect 3873 579 3887 593
rect 3953 582 3967 596
rect 4013 619 4027 633
rect 4053 619 4067 633
rect 4273 676 4287 690
rect 4413 676 4427 690
rect 4193 639 4207 653
rect 4253 647 4267 661
rect 4173 619 4187 633
rect 4213 619 4227 633
rect 3953 544 3967 558
rect 4093 550 4107 564
rect 4273 582 4287 596
rect 4333 619 4347 633
rect 4373 619 4387 633
rect 4473 639 4487 653
rect 4493 627 4507 641
rect 4273 544 4287 558
rect 4413 550 4427 564
rect 4533 619 4547 633
rect 4553 627 4567 641
rect 4573 619 4587 633
rect 4593 627 4607 641
rect 4613 619 4627 633
rect 4673 619 4687 633
rect 4693 627 4707 641
rect 4713 639 4727 653
rect 4733 627 4747 641
rect 4773 633 4787 647
rect 4793 619 4807 633
rect 4813 627 4827 641
rect 4833 619 4847 633
rect 4773 599 4787 613
rect 4753 573 4767 587
rect 4853 607 4867 621
rect 4953 627 4967 641
rect 4973 639 4987 653
rect 4873 599 4887 613
rect 4893 607 4907 621
rect 5013 619 5027 633
rect 5033 627 5047 641
rect 5253 676 5267 690
rect 5393 676 5407 690
rect 5073 619 5087 633
rect 5093 627 5107 641
rect 5233 647 5247 661
rect 5113 599 5127 613
rect 5153 599 5167 613
rect 5173 607 5187 621
rect 5133 579 5147 593
rect 5253 582 5267 596
rect 5313 619 5327 633
rect 5353 619 5367 633
rect 5453 627 5467 641
rect 5473 619 5487 633
rect 5513 627 5527 641
rect 5533 619 5547 633
rect 5693 653 5707 667
rect 5573 627 5587 641
rect 5673 639 5687 653
rect 5253 544 5267 558
rect 5393 550 5407 564
rect 5593 619 5607 633
rect 5653 619 5667 633
rect 5693 619 5707 633
rect 5913 653 5927 667
rect 5753 639 5767 653
rect 5833 639 5847 653
rect 5893 639 5907 653
rect 5733 619 5747 633
rect 5713 593 5727 607
rect 5773 619 5787 633
rect 5813 619 5827 633
rect 5853 619 5867 633
rect 5873 619 5887 633
rect 5913 619 5927 633
rect 6353 676 6367 690
rect 5993 639 6007 653
rect 5973 619 5987 633
rect 5953 593 5967 607
rect 6013 619 6027 633
rect 6033 619 6047 633
rect 6053 627 6067 641
rect 6073 619 6087 633
rect 6133 619 6147 633
rect 6153 627 6167 641
rect 6173 619 6187 633
rect 6093 599 6107 613
rect 6193 599 6207 613
rect 6253 607 6267 621
rect 6273 599 6287 613
rect 6293 607 6307 621
rect 6493 676 6507 690
rect 6393 619 6407 633
rect 6433 619 6447 633
rect 6513 647 6527 661
rect 6493 582 6507 596
rect 6553 639 6567 653
rect 6573 627 6587 641
rect 6613 639 6627 653
rect 6633 627 6647 641
rect 6353 550 6367 564
rect 6493 544 6507 558
rect 53 422 67 436
rect 193 416 207 430
rect 53 384 67 398
rect 33 319 47 333
rect 113 347 127 361
rect 153 347 167 361
rect 53 290 67 304
rect 193 290 207 304
rect 293 416 307 430
rect 433 422 447 436
rect 333 347 347 361
rect 373 347 387 361
rect 433 384 447 398
rect 513 387 527 401
rect 493 367 507 381
rect 533 367 547 381
rect 573 393 587 407
rect 553 359 567 373
rect 453 319 467 333
rect 293 290 307 304
rect 433 290 447 304
rect 593 347 607 361
rect 633 347 647 361
rect 693 347 707 361
rect 613 327 627 341
rect 593 313 607 327
rect 733 347 747 361
rect 753 359 767 373
rect 773 367 787 381
rect 713 327 727 341
rect 793 359 807 373
rect 933 416 947 430
rect 1073 422 1087 436
rect 853 339 867 353
rect 873 327 887 341
rect 973 347 987 361
rect 1013 347 1027 361
rect 1073 384 1087 398
rect 1093 319 1107 333
rect 933 290 947 304
rect 1153 347 1167 361
rect 1193 347 1207 361
rect 1213 347 1227 361
rect 1253 347 1267 361
rect 1293 347 1307 361
rect 1073 290 1087 304
rect 1333 347 1347 361
rect 1493 367 1507 381
rect 1393 339 1407 353
rect 1433 347 1447 361
rect 1413 327 1427 341
rect 1453 339 1467 353
rect 1473 347 1487 361
rect 1733 416 1747 430
rect 1873 422 1887 436
rect 1653 367 1667 381
rect 1553 339 1567 353
rect 1593 347 1607 361
rect 1573 327 1587 341
rect 1613 339 1627 353
rect 1633 347 1647 361
rect 1773 347 1787 361
rect 1813 347 1827 361
rect 1873 384 1887 398
rect 2113 367 2127 381
rect 1953 339 1967 353
rect 1893 319 1907 333
rect 1733 290 1747 304
rect 1873 290 1887 304
rect 1973 327 1987 341
rect 2013 339 2027 353
rect 2053 347 2067 361
rect 2033 327 2047 341
rect 2073 339 2087 353
rect 2093 347 2107 361
rect 2193 373 2207 387
rect 2153 327 2167 341
rect 2173 339 2187 353
rect 2353 367 2367 381
rect 2213 347 2227 361
rect 2233 339 2247 353
rect 2253 347 2267 361
rect 2273 339 2287 353
rect 2293 347 2307 361
rect 2333 353 2347 367
rect 2553 416 2567 430
rect 2693 422 2707 436
rect 2193 293 2207 307
rect 2293 313 2307 327
rect 2373 347 2387 361
rect 2393 339 2407 353
rect 2413 347 2427 361
rect 2433 347 2447 361
rect 2473 347 2487 361
rect 2453 327 2467 341
rect 2593 347 2607 361
rect 2633 347 2647 361
rect 2693 384 2707 398
rect 2773 367 2787 381
rect 2973 416 2987 430
rect 3113 422 3127 436
rect 2713 319 2727 333
rect 2793 347 2807 361
rect 2813 339 2827 353
rect 2833 347 2847 361
rect 2853 347 2867 361
rect 2893 347 2907 361
rect 2873 327 2887 341
rect 2553 290 2567 304
rect 2693 290 2707 304
rect 3013 347 3027 361
rect 3053 347 3067 361
rect 3113 384 3127 398
rect 3173 359 3187 373
rect 3193 367 3207 381
rect 3133 319 3147 333
rect 2973 290 2987 304
rect 3213 359 3227 373
rect 3273 367 3287 381
rect 3293 347 3307 361
rect 3313 339 3327 353
rect 3333 347 3347 361
rect 3353 347 3367 361
rect 3593 367 3607 381
rect 3393 347 3407 361
rect 3453 347 3467 361
rect 3373 327 3387 341
rect 3113 290 3127 304
rect 3473 339 3487 353
rect 3493 327 3507 341
rect 3513 339 3527 353
rect 3533 347 3547 361
rect 3553 339 3567 353
rect 3573 347 3587 361
rect 3633 347 3647 361
rect 3673 347 3687 361
rect 3653 327 3667 341
rect 3673 313 3687 327
rect 3713 373 3727 387
rect 3713 339 3727 353
rect 3733 327 3747 341
rect 3753 339 3767 353
rect 3773 347 3787 361
rect 3833 347 3847 361
rect 3953 367 3967 381
rect 4053 387 4067 401
rect 4153 393 4167 407
rect 4213 422 4227 436
rect 4353 416 4367 430
rect 3873 347 3887 361
rect 3893 347 3907 361
rect 3853 327 3867 341
rect 3913 339 3927 353
rect 3933 347 3947 361
rect 4013 359 4027 373
rect 4033 367 4047 381
rect 4073 367 4087 381
rect 4093 347 4107 361
rect 4133 347 4147 361
rect 4113 327 4127 341
rect 4133 313 4147 327
rect 4213 384 4227 398
rect 4193 319 4207 333
rect 4273 347 4287 361
rect 4313 347 4327 361
rect 4213 290 4227 304
rect 4413 347 4427 361
rect 4513 367 4527 381
rect 4453 347 4467 361
rect 4533 347 4547 361
rect 4433 327 4447 341
rect 4353 290 4367 304
rect 4553 339 4567 353
rect 4573 347 4587 361
rect 4593 347 4607 361
rect 4633 347 4647 361
rect 4693 347 4707 361
rect 4613 327 4627 341
rect 4713 339 4727 353
rect 4733 347 4747 361
rect 4753 339 4767 353
rect 4773 347 4787 361
rect 4893 416 4907 430
rect 5033 422 5047 436
rect 4813 339 4827 353
rect 4833 327 4847 341
rect 4933 347 4947 361
rect 4973 347 4987 361
rect 5033 384 5047 398
rect 5113 347 5127 361
rect 5053 319 5067 333
rect 4893 290 4907 304
rect 5033 290 5047 304
rect 5133 339 5147 353
rect 5153 327 5167 341
rect 5173 339 5187 353
rect 5193 347 5207 361
rect 5253 373 5267 387
rect 5233 347 5247 361
rect 5213 327 5227 341
rect 5233 313 5247 327
rect 5293 367 5307 381
rect 5313 347 5327 361
rect 5333 339 5347 353
rect 5353 347 5367 361
rect 5373 347 5387 361
rect 5573 387 5587 401
rect 5553 367 5567 381
rect 5593 367 5607 381
rect 5413 347 5427 361
rect 5393 327 5407 341
rect 5453 339 5467 353
rect 5473 327 5487 341
rect 5493 339 5507 353
rect 5513 347 5527 361
rect 5613 359 5627 373
rect 5713 367 5727 381
rect 5653 347 5667 361
rect 5673 339 5687 353
rect 5693 347 5707 361
rect 5773 359 5787 373
rect 5793 367 5807 381
rect 5813 359 5827 373
rect 5853 367 5867 381
rect 5993 367 6007 381
rect 6133 393 6147 407
rect 6093 367 6107 381
rect 5873 347 5887 361
rect 5893 339 5907 353
rect 5913 347 5927 361
rect 5933 347 5947 361
rect 5953 339 5967 353
rect 5973 347 5987 361
rect 6033 347 6047 361
rect 6053 339 6067 353
rect 6073 347 6087 361
rect 6293 393 6307 407
rect 6453 416 6467 430
rect 6593 422 6607 436
rect 6153 347 6167 361
rect 6193 347 6207 361
rect 6233 347 6247 361
rect 6273 347 6287 361
rect 6173 327 6187 341
rect 6253 327 6267 341
rect 6313 347 6327 361
rect 6333 339 6347 353
rect 6353 347 6367 361
rect 6153 313 6167 327
rect 6293 313 6307 327
rect 6373 339 6387 353
rect 6393 347 6407 361
rect 6493 347 6507 361
rect 6533 347 6547 361
rect 6593 384 6607 398
rect 6613 319 6627 333
rect 6453 290 6467 304
rect 6593 290 6607 304
rect 53 196 67 210
rect 193 196 207 210
rect 33 167 47 181
rect 53 102 67 116
rect 113 139 127 153
rect 153 139 167 153
rect 53 64 67 78
rect 193 70 207 84
rect 293 196 307 210
rect 433 196 447 210
rect 273 167 287 181
rect 293 102 307 116
rect 353 139 367 153
rect 393 139 407 153
rect 513 139 527 153
rect 553 139 567 153
rect 573 139 587 153
rect 613 139 627 153
rect 293 64 307 78
rect 433 70 447 84
rect 773 196 787 210
rect 673 139 687 153
rect 913 196 927 210
rect 753 167 767 181
rect 713 139 727 153
rect 773 102 787 116
rect 833 139 847 153
rect 873 139 887 153
rect 973 139 987 153
rect 1013 139 1027 153
rect 773 64 787 78
rect 913 70 927 84
rect 1073 127 1087 141
rect 1273 196 1287 210
rect 1093 119 1107 133
rect 1113 127 1127 141
rect 1173 139 1187 153
rect 1193 147 1207 161
rect 1213 139 1227 153
rect 1153 119 1167 133
rect 1413 196 1427 210
rect 1313 139 1327 153
rect 1353 139 1367 153
rect 1433 167 1447 181
rect 1413 102 1427 116
rect 1493 147 1507 161
rect 1513 159 1527 173
rect 1273 70 1287 84
rect 1413 64 1427 78
rect 1533 127 1547 141
rect 1553 119 1567 133
rect 1573 127 1587 141
rect 1653 139 1667 153
rect 1673 147 1687 161
rect 1713 159 1727 173
rect 2153 196 2167 210
rect 1693 139 1707 153
rect 1733 147 1747 161
rect 1633 119 1647 133
rect 1773 127 1787 141
rect 1793 119 1807 133
rect 1813 127 1827 141
rect 1853 127 1867 141
rect 1873 119 1887 133
rect 1893 127 1907 141
rect 1933 127 1947 141
rect 1953 119 1967 133
rect 1973 127 1987 141
rect 2053 139 2067 153
rect 2073 147 2087 161
rect 2093 139 2107 153
rect 2033 119 2047 133
rect 2293 196 2307 210
rect 2193 139 2207 153
rect 2233 139 2247 153
rect 2313 167 2327 181
rect 2293 102 2307 116
rect 2353 127 2367 141
rect 2373 119 2387 133
rect 2393 127 2407 141
rect 2453 127 2467 141
rect 2713 196 2727 210
rect 2473 119 2487 133
rect 2493 127 2507 141
rect 2553 139 2567 153
rect 2573 147 2587 161
rect 2593 139 2607 153
rect 2633 147 2647 161
rect 2653 159 2667 173
rect 2533 119 2547 133
rect 2153 70 2167 84
rect 2293 64 2307 78
rect 2853 196 2867 210
rect 2753 139 2767 153
rect 2793 139 2807 153
rect 2873 167 2887 181
rect 2853 102 2867 116
rect 2953 139 2967 153
rect 2973 147 2987 161
rect 3053 159 3067 173
rect 2993 139 3007 153
rect 3033 139 3047 153
rect 2933 119 2947 133
rect 3073 139 3087 153
rect 3113 139 3127 153
rect 3133 147 3147 161
rect 3313 196 3327 210
rect 3453 196 3467 210
rect 3153 139 3167 153
rect 3173 147 3187 161
rect 3193 139 3207 153
rect 3233 147 3247 161
rect 3253 159 3267 173
rect 3293 167 3307 181
rect 2713 70 2727 84
rect 2853 64 2867 78
rect 3313 102 3327 116
rect 3373 139 3387 153
rect 3413 139 3427 153
rect 3533 127 3547 141
rect 3833 196 3847 210
rect 3973 196 3987 210
rect 3553 119 3567 133
rect 3573 127 3587 141
rect 3633 139 3647 153
rect 3653 147 3667 161
rect 3673 139 3687 153
rect 3693 139 3707 153
rect 3713 147 3727 161
rect 3733 139 3747 153
rect 3813 167 3827 181
rect 3613 119 3627 133
rect 3313 64 3327 78
rect 3453 70 3467 84
rect 3753 119 3767 133
rect 3833 102 3847 116
rect 3893 139 3907 153
rect 3933 139 3947 153
rect 4353 196 4367 210
rect 4033 139 4047 153
rect 4053 147 4067 161
rect 4073 139 4087 153
rect 4133 139 4147 153
rect 4153 147 4167 161
rect 4173 139 4187 153
rect 4093 119 4107 133
rect 4193 119 4207 133
rect 4233 127 4247 141
rect 4493 196 4507 210
rect 4333 167 4347 181
rect 4253 119 4267 133
rect 4273 127 4287 141
rect 3833 64 3847 78
rect 3973 70 3987 84
rect 4353 102 4367 116
rect 4413 139 4427 153
rect 4453 139 4467 153
rect 4873 196 4887 210
rect 4553 139 4567 153
rect 4573 147 4587 161
rect 4593 139 4607 153
rect 4653 139 4667 153
rect 4673 147 4687 161
rect 4693 139 4707 153
rect 4613 119 4627 133
rect 4713 119 4727 133
rect 4753 127 4767 141
rect 5013 196 5027 210
rect 4853 167 4867 181
rect 4773 119 4787 133
rect 4793 127 4807 141
rect 4353 64 4367 78
rect 4493 70 4507 84
rect 4873 102 4887 116
rect 4933 139 4947 153
rect 4973 139 4987 153
rect 5393 196 5407 210
rect 5113 139 5127 153
rect 5133 147 5147 161
rect 5153 139 5167 153
rect 5173 139 5187 153
rect 5193 147 5207 161
rect 5213 139 5227 153
rect 5093 119 5107 133
rect 5233 119 5247 133
rect 5273 127 5287 141
rect 5533 196 5547 210
rect 5373 167 5387 181
rect 5293 119 5307 133
rect 5313 127 5327 141
rect 4873 64 4887 78
rect 5013 70 5027 84
rect 5393 102 5407 116
rect 5453 139 5467 153
rect 5493 139 5507 153
rect 5393 64 5407 78
rect 5533 70 5547 84
rect 5633 196 5647 210
rect 5773 196 5787 210
rect 5613 167 5627 181
rect 5633 102 5647 116
rect 5693 139 5707 153
rect 5733 139 5747 153
rect 5633 64 5647 78
rect 5773 70 5787 84
rect 5873 196 5887 210
rect 6013 196 6027 210
rect 5853 167 5867 181
rect 5873 102 5887 116
rect 5933 139 5947 153
rect 5973 139 5987 153
rect 6093 139 6107 153
rect 6113 147 6127 161
rect 6133 139 6147 153
rect 6153 147 6167 161
rect 6173 139 6187 153
rect 6253 139 6267 153
rect 6273 147 6287 161
rect 6453 196 6467 210
rect 6593 196 6607 210
rect 6293 139 6307 153
rect 6313 147 6327 161
rect 6333 139 6347 153
rect 6373 147 6387 161
rect 6393 159 6407 173
rect 6433 167 6447 181
rect 6193 119 6207 133
rect 5873 64 5887 78
rect 6013 70 6027 84
rect 6453 102 6467 116
rect 6513 139 6527 153
rect 6553 139 6567 153
rect 6453 64 6467 78
rect 6593 70 6607 84
<< metal2 >>
rect 56 6324 64 6436
rect 136 6407 143 6413
rect 133 6393 147 6407
rect 57 6158 65 6182
rect 57 6064 65 6144
rect 156 6143 163 6413
rect 195 6356 203 6436
rect 447 6416 463 6423
rect 213 6393 227 6407
rect 216 6367 223 6393
rect 313 6373 327 6387
rect 456 6403 463 6416
rect 456 6396 483 6403
rect 195 6318 203 6342
rect 316 6187 323 6373
rect 393 6353 407 6367
rect 396 6347 403 6353
rect 416 6347 423 6393
rect 136 6136 163 6143
rect 113 6103 127 6107
rect 136 6103 143 6136
rect 113 6096 143 6103
rect 113 6093 127 6096
rect 76 5927 83 6093
rect 196 6064 204 6176
rect 396 6167 403 6313
rect 436 6163 443 6393
rect 476 6387 483 6396
rect 536 6387 543 6393
rect 473 6373 487 6387
rect 533 6373 547 6387
rect 553 6363 567 6367
rect 576 6363 583 6393
rect 616 6387 623 6393
rect 553 6356 583 6363
rect 637 6356 645 6436
rect 696 6407 703 6413
rect 736 6407 743 6433
rect 693 6393 707 6407
rect 733 6393 747 6407
rect 553 6353 567 6356
rect 637 6318 645 6342
rect 416 6156 443 6163
rect 416 6147 423 6156
rect 33 5923 47 5927
rect 73 5923 87 5927
rect 16 5916 47 5923
rect 16 5887 23 5916
rect 33 5913 47 5916
rect 56 5916 87 5923
rect 56 5887 63 5916
rect 73 5913 87 5916
rect 116 5907 123 6053
rect 113 5893 127 5907
rect 133 5873 147 5887
rect 173 5873 187 5887
rect 236 5887 243 6113
rect 393 6113 407 6127
rect 376 6067 383 6093
rect 396 6067 403 6113
rect 433 6093 447 6107
rect 473 6103 487 6107
rect 496 6103 503 6293
rect 516 6127 523 6173
rect 273 5923 287 5927
rect 256 5916 287 5923
rect 213 5873 227 5887
rect 136 5867 143 5873
rect 73 5623 87 5627
rect 73 5616 103 5623
rect 73 5613 87 5616
rect 33 5433 47 5447
rect 36 5427 43 5433
rect 57 5396 65 5476
rect 96 5427 103 5616
rect 113 5613 127 5627
rect 153 5623 167 5627
rect 176 5623 183 5873
rect 216 5867 223 5873
rect 217 5678 225 5702
rect 193 5623 207 5627
rect 153 5616 207 5623
rect 153 5613 167 5616
rect 193 5613 207 5616
rect 116 5607 123 5613
rect 217 5584 225 5664
rect 256 5627 263 5916
rect 273 5913 287 5916
rect 293 5893 307 5907
rect 396 5907 403 5953
rect 416 5947 423 6073
rect 436 5967 443 6093
rect 473 6096 503 6103
rect 473 6093 487 6096
rect 593 6093 607 6107
rect 633 6093 647 6107
rect 516 6047 523 6093
rect 556 6087 563 6093
rect 596 6083 603 6093
rect 636 6083 643 6093
rect 576 6076 603 6083
rect 616 6076 643 6083
rect 436 5947 443 5953
rect 433 5933 447 5947
rect 416 5927 423 5933
rect 296 5887 303 5893
rect 336 5887 343 5893
rect 393 5893 407 5907
rect 453 5893 467 5907
rect 456 5887 463 5893
rect 273 5613 287 5627
rect 116 5447 123 5453
rect 113 5433 127 5447
rect 57 5358 65 5382
rect 137 5198 145 5222
rect 116 5147 123 5153
rect 137 5104 145 5184
rect 176 5143 183 5453
rect 196 5364 204 5476
rect 276 5467 283 5613
rect 296 5603 303 5873
rect 496 5847 503 5993
rect 536 5947 543 5973
rect 533 5933 547 5947
rect 516 5927 523 5933
rect 556 5927 563 6073
rect 576 5963 583 6076
rect 616 6047 623 6076
rect 576 5956 603 5963
rect 596 5947 603 5956
rect 553 5913 567 5927
rect 616 5927 623 5993
rect 656 5987 663 6093
rect 656 5947 663 5973
rect 676 5947 683 6353
rect 776 6324 784 6436
rect 833 6423 847 6427
rect 816 6416 847 6423
rect 816 6403 823 6416
rect 796 6396 823 6403
rect 833 6413 847 6416
rect 936 6407 943 6433
rect 1053 6423 1067 6427
rect 1053 6416 1083 6423
rect 1053 6413 1067 6416
rect 893 6403 907 6407
rect 796 6387 803 6396
rect 876 6396 907 6403
rect 876 6387 883 6396
rect 893 6393 907 6396
rect 853 6373 867 6387
rect 913 6373 927 6387
rect 933 6393 947 6407
rect 973 6403 987 6407
rect 953 6373 967 6387
rect 973 6396 1003 6403
rect 973 6393 987 6396
rect 816 6347 823 6373
rect 856 6367 863 6373
rect 916 6367 923 6373
rect 756 6127 763 6153
rect 816 6127 823 6333
rect 956 6287 963 6373
rect 836 6143 843 6153
rect 836 6136 863 6143
rect 713 6113 727 6127
rect 716 6107 723 6113
rect 753 6113 767 6127
rect 773 6103 787 6107
rect 793 6103 807 6107
rect 773 6096 807 6103
rect 833 6103 847 6107
rect 856 6103 863 6136
rect 773 6093 787 6096
rect 793 6093 807 6096
rect 736 6083 743 6093
rect 716 6076 743 6083
rect 696 6047 703 6073
rect 613 5913 627 5927
rect 653 5923 667 5927
rect 647 5916 667 5923
rect 653 5913 667 5916
rect 296 5596 323 5603
rect 293 5393 307 5407
rect 296 5387 303 5393
rect 316 5367 323 5596
rect 356 5584 364 5696
rect 536 5667 543 5893
rect 636 5887 643 5913
rect 673 5893 687 5907
rect 716 5907 723 6076
rect 713 5893 727 5907
rect 436 5547 443 5613
rect 473 5613 487 5627
rect 516 5643 523 5653
rect 533 5643 547 5647
rect 516 5636 547 5643
rect 533 5633 547 5636
rect 456 5587 463 5593
rect 476 5583 483 5613
rect 553 5613 567 5627
rect 476 5576 503 5583
rect 193 5143 207 5147
rect 176 5136 207 5143
rect 76 4967 83 5013
rect 73 4953 87 4967
rect 176 4707 183 5136
rect 193 5133 207 5136
rect 233 5133 247 5147
rect 196 5127 203 5133
rect 236 5107 243 5133
rect 276 5104 284 5216
rect 336 5207 343 5473
rect 373 5413 387 5427
rect 476 5427 483 5553
rect 496 5507 503 5576
rect 556 5547 563 5613
rect 413 5413 427 5427
rect 376 5367 383 5413
rect 416 5407 423 5413
rect 473 5413 487 5427
rect 493 5403 507 5407
rect 516 5403 523 5453
rect 536 5447 543 5533
rect 533 5433 547 5447
rect 493 5396 523 5403
rect 493 5393 507 5396
rect 536 5367 543 5393
rect 576 5387 583 5853
rect 636 5687 643 5853
rect 613 5633 627 5647
rect 596 5547 603 5613
rect 616 5527 623 5633
rect 616 5463 623 5493
rect 636 5483 643 5613
rect 656 5603 663 5873
rect 676 5847 683 5893
rect 736 5727 743 5913
rect 676 5667 683 5693
rect 713 5663 727 5667
rect 696 5656 727 5663
rect 756 5663 763 5973
rect 776 5947 783 6073
rect 796 5987 803 6093
rect 833 6096 863 6103
rect 876 6103 883 6273
rect 996 6167 1003 6396
rect 1076 6403 1083 6416
rect 1093 6403 1107 6407
rect 1076 6396 1107 6403
rect 1076 6307 1083 6396
rect 1093 6393 1107 6396
rect 1117 6356 1125 6436
rect 1176 6407 1183 6413
rect 1216 6407 1223 6433
rect 1173 6393 1187 6407
rect 1213 6393 1227 6407
rect 1117 6318 1125 6342
rect 893 6103 907 6107
rect 876 6096 907 6103
rect 833 6093 847 6096
rect 893 6093 907 6096
rect 813 6073 827 6087
rect 816 6047 823 6073
rect 796 5947 803 5953
rect 836 5947 843 6093
rect 1033 6123 1047 6127
rect 1056 6123 1063 6153
rect 1033 6116 1063 6123
rect 1033 6113 1047 6116
rect 933 6073 947 6087
rect 993 6093 1007 6107
rect 973 6073 987 6087
rect 936 6067 943 6073
rect 896 5967 903 6033
rect 793 5933 807 5947
rect 833 5933 847 5947
rect 773 5893 787 5907
rect 856 5927 863 5933
rect 853 5913 867 5927
rect 776 5867 783 5893
rect 816 5687 823 5873
rect 876 5867 883 5913
rect 896 5667 903 5953
rect 976 5927 983 6073
rect 996 6067 1003 6093
rect 996 5907 1003 5953
rect 1016 5927 1023 6113
rect 1113 6083 1127 6087
rect 1096 6076 1127 6083
rect 1096 5947 1103 6076
rect 1113 6073 1127 6076
rect 1093 5933 1107 5947
rect 993 5893 1007 5907
rect 953 5873 967 5887
rect 773 5663 787 5667
rect 756 5656 787 5663
rect 813 5663 827 5667
rect 853 5663 867 5667
rect 656 5596 683 5603
rect 636 5476 663 5483
rect 633 5463 647 5467
rect 616 5456 647 5463
rect 633 5453 647 5456
rect 656 5447 663 5476
rect 676 5387 683 5596
rect 696 5587 703 5656
rect 713 5653 727 5656
rect 773 5653 787 5656
rect 813 5656 867 5663
rect 813 5653 827 5656
rect 733 5613 747 5627
rect 736 5607 743 5613
rect 696 5447 703 5493
rect 716 5467 723 5473
rect 713 5453 727 5467
rect 693 5433 707 5447
rect 736 5447 743 5533
rect 733 5433 747 5447
rect 796 5427 803 5453
rect 816 5443 823 5613
rect 836 5607 843 5656
rect 853 5653 867 5656
rect 873 5633 887 5647
rect 893 5653 907 5667
rect 876 5627 883 5633
rect 916 5527 923 5713
rect 956 5707 963 5873
rect 976 5847 983 5893
rect 1036 5687 1043 5893
rect 1096 5867 1103 5893
rect 973 5613 987 5627
rect 953 5593 967 5607
rect 956 5547 963 5593
rect 976 5547 983 5613
rect 996 5607 1003 5633
rect 1013 5593 1027 5607
rect 816 5436 843 5443
rect 836 5427 843 5436
rect 876 5427 883 5473
rect 933 5463 947 5467
rect 916 5456 947 5463
rect 773 5393 787 5407
rect 793 5413 807 5427
rect 813 5403 827 5407
rect 813 5396 843 5403
rect 813 5393 827 5396
rect 376 5187 383 5193
rect 333 5183 347 5187
rect 316 5176 347 5183
rect 316 5167 323 5176
rect 333 5173 347 5176
rect 373 5173 387 5187
rect 416 5167 423 5353
rect 496 5167 503 5173
rect 193 4913 207 4927
rect 276 4927 283 4953
rect 297 4916 305 4996
rect 196 4907 203 4913
rect 297 4878 305 4902
rect 176 4687 183 4693
rect 33 4683 47 4687
rect 16 4676 47 4683
rect 16 4447 23 4676
rect 33 4673 47 4676
rect 173 4673 187 4687
rect 273 4653 287 4667
rect 253 4633 267 4647
rect 256 4603 263 4633
rect 276 4627 283 4653
rect 296 4643 303 4773
rect 336 4687 343 5133
rect 356 4967 363 5113
rect 353 4953 367 4967
rect 416 4787 423 5153
rect 433 5133 447 5147
rect 493 5153 507 5167
rect 436 5107 443 5133
rect 516 5127 523 5213
rect 576 5187 583 5213
rect 596 5207 603 5373
rect 573 5173 587 5187
rect 436 4884 444 4996
rect 556 4987 563 4993
rect 553 4973 567 4987
rect 573 4933 587 4947
rect 556 4927 563 4933
rect 576 4927 583 4933
rect 596 4907 603 5193
rect 616 5167 623 5353
rect 636 5104 644 5216
rect 616 4967 623 4993
rect 636 4947 643 4993
rect 696 4967 703 5373
rect 713 5133 727 5147
rect 716 5127 723 5133
rect 736 5127 743 5393
rect 776 5387 783 5393
rect 776 5367 783 5373
rect 775 5198 783 5222
rect 816 5207 823 5373
rect 775 5104 783 5184
rect 796 5147 803 5173
rect 793 5133 807 5147
rect 736 4967 743 4993
rect 816 4987 823 5193
rect 836 5187 843 5396
rect 853 5393 867 5407
rect 873 5413 887 5427
rect 893 5403 907 5407
rect 916 5403 923 5456
rect 933 5453 947 5456
rect 953 5413 967 5427
rect 976 5423 983 5513
rect 996 5463 1003 5593
rect 1016 5587 1023 5593
rect 1056 5587 1063 5853
rect 1073 5593 1087 5607
rect 1076 5527 1083 5593
rect 1116 5547 1123 5673
rect 1136 5663 1143 6093
rect 1173 6093 1187 6107
rect 1153 6073 1167 6087
rect 1156 6047 1163 6073
rect 1176 6067 1183 6093
rect 1196 6007 1203 6373
rect 1256 6324 1264 6436
rect 1296 6303 1303 6413
rect 1356 6407 1363 6433
rect 1333 6373 1347 6387
rect 1353 6393 1367 6407
rect 1393 6403 1407 6407
rect 1393 6396 1413 6403
rect 1393 6393 1407 6396
rect 1473 6403 1487 6407
rect 1467 6396 1487 6403
rect 1513 6403 1527 6407
rect 1473 6393 1487 6396
rect 1453 6383 1467 6387
rect 1436 6376 1467 6383
rect 1336 6367 1343 6373
rect 1436 6367 1443 6376
rect 1453 6373 1467 6376
rect 1513 6396 1543 6403
rect 1513 6393 1527 6396
rect 1536 6367 1543 6396
rect 1613 6403 1627 6407
rect 1596 6396 1627 6403
rect 1596 6387 1603 6396
rect 1613 6393 1627 6396
rect 1296 6296 1323 6303
rect 1216 6123 1223 6153
rect 1233 6123 1247 6127
rect 1216 6116 1247 6123
rect 1233 6113 1247 6116
rect 1253 6093 1267 6107
rect 1236 5967 1243 6093
rect 1256 6007 1263 6093
rect 1156 5903 1163 5953
rect 1193 5943 1207 5947
rect 1193 5936 1223 5943
rect 1193 5933 1207 5936
rect 1216 5927 1223 5936
rect 1233 5913 1247 5927
rect 1173 5903 1187 5907
rect 1156 5896 1187 5903
rect 1173 5893 1187 5896
rect 1216 5683 1223 5913
rect 1236 5707 1243 5913
rect 1257 5876 1265 5956
rect 1316 5927 1323 6296
rect 1436 6267 1443 6353
rect 1333 6123 1347 6127
rect 1356 6123 1363 6153
rect 1393 6123 1407 6127
rect 1333 6116 1363 6123
rect 1376 6116 1407 6123
rect 1333 6113 1347 6116
rect 1353 6073 1367 6087
rect 1356 6047 1363 6073
rect 1376 6067 1383 6116
rect 1393 6113 1407 6116
rect 1473 6093 1487 6107
rect 1513 6093 1527 6107
rect 1476 6047 1483 6093
rect 1516 6067 1523 6093
rect 1576 6067 1583 6353
rect 1596 6147 1603 6373
rect 1616 6127 1623 6153
rect 1613 6113 1627 6127
rect 1636 6107 1643 6433
rect 1676 6427 1683 6433
rect 1673 6423 1687 6427
rect 1673 6416 1703 6423
rect 1673 6413 1687 6416
rect 1696 6403 1703 6416
rect 1713 6403 1727 6407
rect 1696 6396 1727 6403
rect 1713 6393 1727 6396
rect 1737 6356 1745 6436
rect 1796 6407 1803 6413
rect 1793 6393 1807 6407
rect 1737 6318 1745 6342
rect 1716 6127 1723 6153
rect 1756 6127 1763 6373
rect 1796 6147 1803 6353
rect 1876 6324 1884 6436
rect 1933 6403 1947 6407
rect 1916 6396 1947 6403
rect 1916 6387 1923 6396
rect 1933 6393 1947 6396
rect 1953 6373 1967 6387
rect 1996 6387 2003 6393
rect 1993 6373 2007 6387
rect 1956 6247 1963 6373
rect 2033 6353 2047 6367
rect 2133 6383 2147 6387
rect 2116 6376 2147 6383
rect 2016 6127 2023 6273
rect 2036 6267 2043 6353
rect 2056 6127 2063 6133
rect 2076 6127 2083 6153
rect 2096 6143 2103 6313
rect 2116 6267 2123 6376
rect 2133 6373 2147 6376
rect 2253 6373 2267 6387
rect 2293 6373 2307 6387
rect 2096 6136 2123 6143
rect 1653 6093 1667 6107
rect 1656 6027 1663 6093
rect 1733 6093 1747 6107
rect 1673 6073 1687 6087
rect 1676 6047 1683 6073
rect 1696 6027 1703 6073
rect 1716 6003 1723 6093
rect 1696 5996 1723 6003
rect 1313 5923 1327 5927
rect 1296 5916 1327 5923
rect 1257 5838 1265 5862
rect 1216 5676 1243 5683
rect 1136 5656 1163 5663
rect 1013 5463 1027 5467
rect 996 5456 1027 5463
rect 1013 5453 1027 5456
rect 993 5423 1007 5427
rect 976 5416 1007 5423
rect 993 5413 1007 5416
rect 1033 5413 1047 5427
rect 893 5396 923 5403
rect 893 5393 907 5396
rect 856 5367 863 5393
rect 916 5387 923 5396
rect 956 5403 963 5413
rect 1016 5407 1023 5413
rect 1036 5407 1043 5413
rect 956 5396 973 5403
rect 936 5227 943 5393
rect 876 5187 883 5193
rect 873 5173 887 5187
rect 1016 5163 1023 5273
rect 1076 5187 1083 5473
rect 1096 5403 1103 5533
rect 1136 5463 1143 5593
rect 1156 5487 1163 5656
rect 1173 5613 1187 5627
rect 1176 5567 1183 5613
rect 1213 5613 1227 5627
rect 1193 5593 1207 5607
rect 1196 5587 1203 5593
rect 1216 5587 1223 5613
rect 1236 5607 1243 5676
rect 1296 5647 1303 5916
rect 1313 5913 1327 5916
rect 1396 5844 1404 5956
rect 1476 5907 1483 5913
rect 1656 5907 1663 5993
rect 1696 5947 1703 5996
rect 1736 5987 1743 6093
rect 1776 6087 1783 6093
rect 1796 6087 1803 6113
rect 1813 6093 1827 6107
rect 1853 6093 1867 6107
rect 1716 5927 1723 5973
rect 1756 5927 1763 6053
rect 1776 5967 1783 6053
rect 1773 5943 1787 5947
rect 1796 5943 1803 5993
rect 1816 5987 1823 6093
rect 1773 5936 1803 5943
rect 1773 5933 1787 5936
rect 1453 5873 1467 5887
rect 1473 5893 1487 5907
rect 1456 5847 1463 5873
rect 1536 5867 1543 5893
rect 1613 5903 1627 5907
rect 1613 5896 1643 5903
rect 1613 5893 1627 5896
rect 1497 5678 1505 5702
rect 1413 5643 1427 5647
rect 1253 5593 1267 5607
rect 1256 5567 1263 5593
rect 1116 5456 1143 5463
rect 1116 5447 1123 5456
rect 1113 5433 1127 5447
rect 1193 5443 1207 5447
rect 1173 5413 1187 5427
rect 1193 5436 1223 5443
rect 1193 5433 1207 5436
rect 1176 5407 1183 5413
rect 1096 5396 1123 5403
rect 1116 5167 1123 5396
rect 1033 5163 1047 5167
rect 1016 5156 1047 5163
rect 1033 5153 1047 5156
rect 993 5133 1007 5147
rect 1053 5133 1067 5147
rect 996 5127 1003 5133
rect 1016 5107 1023 5133
rect 1056 5127 1063 5133
rect 1116 5087 1123 5153
rect 1133 5133 1147 5147
rect 1193 5133 1207 5147
rect 1136 5107 1143 5133
rect 1196 5087 1203 5133
rect 853 4953 867 4967
rect 633 4933 647 4947
rect 676 4903 683 4913
rect 736 4903 743 4933
rect 656 4896 683 4903
rect 696 4896 743 4903
rect 473 4683 487 4687
rect 456 4676 487 4683
rect 296 4636 323 4643
rect 256 4596 283 4603
rect 76 4467 83 4513
rect 136 4487 143 4553
rect 133 4473 147 4487
rect 216 4487 223 4513
rect 256 4487 263 4573
rect 276 4487 283 4596
rect 213 4473 227 4487
rect 253 4473 267 4487
rect 273 4463 287 4467
rect 296 4463 303 4593
rect 316 4487 323 4636
rect 413 4633 427 4647
rect 336 4607 343 4613
rect 336 4487 343 4533
rect 356 4507 363 4613
rect 376 4507 383 4633
rect 333 4473 347 4487
rect 396 4487 403 4573
rect 416 4547 423 4633
rect 456 4567 463 4676
rect 473 4673 487 4676
rect 516 4647 523 4673
rect 573 4653 587 4667
rect 576 4647 583 4653
rect 596 4623 603 4893
rect 616 4887 623 4893
rect 636 4707 643 4853
rect 633 4693 647 4707
rect 656 4647 663 4896
rect 696 4887 703 4896
rect 756 4887 763 4933
rect 773 4913 787 4927
rect 836 4927 843 4953
rect 856 4947 863 4953
rect 877 4916 885 4996
rect 896 4947 903 5013
rect 976 4967 983 4993
rect 933 4963 947 4967
rect 933 4956 963 4963
rect 933 4953 947 4956
rect 956 4947 963 4956
rect 973 4953 987 4967
rect 776 4907 783 4913
rect 736 4747 743 4873
rect 673 4663 687 4667
rect 693 4663 707 4667
rect 673 4656 707 4663
rect 733 4663 747 4667
rect 756 4663 763 4853
rect 836 4707 843 4893
rect 877 4878 885 4902
rect 1016 4884 1024 4996
rect 1036 4843 1043 5073
rect 1016 4836 1043 4843
rect 977 4718 985 4742
rect 873 4703 887 4707
rect 856 4696 887 4703
rect 673 4653 687 4656
rect 693 4653 707 4656
rect 576 4616 603 4623
rect 416 4527 423 4533
rect 436 4487 443 4533
rect 456 4487 463 4553
rect 496 4507 503 4533
rect 493 4493 507 4507
rect 373 4483 387 4487
rect 393 4483 407 4487
rect 273 4456 303 4463
rect 273 4453 287 4456
rect 373 4476 407 4483
rect 373 4473 387 4476
rect 393 4473 407 4476
rect 516 4487 523 4493
rect 453 4463 467 4467
rect 453 4456 483 4463
rect 453 4453 467 4456
rect 16 3023 23 4433
rect 96 4203 103 4313
rect 156 4247 163 4453
rect 196 4223 203 4453
rect 316 4443 323 4453
rect 316 4436 343 4443
rect 336 4407 343 4436
rect 196 4216 223 4223
rect 156 4207 163 4213
rect 216 4207 223 4216
rect 113 4203 127 4207
rect 96 4196 127 4203
rect 113 4193 127 4196
rect 73 4173 87 4187
rect 133 4173 147 4187
rect 153 4193 167 4207
rect 193 4173 207 4187
rect 213 4193 227 4207
rect 253 4193 267 4207
rect 256 4187 263 4193
rect 233 4173 247 4187
rect 76 4167 83 4173
rect 136 4163 143 4173
rect 196 4163 203 4173
rect 136 4156 203 4163
rect 236 4147 243 4173
rect 276 4167 283 4193
rect 336 4144 344 4256
rect 356 4127 363 4453
rect 416 4443 423 4453
rect 376 4436 423 4443
rect 376 4407 383 4436
rect 476 4427 483 4456
rect 553 4453 567 4467
rect 376 4227 383 4393
rect 556 4267 563 4453
rect 475 4238 483 4262
rect 576 4247 583 4616
rect 653 4483 667 4487
rect 633 4453 647 4467
rect 653 4476 683 4483
rect 653 4473 667 4476
rect 373 4173 387 4187
rect 436 4187 443 4213
rect 413 4173 427 4187
rect 376 4147 383 4173
rect 416 4167 423 4173
rect 33 4003 47 4007
rect 33 3996 63 4003
rect 33 3993 47 3996
rect 56 3967 63 3996
rect 116 3967 123 3993
rect 137 3956 145 4036
rect 196 4007 203 4013
rect 193 3993 207 4007
rect 137 3918 145 3942
rect 276 3924 284 4036
rect 416 3987 423 4113
rect 456 4027 463 4153
rect 475 4144 483 4224
rect 533 4223 547 4227
rect 516 4216 547 4223
rect 493 4183 507 4187
rect 516 4183 523 4216
rect 533 4213 547 4216
rect 493 4176 523 4183
rect 493 4173 507 4176
rect 493 3973 507 3987
rect 373 3953 387 3967
rect 376 3947 383 3953
rect 297 3758 305 3782
rect 196 3747 203 3753
rect 193 3733 207 3747
rect 233 3743 247 3747
rect 73 3693 87 3707
rect 113 3693 127 3707
rect 233 3736 263 3743
rect 233 3733 247 3736
rect 256 3707 263 3736
rect 273 3703 287 3707
rect 267 3696 287 3703
rect 273 3693 287 3696
rect 76 3667 83 3693
rect 116 3687 123 3693
rect 297 3664 305 3744
rect 353 3693 367 3707
rect 356 3687 363 3693
rect 416 3607 423 3973
rect 496 3967 503 3973
rect 516 3943 523 4176
rect 556 3987 563 4013
rect 553 3973 567 3987
rect 596 3947 603 4233
rect 616 4027 623 4453
rect 636 4407 643 4453
rect 636 4227 643 4393
rect 676 4223 683 4476
rect 696 4403 703 4653
rect 733 4656 763 4663
rect 733 4653 747 4656
rect 793 4653 807 4667
rect 796 4647 803 4653
rect 816 4647 823 4673
rect 713 4633 727 4647
rect 716 4627 723 4633
rect 856 4627 863 4696
rect 873 4693 887 4696
rect 936 4663 943 4693
rect 953 4663 967 4667
rect 936 4656 967 4663
rect 953 4653 967 4656
rect 736 4527 743 4533
rect 736 4507 743 4513
rect 776 4507 783 4573
rect 733 4493 747 4507
rect 773 4493 787 4507
rect 713 4453 727 4467
rect 796 4487 803 4513
rect 793 4473 807 4487
rect 716 4427 723 4453
rect 816 4407 823 4613
rect 896 4507 903 4653
rect 977 4624 985 4704
rect 916 4507 923 4533
rect 913 4493 927 4507
rect 696 4396 723 4403
rect 656 4216 683 4223
rect 656 4207 663 4216
rect 696 4207 703 4253
rect 716 4223 723 4396
rect 716 4216 733 4223
rect 756 4207 763 4253
rect 837 4238 845 4262
rect 633 4173 647 4187
rect 653 4193 667 4207
rect 673 4173 687 4187
rect 693 4193 707 4207
rect 713 4173 727 4187
rect 753 4193 767 4207
rect 636 4167 643 4173
rect 676 4147 683 4173
rect 636 3987 643 3993
rect 613 3953 627 3967
rect 676 3963 683 4113
rect 716 4107 723 4173
rect 747 4156 763 4163
rect 696 4007 703 4033
rect 736 4007 743 4013
rect 693 3993 707 4007
rect 676 3956 703 3963
rect 616 3947 623 3953
rect 516 3936 573 3943
rect 436 3664 444 3776
rect 456 3627 463 3913
rect 576 3763 583 3773
rect 596 3767 603 3933
rect 516 3756 583 3763
rect 516 3743 523 3756
rect 496 3736 523 3743
rect 116 3487 123 3513
rect 137 3476 145 3556
rect 196 3527 203 3533
rect 236 3527 243 3573
rect 193 3513 207 3527
rect 233 3513 247 3527
rect 137 3438 145 3462
rect 216 3447 223 3493
rect 276 3444 284 3556
rect 416 3527 423 3553
rect 456 3527 463 3593
rect 476 3547 483 3673
rect 496 3647 503 3736
rect 536 3727 543 3733
rect 576 3727 583 3733
rect 533 3713 547 3727
rect 556 3647 563 3673
rect 137 3278 145 3302
rect 116 3227 123 3233
rect 137 3184 145 3264
rect 193 3213 207 3227
rect 33 3023 47 3027
rect 16 3016 47 3023
rect 33 3013 47 3016
rect 196 3027 203 3213
rect 276 3184 284 3296
rect 173 3023 187 3027
rect 173 3016 193 3023
rect 173 3013 187 3016
rect 273 3043 287 3047
rect 273 3036 303 3043
rect 273 3033 287 3036
rect 36 2783 43 3013
rect 296 2947 303 3036
rect 36 2776 63 2783
rect 13 2713 27 2727
rect 16 2563 23 2713
rect 56 2647 63 2776
rect 133 2733 147 2747
rect 136 2727 143 2733
rect 33 2563 47 2567
rect 16 2556 47 2563
rect 33 2553 47 2556
rect 57 2516 65 2596
rect 116 2567 123 2593
rect 113 2553 127 2567
rect 57 2478 65 2502
rect 136 2363 143 2713
rect 196 2704 204 2816
rect 273 2733 287 2747
rect 156 2587 163 2693
rect 153 2563 167 2567
rect 153 2556 183 2563
rect 153 2553 167 2556
rect 116 2356 143 2363
rect 56 2224 64 2336
rect 56 2107 63 2173
rect 53 2093 67 2107
rect 116 2103 123 2356
rect 133 2263 147 2267
rect 156 2263 163 2513
rect 133 2256 163 2263
rect 133 2253 147 2256
rect 176 2187 183 2556
rect 196 2484 204 2596
rect 195 2318 203 2342
rect 195 2224 203 2304
rect 236 2247 243 2273
rect 216 2127 223 2213
rect 96 2096 123 2103
rect 33 2083 47 2087
rect 16 2076 47 2083
rect 73 2083 87 2087
rect 96 2083 103 2096
rect 16 2043 23 2076
rect 33 2073 47 2076
rect 73 2076 103 2083
rect 73 2073 87 2076
rect 16 2036 43 2043
rect 36 1807 43 2036
rect 56 2007 63 2053
rect 76 1987 83 2033
rect 96 2027 103 2076
rect 136 2067 143 2093
rect 113 2033 127 2047
rect 133 2053 147 2067
rect 116 2007 123 2033
rect 96 1847 103 1993
rect 156 1907 163 2013
rect 176 2007 183 2073
rect 216 2067 223 2093
rect 213 2053 227 2067
rect 236 2063 243 2213
rect 256 2083 263 2633
rect 276 2607 283 2733
rect 316 2663 323 3513
rect 453 3513 467 3527
rect 376 3267 383 3273
rect 373 3253 387 3267
rect 416 3247 423 3293
rect 456 3247 463 3253
rect 476 3247 483 3533
rect 516 3527 523 3573
rect 556 3547 563 3573
rect 553 3533 567 3547
rect 513 3513 527 3527
rect 573 3493 587 3507
rect 576 3467 583 3493
rect 596 3487 603 3753
rect 616 3747 623 3753
rect 656 3747 663 3773
rect 676 3747 683 3773
rect 696 3763 703 3956
rect 756 3927 763 4156
rect 773 4153 787 4167
rect 776 4127 783 4153
rect 796 4107 803 4213
rect 816 4187 823 4213
rect 813 4173 827 4187
rect 837 4144 845 4224
rect 797 3956 805 4036
rect 856 4007 863 4173
rect 876 4127 883 4213
rect 896 4167 903 4173
rect 896 4007 903 4053
rect 853 4003 867 4007
rect 836 3996 867 4003
rect 776 3787 783 3953
rect 797 3918 805 3942
rect 696 3756 723 3763
rect 716 3747 723 3756
rect 613 3733 627 3747
rect 633 3713 647 3727
rect 653 3733 667 3747
rect 673 3733 687 3747
rect 693 3713 707 3727
rect 713 3733 727 3747
rect 736 3727 743 3733
rect 636 3627 643 3713
rect 696 3687 703 3713
rect 736 3647 743 3713
rect 756 3703 763 3773
rect 776 3747 783 3753
rect 816 3747 823 3773
rect 773 3733 787 3747
rect 813 3733 827 3747
rect 836 3707 843 3996
rect 853 3993 867 3996
rect 893 3993 907 4007
rect 856 3707 863 3773
rect 877 3758 885 3782
rect 756 3696 783 3703
rect 696 3527 703 3633
rect 736 3527 743 3553
rect 756 3527 763 3553
rect 776 3527 783 3696
rect 877 3664 885 3744
rect 896 3667 903 3693
rect 916 3667 923 4453
rect 933 4173 947 4187
rect 936 4147 943 4173
rect 936 3924 944 4036
rect 933 3693 947 3707
rect 936 3687 943 3693
rect 796 3527 803 3533
rect 733 3513 747 3527
rect 613 3473 627 3487
rect 653 3483 667 3487
rect 653 3476 683 3483
rect 653 3473 667 3476
rect 496 3267 503 3293
rect 536 3267 543 3273
rect 576 3267 583 3293
rect 596 3287 603 3473
rect 616 3467 623 3473
rect 676 3467 683 3476
rect 533 3253 547 3267
rect 496 3247 503 3253
rect 453 3233 467 3247
rect 493 3233 507 3247
rect 553 3233 567 3247
rect 573 3253 587 3267
rect 596 3247 603 3273
rect 616 3247 623 3313
rect 636 3287 643 3293
rect 656 3287 663 3453
rect 716 3283 723 3513
rect 753 3513 767 3527
rect 793 3513 807 3527
rect 776 3467 783 3493
rect 816 3483 823 3513
rect 856 3507 863 3573
rect 916 3507 923 3653
rect 956 3567 963 4593
rect 976 4507 983 4513
rect 973 4503 987 4507
rect 996 4503 1003 4793
rect 973 4496 1003 4503
rect 973 4493 987 4496
rect 1016 4443 1023 4836
rect 1033 4653 1047 4667
rect 1036 4647 1043 4653
rect 1056 4507 1063 5033
rect 1096 4967 1103 4973
rect 1136 4967 1143 5033
rect 1176 4967 1183 4993
rect 1196 4983 1203 5013
rect 1216 5007 1223 5436
rect 1233 5433 1247 5447
rect 1236 5387 1243 5433
rect 1257 5396 1265 5476
rect 1296 5467 1303 5633
rect 1353 5613 1367 5627
rect 1413 5636 1433 5643
rect 1413 5633 1427 5636
rect 1356 5607 1363 5613
rect 1436 5607 1443 5633
rect 1473 5623 1487 5627
rect 1456 5616 1487 5623
rect 1393 5593 1407 5607
rect 1396 5587 1403 5593
rect 1456 5587 1463 5616
rect 1473 5613 1487 5616
rect 1497 5584 1505 5664
rect 1553 5613 1567 5627
rect 1556 5607 1563 5613
rect 1316 5447 1323 5453
rect 1313 5433 1327 5447
rect 1257 5358 1265 5382
rect 1396 5364 1404 5476
rect 1616 5463 1623 5833
rect 1636 5787 1643 5896
rect 1653 5893 1667 5907
rect 1713 5913 1727 5927
rect 1753 5913 1767 5927
rect 1716 5776 1733 5783
rect 1636 5584 1644 5696
rect 1716 5647 1723 5776
rect 1776 5663 1783 5893
rect 1816 5867 1823 5953
rect 1856 5907 1863 6093
rect 1913 6073 1927 6087
rect 1916 6067 1923 6073
rect 1916 5947 1923 5973
rect 1913 5933 1927 5947
rect 1853 5893 1867 5907
rect 1876 5887 1883 5913
rect 1776 5656 1803 5663
rect 1676 5623 1683 5633
rect 1693 5623 1707 5627
rect 1676 5616 1707 5623
rect 1713 5633 1727 5647
rect 1693 5613 1707 5616
rect 1773 5623 1787 5627
rect 1796 5623 1803 5656
rect 1876 5647 1883 5673
rect 1896 5667 1903 5813
rect 1833 5633 1847 5647
rect 1836 5627 1843 5633
rect 1773 5616 1803 5623
rect 1773 5613 1787 5616
rect 1853 5613 1867 5627
rect 1873 5633 1887 5647
rect 1776 5467 1783 5593
rect 1596 5456 1623 5463
rect 1536 5427 1543 5433
rect 1596 5427 1603 5456
rect 1656 5447 1663 5453
rect 1473 5393 1487 5407
rect 1533 5413 1547 5427
rect 1593 5413 1607 5427
rect 1616 5407 1623 5433
rect 1736 5447 1743 5453
rect 1633 5423 1647 5427
rect 1633 5416 1663 5423
rect 1633 5413 1647 5416
rect 1656 5407 1663 5416
rect 1257 5198 1265 5222
rect 1236 5147 1243 5153
rect 1257 5104 1265 5184
rect 1313 5133 1327 5147
rect 1353 5143 1367 5147
rect 1376 5143 1383 5173
rect 1353 5136 1383 5143
rect 1353 5133 1367 5136
rect 1316 5127 1323 5133
rect 1213 4983 1227 4987
rect 1196 4976 1227 4983
rect 1236 4983 1243 5093
rect 1256 5007 1263 5013
rect 1236 4976 1263 4983
rect 1213 4973 1227 4976
rect 1093 4953 1107 4967
rect 1133 4953 1147 4967
rect 1173 4953 1187 4967
rect 1156 4927 1163 4953
rect 1233 4933 1247 4947
rect 1236 4927 1243 4933
rect 1116 4624 1124 4736
rect 1156 4587 1163 4913
rect 1053 4453 1067 4467
rect 1056 4447 1063 4453
rect 996 4436 1023 4443
rect 976 4144 984 4256
rect 973 3693 987 3707
rect 976 3627 983 3693
rect 833 3483 847 3487
rect 816 3476 847 3483
rect 833 3473 847 3476
rect 873 3473 887 3487
rect 716 3276 743 3283
rect 613 3233 627 3247
rect 556 3227 563 3233
rect 336 2964 344 3076
rect 376 3047 383 3093
rect 373 3033 387 3047
rect 456 3027 463 3193
rect 516 3187 523 3213
rect 335 2798 343 2822
rect 335 2704 343 2784
rect 413 2763 427 2767
rect 413 2756 443 2763
rect 413 2753 427 2756
rect 353 2743 367 2747
rect 353 2736 383 2743
rect 353 2733 367 2736
rect 376 2723 383 2736
rect 436 2727 443 2756
rect 456 2727 463 3013
rect 475 2996 483 3076
rect 493 3033 507 3047
rect 496 3007 503 3033
rect 516 3007 523 3053
rect 556 3047 563 3193
rect 576 3047 583 3213
rect 636 3227 643 3253
rect 673 3253 687 3267
rect 593 3193 607 3207
rect 596 3187 603 3193
rect 676 3187 683 3253
rect 736 3227 743 3276
rect 793 3263 807 3267
rect 773 3233 787 3247
rect 793 3256 823 3263
rect 793 3253 807 3256
rect 676 3047 683 3053
rect 636 3027 643 3033
rect 696 3027 703 3213
rect 756 3167 763 3213
rect 736 3047 743 3093
rect 756 3063 763 3093
rect 776 3087 783 3233
rect 816 3227 823 3256
rect 836 3243 843 3313
rect 876 3307 883 3473
rect 896 3247 903 3313
rect 916 3267 923 3493
rect 956 3267 963 3553
rect 996 3487 1003 4436
rect 1056 4387 1063 4433
rect 1076 4227 1083 4233
rect 1033 4223 1047 4227
rect 1016 4216 1047 4223
rect 1016 4207 1023 4216
rect 1033 4213 1047 4216
rect 1073 4213 1087 4227
rect 1116 4207 1123 4573
rect 1176 4463 1183 4913
rect 1216 4907 1223 4913
rect 1236 4887 1243 4913
rect 1256 4807 1263 4976
rect 1316 4967 1323 5113
rect 1396 5104 1404 5216
rect 1476 5187 1483 5393
rect 1516 5187 1523 5193
rect 1473 5173 1487 5187
rect 1513 5173 1527 5187
rect 1573 5183 1587 5187
rect 1573 5176 1603 5183
rect 1573 5173 1587 5176
rect 1356 4987 1363 4993
rect 1356 4967 1363 4973
rect 1396 4967 1403 5033
rect 1353 4953 1367 4967
rect 1393 4953 1407 4967
rect 1313 4923 1327 4927
rect 1336 4923 1343 4933
rect 1313 4916 1343 4923
rect 1313 4913 1327 4916
rect 1413 4913 1427 4927
rect 1453 4913 1467 4927
rect 1496 4923 1503 4973
rect 1513 4923 1527 4927
rect 1496 4916 1527 4923
rect 1513 4913 1527 4916
rect 1553 4913 1567 4927
rect 1316 4907 1323 4913
rect 1416 4907 1423 4913
rect 1456 4887 1463 4913
rect 1556 4887 1563 4913
rect 1236 4687 1243 4693
rect 1276 4687 1283 4873
rect 1296 4707 1303 4713
rect 1336 4707 1343 4773
rect 1356 4707 1363 4753
rect 1396 4747 1403 4773
rect 1396 4707 1403 4713
rect 1293 4693 1307 4707
rect 1233 4673 1247 4687
rect 1333 4693 1347 4707
rect 1353 4693 1367 4707
rect 1393 4693 1407 4707
rect 1253 4663 1267 4667
rect 1253 4656 1283 4663
rect 1253 4653 1267 4656
rect 1276 4627 1283 4656
rect 1236 4507 1243 4513
rect 1236 4487 1243 4493
rect 1276 4487 1283 4613
rect 1356 4587 1363 4653
rect 1376 4567 1383 4673
rect 1396 4507 1403 4653
rect 1416 4507 1423 4753
rect 1436 4687 1443 4733
rect 1556 4687 1563 4733
rect 1576 4727 1583 4993
rect 1596 4987 1603 5176
rect 1616 5007 1623 5333
rect 1676 5327 1683 5373
rect 1716 5307 1723 5433
rect 1816 5347 1823 5533
rect 1836 5447 1843 5453
rect 1856 5447 1863 5613
rect 1916 5607 1923 5873
rect 1936 5667 1943 5873
rect 1956 5863 1963 5893
rect 1976 5887 1983 6113
rect 1993 6093 2007 6107
rect 2013 6113 2027 6127
rect 2053 6113 2067 6127
rect 1996 6087 2003 6093
rect 2073 6073 2087 6087
rect 2076 6047 2083 6073
rect 2116 6047 2123 6136
rect 2136 6103 2143 6133
rect 2196 6127 2203 6133
rect 2236 6127 2243 6353
rect 2256 6307 2263 6373
rect 2276 6347 2283 6373
rect 2296 6367 2303 6373
rect 2316 6187 2323 6433
rect 2496 6427 2503 6433
rect 2493 6413 2507 6427
rect 2356 6387 2363 6393
rect 2353 6373 2367 6387
rect 2513 6403 2527 6407
rect 2513 6396 2543 6403
rect 2513 6393 2527 6396
rect 2373 6353 2387 6367
rect 2376 6347 2383 6353
rect 2136 6096 2163 6103
rect 2156 6083 2163 6096
rect 2193 6113 2207 6127
rect 2253 6123 2267 6127
rect 2253 6116 2283 6123
rect 2253 6113 2267 6116
rect 2213 6093 2227 6107
rect 2216 6083 2223 6093
rect 2156 6076 2183 6083
rect 1996 5927 2003 5933
rect 2016 5927 2023 5953
rect 2056 5927 2063 5933
rect 2013 5913 2027 5927
rect 2033 5893 2047 5907
rect 2053 5913 2067 5927
rect 2136 5923 2143 6073
rect 2136 5916 2163 5923
rect 1956 5856 1983 5863
rect 1956 5827 1963 5833
rect 1976 5667 1983 5856
rect 2036 5847 2043 5893
rect 2133 5873 2147 5887
rect 1996 5707 2003 5833
rect 1933 5653 1947 5667
rect 1996 5647 2003 5673
rect 2016 5647 2023 5653
rect 2013 5633 2027 5647
rect 1833 5433 1847 5447
rect 1876 5427 1883 5553
rect 1896 5447 1903 5453
rect 1916 5447 1923 5593
rect 1893 5433 1907 5447
rect 1956 5427 1963 5433
rect 1953 5413 1967 5427
rect 1973 5403 1987 5407
rect 1996 5403 2003 5473
rect 2036 5463 2043 5693
rect 2136 5687 2143 5873
rect 2096 5647 2103 5673
rect 2156 5663 2163 5916
rect 2176 5687 2183 6076
rect 2196 6076 2223 6083
rect 2196 6047 2203 6076
rect 2247 6076 2263 6083
rect 2196 5927 2203 5993
rect 2216 5947 2223 6053
rect 2236 5947 2243 5953
rect 2256 5947 2263 6076
rect 2276 6047 2283 6116
rect 2233 5933 2247 5947
rect 2193 5913 2207 5927
rect 2276 5927 2283 6033
rect 2296 5947 2303 6133
rect 2356 6127 2363 6333
rect 2416 6147 2423 6353
rect 2536 6327 2543 6396
rect 2576 6387 2583 6393
rect 2716 6387 2723 6413
rect 2896 6387 2903 6433
rect 3096 6423 3103 6453
rect 3196 6436 3243 6443
rect 3016 6416 3103 6423
rect 2573 6373 2587 6387
rect 2593 6353 2607 6367
rect 2333 6093 2347 6107
rect 2353 6113 2367 6127
rect 2453 6133 2467 6147
rect 2433 6113 2447 6127
rect 2316 5943 2323 6093
rect 2336 5987 2343 6093
rect 2436 6067 2443 6113
rect 2316 5936 2343 5943
rect 2273 5913 2287 5927
rect 2336 5907 2343 5936
rect 2356 5927 2363 5953
rect 2236 5827 2243 5893
rect 2156 5656 2183 5663
rect 2136 5647 2143 5653
rect 2176 5647 2183 5656
rect 2073 5613 2087 5627
rect 2093 5633 2107 5647
rect 2133 5633 2147 5647
rect 2076 5567 2083 5613
rect 2113 5593 2127 5607
rect 2116 5587 2123 5593
rect 2216 5587 2223 5673
rect 2236 5667 2243 5813
rect 2276 5667 2283 5673
rect 2296 5667 2303 5893
rect 2376 5847 2383 5993
rect 2416 5907 2423 6053
rect 2456 5947 2463 6133
rect 2536 6127 2543 6173
rect 2596 6167 2603 6353
rect 2636 6307 2643 6373
rect 2653 6353 2667 6367
rect 2636 6127 2643 6293
rect 2656 6287 2663 6353
rect 2776 6347 2783 6353
rect 2796 6327 2803 6373
rect 2893 6373 2907 6387
rect 2933 6383 2947 6387
rect 2916 6376 2947 6383
rect 2696 6147 2703 6153
rect 2693 6133 2707 6147
rect 2573 6123 2587 6127
rect 2573 6116 2603 6123
rect 2573 6113 2587 6116
rect 2553 6073 2567 6087
rect 2556 5947 2563 6073
rect 2596 6067 2603 6116
rect 2713 6113 2727 6127
rect 2816 6127 2823 6133
rect 2856 6127 2863 6273
rect 2896 6167 2903 6333
rect 2916 6287 2923 6376
rect 2933 6373 2947 6376
rect 3016 6387 3023 6416
rect 3096 6407 3103 6416
rect 3036 6387 3043 6393
rect 3093 6393 3107 6407
rect 2956 6187 2963 6353
rect 2753 6113 2767 6127
rect 2653 6093 2667 6107
rect 2656 6087 2663 6093
rect 2716 6047 2723 6113
rect 2756 6107 2763 6113
rect 2813 6113 2827 6127
rect 2833 6093 2847 6107
rect 2853 6113 2867 6127
rect 2873 6103 2887 6107
rect 2896 6103 2903 6153
rect 2973 6133 2987 6147
rect 2873 6096 2903 6103
rect 2956 6107 2963 6113
rect 2873 6093 2887 6096
rect 2393 5873 2407 5887
rect 2413 5893 2427 5907
rect 2516 5887 2523 5933
rect 2533 5903 2547 5907
rect 2533 5896 2563 5903
rect 2533 5893 2547 5896
rect 2513 5873 2527 5887
rect 2396 5867 2403 5873
rect 2556 5867 2563 5896
rect 2633 5893 2647 5907
rect 2596 5883 2603 5893
rect 2576 5876 2603 5883
rect 2396 5847 2403 5853
rect 2253 5633 2267 5647
rect 2273 5653 2287 5667
rect 2356 5647 2363 5653
rect 2353 5633 2367 5647
rect 2256 5627 2263 5633
rect 2376 5623 2383 5713
rect 2576 5687 2583 5876
rect 2416 5647 2423 5673
rect 2393 5623 2407 5627
rect 2376 5616 2407 5623
rect 2413 5633 2427 5647
rect 2393 5613 2407 5616
rect 2216 5467 2223 5513
rect 2016 5456 2043 5463
rect 2016 5427 2023 5456
rect 2213 5453 2227 5467
rect 2076 5447 2083 5453
rect 1973 5396 2003 5403
rect 2013 5413 2027 5427
rect 2053 5413 2067 5427
rect 2073 5433 2087 5447
rect 2056 5403 2063 5413
rect 2093 5403 2107 5407
rect 2056 5396 2107 5403
rect 2156 5407 2163 5453
rect 2193 5413 2207 5427
rect 1973 5393 1987 5396
rect 1657 5198 1665 5222
rect 1657 5104 1665 5184
rect 1713 5133 1727 5147
rect 1676 5007 1683 5133
rect 1716 5127 1723 5133
rect 1656 4967 1663 4973
rect 1633 4933 1647 4947
rect 1653 4953 1667 4967
rect 1453 4673 1467 4687
rect 1456 4667 1463 4673
rect 1513 4653 1527 4667
rect 1436 4647 1443 4653
rect 1516 4627 1523 4653
rect 1573 4653 1587 4667
rect 1576 4627 1583 4653
rect 1193 4463 1207 4467
rect 1176 4456 1207 4463
rect 1233 4473 1247 4487
rect 1436 4487 1443 4493
rect 1193 4453 1207 4456
rect 1333 4453 1347 4467
rect 1336 4447 1343 4453
rect 1157 4238 1165 4262
rect 1276 4227 1283 4253
rect 1016 4187 1023 4193
rect 1076 4007 1083 4033
rect 1116 4007 1123 4193
rect 1157 4144 1165 4224
rect 1213 4173 1227 4187
rect 1253 4173 1267 4187
rect 1216 4167 1223 4173
rect 1256 4127 1263 4173
rect 1296 4144 1304 4256
rect 1376 4243 1383 4473
rect 1433 4473 1447 4487
rect 1456 4427 1463 4473
rect 1496 4467 1503 4493
rect 1493 4453 1507 4467
rect 1533 4433 1547 4447
rect 1573 4433 1587 4447
rect 1536 4423 1543 4433
rect 1576 4427 1583 4433
rect 1487 4416 1543 4423
rect 1496 4327 1503 4416
rect 1376 4236 1403 4243
rect 1396 4227 1403 4236
rect 1256 4007 1263 4053
rect 1316 4047 1323 4213
rect 1393 4213 1407 4227
rect 1456 4207 1463 4313
rect 1453 4193 1467 4207
rect 1476 4187 1483 4213
rect 1556 4207 1563 4233
rect 1596 4207 1603 4893
rect 1616 4767 1623 4913
rect 1636 4707 1643 4933
rect 1676 4923 1683 4973
rect 1693 4923 1707 4927
rect 1676 4916 1707 4923
rect 1693 4913 1707 4916
rect 1733 4913 1747 4927
rect 1736 4907 1743 4913
rect 1676 4867 1683 4893
rect 1653 4653 1667 4667
rect 1656 4607 1663 4653
rect 1676 4623 1683 4793
rect 1696 4687 1703 4733
rect 1756 4703 1763 5113
rect 1796 5104 1804 5216
rect 1856 5143 1863 5373
rect 1936 5347 1943 5393
rect 2056 5367 2063 5396
rect 2093 5393 2107 5396
rect 2176 5347 2183 5413
rect 2196 5407 2203 5413
rect 2216 5367 2223 5393
rect 1896 5167 1903 5173
rect 1873 5143 1887 5147
rect 1856 5136 1887 5143
rect 1893 5153 1907 5167
rect 1873 5133 1887 5136
rect 2016 5147 2023 5173
rect 1973 5113 1987 5127
rect 1936 4987 1943 5113
rect 1956 4963 1963 4993
rect 1976 4987 1983 5113
rect 1996 4987 2003 5093
rect 2036 5027 2043 5173
rect 2196 5167 2203 5313
rect 2036 4967 2043 4993
rect 2116 4967 2123 5113
rect 2216 5047 2223 5333
rect 2236 5187 2243 5573
rect 2256 5427 2263 5513
rect 2276 5447 2283 5473
rect 2356 5467 2363 5473
rect 2353 5453 2367 5467
rect 2316 5447 2323 5453
rect 2273 5433 2287 5447
rect 2253 5413 2267 5427
rect 2313 5433 2327 5447
rect 2376 5447 2383 5453
rect 2296 5207 2303 5413
rect 2356 5367 2363 5413
rect 2396 5347 2403 5613
rect 2436 5467 2443 5673
rect 2596 5667 2603 5833
rect 2616 5707 2623 5893
rect 2636 5867 2643 5893
rect 2653 5873 2667 5887
rect 2716 5887 2723 5933
rect 2776 5907 2783 5933
rect 2796 5907 2803 6093
rect 2836 6087 2843 6093
rect 2816 5907 2823 5913
rect 2876 5907 2883 5933
rect 2896 5927 2903 6073
rect 2976 6067 2983 6133
rect 2993 6113 3007 6127
rect 3076 6143 3083 6373
rect 3116 6307 3123 6433
rect 3153 6423 3167 6427
rect 3176 6423 3183 6433
rect 3196 6427 3203 6436
rect 3236 6427 3243 6436
rect 3256 6427 3263 6433
rect 3153 6416 3183 6423
rect 3153 6413 3167 6416
rect 3156 6347 3163 6373
rect 3176 6287 3183 6416
rect 3253 6413 3267 6427
rect 3193 6373 3207 6387
rect 3376 6407 3383 6413
rect 3233 6383 3247 6387
rect 3233 6376 3263 6383
rect 3233 6373 3247 6376
rect 3196 6367 3203 6373
rect 3076 6136 3103 6143
rect 3096 6127 3103 6136
rect 3116 6127 3123 6253
rect 3136 6127 3143 6193
rect 3236 6167 3243 6273
rect 3256 6267 3263 6376
rect 3373 6393 3387 6407
rect 3396 6387 3403 6433
rect 3456 6407 3463 6453
rect 3736 6436 3783 6443
rect 3453 6393 3467 6407
rect 3393 6373 3407 6387
rect 3473 6373 3487 6387
rect 3276 6207 3283 6373
rect 3476 6327 3483 6373
rect 3176 6147 3183 6153
rect 3173 6133 3187 6147
rect 2916 5907 2923 5913
rect 2656 5867 2663 5873
rect 2736 5707 2743 5893
rect 2773 5893 2787 5907
rect 2813 5893 2827 5907
rect 2873 5893 2887 5907
rect 2913 5893 2927 5907
rect 2676 5687 2683 5693
rect 2816 5667 2823 5693
rect 2513 5663 2527 5667
rect 2496 5656 2527 5663
rect 2553 5663 2567 5667
rect 2453 5613 2467 5627
rect 2456 5507 2463 5613
rect 2447 5456 2453 5463
rect 2476 5463 2483 5533
rect 2496 5527 2503 5656
rect 2513 5653 2527 5656
rect 2533 5633 2547 5647
rect 2553 5656 2583 5663
rect 2553 5653 2567 5656
rect 2536 5623 2543 5633
rect 2576 5627 2583 5656
rect 2593 5653 2607 5667
rect 2633 5653 2647 5667
rect 2693 5663 2707 5667
rect 2613 5633 2627 5647
rect 2536 5616 2563 5623
rect 2556 5607 2563 5616
rect 2616 5607 2623 5633
rect 2536 5467 2543 5533
rect 2476 5456 2503 5463
rect 2496 5447 2503 5456
rect 2596 5463 2603 5533
rect 2636 5527 2643 5653
rect 2653 5643 2667 5647
rect 2676 5656 2707 5663
rect 2676 5643 2683 5656
rect 2653 5636 2683 5643
rect 2693 5653 2707 5656
rect 2733 5653 2747 5667
rect 2653 5633 2667 5636
rect 2713 5633 2727 5647
rect 2656 5627 2663 5633
rect 2716 5623 2723 5633
rect 2736 5627 2743 5653
rect 2793 5633 2807 5647
rect 2813 5653 2827 5667
rect 2696 5616 2723 5623
rect 2676 5607 2683 5613
rect 2433 5413 2447 5427
rect 2493 5433 2507 5447
rect 2576 5456 2603 5463
rect 2576 5447 2583 5456
rect 2616 5447 2623 5473
rect 2513 5413 2527 5427
rect 2573 5433 2587 5447
rect 2613 5433 2627 5447
rect 2636 5427 2643 5433
rect 2633 5413 2647 5427
rect 2436 5203 2443 5413
rect 2516 5387 2523 5413
rect 2656 5387 2663 5473
rect 2696 5427 2703 5616
rect 2673 5393 2687 5407
rect 2693 5413 2707 5427
rect 2396 5196 2443 5203
rect 2256 5143 2263 5193
rect 2376 5187 2383 5193
rect 2333 5183 2347 5187
rect 2316 5176 2347 5183
rect 2273 5143 2287 5147
rect 2256 5136 2287 5143
rect 2273 5133 2287 5136
rect 2293 5123 2307 5127
rect 2316 5123 2323 5176
rect 2333 5173 2347 5176
rect 2353 5153 2367 5167
rect 2373 5173 2387 5187
rect 2396 5167 2403 5196
rect 2453 5173 2467 5187
rect 2456 5167 2463 5173
rect 2496 5167 2503 5173
rect 2596 5167 2603 5173
rect 2433 5153 2447 5167
rect 2473 5163 2487 5167
rect 2473 5156 2493 5163
rect 2473 5153 2487 5156
rect 2356 5147 2363 5153
rect 2436 5147 2443 5153
rect 2513 5143 2527 5147
rect 2507 5136 2527 5143
rect 2513 5133 2527 5136
rect 2276 5116 2323 5123
rect 1973 4963 1987 4967
rect 1956 4956 1987 4963
rect 1973 4953 1987 4956
rect 1853 4913 1867 4927
rect 1916 4927 1923 4933
rect 1736 4696 1763 4703
rect 1796 4703 1803 4913
rect 1856 4807 1863 4913
rect 1896 4847 1903 4893
rect 1796 4696 1813 4703
rect 1676 4616 1703 4623
rect 1616 4247 1623 4493
rect 1656 4487 1663 4513
rect 1696 4487 1703 4616
rect 1736 4507 1743 4696
rect 1793 4653 1807 4667
rect 1796 4647 1803 4653
rect 1816 4647 1823 4673
rect 1893 4673 1907 4687
rect 1773 4633 1787 4647
rect 1896 4643 1903 4673
rect 1876 4636 1903 4643
rect 1653 4473 1667 4487
rect 1693 4473 1707 4487
rect 1756 4267 1763 4633
rect 1776 4627 1783 4633
rect 1776 4404 1784 4516
rect 1816 4487 1823 4613
rect 1876 4567 1883 4636
rect 1916 4563 1923 4893
rect 1936 4827 1943 4953
rect 2053 4943 2067 4947
rect 2036 4936 2067 4943
rect 1936 4687 1943 4713
rect 1956 4667 1963 4873
rect 1976 4867 1983 4913
rect 1977 4718 1985 4742
rect 1953 4653 1967 4667
rect 1977 4624 1985 4704
rect 1896 4556 1923 4563
rect 1813 4473 1827 4487
rect 1636 4207 1643 4213
rect 1656 4207 1663 4233
rect 1676 4227 1683 4253
rect 1676 4207 1683 4213
rect 1553 4193 1567 4207
rect 1573 4173 1587 4187
rect 1613 4173 1627 4187
rect 1633 4193 1647 4207
rect 1673 4193 1687 4207
rect 1433 4163 1447 4167
rect 1416 4156 1447 4163
rect 1253 3993 1267 4007
rect 1073 3953 1087 3967
rect 1113 3953 1127 3967
rect 1076 3947 1083 3953
rect 1016 3664 1024 3776
rect 1056 3647 1063 3933
rect 1116 3827 1123 3953
rect 1136 3943 1143 3993
rect 1313 3973 1327 3987
rect 1316 3967 1323 3973
rect 1193 3953 1207 3967
rect 1377 3956 1385 4036
rect 1136 3936 1163 3943
rect 1076 3727 1083 3813
rect 1116 3727 1123 3733
rect 1113 3713 1127 3727
rect 1156 3707 1163 3936
rect 1196 3767 1203 3953
rect 1377 3918 1385 3942
rect 1416 3907 1423 4156
rect 1433 4153 1447 4156
rect 1436 4007 1443 4013
rect 1433 3993 1447 4007
rect 1456 3763 1463 4033
rect 1473 4003 1487 4007
rect 1496 4003 1503 4173
rect 1473 3996 1503 4003
rect 1473 3993 1487 3996
rect 1516 3924 1524 4036
rect 1536 3947 1543 4153
rect 1576 4147 1583 4173
rect 1616 4127 1623 4173
rect 1696 4163 1703 4253
rect 1776 4227 1783 4233
rect 1733 4193 1747 4207
rect 1773 4213 1787 4227
rect 1676 4156 1703 4163
rect 1616 3987 1623 4073
rect 1656 4007 1663 4033
rect 1653 3993 1667 4007
rect 1613 3973 1627 3987
rect 1536 3883 1543 3933
rect 1516 3876 1543 3883
rect 1436 3756 1463 3763
rect 1196 3747 1203 3753
rect 1193 3733 1207 3747
rect 1133 3693 1147 3707
rect 1093 3673 1107 3687
rect 1096 3647 1103 3673
rect 1136 3647 1143 3693
rect 1156 3623 1163 3693
rect 1136 3616 1163 3623
rect 1036 3547 1043 3553
rect 1033 3533 1047 3547
rect 1116 3527 1123 3553
rect 1073 3523 1087 3527
rect 1013 3493 1027 3507
rect 1056 3516 1087 3523
rect 1016 3327 1023 3493
rect 1056 3447 1063 3516
rect 1073 3513 1087 3516
rect 1113 3513 1127 3527
rect 1136 3507 1143 3616
rect 1156 3527 1163 3573
rect 1176 3567 1183 3733
rect 1213 3713 1227 3727
rect 1216 3687 1223 3713
rect 1253 3693 1267 3707
rect 1316 3707 1323 3733
rect 1416 3727 1423 3733
rect 1293 3693 1307 3707
rect 1413 3713 1427 3727
rect 1256 3667 1263 3693
rect 1296 3687 1303 3693
rect 1176 3527 1183 3553
rect 1196 3527 1203 3533
rect 1153 3513 1167 3527
rect 1193 3513 1207 3527
rect 1257 3476 1265 3556
rect 1257 3438 1265 3462
rect 853 3243 867 3247
rect 836 3236 867 3243
rect 853 3233 867 3236
rect 893 3233 907 3247
rect 976 3223 983 3273
rect 1116 3263 1123 3313
rect 1096 3256 1123 3263
rect 993 3223 1007 3227
rect 976 3216 1007 3223
rect 1033 3223 1047 3227
rect 1056 3223 1063 3253
rect 1096 3247 1103 3256
rect 976 3207 983 3216
rect 993 3213 1007 3216
rect 1033 3216 1063 3223
rect 1033 3213 1047 3216
rect 1093 3233 1107 3247
rect 1133 3243 1147 3247
rect 1156 3243 1163 3353
rect 1133 3236 1163 3243
rect 1133 3233 1147 3236
rect 1113 3223 1127 3227
rect 1113 3216 1153 3223
rect 1113 3213 1127 3216
rect 1173 3213 1187 3227
rect 1013 3193 1027 3207
rect 796 3067 803 3173
rect 756 3056 783 3063
rect 776 3047 783 3056
rect 733 3033 747 3047
rect 773 3043 787 3047
rect 856 3043 863 3053
rect 896 3043 903 3193
rect 1016 3147 1023 3193
rect 1036 3167 1043 3213
rect 1176 3167 1183 3213
rect 976 3067 983 3073
rect 936 3043 943 3053
rect 716 3027 723 3033
rect 613 2993 627 3007
rect 633 3013 647 3027
rect 713 3013 727 3027
rect 753 3013 767 3027
rect 773 3036 803 3043
rect 773 3033 787 3036
rect 475 2958 483 2982
rect 616 2983 623 2993
rect 676 2987 683 3013
rect 616 2976 653 2983
rect 473 2733 487 2747
rect 476 2727 483 2733
rect 393 2723 407 2727
rect 376 2716 407 2723
rect 393 2713 407 2716
rect 493 2713 507 2727
rect 316 2656 343 2663
rect 276 2587 283 2593
rect 273 2563 287 2567
rect 273 2556 303 2563
rect 273 2553 287 2556
rect 296 2507 303 2556
rect 273 2263 287 2267
rect 296 2263 303 2293
rect 273 2256 303 2263
rect 313 2263 327 2267
rect 336 2263 343 2656
rect 356 2527 363 2553
rect 377 2516 385 2596
rect 436 2567 443 2573
rect 433 2563 447 2567
rect 456 2563 463 2713
rect 496 2687 503 2713
rect 433 2556 463 2563
rect 433 2553 447 2556
rect 377 2478 385 2502
rect 516 2484 524 2596
rect 556 2507 563 2773
rect 576 2704 584 2816
rect 596 2787 603 2973
rect 696 2967 703 2993
rect 756 2967 763 3013
rect 796 3007 803 3036
rect 836 3036 863 3043
rect 876 3036 903 3043
rect 916 3036 943 3043
rect 836 3027 843 3036
rect 813 2993 827 3007
rect 833 3013 847 3027
rect 853 2993 867 3007
rect 816 2987 823 2993
rect 856 2987 863 2993
rect 876 2983 883 3036
rect 916 3027 923 3036
rect 913 3013 927 3027
rect 953 3013 967 3027
rect 933 2993 947 3007
rect 876 2976 903 2983
rect 616 2827 623 2953
rect 715 2798 723 2822
rect 796 2807 803 2973
rect 856 2947 863 2973
rect 816 2807 823 2813
rect 896 2803 903 2976
rect 936 2807 943 2993
rect 956 2967 963 3013
rect 1036 3003 1043 3073
rect 1073 3033 1087 3047
rect 1016 2996 1043 3003
rect 956 2807 963 2953
rect 896 2796 923 2803
rect 613 2733 627 2747
rect 653 2733 667 2747
rect 616 2687 623 2733
rect 656 2727 663 2733
rect 715 2704 723 2784
rect 736 2747 743 2753
rect 733 2733 747 2747
rect 636 2587 643 2593
rect 633 2573 647 2587
rect 613 2533 627 2547
rect 616 2347 623 2533
rect 713 2513 727 2527
rect 716 2507 723 2513
rect 756 2347 763 2793
rect 793 2743 807 2747
rect 816 2743 823 2793
rect 856 2767 863 2793
rect 896 2767 903 2773
rect 793 2736 823 2743
rect 793 2733 807 2736
rect 853 2753 867 2767
rect 893 2753 907 2767
rect 916 2747 923 2796
rect 936 2787 943 2793
rect 933 2773 947 2787
rect 953 2753 967 2767
rect 956 2607 963 2753
rect 813 2523 827 2527
rect 836 2523 843 2593
rect 853 2533 867 2547
rect 976 2543 983 2633
rect 996 2607 1003 2833
rect 1016 2787 1023 2996
rect 1076 2987 1083 3033
rect 1097 2996 1105 3076
rect 1156 3047 1163 3053
rect 1153 3043 1167 3047
rect 1136 3036 1167 3043
rect 1097 2958 1105 2982
rect 1056 2787 1063 2793
rect 1013 2773 1027 2787
rect 1053 2773 1067 2787
rect 1096 2767 1103 2793
rect 1016 2567 1023 2733
rect 1076 2723 1083 2733
rect 1093 2723 1107 2727
rect 1076 2716 1107 2723
rect 1093 2713 1107 2716
rect 1136 2707 1143 3036
rect 1153 3033 1167 3036
rect 1236 2964 1244 3076
rect 1216 2767 1223 2813
rect 1213 2753 1227 2767
rect 993 2543 1007 2547
rect 976 2536 1007 2543
rect 993 2533 1007 2536
rect 856 2527 863 2533
rect 1036 2527 1043 2573
rect 813 2516 843 2523
rect 813 2513 827 2516
rect 1077 2516 1085 2596
rect 1136 2587 1143 2693
rect 1136 2567 1143 2573
rect 1133 2553 1147 2567
rect 1156 2523 1163 2673
rect 1136 2516 1163 2523
rect 376 2307 383 2333
rect 527 2296 563 2303
rect 376 2287 383 2293
rect 416 2287 423 2293
rect 556 2287 563 2296
rect 616 2287 623 2333
rect 957 2318 965 2342
rect 673 2303 687 2307
rect 673 2296 703 2303
rect 673 2293 687 2296
rect 313 2256 343 2263
rect 273 2253 287 2256
rect 313 2253 327 2256
rect 353 2253 367 2267
rect 373 2273 387 2287
rect 316 2147 323 2253
rect 276 2107 283 2133
rect 256 2076 283 2083
rect 253 2063 267 2067
rect 236 2056 267 2063
rect 253 2053 267 2056
rect 117 1838 125 1862
rect 33 1793 47 1807
rect 93 1783 107 1787
rect 53 1763 67 1767
rect 76 1776 107 1783
rect 76 1763 83 1776
rect 53 1756 83 1763
rect 93 1773 107 1776
rect 53 1753 67 1756
rect 117 1744 125 1824
rect 173 1773 187 1787
rect 176 1743 183 1773
rect 196 1767 203 2013
rect 256 1903 263 1993
rect 236 1896 263 1903
rect 156 1736 183 1743
rect 16 1347 23 1613
rect 96 1587 103 1613
rect 156 1587 163 1736
rect 196 1627 203 1753
rect 156 1567 163 1573
rect 176 1447 183 1593
rect 196 1423 203 1613
rect 176 1416 203 1423
rect 176 1347 183 1416
rect 236 1367 243 1896
rect 256 1744 264 1856
rect 253 1583 267 1587
rect 276 1583 283 2076
rect 316 2067 323 2093
rect 356 2087 363 2253
rect 553 2273 567 2287
rect 593 2273 607 2287
rect 573 2253 587 2267
rect 433 2233 447 2247
rect 396 2123 403 2133
rect 387 2116 403 2123
rect 336 2076 353 2083
rect 293 2033 307 2047
rect 313 2053 327 2067
rect 336 2047 343 2076
rect 296 1987 303 2033
rect 376 1967 383 2093
rect 396 2083 403 2116
rect 436 2083 443 2233
rect 476 2223 483 2233
rect 516 2223 523 2233
rect 476 2216 523 2223
rect 496 2123 503 2133
rect 496 2116 513 2123
rect 396 2076 423 2083
rect 436 2076 463 2083
rect 416 2067 423 2076
rect 456 2067 463 2076
rect 413 2053 427 2067
rect 476 2047 483 2113
rect 496 2067 503 2073
rect 493 2053 507 2067
rect 473 2033 487 2047
rect 396 2007 403 2033
rect 313 1773 327 1787
rect 316 1767 323 1773
rect 353 1773 367 1787
rect 396 1783 403 1893
rect 436 1807 443 2033
rect 496 1827 503 1953
rect 556 1843 563 2213
rect 576 2167 583 2253
rect 596 2187 603 2273
rect 653 2253 667 2267
rect 696 2263 703 2296
rect 753 2293 767 2307
rect 676 2256 703 2263
rect 733 2273 747 2287
rect 736 2267 743 2273
rect 656 2247 663 2253
rect 576 2127 583 2133
rect 576 2087 583 2093
rect 573 2073 587 2087
rect 676 2087 683 2256
rect 713 2253 727 2267
rect 716 2247 723 2253
rect 756 2227 763 2293
rect 833 2303 847 2307
rect 816 2296 847 2303
rect 873 2303 887 2307
rect 816 2267 823 2296
rect 833 2293 847 2296
rect 853 2273 867 2287
rect 873 2296 903 2303
rect 873 2293 887 2296
rect 673 2073 687 2087
rect 696 2067 703 2173
rect 693 2053 707 2067
rect 596 1967 603 2053
rect 616 1947 623 2033
rect 536 1836 563 1843
rect 496 1807 503 1813
rect 413 1783 427 1787
rect 396 1776 427 1783
rect 413 1773 427 1776
rect 356 1667 363 1773
rect 493 1793 507 1807
rect 536 1803 543 1836
rect 677 1838 685 1862
rect 596 1807 603 1813
rect 553 1803 567 1807
rect 536 1796 567 1803
rect 433 1753 447 1767
rect 513 1763 527 1767
rect 536 1763 543 1796
rect 553 1793 567 1796
rect 573 1773 587 1787
rect 593 1793 607 1807
rect 613 1783 627 1787
rect 636 1783 643 1833
rect 716 1827 723 2153
rect 736 2067 743 2133
rect 756 2047 763 2093
rect 816 2087 823 2233
rect 836 2127 843 2253
rect 856 2187 863 2273
rect 836 2087 843 2113
rect 833 2073 847 2087
rect 753 2033 767 2047
rect 816 2023 823 2053
rect 796 2016 823 2023
rect 656 1787 663 1793
rect 613 1776 643 1783
rect 613 1773 627 1776
rect 653 1773 667 1787
rect 513 1756 543 1763
rect 513 1753 527 1756
rect 253 1576 283 1583
rect 253 1573 267 1576
rect 276 1387 283 1576
rect 336 1524 344 1636
rect 376 1607 383 1713
rect 373 1593 387 1607
rect 413 1603 427 1607
rect 396 1596 427 1603
rect 396 1567 403 1596
rect 413 1593 427 1596
rect 436 1527 443 1753
rect 456 1567 463 1753
rect 496 1647 503 1693
rect 475 1556 483 1636
rect 13 1293 27 1307
rect 73 1303 87 1307
rect 73 1296 103 1303
rect 73 1293 87 1296
rect 16 1287 23 1293
rect 33 1113 47 1127
rect 36 867 43 1113
rect 57 1076 65 1156
rect 57 1038 65 1062
rect 76 847 83 1273
rect 96 1127 103 1296
rect 113 1293 127 1307
rect 153 1303 167 1307
rect 176 1303 183 1333
rect 116 1287 123 1293
rect 153 1296 183 1303
rect 153 1293 167 1296
rect 116 1127 123 1133
rect 113 1113 127 1127
rect 176 1003 183 1296
rect 196 1247 203 1353
rect 256 1327 263 1353
rect 213 1313 227 1327
rect 216 1307 223 1313
rect 233 1293 247 1307
rect 253 1313 267 1327
rect 196 1044 204 1156
rect 236 1107 243 1293
rect 276 1283 283 1293
rect 256 1276 283 1283
rect 256 1103 263 1276
rect 296 1267 303 1353
rect 456 1343 463 1553
rect 475 1518 483 1542
rect 536 1367 543 1756
rect 576 1667 583 1773
rect 677 1744 685 1824
rect 733 1773 747 1787
rect 756 1783 763 1853
rect 776 1823 783 1973
rect 796 1847 803 2016
rect 836 1907 843 2033
rect 856 1887 863 2053
rect 896 2007 903 2296
rect 933 2263 947 2267
rect 916 2256 947 2263
rect 916 2087 923 2256
rect 933 2253 947 2256
rect 957 2224 965 2304
rect 976 2227 983 2453
rect 996 2287 1003 2513
rect 1077 2478 1085 2502
rect 996 2263 1003 2273
rect 1013 2263 1027 2267
rect 996 2256 1027 2263
rect 1013 2253 1027 2256
rect 1036 2087 1043 2333
rect 1053 2253 1067 2267
rect 1056 2107 1063 2253
rect 1096 2224 1104 2336
rect 916 2047 923 2073
rect 956 2067 963 2073
rect 933 2033 947 2047
rect 953 2053 967 2067
rect 993 2053 1007 2067
rect 1073 2083 1087 2087
rect 1073 2076 1103 2083
rect 1073 2073 1087 2076
rect 996 2043 1003 2053
rect 996 2036 1023 2043
rect 936 2007 943 2033
rect 976 1967 983 2033
rect 776 1816 803 1823
rect 773 1783 787 1787
rect 756 1776 787 1783
rect 773 1773 787 1776
rect 736 1767 743 1773
rect 596 1687 603 1713
rect 716 1627 723 1633
rect 713 1613 727 1627
rect 756 1607 763 1713
rect 693 1573 707 1587
rect 733 1573 747 1587
rect 753 1593 767 1607
rect 653 1563 667 1567
rect 696 1563 703 1573
rect 653 1556 703 1563
rect 653 1553 667 1556
rect 547 1356 563 1363
rect 556 1347 563 1356
rect 456 1336 483 1343
rect 353 1293 367 1307
rect 356 1287 363 1293
rect 416 1307 423 1333
rect 476 1287 483 1336
rect 553 1333 567 1347
rect 333 1273 347 1287
rect 433 1273 447 1287
rect 593 1273 607 1287
rect 296 1147 303 1153
rect 293 1133 307 1147
rect 273 1103 287 1107
rect 256 1096 287 1103
rect 273 1093 287 1096
rect 176 996 203 1003
rect 73 843 87 847
rect 56 836 87 843
rect 13 793 27 807
rect 16 687 23 793
rect 56 667 63 836
rect 73 833 87 836
rect 33 613 47 627
rect 16 343 23 613
rect 36 607 43 613
rect 56 467 63 633
rect 96 627 103 693
rect 116 647 123 893
rect 136 867 143 873
rect 133 853 147 867
rect 153 833 167 847
rect 156 663 163 833
rect 196 687 203 996
rect 237 878 245 902
rect 316 887 323 1273
rect 336 1247 343 1273
rect 356 1263 363 1273
rect 396 1263 403 1273
rect 356 1256 403 1263
rect 436 1247 443 1273
rect 357 1076 365 1156
rect 376 1127 383 1153
rect 357 1038 365 1062
rect 216 827 223 833
rect 213 813 227 827
rect 237 784 245 864
rect 293 813 307 827
rect 296 807 303 813
rect 376 784 384 896
rect 136 656 163 663
rect 136 627 143 656
rect 216 647 223 773
rect 396 747 403 1153
rect 416 1127 423 1133
rect 413 1113 427 1127
rect 436 907 443 1233
rect 476 1147 483 1273
rect 596 1267 603 1273
rect 456 847 463 873
rect 476 847 483 1133
rect 496 1044 504 1156
rect 553 1143 567 1147
rect 536 1136 567 1143
rect 536 887 543 1136
rect 553 1133 567 1136
rect 616 1107 623 1173
rect 636 1127 643 1253
rect 656 1247 663 1513
rect 716 1264 724 1376
rect 736 1327 743 1573
rect 776 1347 783 1553
rect 796 1407 803 1816
rect 816 1744 824 1856
rect 836 1683 843 1853
rect 876 1763 883 1913
rect 996 1827 1003 1993
rect 1016 1947 1023 2036
rect 1096 1967 1103 2076
rect 1116 1987 1123 2113
rect 1016 1907 1023 1933
rect 913 1793 927 1807
rect 916 1767 923 1793
rect 876 1756 903 1763
rect 816 1676 843 1683
rect 776 1267 783 1333
rect 793 1293 807 1307
rect 796 1287 803 1293
rect 716 1127 723 1153
rect 736 1147 743 1253
rect 816 1187 823 1676
rect 836 1524 844 1636
rect 876 1607 883 1733
rect 873 1593 887 1607
rect 855 1358 863 1382
rect 855 1264 863 1344
rect 876 1307 883 1353
rect 896 1307 903 1756
rect 956 1707 963 1793
rect 973 1783 987 1787
rect 996 1783 1003 1813
rect 973 1776 1003 1783
rect 973 1773 987 1776
rect 1056 1763 1063 1953
rect 1136 1827 1143 2516
rect 1176 2287 1183 2373
rect 1173 2273 1187 2287
rect 1153 2233 1167 2247
rect 1196 2243 1203 2713
rect 1216 2484 1224 2596
rect 1176 2236 1203 2243
rect 1156 2187 1163 2233
rect 1156 2004 1164 2116
rect 1176 2047 1183 2236
rect 1236 2103 1243 2593
rect 1256 2387 1263 3313
rect 1276 3267 1283 3293
rect 1296 3283 1303 3573
rect 1336 3567 1343 3653
rect 1313 3523 1327 3527
rect 1353 3523 1367 3527
rect 1376 3523 1383 3553
rect 1313 3516 1343 3523
rect 1313 3513 1327 3516
rect 1336 3507 1343 3516
rect 1353 3516 1383 3523
rect 1353 3513 1367 3516
rect 1396 3444 1404 3556
rect 1436 3547 1443 3756
rect 1496 3747 1503 3753
rect 1516 3747 1523 3876
rect 1473 3713 1487 3727
rect 1493 3733 1507 3747
rect 1553 3743 1567 3747
rect 1553 3736 1583 3743
rect 1553 3733 1567 3736
rect 1476 3607 1483 3713
rect 1536 3687 1543 3713
rect 1576 3667 1583 3736
rect 1676 3723 1683 4156
rect 1696 4007 1703 4133
rect 1736 4127 1743 4193
rect 1796 4187 1803 4193
rect 1756 4027 1763 4153
rect 1836 4047 1843 4513
rect 1856 4487 1863 4493
rect 1896 4487 1903 4556
rect 1853 4473 1867 4487
rect 1856 4083 1863 4433
rect 1896 4303 1903 4473
rect 1915 4436 1923 4516
rect 1956 4447 1963 4473
rect 1996 4467 2003 4833
rect 2036 4827 2043 4936
rect 2053 4933 2067 4936
rect 2113 4953 2127 4967
rect 2136 4947 2143 5033
rect 2156 4967 2163 4973
rect 2216 4967 2223 4993
rect 2236 4987 2243 4993
rect 2276 4987 2283 5116
rect 2293 5113 2307 5116
rect 2336 4987 2343 5013
rect 2233 4973 2247 4987
rect 2333 4973 2347 4987
rect 2153 4953 2167 4967
rect 2213 4953 2227 4967
rect 2313 4963 2327 4967
rect 2173 4923 2187 4927
rect 2196 4923 2203 4953
rect 2253 4933 2267 4947
rect 2296 4956 2327 4963
rect 2356 4967 2363 4973
rect 2256 4927 2263 4933
rect 2296 4927 2303 4956
rect 2313 4953 2327 4956
rect 2353 4953 2367 4967
rect 2376 4943 2383 4993
rect 2456 4987 2463 5073
rect 2453 4973 2467 4987
rect 2416 4947 2423 4973
rect 2496 4963 2503 5133
rect 2593 5153 2607 5167
rect 2533 5113 2547 5127
rect 2616 5127 2623 5233
rect 2636 5143 2643 5353
rect 2676 5307 2683 5393
rect 2676 5187 2683 5293
rect 2736 5247 2743 5493
rect 2756 5403 2763 5513
rect 2796 5427 2803 5633
rect 2836 5627 2843 5693
rect 2876 5647 2883 5713
rect 2853 5613 2867 5627
rect 2873 5633 2887 5647
rect 2913 5643 2927 5647
rect 2936 5643 2943 5993
rect 2956 5967 2963 6053
rect 2996 5967 3003 6113
rect 3073 6093 3087 6107
rect 3093 6113 3107 6127
rect 3133 6113 3147 6127
rect 3233 6123 3247 6127
rect 3256 6123 3263 6193
rect 3436 6147 3443 6273
rect 3496 6167 3503 6313
rect 3516 6187 3523 6373
rect 3536 6347 3543 6413
rect 3573 6373 3587 6387
rect 3636 6387 3643 6393
rect 3633 6373 3647 6387
rect 3576 6367 3583 6373
rect 3693 6363 3707 6367
rect 3716 6363 3723 6413
rect 3736 6407 3743 6436
rect 3776 6423 3783 6436
rect 3933 6423 3947 6427
rect 3776 6416 3883 6423
rect 3756 6387 3763 6413
rect 3876 6407 3883 6416
rect 3916 6416 3947 6423
rect 3693 6356 3723 6363
rect 3793 6373 3807 6387
rect 3853 6373 3867 6387
rect 3873 6393 3887 6407
rect 3893 6383 3907 6387
rect 3916 6383 3923 6416
rect 3933 6413 3947 6416
rect 3893 6376 3923 6383
rect 3893 6373 3907 6376
rect 3693 6353 3707 6356
rect 3596 6347 3603 6353
rect 3516 6167 3523 6173
rect 3596 6167 3603 6333
rect 3776 6267 3783 6353
rect 3796 6347 3803 6373
rect 3796 6243 3803 6333
rect 3776 6236 3803 6243
rect 3433 6133 3447 6147
rect 3296 6127 3303 6133
rect 3376 6127 3383 6133
rect 3233 6116 3263 6123
rect 3233 6113 3247 6116
rect 2976 5907 2983 5953
rect 3016 5927 3023 6073
rect 3036 5927 3043 6053
rect 3076 6047 3083 6093
rect 3273 6093 3287 6107
rect 3293 6113 3307 6127
rect 3276 6083 3283 6093
rect 3256 6076 3283 6083
rect 3373 6113 3387 6127
rect 3576 6147 3583 6153
rect 3453 6113 3467 6127
rect 3533 6133 3547 6147
rect 3513 6113 3527 6127
rect 3136 5963 3143 6053
rect 3136 5956 3203 5963
rect 3136 5936 3183 5943
rect 3096 5927 3103 5933
rect 3016 5907 3023 5913
rect 3076 5907 3083 5913
rect 3116 5907 3123 5933
rect 3136 5927 3143 5936
rect 3176 5927 3183 5936
rect 3196 5923 3203 5956
rect 3196 5916 3223 5923
rect 2973 5893 2987 5907
rect 3013 5903 3027 5907
rect 3013 5896 3043 5903
rect 3013 5893 3027 5896
rect 2996 5887 3003 5893
rect 2993 5873 3007 5887
rect 3036 5847 3043 5896
rect 3053 5873 3067 5887
rect 3073 5893 3087 5907
rect 3113 5893 3127 5907
rect 3156 5887 3163 5913
rect 3056 5867 3063 5873
rect 3193 5883 3207 5887
rect 3216 5883 3223 5916
rect 3256 5907 3263 6076
rect 3313 6073 3327 6087
rect 3456 6087 3463 6113
rect 3516 6107 3523 6113
rect 3393 6073 3407 6087
rect 3316 6067 3323 6073
rect 3396 6027 3403 6073
rect 3516 6003 3523 6073
rect 3536 6027 3543 6133
rect 3553 6113 3567 6127
rect 3573 6133 3587 6147
rect 3556 6067 3563 6113
rect 3596 6107 3603 6133
rect 3636 6127 3643 6133
rect 3716 6127 3723 6133
rect 3633 6113 3647 6127
rect 3713 6113 3727 6127
rect 3756 6087 3763 6133
rect 3776 6107 3783 6236
rect 3816 6167 3823 6353
rect 3856 6347 3863 6373
rect 3916 6327 3923 6376
rect 3953 6383 3967 6387
rect 3976 6383 3983 6413
rect 4096 6407 4103 6433
rect 4093 6393 4107 6407
rect 4153 6403 4167 6407
rect 3953 6376 3983 6383
rect 3953 6373 3967 6376
rect 3993 6353 4007 6367
rect 4136 6396 4167 6403
rect 4033 6363 4047 6367
rect 4033 6356 4063 6363
rect 4033 6353 4047 6356
rect 3836 6147 3843 6273
rect 3996 6267 4003 6353
rect 3896 6147 3903 6253
rect 4036 6147 4043 6333
rect 4056 6287 4063 6356
rect 4076 6307 4083 6373
rect 4136 6367 4143 6396
rect 4153 6393 4167 6396
rect 4336 6387 4343 6473
rect 4396 6387 4403 6493
rect 4436 6387 4443 6433
rect 4556 6427 4563 6433
rect 4553 6413 4567 6427
rect 4496 6387 4503 6393
rect 4113 6353 4127 6367
rect 4173 6353 4187 6367
rect 4273 6353 4287 6367
rect 4333 6373 4347 6387
rect 4393 6373 4407 6387
rect 4433 6373 4447 6387
rect 4493 6373 4507 6387
rect 4676 6407 4683 6453
rect 4756 6427 4763 6493
rect 4653 6373 4667 6387
rect 4673 6393 4687 6407
rect 4736 6376 4753 6383
rect 4576 6367 4583 6373
rect 4116 6347 4123 6353
rect 4176 6347 4183 6353
rect 4276 6267 4283 6353
rect 4556 6343 4563 6353
rect 4596 6343 4603 6353
rect 4556 6336 4603 6343
rect 4616 6327 4623 6373
rect 4636 6367 4643 6373
rect 4656 6367 4663 6373
rect 4716 6347 4723 6353
rect 3813 6113 3827 6127
rect 3833 6133 3847 6147
rect 3873 6113 3887 6127
rect 3893 6133 3907 6147
rect 4176 6127 4183 6193
rect 4336 6147 4343 6153
rect 3953 6113 3967 6127
rect 3693 6073 3707 6087
rect 3516 5996 3543 6003
rect 3376 5927 3383 5953
rect 3193 5876 3223 5883
rect 3373 5913 3387 5927
rect 3396 5907 3403 5933
rect 3193 5873 3207 5876
rect 2913 5636 2943 5643
rect 2913 5633 2927 5636
rect 2893 5613 2907 5627
rect 2856 5507 2863 5613
rect 2896 5467 2903 5613
rect 2956 5547 2963 5833
rect 3076 5707 3083 5853
rect 3176 5807 3183 5853
rect 3296 5847 3303 5893
rect 2976 5667 2983 5693
rect 3196 5683 3203 5833
rect 3156 5676 3203 5683
rect 2973 5653 2987 5667
rect 3013 5653 3027 5667
rect 3016 5607 3023 5653
rect 3056 5647 3063 5653
rect 3033 5633 3047 5647
rect 3036 5627 3043 5633
rect 3036 5567 3043 5613
rect 3156 5627 3163 5676
rect 3416 5667 3423 5933
rect 3473 5893 3487 5907
rect 3513 5893 3527 5907
rect 3476 5887 3483 5893
rect 3436 5667 3443 5793
rect 3516 5683 3523 5893
rect 3536 5867 3543 5996
rect 3556 5907 3563 6013
rect 3656 5927 3663 6073
rect 3696 6027 3703 6073
rect 3676 5947 3683 5973
rect 3753 5943 3767 5947
rect 3696 5936 3767 5943
rect 3553 5893 3567 5907
rect 3676 5907 3683 5933
rect 3696 5907 3703 5936
rect 3753 5933 3767 5936
rect 3716 5907 3723 5913
rect 3796 5927 3803 6093
rect 3333 5653 3347 5667
rect 3173 5633 3187 5647
rect 3176 5587 3183 5633
rect 3193 5613 3207 5627
rect 3233 5613 3247 5627
rect 3196 5607 3203 5613
rect 2956 5447 2963 5473
rect 2953 5433 2967 5447
rect 3016 5447 3023 5513
rect 3036 5463 3043 5533
rect 3036 5456 3083 5463
rect 3076 5447 3083 5456
rect 2993 5443 3007 5447
rect 3013 5443 3027 5447
rect 2773 5403 2787 5407
rect 2756 5396 2787 5403
rect 2793 5413 2807 5427
rect 2833 5423 2847 5427
rect 2833 5416 2863 5423
rect 2833 5413 2847 5416
rect 2816 5407 2823 5413
rect 2773 5393 2787 5396
rect 2856 5307 2863 5416
rect 2913 5393 2927 5407
rect 2653 5143 2667 5147
rect 2636 5136 2667 5143
rect 2696 5143 2703 5213
rect 2756 5167 2763 5193
rect 2713 5143 2727 5147
rect 2696 5136 2727 5143
rect 2653 5133 2667 5136
rect 2713 5133 2727 5136
rect 2773 5133 2787 5147
rect 2776 5127 2783 5133
rect 2796 5127 2803 5213
rect 2916 5207 2923 5393
rect 2936 5307 2943 5433
rect 2993 5436 3027 5443
rect 2993 5433 3007 5436
rect 3013 5433 3027 5436
rect 3073 5423 3087 5427
rect 3073 5416 3103 5423
rect 3073 5413 3087 5416
rect 3036 5307 3043 5393
rect 3096 5383 3103 5416
rect 3116 5403 3123 5553
rect 3196 5467 3203 5473
rect 3236 5467 3243 5613
rect 3196 5447 3203 5453
rect 3193 5433 3207 5447
rect 3156 5427 3163 5433
rect 3133 5403 3147 5407
rect 3116 5396 3147 5403
rect 3153 5413 3167 5427
rect 3256 5427 3263 5633
rect 3336 5607 3343 5653
rect 3353 5633 3367 5647
rect 3433 5653 3447 5667
rect 3356 5627 3363 5633
rect 3293 5593 3307 5607
rect 3276 5447 3283 5593
rect 3296 5587 3303 5593
rect 3416 5547 3423 5653
rect 3516 5676 3543 5683
rect 3453 5643 3467 5647
rect 3453 5636 3483 5643
rect 3453 5633 3467 5636
rect 3476 5627 3483 5636
rect 3493 5633 3507 5647
rect 3496 5627 3503 5633
rect 3516 5627 3523 5676
rect 3536 5667 3543 5676
rect 3616 5667 3623 5873
rect 3636 5847 3643 5893
rect 3653 5873 3667 5887
rect 3673 5893 3687 5907
rect 3773 5893 3787 5907
rect 3793 5913 3807 5927
rect 3696 5887 3703 5893
rect 3693 5873 3707 5887
rect 3776 5887 3783 5893
rect 3656 5867 3663 5873
rect 3533 5653 3547 5667
rect 3573 5653 3587 5667
rect 3253 5413 3267 5427
rect 3356 5427 3363 5533
rect 3376 5447 3383 5473
rect 3373 5433 3387 5447
rect 3133 5393 3147 5396
rect 3173 5393 3187 5407
rect 3436 5447 3443 5473
rect 3433 5433 3447 5447
rect 3456 5427 3463 5613
rect 3576 5607 3583 5653
rect 3593 5633 3607 5647
rect 3596 5587 3603 5633
rect 3616 5627 3623 5653
rect 3636 5647 3643 5653
rect 3633 5633 3647 5647
rect 3676 5627 3683 5853
rect 3816 5827 3823 6113
rect 3836 5883 3843 6013
rect 3856 6007 3863 6093
rect 3876 6087 3883 6113
rect 3856 5927 3863 5953
rect 3853 5883 3867 5887
rect 3836 5876 3867 5883
rect 3896 5887 3903 5953
rect 3913 5903 3927 5907
rect 3936 5903 3943 6013
rect 3956 5967 3963 6113
rect 3973 6093 3987 6107
rect 4013 6103 4027 6107
rect 4033 6103 4047 6107
rect 4013 6096 4047 6103
rect 4093 6123 4107 6127
rect 4093 6116 4123 6123
rect 4093 6113 4107 6116
rect 4013 6093 4027 6096
rect 4033 6093 4047 6096
rect 4073 6093 4087 6107
rect 3976 5987 3983 6093
rect 3996 6047 4003 6073
rect 3956 5947 3963 5953
rect 3996 5947 4003 6013
rect 4016 5947 4023 6093
rect 3993 5933 4007 5947
rect 3913 5896 3943 5903
rect 3913 5893 3927 5896
rect 3853 5873 3867 5876
rect 3893 5873 3907 5887
rect 3936 5887 3943 5896
rect 4016 5887 4023 5893
rect 3956 5876 3973 5883
rect 3936 5847 3943 5873
rect 3956 5867 3963 5876
rect 3736 5647 3743 5653
rect 3693 5633 3707 5647
rect 3696 5607 3703 5633
rect 3733 5633 3747 5647
rect 3753 5623 3767 5627
rect 3776 5623 3783 5653
rect 3753 5616 3783 5623
rect 3753 5613 3767 5616
rect 3833 5623 3847 5627
rect 3853 5623 3867 5627
rect 3653 5593 3667 5607
rect 3476 5467 3483 5473
rect 3473 5453 3487 5467
rect 3576 5447 3583 5453
rect 3616 5447 3623 5593
rect 3656 5567 3663 5593
rect 3573 5443 3587 5447
rect 3507 5436 3523 5443
rect 3516 5407 3523 5436
rect 3556 5436 3587 5443
rect 3076 5376 3103 5383
rect 2833 5183 2847 5187
rect 2816 5176 2847 5183
rect 2536 5107 2543 5113
rect 2596 4967 2603 4993
rect 2636 4967 2643 4973
rect 2496 4956 2523 4963
rect 2393 4943 2407 4947
rect 2376 4936 2407 4943
rect 2393 4933 2407 4936
rect 2516 4947 2523 4956
rect 2593 4953 2607 4967
rect 2173 4916 2203 4923
rect 2173 4913 2187 4916
rect 2493 4913 2507 4927
rect 2513 4933 2527 4947
rect 2573 4943 2587 4947
rect 2533 4913 2547 4927
rect 2556 4936 2587 4943
rect 2496 4907 2503 4913
rect 2033 4653 2047 4667
rect 2036 4507 2043 4653
rect 2056 4527 2063 4873
rect 2496 4847 2503 4893
rect 2536 4887 2543 4913
rect 2556 4827 2563 4936
rect 2573 4933 2587 4936
rect 2613 4933 2627 4947
rect 2633 4953 2647 4967
rect 2676 4947 2683 5013
rect 2736 4967 2743 5093
rect 2816 5087 2823 5176
rect 2833 5173 2847 5176
rect 2853 5153 2867 5167
rect 2913 5183 2927 5187
rect 2896 5176 2927 5183
rect 2836 5107 2843 5133
rect 2856 5127 2863 5153
rect 2896 5067 2903 5176
rect 2913 5173 2927 5176
rect 3033 5163 3047 5167
rect 3033 5156 3063 5163
rect 3033 5153 3047 5156
rect 2996 5127 3003 5133
rect 3016 5127 3023 5153
rect 2973 5123 2987 5127
rect 2956 5116 2987 5123
rect 2956 5067 2963 5116
rect 2973 5113 2987 5116
rect 2733 4953 2747 4967
rect 2756 4947 2763 5053
rect 2796 4987 2803 4993
rect 2793 4973 2807 4987
rect 2816 4967 2823 4973
rect 2856 4967 2863 5053
rect 2936 4987 2943 4993
rect 2853 4953 2867 4967
rect 2616 4927 2623 4933
rect 2776 4927 2783 4933
rect 2896 4927 2903 4973
rect 2936 4947 2943 4973
rect 2956 4967 2963 5013
rect 2976 4987 2983 5093
rect 3056 5087 3063 5156
rect 3076 5143 3083 5376
rect 3176 5347 3183 5393
rect 3096 5187 3103 5273
rect 3136 5167 3143 5193
rect 3176 5187 3183 5213
rect 3093 5143 3107 5147
rect 3076 5136 3107 5143
rect 3093 5133 3107 5136
rect 3153 5143 3167 5147
rect 3236 5143 3243 5173
rect 3153 5136 3243 5143
rect 3153 5133 3167 5136
rect 3116 5047 3123 5133
rect 2996 4967 3003 5033
rect 2953 4953 2967 4967
rect 2933 4933 2947 4947
rect 2993 4953 3007 4967
rect 2916 4907 2923 4933
rect 3016 4907 3023 4953
rect 3036 4947 3043 4993
rect 3096 4967 3103 5033
rect 3033 4933 3047 4947
rect 3093 4953 3107 4967
rect 3116 4956 3133 4963
rect 3116 4947 3123 4956
rect 3176 4967 3183 4973
rect 3173 4953 3187 4967
rect 2927 4816 2943 4823
rect 2073 4663 2087 4667
rect 2096 4663 2103 4753
rect 2073 4656 2103 4663
rect 2073 4653 2087 4656
rect 2116 4624 2124 4736
rect 2236 4707 2243 4733
rect 2396 4707 2403 4713
rect 2233 4693 2247 4707
rect 2267 4696 2283 4703
rect 2276 4687 2283 4696
rect 2273 4673 2287 4687
rect 2296 4647 2303 4673
rect 2393 4693 2407 4707
rect 2416 4663 2423 4713
rect 2436 4707 2443 4733
rect 2717 4718 2725 4742
rect 2316 4627 2323 4653
rect 2376 4656 2423 4663
rect 2376 4647 2383 4656
rect 2433 4653 2447 4667
rect 2473 4663 2487 4667
rect 2496 4663 2503 4693
rect 2516 4687 2523 4713
rect 2556 4687 2563 4693
rect 2436 4587 2443 4653
rect 2473 4656 2503 4663
rect 2513 4673 2527 4687
rect 2553 4673 2567 4687
rect 2473 4653 2487 4656
rect 2456 4627 2463 4633
rect 1973 4443 1987 4447
rect 1967 4436 1987 4443
rect 1993 4453 2007 4467
rect 1973 4433 1987 4436
rect 2013 4433 2027 4447
rect 2097 4436 2105 4516
rect 2156 4487 2163 4493
rect 2153 4473 2167 4487
rect 1915 4398 1923 4422
rect 1896 4296 1923 4303
rect 1897 4238 1905 4262
rect 1876 4187 1883 4213
rect 1873 4173 1887 4187
rect 1897 4144 1905 4224
rect 1856 4076 1883 4083
rect 1693 3993 1707 4007
rect 1716 3823 1723 4013
rect 1833 3993 1847 4007
rect 1733 3953 1747 3967
rect 1836 3967 1843 3993
rect 1857 3956 1865 4036
rect 1736 3947 1743 3953
rect 1857 3918 1865 3942
rect 1716 3816 1743 3823
rect 1717 3758 1725 3782
rect 1593 3693 1607 3707
rect 1633 3703 1647 3707
rect 1656 3716 1683 3723
rect 1656 3703 1663 3716
rect 1693 3703 1707 3707
rect 1596 3647 1603 3693
rect 1633 3696 1663 3703
rect 1676 3696 1707 3703
rect 1633 3693 1647 3696
rect 1613 3673 1627 3687
rect 1496 3547 1503 3633
rect 1493 3533 1507 3547
rect 1473 3523 1487 3527
rect 1456 3516 1487 3523
rect 1296 3276 1323 3283
rect 1316 3267 1323 3276
rect 1273 3253 1287 3267
rect 1313 3263 1327 3267
rect 1313 3256 1343 3263
rect 1313 3253 1327 3256
rect 1336 3147 1343 3256
rect 1376 3227 1383 3293
rect 1397 3278 1405 3302
rect 1373 3213 1387 3227
rect 1397 3184 1405 3264
rect 1296 3107 1303 3133
rect 1296 3003 1303 3093
rect 1393 3033 1407 3047
rect 1336 3027 1343 3033
rect 1396 3027 1403 3033
rect 1313 3003 1327 3007
rect 1296 2996 1327 3003
rect 1333 3013 1347 3027
rect 1396 3007 1403 3013
rect 1313 2993 1327 2996
rect 1417 2996 1425 3076
rect 1316 2787 1323 2993
rect 1316 2767 1323 2773
rect 1336 2767 1343 2973
rect 1417 2958 1425 2982
rect 1276 2567 1283 2753
rect 1313 2753 1327 2767
rect 1376 2747 1383 2813
rect 1333 2713 1347 2727
rect 1336 2667 1343 2713
rect 1436 2603 1443 3513
rect 1456 3387 1463 3516
rect 1473 3513 1487 3516
rect 1577 3476 1585 3556
rect 1616 3527 1623 3673
rect 1676 3667 1683 3696
rect 1693 3693 1707 3696
rect 1717 3664 1725 3744
rect 1736 3707 1743 3816
rect 1836 3707 1843 3773
rect 1813 3703 1827 3707
rect 1796 3696 1827 3703
rect 1676 3647 1683 3653
rect 1636 3527 1643 3533
rect 1633 3513 1647 3527
rect 1453 3213 1467 3227
rect 1516 3227 1523 3473
rect 1577 3438 1585 3462
rect 1716 3444 1724 3556
rect 1736 3547 1743 3693
rect 1796 3627 1803 3696
rect 1813 3693 1827 3696
rect 1736 3507 1743 3533
rect 1816 3527 1823 3673
rect 1793 3523 1807 3527
rect 1776 3516 1807 3523
rect 1776 3483 1783 3516
rect 1793 3513 1807 3516
rect 1776 3476 1803 3483
rect 1456 3067 1463 3213
rect 1536 3184 1544 3296
rect 1633 3263 1647 3267
rect 1633 3256 1663 3263
rect 1633 3253 1647 3256
rect 1476 3047 1483 3053
rect 1516 3047 1523 3073
rect 1473 3033 1487 3047
rect 1513 3033 1527 3047
rect 1536 2803 1543 3053
rect 1556 2964 1564 3076
rect 1596 2807 1603 3233
rect 1656 3207 1663 3256
rect 1673 3223 1687 3227
rect 1696 3223 1703 3253
rect 1776 3247 1783 3293
rect 1673 3216 1703 3223
rect 1673 3213 1687 3216
rect 1713 3213 1727 3227
rect 1716 3207 1723 3213
rect 1796 3167 1803 3476
rect 1836 3287 1843 3673
rect 1856 3664 1864 3776
rect 1876 3687 1883 4076
rect 1916 4043 1923 4296
rect 1953 4173 1967 4187
rect 1956 4167 1963 4173
rect 2016 4147 2023 4433
rect 2097 4398 2105 4422
rect 2036 4144 2044 4256
rect 2133 4223 2147 4227
rect 2133 4216 2163 4223
rect 2133 4213 2147 4216
rect 2156 4147 2163 4216
rect 2176 4167 2183 4493
rect 2196 4487 2203 4513
rect 2193 4473 2207 4487
rect 2236 4404 2244 4516
rect 2296 4507 2303 4573
rect 2293 4493 2307 4507
rect 2356 4487 2363 4573
rect 2376 4507 2383 4573
rect 2476 4523 2483 4653
rect 2596 4647 2603 4673
rect 2693 4663 2707 4667
rect 2653 4643 2667 4647
rect 2676 4656 2707 4663
rect 2676 4643 2683 4656
rect 2653 4636 2683 4643
rect 2693 4653 2707 4656
rect 2653 4633 2667 4636
rect 2656 4607 2663 4633
rect 2717 4624 2725 4704
rect 2773 4653 2787 4667
rect 2456 4516 2483 4523
rect 2373 4493 2387 4507
rect 2353 4473 2367 4487
rect 2396 4487 2403 4513
rect 2456 4507 2463 4516
rect 2516 4507 2523 4513
rect 2453 4493 2467 4507
rect 2393 4473 2407 4487
rect 2513 4493 2527 4507
rect 2473 4483 2487 4487
rect 2473 4476 2503 4483
rect 2576 4483 2583 4513
rect 2593 4483 2607 4487
rect 2473 4473 2487 4476
rect 2496 4467 2503 4476
rect 2576 4476 2607 4483
rect 2593 4473 2607 4476
rect 2617 4436 2625 4516
rect 2716 4487 2723 4493
rect 2673 4483 2687 4487
rect 2673 4476 2703 4483
rect 2673 4473 2687 4476
rect 2696 4427 2703 4476
rect 2713 4473 2727 4487
rect 2617 4398 2625 4422
rect 2756 4404 2764 4516
rect 2776 4427 2783 4653
rect 2736 4267 2743 4313
rect 2253 4173 2267 4187
rect 2256 4147 2263 4173
rect 2316 4144 2324 4256
rect 2455 4238 2463 4262
rect 2393 4173 2407 4187
rect 2396 4167 2403 4173
rect 2455 4144 2463 4224
rect 2676 4207 2683 4253
rect 2796 4243 2803 4633
rect 2856 4624 2864 4736
rect 2936 4687 2943 4816
rect 3057 4718 3065 4742
rect 2896 4663 2903 4673
rect 2913 4663 2927 4667
rect 2896 4656 2927 4663
rect 2933 4673 2947 4687
rect 2973 4683 2987 4687
rect 2996 4683 3003 4713
rect 2973 4676 3003 4683
rect 2973 4673 2987 4676
rect 2913 4653 2927 4656
rect 3033 4663 3047 4667
rect 3016 4656 3047 4663
rect 3016 4623 3023 4656
rect 3033 4653 3047 4656
rect 3057 4624 3065 4704
rect 3016 4616 3043 4623
rect 2856 4487 2863 4493
rect 2833 4453 2847 4467
rect 2853 4473 2867 4487
rect 2836 4327 2843 4453
rect 2913 4433 2927 4447
rect 2953 4443 2967 4447
rect 2976 4443 2983 4533
rect 3036 4507 3043 4616
rect 3076 4607 3083 4933
rect 3196 4927 3203 5013
rect 3216 4967 3223 5093
rect 3256 4967 3263 5253
rect 3313 5173 3327 5187
rect 3316 5087 3323 5173
rect 3336 5067 3343 5153
rect 3356 5127 3363 5193
rect 3376 5167 3383 5173
rect 3373 5153 3387 5167
rect 3416 5123 3423 5353
rect 3456 5167 3463 5193
rect 3453 5153 3467 5167
rect 3416 5116 3443 5123
rect 3436 5107 3443 5116
rect 3473 5123 3487 5127
rect 3516 5123 3523 5233
rect 3536 5187 3543 5253
rect 3556 5167 3563 5436
rect 3573 5433 3587 5436
rect 3593 5413 3607 5427
rect 3613 5433 3627 5447
rect 3636 5427 3643 5473
rect 3656 5427 3663 5433
rect 3633 5413 3647 5427
rect 3596 5387 3603 5413
rect 3596 5187 3603 5373
rect 3656 5267 3663 5413
rect 3676 5327 3683 5533
rect 3716 5467 3723 5553
rect 3713 5453 3727 5467
rect 3736 5463 3743 5593
rect 3796 5547 3803 5613
rect 3833 5616 3867 5623
rect 3913 5643 3927 5647
rect 3936 5643 3943 5733
rect 3913 5636 3943 5643
rect 3913 5633 3927 5636
rect 3956 5627 3963 5853
rect 3976 5647 3983 5753
rect 3973 5633 3987 5647
rect 3833 5613 3847 5616
rect 3853 5613 3867 5616
rect 3813 5593 3827 5607
rect 3816 5587 3823 5593
rect 3836 5467 3843 5613
rect 3993 5593 4007 5607
rect 3996 5547 4003 5593
rect 3916 5467 3923 5513
rect 3736 5456 3803 5463
rect 3796 5447 3803 5456
rect 3913 5453 3927 5467
rect 3773 5413 3787 5427
rect 3793 5433 3807 5447
rect 3833 5443 3847 5447
rect 3856 5443 3863 5453
rect 3833 5436 3863 5443
rect 3833 5433 3847 5436
rect 3936 5447 3943 5533
rect 4016 5467 4023 5793
rect 4036 5687 4043 6073
rect 4056 5987 4063 6073
rect 4076 6067 4083 6093
rect 4096 6047 4103 6093
rect 4116 6087 4123 6116
rect 4153 6103 4167 6107
rect 4136 6096 4167 6103
rect 4076 5923 4083 5973
rect 4076 5916 4093 5923
rect 4116 5923 4123 6053
rect 4136 6027 4143 6096
rect 4153 6093 4167 6096
rect 4173 6073 4187 6087
rect 4256 6107 4263 6133
rect 4333 6133 4347 6147
rect 4376 6143 4383 6153
rect 4393 6143 4407 6147
rect 4376 6136 4407 6143
rect 4213 6073 4227 6087
rect 4156 5947 4163 6073
rect 4176 6047 4183 6073
rect 4216 6067 4223 6073
rect 4116 5916 4143 5923
rect 4053 5873 4067 5887
rect 4096 5887 4103 5893
rect 4093 5873 4107 5887
rect 4136 5887 4143 5916
rect 4173 5893 4187 5907
rect 4213 5893 4227 5907
rect 4176 5887 4183 5893
rect 4056 5827 4063 5873
rect 4056 5647 4063 5713
rect 4096 5647 4103 5753
rect 4116 5667 4123 5853
rect 4156 5707 4163 5773
rect 4033 5613 4047 5627
rect 4053 5633 4067 5647
rect 4073 5613 4087 5627
rect 4093 5633 4107 5647
rect 4113 5623 4127 5627
rect 4136 5623 4143 5693
rect 4196 5667 4203 5893
rect 4216 5807 4223 5893
rect 4256 5887 4263 5913
rect 4293 5873 4307 5887
rect 4236 5647 4243 5673
rect 4256 5667 4263 5773
rect 4276 5727 4283 5853
rect 4296 5847 4303 5873
rect 4316 5687 4323 6093
rect 4376 5927 4383 6136
rect 4393 6133 4407 6136
rect 4413 6093 4427 6107
rect 4416 6087 4423 6093
rect 4436 6067 4443 6193
rect 4456 6123 4463 6173
rect 4496 6147 4503 6313
rect 4516 6127 4523 6193
rect 4556 6167 4563 6193
rect 4473 6123 4487 6127
rect 4456 6116 4487 6123
rect 4473 6113 4487 6116
rect 4513 6113 4527 6127
rect 4533 6103 4547 6107
rect 4556 6103 4563 6153
rect 4596 6147 4603 6293
rect 4636 6127 4643 6213
rect 4716 6147 4723 6253
rect 4736 6167 4743 6376
rect 4796 6387 4803 6433
rect 4896 6407 4903 6493
rect 5456 6476 5503 6483
rect 4833 6373 4847 6387
rect 4876 6387 4883 6393
rect 4873 6373 4887 6387
rect 4836 6363 4843 6373
rect 4836 6356 4863 6363
rect 4856 6343 4863 6356
rect 4856 6336 4883 6343
rect 4876 6327 4883 6336
rect 4896 6287 4903 6373
rect 4916 6327 4923 6453
rect 4936 6387 4943 6433
rect 4956 6407 4963 6413
rect 5016 6407 5023 6453
rect 4953 6393 4967 6407
rect 4993 6403 5007 6407
rect 5013 6403 5027 6407
rect 4933 6373 4947 6387
rect 4973 6373 4987 6387
rect 4993 6396 5027 6403
rect 4993 6393 5007 6396
rect 5013 6393 5027 6396
rect 5033 6373 5047 6387
rect 5073 6383 5087 6387
rect 5073 6376 5103 6383
rect 5073 6373 5087 6376
rect 4976 6307 4983 6373
rect 4996 6327 5003 6353
rect 4673 6133 4687 6147
rect 4676 6127 4683 6133
rect 4533 6096 4563 6103
rect 4533 6093 4547 6096
rect 4633 6113 4647 6127
rect 4653 6113 4667 6127
rect 4693 6113 4707 6127
rect 4713 6133 4727 6147
rect 4656 6107 4663 6113
rect 4436 5927 4443 6013
rect 4456 5927 4463 5953
rect 4453 5913 4467 5927
rect 4333 5873 4347 5887
rect 4433 5903 4447 5907
rect 4416 5896 4447 5903
rect 4373 5873 4387 5887
rect 4336 5707 4343 5873
rect 4356 5787 4363 5853
rect 4376 5767 4383 5873
rect 4396 5807 4403 5893
rect 4416 5867 4423 5896
rect 4433 5893 4447 5896
rect 4533 5923 4547 5927
rect 4516 5916 4547 5923
rect 4573 5923 4587 5927
rect 4593 5923 4607 5927
rect 4456 5747 4463 5873
rect 4253 5653 4267 5667
rect 4153 5633 4167 5647
rect 4156 5627 4163 5633
rect 4113 5616 4143 5623
rect 4113 5613 4127 5616
rect 4273 5633 4287 5647
rect 4356 5647 4363 5653
rect 4313 5633 4327 5647
rect 4353 5633 4367 5647
rect 4213 5613 4227 5627
rect 4036 5607 4043 5613
rect 4036 5587 4043 5593
rect 4076 5567 4083 5613
rect 3956 5447 3963 5453
rect 3776 5387 3783 5413
rect 3616 5167 3623 5253
rect 3636 5187 3643 5233
rect 3473 5116 3523 5123
rect 3593 5143 3607 5147
rect 3587 5136 3607 5143
rect 3613 5153 3627 5167
rect 3633 5143 3647 5147
rect 3593 5133 3607 5136
rect 3633 5136 3653 5143
rect 3633 5133 3647 5136
rect 3473 5113 3487 5116
rect 3553 5113 3567 5127
rect 3316 5043 3323 5053
rect 3316 5036 3343 5043
rect 3276 4967 3283 5033
rect 3213 4953 3227 4967
rect 3233 4933 3247 4947
rect 3236 4927 3243 4933
rect 3336 4927 3343 5036
rect 3376 4967 3383 5073
rect 3416 4967 3423 4973
rect 3373 4953 3387 4967
rect 3413 4953 3427 4967
rect 3436 4947 3443 5033
rect 3313 4913 3327 4927
rect 3113 4653 3127 4667
rect 3033 4493 3047 4507
rect 3096 4487 3103 4653
rect 3116 4647 3123 4653
rect 3176 4543 3183 4913
rect 3196 4624 3204 4736
rect 3297 4718 3305 4742
rect 3316 4707 3323 4913
rect 3276 4667 3283 4693
rect 3273 4653 3287 4667
rect 3297 4624 3305 4704
rect 3353 4653 3367 4667
rect 3356 4647 3363 4653
rect 3156 4536 3183 4543
rect 3073 4453 3087 4467
rect 3093 4473 3107 4487
rect 3156 4483 3163 4536
rect 3173 4483 3187 4487
rect 3156 4476 3187 4483
rect 3173 4473 3187 4476
rect 3113 4463 3127 4467
rect 3113 4456 3143 4463
rect 3113 4453 3127 4456
rect 3016 4447 3023 4453
rect 2953 4436 2983 4443
rect 2953 4433 2967 4436
rect 2916 4327 2923 4433
rect 3076 4323 3083 4453
rect 3136 4407 3143 4456
rect 3197 4436 3205 4516
rect 3253 4483 3267 4487
rect 3253 4476 3283 4483
rect 3253 4473 3267 4476
rect 3276 4427 3283 4476
rect 3197 4398 3205 4422
rect 3067 4316 3083 4323
rect 2796 4236 2823 4243
rect 3177 4238 3185 4262
rect 2753 4223 2767 4227
rect 2613 4203 2627 4207
rect 2536 4147 2543 4173
rect 2573 4173 2587 4187
rect 2613 4196 2643 4203
rect 2613 4193 2627 4196
rect 2553 4153 2567 4167
rect 1896 4036 1923 4043
rect 1896 3747 1903 4036
rect 1916 4007 1923 4013
rect 1913 3993 1927 4007
rect 1996 3924 2004 4036
rect 2093 3963 2107 3967
rect 2116 3963 2123 4133
rect 2216 4007 2223 4133
rect 2556 4027 2563 4153
rect 2576 4087 2583 4173
rect 2636 4183 2643 4196
rect 2653 4183 2667 4187
rect 2636 4176 2667 4183
rect 2673 4193 2687 4207
rect 2713 4193 2727 4207
rect 2736 4216 2767 4223
rect 2716 4187 2723 4193
rect 2653 4173 2667 4176
rect 2693 4173 2707 4187
rect 2593 4153 2607 4167
rect 2596 4147 2603 4153
rect 2576 4027 2583 4033
rect 2433 4023 2447 4027
rect 2433 4016 2463 4023
rect 2433 4013 2447 4016
rect 2093 3956 2123 3963
rect 2213 3993 2227 4007
rect 2336 3987 2343 3993
rect 2093 3953 2107 3956
rect 2253 3953 2267 3967
rect 2293 3953 2307 3967
rect 2333 3973 2347 3987
rect 2353 3963 2367 3967
rect 2376 3963 2383 3993
rect 2353 3956 2383 3963
rect 2353 3953 2367 3956
rect 2256 3947 2263 3953
rect 2296 3847 2303 3953
rect 2456 3947 2463 4016
rect 2573 4013 2587 4027
rect 2556 4007 2563 4013
rect 2553 3993 2567 4007
rect 2596 4007 2603 4013
rect 2593 3993 2607 4007
rect 2616 3987 2623 4013
rect 1896 3707 1903 3733
rect 1876 3283 1883 3653
rect 1916 3607 1923 3753
rect 1976 3747 1983 3753
rect 1953 3713 1967 3727
rect 1973 3733 1987 3747
rect 1956 3587 1963 3713
rect 1993 3693 2007 3707
rect 2056 3707 2063 3833
rect 2147 3736 2163 3743
rect 2096 3727 2103 3733
rect 2156 3727 2163 3736
rect 2093 3713 2107 3727
rect 1996 3607 2003 3693
rect 2013 3673 2027 3687
rect 2153 3713 2167 3727
rect 2193 3723 2207 3727
rect 2236 3723 2243 3833
rect 2296 3787 2303 3833
rect 2376 3727 2383 3753
rect 2396 3727 2403 3773
rect 2416 3727 2423 3933
rect 2576 3727 2583 3793
rect 2616 3767 2623 3973
rect 2636 3847 2643 4033
rect 2656 4007 2663 4173
rect 2696 4167 2703 4173
rect 2736 4167 2743 4216
rect 2753 4213 2767 4216
rect 2816 4207 2823 4236
rect 2716 4027 2723 4073
rect 2653 3993 2667 4007
rect 2713 4013 2727 4027
rect 2253 3723 2267 3727
rect 2193 3716 2223 3723
rect 2236 3716 2267 3723
rect 2193 3713 2207 3716
rect 2173 3693 2187 3707
rect 2073 3673 2087 3687
rect 1916 3547 1923 3573
rect 1913 3533 1927 3547
rect 1936 3483 1943 3553
rect 1956 3507 1963 3573
rect 1976 3527 1983 3553
rect 2016 3527 2023 3673
rect 2076 3647 2083 3673
rect 2056 3547 2063 3553
rect 2053 3533 2067 3547
rect 1973 3513 1987 3527
rect 2013 3523 2027 3527
rect 2033 3523 2047 3527
rect 1916 3476 1943 3483
rect 1953 3493 1967 3507
rect 2013 3516 2047 3523
rect 2013 3513 2027 3516
rect 2033 3513 2047 3516
rect 2096 3487 2103 3553
rect 2156 3547 2163 3673
rect 2176 3627 2183 3693
rect 2153 3533 2167 3547
rect 2196 3527 2203 3693
rect 2216 3687 2223 3716
rect 2253 3713 2267 3716
rect 2273 3693 2287 3707
rect 2313 3693 2327 3707
rect 2353 3693 2367 3707
rect 2373 3713 2387 3727
rect 2276 3687 2283 3693
rect 2193 3513 2207 3527
rect 1876 3276 1903 3283
rect 1896 3247 1903 3276
rect 1916 3247 1923 3476
rect 2236 3327 2243 3613
rect 2296 3527 2303 3673
rect 2316 3547 2323 3693
rect 2356 3687 2363 3693
rect 2453 3723 2467 3727
rect 2453 3716 2483 3723
rect 2453 3713 2467 3716
rect 2476 3687 2483 3716
rect 2553 3693 2567 3707
rect 2636 3723 2643 3813
rect 2716 3747 2723 3933
rect 2756 3927 2763 4173
rect 2776 3987 2783 4173
rect 2816 4027 2823 4193
rect 2873 4173 2887 4187
rect 2953 4203 2967 4207
rect 2953 4196 2983 4203
rect 2953 4193 2967 4196
rect 2876 4167 2883 4173
rect 2976 4183 2983 4196
rect 2993 4183 3007 4187
rect 2976 4176 3007 4183
rect 3033 4183 3047 4187
rect 3056 4183 3063 4193
rect 2993 4173 3007 4176
rect 2933 4153 2947 4167
rect 3033 4176 3063 4183
rect 3153 4183 3167 4187
rect 3033 4173 3047 4176
rect 3113 4163 3127 4167
rect 3136 4176 3167 4183
rect 3136 4163 3143 4176
rect 3113 4156 3143 4163
rect 3153 4173 3167 4176
rect 3113 4153 3127 4156
rect 2916 4047 2923 4153
rect 2936 4127 2943 4153
rect 2916 4007 2923 4033
rect 2936 4027 2943 4053
rect 2933 4013 2947 4027
rect 2913 3993 2927 4007
rect 2956 4007 2963 4013
rect 2793 3973 2807 3987
rect 2796 3967 2803 3973
rect 2953 3993 2967 4007
rect 2976 3967 2983 4053
rect 2996 4007 3003 4033
rect 3016 4027 3023 4153
rect 2993 3993 3007 4007
rect 3136 4007 3143 4156
rect 3177 4144 3185 4224
rect 3233 4183 3247 4187
rect 3256 4183 3263 4413
rect 3336 4404 3344 4516
rect 3356 4427 3363 4633
rect 3436 4624 3444 4736
rect 3456 4527 3463 5113
rect 3476 5087 3483 5113
rect 3556 5067 3563 5113
rect 3476 4884 3484 4996
rect 3513 4963 3527 4967
rect 3513 4956 3543 4963
rect 3513 4953 3527 4956
rect 3496 4687 3503 4953
rect 3536 4947 3543 4956
rect 3576 4787 3583 5133
rect 3513 4673 3527 4687
rect 3376 4467 3383 4513
rect 3396 4487 3403 4493
rect 3393 4473 3407 4487
rect 3233 4176 3263 4183
rect 3233 4173 3247 4176
rect 3273 4173 3287 4187
rect 3276 4167 3283 4173
rect 3316 4144 3324 4256
rect 3396 4207 3403 4333
rect 3416 4227 3423 4253
rect 3436 4227 3443 4433
rect 3393 4193 3407 4207
rect 3413 4173 3427 4187
rect 3476 4183 3483 4453
rect 3496 4347 3503 4493
rect 3516 4487 3523 4673
rect 3573 4653 3587 4667
rect 3576 4647 3583 4653
rect 3576 4487 3583 4493
rect 3553 4453 3567 4467
rect 3573 4473 3587 4487
rect 3496 4227 3503 4333
rect 3516 4247 3523 4393
rect 3556 4367 3563 4453
rect 3596 4427 3603 4953
rect 3615 4916 3623 4996
rect 3633 4953 3647 4967
rect 3636 4907 3643 4953
rect 3656 4947 3663 5033
rect 3676 4967 3683 5273
rect 3696 5127 3703 5193
rect 3816 5167 3823 5393
rect 3713 5153 3727 5167
rect 3716 5147 3723 5153
rect 3773 5143 3787 5147
rect 3793 5143 3807 5147
rect 3773 5136 3807 5143
rect 3773 5133 3787 5136
rect 3793 5133 3807 5136
rect 3673 4953 3687 4967
rect 3615 4878 3623 4902
rect 3656 4867 3663 4913
rect 3716 4727 3723 4913
rect 3673 4703 3687 4707
rect 3656 4696 3687 4703
rect 3713 4703 3727 4707
rect 3736 4703 3743 4793
rect 3756 4767 3763 4973
rect 3776 4707 3783 5093
rect 3796 5087 3803 5133
rect 3816 4983 3823 5053
rect 3836 5007 3843 5133
rect 3856 5087 3863 5413
rect 3876 5307 3883 5433
rect 3933 5433 3947 5447
rect 3973 5413 3987 5427
rect 4016 5427 4023 5433
rect 4013 5413 4027 5427
rect 3896 5283 3903 5393
rect 3876 5276 3903 5283
rect 3876 5207 3883 5276
rect 3916 5207 3923 5413
rect 3976 5387 3983 5413
rect 4036 5407 4043 5453
rect 4116 5427 4123 5453
rect 4073 5393 4087 5407
rect 4133 5423 4147 5427
rect 4156 5423 4163 5593
rect 4196 5427 4203 5573
rect 4216 5527 4223 5613
rect 4236 5567 4243 5633
rect 4276 5587 4283 5633
rect 4133 5416 4163 5423
rect 4133 5413 4147 5416
rect 3956 5227 3963 5333
rect 4016 5267 4023 5333
rect 3876 5187 3883 5193
rect 3873 5173 3887 5187
rect 3913 5183 3927 5187
rect 3913 5176 3933 5183
rect 3913 5173 3927 5176
rect 3796 4976 3823 4983
rect 3796 4967 3803 4976
rect 3793 4953 3807 4967
rect 3816 4847 3823 4913
rect 3836 4827 3843 4913
rect 3856 4887 3863 4933
rect 3636 4687 3643 4693
rect 3633 4673 3647 4687
rect 3656 4667 3663 4696
rect 3673 4693 3687 4696
rect 3713 4696 3743 4703
rect 3713 4693 3727 4696
rect 3736 4647 3743 4696
rect 3773 4653 3787 4667
rect 3813 4663 3827 4667
rect 3836 4663 3843 4793
rect 3856 4767 3863 4833
rect 3876 4807 3883 5113
rect 3896 5007 3903 5053
rect 3936 5027 3943 5173
rect 3956 5107 3963 5213
rect 4016 5187 4023 5233
rect 4036 5187 4043 5293
rect 4056 5187 4063 5393
rect 4076 5387 4083 5393
rect 4096 5227 4103 5353
rect 4127 5276 4143 5283
rect 3993 5153 4007 5167
rect 3996 5147 4003 5153
rect 3916 4967 3923 4993
rect 3916 4947 3923 4953
rect 3913 4933 3927 4947
rect 3936 4927 3943 4973
rect 3956 4967 3963 5073
rect 3996 4987 4003 5053
rect 4016 4987 4023 5133
rect 4036 4987 4043 5053
rect 4096 5047 4103 5113
rect 4033 4973 4047 4987
rect 3993 4963 4007 4967
rect 3976 4956 4007 4963
rect 3933 4913 3947 4927
rect 3976 4867 3983 4956
rect 3993 4953 4007 4956
rect 4076 4947 4083 4993
rect 4096 4967 4103 5033
rect 4116 5007 4123 5253
rect 4093 4953 4107 4967
rect 4013 4933 4027 4947
rect 4113 4933 4127 4947
rect 4016 4927 4023 4933
rect 3996 4807 4003 4913
rect 3856 4687 3863 4753
rect 3813 4656 3843 4663
rect 3813 4653 3827 4656
rect 3696 4636 3713 4643
rect 3636 4404 3644 4516
rect 3493 4213 3507 4227
rect 3533 4223 3547 4227
rect 3533 4216 3563 4223
rect 3533 4213 3547 4216
rect 3476 4176 3503 4183
rect 3416 4167 3423 4173
rect 3156 4007 3163 4113
rect 3176 4027 3183 4033
rect 3173 4013 3187 4027
rect 3153 3993 3167 4007
rect 3216 3963 3223 4033
rect 3276 3987 3283 3993
rect 3196 3956 3223 3963
rect 2653 3723 2667 3727
rect 2636 3716 2667 3723
rect 2653 3713 2667 3716
rect 2693 3713 2707 3727
rect 2713 3733 2727 3747
rect 2433 3673 2447 3687
rect 2533 3673 2547 3687
rect 2313 3533 2327 3547
rect 2333 3523 2347 3527
rect 2333 3516 2363 3523
rect 2333 3513 2347 3516
rect 2356 3487 2363 3516
rect 2397 3476 2405 3556
rect 2436 3547 2443 3673
rect 2496 3547 2503 3653
rect 2536 3627 2543 3673
rect 2556 3567 2563 3693
rect 2453 3523 2467 3527
rect 2493 3523 2507 3527
rect 2436 3516 2467 3523
rect 2436 3507 2443 3516
rect 2453 3513 2467 3516
rect 2476 3516 2507 3523
rect 2397 3438 2405 3462
rect 1833 3233 1847 3247
rect 1873 3233 1887 3247
rect 1933 3243 1947 3247
rect 1927 3236 1947 3243
rect 1933 3233 1947 3236
rect 1836 3227 1843 3233
rect 1716 3047 1723 3073
rect 1756 3047 1763 3093
rect 1713 3033 1727 3047
rect 1696 3027 1703 3033
rect 1693 3013 1707 3027
rect 1753 3033 1767 3047
rect 1776 3027 1783 3073
rect 1816 3067 1823 3213
rect 1813 3053 1827 3067
rect 1836 3047 1843 3053
rect 1536 2796 1563 2803
rect 1556 2767 1563 2796
rect 1616 2787 1623 2793
rect 1613 2773 1627 2787
rect 1456 2727 1463 2753
rect 1513 2733 1527 2747
rect 1596 2747 1603 2773
rect 1633 2753 1647 2767
rect 1496 2607 1503 2713
rect 1416 2596 1443 2603
rect 1376 2587 1383 2593
rect 1373 2573 1387 2587
rect 1393 2563 1407 2567
rect 1416 2563 1423 2596
rect 1293 2513 1307 2527
rect 1393 2556 1423 2563
rect 1393 2553 1407 2556
rect 1296 2507 1303 2513
rect 1416 2507 1423 2556
rect 1496 2527 1503 2593
rect 1516 2587 1523 2733
rect 1536 2727 1543 2733
rect 1573 2733 1587 2747
rect 1576 2703 1583 2733
rect 1556 2696 1583 2703
rect 1536 2567 1543 2613
rect 1556 2587 1563 2696
rect 1596 2667 1603 2713
rect 1576 2567 1583 2633
rect 1616 2627 1623 2713
rect 1636 2647 1643 2753
rect 1676 2743 1683 2793
rect 1693 2743 1707 2747
rect 1676 2736 1707 2743
rect 1733 2743 1747 2747
rect 1756 2743 1763 2773
rect 1693 2733 1707 2736
rect 1733 2736 1763 2743
rect 1733 2733 1747 2736
rect 1776 2723 1783 2913
rect 1856 2787 1863 3233
rect 1876 3203 1883 3233
rect 1953 3213 1967 3227
rect 1913 3203 1927 3207
rect 1956 3203 1963 3213
rect 1876 3196 1927 3203
rect 1913 3193 1927 3196
rect 1936 3196 1963 3203
rect 1916 3167 1923 3193
rect 1876 3047 1883 3073
rect 1936 3047 1943 3196
rect 2036 3184 2044 3296
rect 2175 3278 2183 3302
rect 2276 3267 2283 3333
rect 2073 3213 2087 3227
rect 2113 3223 2127 3227
rect 2096 3216 2127 3223
rect 1956 3047 1963 3053
rect 1996 3047 2003 3093
rect 2076 3047 2083 3213
rect 2096 3067 2103 3216
rect 2113 3213 2127 3216
rect 2175 3184 2183 3264
rect 2196 3227 2203 3253
rect 2253 3233 2267 3247
rect 2273 3253 2287 3267
rect 2193 3213 2207 3227
rect 2256 3087 2263 3233
rect 2313 3213 2327 3227
rect 2316 3187 2323 3213
rect 2333 3193 2347 3207
rect 1873 3033 1887 3047
rect 1953 3033 1967 3047
rect 1993 3033 2007 3047
rect 2073 3033 2087 3047
rect 2093 3023 2107 3027
rect 2093 3016 2113 3023
rect 2093 3013 2107 3016
rect 1896 2787 1903 2993
rect 1916 2767 1923 3013
rect 2056 2887 2063 3013
rect 2076 2967 2083 2993
rect 1936 2767 1943 2773
rect 1996 2767 2003 2773
rect 1793 2753 1807 2767
rect 1756 2716 1783 2723
rect 1533 2553 1547 2567
rect 1516 2547 1523 2553
rect 1513 2533 1527 2547
rect 1553 2533 1567 2547
rect 1573 2553 1587 2567
rect 1556 2527 1563 2533
rect 1636 2484 1644 2596
rect 1256 2224 1264 2336
rect 1395 2318 1403 2342
rect 1293 2263 1307 2267
rect 1316 2263 1323 2293
rect 1293 2256 1323 2263
rect 1293 2253 1307 2256
rect 1333 2253 1347 2267
rect 1336 2247 1343 2253
rect 1395 2224 1403 2304
rect 1413 2263 1427 2267
rect 1436 2263 1443 2413
rect 1413 2256 1443 2263
rect 1413 2253 1427 2256
rect 1436 2247 1443 2256
rect 1216 2096 1243 2103
rect 1176 1927 1183 1973
rect 1156 1807 1163 1873
rect 1196 1847 1203 1873
rect 1216 1867 1223 2096
rect 1233 2083 1247 2087
rect 1233 2076 1263 2083
rect 1233 2073 1247 2076
rect 1236 1867 1243 2033
rect 1256 2007 1263 2076
rect 1276 1847 1283 2173
rect 1295 2036 1303 2116
rect 1356 2107 1363 2133
rect 1456 2107 1463 2473
rect 1536 2287 1543 2313
rect 1533 2273 1547 2287
rect 1593 2253 1607 2267
rect 1496 2107 1503 2113
rect 1353 2103 1367 2107
rect 1313 2083 1327 2087
rect 1336 2096 1367 2103
rect 1336 2083 1343 2096
rect 1313 2076 1343 2083
rect 1353 2093 1367 2096
rect 1413 2083 1427 2087
rect 1313 2073 1327 2076
rect 1373 2063 1387 2067
rect 1396 2076 1427 2083
rect 1396 2063 1403 2076
rect 1373 2056 1403 2063
rect 1413 2073 1427 2076
rect 1373 2053 1387 2056
rect 1433 2053 1447 2067
rect 1516 2067 1523 2153
rect 1295 1998 1303 2022
rect 1356 1987 1363 2053
rect 1436 1967 1443 2053
rect 1093 1803 1107 1807
rect 1093 1796 1123 1803
rect 1093 1793 1107 1796
rect 1116 1783 1123 1796
rect 1133 1783 1147 1787
rect 1116 1776 1147 1783
rect 1153 1793 1167 1807
rect 1116 1767 1123 1776
rect 1133 1773 1147 1776
rect 1073 1763 1087 1767
rect 1056 1756 1087 1763
rect 1073 1753 1087 1756
rect 1136 1647 1143 1753
rect 1196 1723 1203 1773
rect 1196 1716 1223 1723
rect 1056 1636 1103 1643
rect 913 1603 927 1607
rect 913 1596 943 1603
rect 913 1593 927 1596
rect 916 1367 923 1533
rect 936 1507 943 1596
rect 975 1556 983 1636
rect 1056 1627 1063 1636
rect 1096 1627 1103 1636
rect 993 1593 1007 1607
rect 975 1518 983 1542
rect 996 1527 1003 1593
rect 1176 1607 1183 1653
rect 1053 1573 1067 1587
rect 1153 1573 1167 1587
rect 1173 1593 1187 1607
rect 1056 1567 1063 1573
rect 1076 1427 1083 1573
rect 1156 1547 1163 1573
rect 873 1293 887 1307
rect 733 1133 747 1147
rect 713 1113 727 1127
rect 756 1127 763 1153
rect 816 1143 823 1153
rect 816 1136 863 1143
rect 573 1093 587 1107
rect 613 1103 627 1107
rect 596 1096 627 1103
rect 576 1087 583 1093
rect 496 847 503 873
rect 596 847 603 1096
rect 613 1093 627 1096
rect 636 1087 643 1113
rect 633 1073 647 1087
rect 753 1113 767 1127
rect 673 1073 687 1087
rect 616 1027 623 1033
rect 616 867 623 1013
rect 676 927 683 1073
rect 696 887 703 1093
rect 756 947 763 1073
rect 776 1027 783 1113
rect 796 1107 803 1133
rect 856 1127 863 1136
rect 816 1087 823 1113
rect 836 1107 843 1113
rect 833 1093 847 1107
rect 813 1073 827 1087
rect 853 1073 867 1087
rect 836 1027 843 1053
rect 453 833 467 847
rect 473 803 487 807
rect 456 796 487 803
rect 456 767 463 796
rect 473 793 487 796
rect 93 613 107 627
rect 153 623 167 627
rect 147 616 167 623
rect 153 613 167 616
rect 193 613 207 627
rect 213 633 227 647
rect 196 607 203 613
rect 236 607 243 673
rect 256 667 263 693
rect 273 613 287 627
rect 76 583 83 593
rect 136 583 143 593
rect 76 576 143 583
rect 57 398 65 422
rect 33 343 47 347
rect 16 336 47 343
rect 33 333 47 336
rect 16 163 23 313
rect 57 304 65 384
rect 113 333 127 347
rect 116 327 123 333
rect 33 163 47 167
rect 16 156 47 163
rect 33 153 47 156
rect 57 116 65 196
rect 116 187 123 313
rect 196 304 204 416
rect 256 387 263 613
rect 276 567 283 613
rect 296 463 303 633
rect 316 547 323 653
rect 456 627 463 653
rect 393 613 407 627
rect 356 607 363 613
rect 396 527 403 613
rect 473 593 487 607
rect 416 567 423 573
rect 476 527 483 593
rect 296 456 323 463
rect 296 304 304 416
rect 316 343 323 456
rect 333 343 347 347
rect 316 336 347 343
rect 333 333 347 336
rect 373 333 387 347
rect 376 327 383 333
rect 116 167 123 173
rect 113 153 127 167
rect 57 78 65 102
rect 196 84 204 196
rect 297 116 305 196
rect 356 167 363 173
rect 396 167 403 453
rect 435 398 443 422
rect 435 304 443 384
rect 456 367 463 413
rect 496 403 503 813
rect 553 813 567 827
rect 673 833 687 847
rect 716 843 723 873
rect 796 867 803 893
rect 733 843 747 847
rect 716 836 747 843
rect 733 833 747 836
rect 533 793 547 807
rect 516 427 523 753
rect 536 667 543 793
rect 556 747 563 813
rect 576 807 583 813
rect 593 793 607 807
rect 576 767 583 793
rect 596 627 603 793
rect 676 767 683 833
rect 696 667 703 733
rect 693 653 707 667
rect 736 627 743 813
rect 756 787 763 853
rect 773 833 787 847
rect 793 853 807 867
rect 776 827 783 833
rect 573 593 587 607
rect 613 593 627 607
rect 773 613 787 627
rect 776 607 783 613
rect 556 547 563 573
rect 576 567 583 593
rect 476 396 503 403
rect 456 347 463 353
rect 453 333 467 347
rect 476 327 483 396
rect 556 396 573 403
rect 556 387 563 396
rect 553 373 567 387
rect 596 383 603 593
rect 616 587 623 593
rect 796 587 803 813
rect 816 643 823 933
rect 836 867 843 1013
rect 856 847 863 1073
rect 876 867 883 1253
rect 916 1167 923 1353
rect 976 1347 983 1353
rect 973 1333 987 1347
rect 1053 1343 1067 1347
rect 993 1313 1007 1327
rect 1033 1313 1047 1327
rect 1053 1336 1083 1343
rect 1053 1333 1067 1336
rect 996 1307 1003 1313
rect 976 1147 983 1293
rect 1036 1287 1043 1313
rect 1076 1303 1083 1336
rect 1093 1303 1107 1307
rect 1076 1296 1107 1303
rect 1176 1307 1183 1453
rect 1093 1293 1107 1296
rect 1113 1273 1127 1287
rect 893 1073 907 1087
rect 956 1087 963 1113
rect 993 1093 1007 1107
rect 896 1067 903 1073
rect 896 847 903 893
rect 936 887 943 1053
rect 976 927 983 1093
rect 996 1087 1003 1093
rect 1076 1044 1084 1156
rect 1116 1127 1123 1273
rect 1113 1113 1127 1127
rect 1153 1123 1167 1127
rect 1153 1116 1183 1123
rect 1153 1113 1167 1116
rect 1176 1087 1183 1116
rect 1196 983 1203 1633
rect 1216 1627 1223 1716
rect 1216 1467 1223 1593
rect 1236 1587 1243 1833
rect 1273 1793 1287 1807
rect 1276 1687 1283 1793
rect 1256 1607 1263 1633
rect 1296 1607 1303 1693
rect 1253 1593 1267 1607
rect 1273 1573 1287 1587
rect 1293 1593 1307 1607
rect 1276 1567 1283 1573
rect 1316 1567 1323 1853
rect 1356 1847 1363 1913
rect 1396 1847 1403 1893
rect 1353 1803 1367 1807
rect 1353 1796 1373 1803
rect 1353 1793 1367 1796
rect 1393 1803 1407 1807
rect 1416 1803 1423 1953
rect 1436 1807 1443 1913
rect 1393 1796 1423 1803
rect 1393 1793 1407 1796
rect 1433 1793 1447 1807
rect 1456 1787 1463 1873
rect 1356 1627 1363 1653
rect 1353 1613 1367 1627
rect 1333 1593 1347 1607
rect 1376 1607 1383 1673
rect 1373 1593 1387 1607
rect 1216 1264 1224 1376
rect 1256 1367 1263 1553
rect 1356 1547 1363 1573
rect 1316 1327 1323 1493
rect 1396 1487 1403 1693
rect 1476 1667 1483 1953
rect 1516 1907 1523 2033
rect 1496 1687 1503 1753
rect 1516 1744 1524 1856
rect 1416 1527 1423 1553
rect 1293 1303 1307 1307
rect 1316 1303 1323 1313
rect 1293 1296 1323 1303
rect 1293 1293 1307 1296
rect 1215 1076 1223 1156
rect 1233 1113 1247 1127
rect 1215 1038 1223 1062
rect 1176 976 1203 983
rect 956 863 963 913
rect 1036 887 1043 893
rect 1096 876 1143 883
rect 956 856 983 863
rect 833 813 847 827
rect 853 833 867 847
rect 893 833 907 847
rect 836 767 843 813
rect 936 803 943 853
rect 976 847 983 856
rect 973 833 987 847
rect 1013 833 1027 847
rect 1016 827 1023 833
rect 956 807 963 813
rect 896 796 943 803
rect 856 667 863 673
rect 853 653 867 667
rect 816 636 833 643
rect 876 647 883 653
rect 873 633 887 647
rect 896 607 903 796
rect 636 547 643 573
rect 576 376 603 383
rect 576 307 583 376
rect 593 333 607 347
rect 596 327 603 333
rect 633 333 647 347
rect 613 313 627 327
rect 353 153 367 167
rect 393 153 407 167
rect 297 78 305 102
rect 436 84 444 196
rect 556 167 563 193
rect 576 167 583 193
rect 616 183 623 313
rect 636 307 643 333
rect 676 307 683 393
rect 756 387 763 393
rect 753 373 767 387
rect 793 383 807 387
rect 773 353 787 367
rect 793 376 823 383
rect 793 373 807 376
rect 733 333 747 347
rect 713 313 727 327
rect 716 207 723 313
rect 736 307 743 333
rect 776 327 783 353
rect 616 176 643 183
rect 513 163 527 167
rect 513 156 543 163
rect 513 153 527 156
rect 536 -17 543 156
rect 553 153 567 167
rect 573 153 587 167
rect 636 127 643 176
rect 656 167 663 193
rect 673 163 687 167
rect 673 156 703 163
rect 673 153 687 156
rect 516 -24 543 -17
rect 596 -24 603 113
rect 696 -17 703 156
rect 676 -24 703 -17
rect 736 -24 743 293
rect 816 227 823 376
rect 836 367 843 573
rect 856 387 863 593
rect 916 547 923 673
rect 933 613 947 627
rect 936 567 943 613
rect 873 313 887 327
rect 876 227 883 313
rect 936 304 944 416
rect 777 116 785 196
rect 836 167 843 173
rect 833 153 847 167
rect 873 163 887 167
rect 856 156 887 163
rect 856 127 863 156
rect 873 153 887 156
rect 777 78 785 102
rect 916 84 924 196
rect 956 167 963 733
rect 1016 383 1023 773
rect 1036 647 1043 873
rect 1096 867 1103 876
rect 1113 843 1127 847
rect 1136 843 1143 876
rect 1113 836 1143 843
rect 1113 833 1127 836
rect 1176 827 1183 976
rect 1196 847 1203 913
rect 1236 907 1243 1113
rect 1336 1107 1343 1373
rect 1355 1358 1363 1382
rect 1355 1264 1363 1344
rect 1376 1307 1383 1413
rect 1373 1293 1387 1307
rect 1336 927 1343 1093
rect 1193 833 1207 847
rect 1093 823 1107 827
rect 1093 816 1113 823
rect 1093 813 1107 816
rect 1233 813 1247 827
rect 1276 823 1283 893
rect 1356 847 1363 853
rect 1293 823 1307 827
rect 1276 816 1307 823
rect 1293 813 1307 816
rect 1353 833 1367 847
rect 1393 833 1407 847
rect 1373 813 1387 827
rect 1067 796 1103 803
rect 1096 767 1103 796
rect 1136 767 1143 813
rect 1033 633 1047 647
rect 1116 564 1124 676
rect 1075 398 1083 422
rect 1016 376 1043 383
rect 973 333 987 347
rect 1013 343 1027 347
rect 1036 343 1043 376
rect 1013 336 1043 343
rect 1013 333 1027 336
rect 976 283 983 333
rect 1075 304 1083 384
rect 1093 343 1107 347
rect 1093 336 1123 343
rect 1093 333 1107 336
rect 1116 287 1123 336
rect 1136 327 1143 753
rect 1156 647 1163 813
rect 1236 807 1243 813
rect 1336 803 1343 813
rect 1336 796 1363 803
rect 1153 633 1167 647
rect 1193 643 1207 647
rect 1176 636 1207 643
rect 1153 333 1167 347
rect 976 276 1003 283
rect 976 167 983 193
rect 973 153 987 167
rect 996 107 1003 276
rect 1156 227 1163 333
rect 1013 163 1027 167
rect 1013 156 1043 163
rect 1013 153 1027 156
rect 1036 27 1043 156
rect 1073 113 1087 127
rect 1113 123 1127 127
rect 1136 123 1143 213
rect 1176 187 1183 636
rect 1193 633 1207 636
rect 1255 596 1263 676
rect 1356 667 1363 796
rect 1376 667 1383 813
rect 1396 783 1403 833
rect 1416 807 1423 1393
rect 1436 1327 1443 1433
rect 1456 1247 1463 1633
rect 1516 1587 1523 1673
rect 1536 1647 1543 2213
rect 1596 2207 1603 2253
rect 1616 2107 1623 2313
rect 1636 2307 1643 2393
rect 1656 2327 1663 2653
rect 1676 2567 1683 2613
rect 1716 2567 1723 2693
rect 1673 2553 1687 2567
rect 1713 2553 1727 2567
rect 1756 2547 1763 2716
rect 1796 2647 1803 2753
rect 1933 2753 1947 2767
rect 1856 2727 1863 2733
rect 1973 2733 1987 2747
rect 1993 2753 2007 2767
rect 2033 2753 2047 2767
rect 2013 2733 2027 2747
rect 1873 2713 1887 2727
rect 1775 2516 1783 2596
rect 1836 2587 1843 2633
rect 1833 2573 1847 2587
rect 1793 2563 1807 2567
rect 1816 2563 1823 2573
rect 1793 2556 1823 2563
rect 1793 2553 1807 2556
rect 1853 2543 1867 2547
rect 1876 2543 1883 2713
rect 1896 2587 1903 2593
rect 1853 2536 1883 2543
rect 1853 2533 1867 2536
rect 1775 2478 1783 2502
rect 1656 2287 1663 2293
rect 1633 2253 1647 2267
rect 1653 2273 1667 2287
rect 1636 2127 1643 2253
rect 1696 2207 1703 2273
rect 1656 2123 1663 2193
rect 1696 2187 1703 2193
rect 1656 2116 1683 2123
rect 1556 2067 1563 2093
rect 1676 2087 1683 2116
rect 1716 2103 1723 2293
rect 1736 2267 1743 2433
rect 1753 2253 1767 2267
rect 1756 2187 1763 2253
rect 1716 2096 1743 2103
rect 1593 2053 1607 2067
rect 1613 2073 1627 2087
rect 1673 2073 1687 2087
rect 1693 2053 1707 2067
rect 1736 2067 1743 2096
rect 1756 2087 1763 2173
rect 1776 2107 1783 2153
rect 1773 2093 1787 2107
rect 1753 2073 1767 2087
rect 1796 2087 1803 2213
rect 1816 2107 1823 2533
rect 1936 2487 1943 2633
rect 1976 2587 1983 2733
rect 1996 2567 2003 2613
rect 2016 2587 2023 2733
rect 2036 2723 2043 2753
rect 2056 2747 2063 2793
rect 2116 2767 2123 3013
rect 2153 2993 2167 3007
rect 2236 3023 2243 3053
rect 2296 3047 2303 3053
rect 2253 3023 2267 3027
rect 2236 3016 2267 3023
rect 2293 3033 2307 3047
rect 2336 3043 2343 3193
rect 2376 3187 2383 3353
rect 2316 3036 2343 3043
rect 2136 2767 2143 2993
rect 2156 2967 2163 2993
rect 2216 2987 2223 3013
rect 2236 2987 2243 3016
rect 2253 3013 2267 3016
rect 2316 3003 2323 3036
rect 2333 3003 2347 3007
rect 2316 2996 2347 3003
rect 2333 2993 2347 2996
rect 2196 2967 2203 2973
rect 2256 2947 2263 2993
rect 2036 2716 2063 2723
rect 2036 2627 2043 2653
rect 2036 2567 2043 2573
rect 1973 2533 1987 2547
rect 1993 2553 2007 2567
rect 2033 2553 2047 2567
rect 1976 2507 1983 2533
rect 2056 2507 2063 2716
rect 2076 2707 2083 2753
rect 2133 2723 2147 2727
rect 2116 2716 2147 2723
rect 2116 2687 2123 2716
rect 2133 2713 2147 2716
rect 2087 2596 2103 2603
rect 2096 2587 2103 2596
rect 2093 2573 2107 2587
rect 2076 2567 2083 2573
rect 2073 2553 2087 2567
rect 2113 2553 2127 2567
rect 2136 2547 2143 2693
rect 2176 2647 2183 2813
rect 2176 2567 2183 2593
rect 2153 2533 2167 2547
rect 2173 2553 2187 2567
rect 1833 2253 1847 2267
rect 1896 2223 1903 2373
rect 1916 2303 1923 2393
rect 1916 2296 1943 2303
rect 1936 2287 1943 2296
rect 1976 2287 1983 2493
rect 2056 2287 2063 2353
rect 1913 2253 1927 2267
rect 1933 2273 1947 2287
rect 1953 2253 1967 2267
rect 1916 2247 1923 2253
rect 1956 2243 1963 2253
rect 1936 2236 1963 2243
rect 2053 2243 2067 2247
rect 2076 2243 2083 2273
rect 2053 2236 2083 2243
rect 1936 2223 1943 2236
rect 2053 2233 2067 2236
rect 1896 2216 1943 2223
rect 1836 2187 1843 2193
rect 1793 2073 1807 2087
rect 1553 1773 1567 1787
rect 1576 1783 1583 1993
rect 1636 1967 1643 2053
rect 1593 1783 1607 1787
rect 1576 1776 1607 1783
rect 1593 1773 1607 1776
rect 1556 1727 1563 1773
rect 1596 1647 1603 1773
rect 1616 1627 1623 1873
rect 1655 1838 1663 1862
rect 1536 1607 1543 1613
rect 1533 1593 1547 1607
rect 1593 1603 1607 1607
rect 1576 1596 1607 1603
rect 1476 1427 1483 1553
rect 1496 1547 1503 1573
rect 1436 1087 1443 1093
rect 1496 1067 1503 1533
rect 1576 1507 1583 1596
rect 1593 1593 1607 1596
rect 1636 1587 1643 1753
rect 1655 1744 1663 1824
rect 1676 1787 1683 1973
rect 1716 1943 1723 2033
rect 1696 1936 1723 1943
rect 1673 1773 1687 1787
rect 1676 1703 1683 1713
rect 1696 1707 1703 1936
rect 1736 1867 1743 2053
rect 1796 1807 1803 1953
rect 1816 1847 1823 2073
rect 1836 2067 1843 2173
rect 1916 2127 1923 2153
rect 1936 2147 1943 2153
rect 1956 2147 1963 2213
rect 1936 2087 1943 2133
rect 2056 2087 2063 2153
rect 1833 2053 1847 2067
rect 1893 2073 1907 2087
rect 1933 2073 1947 2087
rect 1953 2053 1967 2067
rect 1976 2076 1993 2083
rect 1876 1887 1883 1973
rect 1956 1887 1963 2053
rect 1976 1947 1983 2076
rect 2013 2053 2027 2067
rect 2053 2073 2067 2087
rect 2073 2053 2087 2067
rect 1996 1987 2003 2033
rect 2016 1987 2023 2053
rect 2076 2007 2083 2053
rect 2096 2027 2103 2533
rect 2156 2523 2163 2533
rect 2136 2516 2163 2523
rect 2116 2224 2124 2336
rect 2136 2107 2143 2516
rect 2196 2303 2203 2733
rect 2216 2704 2224 2816
rect 2236 2743 2243 2793
rect 2253 2743 2267 2747
rect 2236 2736 2267 2743
rect 2253 2733 2267 2736
rect 2276 2667 2283 2773
rect 2293 2733 2307 2747
rect 2296 2727 2303 2733
rect 2296 2707 2303 2713
rect 2213 2533 2227 2547
rect 2216 2527 2223 2533
rect 2256 2447 2263 2573
rect 2296 2567 2303 2593
rect 2273 2533 2287 2547
rect 2293 2553 2307 2567
rect 2276 2487 2283 2533
rect 2316 2527 2323 2893
rect 2336 2607 2343 2853
rect 2355 2798 2363 2822
rect 2376 2807 2383 3073
rect 2355 2704 2363 2784
rect 2376 2747 2383 2793
rect 2373 2733 2387 2747
rect 2376 2587 2383 2633
rect 2367 2556 2383 2563
rect 2176 2296 2203 2303
rect 2176 2263 2183 2296
rect 2193 2263 2207 2267
rect 2176 2256 2207 2263
rect 2193 2253 2207 2256
rect 2133 2053 2147 2067
rect 1916 1807 1923 1873
rect 1733 1803 1747 1807
rect 1733 1796 1763 1803
rect 1733 1793 1747 1796
rect 1756 1783 1763 1796
rect 1773 1783 1787 1787
rect 1756 1776 1787 1783
rect 1793 1793 1807 1807
rect 1773 1773 1787 1776
rect 1893 1783 1907 1787
rect 1876 1776 1907 1783
rect 1933 1783 1947 1787
rect 1956 1783 1963 1853
rect 2016 1827 2023 1893
rect 1713 1753 1727 1767
rect 1656 1696 1683 1703
rect 1656 1607 1663 1696
rect 1716 1623 1723 1753
rect 1756 1627 1763 1633
rect 1696 1616 1723 1623
rect 1653 1593 1667 1607
rect 1613 1573 1627 1587
rect 1673 1573 1687 1587
rect 1516 1044 1524 1156
rect 1536 943 1543 1233
rect 1556 1227 1563 1353
rect 1576 1327 1583 1373
rect 1573 1313 1587 1327
rect 1596 1287 1603 1513
rect 1616 1467 1623 1573
rect 1636 1367 1643 1573
rect 1676 1507 1683 1573
rect 1696 1527 1703 1616
rect 1733 1573 1747 1587
rect 1736 1547 1743 1573
rect 1756 1447 1763 1613
rect 1797 1556 1805 1636
rect 1797 1518 1805 1542
rect 1556 1127 1563 1153
rect 1553 1113 1567 1127
rect 1593 1123 1607 1127
rect 1576 1116 1607 1123
rect 1576 1107 1583 1116
rect 1593 1113 1607 1116
rect 1536 936 1563 943
rect 1456 847 1463 853
rect 1453 833 1467 847
rect 1396 776 1423 783
rect 1356 647 1363 653
rect 1255 558 1263 582
rect 1193 343 1207 347
rect 1193 336 1213 343
rect 1193 333 1207 336
rect 1276 347 1283 633
rect 1353 643 1367 647
rect 1353 636 1383 643
rect 1353 633 1367 636
rect 1376 603 1383 636
rect 1416 627 1423 776
rect 1476 687 1483 793
rect 1536 784 1544 896
rect 1556 707 1563 936
rect 1576 863 1583 1093
rect 1616 1027 1623 1333
rect 1656 1327 1663 1353
rect 1633 1293 1647 1307
rect 1653 1313 1667 1327
rect 1636 1287 1643 1293
rect 1576 856 1603 863
rect 1596 823 1603 856
rect 1636 827 1643 1253
rect 1676 1183 1683 1373
rect 1716 1327 1723 1373
rect 1713 1313 1727 1327
rect 1736 1307 1743 1413
rect 1756 1367 1763 1393
rect 1776 1327 1783 1413
rect 1756 1263 1763 1293
rect 1793 1293 1807 1307
rect 1736 1256 1763 1263
rect 1676 1176 1703 1183
rect 1655 1076 1663 1156
rect 1655 1038 1663 1062
rect 1696 987 1703 1176
rect 1736 1127 1743 1256
rect 1796 1247 1803 1293
rect 1816 1247 1823 1693
rect 1836 1347 1843 1633
rect 1856 1627 1863 1733
rect 1856 1607 1863 1613
rect 1853 1593 1867 1607
rect 1876 1587 1883 1776
rect 1893 1773 1907 1776
rect 1933 1776 1963 1783
rect 1933 1773 1947 1776
rect 1973 1773 1987 1787
rect 1993 1793 2007 1807
rect 2033 1793 2047 1807
rect 1976 1767 1983 1773
rect 2036 1763 2043 1793
rect 2016 1756 2043 1763
rect 1896 1607 1903 1693
rect 1893 1593 1907 1607
rect 1876 1527 1883 1573
rect 1936 1524 1944 1636
rect 1956 1567 1963 1693
rect 1976 1487 1983 1753
rect 2016 1667 2023 1756
rect 2076 1727 2083 1953
rect 2096 1807 2103 1933
rect 2116 1907 2123 2013
rect 2136 1907 2143 2053
rect 2156 1887 2163 2173
rect 2117 1838 2125 1862
rect 2096 1787 2103 1793
rect 2093 1773 2107 1787
rect 2117 1744 2125 1824
rect 2136 1747 2143 1873
rect 2176 1823 2183 2233
rect 2216 2127 2223 2393
rect 2236 2267 2243 2373
rect 2255 2318 2263 2342
rect 2255 2224 2263 2304
rect 2276 2267 2283 2273
rect 2273 2253 2287 2267
rect 2196 2004 2204 2116
rect 2216 1867 2223 2113
rect 2236 2087 2243 2153
rect 2276 2123 2283 2213
rect 2296 2147 2303 2353
rect 2276 2116 2303 2123
rect 2233 2073 2247 2087
rect 2176 1816 2203 1823
rect 2173 1773 2187 1787
rect 2176 1747 2183 1773
rect 2076 1607 2083 1713
rect 2196 1627 2203 1816
rect 2213 1773 2227 1787
rect 2216 1747 2223 1773
rect 2236 1647 2243 1973
rect 2256 1744 2264 1856
rect 2276 1707 2283 2033
rect 2296 2007 2303 2116
rect 2316 2047 2323 2433
rect 2356 2287 2363 2433
rect 2376 2427 2383 2556
rect 2396 2327 2403 3393
rect 2476 3227 2483 3516
rect 2493 3513 2507 3516
rect 2536 3444 2544 3556
rect 2616 3547 2623 3633
rect 2613 3533 2627 3547
rect 2556 3267 2563 3533
rect 2593 3523 2607 3527
rect 2576 3516 2607 3523
rect 2636 3527 2643 3533
rect 2576 3483 2583 3516
rect 2593 3513 2607 3516
rect 2633 3513 2647 3527
rect 2576 3476 2603 3483
rect 2596 3347 2603 3476
rect 2656 3427 2663 3713
rect 2696 3703 2703 3713
rect 2756 3707 2763 3793
rect 2796 3747 2803 3773
rect 2836 3747 2843 3753
rect 2876 3747 2883 3793
rect 2896 3747 2903 3813
rect 2833 3743 2847 3747
rect 2827 3736 2847 3743
rect 2833 3733 2847 3736
rect 2776 3727 2783 3733
rect 2853 3713 2867 3727
rect 2873 3733 2887 3747
rect 2916 3727 2923 3753
rect 2696 3696 2723 3703
rect 2676 3587 2683 3613
rect 2676 3527 2683 3573
rect 2716 3527 2723 3696
rect 2756 3563 2763 3693
rect 2856 3703 2863 3713
rect 2827 3696 2863 3703
rect 2913 3713 2927 3727
rect 2933 3693 2947 3707
rect 2756 3556 2783 3563
rect 2673 3513 2687 3527
rect 2713 3513 2727 3527
rect 2733 3503 2747 3507
rect 2756 3503 2763 3533
rect 2733 3496 2763 3503
rect 2733 3493 2747 3496
rect 2756 3487 2763 3496
rect 2776 3447 2783 3556
rect 2816 3547 2823 3553
rect 2856 3547 2863 3673
rect 2936 3627 2943 3693
rect 2813 3543 2827 3547
rect 2813 3536 2843 3543
rect 2813 3533 2827 3536
rect 2836 3527 2843 3536
rect 2836 3467 2843 3513
rect 2876 3507 2883 3533
rect 2956 3527 2963 3693
rect 2976 3587 2983 3753
rect 3036 3747 3043 3953
rect 3096 3727 3103 3753
rect 3116 3727 3123 3793
rect 3136 3727 3143 3733
rect 3176 3727 3183 3773
rect 2993 3693 3007 3707
rect 3053 3723 3067 3727
rect 3053 3716 3073 3723
rect 3053 3713 3067 3716
rect 3093 3713 3107 3727
rect 3133 3713 3147 3727
rect 3033 3693 3047 3707
rect 2996 3627 3003 3693
rect 3036 3627 3043 3693
rect 3056 3667 3063 3693
rect 3196 3667 3203 3956
rect 3273 3973 3287 3987
rect 3333 3953 3347 3967
rect 3373 3963 3387 3967
rect 3396 3963 3403 4113
rect 3373 3956 3403 3963
rect 3373 3953 3387 3956
rect 3236 3747 3243 3933
rect 3316 3767 3323 3953
rect 3336 3947 3343 3953
rect 3436 3924 3444 4036
rect 3336 3767 3343 3793
rect 3456 3787 3463 4153
rect 3276 3727 3283 3753
rect 3376 3747 3383 3753
rect 3333 3743 3347 3747
rect 3327 3736 3347 3743
rect 3333 3733 3347 3736
rect 3253 3693 3267 3707
rect 3273 3713 3287 3727
rect 3293 3693 3307 3707
rect 3036 3547 3043 3573
rect 3236 3547 3243 3673
rect 3256 3667 3263 3693
rect 3296 3687 3303 3693
rect 3316 3687 3323 3733
rect 3373 3733 3387 3747
rect 3413 3743 3427 3747
rect 3396 3736 3427 3743
rect 3453 3743 3467 3747
rect 2853 3473 2867 3487
rect 2873 3493 2887 3507
rect 2933 3493 2947 3507
rect 2953 3513 2967 3527
rect 2976 3507 2983 3533
rect 2973 3493 2987 3507
rect 2893 3473 2907 3487
rect 2936 3483 2943 3493
rect 2927 3476 2943 3483
rect 2856 3447 2863 3473
rect 2896 3467 2903 3473
rect 2596 3247 2603 3333
rect 2493 3233 2507 3247
rect 2416 3027 2423 3213
rect 2453 3213 2467 3227
rect 2436 2964 2444 3076
rect 2456 3067 2463 3213
rect 2496 3207 2503 3233
rect 2593 3233 2607 3247
rect 2573 3203 2587 3207
rect 2567 3196 2587 3203
rect 2573 3193 2587 3196
rect 2496 2867 2503 3113
rect 2556 3087 2563 3193
rect 2513 3043 2527 3047
rect 2513 3036 2543 3043
rect 2513 3033 2527 3036
rect 2416 2787 2423 2793
rect 2413 2773 2427 2787
rect 2516 2767 2523 2773
rect 2513 2753 2527 2767
rect 2493 2713 2507 2727
rect 2416 2307 2423 2653
rect 2496 2607 2503 2713
rect 2536 2707 2543 3036
rect 2575 2996 2583 3076
rect 2633 3063 2647 3067
rect 2593 3043 2607 3047
rect 2616 3056 2647 3063
rect 2656 3063 2663 3413
rect 2676 3184 2684 3296
rect 2815 3278 2823 3302
rect 2713 3213 2727 3227
rect 2716 3067 2723 3213
rect 2656 3056 2683 3063
rect 2616 3043 2623 3056
rect 2593 3036 2623 3043
rect 2633 3053 2647 3056
rect 2593 3033 2607 3036
rect 2575 2958 2583 2982
rect 2593 2723 2607 2727
rect 2616 2723 2623 2993
rect 2593 2716 2623 2723
rect 2593 2713 2607 2716
rect 2656 2704 2664 2816
rect 2436 2484 2444 2596
rect 2473 2563 2487 2567
rect 2456 2556 2487 2563
rect 2456 2443 2463 2556
rect 2473 2553 2487 2556
rect 2513 2553 2527 2567
rect 2436 2436 2463 2443
rect 2436 2307 2443 2436
rect 2456 2347 2463 2413
rect 2333 2253 2347 2267
rect 2336 2207 2343 2253
rect 2393 2253 2407 2267
rect 2396 2247 2403 2253
rect 2335 2036 2343 2116
rect 2376 2087 2383 2133
rect 2353 2073 2367 2087
rect 2335 1998 2343 2022
rect 2356 1947 2363 2073
rect 2296 1936 2343 1943
rect 2296 1847 2303 1936
rect 2336 1927 2343 1936
rect 2376 1943 2383 2073
rect 2396 2023 2403 2173
rect 2436 2087 2443 2153
rect 2456 2147 2463 2253
rect 2476 2187 2483 2513
rect 2536 2347 2543 2593
rect 2556 2547 2563 2593
rect 2575 2516 2583 2596
rect 2656 2567 2663 2593
rect 2633 2533 2647 2547
rect 2653 2553 2667 2567
rect 2575 2478 2583 2502
rect 2556 2347 2563 2433
rect 2576 2327 2583 2413
rect 2596 2407 2603 2533
rect 2616 2447 2623 2493
rect 2616 2303 2623 2413
rect 2636 2307 2643 2533
rect 2676 2467 2683 3056
rect 2713 3053 2727 3067
rect 2736 3047 2743 3273
rect 2753 3213 2767 3227
rect 2733 3033 2747 3047
rect 2693 2743 2707 2747
rect 2716 2743 2723 2853
rect 2693 2736 2723 2743
rect 2693 2733 2707 2736
rect 2733 2733 2747 2747
rect 2736 2707 2743 2733
rect 2756 2707 2763 3213
rect 2796 3147 2803 3213
rect 2815 3184 2823 3264
rect 2813 3063 2827 3067
rect 2836 3063 2843 3153
rect 2813 3056 2843 3063
rect 2813 3053 2827 3056
rect 2856 3047 2863 3293
rect 2876 3287 2883 3433
rect 2896 3287 2903 3453
rect 2916 3307 2923 3473
rect 3036 3467 3043 3493
rect 3096 3487 3103 3533
rect 3136 3527 3143 3533
rect 3113 3493 3127 3507
rect 3133 3513 3147 3527
rect 3156 3507 3163 3533
rect 3276 3527 3283 3533
rect 3213 3493 3227 3507
rect 3273 3513 3287 3527
rect 3116 3427 3123 3493
rect 2893 3233 2907 3247
rect 2896 3223 2903 3233
rect 2896 3216 2923 3223
rect 2876 3087 2883 3213
rect 2896 3067 2903 3193
rect 2916 3167 2923 3216
rect 2936 3187 2943 3273
rect 2956 3107 2963 3333
rect 2976 3267 2983 3273
rect 3016 3267 3023 3273
rect 3036 3267 3043 3353
rect 3056 3307 3063 3313
rect 3076 3267 3083 3373
rect 2973 3253 2987 3267
rect 3013 3253 3027 3267
rect 3036 3227 3043 3233
rect 3116 3203 3123 3213
rect 3096 3196 3123 3203
rect 2876 3047 2883 3053
rect 2916 3047 2923 3093
rect 2956 3047 2963 3093
rect 3096 3047 3103 3196
rect 3136 3047 3143 3473
rect 3216 3467 3223 3493
rect 3156 3267 3163 3293
rect 3196 3267 3203 3273
rect 3153 3253 3167 3267
rect 3193 3263 3207 3267
rect 3193 3256 3223 3263
rect 3193 3253 3207 3256
rect 3216 3227 3223 3256
rect 3236 3247 3243 3373
rect 3256 3267 3263 3413
rect 3296 3283 3303 3653
rect 3396 3607 3403 3736
rect 3413 3733 3427 3736
rect 3453 3736 3483 3743
rect 3453 3733 3467 3736
rect 3333 3543 3347 3547
rect 3356 3543 3363 3593
rect 3333 3536 3363 3543
rect 3333 3533 3347 3536
rect 3356 3523 3363 3536
rect 3373 3523 3387 3527
rect 3356 3516 3387 3523
rect 3373 3513 3387 3516
rect 3276 3276 3303 3283
rect 3233 3233 3247 3247
rect 3276 3107 3283 3276
rect 3336 3247 3343 3493
rect 3397 3476 3405 3556
rect 3453 3513 3467 3527
rect 3397 3438 3405 3462
rect 3476 3387 3483 3736
rect 3496 3727 3503 4176
rect 3556 4127 3563 4216
rect 3576 4147 3583 4253
rect 3596 4207 3603 4373
rect 3593 4203 3607 4207
rect 3593 4196 3623 4203
rect 3593 4193 3607 4196
rect 3516 4007 3523 4013
rect 3556 4007 3563 4113
rect 3513 3993 3527 4007
rect 3575 3956 3583 4036
rect 3575 3918 3583 3942
rect 3616 3887 3623 4196
rect 3676 4027 3683 4053
rect 3673 4013 3687 4027
rect 3653 3973 3667 3987
rect 3656 3967 3663 3973
rect 3516 3664 3524 3776
rect 3696 3787 3703 4636
rect 3713 4483 3727 4487
rect 3713 4476 3743 4483
rect 3713 4473 3727 4476
rect 3736 4427 3743 4476
rect 3756 4447 3763 4653
rect 3776 4627 3783 4653
rect 3775 4436 3783 4516
rect 3793 4483 3807 4487
rect 3816 4483 3823 4553
rect 3836 4487 3843 4656
rect 3876 4624 3884 4736
rect 3913 4653 3927 4667
rect 3916 4627 3923 4653
rect 3936 4567 3943 4793
rect 3953 4653 3967 4667
rect 3856 4507 3863 4533
rect 3793 4476 3823 4483
rect 3793 4473 3807 4476
rect 3833 4473 3847 4487
rect 3893 4463 3907 4467
rect 3893 4456 3923 4463
rect 3893 4453 3907 4456
rect 3736 4207 3743 4413
rect 3775 4398 3783 4422
rect 3816 4227 3823 4313
rect 3773 4223 3787 4227
rect 3756 4216 3787 4223
rect 3756 4127 3763 4216
rect 3773 4213 3787 4216
rect 3813 4213 3827 4227
rect 3736 3924 3744 4036
rect 3776 4007 3783 4033
rect 3816 4027 3823 4173
rect 3816 4007 3823 4013
rect 3773 3993 3787 4007
rect 3813 3993 3827 4007
rect 3836 3947 3843 4433
rect 3856 4227 3863 4313
rect 3916 4247 3923 4456
rect 3936 4447 3943 4513
rect 3956 4427 3963 4653
rect 3996 4627 4003 4773
rect 4015 4718 4023 4742
rect 4015 4624 4023 4704
rect 4036 4667 4043 4933
rect 4116 4927 4123 4933
rect 4087 4916 4103 4923
rect 4033 4653 4047 4667
rect 4056 4647 4063 4913
rect 3976 4404 3984 4516
rect 3996 4367 4003 4613
rect 4053 4483 4067 4487
rect 4036 4476 4067 4483
rect 4036 4427 4043 4476
rect 4053 4473 4067 4476
rect 4076 4367 4083 4853
rect 4096 4787 4103 4916
rect 4116 4907 4123 4913
rect 4136 4907 4143 5276
rect 4156 5267 4163 5416
rect 4173 5393 4187 5407
rect 4193 5413 4207 5427
rect 4253 5423 4267 5427
rect 4276 5423 4283 5513
rect 4253 5416 4283 5423
rect 4253 5413 4267 5416
rect 4213 5403 4227 5407
rect 4236 5403 4243 5413
rect 4213 5396 4243 5403
rect 4213 5393 4227 5396
rect 4176 5227 4183 5393
rect 4196 5267 4203 5333
rect 4216 5327 4223 5333
rect 4156 5203 4163 5213
rect 4216 5207 4223 5313
rect 4156 5196 4203 5203
rect 4196 5187 4203 5196
rect 4193 5173 4207 5187
rect 4156 4987 4163 5133
rect 4153 4963 4167 4967
rect 4176 4963 4183 5133
rect 4216 5127 4223 5193
rect 4236 5187 4243 5396
rect 4276 5327 4283 5416
rect 4296 5387 4303 5613
rect 4316 5583 4323 5633
rect 4376 5627 4383 5733
rect 4396 5667 4403 5713
rect 4516 5707 4523 5916
rect 4533 5913 4547 5916
rect 4573 5916 4623 5923
rect 4573 5913 4587 5916
rect 4593 5913 4607 5916
rect 4473 5613 4487 5627
rect 4496 5623 4503 5693
rect 4536 5667 4543 5733
rect 4616 5727 4623 5916
rect 4633 5873 4647 5887
rect 4636 5707 4643 5873
rect 4656 5747 4663 5753
rect 4596 5667 4603 5673
rect 4533 5653 4547 5667
rect 4633 5663 4647 5667
rect 4656 5663 4663 5733
rect 4513 5623 4527 5627
rect 4496 5616 4527 5623
rect 4556 5623 4563 5653
rect 4633 5656 4663 5663
rect 4633 5653 4647 5656
rect 4573 5623 4587 5627
rect 4556 5616 4587 5623
rect 4513 5613 4527 5616
rect 4573 5613 4587 5616
rect 4476 5607 4483 5613
rect 4316 5576 4343 5583
rect 4316 5427 4323 5553
rect 4336 5447 4343 5576
rect 4436 5547 4443 5593
rect 4576 5567 4583 5613
rect 4333 5433 4347 5447
rect 4353 5413 4367 5427
rect 4436 5427 4443 5533
rect 4496 5427 4503 5453
rect 4516 5447 4523 5533
rect 4233 5133 4247 5147
rect 4236 5107 4243 5133
rect 4256 5027 4263 5133
rect 4276 5127 4283 5213
rect 4296 5207 4303 5353
rect 4356 5347 4363 5413
rect 4376 5367 4383 5393
rect 4293 5133 4307 5147
rect 4276 5087 4283 5113
rect 4296 5107 4303 5133
rect 4316 5107 4323 5213
rect 4356 5203 4363 5273
rect 4347 5196 4363 5203
rect 4376 5187 4383 5213
rect 4373 5173 4387 5187
rect 4396 5167 4403 5413
rect 4413 5393 4427 5407
rect 4433 5413 4447 5427
rect 4473 5393 4487 5407
rect 4493 5413 4507 5427
rect 4416 5247 4423 5393
rect 4436 5307 4443 5373
rect 4456 5323 4463 5373
rect 4476 5367 4483 5393
rect 4516 5367 4523 5393
rect 4536 5347 4543 5473
rect 4456 5316 4483 5323
rect 4436 5187 4443 5293
rect 4476 5287 4483 5316
rect 4456 5167 4463 5213
rect 4413 5153 4427 5167
rect 4153 4956 4183 4963
rect 4153 4953 4167 4956
rect 4196 4927 4203 4973
rect 4216 4967 4223 4993
rect 4256 4967 4263 5013
rect 4213 4953 4227 4967
rect 4276 4947 4283 5013
rect 4296 4967 4303 5073
rect 4316 4967 4323 5093
rect 4336 5087 4343 5133
rect 4416 5127 4423 5153
rect 4496 5147 4503 5333
rect 4556 5287 4563 5513
rect 4596 5447 4603 5613
rect 4616 5607 4623 5633
rect 4636 5447 4643 5533
rect 4656 5447 4663 5656
rect 4676 5487 4683 6073
rect 4696 6047 4703 6113
rect 4736 6107 4743 6133
rect 4756 6047 4763 6213
rect 4876 6147 4883 6173
rect 4773 6093 4787 6107
rect 4913 6133 4927 6147
rect 5016 6147 5023 6313
rect 5036 6307 5043 6373
rect 5096 6307 5103 6376
rect 5116 6343 5123 6473
rect 5156 6447 5163 6473
rect 5456 6463 5463 6476
rect 5496 6467 5503 6476
rect 5336 6456 5463 6463
rect 5336 6447 5343 6456
rect 5156 6387 5163 6433
rect 5196 6416 5243 6423
rect 5196 6403 5203 6416
rect 5176 6396 5203 6403
rect 5153 6373 5167 6387
rect 5176 6367 5183 6396
rect 5236 6403 5243 6416
rect 5236 6396 5273 6403
rect 5173 6353 5187 6367
rect 5116 6336 5163 6343
rect 5156 6323 5163 6336
rect 5216 6327 5223 6393
rect 5233 6353 5247 6367
rect 5276 6367 5283 6393
rect 5273 6353 5287 6367
rect 5316 6363 5323 6393
rect 5356 6387 5363 6433
rect 5433 6423 5447 6427
rect 5396 6416 5447 6423
rect 5396 6407 5403 6416
rect 5433 6413 5447 6416
rect 5333 6363 5347 6367
rect 5316 6356 5347 6363
rect 5353 6373 5367 6387
rect 5376 6367 5383 6393
rect 5476 6407 5483 6453
rect 5413 6373 5427 6387
rect 5453 6373 5467 6387
rect 5473 6393 5487 6407
rect 5333 6353 5347 6356
rect 5373 6353 5387 6367
rect 5236 6347 5243 6353
rect 5156 6316 5193 6323
rect 4893 6113 4907 6127
rect 4776 6067 4783 6093
rect 4696 5847 4703 5953
rect 4716 5927 4723 5973
rect 4756 5947 4763 5953
rect 4753 5933 4767 5947
rect 4713 5913 4727 5927
rect 4773 5893 4787 5907
rect 4736 5667 4743 5833
rect 4756 5667 4763 5893
rect 4776 5887 4783 5893
rect 4793 5873 4807 5887
rect 4833 5873 4847 5887
rect 4796 5727 4803 5873
rect 4836 5707 4843 5873
rect 4856 5867 4863 5893
rect 4876 5843 4883 6073
rect 4896 6067 4903 6113
rect 4916 6107 4923 6133
rect 4973 6133 4987 6147
rect 4953 6123 4967 6127
rect 4947 6116 4967 6123
rect 4953 6113 4967 6116
rect 4916 6087 4923 6093
rect 4893 5893 4907 5907
rect 4896 5887 4903 5893
rect 4936 5883 4943 6113
rect 4976 5987 4983 6133
rect 4993 6113 5007 6127
rect 5013 6133 5027 6147
rect 4996 6107 5003 6113
rect 5016 5907 5023 5953
rect 5036 5947 5043 6153
rect 5116 6147 5123 6273
rect 5256 6267 5263 6333
rect 5296 6307 5303 6333
rect 5216 6147 5223 6153
rect 5276 6147 5283 6153
rect 5173 6143 5187 6147
rect 5156 6136 5187 6143
rect 5073 6113 5087 6127
rect 5076 6067 5083 6113
rect 5156 6107 5163 6136
rect 5173 6133 5187 6136
rect 5193 6113 5207 6127
rect 5213 6133 5227 6147
rect 5273 6133 5287 6147
rect 5133 6093 5147 6107
rect 5056 5947 5063 5953
rect 4953 5883 4967 5887
rect 4936 5876 4967 5883
rect 5013 5893 5027 5907
rect 5073 5893 5087 5907
rect 4953 5873 4967 5876
rect 4896 5867 4903 5873
rect 5036 5847 5043 5873
rect 4876 5836 4903 5843
rect 4856 5727 4863 5733
rect 4753 5623 4767 5627
rect 4753 5616 4773 5623
rect 4753 5613 4767 5616
rect 4833 5643 4847 5647
rect 4856 5643 4863 5693
rect 4833 5636 4863 5643
rect 4833 5633 4847 5636
rect 4813 5623 4827 5627
rect 4813 5616 4833 5623
rect 4813 5613 4827 5616
rect 4736 5463 4743 5573
rect 4776 5567 4783 5613
rect 4816 5596 4853 5603
rect 4676 5456 4743 5463
rect 4676 5447 4683 5456
rect 4593 5433 4607 5447
rect 4576 5427 4583 5433
rect 4573 5413 4587 5427
rect 4613 5413 4627 5427
rect 4633 5433 4647 5447
rect 4673 5423 4687 5427
rect 4656 5416 4687 5423
rect 4576 5267 4583 5353
rect 4516 5227 4523 5253
rect 4596 5187 4603 5233
rect 4616 5227 4623 5413
rect 4656 5403 4663 5416
rect 4636 5396 4663 5403
rect 4673 5413 4687 5416
rect 4636 5347 4643 5396
rect 4756 5387 4763 5553
rect 4776 5467 4783 5533
rect 4796 5487 4803 5593
rect 4816 5587 4823 5596
rect 4836 5447 4843 5453
rect 4833 5433 4847 5447
rect 4793 5393 4807 5407
rect 4636 5207 4643 5293
rect 4593 5173 4607 5187
rect 4556 5167 4563 5173
rect 4473 5133 4487 5147
rect 4553 5153 4567 5167
rect 4656 5147 4663 5373
rect 4676 5287 4683 5373
rect 4676 5187 4683 5273
rect 4716 5207 4723 5353
rect 4716 5187 4723 5193
rect 4673 5173 4687 5187
rect 4713 5173 4727 5187
rect 4736 5167 4743 5253
rect 4796 5247 4803 5393
rect 4816 5327 4823 5413
rect 4856 5387 4863 5553
rect 4876 5447 4883 5713
rect 4896 5667 4903 5836
rect 4893 5653 4907 5667
rect 4933 5653 4947 5667
rect 4913 5633 4927 5647
rect 4916 5567 4923 5633
rect 4936 5587 4943 5653
rect 4976 5647 4983 5733
rect 5056 5667 5063 5893
rect 5076 5867 5083 5893
rect 5116 5887 5123 6073
rect 5136 5927 5143 6093
rect 5196 6087 5203 6113
rect 5233 6103 5247 6107
rect 5227 6096 5247 6103
rect 5233 6093 5247 6096
rect 5293 6103 5307 6107
rect 5316 6103 5323 6333
rect 5356 6147 5363 6293
rect 5416 6287 5423 6373
rect 5456 6367 5463 6373
rect 5293 6096 5323 6103
rect 5293 6093 5307 6096
rect 5333 6093 5347 6107
rect 5393 6123 5407 6127
rect 5416 6123 5423 6253
rect 5456 6207 5463 6353
rect 5496 6287 5503 6433
rect 5536 6407 5543 6473
rect 5576 6427 5583 6433
rect 5573 6413 5587 6427
rect 5533 6393 5547 6407
rect 5593 6373 5607 6387
rect 5596 6347 5603 6373
rect 5616 6267 5623 6413
rect 5736 6407 5743 6453
rect 5756 6407 5763 6433
rect 5796 6407 5803 6453
rect 5896 6407 5903 6493
rect 6016 6447 6023 6453
rect 6013 6423 6027 6427
rect 6036 6423 6043 6433
rect 6013 6416 6043 6423
rect 6013 6413 6027 6416
rect 5713 6373 5727 6387
rect 5733 6393 5747 6407
rect 5893 6393 5907 6407
rect 5773 6383 5787 6387
rect 5756 6376 5787 6383
rect 5676 6367 5683 6373
rect 5716 6347 5723 6373
rect 5393 6116 5423 6123
rect 5393 6113 5407 6116
rect 5436 6103 5443 6133
rect 5453 6103 5467 6107
rect 5436 6096 5467 6103
rect 5513 6123 5527 6127
rect 5536 6123 5543 6153
rect 5556 6147 5563 6253
rect 5513 6116 5543 6123
rect 5553 6133 5567 6147
rect 5513 6113 5527 6116
rect 5453 6093 5467 6096
rect 5176 5927 5183 6033
rect 5196 5967 5203 5973
rect 5153 5893 5167 5907
rect 5173 5913 5187 5927
rect 5196 5907 5203 5953
rect 5216 5907 5223 6093
rect 5336 6087 5343 6093
rect 5536 6103 5543 6116
rect 5573 6113 5587 6127
rect 5576 6103 5583 6113
rect 5536 6096 5583 6103
rect 5236 5927 5243 5933
rect 5276 5927 5283 6053
rect 5376 5927 5383 5953
rect 5576 5947 5583 6096
rect 5596 6087 5603 6133
rect 5653 6133 5667 6147
rect 5616 6087 5623 6113
rect 5533 5943 5547 5947
rect 5516 5936 5547 5943
rect 5233 5913 5247 5927
rect 5193 5893 5207 5907
rect 5253 5893 5267 5907
rect 5273 5913 5287 5927
rect 5293 5903 5307 5907
rect 5293 5896 5323 5903
rect 5293 5893 5307 5896
rect 5156 5887 5163 5893
rect 5256 5887 5263 5893
rect 5096 5667 5103 5873
rect 5116 5667 5123 5833
rect 5016 5647 5023 5653
rect 4973 5633 4987 5647
rect 4956 5607 4963 5633
rect 5013 5633 5027 5647
rect 5056 5607 5063 5633
rect 5073 5613 5087 5627
rect 5133 5633 5147 5647
rect 5136 5627 5143 5633
rect 4993 5593 5007 5607
rect 4996 5587 5003 5593
rect 4916 5463 4923 5553
rect 4896 5456 4923 5463
rect 4896 5447 4903 5456
rect 4936 5447 4943 5513
rect 4893 5433 4907 5447
rect 4876 5427 4883 5433
rect 4873 5413 4887 5427
rect 4933 5433 4947 5447
rect 4956 5403 4963 5453
rect 5016 5447 5023 5573
rect 4973 5403 4987 5407
rect 4956 5396 4987 5403
rect 4836 5303 4843 5353
rect 4816 5296 4843 5303
rect 4767 5196 4793 5203
rect 4767 5176 4803 5183
rect 4573 5133 4587 5147
rect 4476 5127 4483 5133
rect 4516 5123 4523 5133
rect 4576 5123 4583 5133
rect 4516 5116 4583 5123
rect 4313 4953 4327 4967
rect 4156 4707 4163 4733
rect 4196 4707 4203 4753
rect 4116 4687 4123 4693
rect 4093 4653 4107 4667
rect 4113 4673 4127 4687
rect 4173 4673 4187 4687
rect 4096 4607 4103 4653
rect 4096 4507 4103 4593
rect 4136 4527 4143 4673
rect 4176 4647 4183 4673
rect 4115 4436 4123 4516
rect 4115 4398 4123 4422
rect 3996 4227 4003 4313
rect 4056 4307 4063 4353
rect 4156 4327 4163 4473
rect 4176 4387 4183 4593
rect 4216 4467 4223 4893
rect 4236 4707 4243 4933
rect 4293 4913 4307 4927
rect 4296 4903 4303 4913
rect 4276 4896 4303 4903
rect 4256 4827 4263 4893
rect 4276 4767 4283 4896
rect 4316 4847 4323 4913
rect 4336 4847 4343 5033
rect 4356 5007 4363 5033
rect 4356 4807 4363 4893
rect 4396 4807 4403 4933
rect 4416 4887 4423 5013
rect 4436 4967 4443 5113
rect 4476 5087 4483 5113
rect 4496 5016 4543 5023
rect 4496 5003 4503 5016
rect 4476 4996 4503 5003
rect 4476 4983 4483 4996
rect 4456 4976 4483 4983
rect 4456 4967 4463 4976
rect 4453 4953 4467 4967
rect 4516 4947 4523 4993
rect 4513 4933 4527 4947
rect 4476 4867 4483 4933
rect 4536 4927 4543 5016
rect 4596 4967 4603 5133
rect 4616 5007 4623 5133
rect 4653 4963 4667 4967
rect 4533 4913 4547 4927
rect 4633 4933 4647 4947
rect 4653 4956 4673 4963
rect 4653 4953 4667 4956
rect 4573 4913 4587 4927
rect 4257 4718 4265 4742
rect 4257 4624 4265 4704
rect 4276 4607 4283 4693
rect 4296 4667 4303 4733
rect 4313 4653 4327 4667
rect 4353 4653 4367 4667
rect 4316 4643 4323 4653
rect 4316 4636 4343 4643
rect 4193 4433 4207 4447
rect 4213 4453 4227 4467
rect 4236 4447 4243 4473
rect 4256 4467 4263 4513
rect 4276 4487 4283 4493
rect 4316 4487 4323 4593
rect 4336 4487 4343 4636
rect 4356 4607 4363 4653
rect 4376 4567 4383 4733
rect 4396 4624 4404 4736
rect 4416 4667 4423 4813
rect 4496 4727 4503 4913
rect 4576 4867 4583 4913
rect 4596 4767 4603 4933
rect 4636 4923 4643 4933
rect 4636 4916 4663 4923
rect 4636 4827 4643 4873
rect 4656 4847 4663 4916
rect 4676 4767 4683 4873
rect 4696 4827 4703 5133
rect 4716 4927 4723 4973
rect 4736 4963 4743 5133
rect 4796 5143 4803 5176
rect 4816 5167 4823 5296
rect 4856 5283 4863 5333
rect 4836 5276 4863 5283
rect 4836 5187 4843 5276
rect 4896 5267 4903 5393
rect 4916 5347 4923 5393
rect 4956 5343 4963 5396
rect 4973 5393 4987 5396
rect 5013 5393 5027 5407
rect 4936 5336 4963 5343
rect 4936 5307 4943 5336
rect 4976 5227 4983 5373
rect 5016 5347 5023 5393
rect 4833 5173 4847 5187
rect 4873 5173 4887 5187
rect 4876 5167 4883 5173
rect 4936 5167 4943 5193
rect 4853 5153 4867 5167
rect 4893 5153 4907 5167
rect 4856 5143 4863 5153
rect 4796 5136 4863 5143
rect 4753 5113 4767 5127
rect 4756 4987 4763 5113
rect 4776 4963 4783 5113
rect 4796 4987 4803 5113
rect 4816 5107 4823 5113
rect 4836 4967 4843 5093
rect 4876 5083 4883 5133
rect 4896 5103 4903 5153
rect 4933 5153 4947 5167
rect 4973 5163 4987 5167
rect 4996 5163 5003 5293
rect 5016 5287 5023 5333
rect 5036 5327 5043 5473
rect 5056 5447 5063 5553
rect 5076 5527 5083 5613
rect 5053 5433 5067 5447
rect 5096 5367 5103 5593
rect 5136 5447 5143 5613
rect 5156 5607 5163 5793
rect 5176 5707 5183 5873
rect 5236 5807 5243 5873
rect 5316 5867 5323 5896
rect 5353 5893 5367 5907
rect 5373 5913 5387 5927
rect 5413 5923 5427 5927
rect 5413 5916 5443 5923
rect 5413 5913 5427 5916
rect 5356 5887 5363 5893
rect 5276 5747 5283 5813
rect 5236 5676 5253 5683
rect 5236 5667 5243 5676
rect 5276 5667 5283 5733
rect 5316 5667 5323 5753
rect 5213 5633 5227 5647
rect 5233 5653 5247 5667
rect 5273 5653 5287 5667
rect 5216 5627 5223 5633
rect 5176 5467 5183 5593
rect 5156 5427 5163 5433
rect 5133 5403 5147 5407
rect 5116 5396 5147 5403
rect 5153 5413 5167 5427
rect 5036 5263 5043 5273
rect 5076 5267 5083 5353
rect 5016 5256 5043 5263
rect 5016 5207 5023 5256
rect 5036 5183 5043 5233
rect 5016 5176 5043 5183
rect 5016 5167 5023 5176
rect 4973 5156 5003 5163
rect 4973 5153 4987 5156
rect 4953 5133 4967 5147
rect 4956 5123 4963 5133
rect 4936 5116 4963 5123
rect 4936 5103 4943 5116
rect 4896 5096 4943 5103
rect 4876 5076 4903 5083
rect 4876 5063 4883 5076
rect 4856 5056 4883 5063
rect 4736 4956 4763 4963
rect 4776 4956 4803 4963
rect 4756 4947 4763 4956
rect 4753 4933 4767 4947
rect 4716 4847 4723 4893
rect 4736 4887 4743 4893
rect 4476 4707 4483 4713
rect 4473 4693 4487 4707
rect 4456 4607 4463 4693
rect 4493 4673 4507 4687
rect 4616 4687 4623 4733
rect 4533 4673 4547 4687
rect 4573 4683 4587 4687
rect 4573 4676 4603 4683
rect 4573 4673 4587 4676
rect 4496 4647 4503 4673
rect 4536 4667 4543 4673
rect 4553 4633 4567 4647
rect 4596 4643 4603 4676
rect 4613 4673 4627 4687
rect 4587 4636 4603 4643
rect 4556 4587 4563 4633
rect 4273 4473 4287 4487
rect 4253 4453 4267 4467
rect 4313 4473 4327 4487
rect 4333 4463 4347 4467
rect 4333 4456 4363 4463
rect 4333 4453 4347 4456
rect 4233 4433 4247 4447
rect 4196 4407 4203 4433
rect 4276 4407 4283 4433
rect 3853 4213 3867 4227
rect 3893 4223 3907 4227
rect 3953 4223 3967 4227
rect 3873 4193 3887 4207
rect 3893 4216 3923 4223
rect 3893 4213 3907 4216
rect 3876 4147 3883 4193
rect 3916 4147 3923 4216
rect 3936 4216 3967 4223
rect 3936 4067 3943 4216
rect 3953 4213 3967 4216
rect 3973 4193 3987 4207
rect 3993 4213 4007 4227
rect 3976 4187 3983 4193
rect 4056 4167 4063 4233
rect 4136 4207 4143 4253
rect 4093 4193 4107 4207
rect 4013 4153 4027 4167
rect 4016 4147 4023 4153
rect 3875 3956 3883 4036
rect 3893 4003 3907 4007
rect 3916 4003 3923 4053
rect 3893 3996 3923 4003
rect 3893 3993 3907 3996
rect 3953 3953 3967 3967
rect 3996 3967 4003 3993
rect 4016 3987 4023 4013
rect 4076 4003 4083 4193
rect 4096 4187 4103 4193
rect 4113 4173 4127 4187
rect 4133 4193 4147 4207
rect 4153 4173 4167 4187
rect 4173 4173 4187 4187
rect 4233 4193 4247 4207
rect 4116 4127 4123 4173
rect 4096 4027 4103 4033
rect 4076 3996 4103 4003
rect 4013 3973 4027 3987
rect 3993 3953 4007 3967
rect 4033 3953 4047 3967
rect 4073 3953 4087 3967
rect 3536 3727 3543 3773
rect 3655 3758 3663 3782
rect 3553 3693 3567 3707
rect 3593 3693 3607 3707
rect 3556 3627 3563 3693
rect 3655 3664 3663 3744
rect 3676 3707 3683 3753
rect 3673 3693 3687 3707
rect 3716 3627 3723 3793
rect 3796 3767 3803 3933
rect 3875 3918 3883 3942
rect 3956 3927 3963 3953
rect 4036 3927 4043 3953
rect 4076 3947 4083 3953
rect 4096 3927 4103 3996
rect 4116 3867 4123 4013
rect 4136 3987 4143 4133
rect 4156 4027 4163 4173
rect 4176 4147 4183 4173
rect 4216 4087 4223 4153
rect 4216 4007 4223 4073
rect 4236 4067 4243 4193
rect 4256 4187 4263 4373
rect 4276 4207 4283 4233
rect 4236 4027 4243 4033
rect 4233 4013 4247 4027
rect 4193 4003 4207 4007
rect 4213 4003 4227 4007
rect 4133 3973 4147 3987
rect 4193 3996 4227 4003
rect 4193 3993 4207 3996
rect 4213 3993 4227 3996
rect 3773 3743 3787 3747
rect 3773 3736 3803 3743
rect 3773 3733 3787 3736
rect 3436 3367 3443 3373
rect 3313 3213 3327 3227
rect 3333 3233 3347 3247
rect 3296 3143 3303 3213
rect 3336 3147 3343 3153
rect 3296 3136 3323 3143
rect 3156 3047 3163 3093
rect 2873 3033 2887 3047
rect 2793 3013 2807 3027
rect 2913 3033 2927 3047
rect 2953 3033 2967 3047
rect 3213 3043 3227 3047
rect 3207 3036 3227 3043
rect 3213 3033 3227 3036
rect 2796 3007 2803 3013
rect 2776 2663 2783 2973
rect 2795 2798 2803 2822
rect 2795 2704 2803 2784
rect 2816 2747 2823 2873
rect 2876 2787 2883 2993
rect 2896 2787 2903 2853
rect 2916 2827 2923 2853
rect 2936 2787 2943 2973
rect 2976 2847 2983 3033
rect 2996 2807 3003 3013
rect 3013 2993 3027 3007
rect 3016 2987 3023 2993
rect 3096 2987 3103 3033
rect 3153 2993 3167 3007
rect 3296 3027 3303 3093
rect 3316 3043 3323 3136
rect 3336 3067 3343 3133
rect 3356 3047 3363 3213
rect 3373 3193 3387 3207
rect 3416 3203 3423 3273
rect 3516 3223 3523 3453
rect 3536 3444 3544 3556
rect 3656 3527 3663 3553
rect 3576 3407 3583 3513
rect 3633 3493 3647 3507
rect 3653 3513 3667 3527
rect 3693 3523 3707 3527
rect 3716 3523 3723 3593
rect 3693 3516 3723 3523
rect 3693 3513 3707 3516
rect 3636 3467 3643 3493
rect 3696 3407 3703 3433
rect 3556 3247 3563 3253
rect 3576 3247 3583 3253
rect 3596 3247 3603 3293
rect 3716 3267 3723 3516
rect 3757 3476 3765 3556
rect 3776 3527 3783 3673
rect 3757 3438 3765 3462
rect 3737 3278 3745 3302
rect 3533 3223 3547 3227
rect 3516 3216 3547 3223
rect 3553 3233 3567 3247
rect 3593 3233 3607 3247
rect 3533 3213 3547 3216
rect 3633 3223 3647 3227
rect 3396 3196 3423 3203
rect 3376 3167 3383 3193
rect 3396 3167 3403 3196
rect 3573 3193 3587 3207
rect 3616 3216 3647 3223
rect 3456 3183 3463 3193
rect 3456 3176 3483 3183
rect 3476 3167 3483 3176
rect 3416 3087 3423 3133
rect 3456 3063 3463 3153
rect 3456 3056 3483 3063
rect 3316 3036 3343 3043
rect 3293 3013 3307 3027
rect 3336 3007 3343 3036
rect 3376 3027 3383 3053
rect 3476 3047 3483 3056
rect 3313 2993 3327 3007
rect 3353 2993 3367 3007
rect 3373 3013 3387 3027
rect 3473 3033 3487 3047
rect 3496 3027 3503 3093
rect 3516 3067 3523 3193
rect 3576 3163 3583 3193
rect 3556 3156 3583 3163
rect 3556 3147 3563 3156
rect 3536 3047 3543 3053
rect 3533 3033 3547 3047
rect 3493 3013 3507 3027
rect 3393 2993 3407 3007
rect 3156 2987 3163 2993
rect 3316 2987 3323 2993
rect 3356 2987 3363 2993
rect 3056 2927 3063 2953
rect 3076 2887 3083 2973
rect 3196 2947 3203 2953
rect 2956 2747 2963 2773
rect 2993 2763 3007 2767
rect 3016 2763 3023 2853
rect 3036 2767 3043 2813
rect 2973 2733 2987 2747
rect 2993 2756 3023 2763
rect 2993 2753 3007 2756
rect 3033 2753 3047 2767
rect 2776 2656 2843 2663
rect 2756 2607 2763 2633
rect 2776 2587 2783 2613
rect 2796 2587 2803 2633
rect 2816 2607 2823 2613
rect 2793 2573 2807 2587
rect 2693 2533 2707 2547
rect 2696 2527 2703 2533
rect 2756 2503 2763 2573
rect 2816 2567 2823 2593
rect 2836 2567 2843 2656
rect 2856 2567 2863 2713
rect 2876 2647 2883 2713
rect 2896 2647 2903 2693
rect 2813 2553 2827 2567
rect 2853 2553 2867 2567
rect 2716 2496 2763 2503
rect 2696 2423 2703 2493
rect 2716 2427 2723 2496
rect 2676 2416 2703 2423
rect 2656 2327 2663 2373
rect 2607 2296 2623 2303
rect 2533 2273 2547 2287
rect 2573 2283 2587 2287
rect 2573 2276 2593 2283
rect 2573 2273 2587 2276
rect 2633 2283 2647 2287
rect 2656 2283 2663 2293
rect 2676 2287 2683 2416
rect 2696 2307 2703 2393
rect 2776 2327 2783 2513
rect 2836 2487 2843 2553
rect 2516 2207 2523 2213
rect 2516 2167 2523 2193
rect 2516 2123 2523 2153
rect 2536 2147 2543 2273
rect 2613 2253 2627 2267
rect 2633 2276 2663 2283
rect 2633 2273 2647 2276
rect 2516 2116 2543 2123
rect 2513 2103 2527 2107
rect 2476 2096 2527 2103
rect 2476 2087 2483 2096
rect 2513 2093 2527 2096
rect 2433 2073 2447 2087
rect 2453 2053 2467 2067
rect 2473 2073 2487 2087
rect 2536 2087 2543 2116
rect 2533 2073 2547 2087
rect 2396 2016 2423 2023
rect 2396 1967 2403 1993
rect 2376 1936 2403 1943
rect 2296 1727 2303 1773
rect 2316 1647 2323 1833
rect 2376 1823 2383 1913
rect 2396 1903 2403 1936
rect 2416 1927 2423 2016
rect 2396 1896 2423 1903
rect 2356 1816 2383 1823
rect 2356 1807 2363 1816
rect 2396 1807 2403 1873
rect 2416 1823 2423 1896
rect 2436 1867 2443 2033
rect 2456 1887 2463 2053
rect 2416 1816 2443 1823
rect 2436 1807 2443 1816
rect 2333 1773 2347 1787
rect 2353 1793 2367 1807
rect 2393 1793 2407 1807
rect 2413 1773 2427 1787
rect 2336 1763 2343 1773
rect 2336 1756 2363 1763
rect 2356 1667 2363 1756
rect 2376 1683 2383 1753
rect 2416 1747 2423 1773
rect 2376 1676 2403 1683
rect 2113 1623 2127 1627
rect 2096 1616 2127 1623
rect 1993 1573 2007 1587
rect 2053 1573 2067 1587
rect 2073 1593 2087 1607
rect 2096 1587 2103 1616
rect 2113 1613 2127 1616
rect 2256 1607 2263 1613
rect 2173 1603 2187 1607
rect 2133 1583 2147 1587
rect 2156 1596 2187 1603
rect 2156 1583 2163 1596
rect 2133 1576 2163 1583
rect 2173 1593 2187 1596
rect 2133 1573 2147 1576
rect 2193 1573 2207 1587
rect 2253 1593 2267 1607
rect 2276 1603 2283 1633
rect 2313 1623 2327 1627
rect 2307 1616 2327 1623
rect 2313 1613 2327 1616
rect 2293 1603 2307 1607
rect 2276 1596 2307 1603
rect 1996 1547 2003 1573
rect 1856 1336 1873 1343
rect 1856 1327 1863 1336
rect 1833 1293 1847 1307
rect 1853 1313 1867 1327
rect 1873 1293 1887 1307
rect 1913 1303 1927 1307
rect 1936 1303 1943 1353
rect 1976 1347 1983 1473
rect 1996 1387 2003 1533
rect 2056 1467 2063 1573
rect 2056 1327 2063 1353
rect 2076 1327 2083 1373
rect 2156 1367 2163 1533
rect 2276 1527 2283 1596
rect 2293 1593 2307 1596
rect 2333 1593 2347 1607
rect 2176 1367 2183 1413
rect 2216 1367 2223 1453
rect 2236 1407 2243 1433
rect 2296 1427 2303 1513
rect 2116 1327 2123 1353
rect 2196 1347 2203 1353
rect 2236 1347 2243 1373
rect 2193 1333 2207 1347
rect 1913 1296 1943 1303
rect 1913 1293 1927 1296
rect 1836 1287 1843 1293
rect 1756 1147 1763 1193
rect 1753 1133 1767 1147
rect 1733 1113 1747 1127
rect 1776 1127 1783 1213
rect 1773 1113 1787 1127
rect 1796 1083 1803 1133
rect 1816 1127 1823 1193
rect 1836 1143 1843 1253
rect 1876 1167 1883 1293
rect 1836 1136 1863 1143
rect 1856 1127 1863 1136
rect 1896 1127 1903 1133
rect 1813 1113 1827 1127
rect 1853 1113 1867 1127
rect 1893 1113 1907 1127
rect 1796 1076 1843 1083
rect 1675 878 1683 902
rect 1613 823 1627 827
rect 1596 816 1627 823
rect 1596 787 1603 816
rect 1613 813 1627 816
rect 1675 784 1683 864
rect 1756 847 1763 853
rect 1796 847 1803 1053
rect 1836 947 1843 1076
rect 1876 1047 1883 1093
rect 1916 1087 1923 1153
rect 1936 1127 1943 1253
rect 1956 1207 1963 1313
rect 1993 1313 2007 1327
rect 2013 1293 2027 1307
rect 2053 1313 2067 1327
rect 2113 1313 2127 1327
rect 2133 1293 2147 1307
rect 2176 1303 2183 1333
rect 2233 1333 2247 1347
rect 2176 1296 2203 1303
rect 2033 1273 2047 1287
rect 1956 1127 1963 1153
rect 1996 1147 2003 1273
rect 1996 1127 2003 1133
rect 1953 1113 1967 1127
rect 1973 1093 1987 1107
rect 1993 1113 2007 1127
rect 2016 1083 2023 1273
rect 2036 1267 2043 1273
rect 2136 1243 2143 1293
rect 2116 1236 2143 1243
rect 2036 1147 2043 1193
rect 2056 1147 2063 1233
rect 2116 1223 2123 1236
rect 2096 1216 2123 1223
rect 2096 1167 2103 1216
rect 2116 1147 2123 1173
rect 2156 1163 2163 1293
rect 2136 1156 2163 1163
rect 2036 1107 2043 1133
rect 2096 1127 2103 1133
rect 2136 1127 2143 1156
rect 2093 1123 2107 1127
rect 1996 1076 2023 1083
rect 2033 1093 2047 1107
rect 2073 1093 2087 1107
rect 2093 1116 2123 1123
rect 2093 1113 2107 1116
rect 1876 867 1883 933
rect 1753 833 1767 847
rect 1793 833 1807 847
rect 1853 843 1867 847
rect 1813 813 1827 827
rect 1836 836 1867 843
rect 1816 807 1823 813
rect 1836 803 1843 836
rect 1853 833 1867 836
rect 1873 813 1887 827
rect 1896 823 1903 973
rect 1916 863 1923 933
rect 1916 856 1943 863
rect 1936 847 1943 856
rect 1913 823 1927 827
rect 1896 816 1927 823
rect 1933 833 1947 847
rect 1996 827 2003 1076
rect 2016 987 2023 993
rect 2036 987 2043 1033
rect 2016 867 2023 973
rect 2116 887 2123 1116
rect 2133 1113 2147 1127
rect 2176 1127 2183 1193
rect 2173 1113 2187 1127
rect 2196 1067 2203 1296
rect 2256 1207 2263 1393
rect 2296 1347 2303 1373
rect 2276 1327 2283 1333
rect 2273 1313 2287 1327
rect 2293 1293 2307 1307
rect 2296 1267 2303 1293
rect 2316 1267 2323 1433
rect 2336 1327 2343 1453
rect 2356 1447 2363 1613
rect 2333 1313 2347 1327
rect 2356 1203 2363 1293
rect 2376 1247 2383 1633
rect 2396 1627 2403 1676
rect 2476 1647 2483 1913
rect 2496 1827 2503 1953
rect 2536 1867 2543 2033
rect 2556 1967 2563 2253
rect 2576 1947 2583 2113
rect 2596 2087 2603 2253
rect 2616 2247 2623 2253
rect 2713 2273 2727 2287
rect 2753 2273 2767 2287
rect 2733 2253 2747 2267
rect 2696 2247 2703 2253
rect 2736 2227 2743 2253
rect 2616 2067 2623 2133
rect 2613 2053 2627 2067
rect 2636 2063 2643 2113
rect 2656 2087 2663 2153
rect 2696 2087 2703 2213
rect 2653 2063 2667 2067
rect 2636 2056 2667 2063
rect 2653 2053 2667 2056
rect 2693 2073 2707 2087
rect 2676 2043 2683 2053
rect 2676 2036 2703 2043
rect 2533 1773 2547 1787
rect 2513 1753 2527 1767
rect 2516 1667 2523 1753
rect 2536 1727 2543 1753
rect 2556 1627 2563 1713
rect 2576 1667 2583 1913
rect 2596 1787 2603 1993
rect 2617 1838 2625 1862
rect 2617 1744 2625 1824
rect 2636 1767 2643 1993
rect 2676 1967 2683 2013
rect 2573 1613 2587 1627
rect 2456 1607 2463 1613
rect 2393 1573 2407 1587
rect 2433 1573 2447 1587
rect 2453 1593 2467 1607
rect 2493 1603 2507 1607
rect 2476 1596 2507 1603
rect 2476 1547 2483 1596
rect 2493 1593 2507 1596
rect 2533 1593 2547 1607
rect 2596 1607 2603 1733
rect 2593 1593 2607 1607
rect 2396 1287 2403 1333
rect 2356 1196 2383 1203
rect 2216 1127 2223 1133
rect 2213 1113 2227 1127
rect 2233 1093 2247 1107
rect 2273 1093 2287 1107
rect 2236 987 2243 1093
rect 2276 1047 2283 1093
rect 2316 1087 2323 1133
rect 2137 878 2145 902
rect 2013 853 2027 867
rect 2053 863 2067 867
rect 2053 856 2083 863
rect 2053 853 2067 856
rect 2076 843 2083 856
rect 2076 836 2103 843
rect 1913 813 1927 816
rect 2096 823 2103 836
rect 2113 823 2127 827
rect 2096 816 2127 823
rect 1836 796 1863 803
rect 1393 603 1407 607
rect 1376 596 1407 603
rect 1413 613 1427 627
rect 1393 593 1407 596
rect 1433 593 1447 607
rect 1396 367 1403 393
rect 1436 387 1443 593
rect 1456 367 1463 393
rect 1476 387 1483 633
rect 1516 564 1524 676
rect 1556 647 1563 653
rect 1596 647 1603 773
rect 1553 633 1567 647
rect 1593 633 1607 647
rect 1655 596 1663 676
rect 1673 643 1687 647
rect 1696 643 1703 673
rect 1673 636 1703 643
rect 1673 633 1687 636
rect 1536 523 1543 573
rect 1655 558 1663 582
rect 1516 516 1543 523
rect 1253 333 1267 347
rect 1333 333 1347 347
rect 1393 353 1407 367
rect 1216 227 1223 233
rect 1216 167 1223 213
rect 1256 207 1263 333
rect 1336 227 1343 333
rect 1433 333 1447 347
rect 1453 353 1467 367
rect 1493 353 1507 367
rect 1413 313 1427 327
rect 1113 116 1143 123
rect 1213 153 1227 167
rect 1113 113 1127 116
rect 996 -24 1003 13
rect 1076 -24 1083 113
rect 1276 84 1284 196
rect 1356 167 1363 173
rect 1353 153 1367 167
rect 1396 -17 1403 293
rect 1436 207 1443 333
rect 1496 327 1503 353
rect 1415 116 1423 196
rect 1516 187 1523 516
rect 1556 367 1563 373
rect 1616 367 1623 373
rect 1553 353 1567 367
rect 1593 333 1607 347
rect 1613 353 1627 367
rect 1653 353 1667 367
rect 1573 313 1587 327
rect 1433 163 1447 167
rect 1456 163 1463 173
rect 1433 156 1463 163
rect 1433 153 1447 156
rect 1536 167 1543 233
rect 1556 187 1563 313
rect 1596 227 1603 333
rect 1656 327 1663 353
rect 1676 347 1683 593
rect 1696 467 1703 636
rect 1756 564 1764 676
rect 1836 647 1843 773
rect 1856 747 1863 796
rect 1876 767 1883 813
rect 2096 807 2103 816
rect 2113 813 2127 816
rect 1833 643 1847 647
rect 1816 636 1847 643
rect 1573 113 1587 127
rect 1415 78 1423 102
rect 1576 -17 1583 113
rect 1596 107 1603 153
rect 1616 127 1623 313
rect 1736 304 1744 416
rect 1756 287 1763 413
rect 1816 383 1823 636
rect 1833 633 1847 636
rect 1895 596 1903 676
rect 1913 633 1927 647
rect 1895 558 1903 582
rect 1996 564 2004 676
rect 2076 647 2083 773
rect 2096 767 2103 793
rect 2137 784 2145 864
rect 2156 687 2163 973
rect 2033 643 2047 647
rect 2016 636 2047 643
rect 2016 607 2023 636
rect 2033 633 2047 636
rect 2073 633 2087 647
rect 2135 596 2143 676
rect 2153 633 2167 647
rect 1875 398 1883 422
rect 1816 376 1843 383
rect 1773 333 1787 347
rect 1813 343 1827 347
rect 1836 343 1843 376
rect 1813 336 1843 343
rect 1813 333 1827 336
rect 1776 287 1783 333
rect 1875 304 1883 384
rect 1896 347 1903 393
rect 2096 387 2103 593
rect 2135 558 2143 582
rect 2136 387 2143 393
rect 2176 387 2183 953
rect 2193 813 2207 827
rect 2233 823 2247 827
rect 2256 823 2263 853
rect 2233 816 2263 823
rect 2233 813 2247 816
rect 2196 787 2203 813
rect 2276 784 2284 896
rect 2196 387 2203 393
rect 2216 387 2223 773
rect 2236 564 2244 676
rect 2273 643 2287 647
rect 2256 636 2287 643
rect 2256 607 2263 636
rect 2273 633 2287 636
rect 2296 527 2303 913
rect 2336 907 2343 1193
rect 2356 1044 2364 1156
rect 2376 967 2383 1196
rect 2436 1147 2443 1213
rect 2396 1127 2403 1133
rect 2393 1113 2407 1127
rect 2433 1123 2447 1127
rect 2416 1116 2447 1123
rect 2416 1083 2423 1116
rect 2433 1113 2447 1116
rect 2396 1076 2423 1083
rect 2396 867 2403 1076
rect 2456 1027 2463 1413
rect 2496 1327 2503 1353
rect 2473 1293 2487 1307
rect 2493 1313 2507 1327
rect 2476 1287 2483 1293
rect 2476 1147 2483 1253
rect 2516 1187 2523 1533
rect 2576 1487 2583 1573
rect 2616 1407 2623 1693
rect 2656 1667 2663 1873
rect 2676 1823 2683 1953
rect 2696 1927 2703 2036
rect 2716 1827 2723 2133
rect 2756 2107 2763 2253
rect 2733 2053 2747 2067
rect 2736 1987 2743 2053
rect 2676 1816 2703 1823
rect 2673 1783 2687 1787
rect 2696 1783 2703 1816
rect 2673 1776 2703 1783
rect 2673 1773 2687 1776
rect 2713 1773 2727 1787
rect 2636 1367 2643 1653
rect 2676 1647 2683 1733
rect 2696 1627 2703 1753
rect 2716 1747 2723 1773
rect 2736 1727 2743 1873
rect 2776 1867 2783 2193
rect 2796 1907 2803 2453
rect 2896 2427 2903 2593
rect 2916 2567 2923 2733
rect 2913 2553 2927 2567
rect 2933 2533 2947 2547
rect 2936 2467 2943 2533
rect 2956 2527 2963 2673
rect 2976 2647 2983 2733
rect 3056 2687 3063 2813
rect 3097 2798 3105 2822
rect 3076 2747 3083 2773
rect 3073 2733 3087 2747
rect 3097 2704 3105 2784
rect 2996 2587 3003 2633
rect 3016 2576 3033 2583
rect 3016 2567 3023 2576
rect 2993 2533 3007 2547
rect 3013 2553 3027 2567
rect 3033 2533 3047 2547
rect 2996 2523 3003 2533
rect 3076 2527 3083 2653
rect 3116 2607 3123 2853
rect 3136 2623 3143 2793
rect 3153 2733 3167 2747
rect 3216 2747 3223 2953
rect 3193 2733 3207 2747
rect 3196 2707 3203 2733
rect 3216 2687 3223 2733
rect 3236 2704 3244 2816
rect 3256 2747 3263 2773
rect 3296 2767 3303 2953
rect 3316 2947 3323 2953
rect 3336 2843 3343 2933
rect 3327 2836 3343 2843
rect 3356 2783 3363 2953
rect 3396 2947 3403 2993
rect 3416 2807 3423 2993
rect 3596 2883 3603 2993
rect 3616 2987 3623 3216
rect 3633 3213 3647 3216
rect 3673 3213 3687 3227
rect 3676 3207 3683 3213
rect 3696 3207 3703 3253
rect 3716 3227 3723 3233
rect 3713 3213 3727 3227
rect 3737 3184 3745 3264
rect 3636 3067 3643 3073
rect 3556 2876 3603 2883
rect 3556 2847 3563 2876
rect 3336 2776 3363 2783
rect 3316 2703 3323 2713
rect 3296 2696 3323 2703
rect 3216 2627 3223 2653
rect 3136 2616 3163 2623
rect 3113 2573 3127 2587
rect 2996 2516 3023 2523
rect 2836 2356 2873 2363
rect 2836 2347 2843 2356
rect 2813 2253 2827 2267
rect 2833 2233 2847 2247
rect 2836 2227 2843 2233
rect 2876 2187 2883 2333
rect 2917 2318 2925 2342
rect 2896 2267 2903 2293
rect 2917 2224 2925 2304
rect 2936 2287 2943 2333
rect 2816 2087 2823 2113
rect 2916 2107 2923 2113
rect 2936 2107 2943 2233
rect 2956 2227 2963 2493
rect 2976 2307 2983 2393
rect 2973 2253 2987 2267
rect 2996 2147 3003 2373
rect 3016 2307 3023 2516
rect 3036 2227 3043 2433
rect 3056 2224 3064 2336
rect 3096 2323 3103 2433
rect 3076 2316 3103 2323
rect 3076 2307 3083 2316
rect 3116 2303 3123 2473
rect 3136 2367 3143 2593
rect 3156 2387 3163 2616
rect 3176 2484 3184 2596
rect 3236 2487 3243 2653
rect 3253 2553 3267 2567
rect 3176 2387 3183 2433
rect 3296 2403 3303 2696
rect 3336 2603 3343 2776
rect 3373 2753 3387 2767
rect 3393 2733 3407 2747
rect 3433 2733 3447 2747
rect 3356 2727 3363 2733
rect 3396 2723 3403 2733
rect 3376 2716 3403 2723
rect 3376 2707 3383 2716
rect 3436 2707 3443 2733
rect 3456 2707 3463 2753
rect 3473 2733 3487 2747
rect 3493 2753 3507 2767
rect 3533 2753 3547 2767
rect 3513 2733 3527 2747
rect 3336 2596 3363 2603
rect 3315 2516 3323 2596
rect 3333 2553 3347 2567
rect 3315 2478 3323 2502
rect 3296 2396 3323 2403
rect 3096 2296 3123 2303
rect 3096 2167 3103 2296
rect 3113 2253 3127 2267
rect 3133 2273 3147 2287
rect 3196 2263 3203 2273
rect 3176 2256 3203 2263
rect 3116 2207 3123 2253
rect 3176 2187 3183 2256
rect 2976 2107 2983 2113
rect 2913 2093 2927 2107
rect 3116 2103 3123 2133
rect 3136 2107 3143 2153
rect 3196 2107 3203 2193
rect 3216 2147 3223 2333
rect 3296 2287 3303 2373
rect 3316 2327 3323 2396
rect 3273 2253 3287 2267
rect 3293 2273 3307 2287
rect 3276 2227 3283 2253
rect 3336 2163 3343 2413
rect 3356 2307 3363 2596
rect 3376 2567 3383 2633
rect 3396 2587 3403 2693
rect 3416 2627 3423 2673
rect 3476 2627 3483 2733
rect 3516 2707 3523 2733
rect 3556 2707 3563 2793
rect 3576 2747 3583 2853
rect 3616 2767 3623 2953
rect 3636 2947 3643 3053
rect 3696 3047 3703 3093
rect 3736 3047 3743 3053
rect 3653 3033 3667 3047
rect 3673 3013 3687 3027
rect 3693 3033 3707 3047
rect 3713 3013 3727 3027
rect 3733 3033 3747 3047
rect 3756 3023 3763 3193
rect 3776 3067 3783 3273
rect 3796 3263 3803 3736
rect 3836 3727 3843 3793
rect 3956 3727 3963 3773
rect 3976 3747 3983 3853
rect 4296 3807 4303 4433
rect 4356 4423 4363 4456
rect 4336 4416 4363 4423
rect 4316 4144 4324 4256
rect 4336 4103 4343 4416
rect 4376 4347 4383 4493
rect 4396 4327 4403 4433
rect 4353 4173 4367 4187
rect 4356 4127 4363 4173
rect 4336 4096 4363 4103
rect 4336 4027 4343 4053
rect 4333 4013 4347 4027
rect 4356 3967 4363 4096
rect 4376 4027 4383 4313
rect 4393 4183 4407 4187
rect 4416 4183 4423 4413
rect 4456 4407 4463 4493
rect 4493 4453 4507 4467
rect 4556 4467 4563 4573
rect 4576 4507 4583 4513
rect 4496 4447 4503 4453
rect 4576 4447 4583 4493
rect 4596 4487 4603 4553
rect 4616 4487 4623 4613
rect 4596 4467 4603 4473
rect 4573 4433 4587 4447
rect 4613 4443 4627 4447
rect 4636 4443 4643 4493
rect 4613 4436 4643 4443
rect 4656 4443 4663 4713
rect 4676 4687 4683 4713
rect 4696 4687 4703 4693
rect 4716 4687 4723 4833
rect 4756 4807 4763 4873
rect 4796 4727 4803 4956
rect 4833 4913 4847 4927
rect 4816 4747 4823 4913
rect 4836 4907 4843 4913
rect 4856 4843 4863 5056
rect 4896 5047 4903 5076
rect 4876 4967 4883 5033
rect 4896 4987 4903 4993
rect 4847 4836 4863 4843
rect 4676 4627 4683 4673
rect 4793 4673 4807 4687
rect 4796 4667 4803 4673
rect 4773 4653 4787 4667
rect 4713 4633 4727 4647
rect 4696 4547 4703 4633
rect 4716 4627 4723 4633
rect 4696 4523 4703 4533
rect 4696 4516 4723 4523
rect 4716 4487 4723 4516
rect 4736 4507 4743 4633
rect 4756 4547 4763 4613
rect 4776 4607 4783 4653
rect 4756 4487 4763 4513
rect 4796 4507 4803 4633
rect 4673 4463 4687 4467
rect 4713 4473 4727 4487
rect 4673 4456 4703 4463
rect 4673 4453 4687 4456
rect 4656 4436 4683 4443
rect 4613 4433 4627 4436
rect 4393 4176 4423 4183
rect 4393 4173 4407 4176
rect 4373 3953 4387 3967
rect 4436 3967 4443 4333
rect 4455 4238 4463 4262
rect 4455 4144 4463 4224
rect 4476 4187 4483 4213
rect 4473 4173 4487 4187
rect 4516 4167 4523 4313
rect 4576 4207 4583 4353
rect 4533 4193 4547 4207
rect 4536 4163 4543 4193
rect 4573 4193 4587 4207
rect 4593 4173 4607 4187
rect 4596 4167 4603 4173
rect 4536 4156 4563 4163
rect 4476 4007 4483 4033
rect 4516 4007 4523 4153
rect 4473 3993 4487 4007
rect 4493 3973 4507 3987
rect 4513 3993 4527 4007
rect 4413 3953 4427 3967
rect 4496 3967 4503 3973
rect 3973 3733 3987 3747
rect 4013 3743 4027 3747
rect 3813 3693 3827 3707
rect 3833 3713 3847 3727
rect 3853 3693 3867 3707
rect 3893 3693 3907 3707
rect 4013 3736 4043 3743
rect 4013 3733 4027 3736
rect 3816 3683 3823 3693
rect 3816 3676 3843 3683
rect 3813 3513 3827 3527
rect 3836 3267 3843 3676
rect 3856 3527 3863 3693
rect 3896 3607 3903 3693
rect 3853 3513 3867 3527
rect 3896 3444 3904 3556
rect 3796 3256 3823 3263
rect 3793 3213 3807 3227
rect 3816 3063 3823 3256
rect 3833 3223 3847 3227
rect 3856 3223 3863 3253
rect 3833 3216 3863 3223
rect 3833 3213 3847 3216
rect 3876 3184 3884 3296
rect 3796 3056 3823 3063
rect 3773 3023 3787 3027
rect 3756 3016 3787 3023
rect 3773 3013 3787 3016
rect 3716 2947 3723 3013
rect 3656 2767 3663 2893
rect 3756 2887 3763 2993
rect 3593 2733 3607 2747
rect 3613 2753 3627 2767
rect 3633 2733 3647 2747
rect 3653 2753 3667 2767
rect 3673 2733 3687 2747
rect 3693 2733 3707 2747
rect 3713 2753 3727 2767
rect 3753 2753 3767 2767
rect 3596 2723 3603 2733
rect 3587 2716 3603 2723
rect 3596 2607 3603 2673
rect 3393 2573 3407 2587
rect 3373 2553 3387 2567
rect 3413 2553 3427 2567
rect 3376 2287 3383 2473
rect 3396 2427 3403 2533
rect 3436 2443 3443 2533
rect 3456 2507 3463 2553
rect 3473 2513 3487 2527
rect 3513 2513 3527 2527
rect 3476 2487 3483 2513
rect 3516 2507 3523 2513
rect 3416 2436 3443 2443
rect 3416 2267 3423 2436
rect 3456 2423 3463 2473
rect 3496 2427 3503 2493
rect 3436 2416 3463 2423
rect 3436 2287 3443 2416
rect 3476 2403 3483 2413
rect 3456 2396 3483 2403
rect 3456 2307 3463 2396
rect 3476 2287 3483 2333
rect 3536 2307 3543 2513
rect 3556 2387 3563 2513
rect 3576 2407 3583 2553
rect 3596 2547 3603 2573
rect 3616 2567 3623 2693
rect 3636 2607 3643 2733
rect 3656 2583 3663 2693
rect 3676 2587 3683 2713
rect 3696 2627 3703 2733
rect 3636 2576 3663 2583
rect 3636 2547 3643 2576
rect 3676 2547 3683 2553
rect 3593 2533 3607 2547
rect 3616 2527 3623 2533
rect 3613 2513 3627 2527
rect 3653 2513 3667 2527
rect 3716 2527 3723 2713
rect 3736 2547 3743 2693
rect 3756 2583 3763 2693
rect 3776 2607 3783 2973
rect 3796 2887 3803 3056
rect 3816 2827 3823 2973
rect 3856 2787 3863 3033
rect 3876 2964 3884 3076
rect 3896 3067 3903 3213
rect 3916 3107 3923 3613
rect 4036 3567 4043 3736
rect 4076 3727 4083 3733
rect 4053 3693 4067 3707
rect 4073 3713 4087 3727
rect 4056 3607 4063 3693
rect 3956 3483 3963 3553
rect 3996 3547 4003 3553
rect 3993 3533 4007 3547
rect 4016 3523 4023 3553
rect 4033 3523 4047 3527
rect 4016 3516 4047 3523
rect 4033 3513 4047 3516
rect 3996 3483 4003 3493
rect 3956 3476 4003 3483
rect 4057 3476 4065 3556
rect 4113 3513 4127 3527
rect 4057 3438 4065 3462
rect 3956 3307 3963 3413
rect 3956 3247 3963 3293
rect 4136 3247 4143 3493
rect 4176 3403 4183 3733
rect 4196 3664 4204 3776
rect 4273 3693 4287 3707
rect 4196 3444 4204 3556
rect 4296 3547 4303 3553
rect 4293 3533 4307 3547
rect 4316 3467 4323 3953
rect 4376 3947 4383 3953
rect 4416 3863 4423 3953
rect 4496 3907 4503 3953
rect 4416 3856 4433 3863
rect 4335 3758 4343 3782
rect 4335 3664 4343 3744
rect 4393 3743 4407 3747
rect 4376 3736 4407 3743
rect 4433 3743 4447 3747
rect 4376 3707 4383 3736
rect 4393 3733 4407 3736
rect 4433 3736 4463 3743
rect 4433 3733 4447 3736
rect 4456 3607 4463 3736
rect 4376 3527 4383 3553
rect 4333 3493 4347 3507
rect 4336 3487 4343 3493
rect 4176 3396 4203 3403
rect 3953 3233 3967 3247
rect 3973 3213 3987 3227
rect 3993 3233 4007 3247
rect 4013 3213 4027 3227
rect 3913 3043 3927 3047
rect 3896 3036 3927 3043
rect 3896 3003 3903 3036
rect 3913 3033 3927 3036
rect 3936 3003 3943 3193
rect 3976 3107 3983 3213
rect 4016 3207 4023 3213
rect 4056 3107 4063 3233
rect 4073 3213 4087 3227
rect 4133 3233 4147 3247
rect 4153 3223 4167 3227
rect 4176 3223 4183 3233
rect 4153 3216 4183 3223
rect 4153 3213 4167 3216
rect 4076 3207 4083 3213
rect 4196 3203 4203 3396
rect 4356 3343 4363 3493
rect 4373 3473 4387 3487
rect 4413 3473 4427 3487
rect 4376 3467 4383 3473
rect 4416 3387 4423 3473
rect 4476 3467 4483 3753
rect 4536 3747 4543 3753
rect 4556 3747 4563 4156
rect 4576 3924 4584 4036
rect 4616 4007 4623 4033
rect 4613 3993 4627 4007
rect 4636 4003 4643 4413
rect 4676 4267 4683 4436
rect 4696 4327 4703 4456
rect 4733 4453 4747 4467
rect 4753 4473 4767 4487
rect 4776 4467 4783 4473
rect 4773 4453 4787 4467
rect 4716 4407 4723 4433
rect 4736 4387 4743 4453
rect 4656 4144 4664 4256
rect 4676 4007 4683 4233
rect 4756 4227 4763 4433
rect 4776 4287 4783 4373
rect 4796 4347 4803 4493
rect 4733 4183 4747 4187
rect 4733 4176 4763 4183
rect 4733 4173 4747 4176
rect 4653 4003 4667 4007
rect 4636 3996 4667 4003
rect 4653 3993 4667 3996
rect 4715 3956 4723 4036
rect 4715 3918 4723 3942
rect 4596 3767 4603 3793
rect 4533 3733 4547 3747
rect 4573 3713 4587 3727
rect 4476 3367 4483 3453
rect 4496 3444 4504 3556
rect 4533 3523 4547 3527
rect 4573 3523 4587 3527
rect 4596 3523 4603 3753
rect 4716 3747 4723 3873
rect 4716 3727 4723 3733
rect 4713 3713 4727 3727
rect 4533 3516 4563 3523
rect 4533 3513 4547 3516
rect 4356 3336 4383 3343
rect 4176 3196 4203 3203
rect 3953 3033 3967 3047
rect 3896 2996 3923 3003
rect 3936 2996 3963 3003
rect 3916 2787 3923 2996
rect 3756 2576 3783 2583
rect 3733 2533 3747 2547
rect 3753 2513 3767 2527
rect 3433 2273 3447 2287
rect 3393 2253 3407 2267
rect 3373 2233 3387 2247
rect 3376 2203 3383 2233
rect 3356 2196 3383 2203
rect 3356 2187 3363 2196
rect 3336 2156 3363 2163
rect 3096 2096 3123 2103
rect 2813 2073 2827 2087
rect 2756 1744 2764 1856
rect 2816 1843 2823 1953
rect 2856 1947 2863 2093
rect 2893 2053 2907 2067
rect 2933 2063 2947 2067
rect 2927 2056 2947 2063
rect 2933 2053 2947 2056
rect 2993 2053 3007 2067
rect 3033 2053 3047 2067
rect 3053 2073 3067 2087
rect 2836 1887 2843 1913
rect 2876 1847 2883 1973
rect 2896 1907 2903 2053
rect 2956 2027 2963 2053
rect 2996 2027 3003 2053
rect 3036 2007 3043 2053
rect 2796 1836 2823 1843
rect 2776 1727 2783 1833
rect 2796 1767 2803 1836
rect 2873 1823 2887 1827
rect 2813 1793 2827 1807
rect 2873 1816 2903 1823
rect 2873 1813 2887 1816
rect 2896 1803 2903 1816
rect 2976 1807 2983 1873
rect 3036 1807 3043 1933
rect 3056 1847 3063 2033
rect 3096 1967 3103 2096
rect 3153 2093 3167 2107
rect 3193 2093 3207 2107
rect 3296 2087 3303 2133
rect 3336 2087 3343 2133
rect 3356 2087 3363 2156
rect 3376 2087 3383 2153
rect 3396 2107 3403 2133
rect 3393 2093 3407 2107
rect 3416 2103 3423 2233
rect 3416 2096 3443 2103
rect 3253 2083 3267 2087
rect 3173 2053 3187 2067
rect 3213 2063 3227 2067
rect 3236 2076 3267 2083
rect 3236 2063 3243 2076
rect 3213 2056 3243 2063
rect 3253 2073 3267 2076
rect 3213 2053 3227 2056
rect 3273 2053 3287 2067
rect 3293 2073 3307 2087
rect 3333 2073 3347 2087
rect 3373 2073 3387 2087
rect 3413 2073 3427 2087
rect 3156 2043 3163 2053
rect 3136 2036 3163 2043
rect 3116 1967 3123 2013
rect 2933 1803 2947 1807
rect 2896 1796 2947 1803
rect 2933 1793 2947 1796
rect 2816 1787 2823 1793
rect 2973 1793 2987 1807
rect 3013 1773 3027 1787
rect 2896 1747 2903 1773
rect 2776 1623 2783 1693
rect 2776 1616 2803 1623
rect 2676 1587 2683 1593
rect 2736 1587 2743 1613
rect 2653 1553 2667 1567
rect 2673 1573 2687 1587
rect 2693 1553 2707 1567
rect 2713 1553 2727 1567
rect 2733 1573 2747 1587
rect 2753 1553 2767 1567
rect 2696 1543 2703 1553
rect 2776 1543 2783 1593
rect 2796 1567 2803 1616
rect 2816 1607 2823 1673
rect 2813 1593 2827 1607
rect 2833 1573 2847 1587
rect 2836 1563 2843 1573
rect 2816 1556 2843 1563
rect 2696 1536 2723 1543
rect 2596 1327 2603 1333
rect 2656 1327 2663 1413
rect 2716 1367 2723 1536
rect 2736 1536 2783 1543
rect 2736 1327 2743 1536
rect 2816 1543 2823 1556
rect 2807 1536 2823 1543
rect 2856 1527 2863 1613
rect 2876 1607 2883 1693
rect 2873 1593 2887 1607
rect 2893 1583 2907 1587
rect 2916 1583 2923 1633
rect 2956 1603 2963 1753
rect 2976 1707 2983 1753
rect 3016 1727 3023 1773
rect 3033 1753 3047 1767
rect 2956 1596 2983 1603
rect 2893 1576 2923 1583
rect 2893 1573 2907 1576
rect 2933 1553 2947 1567
rect 2953 1573 2967 1587
rect 2976 1567 2983 1596
rect 2993 1573 3007 1587
rect 2973 1553 2987 1567
rect 2553 1313 2567 1327
rect 2573 1293 2587 1307
rect 2593 1313 2607 1327
rect 2613 1303 2627 1307
rect 2633 1303 2647 1307
rect 2613 1296 2647 1303
rect 2653 1313 2667 1327
rect 2613 1293 2627 1296
rect 2633 1293 2647 1296
rect 2673 1293 2687 1307
rect 2693 1313 2707 1327
rect 2556 1247 2563 1273
rect 2576 1247 2583 1293
rect 2636 1283 2643 1293
rect 2636 1276 2663 1283
rect 2436 967 2443 1013
rect 2476 927 2483 1113
rect 2495 1076 2503 1156
rect 2495 1038 2503 1062
rect 2516 1007 2523 1093
rect 2536 987 2543 1193
rect 2416 867 2423 913
rect 2416 847 2423 853
rect 2376 787 2383 833
rect 2413 833 2427 847
rect 2433 813 2447 827
rect 2473 813 2487 827
rect 2436 807 2443 813
rect 2316 647 2323 773
rect 2476 767 2483 813
rect 2496 687 2503 893
rect 2536 847 2543 913
rect 2556 907 2563 1173
rect 2656 1143 2663 1276
rect 2676 1163 2683 1293
rect 2676 1156 2703 1163
rect 2656 1136 2683 1143
rect 2676 1127 2683 1136
rect 2576 1087 2583 1093
rect 2616 887 2623 1033
rect 2656 1027 2663 1073
rect 2553 813 2567 827
rect 2556 807 2563 813
rect 2516 707 2523 713
rect 2313 633 2327 647
rect 2375 596 2383 676
rect 2393 633 2407 647
rect 2396 607 2403 633
rect 1953 363 1967 367
rect 1936 356 1967 363
rect 1893 333 1907 347
rect 1696 167 1703 193
rect 1716 187 1723 273
rect 1713 173 1727 187
rect 1693 153 1707 167
rect 1756 123 1763 193
rect 1796 147 1803 173
rect 1773 123 1787 127
rect 1756 116 1787 123
rect 1793 133 1807 147
rect 1773 113 1787 116
rect 1813 113 1827 127
rect 1836 123 1843 193
rect 1853 123 1867 127
rect 1836 116 1867 123
rect 1853 113 1867 116
rect 1893 113 1907 127
rect 1916 123 1923 193
rect 1936 167 1943 356
rect 1953 353 1967 356
rect 1973 313 1987 327
rect 2053 333 2067 347
rect 2113 353 2127 367
rect 2033 313 2047 327
rect 1976 187 1983 313
rect 2036 307 2043 313
rect 2056 227 2063 333
rect 2096 167 2103 213
rect 1933 123 1947 127
rect 1916 116 1947 123
rect 2016 127 2023 153
rect 2073 133 2087 147
rect 2093 153 2107 167
rect 1933 113 1947 116
rect 1973 113 1987 127
rect 2076 127 2083 133
rect 1816 -17 1823 113
rect 1896 -17 1903 113
rect 1976 -17 1983 113
rect 2116 107 2123 353
rect 2136 323 2143 373
rect 2236 367 2243 513
rect 2153 323 2167 327
rect 2136 316 2167 323
rect 2196 323 2203 353
rect 2253 333 2267 347
rect 2196 316 2223 323
rect 2153 313 2167 316
rect 2196 247 2203 293
rect 2156 84 2164 196
rect 2216 163 2223 316
rect 2256 287 2263 333
rect 2296 267 2303 313
rect 2316 307 2323 593
rect 2477 596 2485 676
rect 2496 647 2503 673
rect 2375 558 2383 582
rect 2477 558 2485 582
rect 2396 367 2403 373
rect 2353 353 2367 367
rect 2356 327 2363 353
rect 2373 333 2387 347
rect 2393 353 2407 367
rect 2413 333 2427 347
rect 2473 343 2487 347
rect 2496 343 2503 473
rect 2516 347 2523 693
rect 2536 647 2543 773
rect 2533 633 2547 647
rect 2556 487 2563 793
rect 2576 767 2583 813
rect 2576 647 2583 693
rect 2573 633 2587 647
rect 2596 603 2603 873
rect 2673 813 2687 827
rect 2676 787 2683 813
rect 2576 596 2603 603
rect 2236 167 2243 173
rect 2233 163 2247 167
rect 2216 156 2247 163
rect 2233 153 2247 156
rect 2295 116 2303 196
rect 2336 167 2343 293
rect 2376 247 2383 333
rect 2473 336 2503 343
rect 2473 333 2487 336
rect 2453 313 2467 327
rect 2356 167 2363 213
rect 2295 78 2303 102
rect 2336 87 2343 153
rect 2393 113 2407 127
rect 2396 -17 2403 113
rect 2416 107 2423 133
rect 2436 107 2443 313
rect 2456 267 2463 313
rect 2556 304 2564 416
rect 2453 113 2467 127
rect 2493 123 2507 127
rect 2516 123 2523 213
rect 2576 207 2583 596
rect 2616 564 2624 676
rect 2636 667 2643 773
rect 2636 423 2643 653
rect 2616 416 2643 423
rect 2593 333 2607 347
rect 2596 267 2603 333
rect 2616 307 2623 416
rect 2633 343 2647 347
rect 2656 343 2663 753
rect 2633 336 2663 343
rect 2633 333 2647 336
rect 2656 307 2663 336
rect 2676 327 2683 673
rect 2696 647 2703 1156
rect 2716 967 2723 1273
rect 2736 1207 2743 1313
rect 2756 1167 2763 1413
rect 2856 1343 2863 1413
rect 2836 1336 2863 1343
rect 2836 1327 2843 1336
rect 2773 1293 2787 1307
rect 2793 1313 2807 1327
rect 2813 1293 2827 1307
rect 2833 1313 2847 1327
rect 2853 1293 2867 1307
rect 2873 1293 2887 1307
rect 2776 1287 2783 1293
rect 2816 1287 2823 1293
rect 2856 1247 2863 1293
rect 2776 1203 2783 1213
rect 2776 1196 2803 1203
rect 2776 1127 2783 1173
rect 2796 1147 2803 1196
rect 2816 1147 2823 1233
rect 2793 1133 2807 1147
rect 2733 1123 2747 1127
rect 2733 1116 2763 1123
rect 2733 1113 2747 1116
rect 2736 1027 2743 1073
rect 2756 1067 2763 1116
rect 2773 1113 2787 1127
rect 2813 1093 2827 1107
rect 2713 843 2727 847
rect 2713 836 2743 843
rect 2713 833 2727 836
rect 2736 767 2743 836
rect 2756 767 2763 913
rect 2776 727 2783 1073
rect 2796 967 2803 1093
rect 2816 1067 2823 1093
rect 2836 1047 2843 1153
rect 2856 1003 2863 1193
rect 2896 1183 2903 1493
rect 2956 1407 2963 1533
rect 3016 1487 3023 1713
rect 3036 1707 3043 1753
rect 3036 1647 3043 1673
rect 3056 1647 3063 1773
rect 3076 1727 3083 1873
rect 3136 1827 3143 2036
rect 3133 1803 3147 1807
rect 3156 1803 3163 1873
rect 3176 1827 3183 2033
rect 3113 1773 3127 1787
rect 3133 1796 3163 1803
rect 3133 1793 3147 1796
rect 3116 1743 3123 1773
rect 3196 1767 3203 1913
rect 3236 1887 3243 2033
rect 3236 1807 3243 1873
rect 3213 1773 3227 1787
rect 3233 1793 3247 1807
rect 3153 1753 3167 1767
rect 3096 1736 3123 1743
rect 3096 1667 3103 1736
rect 3136 1723 3143 1733
rect 3116 1716 3143 1723
rect 3116 1687 3123 1716
rect 3036 1607 3043 1633
rect 3033 1593 3047 1607
rect 3053 1573 3067 1587
rect 3056 1447 3063 1553
rect 3116 1524 3124 1636
rect 3136 1443 3143 1693
rect 3156 1607 3163 1673
rect 3176 1663 3183 1753
rect 3216 1727 3223 1773
rect 3296 1707 3303 1873
rect 3316 1827 3323 1933
rect 3313 1773 3327 1787
rect 3316 1767 3323 1773
rect 3336 1747 3343 1993
rect 3396 1987 3403 2053
rect 3436 2027 3443 2096
rect 3456 1907 3463 2073
rect 3476 2047 3483 2273
rect 3533 2253 3547 2267
rect 3513 2233 3527 2247
rect 3496 2167 3503 2233
rect 3536 2167 3543 2253
rect 3496 2004 3504 2116
rect 3536 2087 3543 2113
rect 3533 2073 3547 2087
rect 3556 1967 3563 2333
rect 3576 2207 3583 2393
rect 3596 2387 3603 2473
rect 3656 2423 3663 2513
rect 3676 2487 3683 2513
rect 3776 2487 3783 2576
rect 3796 2547 3803 2773
rect 3956 2767 3963 2996
rect 3976 2787 3983 3013
rect 4015 2996 4023 3076
rect 4073 3043 4087 3047
rect 4056 3036 4087 3043
rect 4015 2958 4023 2982
rect 3996 2827 4003 2953
rect 4036 2923 4043 3033
rect 4016 2916 4043 2923
rect 4016 2863 4023 2916
rect 4016 2856 4033 2863
rect 3996 2767 4003 2793
rect 4016 2787 4023 2833
rect 4056 2783 4063 3036
rect 4073 3033 4087 3036
rect 4093 3013 4107 3027
rect 4133 3023 4147 3027
rect 4133 3016 4163 3023
rect 4133 3013 4147 3016
rect 4076 2807 4083 2993
rect 4096 2787 4103 3013
rect 4156 3007 4163 3016
rect 4056 2776 4083 2783
rect 4076 2767 4083 2776
rect 3813 2733 3827 2747
rect 3853 2733 3867 2747
rect 3873 2753 3887 2767
rect 3816 2727 3823 2733
rect 3856 2723 3863 2733
rect 3856 2716 3893 2723
rect 3816 2567 3823 2633
rect 3836 2547 3843 2713
rect 3916 2707 3923 2733
rect 3973 2733 3987 2747
rect 3953 2723 3967 2727
rect 4013 2733 4027 2747
rect 4053 2733 4067 2747
rect 4093 2733 4107 2747
rect 3953 2716 3983 2723
rect 3953 2713 3967 2716
rect 3976 2703 3983 2716
rect 4016 2703 4023 2713
rect 3976 2696 4023 2703
rect 3936 2567 3943 2593
rect 3956 2567 3963 2693
rect 4096 2667 4103 2733
rect 4116 2727 4123 2953
rect 4176 2907 4183 3196
rect 4216 3184 4224 3296
rect 4236 3027 4243 3293
rect 4355 3278 4363 3302
rect 4293 3213 4307 3227
rect 4355 3184 4363 3264
rect 4376 3227 4383 3336
rect 4373 3213 4387 3227
rect 4396 3147 4403 3313
rect 4476 3267 4483 3313
rect 4516 3247 4523 3473
rect 4556 3327 4563 3516
rect 4573 3516 4603 3523
rect 4573 3513 4587 3516
rect 4616 3507 4623 3533
rect 4635 3476 4643 3556
rect 4736 3547 4743 3933
rect 4756 3767 4763 4176
rect 4776 3967 4783 4273
rect 4795 4238 4803 4262
rect 4816 4247 4823 4733
rect 4836 4703 4843 4793
rect 4876 4727 4883 4813
rect 4836 4696 4863 4703
rect 4856 4687 4863 4696
rect 4836 4607 4843 4653
rect 4896 4663 4903 4953
rect 4936 4947 4943 4993
rect 4976 4967 4983 5133
rect 4996 4947 5003 5156
rect 5013 5153 5027 5167
rect 5056 5123 5063 5253
rect 5076 5187 5083 5253
rect 5096 5207 5103 5313
rect 5116 5287 5123 5396
rect 5133 5393 5147 5396
rect 5173 5393 5187 5407
rect 5116 5187 5123 5213
rect 5073 5173 5087 5187
rect 5156 5167 5163 5253
rect 5176 5247 5183 5393
rect 5196 5223 5203 5613
rect 5256 5607 5263 5653
rect 5293 5633 5307 5647
rect 5313 5653 5327 5667
rect 5296 5623 5303 5633
rect 5336 5623 5343 5873
rect 5356 5727 5363 5873
rect 5436 5847 5443 5916
rect 5456 5867 5463 5933
rect 5496 5907 5503 5933
rect 5516 5927 5523 5936
rect 5533 5933 5547 5936
rect 5493 5893 5507 5907
rect 5513 5883 5527 5887
rect 5513 5876 5543 5883
rect 5513 5873 5527 5876
rect 5396 5687 5403 5713
rect 5416 5667 5423 5693
rect 5373 5653 5387 5667
rect 5353 5633 5367 5647
rect 5356 5627 5363 5633
rect 5276 5616 5303 5623
rect 5316 5616 5343 5623
rect 5216 5447 5223 5513
rect 5236 5467 5243 5533
rect 5256 5447 5263 5533
rect 5276 5527 5283 5616
rect 5316 5567 5323 5616
rect 5276 5476 5323 5483
rect 5276 5467 5283 5476
rect 5213 5433 5227 5447
rect 5233 5413 5247 5427
rect 5253 5433 5267 5447
rect 5236 5407 5243 5413
rect 5176 5216 5203 5223
rect 5153 5163 5167 5167
rect 5136 5156 5167 5163
rect 5036 5116 5063 5123
rect 5016 4967 5023 4993
rect 4913 4913 4927 4927
rect 4933 4933 4947 4947
rect 4953 4913 4967 4927
rect 4993 4933 5007 4947
rect 5013 4913 5027 4927
rect 4916 4907 4923 4913
rect 4956 4887 4963 4913
rect 4976 4887 4983 4913
rect 4996 4883 5003 4893
rect 5016 4883 5023 4913
rect 5036 4907 5043 5116
rect 5056 4967 5063 4973
rect 5053 4953 5067 4967
rect 5056 4887 5063 4913
rect 4996 4876 5023 4883
rect 4916 4727 4923 4873
rect 4996 4767 5003 4876
rect 4956 4727 4963 4753
rect 4916 4707 4923 4713
rect 4976 4707 4983 4733
rect 4996 4707 5003 4733
rect 5016 4723 5023 4813
rect 5036 4747 5043 4873
rect 5076 4827 5083 5093
rect 5096 5007 5103 5133
rect 5116 5047 5123 5133
rect 5096 4967 5103 4993
rect 5136 4987 5143 5156
rect 5153 5153 5167 5156
rect 5176 5123 5183 5216
rect 5196 5167 5203 5193
rect 5156 5116 5183 5123
rect 5113 4963 5127 4967
rect 5113 4956 5143 4963
rect 5113 4953 5127 4956
rect 5136 4927 5143 4956
rect 5096 4807 5103 4893
rect 5116 4847 5123 4893
rect 5156 4867 5163 5116
rect 5176 4987 5183 5013
rect 5196 4947 5203 4993
rect 5216 4987 5223 5333
rect 5256 5287 5263 5393
rect 5236 5187 5243 5253
rect 5256 5216 5273 5223
rect 5256 5207 5263 5216
rect 5276 5187 5283 5193
rect 5253 5153 5267 5167
rect 5273 5173 5287 5187
rect 5256 5123 5263 5153
rect 5256 5116 5283 5123
rect 5193 4933 5207 4947
rect 5236 4887 5243 5113
rect 5276 5107 5283 5116
rect 5276 4967 5283 5073
rect 5273 4913 5287 4927
rect 5196 4803 5203 4833
rect 5116 4796 5203 4803
rect 5116 4783 5123 4796
rect 5056 4776 5123 4783
rect 5156 4776 5223 4783
rect 5056 4747 5063 4776
rect 5016 4716 5063 4723
rect 5056 4707 5063 4716
rect 4933 4673 4947 4687
rect 4993 4693 5007 4707
rect 5013 4673 5027 4687
rect 4936 4667 4943 4673
rect 4896 4656 4923 4663
rect 4853 4633 4867 4647
rect 4856 4587 4863 4633
rect 4833 4453 4847 4467
rect 4836 4427 4843 4453
rect 4856 4443 4863 4533
rect 4876 4487 4883 4513
rect 4896 4507 4903 4533
rect 4873 4473 4887 4487
rect 4856 4436 4883 4443
rect 4856 4267 4863 4413
rect 4876 4267 4883 4436
rect 4896 4387 4903 4433
rect 4916 4287 4923 4656
rect 4976 4527 4983 4673
rect 5016 4663 5023 4673
rect 5076 4667 5083 4733
rect 5096 4727 5103 4753
rect 5156 4707 5163 4776
rect 5216 4767 5223 4776
rect 5176 4687 5183 4713
rect 5196 4707 5203 4753
rect 5236 4707 5243 4873
rect 5256 4767 5263 4913
rect 5276 4907 5283 4913
rect 5296 4867 5303 5453
rect 5316 5267 5323 5476
rect 5336 5447 5343 5573
rect 5356 5527 5363 5613
rect 5376 5607 5383 5653
rect 5413 5653 5427 5667
rect 5396 5547 5403 5633
rect 5396 5447 5403 5513
rect 5436 5487 5443 5753
rect 5496 5647 5503 5853
rect 5516 5667 5523 5813
rect 5536 5807 5543 5876
rect 5576 5867 5583 5913
rect 5596 5883 5603 6073
rect 5656 6047 5663 6133
rect 5716 6127 5723 6153
rect 5616 5967 5623 5993
rect 5636 5907 5643 5933
rect 5613 5883 5627 5887
rect 5596 5876 5627 5883
rect 5656 5887 5663 5913
rect 5676 5907 5683 5953
rect 5696 5947 5703 6073
rect 5736 5967 5743 6353
rect 5756 6267 5763 6376
rect 5773 6373 5787 6376
rect 5876 6367 5883 6393
rect 5953 6373 5967 6387
rect 5956 6367 5963 6373
rect 5833 6353 5847 6367
rect 5836 6347 5843 6353
rect 5816 6167 5823 6333
rect 5896 6147 5903 6233
rect 5753 6093 5767 6107
rect 5833 6113 5847 6127
rect 5756 6067 5763 6093
rect 5836 6107 5843 6113
rect 5856 6087 5863 6133
rect 5893 6133 5907 6147
rect 5716 5947 5723 5953
rect 5673 5893 5687 5907
rect 5733 5893 5747 5907
rect 5613 5873 5627 5876
rect 5736 5887 5743 5893
rect 5536 5607 5543 5773
rect 5576 5707 5583 5833
rect 5596 5687 5603 5853
rect 5556 5667 5563 5673
rect 5553 5653 5567 5667
rect 5573 5633 5587 5647
rect 5416 5447 5423 5453
rect 5456 5447 5463 5553
rect 5476 5447 5483 5533
rect 5393 5443 5407 5447
rect 5376 5436 5407 5443
rect 5376 5407 5383 5436
rect 5393 5433 5407 5436
rect 5413 5433 5427 5447
rect 5433 5413 5447 5427
rect 5453 5433 5467 5447
rect 5353 5393 5367 5407
rect 5336 5287 5343 5353
rect 5336 5187 5343 5273
rect 5356 5247 5363 5393
rect 5376 5207 5383 5253
rect 5313 5133 5327 5147
rect 5353 5133 5367 5147
rect 5316 5127 5323 5133
rect 5356 5127 5363 5133
rect 5376 5027 5383 5133
rect 5396 5007 5403 5353
rect 5436 5327 5443 5413
rect 5496 5367 5503 5593
rect 5576 5507 5583 5633
rect 5513 5393 5527 5407
rect 5516 5347 5523 5393
rect 5576 5387 5583 5453
rect 5596 5427 5603 5613
rect 5616 5467 5623 5793
rect 5636 5687 5643 5853
rect 5656 5687 5663 5693
rect 5756 5667 5763 5873
rect 5776 5847 5783 5933
rect 5796 5903 5803 6033
rect 5836 5927 5843 5953
rect 5876 5947 5883 6113
rect 5916 5987 5923 6353
rect 5976 6327 5983 6413
rect 6036 6387 6043 6416
rect 6056 6407 6063 6453
rect 6096 6427 6103 6433
rect 6093 6413 6107 6427
rect 6053 6393 6067 6407
rect 6073 6373 6087 6387
rect 6113 6383 6127 6387
rect 6096 6376 6127 6383
rect 6076 6367 6083 6373
rect 5956 6127 5963 6153
rect 5976 6147 5983 6313
rect 5933 6093 5947 6107
rect 5953 6113 5967 6127
rect 5936 6087 5943 6093
rect 5936 6067 5943 6073
rect 5936 5927 5943 5933
rect 5833 5913 5847 5927
rect 5813 5903 5827 5907
rect 5796 5896 5827 5903
rect 5796 5847 5803 5896
rect 5813 5893 5827 5896
rect 5853 5893 5867 5907
rect 5913 5893 5927 5907
rect 5933 5913 5947 5927
rect 5653 5663 5667 5667
rect 5636 5656 5667 5663
rect 5636 5587 5643 5656
rect 5653 5653 5667 5656
rect 5673 5633 5687 5647
rect 5636 5547 5643 5553
rect 5656 5547 5663 5593
rect 5656 5467 5663 5513
rect 5676 5507 5683 5633
rect 5753 5613 5767 5627
rect 5793 5613 5807 5627
rect 5696 5603 5703 5613
rect 5696 5596 5743 5603
rect 5736 5547 5743 5596
rect 5756 5587 5763 5613
rect 5593 5413 5607 5427
rect 5616 5407 5623 5433
rect 5676 5427 5683 5473
rect 5613 5393 5627 5407
rect 5653 5403 5667 5407
rect 5696 5403 5703 5513
rect 5716 5447 5723 5533
rect 5776 5507 5783 5593
rect 5796 5567 5803 5613
rect 5836 5587 5843 5833
rect 5856 5827 5863 5893
rect 5896 5707 5903 5833
rect 5916 5827 5923 5893
rect 5976 5867 5983 5933
rect 6016 5927 6023 6353
rect 6096 6327 6103 6376
rect 6113 6373 6127 6376
rect 6056 6127 6063 6153
rect 6033 6093 6047 6107
rect 6053 6113 6067 6127
rect 6093 6113 6107 6127
rect 6116 6123 6123 6333
rect 6136 6287 6143 6433
rect 6156 6407 6163 6453
rect 6176 6407 6183 6473
rect 6216 6407 6223 6433
rect 6173 6393 6187 6407
rect 6193 6373 6207 6387
rect 6213 6393 6227 6407
rect 6196 6363 6203 6373
rect 6236 6367 6243 6433
rect 6256 6407 6263 6453
rect 6296 6427 6303 6453
rect 6356 6443 6363 6453
rect 6356 6436 6383 6443
rect 6293 6413 6307 6427
rect 6253 6393 6267 6407
rect 6313 6373 6327 6387
rect 6176 6356 6203 6363
rect 6176 6343 6183 6356
rect 6156 6336 6183 6343
rect 6156 6327 6163 6336
rect 6136 6167 6143 6233
rect 6176 6167 6183 6273
rect 6196 6147 6203 6153
rect 6133 6123 6147 6127
rect 6116 6116 6147 6123
rect 6133 6113 6147 6116
rect 6193 6133 6207 6147
rect 6073 6093 6087 6107
rect 6036 6087 6043 6093
rect 6076 6087 6083 6093
rect 6096 6027 6103 6113
rect 6176 6087 6183 6113
rect 6216 6103 6223 6353
rect 6236 6167 6243 6173
rect 6276 6167 6283 6373
rect 6316 6347 6323 6373
rect 6356 6367 6363 6413
rect 6376 6387 6383 6436
rect 6353 6353 6367 6367
rect 6416 6347 6423 6413
rect 6516 6387 6523 6433
rect 6536 6427 6543 6433
rect 6533 6413 6547 6427
rect 6436 6247 6443 6373
rect 6453 6353 6467 6367
rect 6513 6373 6527 6387
rect 6553 6373 6567 6387
rect 6273 6113 6287 6127
rect 6196 6096 6223 6103
rect 6156 6047 6163 6073
rect 6156 5947 6163 6033
rect 6036 5927 6043 5933
rect 6076 5927 6083 5933
rect 6136 5927 6143 5933
rect 6176 5927 6183 5933
rect 6033 5913 6047 5927
rect 6013 5903 6027 5907
rect 5996 5896 6027 5903
rect 5936 5707 5943 5713
rect 5936 5647 5943 5693
rect 5956 5667 5963 5673
rect 5956 5647 5963 5653
rect 5853 5633 5867 5647
rect 5856 5607 5863 5633
rect 5953 5633 5967 5647
rect 5913 5613 5927 5627
rect 5916 5603 5923 5613
rect 5976 5623 5983 5733
rect 5996 5667 6003 5896
rect 6013 5893 6027 5896
rect 6073 5913 6087 5927
rect 6113 5893 6127 5907
rect 6133 5913 6147 5927
rect 6173 5913 6187 5927
rect 6116 5887 6123 5893
rect 6096 5847 6103 5873
rect 6116 5767 6123 5873
rect 6016 5647 6023 5693
rect 5993 5623 6007 5627
rect 5976 5616 6007 5623
rect 6013 5633 6027 5647
rect 5993 5613 6007 5616
rect 6033 5613 6047 5627
rect 6096 5643 6103 5673
rect 6176 5667 6183 5693
rect 6133 5653 6147 5667
rect 6113 5643 6127 5647
rect 6096 5636 6127 5643
rect 6113 5633 6127 5636
rect 5996 5607 6003 5613
rect 5933 5603 5947 5607
rect 5916 5596 5947 5603
rect 5933 5593 5947 5596
rect 5967 5596 5983 5603
rect 5876 5563 5883 5593
rect 5856 5556 5883 5563
rect 5796 5507 5803 5533
rect 5776 5487 5783 5493
rect 5713 5433 5727 5447
rect 5653 5396 5703 5403
rect 5653 5393 5667 5396
rect 5733 5393 5747 5407
rect 5736 5387 5743 5393
rect 5476 5203 5483 5313
rect 5536 5267 5543 5313
rect 5516 5227 5523 5253
rect 5556 5223 5563 5353
rect 5576 5247 5583 5353
rect 5556 5216 5583 5223
rect 5476 5196 5493 5203
rect 5576 5187 5583 5216
rect 5413 5153 5427 5167
rect 5453 5153 5467 5167
rect 5553 5153 5567 5167
rect 5573 5173 5587 5187
rect 5416 5147 5423 5153
rect 5336 4967 5343 4973
rect 5333 4953 5347 4967
rect 5416 4963 5423 5013
rect 5456 4987 5463 5153
rect 5476 4987 5483 5133
rect 5496 4967 5503 5133
rect 5536 4967 5543 5133
rect 5556 5107 5563 5153
rect 5576 5107 5583 5133
rect 5556 4987 5563 5013
rect 5453 4963 5467 4967
rect 5416 4956 5467 4963
rect 5356 4927 5363 4953
rect 5453 4953 5467 4956
rect 5473 4933 5487 4947
rect 5493 4953 5507 4967
rect 5513 4933 5527 4947
rect 5373 4913 5387 4927
rect 5276 4767 5283 4853
rect 5296 4727 5303 4793
rect 5016 4656 5043 4663
rect 4956 4467 4963 4513
rect 4996 4487 5003 4653
rect 5036 4607 5043 4656
rect 5116 4663 5123 4673
rect 5096 4656 5123 4663
rect 5036 4467 5043 4573
rect 5096 4567 5103 4656
rect 5153 4653 5167 4667
rect 5173 4673 5187 4687
rect 5193 4653 5207 4667
rect 5156 4647 5163 4653
rect 5196 4627 5203 4653
rect 5236 4647 5243 4673
rect 5256 4623 5263 4713
rect 5336 4687 5343 4713
rect 5356 4703 5363 4913
rect 5376 4827 5383 4913
rect 5416 4887 5423 4933
rect 5416 4807 5423 4873
rect 5436 4847 5443 4933
rect 5396 4776 5443 4783
rect 5396 4727 5403 4776
rect 5416 4707 5423 4733
rect 5373 4703 5387 4707
rect 5356 4696 5387 4703
rect 5373 4693 5387 4696
rect 5313 4653 5327 4667
rect 5333 4673 5347 4687
rect 5436 4667 5443 4776
rect 5353 4653 5367 4667
rect 5236 4616 5263 4623
rect 4933 4433 4947 4447
rect 4973 4433 4987 4447
rect 4936 4263 4943 4433
rect 4976 4407 4983 4433
rect 4996 4367 5003 4453
rect 5013 4433 5027 4447
rect 5033 4453 5047 4467
rect 5056 4447 5063 4553
rect 5136 4487 5143 4493
rect 5156 4487 5163 4533
rect 5113 4453 5127 4467
rect 5133 4473 5147 4487
rect 5053 4433 5067 4447
rect 4916 4256 4943 4263
rect 4795 4144 4803 4224
rect 4813 4183 4827 4187
rect 4836 4183 4843 4233
rect 4813 4176 4843 4183
rect 4856 4183 4863 4253
rect 4896 4207 4903 4213
rect 4873 4183 4887 4187
rect 4856 4176 4887 4183
rect 4893 4193 4907 4207
rect 4813 4173 4827 4176
rect 4873 4173 4887 4176
rect 4916 4067 4923 4256
rect 4956 4207 4963 4313
rect 4976 4227 4983 4273
rect 4996 4267 5003 4293
rect 5016 4267 5023 4433
rect 5056 4247 5063 4393
rect 5096 4387 5103 4433
rect 5116 4387 5123 4453
rect 5136 4367 5143 4433
rect 5176 4347 5183 4493
rect 5213 4453 5227 4467
rect 5196 4387 5203 4453
rect 5216 4367 5223 4453
rect 5096 4247 5103 4253
rect 5116 4227 5123 4253
rect 5136 4227 5143 4333
rect 5236 4247 5243 4616
rect 5276 4507 5283 4593
rect 5316 4507 5323 4653
rect 5336 4547 5343 4633
rect 5356 4627 5363 4653
rect 5376 4603 5383 4653
rect 5356 4596 5383 4603
rect 5336 4527 5343 4533
rect 5356 4507 5363 4596
rect 5396 4583 5403 4653
rect 5456 4627 5463 4853
rect 5476 4827 5483 4933
rect 5516 4927 5523 4933
rect 5496 4803 5503 4893
rect 5556 4847 5563 4973
rect 5576 4967 5583 5013
rect 5596 4987 5603 5353
rect 5616 5187 5623 5193
rect 5636 5167 5643 5173
rect 5633 5153 5647 5167
rect 5613 5123 5627 5127
rect 5613 5116 5633 5123
rect 5613 5113 5627 5116
rect 5616 4963 5623 5093
rect 5636 4967 5643 5113
rect 5656 4987 5663 5373
rect 5736 5347 5743 5373
rect 5736 5207 5743 5333
rect 5756 5327 5763 5453
rect 5773 5443 5787 5447
rect 5796 5443 5803 5493
rect 5856 5447 5863 5556
rect 5896 5447 5903 5493
rect 5916 5447 5923 5573
rect 5936 5467 5943 5593
rect 5773 5436 5803 5443
rect 5773 5433 5787 5436
rect 5853 5433 5867 5447
rect 5873 5413 5887 5427
rect 5936 5427 5943 5453
rect 5673 5153 5687 5167
rect 5713 5153 5727 5167
rect 5676 5147 5683 5153
rect 5696 5127 5703 5153
rect 5596 4956 5623 4963
rect 5596 4947 5603 4956
rect 5696 4963 5703 5093
rect 5716 5007 5723 5153
rect 5756 5087 5763 5213
rect 5776 5187 5783 5393
rect 5796 5167 5803 5293
rect 5816 5287 5823 5353
rect 5836 5227 5843 5413
rect 5856 5187 5863 5273
rect 5876 5247 5883 5413
rect 5933 5413 5947 5427
rect 5953 5403 5967 5407
rect 5976 5403 5983 5596
rect 5996 5527 6003 5573
rect 6016 5527 6023 5593
rect 5996 5483 6003 5513
rect 6036 5507 6043 5613
rect 6056 5567 6063 5593
rect 5996 5476 6043 5483
rect 5996 5427 6003 5453
rect 6036 5427 6043 5476
rect 6056 5447 6063 5533
rect 6076 5487 6083 5613
rect 6096 5467 6103 5513
rect 6116 5467 6123 5573
rect 6136 5567 6143 5653
rect 6153 5633 6167 5647
rect 6173 5653 6187 5667
rect 6156 5627 6163 5633
rect 6176 5527 6183 5613
rect 6136 5467 6143 5513
rect 6113 5453 6127 5467
rect 5953 5396 5983 5403
rect 5993 5413 6007 5427
rect 6033 5413 6047 5427
rect 5953 5393 5967 5396
rect 5896 5267 5903 5353
rect 5916 5347 5923 5393
rect 5936 5307 5943 5373
rect 5956 5307 5963 5393
rect 5936 5247 5943 5293
rect 5996 5247 6003 5373
rect 5773 5133 5787 5147
rect 5793 5153 5807 5167
rect 5876 5147 5883 5193
rect 5896 5187 5903 5233
rect 5936 5187 5943 5233
rect 5976 5223 5983 5233
rect 5976 5216 6003 5223
rect 5996 5207 6003 5216
rect 6016 5187 6023 5353
rect 6076 5307 6083 5433
rect 6156 5447 6163 5473
rect 6093 5413 6107 5427
rect 6133 5423 6147 5427
rect 6116 5416 6147 5423
rect 6153 5433 6167 5447
rect 6096 5387 6103 5413
rect 6116 5327 6123 5416
rect 6133 5413 6147 5416
rect 5893 5173 5907 5187
rect 5933 5173 5947 5187
rect 5953 5153 5967 5167
rect 6013 5173 6027 5187
rect 5956 5147 5963 5153
rect 5813 5133 5827 5147
rect 5776 5107 5783 5133
rect 5816 5107 5823 5133
rect 5836 5087 5843 5133
rect 5676 4956 5703 4963
rect 5676 4947 5683 4956
rect 5573 4913 5587 4927
rect 5593 4933 5607 4947
rect 5613 4913 5627 4927
rect 5673 4933 5687 4947
rect 5693 4913 5707 4927
rect 5576 4907 5583 4913
rect 5616 4907 5623 4913
rect 5636 4883 5643 4893
rect 5636 4876 5683 4883
rect 5476 4796 5503 4803
rect 5476 4747 5483 4796
rect 5576 4767 5583 4873
rect 5596 4787 5603 4853
rect 5476 4707 5483 4713
rect 5516 4707 5523 4713
rect 5473 4693 5487 4707
rect 5493 4673 5507 4687
rect 5533 4673 5547 4687
rect 5573 4673 5587 4687
rect 5376 4576 5403 4583
rect 5273 4503 5287 4507
rect 5273 4496 5303 4503
rect 5273 4493 5287 4496
rect 5296 4487 5303 4496
rect 5293 4473 5307 4487
rect 5333 4483 5347 4487
rect 5313 4453 5327 4467
rect 5333 4476 5353 4483
rect 5333 4473 5347 4476
rect 5276 4407 5283 4453
rect 5316 4443 5323 4453
rect 5307 4436 5323 4443
rect 5376 4447 5383 4576
rect 5396 4507 5403 4533
rect 5416 4527 5423 4573
rect 5393 4493 5407 4507
rect 5413 4463 5427 4467
rect 5396 4456 5427 4463
rect 5073 4223 5087 4227
rect 4953 4203 4967 4207
rect 4953 4196 4973 4203
rect 4953 4193 4967 4196
rect 5013 4193 5027 4207
rect 5073 4216 5103 4223
rect 5073 4213 5087 4216
rect 5016 4187 5023 4193
rect 5056 4183 5063 4193
rect 5056 4176 5083 4183
rect 5076 4147 5083 4176
rect 5096 4147 5103 4216
rect 5116 4167 5123 4213
rect 5196 4207 5203 4233
rect 5173 4173 5187 4187
rect 5233 4193 5247 4207
rect 5176 4127 5183 4173
rect 4936 4007 4943 4113
rect 4793 3953 4807 3967
rect 4833 3953 4847 3967
rect 4796 3947 4803 3953
rect 4836 3863 4843 3953
rect 4856 3887 4863 3993
rect 4913 3973 4927 3987
rect 4933 3993 4947 4007
rect 4916 3967 4923 3973
rect 4836 3856 4853 3863
rect 4916 3847 4923 3953
rect 4996 3924 5004 4036
rect 5073 4003 5087 4007
rect 5073 3996 5103 4003
rect 5073 3993 5087 3996
rect 4796 3664 4804 3776
rect 4935 3758 4943 3782
rect 4873 3703 4887 3707
rect 4896 3703 4903 3753
rect 4873 3696 4903 3703
rect 4873 3693 4887 3696
rect 4773 3513 4787 3527
rect 4713 3493 4727 3507
rect 4716 3487 4723 3493
rect 4635 3438 4643 3462
rect 4776 3387 4783 3513
rect 4797 3476 4805 3556
rect 4853 3523 4867 3527
rect 4876 3523 4883 3693
rect 4935 3664 4943 3744
rect 4956 3707 4963 3773
rect 5096 3767 5103 3996
rect 5135 3956 5143 4036
rect 5153 3993 5167 4007
rect 5156 3987 5163 3993
rect 5135 3918 5143 3942
rect 5156 3747 5163 3773
rect 5196 3767 5203 3993
rect 5236 3987 5243 4193
rect 5256 4127 5263 4313
rect 5296 4207 5303 4433
rect 5316 4144 5324 4256
rect 5336 4167 5343 4393
rect 5356 4247 5363 4413
rect 5376 4387 5383 4413
rect 5396 4227 5403 4456
rect 5413 4453 5427 4456
rect 5416 4307 5423 4433
rect 5393 4183 5407 4187
rect 5376 4176 5407 4183
rect 5256 4107 5263 4113
rect 5276 4067 5283 4133
rect 5276 3987 5283 4053
rect 5296 4027 5303 4113
rect 5356 4007 5363 4093
rect 5296 3987 5303 3993
rect 5213 3953 5227 3967
rect 5233 3973 5247 3987
rect 5293 3973 5307 3987
rect 5333 3973 5347 3987
rect 5353 3993 5367 4007
rect 5253 3953 5267 3967
rect 5336 3967 5343 3973
rect 5216 3807 5223 3953
rect 5256 3867 5263 3953
rect 5236 3747 5243 3853
rect 5256 3767 5263 3793
rect 5376 3767 5383 4176
rect 5393 4173 5407 4176
rect 5416 4167 5423 4293
rect 5436 4207 5443 4613
rect 5456 4447 5463 4493
rect 5476 4487 5483 4653
rect 5496 4607 5503 4673
rect 5536 4647 5543 4673
rect 5536 4563 5543 4633
rect 5556 4587 5563 4673
rect 5576 4567 5583 4673
rect 5516 4556 5543 4563
rect 5496 4467 5503 4533
rect 5516 4467 5523 4556
rect 5536 4467 5543 4493
rect 5576 4467 5583 4513
rect 5596 4487 5603 4653
rect 5473 4433 5487 4447
rect 5493 4453 5507 4467
rect 5573 4453 5587 4467
rect 5593 4433 5607 4447
rect 5616 4443 5623 4873
rect 5636 4647 5643 4713
rect 5656 4707 5663 4753
rect 5676 4727 5683 4876
rect 5696 4787 5703 4913
rect 5716 4887 5723 4973
rect 5716 4747 5723 4793
rect 5736 4767 5743 5073
rect 5773 4933 5787 4947
rect 5776 4927 5783 4933
rect 5756 4887 5763 4913
rect 5776 4847 5783 4893
rect 5756 4767 5763 4833
rect 5776 4783 5783 4833
rect 5796 4807 5803 4933
rect 5816 4907 5823 4933
rect 5836 4923 5843 5033
rect 5856 5027 5863 5133
rect 5876 4987 5883 5013
rect 5853 4923 5867 4927
rect 5836 4916 5867 4923
rect 5896 4927 5903 5073
rect 5916 5007 5923 5113
rect 5916 4967 5923 4973
rect 5853 4913 5867 4916
rect 5893 4913 5907 4927
rect 5776 4776 5803 4783
rect 5776 4707 5783 4713
rect 5653 4693 5667 4707
rect 5673 4673 5687 4687
rect 5713 4673 5727 4687
rect 5753 4673 5767 4687
rect 5773 4693 5787 4707
rect 5656 4527 5663 4613
rect 5676 4587 5683 4673
rect 5716 4667 5723 4673
rect 5636 4487 5643 4493
rect 5676 4487 5683 4533
rect 5696 4487 5703 4613
rect 5633 4473 5647 4487
rect 5653 4453 5667 4467
rect 5673 4473 5687 4487
rect 5616 4436 5643 4443
rect 5456 4387 5463 4393
rect 5476 4307 5483 4433
rect 5496 4347 5503 4413
rect 5516 4323 5523 4353
rect 5496 4316 5523 4323
rect 5476 4267 5483 4293
rect 5455 4238 5463 4262
rect 5455 4144 5463 4224
rect 5416 3987 5423 4053
rect 5456 4007 5463 4093
rect 5496 4027 5503 4316
rect 5536 4243 5543 4413
rect 5596 4387 5603 4433
rect 5516 4236 5543 4243
rect 5516 4227 5523 4236
rect 5556 4227 5563 4333
rect 5576 4227 5583 4253
rect 5513 4213 5527 4227
rect 5533 4193 5547 4207
rect 5553 4213 5567 4227
rect 5616 4207 5623 4413
rect 5636 4367 5643 4436
rect 5656 4327 5663 4453
rect 5696 4247 5703 4393
rect 5716 4347 5723 4633
rect 5736 4627 5743 4673
rect 5756 4587 5763 4673
rect 5776 4527 5783 4653
rect 5796 4587 5803 4776
rect 5736 4267 5743 4493
rect 5793 4433 5807 4447
rect 5796 4427 5803 4433
rect 5756 4387 5763 4413
rect 5756 4243 5763 4373
rect 5796 4287 5803 4333
rect 5736 4236 5763 4243
rect 5676 4207 5683 4233
rect 5536 4067 5543 4193
rect 5453 3993 5467 4007
rect 5393 3953 5407 3967
rect 5413 3973 5427 3987
rect 5516 3987 5523 4053
rect 5556 4047 5563 4173
rect 5576 4023 5583 4193
rect 5653 4173 5667 4187
rect 5673 4193 5687 4207
rect 5713 4193 5727 4207
rect 5716 4187 5723 4193
rect 5736 4187 5743 4236
rect 5796 4227 5803 4233
rect 5693 4173 5707 4187
rect 5593 4153 5607 4167
rect 5656 4163 5663 4173
rect 5647 4156 5663 4163
rect 5596 4127 5603 4153
rect 5596 4043 5603 4113
rect 5596 4036 5623 4043
rect 5556 4016 5583 4023
rect 5513 3973 5527 3987
rect 5433 3953 5447 3967
rect 5396 3787 5403 3953
rect 5436 3867 5443 3953
rect 5536 3927 5543 4013
rect 5556 3987 5563 4016
rect 5573 3973 5587 3987
rect 5576 3967 5583 3973
rect 5113 3743 5127 3747
rect 4953 3693 4967 3707
rect 4993 3693 5007 3707
rect 5013 3713 5027 3727
rect 5096 3736 5127 3743
rect 4996 3607 5003 3693
rect 5096 3607 5103 3736
rect 5113 3733 5127 3736
rect 5153 3733 5167 3747
rect 5193 3743 5207 3747
rect 5176 3736 5207 3743
rect 4853 3516 4883 3523
rect 4853 3513 4867 3516
rect 4797 3438 4805 3462
rect 4916 3403 4923 3533
rect 4936 3444 4944 3556
rect 4916 3396 4943 3403
rect 4716 3327 4723 3353
rect 4556 3247 4563 3273
rect 4453 3213 4467 3227
rect 4476 3223 4483 3233
rect 4493 3223 4507 3227
rect 4476 3216 4507 3223
rect 4513 3233 4527 3247
rect 4493 3213 4507 3216
rect 4553 3233 4567 3247
rect 4456 3183 4463 3213
rect 4496 3207 4503 3213
rect 4456 3176 4483 3183
rect 4256 3027 4263 3093
rect 4276 3067 4283 3113
rect 4296 3067 4303 3093
rect 4253 3013 4267 3027
rect 4276 2903 4283 2973
rect 4316 2964 4324 3076
rect 4393 3033 4407 3047
rect 4416 3007 4423 3093
rect 4276 2896 4303 2903
rect 4176 2807 4183 2853
rect 4296 2827 4303 2896
rect 4136 2647 4143 2773
rect 4176 2767 4183 2793
rect 4256 2767 4263 2773
rect 4173 2753 4187 2767
rect 4233 2733 4247 2747
rect 4253 2753 4267 2767
rect 4293 2763 4307 2767
rect 4316 2763 4323 2773
rect 4336 2767 4343 2993
rect 4436 2827 4443 3133
rect 4476 3087 4483 3176
rect 4496 3107 4503 3133
rect 4596 3107 4603 3273
rect 4613 3213 4627 3227
rect 4616 3207 4623 3213
rect 4653 3213 4667 3227
rect 4656 3207 4663 3213
rect 4455 2996 4463 3076
rect 4473 3043 4487 3047
rect 4496 3043 4503 3053
rect 4473 3036 4503 3043
rect 4473 3033 4487 3036
rect 4455 2958 4463 2982
rect 4516 2927 4523 3093
rect 4616 3087 4623 3193
rect 4576 3047 4583 3073
rect 4533 3033 4547 3047
rect 4553 3013 4567 3027
rect 4573 3033 4587 3047
rect 4593 3013 4607 3027
rect 4556 3003 4563 3013
rect 4536 2996 4563 3003
rect 4536 2967 4543 2996
rect 4416 2803 4423 2813
rect 4416 2796 4443 2803
rect 4293 2756 4323 2763
rect 4293 2753 4307 2756
rect 4393 2773 4407 2787
rect 4396 2767 4403 2773
rect 4373 2753 4387 2767
rect 4273 2733 4287 2747
rect 4193 2713 4207 2727
rect 3996 2596 4043 2603
rect 3996 2587 4003 2596
rect 4036 2587 4043 2596
rect 3796 2527 3803 2533
rect 3813 2513 3827 2527
rect 3833 2533 3847 2547
rect 3913 2533 3927 2547
rect 3933 2553 3947 2567
rect 4056 2567 4063 2633
rect 3953 2533 3967 2547
rect 3993 2533 4007 2547
rect 4053 2553 4067 2567
rect 3996 2527 4003 2533
rect 3796 2507 3803 2513
rect 3816 2487 3823 2513
rect 3636 2416 3663 2423
rect 3596 2224 3604 2336
rect 3636 2327 3643 2416
rect 3633 2253 3647 2267
rect 3636 2227 3643 2253
rect 3636 2163 3643 2193
rect 3596 2156 3643 2163
rect 3356 1883 3363 1893
rect 3356 1876 3383 1883
rect 3376 1847 3383 1876
rect 3396 1847 3403 1893
rect 3516 1867 3523 1913
rect 3576 1887 3583 1893
rect 3356 1823 3363 1833
rect 3576 1827 3583 1873
rect 3356 1816 3383 1823
rect 3353 1773 3367 1787
rect 3376 1783 3383 1816
rect 3393 1813 3407 1827
rect 3413 1793 3427 1807
rect 3533 1823 3547 1827
rect 3527 1816 3547 1823
rect 3533 1813 3547 1816
rect 3376 1776 3423 1783
rect 3316 1683 3323 1713
rect 3296 1676 3323 1683
rect 3176 1656 3203 1663
rect 3196 1607 3203 1656
rect 3153 1593 3167 1607
rect 3193 1593 3207 1607
rect 3116 1436 3143 1443
rect 2913 1293 2927 1307
rect 2887 1176 2903 1183
rect 2916 1167 2923 1293
rect 2936 1227 2943 1333
rect 2956 1327 2963 1373
rect 2976 1347 2983 1413
rect 3116 1367 3123 1436
rect 2996 1327 3003 1333
rect 2973 1303 2987 1307
rect 2956 1296 2987 1303
rect 2993 1313 3007 1327
rect 2956 1287 2963 1296
rect 2973 1293 2987 1296
rect 3053 1293 3067 1307
rect 2887 1156 2903 1163
rect 2896 1143 2903 1156
rect 2896 1136 2923 1143
rect 2876 1127 2883 1133
rect 2916 1127 2923 1136
rect 2873 1113 2887 1127
rect 2893 1093 2907 1107
rect 2913 1113 2927 1127
rect 2953 1123 2967 1127
rect 2976 1123 2983 1233
rect 2933 1093 2947 1107
rect 2953 1116 2983 1123
rect 2953 1113 2967 1116
rect 2896 1083 2903 1093
rect 2896 1076 2923 1083
rect 2816 996 2863 1003
rect 2736 647 2743 693
rect 2776 647 2783 693
rect 2693 633 2707 647
rect 2733 633 2747 647
rect 2695 398 2703 422
rect 2695 304 2703 384
rect 2716 347 2723 353
rect 2736 347 2743 493
rect 2796 387 2803 833
rect 2816 807 2823 996
rect 2836 803 2843 973
rect 2856 847 2863 933
rect 2853 833 2867 847
rect 2876 843 2883 853
rect 2916 847 2923 1076
rect 2936 1067 2943 1093
rect 2976 847 2983 1116
rect 2996 1047 3003 1113
rect 3016 1044 3024 1156
rect 3036 1047 3043 1273
rect 3056 1247 3063 1293
rect 3076 1007 3083 1333
rect 3113 1273 3127 1287
rect 3096 1127 3103 1133
rect 3093 1113 3107 1127
rect 3116 1087 3123 1273
rect 3136 1187 3143 1393
rect 3216 1347 3223 1613
rect 3255 1556 3263 1636
rect 3273 1593 3287 1607
rect 3296 1567 3303 1676
rect 3376 1647 3383 1753
rect 3236 1367 3243 1553
rect 3316 1543 3323 1633
rect 3373 1553 3387 1567
rect 3376 1543 3383 1553
rect 3255 1518 3263 1542
rect 3316 1536 3383 1543
rect 3396 1527 3403 1613
rect 3416 1607 3423 1776
rect 3453 1773 3467 1787
rect 3516 1767 3523 1813
rect 3553 1793 3567 1807
rect 3573 1813 3587 1827
rect 3556 1667 3563 1793
rect 3596 1763 3603 2156
rect 3656 2147 3663 2273
rect 3673 2253 3687 2267
rect 3616 2007 3623 2093
rect 3635 2036 3643 2116
rect 3676 2087 3683 2253
rect 3696 2167 3703 2473
rect 3716 2207 3723 2473
rect 3735 2318 3743 2342
rect 3776 2307 3783 2413
rect 3896 2407 3903 2513
rect 3836 2307 3843 2393
rect 3735 2224 3743 2304
rect 3776 2207 3783 2293
rect 3813 2273 3827 2287
rect 3856 2283 3863 2393
rect 3936 2307 3943 2333
rect 3873 2283 3887 2287
rect 3856 2276 3887 2283
rect 3716 2107 3723 2133
rect 3733 2103 3747 2107
rect 3733 2096 3753 2103
rect 3733 2093 3747 2096
rect 3653 2073 3667 2087
rect 3713 2073 3727 2087
rect 3656 2047 3663 2073
rect 3753 2073 3767 2087
rect 3776 2067 3783 2173
rect 3816 2107 3823 2253
rect 3856 2167 3863 2276
rect 3873 2273 3887 2276
rect 3896 2267 3903 2293
rect 3913 2273 3927 2287
rect 3933 2293 3947 2307
rect 3796 2087 3803 2093
rect 3836 2087 3843 2113
rect 3876 2107 3883 2253
rect 3916 2227 3923 2273
rect 3793 2073 3807 2087
rect 3833 2073 3847 2087
rect 3853 2053 3867 2067
rect 3635 1998 3643 2022
rect 3676 1847 3683 2013
rect 3613 1773 3627 1787
rect 3633 1793 3647 1807
rect 3673 1793 3687 1807
rect 3653 1783 3667 1787
rect 3653 1776 3673 1783
rect 3653 1773 3667 1776
rect 3696 1767 3703 1993
rect 3716 1827 3723 1973
rect 3736 1967 3743 2053
rect 3756 1987 3763 2033
rect 3733 1813 3747 1827
rect 3753 1793 3767 1807
rect 3596 1756 3623 1763
rect 3516 1636 3583 1643
rect 3476 1607 3483 1633
rect 3516 1623 3523 1636
rect 3576 1627 3583 1636
rect 3496 1616 3523 1623
rect 3496 1607 3503 1616
rect 3536 1607 3543 1613
rect 3453 1573 3467 1587
rect 3473 1593 3487 1607
rect 3493 1593 3507 1607
rect 3533 1593 3547 1607
rect 3573 1603 3587 1607
rect 3596 1603 3603 1653
rect 3553 1573 3567 1587
rect 3573 1596 3603 1603
rect 3573 1593 3587 1596
rect 3256 1407 3263 1413
rect 3256 1343 3263 1393
rect 3236 1336 3263 1343
rect 3236 1327 3243 1336
rect 3153 1293 3167 1307
rect 3173 1313 3187 1327
rect 3213 1293 3227 1307
rect 3233 1313 3247 1327
rect 3156 1203 3163 1293
rect 3196 1203 3203 1213
rect 3156 1196 3203 1203
rect 3216 1167 3223 1293
rect 2893 843 2907 847
rect 2876 836 2907 843
rect 2893 833 2907 836
rect 2836 796 2863 803
rect 2816 707 2823 773
rect 2836 667 2843 673
rect 2833 653 2847 667
rect 2856 607 2863 796
rect 2913 793 2927 807
rect 2916 727 2923 793
rect 2976 787 2983 833
rect 2996 823 3003 993
rect 3096 887 3103 953
rect 3116 927 3123 1073
rect 3136 1003 3143 1153
rect 3155 1076 3163 1156
rect 3236 1147 3243 1273
rect 3276 1207 3283 1413
rect 3296 1264 3304 1376
rect 3316 1227 3323 1453
rect 3173 1123 3187 1127
rect 3256 1123 3263 1173
rect 3356 1147 3363 1493
rect 3376 1427 3383 1513
rect 3456 1487 3463 1573
rect 3396 1347 3403 1413
rect 3435 1358 3443 1382
rect 3396 1307 3403 1333
rect 3373 1293 3387 1307
rect 3376 1283 3383 1293
rect 3376 1276 3403 1283
rect 3376 1127 3383 1253
rect 3396 1207 3403 1276
rect 3435 1264 3443 1344
rect 3456 1307 3463 1333
rect 3453 1293 3467 1307
rect 3476 1187 3483 1453
rect 3496 1227 3503 1433
rect 3576 1327 3583 1553
rect 3596 1447 3603 1553
rect 3616 1507 3623 1756
rect 3796 1727 3803 1853
rect 3816 1827 3823 1893
rect 3816 1807 3823 1813
rect 3836 1807 3843 1953
rect 3856 1847 3863 2053
rect 3896 2047 3903 2193
rect 3936 2107 3943 2253
rect 3956 2247 3963 2493
rect 4016 2487 4023 2533
rect 3976 2287 3983 2433
rect 3973 2273 3987 2287
rect 3976 2207 3983 2233
rect 3996 2203 4003 2253
rect 4016 2227 4023 2373
rect 4036 2307 4043 2513
rect 4076 2467 4083 2593
rect 4113 2553 4127 2567
rect 4153 2553 4167 2567
rect 4056 2407 4063 2453
rect 4053 2253 4067 2267
rect 4056 2243 4063 2253
rect 4036 2236 4063 2243
rect 4036 2207 4043 2236
rect 3996 2196 4023 2203
rect 4016 2187 4023 2196
rect 3956 2087 3963 2093
rect 3996 2087 4003 2173
rect 4016 2107 4023 2113
rect 4036 2107 4043 2153
rect 3953 2073 3967 2087
rect 3973 2053 3987 2067
rect 3993 2073 4007 2087
rect 4016 2083 4023 2093
rect 4056 2083 4063 2193
rect 4076 2167 4083 2413
rect 4096 2287 4103 2513
rect 4116 2307 4123 2493
rect 4093 2273 4107 2287
rect 4136 2243 4143 2433
rect 4156 2287 4163 2413
rect 4176 2387 4183 2713
rect 4196 2647 4203 2713
rect 4196 2607 4203 2633
rect 4216 2607 4223 2713
rect 4196 2567 4203 2573
rect 4236 2567 4243 2613
rect 4256 2587 4263 2713
rect 4276 2687 4283 2733
rect 4296 2723 4303 2733
rect 4336 2727 4343 2733
rect 4296 2716 4323 2723
rect 4193 2553 4207 2567
rect 4213 2533 4227 2547
rect 4233 2553 4247 2567
rect 4253 2533 4267 2547
rect 4296 2547 4303 2593
rect 4216 2467 4223 2533
rect 4236 2403 4243 2493
rect 4256 2467 4263 2473
rect 4216 2396 4243 2403
rect 4153 2273 4167 2287
rect 4173 2253 4187 2267
rect 4176 2247 4183 2253
rect 4116 2236 4143 2243
rect 4096 2087 4103 2213
rect 4016 2076 4043 2083
rect 4056 2076 4083 2083
rect 4036 2067 4043 2076
rect 4076 2067 4083 2076
rect 3907 2016 3923 2023
rect 3896 1907 3903 1993
rect 3916 1967 3923 2016
rect 3936 1987 3943 2053
rect 3976 2043 3983 2053
rect 3967 2036 3983 2043
rect 4073 2053 4087 2067
rect 4093 2033 4107 2047
rect 3996 1947 4003 2033
rect 4096 2027 4103 2033
rect 4116 2023 4123 2236
rect 4136 2107 4143 2213
rect 4196 2127 4203 2353
rect 4216 2287 4223 2396
rect 4236 2307 4243 2373
rect 4213 2273 4227 2287
rect 4233 2253 4247 2267
rect 4236 2187 4243 2253
rect 4256 2247 4263 2453
rect 4296 2303 4303 2413
rect 4316 2387 4323 2716
rect 4356 2667 4363 2733
rect 4376 2727 4383 2753
rect 4396 2747 4403 2753
rect 4436 2727 4443 2796
rect 4476 2704 4484 2816
rect 4496 2707 4503 2893
rect 4556 2847 4563 2973
rect 4596 2887 4603 3013
rect 4636 3007 4643 3093
rect 4676 3087 4683 3273
rect 4716 3247 4723 3313
rect 4733 3213 4747 3227
rect 4696 3007 4703 3193
rect 4736 3087 4743 3213
rect 4756 3203 4763 3373
rect 4816 3223 4823 3273
rect 4896 3247 4903 3353
rect 4833 3223 4847 3227
rect 4816 3216 4847 3223
rect 4833 3213 4847 3216
rect 4873 3213 4887 3227
rect 4893 3233 4907 3247
rect 4773 3203 4787 3207
rect 4756 3196 4787 3203
rect 4773 3193 4787 3196
rect 4876 3203 4883 3213
rect 4876 3196 4913 3203
rect 4716 3047 4723 3053
rect 4713 3033 4727 3047
rect 4733 3013 4747 3027
rect 4516 2787 4523 2813
rect 4615 2798 4623 2822
rect 4513 2733 4527 2747
rect 4553 2733 4567 2747
rect 4336 2484 4344 2596
rect 4356 2367 4363 2633
rect 4376 2567 4383 2613
rect 4373 2553 4387 2567
rect 4396 2487 4403 2693
rect 4416 2607 4423 2653
rect 4413 2553 4427 2567
rect 4416 2387 4423 2513
rect 4436 2427 4443 2693
rect 4516 2687 4523 2733
rect 4576 2723 4583 2773
rect 4556 2716 4583 2723
rect 4536 2663 4543 2693
rect 4516 2656 4543 2663
rect 4516 2627 4523 2656
rect 4556 2643 4563 2716
rect 4615 2704 4623 2784
rect 4536 2636 4563 2643
rect 4475 2516 4483 2596
rect 4475 2478 4483 2502
rect 4296 2296 4323 2303
rect 4276 2287 4283 2293
rect 4273 2273 4287 2287
rect 4256 2163 4263 2193
rect 4236 2156 4263 2163
rect 4173 2093 4187 2107
rect 4153 2073 4167 2087
rect 4236 2087 4243 2156
rect 4176 2027 4183 2053
rect 4116 2016 4143 2023
rect 4036 1847 4043 1933
rect 4056 1927 4063 2013
rect 4056 1907 4063 1913
rect 3813 1793 3827 1807
rect 3833 1753 3847 1767
rect 3656 1607 3663 1713
rect 3676 1667 3683 1693
rect 3653 1593 3667 1607
rect 3633 1573 3647 1587
rect 3673 1573 3687 1587
rect 3716 1583 3723 1653
rect 3753 1613 3767 1627
rect 3733 1583 3747 1587
rect 3716 1576 3747 1583
rect 3733 1573 3747 1576
rect 3716 1487 3723 1533
rect 3696 1447 3703 1473
rect 3656 1327 3663 1333
rect 3553 1293 3567 1307
rect 3593 1303 3607 1307
rect 3576 1296 3607 1303
rect 3576 1287 3583 1296
rect 3593 1293 3607 1296
rect 3633 1293 3647 1307
rect 3653 1313 3667 1327
rect 3673 1303 3687 1307
rect 3696 1303 3703 1433
rect 3756 1427 3763 1553
rect 3716 1367 3723 1413
rect 3776 1407 3783 1713
rect 3816 1627 3823 1633
rect 3836 1627 3843 1753
rect 3856 1723 3863 1753
rect 3876 1747 3883 1793
rect 3933 1773 3947 1787
rect 3973 1773 3987 1787
rect 3976 1727 3983 1773
rect 3856 1716 3883 1723
rect 3876 1707 3883 1716
rect 3813 1613 3827 1627
rect 3793 1593 3807 1607
rect 3816 1507 3823 1573
rect 3856 1567 3863 1693
rect 3876 1607 3883 1633
rect 3916 1607 3923 1633
rect 3996 1627 4003 1813
rect 4036 1807 4043 1833
rect 4076 1807 4083 1993
rect 4096 1867 4103 2013
rect 4013 1773 4027 1787
rect 4033 1793 4047 1807
rect 4053 1773 4067 1787
rect 4073 1793 4087 1807
rect 4093 1773 4107 1787
rect 4016 1667 4023 1773
rect 4056 1687 4063 1773
rect 4096 1747 4103 1773
rect 3873 1593 3887 1607
rect 3893 1573 3907 1587
rect 3913 1593 3927 1607
rect 3953 1603 3967 1607
rect 3933 1573 3947 1587
rect 3953 1596 3983 1603
rect 3953 1593 3967 1596
rect 3976 1583 3983 1596
rect 3993 1583 4007 1587
rect 3976 1576 4007 1583
rect 3993 1573 4007 1576
rect 3716 1307 3723 1313
rect 3673 1296 3703 1303
rect 3673 1293 3687 1296
rect 3753 1313 3767 1327
rect 3773 1293 3787 1307
rect 3313 1123 3327 1127
rect 3173 1116 3263 1123
rect 3296 1116 3327 1123
rect 3173 1113 3187 1116
rect 3196 1083 3203 1093
rect 3213 1083 3227 1087
rect 3196 1076 3227 1083
rect 3213 1073 3227 1076
rect 3155 1038 3163 1062
rect 3136 996 3163 1003
rect 3136 847 3143 953
rect 3156 847 3163 996
rect 3176 967 3183 1073
rect 3216 1007 3223 1073
rect 3196 847 3203 953
rect 3013 823 3027 827
rect 2996 816 3027 823
rect 3073 843 3087 847
rect 3073 836 3103 843
rect 3073 833 3087 836
rect 3013 813 3027 816
rect 3053 793 3067 807
rect 2916 667 2923 713
rect 2936 667 2943 693
rect 2996 687 3003 793
rect 3056 727 3063 793
rect 2913 653 2927 667
rect 2876 647 2883 653
rect 2873 633 2887 647
rect 3016 647 3023 653
rect 3056 647 3063 693
rect 3096 687 3103 836
rect 3113 813 3127 827
rect 3133 833 3147 847
rect 3173 813 3187 827
rect 3193 833 3207 847
rect 3116 707 3123 813
rect 3176 807 3183 813
rect 2973 613 2987 627
rect 3013 633 3027 647
rect 3033 613 3047 627
rect 3053 633 3067 647
rect 3076 627 3083 633
rect 3073 613 3087 627
rect 2976 547 2983 613
rect 3036 603 3043 613
rect 3036 596 3063 603
rect 3096 603 3103 653
rect 3116 643 3123 653
rect 3156 647 3163 753
rect 3216 743 3223 993
rect 3256 863 3263 1073
rect 3276 1027 3283 1093
rect 3296 1087 3303 1116
rect 3313 1113 3327 1116
rect 3333 1093 3347 1107
rect 3373 1113 3387 1127
rect 3393 1093 3407 1107
rect 3473 1093 3487 1107
rect 3336 1087 3343 1093
rect 3316 1047 3323 1073
rect 3256 856 3283 863
rect 3233 813 3247 827
rect 3236 787 3243 813
rect 3196 736 3223 743
rect 3116 636 3143 643
rect 3136 627 3143 636
rect 3113 603 3127 607
rect 3096 596 3127 603
rect 3133 613 3147 627
rect 3153 603 3167 607
rect 3176 603 3183 693
rect 3196 667 3203 736
rect 3196 627 3203 633
rect 3236 627 3243 733
rect 3016 583 3023 593
rect 3007 576 3023 583
rect 2713 333 2727 347
rect 2756 323 2763 373
rect 2816 367 2823 373
rect 2773 353 2787 367
rect 2776 347 2783 353
rect 2793 333 2807 347
rect 2813 353 2827 367
rect 2833 333 2847 347
rect 2853 333 2867 347
rect 2756 316 2783 323
rect 2596 167 2603 213
rect 2656 187 2663 193
rect 2653 173 2667 187
rect 2493 116 2523 123
rect 2593 153 2607 167
rect 2616 127 2623 153
rect 2493 113 2507 116
rect 1396 -24 1423 -17
rect 1556 -24 1583 -17
rect 1796 -24 1823 -17
rect 1876 -24 1903 -17
rect 1956 -24 1983 -17
rect 2376 -24 2403 -17
rect 2456 -24 2463 113
rect 2716 84 2724 196
rect 2753 163 2767 167
rect 2736 156 2767 163
rect 2736 127 2743 156
rect 2753 153 2767 156
rect 2776 47 2783 316
rect 2796 267 2803 333
rect 2836 247 2843 333
rect 2856 327 2863 333
rect 2893 333 2907 347
rect 2936 327 2943 373
rect 2856 287 2863 313
rect 2976 304 2984 416
rect 2996 387 3003 573
rect 3016 567 3023 576
rect 3056 547 3063 596
rect 3113 593 3127 596
rect 3153 596 3183 603
rect 3193 613 3207 627
rect 3233 613 3247 627
rect 3153 593 3167 596
rect 3213 593 3227 607
rect 3253 593 3267 607
rect 3013 333 3027 347
rect 3016 267 3023 333
rect 2796 167 2803 173
rect 2793 153 2807 167
rect 2855 116 2863 196
rect 2873 163 2887 167
rect 2896 163 2903 193
rect 2996 167 3003 193
rect 3036 167 3043 473
rect 3053 333 3067 347
rect 3056 307 3063 333
rect 2873 156 2903 163
rect 2873 153 2887 156
rect 2896 127 2903 156
rect 2933 143 2947 147
rect 2916 136 2947 143
rect 2916 107 2923 136
rect 2933 133 2947 136
rect 2973 133 2987 147
rect 2993 153 3007 167
rect 3033 153 3047 167
rect 3076 167 3083 273
rect 3096 247 3103 413
rect 3115 398 3123 422
rect 3115 304 3123 384
rect 3156 383 3163 593
rect 3176 567 3183 573
rect 3256 507 3263 593
rect 3276 403 3283 856
rect 3316 847 3323 953
rect 3376 947 3383 1053
rect 3396 967 3403 1093
rect 3396 847 3403 933
rect 3436 867 3443 1013
rect 3456 927 3463 1013
rect 3476 867 3483 913
rect 3433 853 3447 867
rect 3293 813 3307 827
rect 3313 833 3327 847
rect 3353 833 3367 847
rect 3296 707 3303 813
rect 3336 727 3343 833
rect 3356 727 3363 833
rect 3393 833 3407 847
rect 3453 833 3467 847
rect 3473 853 3487 867
rect 3496 843 3503 1033
rect 3516 887 3523 1213
rect 3536 887 3543 1153
rect 3556 967 3563 1073
rect 3576 987 3583 1233
rect 3596 1167 3603 1273
rect 3596 1127 3603 1133
rect 3593 1113 3607 1127
rect 3616 1027 3623 1273
rect 3636 1127 3643 1293
rect 3776 1283 3783 1293
rect 3756 1276 3783 1283
rect 3676 1183 3683 1273
rect 3696 1207 3703 1273
rect 3676 1176 3703 1183
rect 3696 1167 3703 1176
rect 3656 1044 3664 1156
rect 3676 1107 3683 1153
rect 3576 847 3583 873
rect 3513 843 3527 847
rect 3496 836 3527 843
rect 3513 833 3527 836
rect 3413 813 3427 827
rect 3296 667 3303 693
rect 3293 653 3307 667
rect 3336 607 3343 653
rect 3356 647 3363 653
rect 3396 647 3403 673
rect 3416 667 3423 813
rect 3456 727 3463 833
rect 3573 833 3587 847
rect 3533 813 3547 827
rect 3496 647 3503 773
rect 3536 767 3543 813
rect 3556 787 3563 833
rect 3553 653 3567 667
rect 3353 633 3367 647
rect 3393 633 3407 647
rect 3396 467 3403 573
rect 3256 396 3283 403
rect 3173 383 3187 387
rect 3156 376 3187 383
rect 3213 383 3227 387
rect 3133 343 3147 347
rect 3156 343 3163 376
rect 3173 373 3187 376
rect 3213 376 3243 383
rect 3213 373 3227 376
rect 3133 336 3163 343
rect 3133 333 3147 336
rect 3236 247 3243 376
rect 3116 167 3123 193
rect 3156 167 3163 193
rect 3256 187 3263 396
rect 3316 367 3323 393
rect 3293 333 3307 347
rect 3313 353 3327 367
rect 3333 333 3347 347
rect 3353 333 3367 347
rect 3393 343 3407 347
rect 3416 343 3423 473
rect 3436 467 3443 633
rect 3533 613 3547 627
rect 3573 613 3587 627
rect 3476 367 3483 493
rect 3496 367 3503 593
rect 3536 387 3543 613
rect 3576 507 3583 613
rect 3616 547 3623 913
rect 3636 647 3643 1013
rect 3716 1007 3723 1213
rect 3736 1127 3743 1253
rect 3756 1227 3763 1276
rect 3796 1267 3803 1493
rect 3896 1443 3903 1573
rect 4076 1524 4084 1636
rect 3876 1436 3903 1443
rect 3856 1403 3863 1433
rect 3816 1396 3863 1403
rect 3816 1327 3823 1396
rect 3876 1347 3883 1436
rect 3956 1387 3963 1433
rect 3897 1358 3905 1382
rect 3813 1313 3827 1327
rect 3873 1303 3887 1307
rect 3833 1283 3847 1287
rect 3816 1276 3847 1283
rect 3816 1167 3823 1276
rect 3833 1273 3847 1276
rect 3856 1296 3887 1303
rect 3733 1123 3747 1127
rect 3733 1116 3763 1123
rect 3733 1113 3747 1116
rect 3656 847 3663 933
rect 3653 833 3667 847
rect 3696 823 3703 913
rect 3713 823 3727 827
rect 3696 816 3727 823
rect 3713 813 3727 816
rect 3673 793 3687 807
rect 3656 667 3663 793
rect 3676 767 3683 793
rect 3716 667 3723 793
rect 3756 747 3763 1116
rect 3776 1067 3783 1153
rect 3795 1076 3803 1156
rect 3776 867 3783 1053
rect 3795 1038 3803 1062
rect 3796 847 3803 953
rect 3836 867 3843 1253
rect 3856 1187 3863 1296
rect 3873 1293 3887 1296
rect 3897 1264 3905 1344
rect 3876 1127 3883 1153
rect 3853 1093 3867 1107
rect 3856 967 3863 1093
rect 3896 1047 3903 1153
rect 3916 1147 3923 1333
rect 3953 1293 3967 1307
rect 3956 1287 3963 1293
rect 3936 1127 3943 1173
rect 3913 1093 3927 1107
rect 3916 1027 3923 1093
rect 3956 1047 3963 1113
rect 3773 813 3787 827
rect 3793 833 3807 847
rect 3776 767 3783 813
rect 3856 784 3864 896
rect 3876 823 3883 873
rect 3916 827 3923 933
rect 3893 823 3907 827
rect 3876 816 3907 823
rect 3893 813 3907 816
rect 3933 813 3947 827
rect 3653 653 3667 667
rect 3673 633 3687 647
rect 3753 643 3767 647
rect 3753 636 3773 643
rect 3753 633 3767 636
rect 3576 427 3583 493
rect 3636 407 3643 513
rect 3516 367 3523 373
rect 3556 367 3563 393
rect 3656 367 3663 613
rect 3796 607 3803 753
rect 3816 707 3823 753
rect 3856 627 3863 713
rect 3876 627 3883 773
rect 3936 747 3943 813
rect 3956 787 3963 913
rect 3976 907 3983 1373
rect 4016 1247 4023 1513
rect 4096 1487 4103 1693
rect 4116 1607 4123 1633
rect 4113 1593 4127 1607
rect 4136 1563 4143 2016
rect 4156 1947 4163 1993
rect 4176 1947 4183 1973
rect 4176 1807 4183 1893
rect 4216 1887 4223 1913
rect 4236 1907 4243 2073
rect 4256 2004 4264 2116
rect 4276 2047 4283 2133
rect 4296 2087 4303 2173
rect 4293 2073 4307 2087
rect 4236 1807 4243 1873
rect 4256 1863 4263 1953
rect 4256 1856 4273 1863
rect 4296 1827 4303 1973
rect 4316 1823 4323 2296
rect 4336 2107 4343 2233
rect 4376 2227 4383 2253
rect 4396 2227 4403 2373
rect 4496 2287 4503 2493
rect 4536 2367 4543 2636
rect 4556 2607 4563 2613
rect 4556 2583 4563 2593
rect 4573 2583 4587 2587
rect 4556 2576 4587 2583
rect 4573 2573 4587 2576
rect 4656 2567 4663 2993
rect 4716 2887 4723 2993
rect 4736 2987 4743 3013
rect 4756 2923 4763 3133
rect 4856 3107 4863 3193
rect 4796 3063 4803 3093
rect 4776 3056 4803 3063
rect 4776 3047 4783 3056
rect 4856 3047 4863 3053
rect 4773 3033 4787 3047
rect 4793 3013 4807 3027
rect 4853 3033 4867 3047
rect 4873 3013 4887 3027
rect 4796 3007 4803 3013
rect 4776 2943 4783 2993
rect 4776 2936 4803 2943
rect 4756 2916 4783 2923
rect 4776 2887 4783 2916
rect 4696 2767 4703 2853
rect 4796 2843 4803 2936
rect 4816 2923 4823 2973
rect 4836 2947 4843 3013
rect 4916 2927 4923 3053
rect 4936 2927 4943 3396
rect 4956 3267 4963 3513
rect 4976 3247 4983 3413
rect 4996 3287 5003 3593
rect 5016 3527 5023 3533
rect 5056 3527 5063 3573
rect 5096 3527 5103 3593
rect 5153 3543 5167 3547
rect 5176 3543 5183 3736
rect 5193 3733 5207 3736
rect 5213 3713 5227 3727
rect 5233 3733 5247 3747
rect 5336 3727 5343 3733
rect 5216 3687 5223 3713
rect 5333 3713 5347 3727
rect 5236 3567 5243 3673
rect 5356 3667 5363 3713
rect 5153 3536 5183 3543
rect 5153 3533 5167 3536
rect 5013 3513 5027 3527
rect 5033 3493 5047 3507
rect 5053 3513 5067 3527
rect 5093 3513 5107 3527
rect 5176 3523 5183 3536
rect 5193 3523 5207 3527
rect 5176 3516 5207 3523
rect 5193 3513 5207 3516
rect 4996 3267 5003 3273
rect 4996 3247 5003 3253
rect 4953 3243 4967 3247
rect 4953 3236 4973 3243
rect 4953 3233 4967 3236
rect 4993 3233 5007 3247
rect 5013 3223 5027 3227
rect 5036 3223 5043 3493
rect 5217 3476 5225 3556
rect 5276 3527 5283 3533
rect 5316 3527 5323 3573
rect 5273 3513 5287 3527
rect 5313 3513 5327 3527
rect 5217 3438 5225 3462
rect 5097 3278 5105 3302
rect 5073 3223 5087 3227
rect 5013 3216 5043 3223
rect 5056 3216 5087 3223
rect 5013 3213 5027 3216
rect 4973 3193 4987 3207
rect 5056 3167 5063 3216
rect 5073 3213 5087 3216
rect 5097 3184 5105 3264
rect 4976 3116 5023 3123
rect 4976 3107 4983 3116
rect 4996 3047 5003 3093
rect 5016 3067 5023 3116
rect 5036 3047 5043 3133
rect 5116 3067 5123 3093
rect 5113 3053 5127 3067
rect 4993 3033 5007 3047
rect 5013 3013 5027 3027
rect 5033 3033 5047 3047
rect 5073 3043 5087 3047
rect 5053 3013 5067 3027
rect 5073 3036 5103 3043
rect 5073 3033 5087 3036
rect 4816 2916 4843 2923
rect 4796 2836 4823 2843
rect 4816 2787 4823 2836
rect 4836 2827 4843 2916
rect 4956 2903 4963 2993
rect 4976 2967 4983 3013
rect 4936 2896 4963 2903
rect 4693 2753 4707 2767
rect 4733 2733 4747 2747
rect 4773 2733 4787 2747
rect 4813 2733 4827 2747
rect 4833 2753 4847 2767
rect 4873 2753 4887 2767
rect 4853 2733 4867 2747
rect 4776 2727 4783 2733
rect 4753 2713 4767 2727
rect 4676 2587 4683 2713
rect 4736 2647 4743 2713
rect 4816 2707 4823 2713
rect 4736 2567 4743 2593
rect 4553 2533 4567 2547
rect 4653 2553 4667 2567
rect 4673 2533 4687 2547
rect 4693 2553 4707 2567
rect 4713 2533 4727 2547
rect 4733 2553 4747 2567
rect 4556 2527 4563 2533
rect 4516 2303 4523 2333
rect 4516 2296 4543 2303
rect 4433 2253 4447 2267
rect 4473 2253 4487 2267
rect 4536 2267 4543 2296
rect 4556 2287 4563 2493
rect 4576 2427 4583 2533
rect 4676 2507 4683 2533
rect 4716 2523 4723 2533
rect 4716 2516 4743 2523
rect 4553 2273 4567 2287
rect 4513 2253 4527 2267
rect 4573 2253 4587 2267
rect 4453 2233 4467 2247
rect 4456 2167 4463 2233
rect 4376 2087 4383 2133
rect 4395 2036 4403 2116
rect 4456 2107 4463 2133
rect 4496 2107 4503 2233
rect 4536 2127 4543 2153
rect 4453 2093 4467 2107
rect 4436 2027 4443 2093
rect 4556 2087 4563 2193
rect 4576 2147 4583 2253
rect 4596 2247 4603 2353
rect 4633 2253 4647 2267
rect 4596 2087 4603 2193
rect 4636 2147 4643 2253
rect 4676 2147 4683 2393
rect 4736 2347 4743 2516
rect 4756 2387 4763 2613
rect 4796 2567 4803 2633
rect 4773 2533 4787 2547
rect 4793 2553 4807 2567
rect 4776 2527 4783 2533
rect 4816 2423 4823 2473
rect 4796 2416 4823 2423
rect 4716 2287 4723 2333
rect 4756 2303 4763 2373
rect 4736 2296 4763 2303
rect 4736 2287 4743 2296
rect 4693 2253 4707 2267
rect 4713 2273 4727 2287
rect 4733 2273 4747 2287
rect 4716 2127 4723 2213
rect 4776 2207 4783 2353
rect 4796 2287 4803 2416
rect 4793 2273 4807 2287
rect 4513 2083 4527 2087
rect 4473 2063 4487 2067
rect 4496 2076 4527 2083
rect 4496 2063 4503 2076
rect 4473 2056 4503 2063
rect 4513 2073 4527 2076
rect 4473 2053 4487 2056
rect 4533 2053 4547 2067
rect 4553 2073 4567 2087
rect 4573 2053 4587 2067
rect 4593 2073 4607 2087
rect 4395 1998 4403 2022
rect 4436 1967 4443 1993
rect 4336 1847 4343 1913
rect 4316 1816 4343 1823
rect 4153 1773 4167 1787
rect 4193 1773 4207 1787
rect 4213 1773 4227 1787
rect 4233 1793 4247 1807
rect 4273 1803 4287 1807
rect 4273 1796 4293 1803
rect 4273 1793 4287 1796
rect 4253 1773 4267 1787
rect 4173 1753 4187 1767
rect 4156 1687 4163 1753
rect 4176 1747 4183 1753
rect 4196 1707 4203 1773
rect 4216 1683 4223 1773
rect 4256 1727 4263 1773
rect 4196 1676 4223 1683
rect 4153 1603 4167 1607
rect 4176 1603 4183 1673
rect 4153 1596 4183 1603
rect 4153 1593 4167 1596
rect 4136 1556 4163 1563
rect 4036 1264 4044 1376
rect 4056 1207 4063 1473
rect 4056 1167 4063 1193
rect 4076 1147 4083 1393
rect 4156 1387 4163 1556
rect 4196 1507 4203 1676
rect 4215 1556 4223 1636
rect 4256 1587 4263 1693
rect 4215 1518 4223 1542
rect 4256 1447 4263 1573
rect 4276 1443 4283 1773
rect 4296 1747 4303 1773
rect 4296 1607 4303 1633
rect 4293 1593 4307 1607
rect 4313 1573 4327 1587
rect 4316 1527 4323 1573
rect 4336 1567 4343 1816
rect 4356 1807 4363 1853
rect 4396 1823 4403 1933
rect 4456 1867 4463 2053
rect 4536 2047 4543 2053
rect 4576 2047 4583 2053
rect 4616 2047 4623 2093
rect 4633 2073 4647 2087
rect 4476 1887 4483 1933
rect 4387 1816 4403 1823
rect 4353 1793 4367 1807
rect 4393 1783 4407 1787
rect 4376 1776 4407 1783
rect 4413 1793 4427 1807
rect 4453 1793 4467 1807
rect 4356 1627 4363 1753
rect 4376 1727 4383 1776
rect 4393 1773 4407 1776
rect 4456 1767 4463 1793
rect 4476 1787 4483 1833
rect 4396 1747 4403 1753
rect 4353 1593 4367 1607
rect 4373 1573 4387 1587
rect 4376 1547 4383 1573
rect 4396 1487 4403 1653
rect 4416 1607 4423 1633
rect 4413 1593 4427 1607
rect 4433 1573 4447 1587
rect 4276 1436 4303 1443
rect 4137 1358 4145 1382
rect 4113 1293 4127 1307
rect 4096 1263 4103 1293
rect 4137 1264 4145 1344
rect 4096 1256 4123 1263
rect 4096 1147 4103 1173
rect 4116 1147 4123 1256
rect 4156 1187 4163 1213
rect 4176 1167 4183 1433
rect 4236 1347 4243 1413
rect 4193 1293 4207 1307
rect 4233 1293 4247 1307
rect 4196 1287 4203 1293
rect 4236 1227 4243 1293
rect 4156 1147 4163 1153
rect 4093 1133 4107 1147
rect 3996 1127 4003 1133
rect 3993 1113 4007 1127
rect 4013 1093 4027 1107
rect 3995 878 4003 902
rect 4016 867 4023 1093
rect 4036 1027 4043 1133
rect 4196 1127 4203 1133
rect 4193 1113 4207 1127
rect 4213 1093 4227 1107
rect 3995 784 4003 864
rect 4036 807 4043 993
rect 4056 847 4063 953
rect 4116 847 4123 1033
rect 4136 927 4143 1053
rect 4176 967 4183 1093
rect 4216 927 4223 1093
rect 4256 907 4263 1433
rect 4276 1264 4284 1376
rect 4296 1267 4303 1436
rect 4336 1367 4343 1473
rect 4316 1227 4323 1353
rect 4416 1347 4423 1473
rect 4436 1347 4443 1573
rect 4456 1427 4463 1693
rect 4476 1667 4483 1753
rect 4496 1707 4503 2033
rect 4536 1947 4543 2033
rect 4553 1773 4567 1787
rect 4576 1783 4583 1833
rect 4636 1823 4643 1933
rect 4656 1847 4663 2053
rect 4696 1947 4703 2053
rect 4716 1887 4723 2113
rect 4756 2087 4763 2173
rect 4816 2103 4823 2193
rect 4836 2127 4843 2693
rect 4856 2687 4863 2733
rect 4876 2647 4883 2733
rect 4896 2687 4903 2893
rect 4936 2827 4943 2896
rect 4916 2727 4923 2793
rect 4936 2787 4943 2813
rect 4933 2733 4947 2747
rect 4916 2667 4923 2693
rect 4853 2553 4867 2567
rect 4877 2516 4885 2596
rect 4856 2303 4863 2513
rect 4877 2478 4885 2502
rect 4896 2367 4903 2593
rect 4856 2296 4883 2303
rect 4876 2287 4883 2296
rect 4853 2253 4867 2267
rect 4856 2223 4863 2253
rect 4893 2253 4907 2267
rect 4873 2233 4887 2247
rect 4916 2243 4923 2653
rect 4976 2567 4983 2673
rect 4973 2553 4987 2567
rect 4956 2447 4963 2553
rect 4996 2443 5003 2913
rect 5016 2847 5023 3013
rect 5036 2787 5043 2993
rect 5056 2787 5063 2893
rect 5096 2867 5103 3036
rect 5133 3013 5147 3027
rect 5116 2767 5123 2773
rect 5136 2767 5143 3013
rect 5156 3007 5163 3133
rect 5176 3047 5183 3253
rect 5193 3223 5207 3227
rect 5216 3223 5223 3273
rect 5193 3216 5223 3223
rect 5193 3213 5207 3216
rect 5236 3184 5244 3296
rect 5173 3033 5187 3047
rect 5216 3047 5223 3173
rect 5256 3143 5263 3233
rect 5276 3227 5283 3453
rect 5356 3444 5364 3556
rect 5376 3427 5383 3733
rect 5433 3513 5447 3527
rect 5436 3507 5443 3513
rect 5457 3476 5465 3556
rect 5457 3438 5465 3462
rect 5236 3136 5263 3143
rect 5213 3033 5227 3047
rect 5236 3003 5243 3136
rect 5276 3047 5283 3213
rect 5296 3167 5303 3353
rect 5316 3247 5323 3313
rect 5496 3307 5503 3913
rect 5556 3887 5563 3953
rect 5616 3867 5623 4036
rect 5636 3967 5643 4153
rect 5696 4127 5703 4173
rect 5656 3924 5664 4036
rect 5696 4007 5703 4093
rect 5693 3993 5707 4007
rect 5733 4003 5747 4007
rect 5676 3967 5683 3993
rect 5716 3996 5747 4003
rect 5557 3758 5565 3782
rect 5516 3727 5523 3753
rect 5516 3547 5523 3713
rect 5557 3664 5565 3744
rect 5596 3703 5603 3753
rect 5613 3703 5627 3707
rect 5596 3696 5627 3703
rect 5613 3693 5627 3696
rect 5516 3527 5523 3533
rect 5513 3513 5527 3527
rect 5553 3523 5567 3527
rect 5553 3516 5583 3523
rect 5553 3513 5567 3516
rect 5576 3507 5583 3516
rect 5476 3283 5483 3293
rect 5476 3276 5503 3283
rect 5496 3267 5503 3276
rect 5416 3247 5423 3253
rect 5313 3233 5327 3247
rect 5413 3233 5427 3247
rect 5373 3213 5387 3227
rect 5376 3207 5383 3213
rect 5336 3167 5343 3193
rect 5376 3167 5383 3193
rect 5216 2996 5243 3003
rect 5156 2827 5163 2973
rect 5176 2783 5183 2973
rect 5216 2847 5223 2996
rect 5236 2807 5243 2913
rect 5256 2807 5263 3013
rect 5176 2776 5193 2783
rect 5073 2753 5087 2767
rect 5113 2753 5127 2767
rect 5173 2733 5187 2747
rect 5176 2727 5183 2733
rect 5133 2713 5147 2727
rect 5036 2667 5043 2713
rect 5016 2484 5024 2596
rect 5036 2447 5043 2573
rect 4996 2436 5023 2443
rect 4936 2287 4943 2333
rect 4933 2273 4947 2287
rect 4953 2253 4967 2267
rect 4976 2243 4983 2433
rect 4996 2287 5003 2373
rect 5016 2307 5023 2436
rect 4993 2273 5007 2287
rect 5013 2253 5027 2267
rect 5016 2243 5023 2253
rect 4896 2236 4923 2243
rect 4956 2236 4983 2243
rect 4996 2236 5023 2243
rect 4856 2216 4883 2223
rect 4876 2207 4883 2216
rect 4876 2147 4883 2193
rect 4853 2103 4867 2107
rect 4816 2096 4867 2103
rect 4753 2073 4767 2087
rect 4773 2053 4787 2067
rect 4756 2027 4763 2033
rect 4636 1816 4663 1823
rect 4656 1807 4663 1816
rect 4593 1783 4607 1787
rect 4576 1776 4607 1783
rect 4593 1773 4607 1776
rect 4633 1773 4647 1787
rect 4653 1793 4667 1807
rect 4516 1627 4523 1653
rect 4536 1607 4543 1733
rect 4556 1667 4563 1773
rect 4576 1643 4583 1713
rect 4596 1687 4603 1753
rect 4636 1687 4643 1773
rect 4696 1747 4703 1853
rect 4716 1823 4723 1833
rect 4716 1816 4743 1823
rect 4736 1807 4743 1816
rect 4756 1807 4763 2013
rect 4816 2007 4823 2096
rect 4853 2093 4867 2096
rect 4876 2087 4883 2133
rect 4896 2107 4903 2236
rect 4956 2107 4963 2236
rect 4976 2187 4983 2213
rect 4996 2167 5003 2236
rect 4873 2073 4887 2087
rect 4913 2053 4927 2067
rect 4933 2073 4947 2087
rect 4953 2053 4967 2067
rect 4856 1907 4863 2053
rect 4876 1907 4883 1933
rect 4797 1838 4805 1862
rect 4773 1783 4787 1787
rect 4733 1763 4747 1767
rect 4756 1776 4787 1783
rect 4756 1763 4763 1776
rect 4733 1756 4763 1763
rect 4773 1773 4787 1776
rect 4733 1753 4747 1756
rect 4556 1636 4583 1643
rect 4473 1593 4487 1607
rect 4493 1583 4507 1587
rect 4513 1583 4527 1587
rect 4493 1576 4527 1583
rect 4493 1573 4507 1576
rect 4513 1573 4527 1576
rect 4496 1547 4503 1573
rect 4476 1523 4483 1533
rect 4476 1516 4503 1523
rect 4496 1427 4503 1516
rect 4556 1507 4563 1636
rect 4596 1607 4603 1653
rect 4716 1627 4723 1653
rect 4716 1607 4723 1613
rect 4573 1573 4587 1587
rect 4593 1593 4607 1607
rect 4633 1573 4647 1587
rect 4713 1593 4727 1607
rect 4336 1307 4343 1333
rect 4456 1327 4463 1353
rect 4433 1293 4447 1307
rect 4453 1313 4467 1327
rect 4473 1303 4487 1307
rect 4473 1296 4503 1303
rect 4473 1293 4487 1296
rect 4373 1273 4387 1287
rect 4296 1203 4303 1213
rect 4356 1203 4363 1273
rect 4296 1196 4363 1203
rect 4276 1156 4323 1163
rect 4276 1147 4283 1156
rect 4273 1113 4287 1127
rect 4316 1127 4323 1156
rect 4396 1147 4403 1293
rect 4436 1287 4443 1293
rect 4313 1113 4327 1127
rect 4356 1047 4363 1133
rect 4436 1127 4443 1253
rect 4496 1247 4503 1296
rect 4527 1276 4543 1283
rect 4476 1127 4483 1213
rect 4516 1147 4523 1233
rect 4536 1147 4543 1276
rect 4513 1133 4527 1147
rect 4433 1123 4447 1127
rect 4413 1093 4427 1107
rect 4433 1116 4463 1123
rect 4433 1113 4447 1116
rect 4456 1107 4463 1116
rect 4473 1113 4487 1127
rect 4533 1093 4547 1107
rect 4316 927 4323 1033
rect 4336 927 4343 973
rect 4416 967 4423 1093
rect 4456 987 4463 1073
rect 4256 867 4263 873
rect 4053 833 4067 847
rect 4113 833 4127 847
rect 4076 767 4083 813
rect 3896 667 3903 693
rect 3896 627 3903 653
rect 3833 593 3847 607
rect 3853 613 3867 627
rect 3893 613 3907 627
rect 3873 593 3887 607
rect 3756 567 3763 593
rect 3836 567 3843 593
rect 3676 407 3683 553
rect 3716 536 3783 543
rect 3716 527 3723 536
rect 3716 387 3723 473
rect 3736 387 3743 513
rect 3296 267 3303 333
rect 3336 227 3343 333
rect 3356 287 3363 333
rect 3393 336 3423 343
rect 3393 333 3407 336
rect 3473 353 3487 367
rect 3513 353 3527 367
rect 3533 333 3547 347
rect 3553 353 3567 367
rect 3593 353 3607 367
rect 3573 333 3587 347
rect 3536 327 3543 333
rect 3373 313 3387 327
rect 3376 267 3383 313
rect 3253 183 3267 187
rect 3253 176 3283 183
rect 3253 173 3267 176
rect 3073 153 3087 167
rect 3113 153 3127 167
rect 3153 153 3167 167
rect 3193 163 3207 167
rect 3173 133 3187 147
rect 3193 156 3223 163
rect 3193 153 3207 156
rect 3216 143 3223 156
rect 3276 163 3283 176
rect 3293 163 3307 167
rect 3276 156 3307 163
rect 3293 153 3307 156
rect 3233 143 3247 147
rect 3216 136 3247 143
rect 3233 133 3247 136
rect 2855 78 2863 102
rect 2976 47 2983 133
rect 3176 107 3183 133
rect 3317 116 3325 196
rect 3373 163 3387 167
rect 3396 163 3403 293
rect 3416 267 3423 313
rect 3416 167 3423 193
rect 3373 156 3403 163
rect 3373 153 3387 156
rect 3413 153 3427 167
rect 3317 78 3325 102
rect 3456 84 3464 196
rect 3496 127 3503 313
rect 3536 267 3543 293
rect 3516 123 3523 233
rect 3556 167 3563 313
rect 3576 227 3583 333
rect 3596 307 3603 353
rect 3713 363 3727 367
rect 3736 363 3743 373
rect 3756 367 3763 413
rect 3776 387 3783 536
rect 3673 333 3687 347
rect 3713 356 3743 363
rect 3713 353 3727 356
rect 3753 353 3767 367
rect 3676 327 3683 333
rect 3773 343 3787 347
rect 3796 343 3803 373
rect 3856 367 3863 453
rect 3916 407 3923 673
rect 3957 596 3965 676
rect 3957 558 3965 582
rect 3936 387 3943 493
rect 3976 367 3983 713
rect 3996 643 4003 733
rect 4016 647 4023 653
rect 4056 647 4063 753
rect 4096 743 4103 833
rect 4156 803 4163 853
rect 4216 847 4223 853
rect 4213 833 4227 847
rect 4076 736 4103 743
rect 4136 796 4163 803
rect 4013 643 4027 647
rect 3996 636 4027 643
rect 3773 336 3803 343
rect 3773 333 3787 336
rect 3833 333 3847 347
rect 3933 333 3947 347
rect 3653 313 3667 327
rect 3853 313 3867 327
rect 3596 167 3603 173
rect 3616 167 3623 193
rect 3636 167 3643 213
rect 3656 207 3663 313
rect 3756 187 3763 293
rect 3633 153 3647 167
rect 3533 123 3547 127
rect 3516 116 3547 123
rect 3573 123 3587 127
rect 3596 123 3603 153
rect 3533 113 3547 116
rect 3573 116 3603 123
rect 3653 133 3667 147
rect 3693 153 3707 167
rect 3756 147 3763 173
rect 3753 133 3767 147
rect 3656 127 3663 133
rect 3573 113 3587 116
rect 3776 87 3783 313
rect 3796 147 3803 313
rect 3856 287 3863 313
rect 3876 207 3883 333
rect 3896 267 3903 293
rect 3936 267 3943 333
rect 3956 287 3963 333
rect 3996 307 4003 636
rect 4013 633 4027 636
rect 4053 633 4067 647
rect 4076 527 4083 736
rect 4096 564 4104 676
rect 4016 387 4023 493
rect 4136 427 4143 796
rect 4176 763 4183 793
rect 4156 756 4183 763
rect 4156 507 4163 756
rect 4196 667 4203 693
rect 4193 653 4207 667
rect 4173 633 4187 647
rect 4213 633 4227 647
rect 4156 407 4163 473
rect 4013 373 4027 387
rect 4053 373 4067 387
rect 4073 353 4087 367
rect 4076 327 4083 353
rect 4093 333 4107 347
rect 3813 153 3827 167
rect 3816 127 3823 153
rect 3837 116 3845 196
rect 3896 167 3903 253
rect 3936 167 3943 213
rect 4096 207 4103 333
rect 4133 333 4147 347
rect 4136 327 4143 333
rect 4113 313 4127 327
rect 3893 153 3907 167
rect 3933 153 3947 167
rect 3837 78 3845 102
rect 3976 84 3984 196
rect 4033 163 4047 167
rect 4016 156 4047 163
rect 4016 87 4023 156
rect 4033 153 4047 156
rect 4096 147 4103 173
rect 4116 147 4123 313
rect 4176 227 4183 533
rect 4196 347 4203 593
rect 4217 398 4225 422
rect 4217 304 4225 384
rect 4236 287 4243 773
rect 4256 707 4263 833
rect 4313 813 4327 827
rect 4316 807 4323 813
rect 4256 227 4263 633
rect 4277 596 4285 676
rect 4336 667 4343 793
rect 4356 667 4363 893
rect 4376 747 4383 953
rect 4496 947 4503 1093
rect 4516 1007 4523 1073
rect 4433 853 4447 867
rect 4413 833 4427 847
rect 4453 843 4467 847
rect 4436 836 4467 843
rect 4336 647 4343 653
rect 4356 647 4363 653
rect 4376 647 4383 693
rect 4333 633 4347 647
rect 4373 633 4387 647
rect 4277 558 4285 582
rect 4273 333 4287 347
rect 4276 307 4283 333
rect 4296 327 4303 493
rect 4313 333 4327 347
rect 4316 267 4323 333
rect 4176 167 4183 193
rect 4216 167 4223 213
rect 4093 133 4107 147
rect 4173 153 4187 167
rect 4056 67 4063 133
rect 4216 123 4223 153
rect 4233 123 4247 127
rect 4216 116 4247 123
rect 4273 123 4287 127
rect 4296 123 4303 233
rect 4336 203 4343 453
rect 4396 423 4403 813
rect 4416 727 4423 833
rect 4436 767 4443 836
rect 4453 833 4467 836
rect 4416 564 4424 676
rect 4376 416 4403 423
rect 4356 304 4364 416
rect 4233 113 4247 116
rect 4273 116 4303 123
rect 4316 196 4343 203
rect 4273 113 4287 116
rect 4316 47 4323 196
rect 4357 116 4365 196
rect 4357 78 4365 102
rect 4376 87 4383 416
rect 4396 307 4403 393
rect 4436 387 4443 733
rect 4456 627 4463 733
rect 4516 567 4523 953
rect 4536 887 4543 1093
rect 4556 1067 4563 1493
rect 4576 1347 4583 1573
rect 4636 1507 4643 1573
rect 4736 1563 4743 1733
rect 4756 1647 4763 1756
rect 4797 1744 4805 1824
rect 4816 1667 4823 1833
rect 4876 1787 4883 1853
rect 4896 1823 4903 2033
rect 4956 2007 4963 2053
rect 5016 2043 5023 2213
rect 5036 2087 5043 2413
rect 5056 2227 5063 2613
rect 5076 2607 5083 2713
rect 5073 2573 5087 2587
rect 5116 2367 5123 2633
rect 5176 2567 5183 2673
rect 5196 2667 5203 2753
rect 5213 2733 5227 2747
rect 5236 2707 5243 2773
rect 5253 2733 5267 2747
rect 5256 2647 5263 2733
rect 5276 2727 5283 2993
rect 5296 2964 5304 3076
rect 5316 3067 5323 3093
rect 5376 3063 5383 3113
rect 5396 3087 5403 3233
rect 5376 3056 5403 3063
rect 5333 3043 5347 3047
rect 5316 3036 5347 3043
rect 5316 2987 5323 3036
rect 5333 3033 5347 3036
rect 5396 3003 5403 3056
rect 5376 2996 5403 3003
rect 5293 2733 5307 2747
rect 5333 2743 5347 2747
rect 5333 2736 5353 2743
rect 5333 2733 5347 2736
rect 5236 2616 5283 2623
rect 5236 2603 5243 2616
rect 5276 2607 5283 2616
rect 5216 2596 5243 2603
rect 5216 2567 5223 2596
rect 5153 2533 5167 2547
rect 5173 2553 5187 2567
rect 5213 2553 5227 2567
rect 5236 2547 5243 2573
rect 5296 2567 5303 2573
rect 5293 2553 5307 2567
rect 5316 2547 5323 2573
rect 5336 2547 5343 2713
rect 5356 2587 5363 2713
rect 5376 2687 5383 2996
rect 5416 2987 5423 3133
rect 5435 2996 5443 3076
rect 5435 2958 5443 2982
rect 5456 2827 5463 2953
rect 5476 2947 5483 3253
rect 5513 3203 5527 3207
rect 5536 3203 5543 3353
rect 5513 3196 5543 3203
rect 5513 3193 5527 3196
rect 5556 3167 5563 3473
rect 5596 3444 5604 3556
rect 5616 3347 5623 3513
rect 5636 3467 5643 3913
rect 5696 3664 5704 3776
rect 5716 3767 5723 3996
rect 5733 3993 5747 3996
rect 5756 3567 5763 4213
rect 5816 4167 5823 4813
rect 5836 4803 5843 4893
rect 5876 4867 5883 4893
rect 5856 4827 5863 4853
rect 5916 4847 5923 4873
rect 5936 4847 5943 5113
rect 5976 4967 5983 5073
rect 6016 5047 6023 5133
rect 6036 4987 6043 5293
rect 6096 5207 6103 5253
rect 6096 5187 6103 5193
rect 6093 5173 6107 5187
rect 6056 5087 6063 5133
rect 6116 5127 6123 5293
rect 6136 5107 6143 5393
rect 6176 5387 6183 5453
rect 6196 5407 6203 6096
rect 6236 6067 6243 6093
rect 6216 5807 6223 5973
rect 6236 5947 6243 6053
rect 6256 6027 6263 6113
rect 6276 6067 6283 6113
rect 6316 6047 6323 6173
rect 6456 6167 6463 6353
rect 6556 6287 6563 6373
rect 6576 6347 6583 6413
rect 6596 6407 6603 6433
rect 6636 6407 6643 6413
rect 6593 6393 6607 6407
rect 6613 6373 6627 6387
rect 6633 6393 6647 6407
rect 6616 6367 6623 6373
rect 6353 6143 6367 6147
rect 6336 6136 6367 6143
rect 6336 6007 6343 6136
rect 6353 6133 6367 6136
rect 6413 6113 6427 6127
rect 6273 5873 6287 5887
rect 6216 5447 6223 5673
rect 6236 5647 6243 5653
rect 6256 5647 6263 5793
rect 6276 5787 6283 5873
rect 6316 5867 6323 5953
rect 6336 5927 6343 5973
rect 6333 5873 6347 5887
rect 6376 5883 6383 6073
rect 6416 6047 6423 6113
rect 6436 6083 6443 6133
rect 6516 6127 6523 6133
rect 6513 6113 6527 6127
rect 6436 6076 6463 6083
rect 6396 5927 6403 5953
rect 6436 5927 6443 6013
rect 6456 5927 6463 6076
rect 6613 6123 6627 6127
rect 6613 6116 6643 6123
rect 6613 6113 6627 6116
rect 6533 6073 6547 6087
rect 6593 6073 6607 6087
rect 6536 6067 6543 6073
rect 6476 5927 6483 5933
rect 6393 5913 6407 5927
rect 6413 5893 6427 5907
rect 6433 5913 6447 5927
rect 6496 5907 6503 6053
rect 6576 5907 6583 6033
rect 6596 5987 6603 6073
rect 6636 5947 6643 6116
rect 6453 5903 6467 5907
rect 6493 5903 6507 5907
rect 6453 5896 6507 5903
rect 6453 5893 6467 5896
rect 6376 5876 6393 5883
rect 6336 5787 6343 5873
rect 6276 5647 6283 5693
rect 6336 5667 6343 5753
rect 6356 5707 6363 5873
rect 6376 5683 6383 5813
rect 6416 5767 6423 5893
rect 6456 5707 6463 5853
rect 6476 5687 6483 5896
rect 6493 5893 6507 5896
rect 6516 5887 6523 5893
rect 6513 5873 6527 5887
rect 6633 5873 6647 5887
rect 6496 5727 6503 5833
rect 6356 5676 6383 5683
rect 6356 5667 6363 5676
rect 6316 5647 6323 5653
rect 6393 5653 6407 5667
rect 6233 5633 6247 5647
rect 6253 5593 6267 5607
rect 6293 5593 6307 5607
rect 6256 5467 6263 5593
rect 6276 5527 6283 5593
rect 6296 5587 6303 5593
rect 6296 5547 6303 5573
rect 6236 5447 6243 5453
rect 6276 5447 6283 5473
rect 6296 5467 6303 5493
rect 6316 5467 6323 5593
rect 6356 5567 6363 5593
rect 6336 5447 6343 5533
rect 6233 5433 6247 5447
rect 6273 5443 6287 5447
rect 6293 5443 6307 5447
rect 6216 5427 6223 5433
rect 6273 5436 6307 5443
rect 6273 5433 6287 5436
rect 6293 5433 6307 5436
rect 6333 5433 6347 5447
rect 6356 5427 6363 5433
rect 6176 5167 6183 5193
rect 6196 5187 6203 5213
rect 6236 5187 6243 5393
rect 6256 5167 6263 5193
rect 6276 5187 6283 5213
rect 6153 5133 6167 5147
rect 6173 5153 6187 5167
rect 6213 5163 6227 5167
rect 6213 5156 6243 5163
rect 6213 5153 6227 5156
rect 6156 5107 6163 5133
rect 6236 5147 6243 5156
rect 6253 5153 6267 5167
rect 6236 5107 6243 5113
rect 6116 5087 6123 5093
rect 6076 5027 6083 5073
rect 6096 4967 6103 5013
rect 6116 4967 6123 5033
rect 6013 4963 6027 4967
rect 6007 4956 6027 4963
rect 6013 4953 6027 4956
rect 5953 4913 5967 4927
rect 6033 4933 6047 4947
rect 6073 4933 6087 4947
rect 6093 4953 6107 4967
rect 5956 4907 5963 4913
rect 5836 4796 5863 4803
rect 5836 4687 5843 4693
rect 5856 4687 5863 4796
rect 5996 4787 6003 4913
rect 6016 4827 6023 4913
rect 6036 4907 6043 4933
rect 6076 4927 6083 4933
rect 5893 4693 5907 4707
rect 5833 4673 5847 4687
rect 5873 4673 5887 4687
rect 5853 4643 5867 4647
rect 5876 4643 5883 4673
rect 5853 4636 5883 4643
rect 5853 4633 5867 4636
rect 5856 4607 5863 4633
rect 5896 4567 5903 4693
rect 5956 4687 5963 4773
rect 6016 4707 6023 4753
rect 6013 4693 6027 4707
rect 5976 4667 5983 4693
rect 5993 4653 6007 4667
rect 5916 4527 5923 4653
rect 5853 4463 5867 4467
rect 5876 4463 5883 4473
rect 5896 4467 5903 4513
rect 5936 4487 5943 4533
rect 5996 4527 6003 4653
rect 6016 4507 6023 4553
rect 6013 4493 6027 4507
rect 6036 4503 6043 4873
rect 6056 4707 6063 4913
rect 6116 4863 6123 4933
rect 6136 4923 6143 5053
rect 6276 5047 6283 5093
rect 6156 4967 6163 4993
rect 6196 4947 6203 4993
rect 6216 4947 6223 5013
rect 6236 4967 6243 4973
rect 6276 4967 6283 4993
rect 6296 4987 6303 5393
rect 6376 5387 6383 5593
rect 6396 5587 6403 5653
rect 6413 5633 6427 5647
rect 6456 5643 6463 5673
rect 6536 5667 6543 5693
rect 6493 5653 6507 5667
rect 6473 5643 6487 5647
rect 6456 5636 6487 5643
rect 6473 5633 6487 5636
rect 6416 5527 6423 5633
rect 6456 5607 6463 5613
rect 6496 5587 6503 5653
rect 6513 5633 6527 5647
rect 6533 5653 6547 5667
rect 6556 5643 6563 5833
rect 6576 5687 6583 5873
rect 6596 5827 6603 5853
rect 6616 5687 6623 5713
rect 6636 5667 6643 5873
rect 6656 5807 6663 6313
rect 6633 5663 6647 5667
rect 6573 5643 6587 5647
rect 6556 5636 6587 5643
rect 6573 5633 6587 5636
rect 6613 5633 6627 5647
rect 6633 5656 6663 5663
rect 6633 5653 6647 5656
rect 6396 5427 6403 5453
rect 6416 5447 6423 5473
rect 6436 5447 6443 5553
rect 6516 5527 6523 5633
rect 6476 5447 6483 5453
rect 6433 5433 6447 5447
rect 6473 5433 6487 5447
rect 6316 5187 6323 5273
rect 6356 5227 6363 5353
rect 6376 5227 6383 5233
rect 6396 5207 6403 5393
rect 6416 5227 6423 5353
rect 6436 5203 6443 5233
rect 6496 5207 6503 5453
rect 6516 5447 6523 5493
rect 6536 5487 6543 5613
rect 6556 5467 6563 5613
rect 6576 5447 6583 5453
rect 6536 5436 6553 5443
rect 6536 5427 6543 5436
rect 6596 5407 6603 5633
rect 6616 5547 6623 5633
rect 6636 5463 6643 5493
rect 6656 5467 6663 5656
rect 6676 5467 6683 6333
rect 6696 6327 6703 6433
rect 6616 5456 6643 5463
rect 6616 5447 6623 5456
rect 6613 5433 6627 5447
rect 6673 5423 6687 5427
rect 6656 5416 6687 5423
rect 6416 5196 6443 5203
rect 6396 5187 6403 5193
rect 6416 5187 6423 5196
rect 6313 5173 6327 5187
rect 6316 4967 6323 5133
rect 6356 5127 6363 5173
rect 6413 5173 6427 5187
rect 6373 5153 6387 5167
rect 6516 5167 6523 5213
rect 6376 5147 6383 5153
rect 6376 5127 6383 5133
rect 6233 4953 6247 4967
rect 6153 4923 6167 4927
rect 6136 4916 6167 4923
rect 6213 4933 6227 4947
rect 6273 4953 6287 4967
rect 6296 4947 6303 4953
rect 6293 4933 6307 4947
rect 6153 4913 6167 4916
rect 6136 4887 6143 4893
rect 6116 4856 6143 4863
rect 6136 4747 6143 4856
rect 6156 4747 6163 4793
rect 6096 4687 6103 4733
rect 6073 4653 6087 4667
rect 6093 4673 6107 4687
rect 6133 4683 6147 4687
rect 6156 4683 6163 4713
rect 6133 4676 6163 4683
rect 6133 4673 6147 4676
rect 6056 4527 6063 4653
rect 6076 4643 6083 4653
rect 6076 4636 6103 4643
rect 6036 4496 6063 4503
rect 5996 4487 6003 4493
rect 5853 4456 5883 4463
rect 5853 4453 5867 4456
rect 5893 4453 5907 4467
rect 5973 4453 5987 4467
rect 5993 4473 6007 4487
rect 5976 4447 5983 4453
rect 5856 4247 5863 4413
rect 5916 4407 5923 4433
rect 5876 4263 5883 4393
rect 5876 4256 5903 4263
rect 5896 4243 5903 4256
rect 5896 4236 5923 4243
rect 5916 4227 5923 4236
rect 5853 4193 5867 4207
rect 5893 4193 5907 4207
rect 5913 4213 5927 4227
rect 5836 4147 5843 4173
rect 5776 3947 5783 4093
rect 5856 4067 5863 4193
rect 5795 3956 5803 4036
rect 5856 4027 5863 4053
rect 5853 4013 5867 4027
rect 5876 4023 5883 4193
rect 5896 4107 5903 4193
rect 5916 4127 5923 4133
rect 5936 4123 5943 4233
rect 5956 4207 5963 4213
rect 5996 4207 6003 4353
rect 6016 4327 6023 4453
rect 6036 4447 6043 4453
rect 6056 4347 6063 4496
rect 6076 4387 6083 4553
rect 6096 4507 6103 4636
rect 6136 4627 6143 4673
rect 6156 4527 6163 4653
rect 6113 4503 6127 4507
rect 6113 4496 6143 4503
rect 6113 4493 6127 4496
rect 6136 4467 6143 4496
rect 6176 4483 6183 4773
rect 6196 4707 6203 4713
rect 6193 4693 6207 4707
rect 6256 4687 6263 4713
rect 6276 4687 6283 4873
rect 6296 4807 6303 4873
rect 6296 4747 6303 4753
rect 6296 4687 6303 4733
rect 6316 4707 6323 4953
rect 6336 4927 6343 5033
rect 6396 5027 6403 5153
rect 6436 5147 6443 5153
rect 6416 4947 6423 4953
rect 6413 4933 6427 4947
rect 6336 4747 6343 4893
rect 6436 4803 6443 4993
rect 6476 4967 6483 5153
rect 6536 5107 6543 5373
rect 6556 5227 6563 5353
rect 6596 5207 6603 5393
rect 6636 5367 6643 5413
rect 6656 5407 6663 5416
rect 6673 5413 6687 5416
rect 6676 5207 6683 5393
rect 6556 5167 6563 5193
rect 6696 5187 6703 5893
rect 6716 5207 6723 6353
rect 6593 5153 6607 5167
rect 6693 5183 6707 5187
rect 6673 5153 6687 5167
rect 6693 5176 6723 5183
rect 6693 5173 6707 5176
rect 6556 5007 6563 5133
rect 6596 5107 6603 5153
rect 6453 4913 6467 4927
rect 6496 4927 6503 4993
rect 6576 4987 6583 5093
rect 6616 5007 6623 5153
rect 6516 4947 6523 4953
rect 6556 4947 6563 4953
rect 6513 4933 6527 4947
rect 6553 4933 6567 4947
rect 6573 4923 6587 4927
rect 6596 4923 6603 4993
rect 6636 4983 6643 5153
rect 6656 5007 6663 5133
rect 6676 5127 6683 5153
rect 6716 5147 6723 5176
rect 6653 4983 6667 4987
rect 6636 4976 6683 4983
rect 6653 4973 6667 4976
rect 6616 4943 6623 4973
rect 6633 4943 6647 4947
rect 6616 4936 6647 4943
rect 6633 4933 6647 4936
rect 6636 4927 6643 4933
rect 6573 4916 6603 4923
rect 6573 4913 6587 4916
rect 6456 4867 6463 4913
rect 6436 4796 6463 4803
rect 6253 4673 6267 4687
rect 6293 4673 6307 4687
rect 6313 4653 6327 4667
rect 6156 4476 6183 4483
rect 6093 4453 6107 4467
rect 6133 4463 6147 4467
rect 6116 4456 6147 4463
rect 6096 4407 6103 4453
rect 6116 4427 6123 4456
rect 6133 4453 6147 4456
rect 6156 4447 6163 4476
rect 6153 4433 6167 4447
rect 6193 4433 6207 4447
rect 6196 4427 6203 4433
rect 6216 4367 6223 4573
rect 6236 4427 6243 4593
rect 6276 4587 6283 4633
rect 6316 4547 6323 4653
rect 6336 4607 6343 4733
rect 6356 4727 6363 4753
rect 6416 4707 6423 4713
rect 6353 4673 6367 4687
rect 6393 4683 6407 4687
rect 6376 4676 6407 4683
rect 6413 4693 6427 4707
rect 6356 4587 6363 4673
rect 6376 4627 6383 4676
rect 6393 4673 6407 4676
rect 6436 4667 6443 4713
rect 6376 4563 6383 4593
rect 6356 4556 6383 4563
rect 6256 4507 6263 4533
rect 6256 4467 6263 4493
rect 6316 4487 6323 4533
rect 6356 4527 6363 4556
rect 6253 4453 6267 4467
rect 6293 4453 6307 4467
rect 6313 4473 6327 4487
rect 6336 4467 6343 4493
rect 6333 4453 6347 4467
rect 6296 4443 6303 4453
rect 6276 4436 6303 4443
rect 6276 4387 6283 4436
rect 6356 4447 6363 4473
rect 6376 4467 6383 4513
rect 6396 4487 6403 4653
rect 6436 4487 6443 4633
rect 6456 4627 6463 4796
rect 6476 4707 6483 4793
rect 6496 4707 6503 4773
rect 6473 4653 6487 4667
rect 6516 4663 6523 4733
rect 6536 4703 6543 4913
rect 6616 4747 6623 4913
rect 6636 4747 6643 4833
rect 6676 4727 6683 4976
rect 6536 4696 6563 4703
rect 6556 4667 6563 4696
rect 6613 4693 6627 4707
rect 6593 4673 6607 4687
rect 6533 4663 6547 4667
rect 6516 4656 6547 4663
rect 6533 4653 6547 4656
rect 6456 4527 6463 4613
rect 6476 4607 6483 4653
rect 6476 4503 6483 4553
rect 6456 4496 6483 4503
rect 6456 4467 6463 4496
rect 6496 4483 6503 4513
rect 6476 4476 6503 4483
rect 6476 4467 6483 4476
rect 6516 4467 6523 4633
rect 6556 4567 6563 4633
rect 6576 4487 6583 4513
rect 6373 4453 6387 4467
rect 6353 4433 6367 4447
rect 6473 4453 6487 4467
rect 6573 4473 6587 4487
rect 6596 4467 6603 4673
rect 6616 4627 6623 4693
rect 6633 4683 6647 4687
rect 6656 4683 6663 4713
rect 6633 4676 6663 4683
rect 6633 4673 6647 4676
rect 6616 4487 6623 4533
rect 6493 4433 6507 4447
rect 6036 4207 6043 4213
rect 6033 4193 6047 4207
rect 6053 4173 6067 4187
rect 5936 4116 5963 4123
rect 5876 4016 5903 4023
rect 5836 3967 5843 4013
rect 5873 3973 5887 3987
rect 5795 3918 5803 3942
rect 5856 3887 5863 3953
rect 5876 3947 5883 3973
rect 5896 3967 5903 4016
rect 5956 3987 5963 4116
rect 6016 4007 6023 4153
rect 6056 4107 6063 4173
rect 5953 3973 5967 3987
rect 5993 3983 6007 3987
rect 5993 3976 6023 3983
rect 5993 3973 6007 3976
rect 5796 3727 5803 3873
rect 5896 3756 5963 3763
rect 5896 3747 5903 3756
rect 5853 3743 5867 3747
rect 5833 3713 5847 3727
rect 5853 3736 5883 3743
rect 5853 3733 5867 3736
rect 5836 3687 5843 3713
rect 5793 3673 5807 3687
rect 5796 3627 5803 3673
rect 5876 3587 5883 3736
rect 5893 3733 5907 3747
rect 5656 3527 5663 3533
rect 5696 3527 5703 3553
rect 5673 3493 5687 3507
rect 5693 3513 5707 3527
rect 5716 3507 5723 3513
rect 5676 3487 5683 3493
rect 5576 3184 5584 3296
rect 5613 3213 5627 3227
rect 5516 3047 5523 3113
rect 5513 3043 5527 3047
rect 5496 3036 5527 3043
rect 5556 3047 5563 3133
rect 5576 3047 5583 3053
rect 5616 3047 5623 3213
rect 5636 3047 5643 3413
rect 5676 3327 5683 3473
rect 5696 3347 5703 3373
rect 5653 3213 5667 3227
rect 5656 3067 5663 3213
rect 5496 2927 5503 3036
rect 5513 3033 5527 3036
rect 5553 3033 5567 3047
rect 5573 3033 5587 3047
rect 5593 3013 5607 3027
rect 5613 3033 5627 3047
rect 5633 3023 5647 3027
rect 5633 3016 5653 3023
rect 5633 3013 5647 3016
rect 5536 3003 5543 3013
rect 5596 3007 5603 3013
rect 5536 2996 5563 3003
rect 5516 2883 5523 2973
rect 5496 2876 5523 2883
rect 5496 2807 5503 2876
rect 5396 2767 5403 2773
rect 5436 2767 5443 2773
rect 5413 2743 5427 2747
rect 5396 2736 5427 2743
rect 5433 2753 5447 2767
rect 5396 2667 5403 2736
rect 5413 2733 5427 2736
rect 5453 2733 5467 2747
rect 5456 2723 5463 2733
rect 5436 2716 5463 2723
rect 5436 2707 5443 2716
rect 5476 2687 5483 2713
rect 5376 2587 5383 2593
rect 5373 2573 5387 2587
rect 5353 2553 5367 2567
rect 5313 2533 5327 2547
rect 5393 2553 5407 2567
rect 5156 2507 5163 2533
rect 5196 2447 5203 2493
rect 5156 2327 5163 2353
rect 5176 2287 5183 2313
rect 5093 2273 5107 2287
rect 5133 2273 5147 2287
rect 5173 2273 5187 2287
rect 5113 2233 5127 2247
rect 5153 2233 5167 2247
rect 5156 2223 5163 2233
rect 5136 2216 5163 2223
rect 5056 2127 5063 2193
rect 5096 2147 5103 2213
rect 5136 2167 5143 2216
rect 5116 2087 5123 2133
rect 5156 2087 5163 2193
rect 5196 2147 5203 2433
rect 5256 2303 5263 2353
rect 5236 2296 5263 2303
rect 5236 2287 5243 2296
rect 5276 2287 5283 2313
rect 5296 2307 5303 2453
rect 5233 2273 5247 2287
rect 5253 2253 5267 2267
rect 5273 2273 5287 2287
rect 5293 2253 5307 2267
rect 5176 2107 5183 2133
rect 5173 2093 5187 2107
rect 5056 2067 5063 2073
rect 5033 2043 5047 2047
rect 5016 2036 5047 2043
rect 5053 2053 5067 2067
rect 5033 2033 5047 2036
rect 5073 2033 5087 2047
rect 4936 1927 4943 1993
rect 4976 1947 4983 2033
rect 5036 2027 5043 2033
rect 4976 1887 4983 1933
rect 4896 1816 4923 1823
rect 4853 1773 4867 1787
rect 4893 1773 4907 1787
rect 4856 1767 4863 1773
rect 4896 1743 4903 1773
rect 4916 1767 4923 1816
rect 4876 1736 4903 1743
rect 4876 1687 4883 1736
rect 4896 1687 4903 1713
rect 4773 1603 4787 1607
rect 4753 1573 4767 1587
rect 4773 1596 4803 1603
rect 4773 1593 4787 1596
rect 4716 1556 4743 1563
rect 4756 1563 4763 1573
rect 4796 1567 4803 1596
rect 4756 1556 4783 1563
rect 4656 1527 4663 1553
rect 4596 1427 4603 1493
rect 4716 1367 4723 1556
rect 4616 1347 4623 1353
rect 4616 1207 4623 1313
rect 4636 1267 4643 1353
rect 4736 1343 4743 1533
rect 4776 1407 4783 1556
rect 4736 1336 4763 1343
rect 4716 1327 4723 1333
rect 4653 1293 4667 1307
rect 4673 1313 4687 1327
rect 4693 1293 4707 1307
rect 4713 1313 4727 1327
rect 4656 1287 4663 1293
rect 4576 1127 4583 1153
rect 4576 867 4583 1073
rect 4596 1044 4604 1156
rect 4616 927 4623 1133
rect 4656 1027 4663 1193
rect 4676 947 4683 1033
rect 4656 887 4663 933
rect 4676 867 4683 893
rect 4633 863 4647 867
rect 4533 813 4547 827
rect 4616 856 4647 863
rect 4573 823 4587 827
rect 4573 816 4593 823
rect 4573 813 4587 816
rect 4536 807 4543 813
rect 4616 807 4623 856
rect 4633 853 4647 856
rect 4673 853 4687 867
rect 4656 787 4663 813
rect 4536 647 4543 773
rect 4576 647 4583 693
rect 4616 647 4623 653
rect 4573 633 4587 647
rect 4613 633 4627 647
rect 4496 527 4503 553
rect 4413 333 4427 347
rect 4453 343 4467 347
rect 4476 343 4483 473
rect 4516 467 4523 553
rect 4496 347 4503 433
rect 4556 367 4563 453
rect 4453 336 4483 343
rect 4453 333 4467 336
rect 4433 313 4447 327
rect 4416 167 4423 293
rect 4413 153 4427 167
rect 4436 127 4443 313
rect 4456 167 4463 193
rect 4453 153 4467 167
rect 4496 84 4504 196
rect 4516 107 4523 353
rect 4533 333 4547 347
rect 4553 353 4567 367
rect 4593 333 4607 347
rect 4536 287 4543 333
rect 4556 167 4563 313
rect 4576 307 4583 333
rect 4596 227 4603 333
rect 4633 333 4647 347
rect 4636 267 4643 333
rect 4656 267 4663 753
rect 4696 667 4703 1293
rect 4716 867 4723 1273
rect 4736 1203 4743 1293
rect 4756 1287 4763 1336
rect 4773 1293 4787 1307
rect 4776 1287 4783 1293
rect 4796 1283 4803 1533
rect 4816 1347 4823 1433
rect 4856 1387 4863 1653
rect 4916 1647 4923 1753
rect 4936 1744 4944 1856
rect 5016 1827 5023 2013
rect 5096 2007 5103 2073
rect 4993 1803 5007 1807
rect 5016 1803 5023 1813
rect 5036 1807 5043 1913
rect 4993 1796 5023 1803
rect 4993 1793 5007 1796
rect 4976 1747 4983 1793
rect 5033 1793 5047 1807
rect 5013 1753 5027 1767
rect 4873 1573 4887 1587
rect 4933 1573 4947 1587
rect 4996 1567 5003 1753
rect 5016 1667 5023 1753
rect 4916 1347 4923 1553
rect 5016 1547 5023 1573
rect 5037 1556 5045 1636
rect 5056 1607 5063 1633
rect 5037 1518 5045 1542
rect 5016 1483 5023 1493
rect 5016 1476 5053 1483
rect 4936 1387 4943 1413
rect 4956 1387 4963 1393
rect 5076 1387 5083 1913
rect 5116 1847 5123 2033
rect 5136 1827 5143 2053
rect 5156 1827 5163 1973
rect 5216 1967 5223 2133
rect 5233 2053 5247 2067
rect 5236 1847 5243 2053
rect 5256 2007 5263 2113
rect 5093 1773 5107 1787
rect 5133 1783 5147 1787
rect 5156 1783 5163 1813
rect 5096 1767 5103 1773
rect 5133 1776 5163 1783
rect 5133 1773 5147 1776
rect 5173 1773 5187 1787
rect 5233 1793 5247 1807
rect 5236 1787 5243 1793
rect 5213 1773 5227 1787
rect 5176 1767 5183 1773
rect 5196 1743 5203 1753
rect 5176 1736 5203 1743
rect 5096 1667 5103 1733
rect 5116 1587 5123 1733
rect 5176 1687 5183 1736
rect 4956 1363 4963 1373
rect 5116 1367 5123 1573
rect 5156 1467 5163 1593
rect 5176 1524 5184 1636
rect 5196 1483 5203 1713
rect 5216 1687 5223 1773
rect 5236 1663 5243 1753
rect 5256 1747 5263 1993
rect 5276 1987 5283 2213
rect 5296 2107 5303 2193
rect 5316 2167 5323 2353
rect 5336 2187 5343 2533
rect 5376 2447 5383 2533
rect 5376 2287 5383 2313
rect 5353 2253 5367 2267
rect 5373 2273 5387 2287
rect 5356 2187 5363 2253
rect 5336 2087 5343 2133
rect 5376 2087 5383 2133
rect 5396 2107 5403 2393
rect 5416 2347 5423 2633
rect 5436 2367 5443 2673
rect 5476 2587 5483 2653
rect 5516 2647 5523 2833
rect 5536 2767 5543 2793
rect 5556 2787 5563 2996
rect 5636 2947 5643 2953
rect 5533 2753 5547 2767
rect 5576 2687 5583 2793
rect 5576 2607 5583 2613
rect 5473 2573 5487 2587
rect 5453 2553 5467 2567
rect 5416 2307 5423 2333
rect 5436 2287 5443 2333
rect 5456 2287 5463 2293
rect 5453 2273 5467 2287
rect 5473 2253 5487 2267
rect 5416 2207 5423 2253
rect 5436 2187 5443 2213
rect 5476 2207 5483 2253
rect 5496 2203 5503 2513
rect 5533 2253 5547 2267
rect 5536 2227 5543 2253
rect 5496 2196 5523 2203
rect 5516 2167 5523 2196
rect 5556 2123 5563 2573
rect 5576 2287 5583 2593
rect 5596 2527 5603 2933
rect 5616 2704 5624 2816
rect 5636 2523 5643 2753
rect 5653 2733 5667 2747
rect 5656 2707 5663 2733
rect 5676 2707 5683 3293
rect 5715 3278 5723 3302
rect 5736 3267 5743 3533
rect 5756 3527 5763 3533
rect 5796 3527 5803 3573
rect 5753 3513 5767 3527
rect 5773 3493 5787 3507
rect 5793 3513 5807 3527
rect 5813 3503 5827 3507
rect 5813 3496 5833 3503
rect 5813 3493 5827 3496
rect 5776 3487 5783 3493
rect 5696 3043 5703 3253
rect 5715 3184 5723 3264
rect 5756 3247 5763 3433
rect 5836 3307 5843 3493
rect 5856 3387 5863 3553
rect 5896 3487 5903 3493
rect 5916 3483 5923 3693
rect 5956 3687 5963 3756
rect 6016 3727 6023 3976
rect 6036 3867 6043 3993
rect 6057 3956 6065 4036
rect 6057 3918 6065 3942
rect 6076 3847 6083 4173
rect 6096 4127 6103 4313
rect 6113 4173 6127 4187
rect 6113 4003 6127 4007
rect 6096 3996 6127 4003
rect 6076 3787 6083 3833
rect 6096 3767 6103 3996
rect 6113 3993 6127 3996
rect 6136 3907 6143 4213
rect 6176 4147 6183 4233
rect 6236 4227 6243 4373
rect 6213 4193 6227 4207
rect 6233 4213 6247 4227
rect 6216 4147 6223 4193
rect 6156 4007 6163 4013
rect 6176 4007 6183 4113
rect 6153 3993 6167 4007
rect 6196 3924 6204 4036
rect 5993 3723 6007 3727
rect 5976 3716 6007 3723
rect 5936 3547 5943 3673
rect 5976 3567 5983 3716
rect 5993 3713 6007 3716
rect 6033 3693 6047 3707
rect 6013 3673 6027 3687
rect 6016 3667 6023 3673
rect 6036 3647 6043 3693
rect 6073 3693 6087 3707
rect 6076 3687 6083 3693
rect 5936 3527 5943 3533
rect 5933 3513 5947 3527
rect 5993 3493 6007 3507
rect 6056 3507 6063 3533
rect 5916 3476 5943 3483
rect 5836 3287 5843 3293
rect 5793 3233 5807 3247
rect 5733 3223 5747 3227
rect 5733 3216 5763 3223
rect 5733 3213 5747 3216
rect 5696 3036 5723 3043
rect 5716 3027 5723 3036
rect 5693 2993 5707 3007
rect 5713 3013 5727 3027
rect 5736 3007 5743 3113
rect 5756 3067 5763 3216
rect 5776 3147 5783 3233
rect 5796 3167 5803 3233
rect 5876 3243 5883 3333
rect 5893 3243 5907 3247
rect 5853 3223 5867 3227
rect 5876 3236 5907 3243
rect 5876 3223 5883 3236
rect 5853 3216 5883 3223
rect 5893 3233 5907 3236
rect 5853 3213 5867 3216
rect 5756 3027 5763 3053
rect 5836 3047 5843 3173
rect 5876 3107 5883 3216
rect 5913 3193 5927 3207
rect 5916 3167 5923 3193
rect 5936 3127 5943 3476
rect 5976 3367 5983 3473
rect 5996 3367 6003 3493
rect 6053 3493 6067 3507
rect 6073 3473 6087 3487
rect 6036 3427 6043 3473
rect 6076 3367 6083 3473
rect 5976 3247 5983 3353
rect 6016 3247 6023 3353
rect 6096 3287 6103 3713
rect 6056 3247 6063 3273
rect 5953 3213 5967 3227
rect 5973 3233 5987 3247
rect 6013 3233 6027 3247
rect 5956 3147 5963 3213
rect 6053 3233 6067 3247
rect 6116 3227 6123 3773
rect 6156 3727 6163 3893
rect 6216 3727 6223 3993
rect 6256 3787 6263 4313
rect 6296 4227 6303 4413
rect 6316 4407 6323 4433
rect 6496 4427 6503 4433
rect 6316 4227 6323 4333
rect 6416 4227 6423 4333
rect 6436 4287 6443 4393
rect 6516 4327 6523 4433
rect 6556 4387 6563 4453
rect 6313 4213 6327 4227
rect 6276 4163 6283 4173
rect 6336 4167 6343 4213
rect 6413 4213 6427 4227
rect 6436 4207 6443 4253
rect 6456 4227 6463 4293
rect 6353 4173 6367 4187
rect 6356 4167 6363 4173
rect 6276 4156 6303 4163
rect 6296 4083 6303 4156
rect 6436 4163 6443 4173
rect 6453 4163 6467 4167
rect 6436 4156 6467 4163
rect 6453 4153 6467 4156
rect 6296 4076 6323 4083
rect 6297 3956 6305 4036
rect 6297 3918 6305 3942
rect 6316 3747 6323 4076
rect 6353 4003 6367 4007
rect 6393 4003 6407 4007
rect 6353 3996 6383 4003
rect 6353 3993 6367 3996
rect 6337 3758 6345 3782
rect 6376 3767 6383 3996
rect 6393 3996 6423 4003
rect 6393 3993 6407 3996
rect 6416 3967 6423 3996
rect 6436 3924 6444 4036
rect 6496 3807 6503 4273
rect 6516 4187 6523 4213
rect 6556 4207 6563 4233
rect 6576 4207 6583 4413
rect 6676 4267 6683 4693
rect 6696 4247 6703 5113
rect 6596 4207 6603 4213
rect 6633 4213 6647 4227
rect 6673 4223 6687 4227
rect 6533 4173 6547 4187
rect 6536 4087 6543 4173
rect 6636 4183 6643 4213
rect 6653 4193 6667 4207
rect 6673 4216 6703 4223
rect 6673 4213 6687 4216
rect 6656 4187 6663 4193
rect 6616 4176 6643 4183
rect 6616 4167 6623 4176
rect 6513 3993 6527 4007
rect 6537 3956 6545 4036
rect 6636 4007 6643 4153
rect 6593 4003 6607 4007
rect 6576 3996 6607 4003
rect 6537 3918 6545 3942
rect 6576 3927 6583 3996
rect 6593 3993 6607 3996
rect 6633 3993 6647 4007
rect 6276 3727 6283 3733
rect 6133 3693 6147 3707
rect 6136 3647 6143 3693
rect 6153 3673 6167 3687
rect 6136 3543 6143 3633
rect 6156 3627 6163 3673
rect 6176 3667 6183 3693
rect 6253 3693 6267 3707
rect 6153 3543 6167 3547
rect 6136 3536 6167 3543
rect 6153 3533 6167 3536
rect 6176 3523 6183 3653
rect 6196 3547 6203 3673
rect 6236 3647 6243 3673
rect 6193 3523 6207 3527
rect 6176 3516 6207 3523
rect 6133 3493 6147 3507
rect 6193 3513 6207 3516
rect 6216 3503 6223 3633
rect 6256 3607 6263 3693
rect 6256 3527 6263 3533
rect 6233 3503 6247 3507
rect 6216 3496 6247 3503
rect 6253 3513 6267 3527
rect 6233 3493 6247 3496
rect 6136 3427 6143 3493
rect 6136 3287 6143 3293
rect 6156 3267 6163 3293
rect 6196 3267 6203 3353
rect 6153 3263 6167 3267
rect 6136 3256 6167 3263
rect 6073 3213 6087 3227
rect 6136 3223 6143 3256
rect 6153 3253 6167 3256
rect 6173 3233 6187 3247
rect 6193 3253 6207 3267
rect 6136 3216 6163 3223
rect 5993 3193 6007 3207
rect 5996 3147 6003 3193
rect 6076 3127 6083 3213
rect 5856 3067 5863 3093
rect 5876 3076 6003 3083
rect 5876 3047 5883 3076
rect 5893 3063 5907 3067
rect 5893 3056 5943 3063
rect 5893 3053 5907 3056
rect 5793 3033 5807 3047
rect 5753 3013 5767 3027
rect 5813 3013 5827 3027
rect 5833 3033 5847 3047
rect 5853 3013 5867 3027
rect 5873 3033 5887 3047
rect 5936 3047 5943 3056
rect 5976 3047 5983 3053
rect 5953 3013 5967 3027
rect 5973 3033 5987 3047
rect 5996 3027 6003 3076
rect 6116 3067 6123 3193
rect 6136 3187 6143 3193
rect 6136 3067 6143 3173
rect 6156 3147 6163 3216
rect 6176 3087 6183 3233
rect 6216 3107 6223 3313
rect 6236 3267 6243 3373
rect 6256 3307 6263 3433
rect 6256 3267 6263 3273
rect 6256 3247 6263 3253
rect 6276 3247 6283 3713
rect 6296 3543 6303 3733
rect 6337 3664 6345 3744
rect 6376 3703 6383 3753
rect 6393 3703 6407 3707
rect 6376 3696 6407 3703
rect 6393 3693 6407 3696
rect 6356 3667 6363 3693
rect 6416 3647 6423 3773
rect 6456 3607 6463 3793
rect 6656 3787 6663 4133
rect 6696 4047 6703 4216
rect 6676 3924 6684 4036
rect 6476 3664 6484 3776
rect 6296 3536 6323 3543
rect 6293 3493 6307 3507
rect 6296 3447 6303 3493
rect 6296 3287 6303 3413
rect 6296 3247 6303 3273
rect 6253 3233 6267 3247
rect 6293 3233 6307 3247
rect 6236 3203 6243 3213
rect 6236 3196 6263 3203
rect 6256 3167 6263 3196
rect 6133 3053 6147 3067
rect 6013 3013 6027 3027
rect 6093 3033 6107 3047
rect 5733 2993 5747 3007
rect 5696 2947 5703 2993
rect 5716 2887 5723 2933
rect 5755 2798 5763 2822
rect 5693 2733 5707 2747
rect 5696 2683 5703 2733
rect 5716 2683 5723 2773
rect 5755 2704 5763 2784
rect 5796 2687 5803 2993
rect 5816 2807 5823 3013
rect 5856 2987 5863 3013
rect 5833 2733 5847 2747
rect 5836 2727 5843 2733
rect 5856 2687 5863 2813
rect 5876 2767 5883 2793
rect 5873 2753 5887 2767
rect 5893 2733 5907 2747
rect 5896 2723 5903 2733
rect 5876 2716 5903 2723
rect 5696 2676 5723 2683
rect 5656 2547 5663 2673
rect 5716 2547 5723 2676
rect 5876 2667 5883 2716
rect 5916 2707 5923 2953
rect 5956 2847 5963 3013
rect 5936 2767 5943 2833
rect 5933 2753 5947 2767
rect 5953 2733 5967 2747
rect 5956 2727 5963 2733
rect 5976 2727 5983 2853
rect 6016 2807 6023 3013
rect 6176 3007 6183 3053
rect 6196 3047 6203 3093
rect 6193 3033 6207 3047
rect 6236 3047 6243 3073
rect 6256 3067 6263 3073
rect 6253 3053 6267 3067
rect 6233 3033 6247 3047
rect 6056 2767 6063 2833
rect 6053 2763 6067 2767
rect 6036 2756 6067 2763
rect 5756 2587 5763 2633
rect 5753 2573 5767 2587
rect 5736 2567 5743 2573
rect 5733 2553 5747 2567
rect 5776 2567 5783 2613
rect 5816 2587 5823 2633
rect 5836 2567 5843 2633
rect 5793 2553 5807 2567
rect 5813 2533 5827 2547
rect 5833 2553 5847 2567
rect 5853 2543 5867 2547
rect 5853 2536 5883 2543
rect 5853 2533 5867 2536
rect 5636 2516 5663 2523
rect 5616 2307 5623 2373
rect 5636 2287 5643 2373
rect 5656 2347 5663 2516
rect 5676 2427 5683 2533
rect 5836 2487 5843 2513
rect 5573 2273 5587 2287
rect 5633 2273 5647 2287
rect 5536 2116 5563 2123
rect 5436 2087 5443 2113
rect 5536 2087 5543 2116
rect 5576 2107 5583 2233
rect 5656 2127 5663 2233
rect 5676 2207 5683 2413
rect 5716 2307 5723 2393
rect 5736 2327 5743 2433
rect 5776 2367 5783 2453
rect 5876 2447 5883 2536
rect 5796 2347 5803 2413
rect 5816 2307 5823 2353
rect 5836 2327 5843 2373
rect 5713 2293 5727 2307
rect 5753 2293 5767 2307
rect 5756 2287 5763 2293
rect 5813 2293 5827 2307
rect 5733 2273 5747 2287
rect 5773 2273 5787 2287
rect 5736 2267 5743 2273
rect 5716 2107 5723 2253
rect 5776 2247 5783 2273
rect 5856 2227 5863 2293
rect 5756 2187 5763 2213
rect 5876 2207 5883 2233
rect 5896 2227 5903 2693
rect 5916 2627 5923 2693
rect 5956 2567 5963 2613
rect 5976 2587 5983 2633
rect 5996 2587 6003 2613
rect 5933 2533 5947 2547
rect 5953 2553 5967 2567
rect 5973 2533 5987 2547
rect 5916 2307 5923 2493
rect 5936 2487 5943 2533
rect 5936 2287 5943 2313
rect 5916 2223 5923 2233
rect 5916 2216 5943 2223
rect 5756 2107 5763 2173
rect 5753 2093 5767 2107
rect 5293 2073 5307 2087
rect 5313 2053 5327 2067
rect 5333 2073 5347 2087
rect 5373 2073 5387 2087
rect 5413 2053 5427 2067
rect 5433 2073 5447 2087
rect 5473 2073 5487 2087
rect 5533 2083 5547 2087
rect 5516 2076 5547 2083
rect 5356 2003 5363 2053
rect 5336 1996 5363 2003
rect 5336 1947 5343 1996
rect 5333 1823 5347 1827
rect 5333 1816 5363 1823
rect 5333 1813 5347 1816
rect 5356 1787 5363 1816
rect 5373 1773 5387 1787
rect 5216 1656 5243 1663
rect 5216 1607 5223 1656
rect 5256 1647 5263 1673
rect 5236 1507 5243 1613
rect 5256 1527 5263 1593
rect 5277 1556 5285 1636
rect 5277 1518 5285 1542
rect 5176 1476 5203 1483
rect 4936 1356 4963 1363
rect 4936 1347 4943 1356
rect 4853 1343 4867 1347
rect 4836 1336 4867 1343
rect 4813 1293 4827 1307
rect 4796 1276 4823 1283
rect 4816 1247 4823 1276
rect 4736 1196 4763 1203
rect 4756 1187 4763 1196
rect 4735 1076 4743 1156
rect 4776 1147 4783 1213
rect 4796 1187 4803 1233
rect 4836 1227 4843 1336
rect 4853 1333 4867 1336
rect 4873 1313 4887 1327
rect 4893 1333 4907 1347
rect 4933 1333 4947 1347
rect 4876 1283 4883 1313
rect 4876 1276 4893 1283
rect 4836 1127 4843 1153
rect 4876 1127 4883 1133
rect 4753 1123 4767 1127
rect 4753 1116 4783 1123
rect 4753 1113 4767 1116
rect 4735 1038 4743 1062
rect 4756 1047 4763 1093
rect 4776 1023 4783 1116
rect 4813 1093 4827 1107
rect 4833 1113 4847 1127
rect 4873 1113 4887 1127
rect 4816 1087 4823 1093
rect 4756 1016 4783 1023
rect 4716 827 4723 853
rect 4736 847 4743 893
rect 4756 887 4763 1016
rect 4796 907 4803 1073
rect 4816 947 4823 1073
rect 4896 1027 4903 1233
rect 4916 1227 4923 1333
rect 4973 1333 4987 1347
rect 4936 1247 4943 1293
rect 4756 847 4763 873
rect 4796 847 4803 893
rect 4733 833 4747 847
rect 4716 807 4723 813
rect 4793 833 4807 847
rect 4813 823 4827 827
rect 4813 816 4833 823
rect 4813 813 4827 816
rect 4716 707 4723 733
rect 4716 667 4723 693
rect 4736 667 4743 793
rect 4856 707 4863 993
rect 4876 887 4883 1013
rect 4916 1007 4923 1173
rect 4956 1163 4963 1293
rect 4936 1156 4963 1163
rect 4936 1127 4943 1156
rect 4933 1113 4947 1127
rect 4976 1127 4983 1213
rect 4996 1187 5003 1353
rect 5176 1347 5183 1476
rect 5013 1293 5027 1307
rect 5053 1293 5067 1307
rect 5036 1247 5043 1273
rect 5056 1167 5063 1293
rect 4973 1113 4987 1127
rect 4913 863 4927 867
rect 4913 856 4943 863
rect 4913 853 4927 856
rect 4936 803 4943 856
rect 4956 847 4963 1033
rect 4996 967 5003 1133
rect 5016 1107 5023 1153
rect 5096 1147 5103 1253
rect 5116 1227 5123 1333
rect 5156 1327 5163 1333
rect 5196 1327 5203 1453
rect 5236 1347 5243 1493
rect 5256 1367 5263 1493
rect 5316 1447 5323 1673
rect 5356 1623 5363 1693
rect 5376 1687 5383 1773
rect 5356 1616 5383 1623
rect 5376 1607 5383 1616
rect 5373 1593 5387 1607
rect 5356 1503 5363 1573
rect 5356 1496 5383 1503
rect 5376 1487 5383 1496
rect 5133 1293 5147 1307
rect 5153 1313 5167 1327
rect 5173 1293 5187 1307
rect 5213 1293 5227 1307
rect 5276 1307 5283 1413
rect 5316 1347 5323 1393
rect 5356 1367 5363 1473
rect 5313 1343 5327 1347
rect 5296 1336 5327 1343
rect 5353 1343 5367 1347
rect 5376 1343 5383 1413
rect 5396 1407 5403 2013
rect 5416 1987 5423 2053
rect 5496 2043 5503 2073
rect 5476 2036 5503 2043
rect 5456 1867 5463 2013
rect 5436 1747 5443 1833
rect 5476 1827 5483 2036
rect 5516 2023 5523 2076
rect 5533 2073 5547 2076
rect 5596 2067 5603 2093
rect 5653 2073 5667 2087
rect 5693 2083 5707 2087
rect 5693 2076 5723 2083
rect 5693 2073 5707 2076
rect 5716 2063 5723 2076
rect 5796 2067 5803 2133
rect 5856 2083 5863 2173
rect 5873 2083 5887 2087
rect 5856 2076 5887 2083
rect 5873 2073 5887 2076
rect 5733 2063 5747 2067
rect 5716 2056 5747 2063
rect 5733 2053 5747 2056
rect 5496 2016 5523 2023
rect 5496 1887 5503 2016
rect 5536 1927 5543 2033
rect 5556 2007 5563 2053
rect 5576 1983 5583 2033
rect 5556 1976 5583 1983
rect 5556 1887 5563 1976
rect 5473 1803 5487 1807
rect 5456 1796 5487 1803
rect 5416 1524 5424 1636
rect 5436 1487 5443 1633
rect 5456 1587 5463 1796
rect 5473 1793 5487 1796
rect 5476 1643 5483 1693
rect 5516 1663 5523 1833
rect 5536 1827 5543 1853
rect 5533 1773 5547 1787
rect 5536 1687 5543 1773
rect 5576 1727 5583 1873
rect 5596 1867 5603 2033
rect 5676 1923 5683 2053
rect 5727 2036 5743 2043
rect 5656 1916 5683 1923
rect 5656 1907 5663 1916
rect 5656 1827 5663 1893
rect 5676 1827 5683 1893
rect 5696 1847 5703 2013
rect 5736 1827 5743 2036
rect 5756 1987 5763 2053
rect 5773 2033 5787 2047
rect 5813 2033 5827 2047
rect 5776 2007 5783 2033
rect 5776 1827 5783 1993
rect 5613 1773 5627 1787
rect 5633 1793 5647 1807
rect 5693 1793 5707 1807
rect 5816 1823 5823 1973
rect 5856 1907 5863 2053
rect 5876 1927 5883 2053
rect 5897 2036 5905 2116
rect 5897 1998 5905 2022
rect 5896 1867 5903 1953
rect 5916 1927 5923 2193
rect 5936 2183 5943 2216
rect 5956 2207 5963 2493
rect 5976 2447 5983 2533
rect 6016 2447 6023 2713
rect 6036 2607 6043 2756
rect 6053 2753 6067 2756
rect 6096 2747 6103 2793
rect 6056 2667 6063 2713
rect 6056 2587 6063 2653
rect 6076 2507 6083 2673
rect 6096 2627 6103 2713
rect 6156 2703 6163 2813
rect 6216 2787 6223 2993
rect 6296 2987 6303 3153
rect 6213 2773 6227 2787
rect 6276 2783 6283 2833
rect 6296 2807 6303 2973
rect 6276 2776 6303 2783
rect 6176 2747 6183 2773
rect 6296 2767 6303 2776
rect 6193 2733 6207 2747
rect 6253 2733 6267 2747
rect 6293 2753 6307 2767
rect 6136 2696 6163 2703
rect 6117 2516 6125 2596
rect 6117 2478 6125 2502
rect 6116 2287 6123 2433
rect 5993 2273 6007 2287
rect 6013 2253 6027 2267
rect 6053 2253 6067 2267
rect 5936 2176 5963 2183
rect 5936 2087 5943 2153
rect 5956 2127 5963 2176
rect 5956 2087 5963 2113
rect 5953 2073 5967 2087
rect 5816 1816 5843 1823
rect 5836 1807 5843 1816
rect 5653 1773 5667 1787
rect 5596 1747 5603 1773
rect 5616 1767 5623 1773
rect 5636 1687 5643 1753
rect 5656 1687 5663 1773
rect 5696 1747 5703 1793
rect 5516 1656 5543 1663
rect 5476 1636 5523 1643
rect 5476 1607 5483 1613
rect 5516 1607 5523 1636
rect 5536 1627 5543 1656
rect 5616 1607 5623 1633
rect 5473 1593 5487 1607
rect 5513 1593 5527 1607
rect 5533 1573 5547 1587
rect 5613 1593 5627 1607
rect 5536 1527 5543 1573
rect 5556 1543 5563 1553
rect 5556 1536 5583 1543
rect 5507 1516 5523 1523
rect 5416 1343 5423 1473
rect 5136 1287 5143 1293
rect 5147 1276 5163 1283
rect 5116 1167 5123 1213
rect 5156 1187 5163 1276
rect 5176 1227 5183 1293
rect 5216 1267 5223 1293
rect 5256 1247 5263 1293
rect 5276 1183 5283 1293
rect 5296 1187 5303 1336
rect 5313 1333 5327 1336
rect 5353 1336 5383 1343
rect 5396 1336 5423 1343
rect 5353 1333 5367 1336
rect 5396 1327 5403 1336
rect 5436 1327 5443 1393
rect 5336 1303 5343 1313
rect 5316 1296 5343 1303
rect 5316 1207 5323 1296
rect 5393 1313 5407 1327
rect 5413 1293 5427 1307
rect 5256 1176 5283 1183
rect 5116 1127 5123 1153
rect 5073 1123 5087 1127
rect 5053 1093 5067 1107
rect 5073 1116 5103 1123
rect 5073 1113 5087 1116
rect 5096 1083 5103 1116
rect 5113 1113 5127 1127
rect 5156 1127 5163 1173
rect 5176 1127 5183 1153
rect 5193 1133 5207 1147
rect 5153 1113 5167 1127
rect 5173 1113 5187 1127
rect 5213 1113 5227 1127
rect 5096 1076 5123 1083
rect 5116 1067 5123 1076
rect 4953 833 4967 847
rect 4936 796 4963 803
rect 4713 653 4727 667
rect 4693 613 4707 627
rect 4696 607 4703 613
rect 4756 607 4763 653
rect 4836 647 4843 653
rect 4776 627 4783 633
rect 4773 613 4787 627
rect 4833 633 4847 647
rect 4876 627 4883 653
rect 4873 613 4887 627
rect 4916 583 4923 653
rect 4767 576 4923 583
rect 4936 527 4943 773
rect 4956 767 4963 796
rect 4756 387 4763 493
rect 4756 367 4763 373
rect 4693 333 4707 347
rect 4733 333 4747 347
rect 4753 353 4767 367
rect 4813 363 4827 367
rect 4773 343 4787 347
rect 4796 356 4827 363
rect 4796 343 4803 356
rect 4773 336 4803 343
rect 4813 353 4827 356
rect 4773 333 4787 336
rect 4696 287 4703 333
rect 4736 323 4743 333
rect 4736 316 4773 323
rect 4833 313 4847 327
rect 4836 267 4843 313
rect 4876 287 4883 513
rect 4896 304 4904 416
rect 4976 407 4983 533
rect 4956 343 4963 393
rect 4973 343 4987 347
rect 4956 336 4987 343
rect 4956 283 4963 336
rect 4973 333 4987 336
rect 4936 276 4963 283
rect 4616 187 4623 193
rect 4553 153 4567 167
rect 4573 133 4587 147
rect 4616 147 4623 173
rect 4613 133 4627 147
rect 4576 107 4583 133
rect 4576 67 4583 93
rect 4636 67 4643 253
rect 4696 167 4703 173
rect 4673 133 4687 147
rect 4693 153 4707 167
rect 4676 127 4683 133
rect 4753 113 4767 127
rect 4793 123 4807 127
rect 4816 123 4823 233
rect 4853 153 4867 167
rect 4793 116 4823 123
rect 4793 113 4807 116
rect 4756 87 4763 113
rect 4856 87 4863 153
rect 4877 116 4885 196
rect 4936 167 4943 276
rect 4976 267 4983 313
rect 4996 307 5003 933
rect 5016 847 5023 1013
rect 5096 907 5103 1053
rect 5116 947 5123 1053
rect 5176 847 5183 913
rect 5013 833 5027 847
rect 5033 813 5047 827
rect 5093 813 5107 827
rect 5173 833 5187 847
rect 5036 787 5043 813
rect 5096 767 5103 813
rect 5156 727 5163 733
rect 5033 613 5047 627
rect 5016 267 5023 593
rect 5036 527 5043 613
rect 5056 607 5063 633
rect 5156 627 5163 713
rect 5153 613 5167 627
rect 5133 593 5147 607
rect 5173 593 5187 607
rect 5096 527 5103 593
rect 5176 583 5183 593
rect 5156 576 5183 583
rect 5035 398 5043 422
rect 5035 304 5043 384
rect 5056 367 5063 433
rect 5136 427 5143 533
rect 5156 467 5163 576
rect 5196 427 5203 853
rect 5216 847 5223 973
rect 5236 947 5243 1173
rect 5256 1127 5263 1176
rect 5253 1113 5267 1127
rect 5293 1113 5307 1127
rect 5336 1123 5343 1253
rect 5356 1187 5363 1293
rect 5353 1123 5367 1127
rect 5336 1116 5367 1123
rect 5256 947 5263 1073
rect 5276 847 5283 1093
rect 5213 833 5227 847
rect 5233 633 5247 647
rect 5236 527 5243 633
rect 5257 596 5265 676
rect 5257 558 5265 582
rect 5276 547 5283 833
rect 5296 827 5303 1073
rect 5336 927 5343 1116
rect 5353 1113 5367 1116
rect 5316 647 5323 873
rect 5313 633 5327 647
rect 5296 603 5303 633
rect 5336 627 5343 913
rect 5356 887 5363 1013
rect 5376 987 5383 1213
rect 5396 1127 5403 1233
rect 5416 1207 5423 1293
rect 5456 1267 5463 1273
rect 5476 1227 5483 1453
rect 5496 1427 5503 1453
rect 5516 1427 5523 1516
rect 5496 1347 5503 1353
rect 5527 1336 5543 1343
rect 5536 1327 5543 1336
rect 5556 1327 5563 1493
rect 5576 1387 5583 1536
rect 5596 1327 5603 1453
rect 5616 1347 5623 1513
rect 5636 1507 5643 1673
rect 5656 1627 5663 1653
rect 5676 1627 5683 1713
rect 5653 1573 5667 1587
rect 5696 1563 5703 1673
rect 5716 1607 5723 1733
rect 5736 1607 5743 1793
rect 5773 1773 5787 1787
rect 5793 1793 5807 1807
rect 5813 1773 5827 1787
rect 5833 1793 5847 1807
rect 5853 1773 5867 1787
rect 5873 1773 5887 1787
rect 5776 1767 5783 1773
rect 5756 1607 5763 1673
rect 5816 1667 5823 1773
rect 5856 1763 5863 1773
rect 5836 1756 5863 1763
rect 5836 1707 5843 1756
rect 5796 1607 5803 1633
rect 5856 1627 5863 1733
rect 5896 1707 5903 1793
rect 5936 1787 5943 2033
rect 5913 1773 5927 1787
rect 5916 1667 5923 1773
rect 5956 1767 5963 1853
rect 5976 1847 5983 2233
rect 6016 2227 6023 2253
rect 6036 2183 6043 2233
rect 6056 2227 6063 2253
rect 6036 2176 6063 2183
rect 5993 2073 6007 2087
rect 6016 2067 6023 2093
rect 6036 2004 6044 2116
rect 6056 2087 6063 2176
rect 6076 1963 6083 2273
rect 6113 2273 6127 2287
rect 6136 2243 6143 2696
rect 6156 2347 6163 2633
rect 6176 2567 6183 2733
rect 6196 2647 6203 2733
rect 6256 2727 6263 2733
rect 6173 2553 6187 2567
rect 6116 2236 6143 2243
rect 6096 2167 6103 2233
rect 6096 2027 6103 2073
rect 6116 2007 6123 2236
rect 6196 2227 6203 2533
rect 6256 2484 6264 2596
rect 6296 2447 6303 2693
rect 6296 2287 6303 2353
rect 6316 2327 6323 3536
rect 6336 3327 6343 3593
rect 6393 3543 6407 3547
rect 6393 3536 6423 3543
rect 6393 3533 6407 3536
rect 6416 3523 6423 3536
rect 6433 3523 6447 3527
rect 6416 3516 6447 3523
rect 6433 3513 6447 3516
rect 6373 3493 6387 3507
rect 6376 3367 6383 3493
rect 6457 3476 6465 3556
rect 6457 3438 6465 3462
rect 6336 3267 6343 3273
rect 6333 3253 6347 3267
rect 6353 3233 6367 3247
rect 6356 3207 6363 3233
rect 6453 3233 6467 3247
rect 6356 3187 6363 3193
rect 6376 3187 6383 3213
rect 6456 3207 6463 3233
rect 6356 3067 6363 3173
rect 6336 2827 6343 2993
rect 6336 2767 6343 2813
rect 6333 2753 6347 2767
rect 6353 2743 6367 2747
rect 6376 2743 6383 2933
rect 6396 2787 6403 2793
rect 6393 2773 6407 2787
rect 6353 2736 6383 2743
rect 6353 2733 6367 2736
rect 6413 2733 6427 2747
rect 6356 2727 6363 2733
rect 6336 2567 6343 2613
rect 6376 2567 6383 2613
rect 6416 2587 6423 2733
rect 6436 2583 6443 3153
rect 6456 3063 6463 3133
rect 6476 3087 6483 3233
rect 6496 3127 6503 3773
rect 6516 3527 6523 3753
rect 6533 3693 6547 3707
rect 6593 3713 6607 3727
rect 6673 3743 6687 3747
rect 6653 3713 6667 3727
rect 6673 3736 6703 3743
rect 6673 3733 6687 3736
rect 6536 3627 6543 3693
rect 6596 3607 6603 3713
rect 6513 3513 6527 3527
rect 6553 3523 6567 3527
rect 6536 3516 6567 3523
rect 6536 3467 6543 3516
rect 6553 3513 6567 3516
rect 6537 3278 6545 3302
rect 6516 3227 6523 3253
rect 6537 3184 6545 3264
rect 6556 3247 6563 3273
rect 6556 3187 6563 3213
rect 6576 3167 6583 3593
rect 6596 3444 6604 3556
rect 6596 3267 6603 3393
rect 6593 3213 6607 3227
rect 6616 3223 6623 3273
rect 6636 3267 6643 3633
rect 6633 3223 6647 3227
rect 6616 3216 6647 3223
rect 6633 3213 6647 3216
rect 6496 3067 6503 3093
rect 6473 3063 6487 3067
rect 6456 3056 6487 3063
rect 6473 3053 6487 3056
rect 6496 2863 6503 3013
rect 6496 2856 6523 2863
rect 6497 2798 6505 2822
rect 6473 2743 6487 2747
rect 6456 2736 6487 2743
rect 6456 2707 6463 2736
rect 6473 2733 6487 2736
rect 6497 2704 6505 2784
rect 6516 2727 6523 2856
rect 6436 2576 6463 2583
rect 6333 2553 6347 2567
rect 6353 2533 6367 2547
rect 6373 2553 6387 2567
rect 6393 2533 6407 2547
rect 6396 2407 6403 2533
rect 6316 2287 6323 2313
rect 6336 2287 6343 2353
rect 6376 2307 6383 2333
rect 6396 2287 6403 2353
rect 6416 2307 6423 2453
rect 6436 2427 6443 2533
rect 6436 2347 6443 2393
rect 6456 2347 6463 2576
rect 6476 2347 6483 2533
rect 6496 2527 6503 2653
rect 6516 2587 6523 2693
rect 6536 2587 6543 3113
rect 6556 3047 6563 3133
rect 6596 3067 6603 3213
rect 6553 3033 6567 3047
rect 6593 3043 6607 3047
rect 6616 3043 6623 3193
rect 6636 3087 6643 3153
rect 6593 3036 6623 3043
rect 6593 3033 6607 3036
rect 6613 3023 6627 3027
rect 6613 3016 6643 3023
rect 6613 3013 6627 3016
rect 6576 2747 6583 2993
rect 6636 2987 6643 3016
rect 6593 2743 6607 2747
rect 6593 2736 6623 2743
rect 6593 2733 6607 2736
rect 6513 2573 6527 2587
rect 6576 2583 6583 2713
rect 6556 2576 6583 2583
rect 6556 2383 6563 2576
rect 6616 2567 6623 2736
rect 6636 2704 6644 2816
rect 6656 2583 6663 3713
rect 6676 3184 6684 3296
rect 6696 2667 6703 3736
rect 6656 2576 6683 2583
rect 6613 2553 6627 2567
rect 6633 2533 6647 2547
rect 6536 2376 6563 2383
rect 6476 2307 6483 2313
rect 6473 2293 6487 2307
rect 6213 2253 6227 2267
rect 6273 2253 6287 2267
rect 6293 2273 6307 2287
rect 6333 2273 6347 2287
rect 6136 2004 6144 2116
rect 6076 1956 6123 1963
rect 6076 1947 6083 1956
rect 5993 1773 6007 1787
rect 6013 1793 6027 1807
rect 6033 1773 6047 1787
rect 5853 1613 5867 1627
rect 5836 1607 5843 1613
rect 5753 1593 5767 1607
rect 5793 1603 5807 1607
rect 5773 1573 5787 1587
rect 5793 1596 5823 1603
rect 5793 1593 5807 1596
rect 5696 1556 5723 1563
rect 5533 1313 5547 1327
rect 5593 1313 5607 1327
rect 5613 1293 5627 1307
rect 5416 1127 5423 1173
rect 5393 1113 5407 1127
rect 5413 1113 5427 1127
rect 5456 1127 5463 1153
rect 5453 1113 5467 1127
rect 5416 907 5423 1073
rect 5356 847 5363 873
rect 5396 847 5403 853
rect 5436 847 5443 893
rect 5353 833 5367 847
rect 5393 833 5407 847
rect 5453 813 5467 827
rect 5356 687 5363 793
rect 5296 596 5323 603
rect 5136 367 5143 413
rect 5176 383 5183 393
rect 5196 383 5203 413
rect 5236 387 5243 453
rect 5256 387 5263 473
rect 5316 387 5323 596
rect 5396 564 5404 676
rect 5176 376 5203 383
rect 5176 367 5183 376
rect 5336 367 5343 393
rect 5356 387 5363 433
rect 5416 387 5423 733
rect 5436 587 5443 773
rect 5456 767 5463 813
rect 5476 807 5483 1173
rect 5516 1163 5523 1273
rect 5636 1227 5643 1473
rect 5656 1327 5663 1353
rect 5676 1343 5683 1433
rect 5696 1427 5703 1513
rect 5716 1387 5723 1556
rect 5736 1467 5743 1513
rect 5676 1336 5703 1343
rect 5653 1313 5667 1327
rect 5673 1293 5687 1307
rect 5496 1156 5523 1163
rect 5496 1127 5503 1156
rect 5513 1143 5527 1147
rect 5513 1136 5533 1143
rect 5513 1133 5527 1136
rect 5493 1113 5507 1127
rect 5556 1087 5563 1213
rect 5593 1133 5607 1147
rect 5573 1093 5587 1107
rect 5613 1093 5627 1107
rect 5576 1087 5583 1093
rect 5496 787 5503 1073
rect 5576 867 5583 1073
rect 5616 907 5623 1093
rect 5553 813 5567 827
rect 5613 833 5627 847
rect 5533 793 5547 807
rect 5536 647 5543 793
rect 5556 727 5563 813
rect 5616 787 5623 833
rect 5636 827 5643 1033
rect 5656 1007 5663 1253
rect 5676 1227 5683 1293
rect 5696 1247 5703 1336
rect 5716 1327 5723 1353
rect 5736 1347 5743 1393
rect 5713 1313 5727 1327
rect 5716 1163 5723 1233
rect 5696 1156 5723 1163
rect 5696 1127 5703 1156
rect 5736 1143 5743 1293
rect 5756 1267 5763 1413
rect 5776 1407 5783 1453
rect 5796 1367 5803 1553
rect 5816 1487 5823 1596
rect 5833 1593 5847 1607
rect 5876 1607 5883 1613
rect 5873 1593 5887 1607
rect 5896 1567 5903 1653
rect 5976 1627 5983 1773
rect 5996 1767 6003 1773
rect 6036 1663 6043 1693
rect 6056 1667 6063 1893
rect 6116 1867 6123 1956
rect 6156 1887 6163 2213
rect 6176 1887 6183 1973
rect 6096 1807 6103 1853
rect 6176 1807 6183 1853
rect 6196 1827 6203 2193
rect 6216 2187 6223 2253
rect 6276 2247 6283 2253
rect 6236 2167 6243 2233
rect 6216 2087 6223 2113
rect 6236 2087 6243 2133
rect 6213 2073 6227 2087
rect 6073 1773 6087 1787
rect 6093 1793 6107 1807
rect 6113 1773 6127 1787
rect 6173 1793 6187 1807
rect 6216 1787 6223 1973
rect 6256 1927 6263 2233
rect 6336 2147 6343 2233
rect 6275 2036 6283 2116
rect 6336 2103 6343 2133
rect 6356 2127 6363 2273
rect 6393 2273 6407 2287
rect 6413 2253 6427 2267
rect 6376 2247 6383 2253
rect 6416 2247 6423 2253
rect 6316 2096 6343 2103
rect 6275 1998 6283 2022
rect 6296 1963 6303 2053
rect 6276 1956 6303 1963
rect 6236 1807 6243 1913
rect 6276 1807 6283 1956
rect 6316 1847 6323 2096
rect 6356 2087 6363 2113
rect 6333 2053 6347 2067
rect 6353 2073 6367 2087
rect 6336 1967 6343 2053
rect 6336 1827 6343 1953
rect 6376 1827 6383 2173
rect 6396 2107 6403 2153
rect 6436 2127 6443 2253
rect 6456 2187 6463 2293
rect 6536 2263 6543 2376
rect 6576 2287 6583 2513
rect 6596 2307 6603 2333
rect 6596 2287 6603 2293
rect 6516 2256 6543 2263
rect 6593 2273 6607 2287
rect 6476 2207 6483 2233
rect 6496 2163 6503 2213
rect 6476 2156 6503 2163
rect 6416 2087 6423 2093
rect 6393 2053 6407 2067
rect 6413 2073 6427 2087
rect 6396 2043 6403 2053
rect 6396 2036 6423 2043
rect 6416 2007 6423 2036
rect 6436 1867 6443 2113
rect 6476 2107 6483 2156
rect 6516 2127 6523 2256
rect 6613 2263 6627 2267
rect 6636 2263 6643 2533
rect 6656 2287 6663 2433
rect 6676 2343 6683 2576
rect 6696 2567 6703 2613
rect 6676 2336 6703 2343
rect 6676 2287 6683 2313
rect 6673 2273 6687 2287
rect 6613 2256 6643 2263
rect 6613 2253 6627 2256
rect 6573 2233 6587 2247
rect 6653 2233 6667 2247
rect 6536 2107 6543 2233
rect 6576 2227 6583 2233
rect 6473 2093 6487 2107
rect 6493 2053 6507 2067
rect 6496 2047 6503 2053
rect 6496 1947 6503 2033
rect 6296 1807 6303 1813
rect 6233 1793 6247 1807
rect 6193 1773 6207 1787
rect 6293 1793 6307 1807
rect 6353 1803 6367 1807
rect 6253 1783 6267 1787
rect 6253 1776 6283 1783
rect 6253 1773 6267 1776
rect 6076 1747 6083 1773
rect 6116 1687 6123 1773
rect 6016 1656 6043 1663
rect 5976 1607 5983 1613
rect 6016 1607 6023 1656
rect 6056 1607 6063 1653
rect 6013 1593 6027 1607
rect 5913 1553 5927 1567
rect 5976 1567 5983 1593
rect 6033 1573 6047 1587
rect 6053 1593 6067 1607
rect 6076 1587 6083 1673
rect 6116 1627 6123 1653
rect 6136 1647 6143 1753
rect 6113 1613 6127 1627
rect 6133 1593 6147 1607
rect 5836 1467 5843 1553
rect 5816 1367 5823 1393
rect 5793 1343 5807 1347
rect 5776 1336 5807 1343
rect 5776 1307 5783 1336
rect 5793 1333 5807 1336
rect 5813 1313 5827 1327
rect 5776 1243 5783 1273
rect 5796 1247 5803 1293
rect 5816 1267 5823 1313
rect 5856 1303 5863 1473
rect 5896 1407 5903 1553
rect 5916 1543 5923 1553
rect 5916 1536 5943 1543
rect 5936 1523 5943 1536
rect 5936 1516 5953 1523
rect 5916 1503 5923 1513
rect 5916 1496 5943 1503
rect 5896 1347 5903 1393
rect 5916 1367 5923 1413
rect 5936 1367 5943 1496
rect 5976 1407 5983 1533
rect 5996 1527 6003 1533
rect 6036 1467 6043 1573
rect 6116 1527 6123 1553
rect 5916 1336 5963 1343
rect 5916 1327 5923 1336
rect 5956 1327 5963 1336
rect 5836 1296 5863 1303
rect 5716 1136 5743 1143
rect 5756 1236 5783 1243
rect 5693 1113 5707 1127
rect 5656 907 5663 933
rect 5676 927 5683 1093
rect 5696 907 5703 1073
rect 5716 907 5723 1136
rect 5733 1093 5747 1107
rect 5736 1067 5743 1093
rect 5756 1047 5763 1236
rect 5836 1187 5843 1296
rect 5893 1293 5907 1307
rect 5913 1313 5927 1327
rect 5876 1267 5883 1293
rect 5896 1287 5903 1293
rect 5816 1147 5823 1153
rect 5813 1133 5827 1147
rect 5856 1143 5863 1233
rect 5776 1107 5783 1133
rect 5793 1113 5807 1127
rect 5836 1136 5863 1143
rect 5836 1127 5843 1136
rect 5896 1127 5903 1153
rect 5916 1127 5923 1233
rect 5936 1127 5943 1293
rect 6013 1293 6027 1307
rect 6033 1313 6047 1327
rect 6053 1293 6067 1307
rect 5993 1273 6007 1287
rect 5996 1227 6003 1273
rect 6016 1267 6023 1293
rect 6056 1283 6063 1293
rect 6036 1276 6063 1283
rect 6036 1247 6043 1276
rect 5833 1113 5847 1127
rect 5893 1113 5907 1127
rect 5913 1103 5927 1107
rect 5913 1096 5943 1103
rect 5913 1093 5927 1096
rect 5816 1047 5823 1093
rect 5936 1087 5943 1096
rect 5836 927 5843 1073
rect 5856 1047 5863 1073
rect 5876 887 5883 1073
rect 5956 1067 5963 1093
rect 6016 1103 6023 1153
rect 6036 1127 6043 1193
rect 6056 1127 6063 1253
rect 6076 1147 6083 1313
rect 6096 1207 6103 1513
rect 6116 1367 6123 1433
rect 6136 1343 6143 1553
rect 6156 1427 6163 1733
rect 6196 1727 6203 1773
rect 6236 1707 6243 1753
rect 6256 1683 6263 1753
rect 6236 1676 6263 1683
rect 6176 1607 6183 1633
rect 6216 1607 6223 1673
rect 6236 1667 6243 1676
rect 6256 1607 6263 1653
rect 6173 1593 6187 1607
rect 6213 1593 6227 1607
rect 6253 1593 6267 1607
rect 6236 1567 6243 1573
rect 6276 1567 6283 1776
rect 6313 1773 6327 1787
rect 6336 1796 6367 1803
rect 6316 1767 6323 1773
rect 6296 1647 6303 1753
rect 6316 1747 6323 1753
rect 6336 1727 6343 1796
rect 6353 1793 6367 1796
rect 6396 1707 6403 1853
rect 6436 1807 6443 1813
rect 6433 1793 6447 1807
rect 6456 1783 6463 1893
rect 6536 1867 6543 2093
rect 6556 2087 6563 2133
rect 6596 2107 6603 2173
rect 6553 2073 6567 2087
rect 6593 2083 6607 2087
rect 6636 2083 6643 2193
rect 6573 2053 6587 2067
rect 6593 2076 6643 2083
rect 6593 2073 6607 2076
rect 6496 1807 6503 1813
rect 6473 1783 6487 1787
rect 6456 1776 6487 1783
rect 6493 1793 6507 1807
rect 6556 1787 6563 2033
rect 6576 2007 6583 2053
rect 6656 2007 6663 2113
rect 6576 1987 6583 1993
rect 6473 1773 6487 1776
rect 6313 1573 6327 1587
rect 6316 1567 6323 1573
rect 6127 1336 6143 1343
rect 6136 1327 6143 1336
rect 6176 1327 6183 1373
rect 6196 1347 6203 1513
rect 6256 1327 6263 1413
rect 6277 1358 6285 1382
rect 6133 1313 6147 1327
rect 6173 1313 6187 1327
rect 6193 1303 6207 1307
rect 6253 1303 6267 1307
rect 6193 1296 6223 1303
rect 6193 1293 6207 1296
rect 6116 1247 6123 1273
rect 6116 1147 6123 1173
rect 6053 1113 6067 1127
rect 6033 1103 6047 1107
rect 6016 1096 6047 1103
rect 6033 1093 6047 1096
rect 6073 1093 6087 1107
rect 6116 1107 6123 1113
rect 6113 1093 6127 1107
rect 6013 1073 6027 1087
rect 6076 1083 6083 1093
rect 6076 1076 6103 1083
rect 5936 887 5943 1053
rect 5656 867 5663 873
rect 5653 853 5667 867
rect 5673 833 5687 847
rect 5473 643 5487 647
rect 5453 613 5467 627
rect 5473 636 5503 643
rect 5473 633 5487 636
rect 5456 567 5463 613
rect 5436 447 5443 553
rect 5476 443 5483 533
rect 5496 487 5503 636
rect 5573 613 5587 627
rect 5476 436 5503 443
rect 5133 353 5147 367
rect 5173 353 5187 367
rect 5193 333 5207 347
rect 5096 207 5103 293
rect 4976 167 4983 173
rect 4933 153 4947 167
rect 4973 153 4987 167
rect 4877 78 4885 102
rect 5016 84 5024 196
rect 5096 147 5103 193
rect 5156 167 5163 313
rect 5196 227 5203 333
rect 5233 333 5247 347
rect 5333 353 5347 367
rect 5373 333 5387 347
rect 5236 327 5243 333
rect 5213 313 5227 327
rect 5216 187 5223 313
rect 5256 167 5263 253
rect 5336 247 5343 273
rect 5093 133 5107 147
rect 5133 133 5147 147
rect 5153 153 5167 167
rect 5136 127 5143 133
rect 5256 123 5263 153
rect 5273 123 5287 127
rect 5256 116 5287 123
rect 5313 123 5327 127
rect 5336 123 5343 233
rect 5376 227 5383 333
rect 5413 333 5427 347
rect 5436 327 5443 393
rect 5456 367 5463 413
rect 5496 367 5503 436
rect 5453 353 5467 367
rect 5493 353 5507 367
rect 5536 363 5543 593
rect 5576 587 5583 613
rect 5616 427 5623 693
rect 5636 567 5643 793
rect 5676 787 5683 833
rect 5676 667 5683 693
rect 5696 667 5703 813
rect 5716 727 5723 873
rect 5893 853 5907 867
rect 5913 833 5927 847
rect 5773 823 5787 827
rect 5773 816 5803 823
rect 5773 813 5787 816
rect 5776 723 5783 793
rect 5796 787 5803 816
rect 5876 747 5883 833
rect 5916 807 5923 833
rect 5936 747 5943 873
rect 5956 847 5963 1053
rect 5976 784 5984 896
rect 5756 716 5783 723
rect 5756 667 5763 716
rect 5856 683 5863 713
rect 5896 703 5903 733
rect 5836 676 5863 683
rect 5876 696 5903 703
rect 5836 667 5843 676
rect 5673 653 5687 667
rect 5753 653 5767 667
rect 5653 633 5667 647
rect 5693 643 5707 647
rect 5693 636 5723 643
rect 5693 633 5707 636
rect 5716 627 5723 636
rect 5733 633 5747 647
rect 5833 653 5847 667
rect 5773 633 5787 647
rect 5813 643 5827 647
rect 5796 636 5827 643
rect 5856 647 5863 653
rect 5876 647 5883 696
rect 5896 667 5903 673
rect 5916 667 5923 713
rect 5893 653 5907 667
rect 5573 373 5587 387
rect 5553 363 5567 367
rect 5536 356 5567 363
rect 5553 353 5567 356
rect 5473 313 5487 327
rect 5476 267 5483 313
rect 5273 113 5287 116
rect 5313 116 5343 123
rect 5397 116 5405 196
rect 5456 167 5463 173
rect 5453 153 5467 167
rect 5313 113 5327 116
rect 5136 107 5143 113
rect 5397 78 5405 102
rect 5536 84 5544 196
rect 5556 167 5563 353
rect 5636 243 5643 553
rect 5696 427 5703 593
rect 5796 487 5803 636
rect 5813 633 5827 636
rect 5873 633 5887 647
rect 5896 487 5903 613
rect 5936 567 5943 713
rect 5956 627 5963 693
rect 5996 667 6003 853
rect 6013 813 6027 827
rect 6036 823 6043 1013
rect 6076 847 6083 1053
rect 6096 967 6103 1076
rect 6116 987 6123 1033
rect 6053 823 6067 827
rect 6036 816 6067 823
rect 6053 813 6067 816
rect 6016 787 6023 813
rect 6056 807 6063 813
rect 6056 707 6063 733
rect 5993 653 6007 667
rect 6076 663 6083 833
rect 6096 683 6103 913
rect 6115 878 6123 902
rect 6115 784 6123 864
rect 6136 827 6143 1173
rect 6156 927 6163 1193
rect 6176 1127 6183 1273
rect 6196 1187 6203 1273
rect 6216 1163 6223 1296
rect 6236 1296 6267 1303
rect 6236 1227 6243 1296
rect 6253 1293 6267 1296
rect 6277 1264 6285 1344
rect 6196 1156 6223 1163
rect 6196 1147 6203 1156
rect 6193 1133 6207 1147
rect 6173 1113 6187 1127
rect 6236 1127 6243 1193
rect 6256 1147 6263 1193
rect 6276 1187 6283 1213
rect 6253 1133 6267 1147
rect 6213 1123 6227 1127
rect 6233 1123 6247 1127
rect 6213 1116 6247 1123
rect 6213 1113 6227 1116
rect 6233 1113 6247 1116
rect 6256 967 6263 1093
rect 6296 867 6303 1533
rect 6336 1343 6343 1633
rect 6356 1607 6363 1633
rect 6396 1627 6403 1633
rect 6353 1593 6367 1607
rect 6413 1583 6427 1587
rect 6436 1583 6443 1653
rect 6413 1576 6443 1583
rect 6413 1573 6427 1576
rect 6416 1467 6423 1573
rect 6316 1336 6343 1343
rect 6316 867 6323 1336
rect 6333 1293 6347 1307
rect 6356 1303 6363 1353
rect 6373 1303 6387 1307
rect 6356 1296 6387 1303
rect 6373 1293 6387 1296
rect 6336 1287 6343 1293
rect 6336 1167 6343 1273
rect 6416 1264 6424 1376
rect 6333 1113 6347 1127
rect 6336 1067 6343 1113
rect 6357 1076 6365 1156
rect 6396 1087 6403 1173
rect 6456 1163 6463 1693
rect 6497 1556 6505 1636
rect 6497 1518 6505 1542
rect 6516 1427 6523 1753
rect 6553 1603 6567 1607
rect 6536 1596 6567 1603
rect 6536 1407 6543 1596
rect 6553 1593 6567 1596
rect 6517 1358 6525 1382
rect 6517 1264 6525 1344
rect 6536 1287 6543 1393
rect 6556 1263 6563 1413
rect 6576 1343 6583 1853
rect 6636 1827 6643 1833
rect 6633 1813 6647 1827
rect 6596 1607 6603 1673
rect 6593 1593 6607 1607
rect 6636 1524 6644 1636
rect 6656 1587 6663 1953
rect 6676 1447 6683 2233
rect 6696 2067 6703 2336
rect 6716 2327 6723 5113
rect 6716 1947 6723 2293
rect 6736 2107 6743 6373
rect 6576 1336 6603 1343
rect 6573 1293 6587 1307
rect 6576 1287 6583 1293
rect 6536 1256 6563 1263
rect 6456 1156 6483 1163
rect 6416 1127 6423 1153
rect 6456 1127 6463 1133
rect 6413 1123 6427 1127
rect 6413 1116 6443 1123
rect 6413 1113 6427 1116
rect 6357 1038 6365 1062
rect 6436 1027 6443 1116
rect 6453 1113 6467 1127
rect 6456 887 6463 1013
rect 6476 1007 6483 1156
rect 6496 1044 6504 1156
rect 6156 856 6203 863
rect 6156 727 6163 856
rect 6196 847 6203 856
rect 6173 813 6187 827
rect 6193 833 6207 847
rect 6233 833 6247 847
rect 6236 827 6243 833
rect 6213 813 6227 827
rect 6176 767 6183 813
rect 6216 787 6223 813
rect 6096 676 6123 683
rect 6116 667 6123 676
rect 6076 656 6103 663
rect 6013 633 6027 647
rect 6033 633 6047 647
rect 6053 613 6067 627
rect 6096 627 6103 656
rect 6176 647 6183 653
rect 6196 647 6203 673
rect 6173 633 6187 647
rect 5676 367 5683 413
rect 5673 353 5687 367
rect 5693 333 5707 347
rect 5636 236 5663 243
rect 5637 116 5645 196
rect 5656 127 5663 236
rect 5696 203 5703 333
rect 5696 196 5723 203
rect 5696 167 5703 173
rect 5693 153 5707 167
rect 5716 163 5723 196
rect 5736 183 5743 413
rect 5816 387 5823 413
rect 5773 383 5787 387
rect 5756 376 5787 383
rect 5756 287 5763 376
rect 5773 373 5787 376
rect 5813 373 5827 387
rect 5896 367 5903 453
rect 5936 383 5943 553
rect 5956 467 5963 593
rect 5976 387 5983 593
rect 6036 387 6043 573
rect 6056 567 6063 613
rect 6216 583 6223 633
rect 6236 607 6243 753
rect 6256 647 6263 853
rect 6393 863 6407 867
rect 6376 856 6407 863
rect 6433 863 6447 867
rect 6273 813 6287 827
rect 6276 787 6283 813
rect 6356 747 6363 853
rect 6316 627 6323 733
rect 6253 593 6267 607
rect 6293 603 6307 607
rect 6316 603 6323 613
rect 6293 596 6323 603
rect 6293 593 6307 596
rect 6256 587 6263 593
rect 6216 576 6243 583
rect 6116 487 6123 493
rect 5936 376 5963 383
rect 5956 367 5963 376
rect 6056 367 6063 433
rect 5893 353 5907 367
rect 5933 333 5947 347
rect 5953 353 5967 367
rect 5816 207 5823 333
rect 5936 267 5943 333
rect 5936 247 5943 253
rect 5736 176 5763 183
rect 5756 167 5763 176
rect 5733 163 5747 167
rect 5716 156 5747 163
rect 5733 153 5747 156
rect 5637 78 5645 102
rect 5776 84 5784 196
rect 5877 116 5885 196
rect 5936 167 5943 173
rect 5956 167 5963 313
rect 5996 307 6003 353
rect 6033 333 6047 347
rect 6093 363 6107 367
rect 6116 363 6123 473
rect 6136 407 6143 413
rect 6236 407 6243 576
rect 6256 367 6263 573
rect 6336 447 6343 693
rect 6356 564 6364 676
rect 6376 587 6383 856
rect 6393 853 6407 856
rect 6433 856 6453 863
rect 6433 853 6447 856
rect 6396 647 6403 653
rect 6436 647 6443 793
rect 6393 633 6407 647
rect 6433 643 6447 647
rect 6433 636 6463 643
rect 6433 633 6447 636
rect 6276 383 6283 433
rect 6316 387 6323 413
rect 6276 376 6303 383
rect 6093 356 6123 363
rect 6093 353 6107 356
rect 6073 333 6087 347
rect 5976 167 5983 193
rect 5933 153 5947 167
rect 5973 153 5987 167
rect 5996 147 6003 293
rect 5877 78 5885 102
rect 6016 84 6024 196
rect 6056 67 6063 313
rect 6076 267 6083 333
rect 6096 167 6103 273
rect 6116 227 6123 356
rect 6136 307 6143 353
rect 6193 333 6207 347
rect 6233 333 6247 347
rect 6273 343 6287 347
rect 6296 343 6303 376
rect 6376 367 6383 473
rect 6396 387 6403 593
rect 6456 467 6463 636
rect 6236 327 6243 333
rect 6273 336 6303 343
rect 6273 333 6287 336
rect 6353 333 6367 347
rect 6373 353 6387 367
rect 6173 313 6187 327
rect 6253 313 6267 327
rect 6356 323 6363 333
rect 6416 323 6423 333
rect 6356 316 6423 323
rect 6156 267 6163 313
rect 6176 207 6183 313
rect 6236 307 6243 313
rect 6093 153 6107 167
rect 6153 133 6167 147
rect 6196 147 6203 213
rect 6156 127 6163 133
rect 6216 127 6223 293
rect 6256 267 6263 313
rect 6276 287 6283 313
rect 6296 207 6303 313
rect 6316 267 6323 313
rect 6456 304 6464 416
rect 6476 307 6483 953
rect 6496 784 6504 896
rect 6516 687 6523 1153
rect 6536 867 6543 1256
rect 6556 1147 6563 1233
rect 6596 1167 6603 1336
rect 6613 1293 6627 1307
rect 6616 1143 6623 1293
rect 6656 1264 6664 1376
rect 6676 1327 6683 1433
rect 6596 1136 6623 1143
rect 6596 1127 6603 1136
rect 6636 1127 6643 1173
rect 6573 1093 6587 1107
rect 6593 1113 6607 1127
rect 6633 1113 6647 1127
rect 6656 1107 6663 1193
rect 6556 783 6563 1073
rect 6576 987 6583 1093
rect 6656 987 6663 1073
rect 6573 813 6587 827
rect 6576 807 6583 813
rect 6556 776 6583 783
rect 6495 596 6503 676
rect 6513 633 6527 647
rect 6516 627 6523 633
rect 6495 558 6503 582
rect 6516 343 6523 453
rect 6536 387 6543 673
rect 6556 667 6563 673
rect 6576 667 6583 776
rect 6553 653 6567 667
rect 6596 487 6603 973
rect 6676 907 6683 1293
rect 6696 1267 6703 1873
rect 6716 1027 6723 1313
rect 6736 1227 6743 1913
rect 6736 1067 6743 1213
rect 6616 667 6623 893
rect 6635 878 6643 902
rect 6635 784 6643 864
rect 6656 827 6663 853
rect 6653 813 6667 827
rect 6613 653 6627 667
rect 6633 623 6647 627
rect 6656 623 6663 653
rect 6633 616 6663 623
rect 6633 613 6647 616
rect 6595 398 6603 422
rect 6533 343 6547 347
rect 6516 336 6547 343
rect 6236 107 6243 193
rect 6396 187 6403 193
rect 6393 173 6407 187
rect 6273 133 6287 147
rect 6333 163 6347 167
rect 6333 156 6363 163
rect 6333 153 6347 156
rect 6356 143 6363 156
rect 6416 163 6423 193
rect 6433 163 6447 167
rect 6416 156 6447 163
rect 6433 153 6447 156
rect 6373 143 6387 147
rect 6356 136 6387 143
rect 6373 133 6387 136
rect 6276 107 6283 133
rect 6457 116 6465 196
rect 6516 187 6523 336
rect 6533 333 6547 336
rect 6595 304 6603 384
rect 6616 347 6623 373
rect 6613 333 6627 347
rect 6716 247 6723 973
rect 6516 167 6523 173
rect 6513 153 6527 167
rect 6457 78 6465 102
rect 6596 84 6604 196
<< m3contact >>
rect 4393 6493 4407 6507
rect 4753 6493 4767 6507
rect 4893 6493 4907 6507
rect 5893 6493 5907 6507
rect 4333 6473 4347 6487
rect 3093 6453 3107 6467
rect 3453 6453 3467 6467
rect 133 6413 147 6427
rect 153 6413 167 6427
rect 93 6393 107 6407
rect 33 6093 47 6107
rect 293 6393 307 6407
rect 273 6373 287 6387
rect 333 6393 347 6407
rect 413 6393 427 6407
rect 433 6393 447 6407
rect 213 6353 227 6367
rect 353 6353 367 6367
rect 373 6373 387 6387
rect 393 6333 407 6347
rect 413 6333 427 6347
rect 73 6093 87 6107
rect 153 6093 167 6107
rect 113 6053 127 6067
rect 313 6173 327 6187
rect 393 6153 407 6167
rect 533 6393 547 6407
rect 573 6393 587 6407
rect 613 6393 627 6407
rect 453 6353 467 6367
rect 493 6353 507 6367
rect 513 6353 527 6367
rect 613 6373 627 6387
rect 733 6433 747 6447
rect 693 6413 707 6427
rect 673 6353 687 6367
rect 493 6293 507 6307
rect 373 6133 387 6147
rect 233 6113 247 6127
rect 13 5873 27 5887
rect 53 5873 67 5887
rect 93 5873 107 5887
rect 193 5893 207 5907
rect 273 6093 287 6107
rect 293 6113 307 6127
rect 333 6113 347 6127
rect 413 6133 427 6147
rect 373 6093 387 6107
rect 313 6073 327 6087
rect 513 6173 527 6187
rect 533 6133 547 6147
rect 513 6113 527 6127
rect 553 6113 567 6127
rect 573 6133 587 6147
rect 413 6073 427 6087
rect 373 6053 387 6067
rect 393 6053 407 6067
rect 393 5953 407 5967
rect 313 5933 327 5947
rect 233 5873 247 5887
rect 133 5853 147 5867
rect 33 5613 47 5627
rect 33 5413 47 5427
rect 213 5853 227 5867
rect 113 5593 127 5607
rect 513 6093 527 6107
rect 553 6093 567 6107
rect 613 6113 627 6127
rect 653 6113 667 6127
rect 653 6093 667 6107
rect 453 6073 467 6087
rect 553 6073 567 6087
rect 513 6033 527 6047
rect 493 5993 507 6007
rect 433 5953 447 5967
rect 413 5933 427 5947
rect 413 5913 427 5927
rect 333 5893 347 5907
rect 293 5873 307 5887
rect 333 5873 347 5887
rect 373 5873 387 5887
rect 413 5873 427 5887
rect 453 5873 467 5887
rect 253 5613 267 5627
rect 113 5453 127 5467
rect 173 5453 187 5467
rect 93 5413 107 5427
rect 153 5433 167 5447
rect 33 5133 47 5147
rect 113 5153 127 5167
rect 73 5133 87 5147
rect 113 5133 127 5147
rect 533 5973 547 5987
rect 513 5933 527 5947
rect 513 5913 527 5927
rect 613 6033 627 6047
rect 613 5993 627 6007
rect 593 5933 607 5947
rect 533 5893 547 5907
rect 573 5913 587 5927
rect 653 5973 667 5987
rect 933 6433 947 6447
rect 793 6373 807 6387
rect 813 6373 827 6387
rect 873 6373 887 6387
rect 853 6353 867 6367
rect 913 6353 927 6367
rect 813 6333 827 6347
rect 753 6153 767 6167
rect 873 6273 887 6287
rect 953 6273 967 6287
rect 833 6153 847 6167
rect 713 6093 727 6107
rect 733 6093 747 6107
rect 813 6113 827 6127
rect 693 6073 707 6087
rect 693 6033 707 6047
rect 673 5933 687 5947
rect 633 5913 647 5927
rect 493 5833 507 5847
rect 313 5613 327 5627
rect 273 5453 287 5467
rect 253 5393 267 5407
rect 273 5413 287 5427
rect 293 5373 307 5387
rect 693 5913 707 5927
rect 773 6073 787 6087
rect 753 5973 767 5987
rect 733 5913 747 5927
rect 633 5873 647 5887
rect 653 5873 667 5887
rect 573 5853 587 5867
rect 513 5653 527 5667
rect 533 5653 547 5667
rect 433 5613 447 5627
rect 493 5633 507 5647
rect 453 5593 467 5607
rect 453 5573 467 5587
rect 513 5593 527 5607
rect 473 5553 487 5567
rect 433 5533 447 5547
rect 333 5473 347 5487
rect 313 5353 327 5367
rect 73 5013 87 5027
rect 33 4953 47 4967
rect 113 4953 127 4967
rect 153 4953 167 4967
rect 193 5113 207 5127
rect 233 5093 247 5107
rect 393 5453 407 5467
rect 353 5433 367 5447
rect 533 5533 547 5547
rect 553 5533 567 5547
rect 493 5493 507 5507
rect 513 5453 527 5467
rect 413 5393 427 5407
rect 453 5393 467 5407
rect 533 5393 547 5407
rect 553 5393 567 5407
rect 633 5673 647 5687
rect 593 5653 607 5667
rect 633 5653 647 5667
rect 593 5613 607 5627
rect 593 5533 607 5547
rect 633 5613 647 5627
rect 613 5513 627 5527
rect 613 5493 627 5507
rect 673 5833 687 5847
rect 733 5713 747 5727
rect 673 5693 687 5707
rect 673 5653 687 5667
rect 1033 6373 1047 6387
rect 1213 6433 1227 6447
rect 1173 6413 1187 6427
rect 1193 6373 1207 6387
rect 1073 6293 1087 6307
rect 993 6153 1007 6167
rect 1053 6153 1067 6167
rect 913 6113 927 6127
rect 953 6113 967 6127
rect 813 6033 827 6047
rect 793 5973 807 5987
rect 793 5953 807 5967
rect 1013 6113 1027 6127
rect 933 6053 947 6067
rect 893 6033 907 6047
rect 893 5953 907 5967
rect 773 5933 787 5947
rect 853 5933 867 5947
rect 813 5913 827 5927
rect 873 5913 887 5927
rect 813 5873 827 5887
rect 773 5853 787 5867
rect 873 5853 887 5867
rect 813 5673 827 5687
rect 993 6053 1007 6067
rect 993 5953 1007 5967
rect 973 5913 987 5927
rect 1093 6113 1107 6127
rect 1133 6093 1147 6107
rect 1013 5913 1027 5927
rect 913 5873 927 5887
rect 933 5893 947 5907
rect 973 5893 987 5907
rect 1033 5893 1047 5907
rect 1053 5913 1067 5927
rect 1073 5913 1087 5927
rect 1113 5913 1127 5927
rect 1093 5893 1107 5907
rect 913 5713 927 5727
rect 673 5613 687 5627
rect 593 5433 607 5447
rect 613 5433 627 5447
rect 653 5433 667 5447
rect 793 5633 807 5647
rect 813 5613 827 5627
rect 733 5593 747 5607
rect 693 5573 707 5587
rect 733 5533 747 5547
rect 693 5493 707 5507
rect 713 5473 727 5487
rect 793 5453 807 5467
rect 873 5613 887 5627
rect 833 5593 847 5607
rect 973 5833 987 5847
rect 953 5693 967 5707
rect 1053 5853 1067 5867
rect 1093 5853 1107 5867
rect 1033 5673 1047 5687
rect 933 5613 947 5627
rect 993 5633 1007 5647
rect 1033 5633 1047 5647
rect 993 5593 1007 5607
rect 953 5533 967 5547
rect 973 5533 987 5547
rect 913 5513 927 5527
rect 973 5513 987 5527
rect 873 5473 887 5487
rect 913 5473 927 5487
rect 733 5393 747 5407
rect 833 5413 847 5427
rect 573 5373 587 5387
rect 593 5373 607 5387
rect 673 5373 687 5387
rect 693 5373 707 5387
rect 373 5353 387 5367
rect 413 5353 427 5367
rect 533 5353 547 5367
rect 333 5193 347 5207
rect 373 5193 387 5207
rect 313 5153 327 5167
rect 353 5153 367 5167
rect 513 5213 527 5227
rect 573 5213 587 5227
rect 493 5173 507 5187
rect 413 5153 427 5167
rect 333 5133 347 5147
rect 273 4953 287 4967
rect 213 4933 227 4947
rect 233 4913 247 4927
rect 273 4913 287 4927
rect 193 4893 207 4907
rect 293 4773 307 4787
rect 173 4693 187 4707
rect 233 4653 247 4667
rect 353 5113 367 5127
rect 393 4953 407 4967
rect 453 5153 467 5167
rect 613 5353 627 5367
rect 593 5193 607 5207
rect 533 5173 547 5187
rect 553 5153 567 5167
rect 473 5113 487 5127
rect 513 5113 527 5127
rect 433 5093 447 5107
rect 553 4993 567 5007
rect 513 4953 527 4967
rect 533 4933 547 4947
rect 553 4933 567 4947
rect 573 4913 587 4927
rect 613 5153 627 5167
rect 673 5133 687 5147
rect 613 4993 627 5007
rect 633 4993 647 5007
rect 613 4953 627 4967
rect 773 5373 787 5387
rect 813 5373 827 5387
rect 773 5353 787 5367
rect 813 5193 827 5207
rect 713 5113 727 5127
rect 733 5113 747 5127
rect 793 5173 807 5187
rect 733 4993 747 5007
rect 1113 5673 1127 5687
rect 1093 5613 1107 5627
rect 1013 5573 1027 5587
rect 1053 5573 1067 5587
rect 1173 6053 1187 6067
rect 1153 6033 1167 6047
rect 1353 6433 1367 6447
rect 1633 6433 1647 6447
rect 1673 6433 1687 6447
rect 1293 6413 1307 6427
rect 1313 6393 1327 6407
rect 1373 6373 1387 6387
rect 1493 6373 1507 6387
rect 1333 6353 1347 6367
rect 1433 6353 1447 6367
rect 1553 6393 1567 6407
rect 1593 6373 1607 6387
rect 1533 6353 1547 6367
rect 1573 6353 1587 6367
rect 1213 6153 1227 6167
rect 1233 6093 1247 6107
rect 1273 6113 1287 6127
rect 1293 6093 1307 6107
rect 1193 5993 1207 6007
rect 1253 5993 1267 6007
rect 1153 5953 1167 5967
rect 1233 5953 1247 5967
rect 1213 5913 1227 5927
rect 1353 6153 1367 6167
rect 1433 6093 1447 6107
rect 1413 6073 1427 6087
rect 1453 6073 1467 6087
rect 1373 6053 1387 6067
rect 1553 6093 1567 6107
rect 1533 6073 1547 6087
rect 1613 6153 1627 6167
rect 1593 6133 1607 6147
rect 1653 6373 1667 6387
rect 1793 6413 1807 6427
rect 1753 6373 1767 6387
rect 1833 6393 1847 6407
rect 1713 6153 1727 6167
rect 1793 6353 1807 6367
rect 2313 6433 2327 6447
rect 2493 6433 2507 6447
rect 2893 6433 2907 6447
rect 2273 6413 2287 6427
rect 1913 6373 1927 6387
rect 1973 6393 1987 6407
rect 1993 6393 2007 6407
rect 2153 6393 2167 6407
rect 2053 6373 2067 6387
rect 2073 6353 2087 6367
rect 2013 6273 2027 6287
rect 1893 6233 1907 6247
rect 1953 6233 1967 6247
rect 2093 6313 2107 6327
rect 2033 6253 2047 6267
rect 2073 6153 2087 6167
rect 2053 6133 2067 6147
rect 2173 6373 2187 6387
rect 2193 6393 2207 6407
rect 2233 6393 2247 6407
rect 2273 6373 2287 6387
rect 2233 6353 2247 6367
rect 2113 6253 2127 6267
rect 2133 6153 2147 6167
rect 1633 6093 1647 6107
rect 1753 6113 1767 6127
rect 1593 6073 1607 6087
rect 1513 6053 1527 6067
rect 1573 6053 1587 6067
rect 1353 6033 1367 6047
rect 1473 6033 1487 6047
rect 1693 6093 1707 6107
rect 1713 6093 1727 6107
rect 1793 6113 1807 6127
rect 1673 6033 1687 6047
rect 1653 6013 1667 6027
rect 1693 6013 1707 6027
rect 1653 5993 1667 6007
rect 1233 5693 1247 5707
rect 1133 5633 1147 5647
rect 1133 5593 1147 5607
rect 1093 5533 1107 5547
rect 1113 5533 1127 5547
rect 1073 5513 1087 5527
rect 1073 5473 1087 5487
rect 1013 5413 1027 5427
rect 1053 5433 1067 5447
rect 1033 5393 1047 5407
rect 913 5373 927 5387
rect 853 5353 867 5367
rect 933 5213 947 5227
rect 873 5193 887 5207
rect 833 5173 847 5187
rect 853 5153 867 5167
rect 933 5153 947 5167
rect 953 5133 967 5147
rect 973 5153 987 5167
rect 1353 5913 1367 5927
rect 1473 5913 1487 5927
rect 1633 5913 1647 5927
rect 1773 6093 1787 6107
rect 1833 6113 1847 6127
rect 1873 6113 1887 6127
rect 1933 6113 1947 6127
rect 1973 6113 1987 6127
rect 1753 6073 1767 6087
rect 1773 6073 1787 6087
rect 1793 6073 1807 6087
rect 1753 6053 1767 6067
rect 1713 5973 1727 5987
rect 1733 5973 1747 5987
rect 1693 5933 1707 5947
rect 1793 5993 1807 6007
rect 1773 5953 1787 5967
rect 1813 5973 1827 5987
rect 1813 5953 1827 5967
rect 1673 5913 1687 5927
rect 1533 5893 1547 5907
rect 1493 5873 1507 5887
rect 1553 5873 1567 5887
rect 1573 5893 1587 5907
rect 1593 5873 1607 5887
rect 1533 5853 1547 5867
rect 1453 5833 1467 5847
rect 1273 5633 1287 5647
rect 1293 5633 1307 5647
rect 1233 5593 1247 5607
rect 1193 5573 1207 5587
rect 1213 5573 1227 5587
rect 1173 5553 1187 5567
rect 1253 5553 1267 5567
rect 1153 5473 1167 5487
rect 1133 5413 1147 5427
rect 1153 5433 1167 5447
rect 1073 5173 1087 5187
rect 1173 5393 1187 5407
rect 1153 5173 1167 5187
rect 1013 5133 1027 5147
rect 1073 5153 1087 5167
rect 1113 5153 1127 5167
rect 1093 5133 1107 5147
rect 993 5113 1007 5127
rect 1053 5113 1067 5127
rect 1013 5093 1027 5107
rect 1133 5093 1147 5107
rect 1033 5073 1047 5087
rect 1113 5073 1127 5087
rect 1193 5073 1207 5087
rect 893 5013 907 5027
rect 813 4973 827 4987
rect 693 4953 707 4967
rect 833 4953 847 4967
rect 613 4913 627 4927
rect 653 4913 667 4927
rect 673 4913 687 4927
rect 693 4933 707 4947
rect 733 4933 747 4947
rect 753 4933 767 4947
rect 713 4913 727 4927
rect 593 4893 607 4907
rect 413 4773 427 4787
rect 313 4673 327 4687
rect 333 4673 347 4687
rect 353 4653 367 4667
rect 373 4653 387 4667
rect 393 4673 407 4687
rect 433 4673 447 4687
rect 273 4613 287 4627
rect 253 4573 267 4587
rect 133 4553 147 4567
rect 73 4513 87 4527
rect 53 4493 67 4507
rect 113 4493 127 4507
rect 93 4473 107 4487
rect 213 4513 227 4527
rect 193 4493 207 4507
rect 33 4453 47 4467
rect 73 4453 87 4467
rect 293 4593 307 4607
rect 153 4453 167 4467
rect 173 4453 187 4467
rect 193 4453 207 4467
rect 233 4453 247 4467
rect 273 4473 287 4487
rect 333 4633 347 4647
rect 373 4633 387 4647
rect 353 4613 367 4627
rect 333 4593 347 4607
rect 333 4533 347 4547
rect 393 4573 407 4587
rect 353 4493 367 4507
rect 373 4493 387 4507
rect 313 4473 327 4487
rect 513 4673 527 4687
rect 533 4653 547 4667
rect 493 4633 507 4647
rect 513 4633 527 4647
rect 553 4633 567 4647
rect 573 4633 587 4647
rect 613 4873 627 4887
rect 633 4853 647 4867
rect 613 4653 627 4667
rect 793 4933 807 4947
rect 853 4933 867 4947
rect 813 4913 827 4927
rect 833 4913 847 4927
rect 973 4993 987 5007
rect 893 4933 907 4947
rect 953 4933 967 4947
rect 773 4893 787 4907
rect 833 4893 847 4907
rect 693 4873 707 4887
rect 753 4873 767 4887
rect 753 4853 767 4867
rect 733 4733 747 4747
rect 1053 5033 1067 5047
rect 1133 5033 1147 5047
rect 993 4793 1007 4807
rect 833 4693 847 4707
rect 653 4633 667 4647
rect 453 4553 467 4567
rect 413 4533 427 4547
rect 433 4533 447 4547
rect 413 4513 427 4527
rect 493 4533 507 4547
rect 513 4493 527 4507
rect 313 4453 327 4467
rect 353 4453 367 4467
rect 413 4453 427 4467
rect 433 4473 447 4487
rect 453 4473 467 4487
rect 513 4473 527 4487
rect 13 4433 27 4447
rect 153 4233 167 4247
rect 153 4213 167 4227
rect 333 4393 347 4407
rect 33 4173 47 4187
rect 173 4173 187 4187
rect 273 4193 287 4207
rect 253 4173 267 4187
rect 73 4153 87 4167
rect 273 4153 287 4167
rect 233 4133 247 4147
rect 473 4413 487 4427
rect 373 4393 387 4407
rect 553 4253 567 4267
rect 613 4493 627 4507
rect 593 4453 607 4467
rect 613 4453 627 4467
rect 593 4253 607 4267
rect 373 4213 387 4227
rect 433 4213 447 4227
rect 573 4233 587 4247
rect 593 4233 607 4247
rect 433 4173 447 4187
rect 413 4153 427 4167
rect 453 4153 467 4167
rect 373 4133 387 4147
rect 353 4113 367 4127
rect 413 4113 427 4127
rect 73 3993 87 4007
rect 113 3993 127 4007
rect 53 3953 67 3967
rect 113 3953 127 3967
rect 193 4013 207 4027
rect 233 3993 247 4007
rect 553 4193 567 4207
rect 573 4213 587 4227
rect 453 4013 467 4027
rect 473 4013 487 4027
rect 433 3993 447 4007
rect 333 3953 347 3967
rect 353 3973 367 3987
rect 413 3973 427 3987
rect 453 3973 467 3987
rect 373 3933 387 3947
rect 193 3753 207 3767
rect 33 3693 47 3707
rect 213 3713 227 3727
rect 153 3693 167 3707
rect 253 3693 267 3707
rect 113 3673 127 3687
rect 73 3653 87 3667
rect 393 3693 407 3707
rect 353 3673 367 3687
rect 493 3953 507 3967
rect 553 4013 567 4027
rect 533 3953 547 3967
rect 573 3953 587 3967
rect 633 4393 647 4407
rect 633 4213 647 4227
rect 813 4673 827 4687
rect 833 4653 847 4667
rect 793 4633 807 4647
rect 813 4633 827 4647
rect 893 4673 907 4687
rect 913 4693 927 4707
rect 933 4693 947 4707
rect 893 4653 907 4667
rect 713 4613 727 4627
rect 813 4613 827 4627
rect 853 4613 867 4627
rect 773 4573 787 4587
rect 733 4533 747 4547
rect 733 4513 747 4527
rect 793 4513 807 4527
rect 753 4473 767 4487
rect 713 4413 727 4427
rect 953 4593 967 4607
rect 913 4533 927 4547
rect 833 4493 847 4507
rect 893 4493 907 4507
rect 853 4453 867 4467
rect 893 4473 907 4487
rect 933 4473 947 4487
rect 913 4453 927 4467
rect 693 4253 707 4267
rect 813 4393 827 4407
rect 753 4253 767 4267
rect 793 4213 807 4227
rect 813 4213 827 4227
rect 673 4133 687 4147
rect 673 4113 687 4127
rect 613 4013 627 4027
rect 633 3993 647 4007
rect 633 3973 647 3987
rect 653 3953 667 3967
rect 713 4093 727 4107
rect 693 4033 707 4047
rect 733 4013 747 4027
rect 733 3993 747 4007
rect 593 3933 607 3947
rect 453 3913 467 3927
rect 573 3773 587 3787
rect 653 3773 667 3787
rect 673 3773 687 3787
rect 593 3753 607 3767
rect 473 3673 487 3687
rect 453 3613 467 3627
rect 413 3593 427 3607
rect 453 3593 467 3607
rect 233 3573 247 3587
rect 33 3513 47 3527
rect 73 3513 87 3527
rect 113 3513 127 3527
rect 113 3473 127 3487
rect 193 3533 207 3547
rect 213 3493 227 3507
rect 213 3433 227 3447
rect 413 3553 427 3567
rect 533 3733 547 3747
rect 513 3693 527 3707
rect 573 3713 587 3727
rect 553 3673 567 3687
rect 493 3633 507 3647
rect 553 3633 567 3647
rect 513 3573 527 3587
rect 553 3573 567 3587
rect 473 3533 487 3547
rect 313 3513 327 3527
rect 413 3513 427 3527
rect 33 3213 47 3227
rect 113 3233 127 3247
rect 73 3213 87 3227
rect 113 3213 127 3227
rect 233 3213 247 3227
rect 233 3033 247 3047
rect 193 3013 207 3027
rect 293 2933 307 2947
rect 33 2753 47 2767
rect 93 2733 107 2747
rect 113 2713 127 2727
rect 133 2713 147 2727
rect 53 2633 67 2647
rect 113 2593 127 2607
rect 153 2693 167 2707
rect 233 2733 247 2747
rect 253 2633 267 2647
rect 153 2573 167 2587
rect 153 2513 167 2527
rect 93 2253 107 2267
rect 53 2173 67 2187
rect 73 2093 87 2107
rect 233 2273 247 2287
rect 213 2253 227 2267
rect 233 2233 247 2247
rect 213 2213 227 2227
rect 233 2213 247 2227
rect 173 2173 187 2187
rect 213 2113 227 2127
rect 133 2093 147 2107
rect 173 2093 187 2107
rect 213 2093 227 2107
rect 53 2053 67 2067
rect 73 2033 87 2047
rect 53 1993 67 2007
rect 173 2073 187 2087
rect 153 2033 167 2047
rect 93 2013 107 2027
rect 113 1993 127 2007
rect 73 1973 87 1987
rect 193 2033 207 2047
rect 333 3473 347 3487
rect 353 3493 367 3507
rect 373 3473 387 3487
rect 413 3293 427 3307
rect 373 3273 387 3287
rect 333 3253 347 3267
rect 353 3233 367 3247
rect 453 3253 467 3267
rect 533 3493 547 3507
rect 773 4113 787 4127
rect 873 4213 887 4227
rect 853 4173 867 4187
rect 793 4093 807 4107
rect 773 3993 787 4007
rect 773 3953 787 3967
rect 893 4173 907 4187
rect 893 4153 907 4167
rect 873 4113 887 4127
rect 893 4053 907 4067
rect 753 3913 767 3927
rect 753 3773 767 3787
rect 773 3773 787 3787
rect 813 3773 827 3787
rect 733 3733 747 3747
rect 733 3713 747 3727
rect 693 3673 707 3687
rect 773 3753 787 3767
rect 793 3713 807 3727
rect 853 3773 867 3787
rect 693 3633 707 3647
rect 733 3633 747 3647
rect 633 3613 647 3627
rect 733 3553 747 3567
rect 753 3553 767 3567
rect 833 3693 847 3707
rect 853 3693 867 3707
rect 893 3693 907 3707
rect 933 4133 947 4147
rect 933 3673 947 3687
rect 893 3653 907 3667
rect 913 3653 927 3667
rect 853 3573 867 3587
rect 793 3533 807 3547
rect 693 3513 707 3527
rect 713 3513 727 3527
rect 593 3473 607 3487
rect 633 3493 647 3507
rect 573 3453 587 3467
rect 493 3293 507 3307
rect 573 3293 587 3307
rect 613 3453 627 3467
rect 653 3453 667 3467
rect 673 3453 687 3467
rect 613 3313 627 3327
rect 593 3273 607 3287
rect 413 3233 427 3247
rect 433 3213 447 3227
rect 473 3233 487 3247
rect 633 3293 647 3307
rect 653 3273 667 3287
rect 773 3513 787 3527
rect 813 3513 827 3527
rect 773 3493 787 3507
rect 973 4513 987 4527
rect 993 4453 1007 4467
rect 1033 4633 1047 4647
rect 1093 4973 1107 4987
rect 1193 5013 1207 5027
rect 1173 4993 1187 5007
rect 1313 5613 1327 5627
rect 1433 5633 1447 5647
rect 1333 5593 1347 5607
rect 1353 5593 1367 5607
rect 1433 5593 1447 5607
rect 1393 5573 1407 5587
rect 1453 5573 1467 5587
rect 1593 5613 1607 5627
rect 1553 5593 1567 5607
rect 1293 5453 1307 5467
rect 1313 5453 1327 5467
rect 1353 5433 1367 5447
rect 1233 5373 1247 5387
rect 1693 5893 1707 5907
rect 1793 5913 1807 5927
rect 1773 5893 1787 5907
rect 1913 6053 1927 6067
rect 1913 5973 1927 5987
rect 1873 5913 1887 5927
rect 1833 5873 1847 5887
rect 1953 5913 1967 5927
rect 1893 5893 1907 5907
rect 1933 5893 1947 5907
rect 1953 5893 1967 5907
rect 1873 5873 1887 5887
rect 1913 5873 1927 5887
rect 1933 5873 1947 5887
rect 1813 5853 1827 5867
rect 1893 5813 1907 5827
rect 1873 5673 1887 5687
rect 1673 5633 1687 5647
rect 1733 5613 1747 5627
rect 1753 5633 1767 5647
rect 1893 5653 1907 5667
rect 1833 5613 1847 5627
rect 1893 5613 1907 5627
rect 1773 5593 1787 5607
rect 1813 5533 1827 5547
rect 1533 5433 1547 5447
rect 1653 5453 1667 5467
rect 1693 5453 1707 5467
rect 1733 5453 1747 5467
rect 1773 5453 1787 5467
rect 1493 5413 1507 5427
rect 1513 5393 1527 5407
rect 1573 5393 1587 5407
rect 1713 5433 1727 5447
rect 1753 5433 1767 5447
rect 1613 5393 1627 5407
rect 1673 5413 1687 5427
rect 1653 5393 1667 5407
rect 1693 5393 1707 5407
rect 1233 5153 1247 5167
rect 1233 5133 1247 5147
rect 1233 5093 1247 5107
rect 1373 5173 1387 5187
rect 1313 5113 1327 5127
rect 1213 4993 1227 5007
rect 1253 5013 1267 5027
rect 1153 4953 1167 4967
rect 1193 4933 1207 4947
rect 1153 4913 1167 4927
rect 1173 4913 1187 4927
rect 1233 4913 1247 4927
rect 1073 4653 1087 4667
rect 1113 4573 1127 4587
rect 1153 4573 1167 4587
rect 1053 4493 1067 4507
rect 973 3613 987 3627
rect 953 3553 967 3567
rect 933 3513 947 3527
rect 853 3493 867 3507
rect 913 3493 927 3507
rect 773 3453 787 3467
rect 833 3313 847 3327
rect 633 3253 647 3267
rect 593 3233 607 3247
rect 513 3213 527 3227
rect 553 3213 567 3227
rect 573 3213 587 3227
rect 453 3193 467 3207
rect 473 3193 487 3207
rect 373 3093 387 3107
rect 413 3033 427 3047
rect 553 3193 567 3207
rect 513 3173 527 3187
rect 453 3013 467 3027
rect 513 3053 527 3067
rect 653 3233 667 3247
rect 633 3213 647 3227
rect 633 3193 647 3207
rect 693 3233 707 3247
rect 713 3253 727 3267
rect 753 3253 767 3267
rect 693 3213 707 3227
rect 733 3213 747 3227
rect 753 3213 767 3227
rect 593 3173 607 3187
rect 673 3173 687 3187
rect 673 3073 687 3087
rect 673 3053 687 3067
rect 553 3033 567 3047
rect 573 3033 587 3047
rect 633 3033 647 3047
rect 753 3153 767 3167
rect 733 3093 747 3107
rect 753 3093 767 3107
rect 893 3313 907 3327
rect 873 3293 887 3307
rect 973 3513 987 3527
rect 1053 4433 1067 4447
rect 1053 4373 1067 4387
rect 1073 4233 1087 4247
rect 1013 4193 1027 4207
rect 1053 4193 1067 4207
rect 1213 4893 1227 4907
rect 1233 4873 1247 4887
rect 1673 5373 1687 5387
rect 1613 5333 1627 5347
rect 1513 5193 1527 5207
rect 1493 5153 1507 5167
rect 1533 5173 1547 5187
rect 1553 5153 1567 5167
rect 1393 5033 1407 5047
rect 1353 4993 1367 5007
rect 1353 4973 1367 4987
rect 1573 4993 1587 5007
rect 1493 4973 1507 4987
rect 1313 4953 1327 4967
rect 1273 4913 1287 4927
rect 1293 4933 1307 4947
rect 1333 4933 1347 4947
rect 1433 4933 1447 4947
rect 1533 4933 1547 4947
rect 1313 4893 1327 4907
rect 1413 4893 1427 4907
rect 1273 4873 1287 4887
rect 1453 4873 1467 4887
rect 1553 4873 1567 4887
rect 1253 4793 1267 4807
rect 1233 4693 1247 4707
rect 1333 4773 1347 4787
rect 1393 4773 1407 4787
rect 1293 4713 1307 4727
rect 1353 4753 1367 4767
rect 1413 4753 1427 4767
rect 1193 4673 1207 4687
rect 1213 4653 1227 4667
rect 1273 4673 1287 4687
rect 1313 4673 1327 4687
rect 1373 4673 1387 4687
rect 1353 4653 1367 4667
rect 1273 4613 1287 4627
rect 1233 4513 1247 4527
rect 1233 4493 1247 4507
rect 1353 4573 1367 4587
rect 1393 4653 1407 4667
rect 1373 4553 1387 4567
rect 1553 4733 1567 4747
rect 1673 5313 1687 5327
rect 1733 5413 1747 5427
rect 1773 5413 1787 5427
rect 1793 5433 1807 5447
rect 1833 5453 1847 5467
rect 2073 6113 2087 6127
rect 2093 6113 2107 6127
rect 1993 6073 2007 6087
rect 2033 6073 2047 6087
rect 2133 6133 2147 6147
rect 2193 6133 2207 6147
rect 2293 6353 2307 6367
rect 2273 6333 2287 6347
rect 2253 6293 2267 6307
rect 2433 6413 2447 6427
rect 2353 6393 2367 6407
rect 2413 6393 2427 6407
rect 2713 6413 2727 6427
rect 2333 6353 2347 6367
rect 2453 6393 2467 6407
rect 2473 6393 2487 6407
rect 2413 6353 2427 6367
rect 2353 6333 2367 6347
rect 2373 6333 2387 6347
rect 2293 6133 2307 6147
rect 2153 6113 2167 6127
rect 2173 6093 2187 6107
rect 2233 6113 2247 6127
rect 2073 6033 2087 6047
rect 2113 6033 2127 6047
rect 2013 5953 2027 5967
rect 1993 5933 2007 5947
rect 2053 5933 2067 5947
rect 1993 5893 2007 5907
rect 2073 5893 2087 5907
rect 1973 5873 1987 5887
rect 1953 5813 1967 5827
rect 2113 5893 2127 5907
rect 2093 5873 2107 5887
rect 2033 5833 2047 5847
rect 1993 5693 2007 5707
rect 2033 5693 2047 5707
rect 1993 5673 2007 5687
rect 1953 5633 1967 5647
rect 1973 5653 1987 5667
rect 2013 5653 2027 5667
rect 1993 5633 2007 5647
rect 1913 5593 1927 5607
rect 1993 5593 2007 5607
rect 1873 5553 1887 5567
rect 1853 5433 1867 5447
rect 1893 5453 1907 5467
rect 1993 5473 2007 5487
rect 1913 5433 1927 5447
rect 1953 5433 1967 5447
rect 1873 5413 1887 5427
rect 1853 5393 1867 5407
rect 1933 5393 1947 5407
rect 2093 5673 2107 5687
rect 2133 5673 2147 5687
rect 2133 5653 2147 5667
rect 2233 6073 2247 6087
rect 2213 6053 2227 6067
rect 2193 6033 2207 6047
rect 2193 5993 2207 6007
rect 2233 5953 2247 5967
rect 2273 6033 2287 6047
rect 2213 5933 2227 5947
rect 2253 5933 2267 5947
rect 2573 6393 2587 6407
rect 3113 6433 3127 6447
rect 3173 6433 3187 6447
rect 2953 6393 2967 6407
rect 2553 6353 2567 6367
rect 2633 6373 2647 6387
rect 2533 6313 2547 6327
rect 2533 6173 2547 6187
rect 2413 6133 2427 6147
rect 2313 6113 2327 6127
rect 2373 6093 2387 6107
rect 2293 5933 2307 5947
rect 2413 6053 2427 6067
rect 2433 6053 2447 6067
rect 2373 5993 2387 6007
rect 2333 5973 2347 5987
rect 2353 5953 2367 5967
rect 2213 5893 2227 5907
rect 2233 5893 2247 5907
rect 2253 5893 2267 5907
rect 2293 5893 2307 5907
rect 2313 5913 2327 5927
rect 2353 5913 2367 5927
rect 2333 5893 2347 5907
rect 2233 5813 2247 5827
rect 2173 5673 2187 5687
rect 2213 5673 2227 5687
rect 2173 5633 2187 5647
rect 2153 5613 2167 5627
rect 2193 5613 2207 5627
rect 2173 5593 2187 5607
rect 2273 5673 2287 5687
rect 2673 6373 2687 6387
rect 2713 6373 2727 6387
rect 2693 6353 2707 6367
rect 2733 6353 2747 6367
rect 2753 6373 2767 6387
rect 2793 6373 2807 6387
rect 2773 6353 2787 6367
rect 2633 6293 2647 6307
rect 2593 6153 2607 6167
rect 2773 6333 2787 6347
rect 2833 6353 2847 6367
rect 2853 6373 2867 6387
rect 2873 6353 2887 6367
rect 2893 6333 2907 6347
rect 2793 6313 2807 6327
rect 2653 6273 2667 6287
rect 2853 6273 2867 6287
rect 2693 6153 2707 6167
rect 2473 6113 2487 6127
rect 2513 6093 2527 6107
rect 2533 6113 2547 6127
rect 2633 6113 2647 6127
rect 2613 6093 2627 6107
rect 2733 6133 2747 6147
rect 2813 6133 2827 6147
rect 2973 6373 2987 6387
rect 2993 6393 3007 6407
rect 3033 6393 3047 6407
rect 3053 6393 3067 6407
rect 3013 6373 3027 6387
rect 3033 6373 3047 6387
rect 3073 6373 3087 6387
rect 2953 6353 2967 6367
rect 2913 6273 2927 6287
rect 2953 6173 2967 6187
rect 2893 6153 2907 6167
rect 2633 6073 2647 6087
rect 2653 6073 2667 6087
rect 2593 6053 2607 6067
rect 2753 6093 2767 6107
rect 2793 6093 2807 6107
rect 2913 6113 2927 6127
rect 2953 6113 2967 6127
rect 2713 6033 2727 6047
rect 2453 5933 2467 5947
rect 2513 5933 2527 5947
rect 2553 5933 2567 5947
rect 2613 5933 2627 5947
rect 2713 5933 2727 5947
rect 2773 5933 2787 5947
rect 2433 5873 2447 5887
rect 2473 5873 2487 5887
rect 2493 5893 2507 5907
rect 2573 5913 2587 5927
rect 2393 5853 2407 5867
rect 2593 5893 2607 5907
rect 2613 5893 2627 5907
rect 2553 5853 2567 5867
rect 2373 5833 2387 5847
rect 2393 5833 2407 5847
rect 2373 5713 2387 5727
rect 2233 5653 2247 5667
rect 2293 5653 2307 5667
rect 2353 5653 2367 5667
rect 2253 5613 2267 5627
rect 2593 5833 2607 5847
rect 2413 5673 2427 5687
rect 2433 5673 2447 5687
rect 2113 5573 2127 5587
rect 2213 5573 2227 5587
rect 2233 5573 2247 5587
rect 2073 5553 2087 5567
rect 2213 5513 2227 5527
rect 2073 5453 2087 5467
rect 2153 5453 2167 5467
rect 2033 5433 2047 5447
rect 2113 5413 2127 5427
rect 2173 5413 2187 5427
rect 1853 5373 1867 5387
rect 1813 5333 1827 5347
rect 1633 5133 1647 5147
rect 1673 5133 1687 5147
rect 1753 5133 1767 5147
rect 1713 5113 1727 5127
rect 1753 5113 1767 5127
rect 1613 4993 1627 5007
rect 1593 4973 1607 4987
rect 1653 4973 1667 4987
rect 1673 4973 1687 4987
rect 1613 4953 1627 4967
rect 1593 4933 1607 4947
rect 1613 4913 1627 4927
rect 1593 4893 1607 4907
rect 1573 4713 1587 4727
rect 1433 4673 1447 4687
rect 1453 4653 1467 4667
rect 1473 4653 1487 4667
rect 1493 4673 1507 4687
rect 1553 4673 1567 4687
rect 1533 4653 1547 4667
rect 1433 4633 1447 4647
rect 1553 4633 1567 4647
rect 1513 4613 1527 4627
rect 1573 4613 1587 4627
rect 1353 4493 1367 4507
rect 1413 4493 1427 4507
rect 1493 4493 1507 4507
rect 1273 4473 1287 4487
rect 1373 4473 1387 4487
rect 1393 4473 1407 4487
rect 1333 4433 1347 4447
rect 1353 4433 1367 4447
rect 1273 4253 1287 4267
rect 1113 4193 1127 4207
rect 1013 4173 1027 4187
rect 1073 4033 1087 4047
rect 1133 4173 1147 4187
rect 1273 4213 1287 4227
rect 1213 4153 1227 4167
rect 1453 4473 1467 4487
rect 1473 4433 1487 4447
rect 1513 4433 1527 4447
rect 1553 4453 1567 4467
rect 1453 4413 1467 4427
rect 1573 4413 1587 4427
rect 1453 4313 1467 4327
rect 1493 4313 1507 4327
rect 1313 4213 1327 4227
rect 1353 4213 1367 4227
rect 1253 4113 1267 4127
rect 1253 4053 1267 4067
rect 1133 4013 1147 4027
rect 1373 4193 1387 4207
rect 1553 4233 1567 4247
rect 1473 4213 1487 4227
rect 1613 4753 1627 4767
rect 1713 4933 1727 4947
rect 1733 4893 1747 4907
rect 1673 4853 1687 4867
rect 1633 4693 1647 4707
rect 1613 4653 1627 4667
rect 1633 4633 1647 4647
rect 1693 4733 1707 4747
rect 1733 4713 1747 4727
rect 2133 5393 2147 5407
rect 2153 5393 2167 5407
rect 2053 5353 2067 5367
rect 2193 5393 2207 5407
rect 2213 5393 2227 5407
rect 2213 5353 2227 5367
rect 1933 5333 1947 5347
rect 2173 5333 2187 5347
rect 2213 5333 2227 5347
rect 2193 5313 2207 5327
rect 1893 5173 1907 5187
rect 2013 5173 2027 5187
rect 2033 5173 2047 5187
rect 2073 5173 2087 5187
rect 1913 5133 1927 5147
rect 1933 5153 1947 5167
rect 1953 5133 1967 5147
rect 1993 5153 2007 5167
rect 2013 5133 2027 5147
rect 1933 5113 1947 5127
rect 1953 4993 1967 5007
rect 1933 4973 1947 4987
rect 1793 4953 1807 4967
rect 1773 4933 1787 4947
rect 1813 4933 1827 4947
rect 1833 4953 1847 4967
rect 1933 4953 1947 4967
rect 1993 5093 2007 5107
rect 2133 5173 2147 5187
rect 2053 5133 2067 5147
rect 2153 5153 2167 5167
rect 2173 5173 2187 5187
rect 2193 5153 2207 5167
rect 2113 5133 2127 5147
rect 2113 5113 2127 5127
rect 2033 5013 2047 5027
rect 2033 4993 2047 5007
rect 1973 4973 1987 4987
rect 1993 4973 2007 4987
rect 2253 5513 2267 5527
rect 2273 5473 2287 5487
rect 2353 5473 2367 5487
rect 2313 5453 2327 5467
rect 2373 5453 2387 5467
rect 2293 5413 2307 5427
rect 2333 5433 2347 5447
rect 2373 5433 2387 5447
rect 2353 5413 2367 5427
rect 2353 5353 2367 5367
rect 2673 5893 2687 5907
rect 2953 6093 2967 6107
rect 2833 6073 2847 6087
rect 2893 6073 2907 6087
rect 2933 6073 2947 6087
rect 2873 5933 2887 5947
rect 2813 5913 2827 5927
rect 3013 6133 3027 6147
rect 3253 6433 3267 6447
rect 3393 6433 3407 6447
rect 3133 6373 3147 6387
rect 3153 6373 3167 6387
rect 3153 6333 3167 6347
rect 3113 6293 3127 6307
rect 3193 6413 3207 6427
rect 3213 6413 3227 6427
rect 3233 6413 3247 6427
rect 3373 6413 3387 6427
rect 3193 6353 3207 6367
rect 3173 6273 3187 6287
rect 3233 6273 3247 6287
rect 3113 6253 3127 6267
rect 3133 6193 3147 6207
rect 3273 6373 3287 6387
rect 3293 6393 3307 6407
rect 3333 6393 3347 6407
rect 3353 6373 3367 6387
rect 3493 6413 3507 6427
rect 3533 6413 3547 6427
rect 3593 6413 3607 6427
rect 3713 6413 3727 6427
rect 3513 6373 3527 6387
rect 3253 6253 3267 6267
rect 3473 6313 3487 6327
rect 3493 6313 3507 6327
rect 3433 6273 3447 6287
rect 3253 6193 3267 6207
rect 3273 6193 3287 6207
rect 3173 6153 3187 6167
rect 3233 6153 3247 6167
rect 2953 6053 2967 6067
rect 2973 6053 2987 6067
rect 2933 5993 2947 6007
rect 2893 5913 2907 5927
rect 2913 5913 2927 5927
rect 2733 5893 2747 5907
rect 2693 5873 2707 5887
rect 2713 5873 2727 5887
rect 2633 5853 2647 5867
rect 2653 5853 2667 5867
rect 2753 5873 2767 5887
rect 2793 5893 2807 5907
rect 2793 5873 2807 5887
rect 2853 5873 2867 5887
rect 2893 5893 2907 5907
rect 2893 5873 2907 5887
rect 2873 5713 2887 5727
rect 2613 5693 2627 5707
rect 2673 5693 2687 5707
rect 2733 5693 2747 5707
rect 2813 5693 2827 5707
rect 2833 5693 2847 5707
rect 2473 5533 2487 5547
rect 2453 5493 2467 5507
rect 2433 5453 2447 5467
rect 2453 5453 2467 5467
rect 2573 5613 2587 5627
rect 2613 5593 2627 5607
rect 2533 5533 2547 5547
rect 2593 5533 2607 5547
rect 2493 5513 2507 5527
rect 2533 5453 2547 5467
rect 2653 5613 2667 5627
rect 2753 5633 2767 5647
rect 2773 5653 2787 5667
rect 2673 5593 2687 5607
rect 2633 5513 2647 5527
rect 2613 5473 2627 5487
rect 2653 5473 2667 5487
rect 2553 5413 2567 5427
rect 2593 5413 2607 5427
rect 2633 5433 2647 5447
rect 2393 5333 2407 5347
rect 2253 5193 2267 5207
rect 2293 5193 2307 5207
rect 2373 5193 2387 5207
rect 2733 5613 2747 5627
rect 2753 5513 2767 5527
rect 2733 5493 2747 5507
rect 2713 5393 2727 5407
rect 2513 5373 2527 5387
rect 2653 5373 2667 5387
rect 2633 5353 2647 5367
rect 2613 5233 2627 5247
rect 2233 5173 2247 5187
rect 2233 5153 2247 5167
rect 2413 5173 2427 5187
rect 2393 5153 2407 5167
rect 2493 5173 2507 5187
rect 2593 5173 2607 5187
rect 2453 5153 2467 5167
rect 2493 5153 2507 5167
rect 2353 5133 2367 5147
rect 2433 5133 2447 5147
rect 2493 5133 2507 5147
rect 2133 5033 2147 5047
rect 2213 5033 2227 5047
rect 1793 4913 1807 4927
rect 1873 4933 1887 4947
rect 1913 4933 1927 4947
rect 1893 4913 1907 4927
rect 1913 4893 1927 4907
rect 1893 4833 1907 4847
rect 1813 4793 1827 4807
rect 1853 4793 1867 4807
rect 1693 4673 1707 4687
rect 1713 4673 1727 4687
rect 1693 4633 1707 4647
rect 1653 4593 1667 4607
rect 1653 4513 1667 4527
rect 1613 4493 1627 4507
rect 1753 4653 1767 4667
rect 1813 4673 1827 4687
rect 1833 4653 1847 4667
rect 1853 4673 1867 4687
rect 1873 4653 1887 4667
rect 1793 4633 1807 4647
rect 1813 4633 1827 4647
rect 1733 4493 1747 4507
rect 1773 4613 1787 4627
rect 1873 4553 1887 4567
rect 1953 4933 1967 4947
rect 1993 4933 2007 4947
rect 2013 4953 2027 4967
rect 2073 4953 2087 4967
rect 1973 4913 1987 4927
rect 1953 4873 1967 4887
rect 1933 4813 1947 4827
rect 1933 4713 1947 4727
rect 1933 4673 1947 4687
rect 1973 4853 1987 4867
rect 1993 4833 2007 4847
rect 1833 4513 1847 4527
rect 1673 4253 1687 4267
rect 1693 4253 1707 4267
rect 1753 4253 1767 4267
rect 1613 4233 1627 4247
rect 1653 4233 1667 4247
rect 1633 4213 1647 4227
rect 1673 4213 1687 4227
rect 1513 4193 1527 4207
rect 1473 4173 1487 4187
rect 1493 4173 1507 4187
rect 1533 4173 1547 4187
rect 1593 4193 1607 4207
rect 1653 4193 1667 4207
rect 1313 4033 1327 4047
rect 1293 4013 1307 4027
rect 1073 3993 1087 4007
rect 1113 3993 1127 4007
rect 1133 3993 1147 4007
rect 1013 3953 1027 3967
rect 1033 3973 1047 3987
rect 1053 3953 1067 3967
rect 1093 3973 1107 3987
rect 1053 3933 1067 3947
rect 1073 3933 1087 3947
rect 1153 3953 1167 3967
rect 1173 3973 1187 3987
rect 1273 3973 1287 3987
rect 1353 3993 1367 4007
rect 1313 3953 1327 3967
rect 1133 3913 1147 3927
rect 1073 3813 1087 3827
rect 1113 3813 1127 3827
rect 1113 3733 1127 3747
rect 1073 3713 1087 3727
rect 1453 4033 1467 4047
rect 1433 4013 1447 4027
rect 1413 3893 1427 3907
rect 1193 3753 1207 3767
rect 1533 4153 1547 4167
rect 1573 4133 1587 4147
rect 1653 4153 1667 4167
rect 1773 4233 1787 4247
rect 1713 4213 1727 4227
rect 1753 4213 1767 4227
rect 1793 4193 1807 4207
rect 1813 4213 1827 4227
rect 1613 4113 1627 4127
rect 1613 4073 1627 4087
rect 1653 4033 1667 4047
rect 1593 3953 1607 3967
rect 1633 3953 1647 3967
rect 1533 3933 1547 3947
rect 1173 3733 1187 3747
rect 1153 3693 1167 3707
rect 1053 3633 1067 3647
rect 1093 3633 1107 3647
rect 1133 3633 1147 3647
rect 1033 3553 1047 3567
rect 1113 3553 1127 3567
rect 993 3473 1007 3487
rect 1153 3573 1167 3587
rect 1233 3733 1247 3747
rect 1313 3733 1327 3747
rect 1413 3733 1427 3747
rect 1313 3693 1327 3707
rect 1333 3693 1347 3707
rect 1353 3693 1367 3707
rect 1373 3713 1387 3727
rect 1213 3673 1227 3687
rect 1293 3673 1307 3687
rect 1393 3673 1407 3687
rect 1253 3653 1267 3667
rect 1293 3573 1307 3587
rect 1173 3553 1187 3567
rect 1193 3533 1207 3547
rect 1173 3513 1187 3527
rect 1233 3513 1247 3527
rect 1133 3493 1147 3507
rect 1053 3433 1067 3447
rect 1013 3313 1027 3327
rect 1113 3313 1127 3327
rect 973 3273 987 3287
rect 913 3253 927 3267
rect 953 3253 967 3267
rect 813 3213 827 3227
rect 873 3213 887 3227
rect 913 3213 927 3227
rect 953 3233 967 3247
rect 1053 3253 1067 3267
rect 1073 3213 1087 3227
rect 1253 3313 1267 3327
rect 1153 3213 1167 3227
rect 1193 3233 1207 3247
rect 1233 3233 1247 3247
rect 1213 3213 1227 3227
rect 893 3193 907 3207
rect 933 3193 947 3207
rect 973 3193 987 3207
rect 793 3173 807 3187
rect 773 3073 787 3087
rect 713 3033 727 3047
rect 1033 3153 1047 3167
rect 1173 3153 1187 3167
rect 1013 3133 1027 3147
rect 973 3073 987 3087
rect 1033 3073 1047 3087
rect 933 3053 947 3067
rect 973 3053 987 3067
rect 493 2993 507 3007
rect 513 2993 527 3007
rect 553 2993 567 3007
rect 573 3013 587 3027
rect 593 2993 607 3007
rect 673 3013 687 3027
rect 693 3013 707 3027
rect 653 2993 667 3007
rect 593 2973 607 2987
rect 673 2973 687 2987
rect 553 2773 567 2787
rect 513 2733 527 2747
rect 453 2713 467 2727
rect 273 2593 287 2607
rect 273 2573 287 2587
rect 313 2553 327 2567
rect 293 2493 307 2507
rect 293 2293 307 2307
rect 353 2553 367 2567
rect 353 2513 367 2527
rect 433 2573 447 2587
rect 493 2673 507 2687
rect 473 2553 487 2567
rect 793 2993 807 3007
rect 813 2973 827 2987
rect 853 2973 867 2987
rect 893 2993 907 3007
rect 993 3013 1007 3027
rect 1013 3033 1027 3047
rect 613 2953 627 2967
rect 693 2953 707 2967
rect 753 2953 767 2967
rect 613 2813 627 2827
rect 873 2953 887 2967
rect 853 2933 867 2947
rect 813 2813 827 2827
rect 593 2773 607 2787
rect 753 2793 767 2807
rect 793 2793 807 2807
rect 813 2793 827 2807
rect 853 2793 867 2807
rect 953 2953 967 2967
rect 993 2833 1007 2847
rect 653 2713 667 2727
rect 733 2753 747 2767
rect 613 2673 627 2687
rect 633 2593 647 2607
rect 593 2553 607 2567
rect 653 2533 667 2547
rect 553 2493 567 2507
rect 673 2513 687 2527
rect 693 2533 707 2547
rect 713 2493 727 2507
rect 893 2773 907 2787
rect 833 2733 847 2747
rect 933 2793 947 2807
rect 953 2793 967 2807
rect 973 2773 987 2787
rect 913 2733 927 2747
rect 973 2633 987 2647
rect 833 2593 847 2607
rect 953 2593 967 2607
rect 773 2513 787 2527
rect 793 2533 807 2547
rect 1153 3053 1167 3067
rect 1073 2973 1087 2987
rect 1053 2793 1067 2807
rect 1093 2793 1107 2807
rect 1033 2753 1047 2767
rect 1093 2753 1107 2767
rect 1113 2753 1127 2767
rect 1013 2733 1027 2747
rect 1073 2733 1087 2747
rect 993 2593 1007 2607
rect 1193 3033 1207 3047
rect 1213 2813 1227 2827
rect 1153 2733 1167 2747
rect 1173 2753 1187 2767
rect 1193 2733 1207 2747
rect 1233 2733 1247 2747
rect 1193 2713 1207 2727
rect 1133 2693 1147 2707
rect 1033 2573 1047 2587
rect 1013 2553 1027 2567
rect 1053 2553 1067 2567
rect 853 2513 867 2527
rect 993 2513 1007 2527
rect 1033 2513 1047 2527
rect 1153 2673 1167 2687
rect 1133 2573 1147 2587
rect 1173 2553 1187 2567
rect 973 2453 987 2467
rect 373 2333 387 2347
rect 613 2333 627 2347
rect 753 2333 767 2347
rect 373 2293 387 2307
rect 413 2293 427 2307
rect 513 2293 527 2307
rect 413 2273 427 2287
rect 273 2133 287 2147
rect 313 2133 327 2147
rect 313 2093 327 2107
rect 233 2033 247 2047
rect 193 2013 207 2027
rect 173 1993 187 2007
rect 153 1893 167 1907
rect 93 1833 107 1847
rect 213 1773 227 1787
rect 193 1753 207 1767
rect 13 1613 27 1627
rect 53 1613 67 1627
rect 93 1613 107 1627
rect 33 1593 47 1607
rect 73 1593 87 1607
rect 193 1613 207 1627
rect 173 1593 187 1607
rect 93 1573 107 1587
rect 113 1573 127 1587
rect 153 1573 167 1587
rect 153 1553 167 1567
rect 473 2253 487 2267
rect 513 2253 527 2267
rect 533 2253 547 2267
rect 613 2273 627 2287
rect 473 2233 487 2247
rect 493 2233 507 2247
rect 513 2233 527 2247
rect 393 2133 407 2147
rect 373 2093 387 2107
rect 353 2073 367 2087
rect 353 2053 367 2067
rect 333 2033 347 2047
rect 353 1993 367 2007
rect 293 1973 307 1987
rect 553 2213 567 2227
rect 493 2133 507 2147
rect 473 2113 487 2127
rect 393 2033 407 2047
rect 433 2033 447 2047
rect 453 2053 467 2067
rect 493 2073 507 2087
rect 513 2033 527 2047
rect 533 2033 547 2047
rect 393 1993 407 2007
rect 373 1953 387 1967
rect 393 1893 407 1907
rect 493 1953 507 1967
rect 653 2233 667 2247
rect 593 2173 607 2187
rect 573 2153 587 2167
rect 573 2133 587 2147
rect 593 2093 607 2107
rect 733 2253 747 2267
rect 713 2233 727 2247
rect 773 2273 787 2287
rect 793 2293 807 2307
rect 813 2253 827 2267
rect 833 2253 847 2267
rect 813 2233 827 2247
rect 753 2213 767 2227
rect 693 2173 707 2187
rect 613 2073 627 2087
rect 593 2053 607 2067
rect 633 2073 647 2087
rect 653 2053 667 2067
rect 713 2153 727 2167
rect 613 2033 627 2047
rect 593 1953 607 1967
rect 613 1933 627 1947
rect 493 1813 507 1827
rect 433 1793 447 1807
rect 313 1753 327 1767
rect 333 1753 347 1767
rect 453 1773 467 1787
rect 633 1833 647 1847
rect 593 1813 607 1827
rect 453 1753 467 1767
rect 733 2133 747 2147
rect 753 2093 767 2107
rect 733 2053 747 2067
rect 853 2173 867 2187
rect 833 2113 847 2127
rect 853 2093 867 2107
rect 813 2073 827 2087
rect 773 2053 787 2067
rect 813 2053 827 2067
rect 873 2073 887 2087
rect 853 2053 867 2067
rect 793 2033 807 2047
rect 833 2033 847 2047
rect 773 1973 787 1987
rect 753 1853 767 1867
rect 653 1793 667 1807
rect 373 1713 387 1727
rect 353 1653 367 1667
rect 393 1553 407 1567
rect 493 1693 507 1707
rect 453 1553 467 1567
rect 493 1633 507 1647
rect 493 1593 507 1607
rect 433 1513 447 1527
rect 273 1373 287 1387
rect 193 1353 207 1367
rect 233 1353 247 1367
rect 253 1353 267 1367
rect 293 1353 307 1367
rect 13 1333 27 1347
rect 53 1333 67 1347
rect 173 1333 187 1347
rect 13 1273 27 1287
rect 73 1273 87 1287
rect 33 853 47 867
rect 113 1273 127 1287
rect 133 1273 147 1287
rect 113 1133 127 1147
rect 93 1113 107 1127
rect 153 1113 167 1127
rect 213 1293 227 1307
rect 273 1293 287 1307
rect 193 1233 207 1247
rect 233 1093 247 1107
rect 413 1333 427 1347
rect 713 1813 727 1827
rect 833 1893 847 1907
rect 1033 2333 1047 2347
rect 993 2273 1007 2287
rect 973 2213 987 2227
rect 1113 2113 1127 2127
rect 1053 2093 1067 2107
rect 913 2073 927 2087
rect 953 2073 967 2087
rect 913 2033 927 2047
rect 1013 2073 1027 2087
rect 1033 2073 1047 2087
rect 1053 2053 1067 2067
rect 973 2033 987 2047
rect 893 1993 907 2007
rect 933 1993 947 2007
rect 993 1993 1007 2007
rect 973 1953 987 1967
rect 873 1913 887 1927
rect 853 1873 867 1887
rect 793 1833 807 1847
rect 733 1753 747 1767
rect 593 1713 607 1727
rect 753 1713 767 1727
rect 593 1673 607 1687
rect 573 1653 587 1667
rect 713 1633 727 1647
rect 573 1613 587 1627
rect 553 1573 567 1587
rect 593 1573 607 1587
rect 633 1573 647 1587
rect 613 1553 627 1567
rect 653 1513 667 1527
rect 533 1353 547 1367
rect 313 1293 327 1307
rect 393 1313 407 1327
rect 453 1313 467 1327
rect 413 1293 427 1307
rect 513 1333 527 1347
rect 533 1313 547 1327
rect 573 1313 587 1327
rect 613 1313 627 1327
rect 633 1293 647 1307
rect 313 1273 327 1287
rect 353 1273 367 1287
rect 373 1273 387 1287
rect 393 1273 407 1287
rect 473 1273 487 1287
rect 293 1253 307 1267
rect 293 1153 307 1167
rect 113 893 127 907
rect 33 813 47 827
rect 13 673 27 687
rect 93 693 107 707
rect 13 653 27 667
rect 53 653 67 667
rect 53 633 67 647
rect 13 613 27 627
rect 33 593 47 607
rect 133 873 147 887
rect 173 853 187 867
rect 333 1233 347 1247
rect 433 1233 447 1247
rect 333 1113 347 1127
rect 373 1153 387 1167
rect 393 1153 407 1167
rect 373 1113 387 1127
rect 313 873 327 887
rect 213 833 227 847
rect 213 773 227 787
rect 333 813 347 827
rect 293 793 307 807
rect 193 673 207 687
rect 113 633 127 647
rect 173 653 187 667
rect 413 1133 427 1147
rect 593 1253 607 1267
rect 633 1253 647 1267
rect 613 1173 627 1187
rect 473 1133 487 1147
rect 453 1113 467 1127
rect 433 893 447 907
rect 453 873 467 887
rect 773 1553 787 1567
rect 833 1853 847 1867
rect 1113 1973 1127 1987
rect 1053 1953 1067 1967
rect 1093 1953 1107 1967
rect 1013 1933 1027 1947
rect 1013 1893 1027 1907
rect 893 1813 907 1827
rect 933 1813 947 1827
rect 993 1813 1007 1827
rect 1013 1813 1027 1827
rect 953 1793 967 1807
rect 873 1733 887 1747
rect 793 1393 807 1407
rect 773 1333 787 1347
rect 733 1313 747 1327
rect 753 1293 767 1307
rect 793 1273 807 1287
rect 733 1253 747 1267
rect 773 1253 787 1267
rect 653 1233 667 1247
rect 713 1153 727 1167
rect 873 1353 887 1367
rect 913 1753 927 1767
rect 1033 1773 1047 1787
rect 1173 2373 1187 2387
rect 1233 2593 1247 2607
rect 1153 2173 1167 2187
rect 1273 3293 1287 3307
rect 1333 3553 1347 3567
rect 1373 3553 1387 3567
rect 1333 3493 1347 3507
rect 1493 3753 1507 3767
rect 1453 3733 1467 3747
rect 1513 3733 1527 3747
rect 1533 3713 1547 3727
rect 1533 3673 1547 3687
rect 1693 4133 1707 4147
rect 1793 4173 1807 4187
rect 1753 4153 1767 4167
rect 1733 4113 1747 4127
rect 1853 4493 1867 4507
rect 1893 4473 1907 4487
rect 1853 4433 1867 4447
rect 1933 4473 1947 4487
rect 1953 4473 1967 4487
rect 2093 4933 2107 4947
rect 2213 4993 2227 5007
rect 2233 4993 2247 5007
rect 2153 4973 2167 4987
rect 2453 5073 2467 5087
rect 2333 5013 2347 5027
rect 2373 4993 2387 5007
rect 2273 4973 2287 4987
rect 2353 4973 2367 4987
rect 2193 4953 2207 4967
rect 2133 4933 2147 4947
rect 2413 4973 2427 4987
rect 2433 4953 2447 4967
rect 2553 5133 2567 5147
rect 2673 5293 2687 5307
rect 2833 5613 2847 5627
rect 3113 6113 3127 6127
rect 3213 6133 3227 6147
rect 3193 6113 3207 6127
rect 3553 6393 3567 6407
rect 3633 6393 3647 6407
rect 3613 6373 3627 6387
rect 3573 6353 3587 6367
rect 3593 6353 3607 6367
rect 3673 6373 3687 6387
rect 3653 6353 3667 6367
rect 3753 6413 3767 6427
rect 4093 6433 4107 6447
rect 3733 6393 3747 6407
rect 3773 6393 3787 6407
rect 3753 6373 3767 6387
rect 3813 6393 3827 6407
rect 3833 6393 3847 6407
rect 3973 6413 3987 6427
rect 3773 6353 3787 6367
rect 3533 6333 3547 6347
rect 3593 6333 3607 6347
rect 3513 6173 3527 6187
rect 3813 6353 3827 6367
rect 3793 6333 3807 6347
rect 3773 6253 3787 6267
rect 3493 6153 3507 6167
rect 3513 6153 3527 6167
rect 3293 6133 3307 6147
rect 3373 6133 3387 6147
rect 3013 6073 3027 6087
rect 2973 5953 2987 5967
rect 2993 5953 3007 5967
rect 3033 6053 3047 6067
rect 3333 6113 3347 6127
rect 3113 6073 3127 6087
rect 3473 6133 3487 6147
rect 3573 6153 3587 6167
rect 3493 6113 3507 6127
rect 3133 6053 3147 6067
rect 3073 6033 3087 6047
rect 3093 5933 3107 5947
rect 3113 5933 3127 5947
rect 3013 5913 3027 5927
rect 3033 5913 3047 5927
rect 3073 5913 3087 5927
rect 3153 5913 3167 5927
rect 3173 5913 3187 5927
rect 2953 5873 2967 5887
rect 2993 5893 3007 5907
rect 3093 5873 3107 5887
rect 3133 5893 3147 5907
rect 3173 5893 3187 5907
rect 3053 5853 3067 5867
rect 3073 5853 3087 5867
rect 3153 5873 3167 5887
rect 3513 6093 3527 6107
rect 3453 6073 3467 6087
rect 3513 6073 3527 6087
rect 3313 6053 3327 6067
rect 3393 6013 3407 6027
rect 3593 6133 3607 6147
rect 3633 6133 3647 6147
rect 3713 6133 3727 6147
rect 3753 6133 3767 6147
rect 3593 6093 3607 6107
rect 3673 6113 3687 6127
rect 3733 6093 3747 6107
rect 3853 6333 3867 6347
rect 4013 6373 4027 6387
rect 4073 6373 4087 6387
rect 3913 6313 3927 6327
rect 3833 6273 3847 6287
rect 3813 6153 3827 6167
rect 4033 6333 4047 6347
rect 3893 6253 3907 6267
rect 3993 6253 4007 6267
rect 4673 6453 4687 6467
rect 4433 6433 4447 6447
rect 4553 6433 4567 6447
rect 4493 6393 4507 6407
rect 4633 6413 4647 6427
rect 4133 6353 4147 6367
rect 4193 6373 4207 6387
rect 4213 6353 4227 6367
rect 4293 6373 4307 6387
rect 4313 6353 4327 6367
rect 4373 6353 4387 6367
rect 4413 6353 4427 6367
rect 4473 6353 4487 6367
rect 4533 6373 4547 6387
rect 4573 6373 4587 6387
rect 4793 6433 4807 6447
rect 4693 6413 4707 6427
rect 4733 6413 4747 6427
rect 4753 6413 4767 6427
rect 4613 6373 4627 6387
rect 4633 6373 4647 6387
rect 4713 6373 4727 6387
rect 4513 6353 4527 6367
rect 4553 6353 4567 6367
rect 4573 6353 4587 6367
rect 4113 6333 4127 6347
rect 4173 6333 4187 6347
rect 4073 6293 4087 6307
rect 4053 6273 4067 6287
rect 4653 6353 4667 6367
rect 4713 6333 4727 6347
rect 4493 6313 4507 6327
rect 4613 6313 4627 6327
rect 4273 6253 4287 6267
rect 4173 6193 4187 6207
rect 4433 6193 4447 6207
rect 3793 6133 3807 6147
rect 3853 6133 3867 6147
rect 4033 6133 4047 6147
rect 4333 6153 4347 6167
rect 4373 6153 4387 6167
rect 4253 6133 4267 6147
rect 4293 6133 4307 6147
rect 3773 6093 3787 6107
rect 3793 6093 3807 6107
rect 3593 6073 3607 6087
rect 3613 6073 3627 6087
rect 3653 6073 3667 6087
rect 3753 6073 3767 6087
rect 3553 6053 3567 6067
rect 3533 6013 3547 6027
rect 3553 6013 3567 6027
rect 3373 5953 3387 5967
rect 3393 5933 3407 5947
rect 3413 5933 3427 5947
rect 3493 5933 3507 5947
rect 3273 5913 3287 5927
rect 3253 5893 3267 5907
rect 3293 5893 3307 5907
rect 3313 5913 3327 5927
rect 3333 5913 3347 5927
rect 3353 5893 3367 5907
rect 3393 5893 3407 5907
rect 3173 5853 3187 5867
rect 2953 5833 2967 5847
rect 3033 5833 3047 5847
rect 2853 5493 2867 5507
rect 3193 5833 3207 5847
rect 3293 5833 3307 5847
rect 3173 5793 3187 5807
rect 2973 5693 2987 5707
rect 3073 5693 3087 5707
rect 2993 5633 3007 5647
rect 3053 5653 3067 5667
rect 3053 5633 3067 5647
rect 3033 5613 3047 5627
rect 3093 5633 3107 5647
rect 3013 5593 3027 5607
rect 3453 5913 3467 5927
rect 3473 5873 3487 5887
rect 3433 5793 3447 5807
rect 3693 6013 3707 6027
rect 3673 5973 3687 5987
rect 3673 5933 3687 5947
rect 3573 5913 3587 5927
rect 3593 5893 3607 5907
rect 3613 5913 3627 5927
rect 3653 5913 3667 5927
rect 3713 5913 3727 5927
rect 3633 5893 3647 5907
rect 3613 5873 3627 5887
rect 3533 5853 3547 5867
rect 3113 5613 3127 5627
rect 3153 5613 3167 5627
rect 3073 5593 3087 5607
rect 3213 5633 3227 5647
rect 3253 5633 3267 5647
rect 3273 5633 3287 5647
rect 3313 5633 3327 5647
rect 3193 5593 3207 5607
rect 3173 5573 3187 5587
rect 3033 5553 3047 5567
rect 3113 5553 3127 5567
rect 2953 5533 2967 5547
rect 3033 5533 3047 5547
rect 3013 5513 3027 5527
rect 2953 5473 2967 5487
rect 2893 5453 2907 5467
rect 2973 5453 2987 5467
rect 2933 5433 2947 5447
rect 2813 5413 2827 5427
rect 2813 5393 2827 5407
rect 2873 5393 2887 5407
rect 2893 5413 2907 5427
rect 2853 5293 2867 5307
rect 2733 5233 2747 5247
rect 2693 5213 2707 5227
rect 2793 5213 2807 5227
rect 2673 5173 2687 5187
rect 2753 5193 2767 5207
rect 2753 5153 2767 5167
rect 2733 5133 2747 5147
rect 3033 5413 3047 5427
rect 3053 5433 3067 5447
rect 3073 5433 3087 5447
rect 3033 5393 3047 5407
rect 3193 5473 3207 5487
rect 3193 5453 3207 5467
rect 3233 5453 3247 5467
rect 3153 5433 3167 5447
rect 3213 5413 3227 5427
rect 3233 5433 3247 5447
rect 3373 5653 3387 5667
rect 3413 5653 3427 5667
rect 3353 5613 3367 5627
rect 3273 5593 3287 5607
rect 3333 5593 3347 5607
rect 3293 5573 3307 5587
rect 3473 5653 3487 5667
rect 3693 5893 3707 5907
rect 3713 5893 3727 5907
rect 3733 5893 3747 5907
rect 3773 5873 3787 5887
rect 3653 5853 3667 5867
rect 3673 5853 3687 5867
rect 3633 5833 3647 5847
rect 3553 5633 3567 5647
rect 3453 5613 3467 5627
rect 3493 5613 3507 5627
rect 3353 5533 3367 5547
rect 3413 5533 3427 5547
rect 3273 5433 3287 5447
rect 3313 5433 3327 5447
rect 3373 5473 3387 5487
rect 3433 5473 3447 5487
rect 3413 5453 3427 5467
rect 3353 5413 3367 5427
rect 3393 5433 3407 5447
rect 3613 5653 3627 5667
rect 3633 5653 3647 5667
rect 3573 5593 3587 5607
rect 3613 5613 3627 5627
rect 3853 6093 3867 6107
rect 3833 6013 3847 6027
rect 3873 6073 3887 6087
rect 3933 6013 3947 6027
rect 3853 5993 3867 6007
rect 3853 5953 3867 5967
rect 3893 5953 3907 5967
rect 3853 5913 3867 5927
rect 3873 5893 3887 5907
rect 3993 6113 4007 6127
rect 4053 6113 4067 6127
rect 4093 6093 4107 6107
rect 3993 6073 4007 6087
rect 3993 6033 4007 6047
rect 3993 6013 4007 6027
rect 3973 5973 3987 5987
rect 3953 5953 3967 5967
rect 4033 6073 4047 6087
rect 4053 6073 4067 6087
rect 3953 5933 3967 5947
rect 4013 5933 4027 5947
rect 3953 5913 3967 5927
rect 3973 5893 3987 5907
rect 4013 5893 4027 5907
rect 3933 5873 3947 5887
rect 3953 5853 3967 5867
rect 3933 5833 3947 5847
rect 3813 5813 3827 5827
rect 3933 5733 3947 5747
rect 3733 5653 3747 5667
rect 3773 5653 3787 5667
rect 3673 5613 3687 5627
rect 3713 5613 3727 5627
rect 3793 5613 3807 5627
rect 3613 5593 3627 5607
rect 3693 5593 3707 5607
rect 3733 5593 3747 5607
rect 3593 5573 3607 5587
rect 3473 5473 3487 5487
rect 3573 5453 3587 5467
rect 3653 5553 3667 5567
rect 3713 5553 3727 5567
rect 3673 5533 3687 5547
rect 3633 5473 3647 5487
rect 3493 5433 3507 5447
rect 3453 5413 3467 5427
rect 3533 5413 3547 5427
rect 3333 5393 3347 5407
rect 3513 5393 3527 5407
rect 3033 5293 3047 5307
rect 2913 5193 2927 5207
rect 2573 5113 2587 5127
rect 2613 5113 2627 5127
rect 2753 5113 2767 5127
rect 2773 5113 2787 5127
rect 2793 5113 2807 5127
rect 2533 5093 2547 5107
rect 2733 5093 2747 5107
rect 2673 5013 2687 5027
rect 2593 4993 2607 5007
rect 2633 4973 2647 4987
rect 2413 4933 2427 4947
rect 2253 4913 2267 4927
rect 2293 4913 2307 4927
rect 2493 4893 2507 4907
rect 2533 4873 2547 4887
rect 2493 4833 2507 4847
rect 2873 5173 2887 5187
rect 2833 5133 2847 5147
rect 2853 5113 2867 5127
rect 2833 5093 2847 5107
rect 2813 5073 2827 5087
rect 2933 5153 2947 5167
rect 2953 5173 2967 5187
rect 3013 5153 3027 5167
rect 2993 5133 3007 5147
rect 2993 5113 3007 5127
rect 3013 5113 3027 5127
rect 2973 5093 2987 5107
rect 2753 5053 2767 5067
rect 2853 5053 2867 5067
rect 2893 5053 2907 5067
rect 2953 5053 2967 5067
rect 2693 4953 2707 4967
rect 2673 4933 2687 4947
rect 2713 4933 2727 4947
rect 2793 4993 2807 5007
rect 2813 4973 2827 4987
rect 2953 5013 2967 5027
rect 2933 4993 2947 5007
rect 2893 4973 2907 4987
rect 2933 4973 2947 4987
rect 2753 4933 2767 4947
rect 2773 4933 2787 4947
rect 2813 4953 2827 4967
rect 2833 4933 2847 4947
rect 2873 4933 2887 4947
rect 2613 4913 2627 4927
rect 2773 4913 2787 4927
rect 3413 5353 3427 5367
rect 3173 5333 3187 5347
rect 3093 5273 3107 5287
rect 3253 5253 3267 5267
rect 3173 5213 3187 5227
rect 3133 5193 3147 5207
rect 3093 5173 3107 5187
rect 3113 5173 3127 5187
rect 3173 5173 3187 5187
rect 3133 5153 3147 5167
rect 3193 5153 3207 5167
rect 3213 5173 3227 5187
rect 3233 5173 3247 5187
rect 3113 5133 3127 5147
rect 3053 5073 3067 5087
rect 3213 5093 3227 5107
rect 2993 5033 3007 5047
rect 3093 5033 3107 5047
rect 3113 5033 3127 5047
rect 2973 4973 2987 4987
rect 3033 4993 3047 5007
rect 2913 4933 2927 4947
rect 2973 4933 2987 4947
rect 3013 4953 3027 4967
rect 2893 4913 2907 4927
rect 3193 5013 3207 5027
rect 3153 4973 3167 4987
rect 3173 4973 3187 4987
rect 3053 4953 3067 4967
rect 3073 4933 3087 4947
rect 3133 4953 3147 4967
rect 3113 4933 3127 4947
rect 2913 4893 2927 4907
rect 3013 4893 3027 4907
rect 2093 4753 2107 4767
rect 2233 4733 2247 4747
rect 2433 4733 2447 4747
rect 2393 4713 2407 4727
rect 2413 4713 2427 4727
rect 2193 4693 2207 4707
rect 2213 4673 2227 4687
rect 2253 4693 2267 4707
rect 2353 4693 2367 4707
rect 2293 4673 2307 4687
rect 2373 4673 2387 4687
rect 2313 4653 2327 4667
rect 2513 4713 2527 4727
rect 2433 4693 2447 4707
rect 2293 4633 2307 4647
rect 2333 4633 2347 4647
rect 2373 4633 2387 4647
rect 2313 4613 2327 4627
rect 2453 4633 2467 4647
rect 2453 4613 2467 4627
rect 2293 4573 2307 4587
rect 2353 4573 2367 4587
rect 2373 4573 2387 4587
rect 2433 4573 2447 4587
rect 2053 4513 2067 4527
rect 2033 4493 2047 4507
rect 2073 4473 2087 4487
rect 1953 4433 1967 4447
rect 2193 4513 2207 4527
rect 2153 4493 2167 4507
rect 2173 4493 2187 4507
rect 1873 4213 1887 4227
rect 1833 4033 1847 4047
rect 1713 4013 1727 4027
rect 1753 4013 1767 4027
rect 1753 3973 1767 3987
rect 1773 3953 1787 3967
rect 1833 3953 1847 3967
rect 1733 3933 1747 3947
rect 1573 3653 1587 3667
rect 1493 3633 1507 3647
rect 1593 3633 1607 3647
rect 1473 3593 1487 3607
rect 1433 3533 1447 3547
rect 1433 3513 1447 3527
rect 1373 3293 1387 3307
rect 1293 3233 1307 3247
rect 1293 3133 1307 3147
rect 1333 3133 1347 3147
rect 1293 3093 1307 3107
rect 1333 3033 1347 3047
rect 1393 3013 1407 3027
rect 1353 2993 1367 3007
rect 1393 2993 1407 3007
rect 1333 2973 1347 2987
rect 1313 2773 1327 2787
rect 1373 2813 1387 2827
rect 1273 2753 1287 2767
rect 1293 2733 1307 2747
rect 1333 2753 1347 2767
rect 1353 2753 1367 2767
rect 1393 2753 1407 2767
rect 1373 2733 1387 2747
rect 1413 2713 1427 2727
rect 1333 2653 1347 2667
rect 1373 2593 1387 2607
rect 1513 3513 1527 3527
rect 1553 3513 1567 3527
rect 1513 3473 1527 3487
rect 1673 3653 1687 3667
rect 1833 3773 1847 3787
rect 1733 3693 1747 3707
rect 1773 3693 1787 3707
rect 1673 3633 1687 3647
rect 1633 3533 1647 3547
rect 1613 3513 1627 3527
rect 1673 3513 1687 3527
rect 1833 3693 1847 3707
rect 1813 3673 1827 3687
rect 1833 3673 1847 3687
rect 1793 3613 1807 3627
rect 1733 3533 1747 3547
rect 1733 3493 1747 3507
rect 1813 3513 1827 3527
rect 1493 3213 1507 3227
rect 1513 3213 1527 3227
rect 1773 3293 1787 3307
rect 1593 3233 1607 3247
rect 1513 3073 1527 3087
rect 1453 3053 1467 3067
rect 1473 3053 1487 3067
rect 1533 3053 1547 3067
rect 1613 3213 1627 3227
rect 1693 3253 1707 3267
rect 1733 3233 1747 3247
rect 1773 3233 1787 3247
rect 1653 3193 1667 3207
rect 1713 3193 1727 3207
rect 1753 3193 1767 3207
rect 1813 3473 1827 3487
rect 1993 4173 2007 4187
rect 1953 4153 1967 4167
rect 2013 4133 2027 4147
rect 2093 4213 2107 4227
rect 2113 4193 2127 4207
rect 2393 4513 2407 4527
rect 2593 4673 2607 4687
rect 2633 4673 2647 4687
rect 2573 4653 2587 4667
rect 2533 4633 2547 4647
rect 2593 4633 2607 4647
rect 2813 4653 2827 4667
rect 2653 4593 2667 4607
rect 2313 4453 2327 4467
rect 2513 4513 2527 4527
rect 2573 4513 2587 4527
rect 2433 4473 2447 4487
rect 2493 4453 2507 4467
rect 2533 4453 2547 4467
rect 2713 4493 2727 4507
rect 2693 4413 2707 4427
rect 2793 4633 2807 4647
rect 2773 4413 2787 4427
rect 2193 4193 2207 4207
rect 2213 4173 2227 4187
rect 2233 4193 2247 4207
rect 2173 4153 2187 4167
rect 2113 4133 2127 4147
rect 2153 4133 2167 4147
rect 2213 4133 2227 4147
rect 2253 4133 2267 4147
rect 2673 4253 2687 4267
rect 2733 4253 2747 4267
rect 2353 4173 2367 4187
rect 2393 4153 2407 4167
rect 2993 4713 3007 4727
rect 2893 4673 2907 4687
rect 2953 4653 2967 4667
rect 2973 4533 2987 4547
rect 2853 4493 2867 4507
rect 2813 4473 2827 4487
rect 2873 4453 2887 4467
rect 2933 4453 2947 4467
rect 3353 5193 3367 5207
rect 3273 5173 3287 5187
rect 3293 5153 3307 5167
rect 3333 5153 3347 5167
rect 3313 5073 3327 5087
rect 3373 5173 3387 5187
rect 3353 5113 3367 5127
rect 3393 5113 3407 5127
rect 3533 5253 3547 5267
rect 3513 5233 3527 5247
rect 3453 5193 3467 5207
rect 3433 5133 3447 5147
rect 3493 5153 3507 5167
rect 3453 5113 3467 5127
rect 3533 5173 3547 5187
rect 3653 5433 3667 5447
rect 3653 5413 3667 5427
rect 3593 5373 3607 5387
rect 3873 5633 3887 5647
rect 4013 5793 4027 5807
rect 3973 5753 3987 5767
rect 3893 5613 3907 5627
rect 3953 5613 3967 5627
rect 3813 5573 3827 5587
rect 3793 5533 3807 5547
rect 3933 5533 3947 5547
rect 3993 5533 4007 5547
rect 3913 5513 3927 5527
rect 3693 5433 3707 5447
rect 3833 5453 3847 5467
rect 3853 5453 3867 5467
rect 3733 5433 3747 5447
rect 3753 5433 3767 5447
rect 3813 5413 3827 5427
rect 3873 5433 3887 5447
rect 3893 5433 3907 5447
rect 4073 6053 4087 6067
rect 4173 6113 4187 6127
rect 4113 6073 4127 6087
rect 4113 6053 4127 6067
rect 4093 6033 4107 6047
rect 4053 5973 4067 5987
rect 4073 5973 4087 5987
rect 4193 6093 4207 6107
rect 4233 6113 4247 6127
rect 4153 6073 4167 6087
rect 4313 6113 4327 6127
rect 4253 6093 4267 6107
rect 4313 6093 4327 6107
rect 4353 6093 4367 6107
rect 4133 6013 4147 6027
rect 4213 6053 4227 6067
rect 4173 6033 4187 6047
rect 4153 5933 4167 5947
rect 4193 5933 4207 5947
rect 4073 5893 4087 5907
rect 4113 5893 4127 5907
rect 4153 5913 4167 5927
rect 4253 5913 4267 5927
rect 4193 5893 4207 5907
rect 4233 5893 4247 5907
rect 4133 5873 4147 5887
rect 4173 5873 4187 5887
rect 4113 5853 4127 5867
rect 4053 5813 4067 5827
rect 4093 5753 4107 5767
rect 4053 5713 4067 5727
rect 4033 5673 4047 5687
rect 4153 5773 4167 5787
rect 4133 5693 4147 5707
rect 4113 5653 4127 5667
rect 4273 5893 4287 5907
rect 4253 5873 4267 5887
rect 4273 5853 4287 5867
rect 4213 5793 4227 5807
rect 4253 5773 4267 5787
rect 4233 5673 4247 5687
rect 4193 5653 4207 5667
rect 4293 5833 4307 5847
rect 4273 5713 4287 5727
rect 4413 6073 4427 6087
rect 4453 6173 4467 6187
rect 4593 6293 4607 6307
rect 4513 6193 4527 6207
rect 4553 6193 4567 6207
rect 4493 6133 4507 6147
rect 4553 6153 4567 6167
rect 4493 6093 4507 6107
rect 4713 6253 4727 6267
rect 4633 6213 4647 6227
rect 4593 6133 4607 6147
rect 4753 6373 4767 6387
rect 4773 6393 4787 6407
rect 5113 6473 5127 6487
rect 5153 6473 5167 6487
rect 4913 6453 4927 6467
rect 5013 6453 5027 6467
rect 4813 6393 4827 6407
rect 4793 6373 4807 6387
rect 4853 6393 4867 6407
rect 4893 6373 4907 6387
rect 4933 6433 4947 6447
rect 4953 6413 4967 6427
rect 5053 6393 5067 6407
rect 4993 6353 5007 6367
rect 4993 6313 5007 6327
rect 5013 6313 5027 6327
rect 4973 6293 4987 6307
rect 4893 6273 4907 6287
rect 4753 6213 4767 6227
rect 4733 6153 4747 6167
rect 4573 6093 4587 6107
rect 4593 6113 4607 6127
rect 4673 6113 4687 6127
rect 4733 6133 4747 6147
rect 4653 6093 4667 6107
rect 4613 6073 4627 6087
rect 4673 6073 4687 6087
rect 4433 6053 4447 6067
rect 4433 6013 4447 6027
rect 4453 5953 4467 5967
rect 4553 5933 4567 5947
rect 4373 5913 4387 5927
rect 4433 5913 4447 5927
rect 4353 5893 4367 5907
rect 4393 5893 4407 5907
rect 4353 5853 4367 5867
rect 4353 5773 4367 5787
rect 4473 5893 4487 5907
rect 4493 5913 4507 5927
rect 4453 5873 4467 5887
rect 4413 5853 4427 5867
rect 4393 5793 4407 5807
rect 4373 5753 4387 5767
rect 4373 5733 4387 5747
rect 4453 5733 4467 5747
rect 4333 5693 4347 5707
rect 4313 5673 4327 5687
rect 4173 5613 4187 5627
rect 4193 5633 4207 5647
rect 4233 5633 4247 5647
rect 4293 5653 4307 5667
rect 4353 5653 4367 5667
rect 4033 5593 4047 5607
rect 4033 5573 4047 5587
rect 4153 5593 4167 5607
rect 4073 5553 4087 5567
rect 3953 5453 3967 5467
rect 4013 5453 4027 5467
rect 4033 5453 4047 5467
rect 4113 5453 4127 5467
rect 3853 5413 3867 5427
rect 3813 5393 3827 5407
rect 3773 5373 3787 5387
rect 3673 5313 3687 5327
rect 3613 5253 3627 5267
rect 3653 5253 3667 5267
rect 3593 5173 3607 5187
rect 3633 5233 3647 5247
rect 3653 5213 3667 5227
rect 3633 5173 3647 5187
rect 3553 5153 3567 5167
rect 3533 5133 3547 5147
rect 3573 5133 3587 5147
rect 3653 5153 3667 5167
rect 3433 5093 3447 5107
rect 3373 5073 3387 5087
rect 3313 5053 3327 5067
rect 3333 5053 3347 5067
rect 3273 5033 3287 5047
rect 3253 4953 3267 4967
rect 3273 4953 3287 4967
rect 3173 4913 3187 4927
rect 3193 4913 3207 4927
rect 3233 4913 3247 4927
rect 3273 4913 3287 4927
rect 3293 4933 3307 4947
rect 3433 5033 3447 5047
rect 3413 4973 3427 4987
rect 3353 4933 3367 4947
rect 3393 4933 3407 4947
rect 3433 4933 3447 4947
rect 3333 4913 3347 4927
rect 3093 4653 3107 4667
rect 3153 4653 3167 4667
rect 3073 4593 3087 4607
rect 3113 4633 3127 4647
rect 3273 4693 3287 4707
rect 3313 4693 3327 4707
rect 3393 4653 3407 4667
rect 3353 4633 3367 4647
rect 3013 4453 3027 4467
rect 3053 4473 3067 4487
rect 3013 4433 3027 4447
rect 2833 4313 2847 4327
rect 2913 4313 2927 4327
rect 3293 4473 3307 4487
rect 3133 4393 3147 4407
rect 3253 4413 3267 4427
rect 3273 4413 3287 4427
rect 2473 4173 2487 4187
rect 2533 4173 2547 4187
rect 1913 4013 1927 4027
rect 1953 3993 1967 4007
rect 2053 3953 2067 3967
rect 2073 3973 2087 3987
rect 2533 4133 2547 4147
rect 2713 4173 2727 4187
rect 2593 4133 2607 4147
rect 2573 4073 2587 4087
rect 2573 4033 2587 4047
rect 2633 4033 2647 4047
rect 2173 3993 2187 4007
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 2333 3993 2347 4007
rect 2373 3993 2387 4007
rect 2273 3973 2287 3987
rect 2313 3953 2327 3967
rect 2413 3973 2427 3987
rect 2253 3933 2267 3947
rect 2553 4013 2567 4027
rect 2593 4013 2607 4027
rect 2613 4013 2627 4027
rect 2493 3993 2507 4007
rect 2473 3973 2487 3987
rect 2513 3973 2527 3987
rect 2533 3993 2547 4007
rect 2613 3973 2627 3987
rect 2413 3933 2427 3947
rect 2453 3933 2467 3947
rect 2293 3833 2307 3847
rect 1913 3753 1927 3767
rect 1973 3753 1987 3767
rect 1893 3733 1907 3747
rect 1893 3693 1907 3707
rect 1873 3673 1887 3687
rect 1873 3653 1887 3667
rect 1853 3513 1867 3527
rect 1833 3273 1847 3287
rect 1933 3733 1947 3747
rect 1913 3593 1927 3607
rect 2093 3733 2107 3747
rect 2133 3733 2147 3747
rect 2033 3693 2047 3707
rect 2053 3693 2067 3707
rect 2133 3693 2147 3707
rect 2293 3773 2307 3787
rect 2393 3773 2407 3787
rect 2373 3753 2387 3767
rect 2573 3793 2587 3807
rect 2773 4193 2787 4207
rect 2793 4213 2807 4227
rect 2813 4193 2827 4207
rect 2853 4193 2867 4207
rect 2753 4173 2767 4187
rect 2773 4173 2787 4187
rect 2693 4153 2707 4167
rect 2733 4153 2747 4167
rect 2713 4073 2727 4087
rect 2673 4013 2687 4027
rect 2693 3993 2707 4007
rect 2733 3973 2747 3987
rect 2713 3933 2727 3947
rect 2633 3833 2647 3847
rect 2633 3813 2647 3827
rect 2613 3753 2627 3767
rect 2193 3693 2207 3707
rect 2153 3673 2167 3687
rect 1993 3593 2007 3607
rect 1913 3573 1927 3587
rect 1953 3573 1967 3587
rect 1933 3553 1947 3567
rect 1893 3493 1907 3507
rect 1973 3553 1987 3567
rect 2073 3633 2087 3647
rect 2053 3553 2067 3567
rect 2093 3553 2107 3567
rect 1993 3493 2007 3507
rect 2073 3513 2087 3527
rect 2173 3613 2187 3627
rect 2293 3713 2307 3727
rect 2393 3713 2407 3727
rect 2413 3713 2427 3727
rect 2213 3673 2227 3687
rect 2273 3673 2287 3687
rect 2293 3673 2307 3687
rect 2233 3613 2247 3627
rect 2133 3493 2147 3507
rect 1813 3253 1827 3267
rect 1853 3253 1867 3267
rect 2093 3473 2107 3487
rect 2213 3473 2227 3487
rect 2353 3673 2367 3687
rect 2393 3673 2407 3687
rect 2513 3713 2527 3727
rect 2573 3713 2587 3727
rect 2613 3713 2627 3727
rect 2893 4193 2907 4207
rect 2913 4173 2927 4187
rect 3053 4193 3067 4207
rect 3093 4193 3107 4207
rect 2873 4153 2887 4167
rect 2913 4153 2927 4167
rect 3013 4153 3027 4167
rect 2933 4113 2947 4127
rect 2933 4053 2947 4067
rect 2973 4053 2987 4067
rect 2913 4033 2927 4047
rect 2813 4013 2827 4027
rect 2953 4013 2967 4027
rect 2773 3973 2787 3987
rect 2793 3953 2807 3967
rect 2853 3953 2867 3967
rect 2873 3973 2887 3987
rect 2993 4033 3007 4047
rect 3013 4013 3027 4027
rect 3093 4013 3107 4027
rect 3013 3973 3027 3987
rect 3033 3993 3047 4007
rect 3473 5073 3487 5087
rect 3553 5053 3567 5067
rect 3493 4953 3507 4967
rect 3553 4953 3567 4967
rect 3533 4933 3547 4947
rect 3653 5033 3667 5047
rect 3593 4953 3607 4967
rect 3573 4773 3587 4787
rect 3493 4673 3507 4687
rect 3373 4513 3387 4527
rect 3453 4513 3467 4527
rect 3393 4493 3407 4507
rect 3493 4493 3507 4507
rect 3373 4453 3387 4467
rect 3413 4453 3427 4467
rect 3433 4473 3447 4487
rect 3453 4453 3467 4467
rect 3473 4453 3487 4467
rect 3433 4433 3447 4447
rect 3353 4413 3367 4427
rect 3393 4333 3407 4347
rect 3273 4153 3287 4167
rect 3413 4253 3427 4267
rect 3413 4213 3427 4227
rect 3433 4213 3447 4227
rect 3373 4173 3387 4187
rect 3433 4193 3447 4207
rect 3453 4173 3467 4187
rect 3533 4653 3547 4667
rect 3553 4673 3567 4687
rect 3573 4633 3587 4647
rect 3573 4493 3587 4507
rect 3533 4473 3547 4487
rect 3513 4453 3527 4467
rect 3493 4333 3507 4347
rect 3693 5193 3707 5207
rect 3713 5133 3727 5147
rect 3733 5133 3747 5147
rect 3753 5153 3767 5167
rect 3813 5153 3827 5167
rect 3693 5113 3707 5127
rect 3773 5093 3787 5107
rect 3753 4973 3767 4987
rect 3653 4933 3667 4947
rect 3693 4933 3707 4947
rect 3713 4953 3727 4967
rect 3733 4933 3747 4947
rect 3653 4913 3667 4927
rect 3713 4913 3727 4927
rect 3633 4893 3647 4907
rect 3653 4853 3667 4867
rect 3733 4793 3747 4807
rect 3633 4693 3647 4707
rect 3753 4753 3767 4767
rect 3833 5133 3847 5147
rect 3813 5113 3827 5127
rect 3793 5073 3807 5087
rect 3813 5053 3827 5067
rect 3913 5413 3927 5427
rect 3953 5433 3967 5447
rect 3993 5433 4007 5447
rect 4013 5433 4027 5447
rect 3893 5393 3907 5407
rect 3873 5293 3887 5307
rect 4033 5393 4047 5407
rect 4053 5393 4067 5407
rect 4093 5413 4107 5427
rect 4113 5413 4127 5427
rect 4193 5573 4207 5587
rect 4293 5613 4307 5627
rect 4273 5573 4287 5587
rect 4233 5553 4247 5567
rect 4213 5513 4227 5527
rect 4273 5513 4287 5527
rect 4233 5453 4247 5467
rect 4113 5393 4127 5407
rect 3973 5373 3987 5387
rect 3953 5333 3967 5347
rect 4013 5333 4027 5347
rect 4033 5293 4047 5307
rect 4013 5253 4027 5267
rect 4013 5233 4027 5247
rect 3953 5213 3967 5227
rect 3893 5153 3907 5167
rect 3933 5173 3947 5187
rect 3853 5073 3867 5087
rect 3833 4993 3847 5007
rect 3833 4973 3847 4987
rect 3813 4933 3827 4947
rect 3853 4933 3867 4947
rect 3813 4913 3827 4927
rect 3813 4833 3827 4847
rect 3853 4873 3867 4887
rect 3853 4833 3867 4847
rect 3833 4813 3847 4827
rect 3833 4793 3847 4807
rect 3613 4653 3627 4667
rect 3693 4673 3707 4687
rect 3653 4653 3667 4667
rect 3773 4693 3787 4707
rect 3753 4673 3767 4687
rect 3753 4653 3767 4667
rect 3793 4673 3807 4687
rect 3893 5053 3907 5067
rect 4073 5373 4087 5387
rect 4093 5353 4107 5367
rect 4113 5253 4127 5267
rect 3973 5173 3987 5187
rect 4013 5173 4027 5187
rect 4033 5173 4047 5187
rect 4053 5173 4067 5187
rect 3993 5133 4007 5147
rect 4013 5133 4027 5147
rect 4033 5133 4047 5147
rect 4053 5153 4067 5167
rect 4093 5153 4107 5167
rect 4073 5133 4087 5147
rect 3953 5093 3967 5107
rect 3933 5013 3947 5027
rect 3913 4993 3927 5007
rect 3933 4973 3947 4987
rect 3913 4953 3927 4967
rect 3893 4913 3907 4927
rect 3993 5053 4007 5067
rect 4093 5113 4107 5127
rect 4033 5053 4047 5067
rect 4093 5033 4107 5047
rect 4073 4993 4087 5007
rect 3993 4973 4007 4987
rect 4013 4973 4027 4987
rect 3953 4953 3967 4967
rect 3953 4933 3967 4947
rect 4113 4993 4127 5007
rect 4033 4933 4047 4947
rect 4053 4933 4067 4947
rect 4073 4933 4087 4947
rect 3993 4913 4007 4927
rect 3973 4853 3987 4867
rect 3873 4793 3887 4807
rect 3933 4793 3947 4807
rect 3993 4793 4007 4807
rect 3853 4753 3867 4767
rect 3853 4673 3867 4687
rect 3593 4413 3607 4427
rect 3673 4473 3687 4487
rect 3593 4373 3607 4387
rect 3553 4353 3567 4367
rect 3573 4253 3587 4267
rect 3513 4233 3527 4247
rect 3513 4193 3527 4207
rect 3413 4153 3427 4167
rect 3453 4153 3467 4167
rect 3153 4113 3167 4127
rect 3393 4113 3407 4127
rect 3173 4033 3187 4047
rect 3213 4033 3227 4047
rect 3133 3993 3147 4007
rect 3053 3973 3067 3987
rect 3113 3973 3127 3987
rect 3193 3993 3207 4007
rect 2893 3953 2907 3967
rect 2973 3953 2987 3967
rect 3033 3953 3047 3967
rect 3273 3993 3287 4007
rect 2753 3913 2767 3927
rect 2893 3813 2907 3827
rect 2753 3793 2767 3807
rect 2873 3793 2887 3807
rect 2673 3733 2687 3747
rect 2593 3693 2607 3707
rect 2253 3513 2267 3527
rect 2293 3513 2307 3527
rect 2373 3513 2387 3527
rect 2353 3473 2367 3487
rect 2533 3613 2547 3627
rect 2613 3633 2627 3647
rect 2433 3533 2447 3547
rect 2493 3533 2507 3547
rect 2433 3493 2447 3507
rect 2393 3393 2407 3407
rect 2273 3333 2287 3347
rect 2233 3313 2247 3327
rect 1853 3233 1867 3247
rect 1893 3233 1907 3247
rect 1913 3233 1927 3247
rect 1813 3213 1827 3227
rect 1833 3213 1847 3227
rect 1793 3153 1807 3167
rect 1753 3093 1767 3107
rect 1713 3073 1727 3087
rect 1653 3053 1667 3067
rect 1773 3073 1787 3087
rect 1693 3033 1707 3047
rect 1633 3013 1647 3027
rect 1733 3013 1747 3027
rect 1833 3053 1847 3067
rect 1793 3033 1807 3047
rect 1773 3013 1787 3027
rect 1833 3033 1847 3047
rect 1773 2913 1787 2927
rect 1613 2793 1627 2807
rect 1673 2793 1687 2807
rect 1593 2773 1607 2787
rect 1453 2753 1467 2767
rect 1473 2733 1487 2747
rect 1493 2753 1507 2767
rect 1553 2753 1567 2767
rect 1533 2733 1547 2747
rect 1653 2773 1667 2787
rect 1453 2713 1467 2727
rect 1493 2713 1507 2727
rect 1273 2553 1287 2567
rect 1353 2553 1367 2567
rect 1493 2593 1507 2607
rect 1313 2533 1327 2547
rect 1433 2573 1447 2587
rect 1333 2513 1347 2527
rect 1453 2533 1467 2547
rect 1593 2733 1607 2747
rect 1533 2713 1547 2727
rect 1553 2713 1567 2727
rect 1593 2713 1607 2727
rect 1533 2613 1547 2627
rect 1513 2573 1527 2587
rect 1593 2653 1607 2667
rect 1573 2633 1587 2647
rect 1553 2573 1567 2587
rect 1753 2773 1767 2787
rect 1713 2713 1727 2727
rect 1913 3153 1927 3167
rect 1873 3073 1887 3087
rect 1993 3093 2007 3107
rect 1953 3053 1967 3067
rect 2193 3253 2207 3267
rect 2233 3253 2247 3267
rect 2353 3213 2367 3227
rect 2313 3173 2327 3187
rect 2253 3073 2267 3087
rect 2093 3053 2107 3067
rect 2113 3053 2127 3067
rect 2233 3053 2247 3067
rect 2273 3053 2287 3067
rect 2293 3053 2307 3067
rect 1933 3033 1947 3047
rect 1913 3013 1927 3027
rect 1973 3013 1987 3027
rect 2013 3013 2027 3027
rect 2053 3013 2067 3027
rect 2113 3013 2127 3027
rect 2133 3013 2147 3027
rect 1893 2993 1907 3007
rect 1853 2773 1867 2787
rect 1893 2773 1907 2787
rect 2073 2993 2087 3007
rect 2073 2953 2087 2967
rect 2053 2793 2067 2807
rect 1933 2773 1947 2787
rect 1993 2773 2007 2787
rect 1713 2693 1727 2707
rect 1653 2653 1667 2667
rect 1633 2633 1647 2647
rect 1613 2613 1627 2627
rect 1513 2553 1527 2567
rect 1493 2513 1507 2527
rect 1553 2513 1567 2527
rect 1293 2493 1307 2507
rect 1413 2493 1427 2507
rect 1453 2473 1467 2487
rect 1433 2413 1447 2427
rect 1253 2373 1267 2387
rect 1313 2293 1327 2307
rect 1333 2233 1347 2247
rect 1433 2233 1447 2247
rect 1273 2173 1287 2187
rect 1193 2073 1207 2087
rect 1173 2033 1187 2047
rect 1173 1973 1187 1987
rect 1173 1913 1187 1927
rect 1153 1873 1167 1887
rect 1193 1873 1207 1887
rect 1133 1813 1147 1827
rect 1233 2033 1247 2047
rect 1253 1993 1267 2007
rect 1213 1853 1227 1867
rect 1353 2133 1367 2147
rect 1633 2393 1647 2407
rect 1533 2313 1547 2327
rect 1613 2313 1627 2327
rect 1473 2273 1487 2287
rect 1513 2253 1527 2267
rect 1553 2253 1567 2267
rect 1573 2273 1587 2287
rect 1493 2233 1507 2247
rect 1533 2213 1547 2227
rect 1513 2153 1527 2167
rect 1493 2113 1507 2127
rect 1453 2093 1467 2107
rect 1353 2053 1367 2067
rect 1453 2073 1467 2087
rect 1473 2053 1487 2067
rect 1493 2073 1507 2087
rect 1513 2053 1527 2067
rect 1353 1973 1367 1987
rect 1413 1953 1427 1967
rect 1433 1953 1447 1967
rect 1473 1953 1487 1967
rect 1353 1913 1367 1927
rect 1313 1853 1327 1867
rect 1193 1833 1207 1847
rect 1233 1833 1247 1847
rect 1273 1833 1287 1847
rect 1193 1793 1207 1807
rect 1173 1773 1187 1787
rect 1113 1753 1127 1767
rect 1133 1753 1147 1767
rect 953 1693 967 1707
rect 1173 1653 1187 1667
rect 913 1533 927 1547
rect 1133 1633 1147 1647
rect 1053 1613 1067 1627
rect 1073 1613 1087 1627
rect 1093 1613 1107 1627
rect 1193 1633 1207 1647
rect 1093 1593 1107 1607
rect 1073 1573 1087 1587
rect 1113 1573 1127 1587
rect 1133 1593 1147 1607
rect 1053 1553 1067 1567
rect 933 1493 947 1507
rect 993 1513 1007 1527
rect 1153 1533 1167 1547
rect 1173 1453 1187 1467
rect 1073 1413 1087 1427
rect 913 1353 927 1367
rect 973 1353 987 1367
rect 893 1293 907 1307
rect 873 1253 887 1267
rect 813 1173 827 1187
rect 753 1153 767 1167
rect 813 1153 827 1167
rect 793 1133 807 1147
rect 573 1073 587 1087
rect 493 873 507 887
rect 533 873 547 887
rect 653 1093 667 1107
rect 693 1093 707 1107
rect 613 1013 627 1027
rect 673 913 687 927
rect 753 1073 767 1087
rect 833 1113 847 1127
rect 853 1113 867 1127
rect 793 1093 807 1107
rect 833 1053 847 1067
rect 773 1013 787 1027
rect 833 1013 847 1027
rect 753 933 767 947
rect 813 933 827 947
rect 793 893 807 907
rect 713 873 727 887
rect 613 853 627 867
rect 653 853 667 867
rect 473 833 487 847
rect 493 813 507 827
rect 513 813 527 827
rect 473 773 487 787
rect 453 753 467 767
rect 393 733 407 747
rect 253 693 267 707
rect 233 673 247 687
rect 73 593 87 607
rect 133 613 147 627
rect 253 653 267 667
rect 313 653 327 667
rect 373 653 387 667
rect 453 653 467 667
rect 293 633 307 647
rect 253 613 267 627
rect 113 593 127 607
rect 133 593 147 607
rect 193 593 207 607
rect 233 593 247 607
rect 53 453 67 467
rect 13 313 27 327
rect 153 333 167 347
rect 113 313 127 327
rect 273 553 287 567
rect 333 633 347 647
rect 353 613 367 627
rect 413 613 427 627
rect 353 593 367 607
rect 313 533 327 547
rect 453 613 467 627
rect 433 593 447 607
rect 413 573 427 587
rect 413 553 427 567
rect 393 513 407 527
rect 473 513 487 527
rect 253 373 267 387
rect 393 453 407 467
rect 373 313 387 327
rect 113 173 127 187
rect 153 153 167 167
rect 273 153 287 167
rect 353 173 367 187
rect 453 413 467 427
rect 593 833 607 847
rect 573 813 587 827
rect 693 853 707 867
rect 753 853 767 867
rect 513 753 527 767
rect 613 813 627 827
rect 573 793 587 807
rect 573 753 587 767
rect 553 733 567 747
rect 533 653 547 667
rect 733 813 747 827
rect 673 753 687 767
rect 693 733 707 747
rect 773 813 787 827
rect 793 813 807 827
rect 753 773 767 787
rect 753 653 767 667
rect 533 593 547 607
rect 553 613 567 627
rect 593 613 607 627
rect 593 593 607 607
rect 633 613 647 627
rect 673 613 687 627
rect 713 613 727 627
rect 733 613 747 627
rect 653 593 667 607
rect 773 593 787 607
rect 553 573 567 587
rect 573 553 587 567
rect 553 533 567 547
rect 513 413 527 427
rect 453 353 467 367
rect 513 373 527 387
rect 493 353 507 367
rect 533 353 547 367
rect 613 573 627 587
rect 633 573 647 587
rect 833 853 847 867
rect 933 1333 947 1347
rect 953 1313 967 1327
rect 1013 1333 1027 1347
rect 973 1293 987 1307
rect 993 1293 1007 1307
rect 913 1153 927 1167
rect 1133 1293 1147 1307
rect 1173 1293 1187 1307
rect 1033 1273 1047 1287
rect 973 1133 987 1147
rect 953 1113 967 1127
rect 913 1093 927 1107
rect 973 1093 987 1107
rect 933 1073 947 1087
rect 953 1073 967 1087
rect 893 1053 907 1067
rect 933 1053 947 1067
rect 893 893 907 907
rect 873 853 887 867
rect 993 1073 1007 1087
rect 1173 1073 1187 1087
rect 1213 1613 1227 1627
rect 1213 1593 1227 1607
rect 1253 1813 1267 1827
rect 1293 1813 1307 1827
rect 1293 1693 1307 1707
rect 1273 1673 1287 1687
rect 1253 1633 1267 1647
rect 1233 1573 1247 1587
rect 1393 1893 1407 1907
rect 1353 1833 1367 1847
rect 1393 1833 1407 1847
rect 1333 1813 1347 1827
rect 1373 1813 1387 1827
rect 1373 1793 1387 1807
rect 1433 1913 1447 1927
rect 1453 1873 1467 1887
rect 1453 1773 1467 1787
rect 1413 1753 1427 1767
rect 1393 1693 1407 1707
rect 1373 1673 1387 1687
rect 1353 1653 1367 1667
rect 1353 1573 1367 1587
rect 1253 1553 1267 1567
rect 1273 1553 1287 1567
rect 1313 1553 1327 1567
rect 1213 1453 1227 1467
rect 1353 1533 1367 1547
rect 1313 1493 1327 1507
rect 1253 1353 1267 1367
rect 1513 1893 1527 1907
rect 1493 1753 1507 1767
rect 1493 1673 1507 1687
rect 1513 1673 1527 1687
rect 1473 1653 1487 1667
rect 1453 1633 1467 1647
rect 1413 1593 1427 1607
rect 1433 1573 1447 1587
rect 1413 1553 1427 1567
rect 1413 1513 1427 1527
rect 1393 1473 1407 1487
rect 1433 1433 1447 1447
rect 1373 1413 1387 1427
rect 1333 1373 1347 1387
rect 1253 1293 1267 1307
rect 1313 1313 1327 1327
rect 953 913 967 927
rect 973 913 987 927
rect 933 853 947 867
rect 1033 893 1047 907
rect 1033 873 1047 887
rect 873 813 887 827
rect 913 813 927 827
rect 953 813 967 827
rect 993 813 1007 827
rect 833 753 847 767
rect 853 673 867 687
rect 873 653 887 667
rect 833 633 847 647
rect 1013 773 1027 787
rect 953 733 967 747
rect 913 673 927 687
rect 853 593 867 607
rect 893 593 907 607
rect 793 573 807 587
rect 833 573 847 587
rect 633 533 647 547
rect 673 393 687 407
rect 753 393 767 407
rect 473 313 487 327
rect 573 293 587 307
rect 553 193 567 207
rect 573 193 587 207
rect 693 333 707 347
rect 633 293 647 307
rect 673 293 687 307
rect 773 313 787 327
rect 733 293 747 307
rect 653 193 667 207
rect 713 193 727 207
rect 613 153 627 167
rect 653 153 667 167
rect 593 113 607 127
rect 633 113 647 127
rect 713 153 727 167
rect 933 553 947 567
rect 913 533 927 547
rect 853 373 867 387
rect 833 353 847 367
rect 853 353 867 367
rect 813 213 827 227
rect 873 213 887 227
rect 753 153 767 167
rect 833 173 847 187
rect 853 113 867 127
rect 973 633 987 647
rect 993 613 1007 627
rect 1093 853 1107 867
rect 1053 813 1067 827
rect 1073 833 1087 847
rect 1193 913 1207 927
rect 1413 1393 1427 1407
rect 1293 1093 1307 1107
rect 1333 1093 1347 1107
rect 1333 913 1347 927
rect 1233 893 1247 907
rect 1273 893 1287 907
rect 1133 813 1147 827
rect 1173 813 1187 827
rect 1253 833 1267 847
rect 1353 853 1367 867
rect 1333 813 1347 827
rect 1093 753 1107 767
rect 1133 753 1147 767
rect 1233 793 1247 807
rect 1133 313 1147 327
rect 973 193 987 207
rect 953 153 967 167
rect 1113 273 1127 287
rect 1133 213 1147 227
rect 1153 213 1167 227
rect 993 93 1007 107
rect 1093 133 1107 147
rect 1433 1313 1447 1327
rect 1473 1593 1487 1607
rect 1593 2193 1607 2207
rect 1673 2613 1687 2627
rect 1813 2733 1827 2747
rect 1833 2753 1847 2767
rect 1853 2733 1867 2747
rect 1913 2753 1927 2767
rect 1893 2733 1907 2747
rect 1853 2713 1867 2727
rect 1793 2633 1807 2647
rect 1833 2633 1847 2647
rect 1753 2533 1767 2547
rect 1813 2573 1827 2587
rect 1813 2533 1827 2547
rect 1933 2633 1947 2647
rect 1893 2593 1907 2607
rect 1893 2573 1907 2587
rect 1913 2533 1927 2547
rect 1733 2433 1747 2447
rect 1653 2313 1667 2327
rect 1633 2293 1647 2307
rect 1653 2293 1667 2307
rect 1713 2293 1727 2307
rect 1693 2273 1707 2287
rect 1673 2253 1687 2267
rect 1653 2193 1667 2207
rect 1693 2193 1707 2207
rect 1633 2113 1647 2127
rect 1693 2173 1707 2187
rect 1553 2093 1567 2107
rect 1613 2093 1627 2107
rect 1733 2253 1747 2267
rect 1793 2253 1807 2267
rect 1773 2233 1787 2247
rect 1793 2213 1807 2227
rect 1753 2173 1767 2187
rect 1573 2073 1587 2087
rect 1553 2053 1567 2067
rect 1633 2053 1647 2067
rect 1653 2053 1667 2067
rect 1713 2073 1727 2087
rect 1773 2153 1787 2167
rect 1993 2613 2007 2627
rect 1973 2573 1987 2587
rect 2133 2993 2147 3007
rect 2173 3013 2187 3027
rect 2213 3013 2227 3027
rect 2373 3173 2387 3187
rect 2373 3073 2387 3087
rect 2193 2993 2207 3007
rect 2253 2993 2267 3007
rect 2353 3033 2367 3047
rect 2213 2973 2227 2987
rect 2153 2953 2167 2967
rect 2193 2953 2207 2967
rect 2253 2933 2267 2947
rect 2313 2893 2327 2907
rect 2173 2813 2187 2827
rect 2073 2753 2087 2767
rect 2053 2733 2067 2747
rect 2033 2653 2047 2667
rect 2033 2613 2047 2627
rect 2013 2573 2027 2587
rect 1953 2553 1967 2567
rect 2013 2533 2027 2547
rect 2093 2733 2107 2747
rect 2113 2753 2127 2767
rect 2133 2753 2147 2767
rect 2153 2753 2167 2767
rect 2073 2693 2087 2707
rect 2133 2693 2147 2707
rect 2113 2673 2127 2687
rect 2073 2573 2087 2587
rect 2093 2533 2107 2547
rect 2193 2733 2207 2747
rect 2173 2633 2187 2647
rect 2173 2593 2187 2607
rect 2133 2533 2147 2547
rect 1973 2493 1987 2507
rect 2053 2493 2067 2507
rect 1933 2473 1947 2487
rect 1913 2393 1927 2407
rect 1893 2373 1907 2387
rect 1873 2253 1887 2267
rect 1853 2233 1867 2247
rect 2053 2353 2067 2367
rect 1973 2273 1987 2287
rect 1993 2253 2007 2267
rect 2033 2273 2047 2287
rect 2053 2273 2067 2287
rect 2073 2273 2087 2287
rect 1913 2233 1927 2247
rect 1953 2213 1967 2227
rect 1833 2193 1847 2207
rect 1833 2173 1847 2187
rect 1813 2093 1827 2107
rect 1733 2053 1747 2067
rect 1813 2073 1827 2087
rect 1573 1993 1587 2007
rect 1713 2033 1727 2047
rect 1673 1973 1687 1987
rect 1633 1953 1647 1967
rect 1613 1873 1627 1887
rect 1553 1713 1567 1727
rect 1533 1633 1547 1647
rect 1593 1633 1607 1647
rect 1633 1753 1647 1767
rect 1533 1613 1547 1627
rect 1613 1613 1627 1627
rect 1493 1573 1507 1587
rect 1513 1573 1527 1587
rect 1553 1573 1567 1587
rect 1473 1553 1487 1567
rect 1493 1533 1507 1547
rect 1473 1413 1487 1427
rect 1453 1233 1467 1247
rect 1433 1093 1447 1107
rect 1433 1073 1447 1087
rect 1673 1713 1687 1727
rect 1793 1953 1807 1967
rect 1733 1853 1747 1867
rect 1913 2153 1927 2167
rect 1933 2153 1947 2167
rect 2053 2153 2067 2167
rect 1933 2133 1947 2147
rect 1953 2133 1967 2147
rect 1913 2113 1927 2127
rect 1853 2073 1867 2087
rect 1873 2053 1887 2067
rect 1873 1973 1887 1987
rect 1993 2073 2007 2087
rect 1993 2033 2007 2047
rect 2233 2793 2247 2807
rect 2273 2773 2287 2787
rect 2293 2713 2307 2727
rect 2293 2693 2307 2707
rect 2273 2653 2287 2667
rect 2293 2593 2307 2607
rect 2253 2573 2267 2587
rect 2233 2553 2247 2567
rect 2213 2513 2227 2527
rect 2333 2853 2347 2867
rect 2373 2793 2387 2807
rect 2373 2633 2387 2647
rect 2333 2593 2347 2607
rect 2373 2573 2387 2587
rect 2333 2533 2347 2547
rect 2353 2553 2367 2567
rect 2313 2513 2327 2527
rect 2273 2473 2287 2487
rect 2253 2433 2267 2447
rect 2313 2433 2327 2447
rect 2353 2433 2367 2447
rect 2213 2393 2227 2407
rect 2153 2253 2167 2267
rect 2173 2233 2187 2247
rect 2153 2173 2167 2187
rect 2133 2093 2147 2107
rect 2113 2073 2127 2087
rect 2093 2013 2107 2027
rect 2113 2013 2127 2027
rect 2073 1993 2087 2007
rect 1993 1973 2007 1987
rect 2013 1973 2027 1987
rect 2073 1953 2087 1967
rect 1973 1933 1987 1947
rect 2013 1893 2027 1907
rect 1873 1873 1887 1887
rect 1913 1873 1927 1887
rect 1953 1873 1967 1887
rect 1813 1833 1827 1847
rect 1953 1853 1967 1867
rect 1813 1773 1827 1787
rect 1833 1793 1847 1807
rect 1853 1773 1867 1787
rect 1913 1793 1927 1807
rect 2013 1813 2027 1827
rect 1693 1693 1707 1707
rect 1853 1733 1867 1747
rect 1813 1693 1827 1707
rect 1753 1633 1767 1647
rect 1633 1573 1647 1587
rect 1593 1513 1607 1527
rect 1573 1493 1587 1507
rect 1573 1373 1587 1387
rect 1553 1353 1567 1367
rect 1533 1233 1547 1247
rect 1493 1053 1507 1067
rect 1613 1453 1627 1467
rect 1753 1613 1767 1627
rect 1713 1593 1727 1607
rect 1733 1533 1747 1547
rect 1693 1513 1707 1527
rect 1673 1493 1687 1507
rect 1773 1593 1787 1607
rect 1753 1433 1767 1447
rect 1733 1413 1747 1427
rect 1773 1413 1787 1427
rect 1673 1373 1687 1387
rect 1713 1373 1727 1387
rect 1633 1353 1647 1367
rect 1653 1353 1667 1367
rect 1613 1333 1627 1347
rect 1593 1273 1607 1287
rect 1553 1213 1567 1227
rect 1553 1153 1567 1167
rect 1573 1093 1587 1107
rect 1453 853 1467 867
rect 1413 793 1427 807
rect 1473 793 1487 807
rect 1353 653 1367 667
rect 1373 653 1387 667
rect 1273 633 1287 647
rect 1313 633 1327 647
rect 1213 333 1227 347
rect 1633 1273 1647 1287
rect 1633 1253 1647 1267
rect 1613 1013 1627 1027
rect 1573 813 1587 827
rect 1693 1293 1707 1307
rect 1753 1393 1767 1407
rect 1753 1353 1767 1367
rect 1773 1313 1787 1327
rect 1733 1293 1747 1307
rect 1753 1293 1767 1307
rect 1773 1273 1787 1287
rect 1673 1113 1687 1127
rect 1833 1633 1847 1647
rect 1853 1613 1867 1627
rect 2013 1773 2027 1787
rect 1913 1753 1927 1767
rect 1973 1753 1987 1767
rect 1893 1693 1907 1707
rect 1953 1693 1967 1707
rect 1873 1573 1887 1587
rect 1873 1513 1887 1527
rect 1953 1553 1967 1567
rect 2093 1933 2107 1947
rect 2113 1893 2127 1907
rect 2133 1893 2147 1907
rect 2133 1873 2147 1887
rect 2153 1873 2167 1887
rect 2093 1793 2107 1807
rect 2233 2373 2247 2387
rect 2293 2353 2307 2367
rect 2233 2253 2247 2267
rect 2273 2273 2287 2287
rect 2273 2213 2287 2227
rect 2233 2153 2247 2167
rect 2213 2113 2227 2127
rect 2293 2133 2307 2147
rect 2273 2073 2287 2087
rect 2273 2033 2287 2047
rect 2233 1973 2247 1987
rect 2213 1853 2227 1867
rect 2133 1733 2147 1747
rect 2173 1733 2187 1747
rect 2073 1713 2087 1727
rect 2013 1653 2027 1667
rect 2213 1733 2227 1747
rect 2373 2413 2387 2427
rect 2413 3213 2427 3227
rect 2553 3553 2567 3567
rect 2553 3533 2567 3547
rect 2633 3533 2647 3547
rect 2793 3773 2807 3787
rect 2833 3753 2847 3767
rect 2913 3753 2927 3767
rect 2973 3753 2987 3767
rect 2773 3733 2787 3747
rect 2813 3733 2827 3747
rect 2773 3713 2787 3727
rect 2893 3733 2907 3747
rect 2673 3613 2687 3627
rect 2673 3573 2687 3587
rect 2753 3693 2767 3707
rect 2893 3693 2907 3707
rect 2953 3713 2967 3727
rect 2953 3693 2967 3707
rect 2793 3673 2807 3687
rect 2853 3673 2867 3687
rect 2753 3533 2767 3547
rect 2693 3493 2707 3507
rect 2753 3473 2767 3487
rect 2813 3553 2827 3567
rect 2933 3613 2947 3627
rect 2853 3533 2867 3547
rect 2873 3533 2887 3547
rect 2833 3513 2847 3527
rect 2793 3493 2807 3507
rect 3113 3793 3127 3807
rect 3093 3753 3107 3767
rect 3033 3733 3047 3747
rect 3173 3773 3187 3787
rect 3133 3733 3147 3747
rect 3013 3713 3027 3727
rect 3073 3713 3087 3727
rect 3113 3713 3127 3727
rect 3053 3693 3067 3707
rect 3173 3713 3187 3727
rect 3153 3693 3167 3707
rect 3113 3673 3127 3687
rect 3253 3953 3267 3967
rect 3293 3953 3307 3967
rect 3313 3953 3327 3967
rect 3353 3973 3367 3987
rect 3233 3933 3247 3947
rect 3333 3933 3347 3947
rect 3333 3793 3347 3807
rect 3473 3993 3487 4007
rect 3453 3773 3467 3787
rect 3273 3753 3287 3767
rect 3313 3753 3327 3767
rect 3333 3753 3347 3767
rect 3373 3753 3387 3767
rect 3233 3733 3247 3747
rect 3313 3733 3327 3747
rect 3213 3693 3227 3707
rect 3233 3713 3247 3727
rect 3233 3673 3247 3687
rect 3053 3653 3067 3667
rect 3193 3653 3207 3667
rect 2993 3613 3007 3627
rect 3033 3613 3047 3627
rect 2973 3573 2987 3587
rect 3033 3573 3047 3587
rect 3353 3713 3367 3727
rect 3293 3673 3307 3687
rect 3313 3673 3327 3687
rect 3253 3653 3267 3667
rect 3293 3653 3307 3667
rect 2973 3533 2987 3547
rect 3033 3533 3047 3547
rect 3093 3533 3107 3547
rect 3133 3533 3147 3547
rect 3153 3533 3167 3547
rect 3233 3533 3247 3547
rect 3273 3533 3287 3547
rect 2913 3513 2927 3527
rect 3013 3493 3027 3507
rect 3033 3493 3047 3507
rect 3053 3493 3067 3507
rect 3073 3513 3087 3527
rect 2913 3473 2927 3487
rect 2833 3453 2847 3467
rect 2893 3453 2907 3467
rect 2773 3433 2787 3447
rect 2853 3433 2867 3447
rect 2873 3433 2887 3447
rect 2653 3413 2667 3427
rect 2593 3333 2607 3347
rect 2553 3253 2567 3267
rect 2473 3213 2487 3227
rect 2433 3193 2447 3207
rect 2413 3013 2427 3027
rect 2513 3213 2527 3227
rect 2533 3233 2547 3247
rect 2553 3213 2567 3227
rect 2493 3193 2507 3207
rect 2553 3193 2567 3207
rect 2493 3113 2507 3127
rect 2453 3053 2467 3067
rect 2473 3033 2487 3047
rect 2553 3073 2567 3087
rect 2493 2853 2507 2867
rect 2413 2793 2427 2807
rect 2433 2753 2447 2767
rect 2453 2773 2467 2787
rect 2513 2773 2527 2787
rect 2413 2653 2427 2667
rect 2393 2313 2407 2327
rect 2733 3273 2747 3287
rect 2853 3293 2867 3307
rect 2653 3013 2667 3027
rect 2613 2993 2627 3007
rect 2573 2753 2587 2767
rect 2533 2693 2547 2707
rect 2493 2593 2507 2607
rect 2533 2593 2547 2607
rect 2553 2593 2567 2607
rect 2473 2513 2487 2527
rect 2453 2413 2467 2427
rect 2413 2293 2427 2307
rect 2433 2293 2447 2307
rect 2353 2273 2367 2287
rect 2373 2253 2387 2267
rect 2413 2273 2427 2287
rect 2453 2273 2467 2287
rect 2433 2253 2447 2267
rect 2453 2253 2467 2267
rect 2353 2233 2367 2247
rect 2393 2233 2407 2247
rect 2333 2193 2347 2207
rect 2393 2173 2407 2187
rect 2373 2133 2387 2147
rect 2313 2033 2327 2047
rect 2373 2073 2387 2087
rect 2293 1993 2307 2007
rect 2353 1933 2367 1947
rect 2433 2153 2447 2167
rect 2553 2533 2567 2547
rect 2653 2593 2667 2607
rect 2593 2553 2607 2567
rect 2593 2533 2607 2547
rect 2553 2433 2567 2447
rect 2573 2413 2587 2427
rect 2533 2333 2547 2347
rect 2553 2333 2567 2347
rect 2613 2493 2627 2507
rect 2613 2433 2627 2447
rect 2613 2413 2627 2427
rect 2593 2393 2607 2407
rect 2573 2313 2587 2327
rect 2513 2293 2527 2307
rect 2553 2293 2567 2307
rect 2693 3033 2707 3047
rect 2793 3213 2807 3227
rect 2713 2853 2727 2867
rect 2833 3213 2847 3227
rect 2833 3153 2847 3167
rect 2793 3133 2807 3147
rect 3193 3513 3207 3527
rect 3153 3493 3167 3507
rect 3233 3513 3247 3527
rect 3253 3493 3267 3507
rect 3093 3473 3107 3487
rect 3033 3453 3047 3467
rect 3133 3473 3147 3487
rect 3113 3413 3127 3427
rect 3073 3373 3087 3387
rect 3033 3353 3047 3367
rect 2953 3333 2967 3347
rect 2913 3293 2927 3307
rect 2873 3273 2887 3287
rect 2893 3273 2907 3287
rect 2933 3273 2947 3287
rect 2873 3253 2887 3267
rect 2913 3253 2927 3267
rect 2873 3213 2887 3227
rect 2893 3193 2907 3207
rect 2873 3073 2887 3087
rect 2933 3173 2947 3187
rect 2913 3153 2927 3167
rect 2973 3273 2987 3287
rect 3013 3273 3027 3287
rect 3053 3313 3067 3327
rect 2993 3233 3007 3247
rect 3033 3253 3047 3267
rect 3073 3253 3087 3267
rect 3053 3233 3067 3247
rect 3033 3213 3047 3227
rect 3073 3213 3087 3227
rect 3093 3233 3107 3247
rect 3113 3213 3127 3227
rect 2913 3093 2927 3107
rect 2953 3093 2967 3107
rect 2873 3053 2887 3067
rect 2893 3053 2907 3067
rect 3213 3453 3227 3467
rect 3253 3413 3267 3427
rect 3233 3373 3247 3387
rect 3153 3293 3167 3307
rect 3193 3273 3207 3287
rect 3173 3233 3187 3247
rect 3433 3713 3447 3727
rect 3353 3593 3367 3607
rect 3393 3593 3407 3607
rect 3313 3493 3327 3507
rect 3333 3493 3347 3507
rect 3213 3213 3227 3227
rect 3253 3193 3267 3207
rect 3573 4133 3587 4147
rect 3553 4113 3567 4127
rect 3513 4013 3527 4027
rect 3553 3993 3567 4007
rect 3593 3993 3607 4007
rect 3673 4053 3687 4067
rect 3653 3953 3667 3967
rect 3613 3873 3627 3887
rect 3493 3713 3507 3727
rect 3533 3773 3547 3787
rect 3733 4633 3747 4647
rect 3773 4613 3787 4627
rect 3813 4553 3827 4567
rect 3753 4433 3767 4447
rect 3913 4613 3927 4627
rect 3993 4773 4007 4787
rect 3933 4553 3947 4567
rect 3853 4533 3867 4547
rect 3933 4513 3947 4527
rect 3853 4493 3867 4507
rect 3853 4453 3867 4467
rect 3873 4473 3887 4487
rect 3733 4413 3747 4427
rect 3833 4433 3847 4447
rect 3813 4313 3827 4327
rect 3733 4193 3747 4207
rect 3793 4193 3807 4207
rect 3813 4173 3827 4187
rect 3753 4113 3767 4127
rect 3773 4033 3787 4047
rect 3813 4013 3827 4027
rect 3853 4313 3867 4327
rect 3933 4433 3947 4447
rect 3993 4613 4007 4627
rect 4053 4913 4067 4927
rect 4073 4853 4087 4867
rect 4053 4633 4067 4647
rect 3953 4413 3967 4427
rect 4013 4473 4027 4487
rect 4033 4413 4047 4427
rect 4113 4913 4127 4927
rect 4233 5413 4247 5427
rect 4153 5253 4167 5267
rect 4193 5333 4207 5347
rect 4213 5333 4227 5347
rect 4213 5313 4227 5327
rect 4193 5253 4207 5267
rect 4173 5213 4187 5227
rect 4213 5193 4227 5207
rect 4153 5173 4167 5187
rect 4173 5153 4187 5167
rect 4153 5133 4167 5147
rect 4173 5133 4187 5147
rect 4153 4973 4167 4987
rect 4393 5713 4407 5727
rect 4533 5733 4547 5747
rect 4493 5693 4507 5707
rect 4513 5693 4527 5707
rect 4393 5653 4407 5667
rect 4413 5633 4427 5647
rect 4373 5613 4387 5627
rect 4433 5613 4447 5627
rect 4453 5633 4467 5647
rect 4653 5913 4667 5927
rect 4613 5713 4627 5727
rect 4653 5753 4667 5767
rect 4653 5733 4667 5747
rect 4633 5693 4647 5707
rect 4593 5673 4607 5687
rect 4553 5653 4567 5667
rect 4593 5653 4607 5667
rect 4613 5633 4627 5647
rect 4593 5613 4607 5627
rect 4333 5593 4347 5607
rect 4433 5593 4447 5607
rect 4473 5593 4487 5607
rect 4313 5553 4327 5567
rect 4573 5553 4587 5567
rect 4433 5533 4447 5547
rect 4513 5533 4527 5547
rect 4313 5413 4327 5427
rect 4373 5433 4387 5447
rect 4493 5453 4507 5467
rect 4553 5513 4567 5527
rect 4533 5473 4547 5487
rect 4513 5433 4527 5447
rect 4393 5413 4407 5427
rect 4293 5373 4307 5387
rect 4293 5353 4307 5367
rect 4273 5313 4287 5327
rect 4273 5213 4287 5227
rect 4233 5173 4247 5187
rect 4253 5173 4267 5187
rect 4253 5133 4267 5147
rect 4213 5113 4227 5127
rect 4233 5093 4247 5107
rect 4373 5393 4387 5407
rect 4373 5353 4387 5367
rect 4353 5333 4367 5347
rect 4353 5273 4367 5287
rect 4313 5213 4327 5227
rect 4273 5113 4287 5127
rect 4373 5213 4387 5227
rect 4333 5173 4347 5187
rect 4353 5153 4367 5167
rect 4453 5393 4467 5407
rect 4513 5393 4527 5407
rect 4433 5373 4447 5387
rect 4453 5373 4467 5387
rect 4473 5353 4487 5367
rect 4513 5353 4527 5367
rect 4493 5333 4507 5347
rect 4533 5333 4547 5347
rect 4433 5293 4447 5307
rect 4413 5233 4427 5247
rect 4473 5273 4487 5287
rect 4453 5213 4467 5227
rect 4433 5173 4447 5187
rect 4393 5153 4407 5167
rect 4333 5133 4347 5147
rect 4293 5093 4307 5107
rect 4313 5093 4327 5107
rect 4273 5073 4287 5087
rect 4293 5073 4307 5087
rect 4253 5013 4267 5027
rect 4273 5013 4287 5027
rect 4213 4993 4227 5007
rect 4193 4973 4207 4987
rect 4253 4953 4267 4967
rect 4433 5133 4447 5147
rect 4453 5153 4467 5167
rect 4613 5593 4627 5607
rect 4633 5533 4647 5547
rect 4733 6093 4747 6107
rect 4873 6173 4887 6187
rect 4873 6133 4887 6147
rect 4793 6113 4807 6127
rect 4833 6113 4847 6127
rect 5533 6473 5547 6487
rect 5473 6453 5487 6467
rect 5493 6453 5507 6467
rect 5153 6433 5167 6447
rect 5213 6433 5227 6447
rect 5333 6433 5347 6447
rect 5353 6433 5367 6447
rect 5133 6353 5147 6367
rect 5213 6393 5227 6407
rect 5193 6373 5207 6387
rect 5253 6373 5267 6387
rect 5293 6373 5307 6387
rect 5373 6393 5387 6407
rect 5393 6393 5407 6407
rect 5493 6433 5507 6447
rect 5393 6373 5407 6387
rect 5233 6333 5247 6347
rect 5253 6333 5267 6347
rect 5293 6333 5307 6347
rect 5313 6333 5327 6347
rect 5213 6313 5227 6327
rect 5033 6293 5047 6307
rect 5093 6293 5107 6307
rect 5113 6273 5127 6287
rect 5033 6153 5047 6167
rect 4813 6073 4827 6087
rect 4873 6073 4887 6087
rect 4773 6053 4787 6067
rect 4693 6033 4707 6047
rect 4753 6033 4767 6047
rect 4713 5973 4727 5987
rect 4693 5953 4707 5967
rect 4753 5953 4767 5967
rect 4733 5893 4747 5907
rect 4753 5893 4767 5907
rect 4693 5833 4707 5847
rect 4733 5833 4747 5847
rect 4773 5873 4787 5887
rect 4813 5893 4827 5907
rect 4853 5893 4867 5907
rect 4793 5713 4807 5727
rect 4853 5853 4867 5867
rect 4933 6113 4947 6127
rect 4913 6093 4927 6107
rect 4913 6073 4927 6087
rect 4893 6053 4907 6067
rect 4913 5933 4927 5947
rect 4893 5873 4907 5887
rect 4993 6093 5007 6107
rect 4973 5973 4987 5987
rect 5013 5953 5027 5967
rect 5293 6293 5307 6307
rect 5253 6253 5267 6267
rect 5213 6153 5227 6167
rect 5273 6153 5287 6167
rect 5113 6133 5127 6147
rect 5093 6093 5107 6107
rect 5113 6113 5127 6127
rect 5153 6093 5167 6107
rect 5113 6073 5127 6087
rect 5073 6053 5087 6067
rect 5053 5953 5067 5967
rect 5033 5933 5047 5947
rect 5053 5933 5067 5947
rect 4973 5893 4987 5907
rect 5033 5893 5047 5907
rect 5053 5893 5067 5907
rect 5093 5913 5107 5927
rect 4993 5873 5007 5887
rect 5033 5873 5047 5887
rect 4893 5853 4907 5867
rect 4853 5733 4867 5747
rect 4873 5713 4887 5727
rect 4833 5693 4847 5707
rect 4853 5693 4867 5707
rect 4733 5653 4747 5667
rect 4753 5653 4767 5667
rect 4693 5633 4707 5647
rect 4713 5613 4727 5627
rect 4733 5633 4747 5647
rect 4773 5613 4787 5627
rect 4793 5633 4807 5647
rect 4733 5573 4747 5587
rect 4673 5473 4687 5487
rect 4793 5593 4807 5607
rect 4753 5553 4767 5567
rect 4773 5553 4787 5567
rect 4673 5433 4687 5447
rect 4693 5433 4707 5447
rect 4553 5273 4567 5287
rect 4513 5253 4527 5267
rect 4573 5253 4587 5267
rect 4593 5233 4607 5247
rect 4713 5413 4727 5427
rect 4733 5433 4747 5447
rect 4773 5533 4787 5547
rect 4853 5593 4867 5607
rect 4813 5573 4827 5587
rect 4853 5553 4867 5567
rect 4793 5473 4807 5487
rect 4773 5453 4787 5467
rect 4833 5453 4847 5467
rect 4773 5433 4787 5447
rect 4813 5413 4827 5427
rect 4673 5373 4687 5387
rect 4753 5373 4767 5387
rect 4633 5333 4647 5347
rect 4633 5293 4647 5307
rect 4613 5213 4627 5227
rect 4553 5173 4567 5187
rect 4513 5153 4527 5167
rect 4493 5133 4507 5147
rect 4533 5133 4547 5147
rect 4613 5153 4627 5167
rect 4633 5173 4647 5187
rect 4713 5353 4727 5367
rect 4673 5273 4687 5287
rect 4733 5253 4747 5267
rect 4693 5153 4707 5167
rect 5033 5833 5047 5847
rect 4973 5733 4987 5747
rect 4893 5573 4907 5587
rect 5213 6093 5227 6107
rect 5353 6293 5367 6307
rect 5453 6353 5467 6367
rect 5413 6273 5427 6287
rect 5413 6253 5427 6267
rect 5353 6133 5367 6147
rect 5353 6113 5367 6127
rect 5733 6453 5747 6467
rect 5793 6453 5807 6467
rect 5573 6433 5587 6447
rect 5613 6413 5627 6427
rect 5653 6413 5667 6427
rect 5553 6373 5567 6387
rect 5593 6333 5607 6347
rect 5493 6273 5507 6287
rect 5693 6413 5707 6427
rect 5633 6373 5647 6387
rect 5753 6433 5767 6447
rect 6173 6473 6187 6487
rect 6013 6453 6027 6467
rect 6053 6453 6067 6467
rect 6153 6453 6167 6467
rect 6033 6433 6047 6447
rect 5933 6413 5947 6427
rect 5973 6413 5987 6427
rect 5673 6373 5687 6387
rect 5753 6393 5767 6407
rect 5793 6393 5807 6407
rect 5873 6393 5887 6407
rect 5673 6353 5687 6367
rect 5733 6353 5747 6367
rect 5713 6333 5727 6347
rect 5553 6253 5567 6267
rect 5613 6253 5627 6267
rect 5453 6193 5467 6207
rect 5533 6153 5547 6167
rect 5433 6133 5447 6147
rect 5373 6093 5387 6107
rect 5473 6113 5487 6127
rect 5593 6133 5607 6147
rect 5713 6153 5727 6167
rect 5193 6073 5207 6087
rect 5173 6033 5187 6047
rect 5193 5973 5207 5987
rect 5193 5953 5207 5967
rect 5133 5913 5147 5927
rect 5333 6073 5347 6087
rect 5493 6073 5507 6087
rect 5273 6053 5287 6067
rect 5233 5933 5247 5947
rect 5373 5953 5387 5967
rect 5613 6113 5627 6127
rect 5633 6113 5647 6127
rect 5593 6073 5607 6087
rect 5613 6073 5627 6087
rect 5453 5933 5467 5947
rect 5493 5933 5507 5947
rect 5213 5893 5227 5907
rect 5333 5913 5347 5927
rect 5093 5873 5107 5887
rect 5113 5873 5127 5887
rect 5153 5873 5167 5887
rect 5173 5873 5187 5887
rect 5233 5873 5247 5887
rect 5253 5873 5267 5887
rect 5073 5853 5087 5867
rect 5113 5833 5127 5847
rect 5153 5793 5167 5807
rect 5013 5653 5027 5667
rect 5093 5653 5107 5667
rect 5113 5653 5127 5667
rect 4953 5633 4967 5647
rect 5053 5633 5067 5647
rect 5033 5613 5047 5627
rect 5093 5633 5107 5647
rect 5113 5613 5127 5627
rect 5133 5613 5147 5627
rect 4953 5593 4967 5607
rect 5053 5593 5067 5607
rect 4933 5573 4947 5587
rect 4993 5573 5007 5587
rect 5013 5573 5027 5587
rect 5053 5573 5067 5587
rect 4913 5553 4927 5567
rect 4933 5513 4947 5527
rect 4953 5453 4967 5467
rect 4873 5433 4887 5447
rect 4913 5413 4927 5427
rect 4893 5393 4907 5407
rect 4913 5393 4927 5407
rect 5053 5553 5067 5567
rect 5033 5473 5047 5487
rect 5013 5433 5027 5447
rect 4993 5413 5007 5427
rect 4853 5373 4867 5387
rect 4833 5353 4847 5367
rect 4813 5313 4827 5327
rect 4853 5333 4867 5347
rect 4793 5233 4807 5247
rect 4733 5153 4747 5167
rect 4773 5153 4787 5167
rect 4593 5133 4607 5147
rect 4613 5133 4627 5147
rect 4653 5133 4667 5147
rect 4693 5133 4707 5147
rect 4413 5113 4427 5127
rect 4433 5113 4447 5127
rect 4473 5113 4487 5127
rect 4333 5073 4347 5087
rect 4333 5033 4347 5047
rect 4353 5033 4367 5047
rect 4293 4953 4307 4967
rect 4233 4933 4247 4947
rect 4173 4913 4187 4927
rect 4193 4913 4207 4927
rect 4113 4893 4127 4907
rect 4133 4893 4147 4907
rect 4213 4893 4227 4907
rect 4093 4773 4107 4787
rect 4193 4753 4207 4767
rect 4153 4733 4167 4747
rect 4113 4693 4127 4707
rect 4153 4693 4167 4707
rect 4133 4673 4147 4687
rect 4193 4693 4207 4707
rect 4093 4593 4107 4607
rect 4173 4633 4187 4647
rect 4173 4593 4187 4607
rect 4093 4493 4107 4507
rect 4133 4513 4147 4527
rect 4133 4473 4147 4487
rect 4153 4473 4167 4487
rect 3993 4353 4007 4367
rect 4053 4353 4067 4367
rect 4073 4353 4087 4367
rect 3993 4313 4007 4327
rect 3913 4233 3927 4247
rect 4253 4913 4267 4927
rect 4273 4933 4287 4947
rect 4313 4913 4327 4927
rect 4253 4893 4267 4907
rect 4253 4813 4267 4827
rect 4413 5013 4427 5027
rect 4353 4993 4367 5007
rect 4373 4953 4387 4967
rect 4393 4933 4407 4947
rect 4353 4913 4367 4927
rect 4353 4893 4367 4907
rect 4313 4833 4327 4847
rect 4333 4833 4347 4847
rect 4473 5073 4487 5087
rect 4513 4993 4527 5007
rect 4433 4953 4447 4967
rect 4433 4933 4447 4947
rect 4473 4933 4487 4947
rect 4493 4953 4507 4967
rect 4413 4873 4427 4887
rect 4493 4913 4507 4927
rect 4653 5113 4667 5127
rect 4613 4993 4627 5007
rect 4593 4953 4607 4967
rect 4613 4953 4627 4967
rect 4553 4933 4567 4947
rect 4593 4933 4607 4947
rect 4673 4933 4687 4947
rect 4473 4853 4487 4867
rect 4353 4793 4367 4807
rect 4393 4793 4407 4807
rect 4273 4753 4287 4767
rect 4293 4733 4307 4747
rect 4373 4733 4387 4747
rect 4233 4693 4247 4707
rect 4233 4653 4247 4667
rect 4273 4693 4287 4707
rect 4293 4653 4307 4667
rect 4273 4593 4287 4607
rect 4313 4593 4327 4607
rect 4253 4513 4267 4527
rect 4233 4473 4247 4487
rect 4273 4493 4287 4507
rect 4353 4593 4367 4607
rect 4573 4853 4587 4867
rect 4633 4873 4647 4887
rect 4653 4833 4667 4847
rect 4633 4813 4647 4827
rect 4713 4973 4727 4987
rect 4913 5333 4927 5347
rect 4973 5373 4987 5387
rect 4933 5293 4947 5307
rect 4893 5253 4907 5267
rect 5013 5333 5027 5347
rect 4993 5293 5007 5307
rect 4933 5193 4947 5207
rect 4873 5153 4887 5167
rect 4873 5133 4887 5147
rect 4773 5113 4787 5127
rect 4753 4973 4767 4987
rect 4813 5093 4827 5107
rect 4833 5093 4847 5107
rect 4793 4973 4807 4987
rect 4913 5133 4927 5147
rect 5093 5593 5107 5607
rect 5073 5513 5087 5527
rect 5073 5393 5087 5407
rect 5393 5893 5407 5907
rect 5333 5873 5347 5887
rect 5353 5873 5367 5887
rect 5313 5853 5327 5867
rect 5273 5813 5287 5827
rect 5233 5793 5247 5807
rect 5313 5753 5327 5767
rect 5273 5733 5287 5747
rect 5193 5653 5207 5667
rect 5173 5633 5187 5647
rect 5253 5653 5267 5667
rect 5213 5613 5227 5627
rect 5153 5593 5167 5607
rect 5173 5593 5187 5607
rect 5173 5453 5187 5467
rect 5113 5433 5127 5447
rect 5133 5433 5147 5447
rect 5153 5433 5167 5447
rect 5073 5353 5087 5367
rect 5093 5353 5107 5367
rect 5033 5313 5047 5327
rect 5013 5273 5027 5287
rect 5033 5273 5047 5287
rect 5093 5313 5107 5327
rect 5053 5253 5067 5267
rect 5073 5253 5087 5267
rect 5033 5233 5047 5247
rect 5013 5193 5027 5207
rect 4733 4913 4747 4927
rect 4773 4913 4787 4927
rect 4713 4893 4727 4907
rect 4733 4873 4747 4887
rect 4753 4873 4767 4887
rect 4713 4833 4727 4847
rect 4693 4813 4707 4827
rect 4593 4753 4607 4767
rect 4673 4753 4687 4767
rect 4613 4733 4627 4747
rect 4473 4713 4487 4727
rect 4493 4713 4507 4727
rect 4453 4693 4467 4707
rect 4413 4653 4427 4667
rect 4513 4693 4527 4707
rect 4653 4713 4667 4727
rect 4673 4713 4687 4727
rect 4533 4653 4547 4667
rect 4493 4633 4507 4647
rect 4573 4633 4587 4647
rect 4633 4653 4647 4667
rect 4453 4593 4467 4607
rect 4613 4613 4627 4627
rect 4553 4573 4567 4587
rect 4373 4553 4387 4567
rect 4373 4493 4387 4507
rect 4413 4493 4427 4507
rect 4453 4493 4467 4507
rect 4513 4493 4527 4507
rect 4293 4453 4307 4467
rect 4333 4473 4347 4487
rect 4273 4433 4287 4447
rect 4293 4433 4307 4447
rect 4193 4393 4207 4407
rect 4273 4393 4287 4407
rect 4173 4373 4187 4387
rect 4253 4373 4267 4387
rect 4073 4313 4087 4327
rect 4153 4313 4167 4327
rect 4053 4293 4067 4307
rect 4133 4253 4147 4267
rect 4053 4233 4067 4247
rect 3873 4133 3887 4147
rect 3913 4133 3927 4147
rect 4033 4193 4047 4207
rect 3973 4173 3987 4187
rect 4073 4193 4087 4207
rect 4053 4153 4067 4167
rect 4013 4133 4027 4147
rect 3913 4053 3927 4067
rect 3933 4053 3947 4067
rect 4013 4013 4027 4027
rect 3993 3993 4007 4007
rect 3793 3933 3807 3947
rect 3833 3933 3847 3947
rect 3973 3973 3987 3987
rect 4093 4173 4107 4187
rect 4193 4193 4207 4207
rect 4213 4173 4227 4187
rect 4133 4133 4147 4147
rect 4113 4113 4127 4127
rect 4093 4033 4107 4047
rect 4113 4013 4127 4027
rect 4053 3973 4067 3987
rect 3713 3793 3727 3807
rect 3693 3773 3707 3787
rect 3673 3753 3687 3767
rect 3533 3713 3547 3727
rect 3953 3913 3967 3927
rect 4033 3913 4047 3927
rect 4093 3913 4107 3927
rect 4213 4153 4227 4167
rect 4173 4133 4187 4147
rect 4213 4073 4227 4087
rect 4153 4013 4167 4027
rect 4273 4233 4287 4247
rect 4273 4193 4287 4207
rect 4253 4173 4267 4187
rect 4233 4053 4247 4067
rect 4233 4033 4247 4047
rect 4153 3993 4167 4007
rect 4173 3973 4187 3987
rect 4253 3993 4267 4007
rect 3973 3853 3987 3867
rect 4113 3853 4127 3867
rect 3833 3793 3847 3807
rect 3793 3753 3807 3767
rect 3733 3733 3747 3747
rect 3753 3713 3767 3727
rect 3773 3673 3787 3687
rect 3553 3613 3567 3627
rect 3713 3613 3727 3627
rect 3713 3593 3727 3607
rect 3493 3513 3507 3527
rect 3513 3453 3527 3467
rect 3433 3373 3447 3387
rect 3473 3373 3487 3387
rect 3413 3273 3427 3287
rect 3293 3233 3307 3247
rect 3353 3213 3367 3227
rect 3393 3233 3407 3247
rect 3333 3153 3347 3167
rect 3153 3093 3167 3107
rect 3273 3093 3287 3107
rect 3293 3093 3307 3107
rect 2853 3033 2867 3047
rect 2853 3013 2867 3027
rect 2893 3013 2907 3027
rect 2933 3013 2947 3027
rect 2973 3033 2987 3047
rect 3093 3033 3107 3047
rect 3133 3033 3147 3047
rect 3153 3033 3167 3047
rect 2793 2993 2807 3007
rect 2873 2993 2887 3007
rect 2773 2973 2787 2987
rect 2733 2693 2747 2707
rect 2753 2693 2767 2707
rect 2813 2873 2827 2887
rect 2933 2973 2947 2987
rect 2893 2853 2907 2867
rect 2913 2853 2927 2867
rect 2913 2813 2927 2827
rect 2993 3013 3007 3027
rect 2973 2833 2987 2847
rect 3033 3013 3047 3027
rect 3073 3013 3087 3027
rect 3053 2993 3067 3007
rect 3013 2973 3027 2987
rect 3113 2993 3127 3007
rect 3133 3013 3147 3027
rect 3193 3013 3207 3027
rect 3233 3013 3247 3027
rect 3253 3033 3267 3047
rect 3333 3133 3347 3147
rect 3453 3213 3467 3227
rect 3493 3213 3507 3227
rect 3653 3553 3667 3567
rect 3573 3513 3587 3527
rect 3613 3513 3627 3527
rect 3673 3493 3687 3507
rect 3633 3453 3647 3467
rect 3693 3433 3707 3447
rect 3573 3393 3587 3407
rect 3693 3393 3707 3407
rect 3593 3293 3607 3307
rect 3553 3253 3567 3267
rect 3733 3513 3747 3527
rect 3773 3513 3787 3527
rect 3693 3253 3707 3267
rect 3713 3253 3727 3267
rect 3773 3273 3787 3287
rect 3573 3233 3587 3247
rect 3453 3193 3467 3207
rect 3473 3193 3487 3207
rect 3513 3193 3527 3207
rect 3373 3153 3387 3167
rect 3393 3153 3407 3167
rect 3453 3153 3467 3167
rect 3473 3153 3487 3167
rect 3413 3133 3427 3147
rect 3373 3053 3387 3067
rect 3493 3093 3507 3107
rect 3273 2993 3287 3007
rect 3353 3033 3367 3047
rect 3433 3033 3447 3047
rect 3333 2993 3347 3007
rect 3453 3013 3467 3027
rect 3553 3133 3567 3147
rect 3533 3053 3547 3067
rect 3593 3033 3607 3047
rect 3573 2993 3587 3007
rect 3593 2993 3607 3007
rect 3073 2973 3087 2987
rect 3093 2973 3107 2987
rect 3153 2973 3167 2987
rect 3313 2973 3327 2987
rect 3053 2953 3067 2967
rect 3053 2913 3067 2927
rect 3213 2953 3227 2967
rect 3293 2953 3307 2967
rect 3193 2933 3207 2947
rect 3073 2873 3087 2887
rect 3013 2853 3027 2867
rect 3113 2853 3127 2867
rect 2993 2793 3007 2807
rect 2873 2773 2887 2787
rect 2893 2773 2907 2787
rect 2933 2773 2947 2787
rect 2953 2773 2967 2787
rect 2813 2733 2827 2747
rect 2853 2733 2867 2747
rect 2873 2753 2887 2767
rect 2913 2753 2927 2767
rect 3033 2813 3047 2827
rect 3053 2813 3067 2827
rect 2893 2733 2907 2747
rect 2913 2733 2927 2747
rect 2953 2733 2967 2747
rect 2853 2713 2867 2727
rect 2873 2713 2887 2727
rect 2753 2633 2767 2647
rect 2793 2633 2807 2647
rect 2773 2613 2787 2627
rect 2753 2593 2767 2607
rect 2813 2613 2827 2627
rect 2813 2593 2827 2607
rect 2753 2573 2767 2587
rect 2773 2573 2787 2587
rect 2713 2553 2727 2567
rect 2693 2513 2707 2527
rect 2693 2493 2707 2507
rect 2773 2553 2787 2567
rect 2893 2693 2907 2707
rect 2873 2633 2887 2647
rect 2893 2633 2907 2647
rect 2893 2593 2907 2607
rect 2833 2553 2847 2567
rect 2773 2513 2787 2527
rect 2673 2453 2687 2467
rect 2653 2373 2667 2387
rect 2653 2313 2667 2327
rect 2633 2293 2647 2307
rect 2653 2293 2667 2307
rect 2553 2273 2567 2287
rect 2713 2413 2727 2427
rect 2693 2393 2707 2407
rect 2873 2533 2887 2547
rect 2833 2473 2847 2487
rect 2793 2453 2807 2467
rect 2773 2313 2787 2327
rect 2693 2293 2707 2307
rect 2513 2193 2527 2207
rect 2473 2173 2487 2187
rect 2513 2153 2527 2167
rect 2453 2133 2467 2147
rect 2553 2253 2567 2267
rect 2673 2273 2687 2287
rect 2533 2133 2547 2147
rect 2413 2053 2427 2067
rect 2493 2073 2507 2087
rect 2433 2033 2447 2047
rect 2393 1993 2407 2007
rect 2393 1953 2407 1967
rect 2333 1913 2347 1927
rect 2373 1913 2387 1927
rect 2293 1833 2307 1847
rect 2313 1833 2327 1847
rect 2293 1773 2307 1787
rect 2293 1713 2307 1727
rect 2273 1693 2287 1707
rect 2413 1913 2427 1927
rect 2393 1873 2407 1887
rect 2533 2033 2547 2047
rect 2493 1953 2507 1967
rect 2473 1913 2487 1927
rect 2453 1873 2467 1887
rect 2433 1853 2447 1867
rect 2373 1773 2387 1787
rect 2433 1793 2447 1807
rect 2453 1793 2467 1807
rect 2373 1753 2387 1767
rect 2433 1753 2447 1767
rect 2413 1733 2427 1747
rect 2353 1653 2367 1667
rect 2233 1633 2247 1647
rect 2273 1633 2287 1647
rect 2313 1633 2327 1647
rect 2373 1633 2387 1647
rect 2013 1593 2027 1607
rect 2193 1613 2207 1627
rect 2093 1573 2107 1587
rect 2213 1593 2227 1607
rect 2233 1573 2247 1587
rect 2353 1613 2367 1627
rect 1993 1533 2007 1547
rect 1973 1473 1987 1487
rect 1933 1353 1947 1367
rect 1833 1333 1847 1347
rect 1873 1333 1887 1347
rect 1893 1313 1907 1327
rect 2153 1533 2167 1547
rect 2053 1453 2067 1467
rect 1993 1373 2007 1387
rect 2073 1373 2087 1387
rect 2053 1353 2067 1367
rect 1973 1333 1987 1347
rect 2273 1513 2287 1527
rect 2293 1513 2307 1527
rect 2213 1453 2227 1467
rect 2173 1413 2187 1427
rect 2233 1433 2247 1447
rect 2333 1453 2347 1467
rect 2313 1433 2327 1447
rect 2293 1413 2307 1427
rect 2233 1393 2247 1407
rect 2253 1393 2267 1407
rect 2233 1373 2247 1387
rect 2113 1353 2127 1367
rect 2153 1353 2167 1367
rect 2193 1353 2207 1367
rect 2213 1353 2227 1367
rect 2173 1333 2187 1347
rect 1953 1313 1967 1327
rect 1833 1273 1847 1287
rect 1833 1253 1847 1267
rect 1793 1233 1807 1247
rect 1813 1233 1827 1247
rect 1773 1213 1787 1227
rect 1753 1193 1767 1207
rect 1813 1193 1827 1207
rect 1793 1133 1807 1147
rect 1933 1253 1947 1267
rect 1873 1153 1887 1167
rect 1913 1153 1927 1167
rect 1893 1133 1907 1147
rect 1833 1093 1847 1107
rect 1873 1093 1887 1107
rect 1793 1053 1807 1067
rect 1693 973 1707 987
rect 1633 813 1647 827
rect 1593 773 1607 787
rect 1753 853 1767 867
rect 1973 1293 1987 1307
rect 2073 1313 2087 1327
rect 2093 1293 2107 1307
rect 2153 1313 2167 1327
rect 2213 1313 2227 1327
rect 1993 1273 2007 1287
rect 2013 1273 2027 1287
rect 1953 1193 1967 1207
rect 1953 1153 1967 1167
rect 1933 1113 1947 1127
rect 1933 1093 1947 1107
rect 1913 1073 1927 1087
rect 2033 1253 2047 1267
rect 2053 1233 2067 1247
rect 2033 1193 2047 1207
rect 2113 1173 2127 1187
rect 2093 1153 2107 1167
rect 2173 1193 2187 1207
rect 2033 1133 2047 1147
rect 2053 1133 2067 1147
rect 2093 1133 2107 1147
rect 2113 1133 2127 1147
rect 2153 1133 2167 1147
rect 2053 1113 2067 1127
rect 1873 1033 1887 1047
rect 1893 973 1907 987
rect 1833 933 1847 947
rect 1873 933 1887 947
rect 1873 853 1887 867
rect 1693 813 1707 827
rect 1733 793 1747 807
rect 1813 793 1827 807
rect 1913 933 1927 947
rect 1973 833 1987 847
rect 2013 993 2027 1007
rect 2013 973 2027 987
rect 2033 973 2047 987
rect 2293 1373 2307 1387
rect 2273 1333 2287 1347
rect 2293 1333 2307 1347
rect 2353 1433 2367 1447
rect 2353 1293 2367 1307
rect 2293 1253 2307 1267
rect 2313 1253 2327 1267
rect 2253 1193 2267 1207
rect 2333 1193 2347 1207
rect 2573 2113 2587 2127
rect 2553 1953 2567 1967
rect 2693 2253 2707 2267
rect 2753 2253 2767 2267
rect 2613 2233 2627 2247
rect 2653 2233 2667 2247
rect 2693 2233 2707 2247
rect 2693 2213 2707 2227
rect 2733 2213 2747 2227
rect 2653 2153 2667 2167
rect 2613 2133 2627 2147
rect 2593 2073 2607 2087
rect 2633 2113 2647 2127
rect 2593 2033 2607 2047
rect 2713 2133 2727 2147
rect 2653 2073 2667 2087
rect 2673 2053 2687 2067
rect 2633 2033 2647 2047
rect 2673 2013 2687 2027
rect 2593 1993 2607 2007
rect 2633 1993 2647 2007
rect 2573 1933 2587 1947
rect 2573 1913 2587 1927
rect 2533 1853 2547 1867
rect 2493 1813 2507 1827
rect 2493 1773 2507 1787
rect 2533 1753 2547 1767
rect 2533 1713 2547 1727
rect 2553 1713 2567 1727
rect 2513 1653 2527 1667
rect 2473 1633 2487 1647
rect 2593 1773 2607 1787
rect 2593 1733 2607 1747
rect 2673 1953 2687 1967
rect 2653 1873 2667 1887
rect 2633 1753 2647 1767
rect 2573 1653 2587 1667
rect 2393 1613 2407 1627
rect 2453 1613 2467 1627
rect 2553 1613 2567 1627
rect 2413 1593 2427 1607
rect 2553 1593 2567 1607
rect 2613 1693 2627 1707
rect 2573 1573 2587 1587
rect 2473 1533 2487 1547
rect 2513 1533 2527 1547
rect 2453 1413 2467 1427
rect 2393 1333 2407 1347
rect 2413 1293 2427 1307
rect 2433 1313 2447 1327
rect 2393 1273 2407 1287
rect 2373 1233 2387 1247
rect 2433 1213 2447 1227
rect 2213 1133 2227 1147
rect 2313 1133 2327 1147
rect 2253 1113 2267 1127
rect 2293 1113 2307 1127
rect 2193 1053 2207 1067
rect 2313 1073 2327 1087
rect 2273 1033 2287 1047
rect 2153 973 2167 987
rect 2233 973 2247 987
rect 2113 873 2127 887
rect 2033 833 2047 847
rect 1953 813 1967 827
rect 1993 813 2007 827
rect 1553 693 1567 707
rect 1473 673 1487 687
rect 1473 633 1487 647
rect 1393 393 1407 407
rect 1453 393 1467 407
rect 1433 373 1447 387
rect 1553 653 1567 667
rect 1833 773 1847 787
rect 1693 673 1707 687
rect 1533 573 1547 587
rect 1673 593 1687 607
rect 1473 373 1487 387
rect 1273 333 1287 347
rect 1293 333 1307 347
rect 1213 233 1227 247
rect 1213 213 1227 227
rect 1173 173 1187 187
rect 1473 333 1487 347
rect 1393 293 1407 307
rect 1333 213 1347 227
rect 1253 193 1267 207
rect 1173 153 1187 167
rect 1153 133 1167 147
rect 1193 133 1207 147
rect 993 13 1007 27
rect 1033 13 1047 27
rect 1353 173 1367 187
rect 1313 153 1327 167
rect 1493 313 1507 327
rect 1433 193 1447 207
rect 1553 373 1567 387
rect 1613 373 1627 387
rect 1633 333 1647 347
rect 1553 313 1567 327
rect 1533 233 1547 247
rect 1453 173 1467 187
rect 1513 173 1527 187
rect 2093 793 2107 807
rect 2073 773 2087 787
rect 1873 753 1887 767
rect 1853 733 1867 747
rect 1793 633 1807 647
rect 1693 453 1707 467
rect 1673 333 1687 347
rect 1613 313 1627 327
rect 1653 313 1667 327
rect 1593 213 1607 227
rect 1553 173 1567 187
rect 1533 153 1547 167
rect 1593 153 1607 167
rect 1493 133 1507 147
rect 1533 113 1547 127
rect 1553 133 1567 147
rect 1753 413 1767 427
rect 2093 753 2107 767
rect 2173 953 2187 967
rect 2013 593 2027 607
rect 2093 593 2107 607
rect 2153 673 2167 687
rect 1893 393 1907 407
rect 2133 393 2147 407
rect 2293 913 2307 927
rect 2253 853 2267 867
rect 2193 773 2207 787
rect 2213 773 2227 787
rect 2193 393 2207 407
rect 2253 593 2267 607
rect 2393 1133 2407 1147
rect 2433 1133 2447 1147
rect 2373 953 2387 967
rect 2333 893 2347 907
rect 2493 1353 2507 1367
rect 2473 1273 2487 1287
rect 2473 1253 2487 1267
rect 2573 1473 2587 1487
rect 2693 1913 2707 1927
rect 2773 2193 2787 2207
rect 2753 2093 2767 2107
rect 2753 2073 2767 2087
rect 2733 1973 2747 1987
rect 2733 1873 2747 1887
rect 2713 1813 2727 1827
rect 2693 1753 2707 1767
rect 2673 1733 2687 1747
rect 2633 1653 2647 1667
rect 2653 1653 2667 1667
rect 2613 1393 2627 1407
rect 2673 1633 2687 1647
rect 2713 1733 2727 1747
rect 2953 2673 2967 2687
rect 3013 2713 3027 2727
rect 3073 2773 3087 2787
rect 3053 2673 3067 2687
rect 3073 2653 3087 2667
rect 2973 2633 2987 2647
rect 2993 2633 3007 2647
rect 2993 2573 3007 2587
rect 3033 2573 3047 2587
rect 2973 2553 2987 2567
rect 3053 2553 3067 2567
rect 2953 2513 2967 2527
rect 3133 2793 3147 2807
rect 3213 2733 3227 2747
rect 3193 2693 3207 2707
rect 3253 2773 3267 2787
rect 3313 2933 3327 2947
rect 3333 2933 3347 2947
rect 3313 2833 3327 2847
rect 3393 2933 3407 2947
rect 3533 2973 3547 2987
rect 3713 3233 3727 3247
rect 3633 3193 3647 3207
rect 3653 3193 3667 3207
rect 3673 3193 3687 3207
rect 3693 3193 3707 3207
rect 3753 3193 3767 3207
rect 3693 3093 3707 3107
rect 3633 3073 3647 3087
rect 3633 3053 3647 3067
rect 3613 2973 3627 2987
rect 3613 2953 3627 2967
rect 3573 2853 3587 2867
rect 3553 2833 3567 2847
rect 3413 2793 3427 2807
rect 3553 2793 3567 2807
rect 3293 2753 3307 2767
rect 3313 2753 3327 2767
rect 3253 2733 3267 2747
rect 3293 2713 3307 2727
rect 3313 2713 3327 2727
rect 3213 2673 3227 2687
rect 3213 2653 3227 2667
rect 3233 2653 3247 2667
rect 3113 2593 3127 2607
rect 3133 2593 3147 2607
rect 3093 2533 3107 2547
rect 2953 2493 2967 2507
rect 2933 2453 2947 2467
rect 2893 2413 2907 2427
rect 2873 2353 2887 2367
rect 2833 2333 2847 2347
rect 2873 2333 2887 2347
rect 2853 2253 2867 2267
rect 2833 2213 2847 2227
rect 2933 2333 2947 2347
rect 2893 2293 2907 2307
rect 2893 2253 2907 2267
rect 2933 2273 2947 2287
rect 2933 2233 2947 2247
rect 2873 2173 2887 2187
rect 2813 2113 2827 2127
rect 2913 2113 2927 2127
rect 2973 2393 2987 2407
rect 2993 2373 3007 2387
rect 2973 2293 2987 2307
rect 2953 2213 2967 2227
rect 3073 2513 3087 2527
rect 3113 2473 3127 2487
rect 3033 2433 3047 2447
rect 3093 2433 3107 2447
rect 3013 2293 3027 2307
rect 3013 2253 3027 2267
rect 3033 2213 3047 2227
rect 3073 2293 3087 2307
rect 3213 2613 3227 2627
rect 3213 2553 3227 2567
rect 3233 2473 3247 2487
rect 3173 2433 3187 2447
rect 3353 2733 3367 2747
rect 3413 2753 3427 2767
rect 3453 2753 3467 2767
rect 3353 2713 3367 2727
rect 3373 2693 3387 2707
rect 3393 2693 3407 2707
rect 3433 2693 3447 2707
rect 3453 2693 3467 2707
rect 3373 2633 3387 2647
rect 3333 2413 3347 2427
rect 3153 2373 3167 2387
rect 3173 2373 3187 2387
rect 3293 2373 3307 2387
rect 3133 2353 3147 2367
rect 3213 2333 3227 2347
rect 3173 2273 3187 2287
rect 3193 2273 3207 2287
rect 3153 2253 3167 2267
rect 3113 2193 3127 2207
rect 3193 2193 3207 2207
rect 3173 2173 3187 2187
rect 3093 2153 3107 2167
rect 3133 2153 3147 2167
rect 2993 2133 3007 2147
rect 3113 2133 3127 2147
rect 2973 2113 2987 2127
rect 2853 2093 2867 2107
rect 2933 2093 2947 2107
rect 3313 2313 3327 2327
rect 3233 2253 3247 2267
rect 3253 2273 3267 2287
rect 3313 2253 3327 2267
rect 3273 2213 3287 2227
rect 3413 2673 3427 2687
rect 3953 3773 3967 3787
rect 4393 4473 4407 4487
rect 4433 4473 4447 4487
rect 4393 4433 4407 4447
rect 4413 4413 4427 4427
rect 4373 4313 4387 4327
rect 4393 4313 4407 4327
rect 4353 4113 4367 4127
rect 4333 4053 4347 4067
rect 4313 3973 4327 3987
rect 4473 4473 4487 4487
rect 4593 4553 4607 4567
rect 4573 4513 4587 4527
rect 4573 4493 4587 4507
rect 4533 4453 4547 4467
rect 4553 4453 4567 4467
rect 4493 4433 4507 4447
rect 4633 4493 4647 4507
rect 4593 4473 4607 4487
rect 4613 4473 4627 4487
rect 4593 4453 4607 4467
rect 4693 4693 4707 4707
rect 4753 4793 4767 4807
rect 4813 4953 4827 4967
rect 4833 4953 4847 4967
rect 4813 4913 4827 4927
rect 4833 4893 4847 4907
rect 4833 4833 4847 4847
rect 4873 5033 4887 5047
rect 4893 5033 4907 5047
rect 4893 4993 4907 5007
rect 4933 4993 4947 5007
rect 4873 4953 4887 4967
rect 4893 4953 4907 4967
rect 4873 4813 4887 4827
rect 4833 4793 4847 4807
rect 4813 4733 4827 4747
rect 4793 4713 4807 4727
rect 4673 4673 4687 4687
rect 4693 4673 4707 4687
rect 4713 4673 4727 4687
rect 4733 4653 4747 4667
rect 4753 4673 4767 4687
rect 4793 4653 4807 4667
rect 4693 4633 4707 4647
rect 4733 4633 4747 4647
rect 4673 4613 4687 4627
rect 4713 4613 4727 4627
rect 4693 4533 4707 4547
rect 4693 4493 4707 4507
rect 4753 4613 4767 4627
rect 4793 4633 4807 4647
rect 4773 4593 4787 4607
rect 4753 4533 4767 4547
rect 4753 4513 4767 4527
rect 4733 4493 4747 4507
rect 4793 4493 4807 4507
rect 4633 4413 4647 4427
rect 4453 4393 4467 4407
rect 4573 4353 4587 4367
rect 4433 4333 4447 4347
rect 4373 4013 4387 4027
rect 4313 3953 4327 3967
rect 4353 3953 4367 3967
rect 4393 3973 4407 3987
rect 4473 4213 4487 4227
rect 4513 4153 4527 4167
rect 4553 4173 4567 4187
rect 4473 4033 4487 4047
rect 4453 3973 4467 3987
rect 4433 3953 4447 3967
rect 4493 3953 4507 3967
rect 4293 3793 4307 3807
rect 3873 3713 3887 3727
rect 3933 3713 3947 3727
rect 3953 3713 3967 3727
rect 3993 3713 4007 3727
rect 3913 3673 3927 3687
rect 3913 3613 3927 3627
rect 3893 3593 3907 3607
rect 3773 3053 3787 3067
rect 3833 3253 3847 3267
rect 3853 3253 3867 3267
rect 3893 3213 3907 3227
rect 3633 2933 3647 2947
rect 3713 2933 3727 2947
rect 3653 2893 3667 2907
rect 3773 2973 3787 2987
rect 3753 2873 3767 2887
rect 3573 2733 3587 2747
rect 3733 2733 3747 2747
rect 3573 2713 3587 2727
rect 3513 2693 3527 2707
rect 3553 2693 3567 2707
rect 3613 2693 3627 2707
rect 3593 2673 3607 2687
rect 3413 2613 3427 2627
rect 3473 2613 3487 2627
rect 3593 2593 3607 2607
rect 3533 2573 3547 2587
rect 3593 2573 3607 2587
rect 3453 2553 3467 2567
rect 3393 2533 3407 2547
rect 3433 2533 3447 2547
rect 3373 2473 3387 2487
rect 3353 2293 3367 2307
rect 3573 2553 3587 2567
rect 3493 2533 3507 2547
rect 3553 2533 3567 2547
rect 3533 2513 3547 2527
rect 3553 2513 3567 2527
rect 3453 2493 3467 2507
rect 3493 2493 3507 2507
rect 3513 2493 3527 2507
rect 3453 2473 3467 2487
rect 3473 2473 3487 2487
rect 3393 2413 3407 2427
rect 3373 2273 3387 2287
rect 3353 2253 3367 2267
rect 3473 2413 3487 2427
rect 3493 2413 3507 2427
rect 3473 2333 3487 2347
rect 3673 2713 3687 2727
rect 3653 2693 3667 2707
rect 3633 2593 3647 2607
rect 3713 2713 3727 2727
rect 3693 2613 3707 2627
rect 3613 2553 3627 2567
rect 3673 2573 3687 2587
rect 3673 2553 3687 2567
rect 3633 2533 3647 2547
rect 3673 2533 3687 2547
rect 3693 2533 3707 2547
rect 3673 2513 3687 2527
rect 3733 2693 3747 2707
rect 3753 2693 3767 2707
rect 3853 3033 3867 3047
rect 3813 3013 3827 3027
rect 3813 2973 3827 2987
rect 3813 2813 3827 2827
rect 3793 2793 3807 2807
rect 4073 3733 4087 3747
rect 4173 3733 4187 3747
rect 4113 3713 4127 3727
rect 4093 3693 4107 3707
rect 4053 3593 4067 3607
rect 3953 3553 3967 3567
rect 3993 3553 4007 3567
rect 4013 3553 4027 3567
rect 4033 3553 4047 3567
rect 3973 3493 3987 3507
rect 3993 3493 4007 3507
rect 4153 3513 4167 3527
rect 4133 3493 4147 3507
rect 3953 3413 3967 3427
rect 3953 3293 3967 3307
rect 4233 3693 4247 3707
rect 4293 3553 4307 3567
rect 4273 3493 4287 3507
rect 4373 3933 4387 3947
rect 4493 3893 4507 3907
rect 4473 3753 4487 3767
rect 4533 3753 4547 3767
rect 4413 3713 4427 3727
rect 4353 3693 4367 3707
rect 4373 3693 4387 3707
rect 4453 3593 4467 3607
rect 4373 3553 4387 3567
rect 4353 3533 4367 3547
rect 4373 3513 4387 3527
rect 4353 3493 4367 3507
rect 4333 3473 4347 3487
rect 4313 3453 4327 3467
rect 3933 3213 3947 3227
rect 4053 3233 4067 3247
rect 3933 3193 3947 3207
rect 3913 3093 3927 3107
rect 3893 3053 3907 3067
rect 4013 3193 4027 3207
rect 4093 3233 4107 3247
rect 4113 3213 4127 3227
rect 4173 3233 4187 3247
rect 4073 3193 4087 3207
rect 4393 3493 4407 3507
rect 4373 3453 4387 3467
rect 4593 4153 4607 4167
rect 4613 4033 4627 4047
rect 4773 4473 4787 4487
rect 4713 4433 4727 4447
rect 4713 4393 4727 4407
rect 4753 4433 4767 4447
rect 4733 4373 4747 4387
rect 4693 4313 4707 4327
rect 4673 4253 4687 4267
rect 4673 4233 4687 4247
rect 4773 4373 4787 4387
rect 4793 4333 4807 4347
rect 4773 4273 4787 4287
rect 4753 4213 4767 4227
rect 4693 4173 4707 4187
rect 4673 3993 4687 4007
rect 4733 3993 4747 4007
rect 4733 3933 4747 3947
rect 4713 3873 4727 3887
rect 4593 3793 4607 3807
rect 4593 3753 4607 3767
rect 4493 3733 4507 3747
rect 4513 3713 4527 3727
rect 4553 3733 4567 3747
rect 4473 3453 4487 3467
rect 4413 3373 4427 3387
rect 4713 3733 4727 3747
rect 4613 3533 4627 3547
rect 4513 3473 4527 3487
rect 3973 3093 3987 3107
rect 4053 3093 4067 3107
rect 3973 3013 3987 3027
rect 3793 2773 3807 2787
rect 3853 2773 3867 2787
rect 3773 2593 3787 2607
rect 3713 2513 3727 2527
rect 3573 2393 3587 2407
rect 3553 2373 3567 2387
rect 3553 2333 3567 2347
rect 3533 2293 3547 2307
rect 3473 2273 3487 2287
rect 3413 2253 3427 2267
rect 3413 2233 3427 2247
rect 3453 2233 3467 2247
rect 3353 2173 3367 2187
rect 3213 2133 3227 2147
rect 3293 2133 3307 2147
rect 3333 2133 3347 2147
rect 2833 2053 2847 2067
rect 2813 1953 2827 1967
rect 2793 1893 2807 1907
rect 2773 1853 2787 1867
rect 2773 1833 2787 1847
rect 2873 2073 2887 2087
rect 2973 2073 2987 2087
rect 2913 2053 2927 2067
rect 3013 2073 3027 2087
rect 2873 1973 2887 1987
rect 2853 1933 2867 1947
rect 2833 1913 2847 1927
rect 2833 1873 2847 1887
rect 2953 2013 2967 2027
rect 2993 2013 3007 2027
rect 3053 2033 3067 2047
rect 3033 1993 3047 2007
rect 3033 1933 3047 1947
rect 2893 1893 2907 1907
rect 2973 1873 2987 1887
rect 2873 1833 2887 1847
rect 2833 1813 2847 1827
rect 2853 1793 2867 1807
rect 3133 2093 3147 2107
rect 3113 2073 3127 2087
rect 3373 2153 3387 2167
rect 3393 2133 3407 2147
rect 3133 2053 3147 2067
rect 3153 2053 3167 2067
rect 3313 2053 3327 2067
rect 3353 2073 3367 2087
rect 3393 2053 3407 2067
rect 3113 2013 3127 2027
rect 3093 1953 3107 1967
rect 3113 1953 3127 1967
rect 3073 1873 3087 1887
rect 3053 1833 3067 1847
rect 2813 1773 2827 1787
rect 2893 1773 2907 1787
rect 2953 1773 2967 1787
rect 2993 1773 3007 1787
rect 3033 1793 3047 1807
rect 2793 1753 2807 1767
rect 2953 1753 2967 1767
rect 2973 1753 2987 1767
rect 2893 1733 2907 1747
rect 2733 1713 2747 1727
rect 2773 1713 2787 1727
rect 2773 1693 2787 1707
rect 2873 1693 2887 1707
rect 2693 1613 2707 1627
rect 2733 1613 2747 1627
rect 2813 1673 2827 1687
rect 2673 1593 2687 1607
rect 2773 1593 2787 1607
rect 2853 1613 2867 1627
rect 2793 1553 2807 1567
rect 2653 1413 2667 1427
rect 2633 1353 2647 1367
rect 2593 1333 2607 1347
rect 2713 1353 2727 1367
rect 2793 1533 2807 1547
rect 2913 1633 2927 1647
rect 3053 1773 3067 1787
rect 3013 1713 3027 1727
rect 2973 1693 2987 1707
rect 2953 1533 2967 1547
rect 2853 1513 2867 1527
rect 2893 1493 2907 1507
rect 2753 1413 2767 1427
rect 2853 1413 2867 1427
rect 2533 1293 2547 1307
rect 2733 1313 2747 1327
rect 2713 1293 2727 1307
rect 2553 1273 2567 1287
rect 2553 1233 2567 1247
rect 2573 1233 2587 1247
rect 2533 1193 2547 1207
rect 2513 1173 2527 1187
rect 2473 1133 2487 1147
rect 2473 1113 2487 1127
rect 2433 1013 2447 1027
rect 2453 1013 2467 1027
rect 2433 953 2447 967
rect 2513 1113 2527 1127
rect 2513 1093 2527 1107
rect 2513 993 2527 1007
rect 2553 1173 2567 1187
rect 2533 973 2547 987
rect 2413 913 2427 927
rect 2473 913 2487 927
rect 2533 913 2547 927
rect 2493 893 2507 907
rect 2373 853 2387 867
rect 2393 853 2407 867
rect 2413 853 2427 867
rect 2353 833 2367 847
rect 2373 833 2387 847
rect 2333 793 2347 807
rect 2393 813 2407 827
rect 2453 833 2467 847
rect 2393 793 2407 807
rect 2433 793 2447 807
rect 2313 773 2327 787
rect 2373 773 2387 787
rect 2473 753 2487 767
rect 2593 1133 2607 1147
rect 2713 1273 2727 1287
rect 2573 1093 2587 1107
rect 2613 1113 2627 1127
rect 2633 1093 2647 1107
rect 2653 1113 2667 1127
rect 2673 1113 2687 1127
rect 2673 1093 2687 1107
rect 2573 1073 2587 1087
rect 2653 1073 2667 1087
rect 2613 1033 2627 1047
rect 2553 893 2567 907
rect 2653 1013 2667 1027
rect 2593 873 2607 887
rect 2613 873 2627 887
rect 2533 833 2547 847
rect 2513 813 2527 827
rect 2573 813 2587 827
rect 2533 793 2547 807
rect 2553 793 2567 807
rect 2533 773 2547 787
rect 2513 713 2527 727
rect 2513 693 2527 707
rect 2313 593 2327 607
rect 2453 633 2467 647
rect 2233 513 2247 527
rect 2293 513 2307 527
rect 2093 373 2107 387
rect 2133 373 2147 387
rect 2173 373 2187 387
rect 2213 373 2227 387
rect 1713 273 1727 287
rect 1753 273 1767 287
rect 1773 273 1787 287
rect 1693 193 1707 207
rect 1753 193 1767 207
rect 1833 193 1847 207
rect 1913 193 1927 207
rect 1653 153 1667 167
rect 1633 133 1647 147
rect 1673 133 1687 147
rect 1733 133 1747 147
rect 1613 113 1627 127
rect 1793 173 1807 187
rect 1873 133 1887 147
rect 2013 353 2027 367
rect 2073 353 2087 367
rect 2093 333 2107 347
rect 2033 293 2047 307
rect 2053 213 2067 227
rect 2093 213 2107 227
rect 1973 173 1987 187
rect 1933 153 1947 167
rect 2013 153 2027 167
rect 2053 153 2067 167
rect 1953 133 1967 147
rect 2033 133 2047 147
rect 2013 113 2027 127
rect 2073 113 2087 127
rect 1593 93 1607 107
rect 2173 353 2187 367
rect 2193 353 2207 367
rect 2213 333 2227 347
rect 2233 353 2247 367
rect 2273 353 2287 367
rect 2293 333 2307 347
rect 2193 233 2207 247
rect 2113 93 2127 107
rect 2193 153 2207 167
rect 2253 273 2267 287
rect 2393 593 2407 607
rect 2493 673 2507 687
rect 2493 633 2507 647
rect 2493 473 2507 487
rect 2393 373 2407 387
rect 2333 353 2347 367
rect 2433 333 2447 347
rect 2573 753 2587 767
rect 2573 693 2587 707
rect 2613 833 2627 847
rect 2633 813 2647 827
rect 2653 833 2667 847
rect 2633 773 2647 787
rect 2673 773 2687 787
rect 2553 473 2567 487
rect 2353 313 2367 327
rect 2313 293 2327 307
rect 2333 293 2347 307
rect 2293 253 2307 267
rect 2233 173 2247 187
rect 2513 333 2527 347
rect 2433 313 2447 327
rect 2373 233 2387 247
rect 2353 213 2367 227
rect 2313 153 2327 167
rect 2333 153 2347 167
rect 2353 153 2367 167
rect 2353 113 2367 127
rect 2373 133 2387 147
rect 2413 133 2427 147
rect 2333 73 2347 87
rect 2453 253 2467 267
rect 2513 213 2527 227
rect 2473 133 2487 147
rect 2653 753 2667 767
rect 2633 653 2647 667
rect 2673 673 2687 687
rect 2733 1193 2747 1207
rect 2773 1273 2787 1287
rect 2813 1273 2827 1287
rect 2813 1233 2827 1247
rect 2853 1233 2867 1247
rect 2773 1213 2787 1227
rect 2773 1173 2787 1187
rect 2753 1153 2767 1167
rect 2853 1193 2867 1207
rect 2833 1153 2847 1167
rect 2813 1133 2827 1147
rect 2733 1073 2747 1087
rect 2793 1093 2807 1107
rect 2773 1073 2787 1087
rect 2753 1053 2767 1067
rect 2733 1013 2747 1027
rect 2713 953 2727 967
rect 2753 913 2767 927
rect 2733 753 2747 767
rect 2753 753 2767 767
rect 2813 1053 2827 1067
rect 2833 1033 2847 1047
rect 2873 1173 2887 1187
rect 3033 1693 3047 1707
rect 3033 1673 3047 1687
rect 3173 2033 3187 2047
rect 3233 2033 3247 2047
rect 3153 1873 3167 1887
rect 3133 1813 3147 1827
rect 3193 1913 3207 1927
rect 3173 1813 3187 1827
rect 3173 1793 3187 1807
rect 3333 1993 3347 2007
rect 3313 1933 3327 1947
rect 3233 1873 3247 1887
rect 3293 1873 3307 1887
rect 3273 1793 3287 1807
rect 3173 1753 3187 1767
rect 3193 1753 3207 1767
rect 3073 1713 3087 1727
rect 3133 1733 3147 1747
rect 3133 1693 3147 1707
rect 3113 1673 3127 1687
rect 3093 1653 3107 1667
rect 3033 1633 3047 1647
rect 3053 1633 3067 1647
rect 3053 1553 3067 1567
rect 3013 1473 3027 1487
rect 3053 1433 3067 1447
rect 3153 1673 3167 1687
rect 3253 1753 3267 1767
rect 3213 1713 3227 1727
rect 3313 1813 3327 1827
rect 3313 1753 3327 1767
rect 3453 2073 3467 2087
rect 3433 2013 3447 2027
rect 3393 1973 3407 1987
rect 3493 2253 3507 2267
rect 3493 2153 3507 2167
rect 3533 2153 3547 2167
rect 3473 2033 3487 2047
rect 3533 2113 3547 2127
rect 4033 3033 4047 3047
rect 3993 2953 4007 2967
rect 4013 2833 4027 2847
rect 3993 2813 4007 2827
rect 3993 2793 4007 2807
rect 3973 2773 3987 2787
rect 4013 2773 4027 2787
rect 4113 3033 4127 3047
rect 4073 2993 4087 3007
rect 4073 2793 4087 2807
rect 4153 2993 4167 3007
rect 4113 2953 4127 2967
rect 4093 2773 4107 2787
rect 3833 2753 3847 2767
rect 3933 2753 3947 2767
rect 3953 2753 3967 2767
rect 3893 2733 3907 2747
rect 3913 2733 3927 2747
rect 3993 2753 4007 2767
rect 3833 2713 3847 2727
rect 3813 2633 3827 2647
rect 3813 2553 3827 2567
rect 4073 2753 4087 2767
rect 3913 2693 3927 2707
rect 3953 2693 3967 2707
rect 3993 2713 4007 2727
rect 4073 2713 4087 2727
rect 3933 2593 3947 2607
rect 4233 3293 4247 3307
rect 4253 3213 4267 3227
rect 4393 3313 4407 3327
rect 4473 3313 4487 3327
rect 4613 3493 4627 3507
rect 4873 4713 4887 4727
rect 4853 4673 4867 4687
rect 4833 4653 4847 4667
rect 4873 4653 4887 4667
rect 4973 4953 4987 4967
rect 5033 5133 5047 5147
rect 5113 5273 5127 5287
rect 5153 5253 5167 5267
rect 5113 5213 5127 5227
rect 5093 5193 5107 5207
rect 5093 5153 5107 5167
rect 5113 5173 5127 5187
rect 5173 5233 5187 5247
rect 5513 5913 5527 5927
rect 5573 5913 5587 5927
rect 5473 5873 5487 5887
rect 5553 5893 5567 5907
rect 5453 5853 5467 5867
rect 5493 5853 5507 5867
rect 5433 5833 5447 5847
rect 5433 5753 5447 5767
rect 5353 5713 5367 5727
rect 5393 5713 5407 5727
rect 5413 5693 5427 5707
rect 5393 5673 5407 5687
rect 5253 5593 5267 5607
rect 5233 5573 5247 5587
rect 5233 5533 5247 5547
rect 5253 5533 5267 5547
rect 5213 5513 5227 5527
rect 5233 5453 5247 5467
rect 5353 5613 5367 5627
rect 5333 5573 5347 5587
rect 5313 5553 5327 5567
rect 5273 5513 5287 5527
rect 5273 5453 5287 5467
rect 5293 5453 5307 5467
rect 5273 5413 5287 5427
rect 5233 5393 5247 5407
rect 5253 5393 5267 5407
rect 5213 5333 5227 5347
rect 5093 5133 5107 5147
rect 5113 5133 5127 5147
rect 5013 4993 5027 5007
rect 5013 4953 5027 4967
rect 4973 4913 4987 4927
rect 4993 4893 5007 4907
rect 4913 4873 4927 4887
rect 4953 4873 4967 4887
rect 4973 4873 4987 4887
rect 5073 5093 5087 5107
rect 5053 4973 5067 4987
rect 5053 4913 5067 4927
rect 5033 4893 5047 4907
rect 5033 4873 5047 4887
rect 5053 4873 5067 4887
rect 5013 4813 5027 4827
rect 4953 4753 4967 4767
rect 4993 4753 5007 4767
rect 4973 4733 4987 4747
rect 4993 4733 5007 4747
rect 4913 4713 4927 4727
rect 5113 5033 5127 5047
rect 5093 4993 5107 5007
rect 5193 5193 5207 5207
rect 5193 5153 5207 5167
rect 5133 4973 5147 4987
rect 5093 4953 5107 4967
rect 5093 4913 5107 4927
rect 5133 4913 5147 4927
rect 5093 4893 5107 4907
rect 5113 4893 5127 4907
rect 5073 4813 5087 4827
rect 5173 5013 5187 5027
rect 5193 4993 5207 5007
rect 5173 4973 5187 4987
rect 5253 5273 5267 5287
rect 5233 5253 5247 5267
rect 5253 5193 5267 5207
rect 5273 5193 5287 5207
rect 5233 5173 5247 5187
rect 5233 5113 5247 5127
rect 5213 4973 5227 4987
rect 5173 4913 5187 4927
rect 5213 4913 5227 4927
rect 5273 5093 5287 5107
rect 5273 5073 5287 5087
rect 5253 4953 5267 4967
rect 5273 4953 5287 4967
rect 5253 4913 5267 4927
rect 5233 4873 5247 4887
rect 5153 4853 5167 4867
rect 5113 4833 5127 4847
rect 5193 4833 5207 4847
rect 5093 4793 5107 4807
rect 5093 4753 5107 4767
rect 5053 4733 5067 4747
rect 4913 4693 4927 4707
rect 4953 4693 4967 4707
rect 4973 4693 4987 4707
rect 5033 4693 5047 4707
rect 5053 4693 5067 4707
rect 5053 4673 5067 4687
rect 4833 4593 4847 4607
rect 4853 4573 4867 4587
rect 4853 4533 4867 4547
rect 4893 4533 4907 4547
rect 4873 4513 4887 4527
rect 4893 4493 4907 4507
rect 4833 4413 4847 4427
rect 4853 4413 4867 4427
rect 4893 4433 4907 4447
rect 4893 4373 4907 4387
rect 4933 4653 4947 4667
rect 4993 4653 5007 4667
rect 5193 4753 5207 4767
rect 5213 4753 5227 4767
rect 5173 4713 5187 4727
rect 5093 4693 5107 4707
rect 5113 4673 5127 4687
rect 5133 4693 5147 4707
rect 5153 4693 5167 4707
rect 5273 4893 5287 4907
rect 5393 5633 5407 5647
rect 5373 5593 5387 5607
rect 5393 5533 5407 5547
rect 5353 5513 5367 5527
rect 5393 5513 5407 5527
rect 5513 5813 5527 5827
rect 5673 6113 5687 6127
rect 5693 6133 5707 6147
rect 5713 6113 5727 6127
rect 5693 6073 5707 6087
rect 5653 6033 5667 6047
rect 5613 5993 5627 6007
rect 5673 5953 5687 5967
rect 5633 5933 5647 5947
rect 5653 5913 5667 5927
rect 5633 5893 5647 5907
rect 5813 6373 5827 6387
rect 5793 6353 5807 6367
rect 5913 6373 5927 6387
rect 5873 6353 5887 6367
rect 5913 6353 5927 6367
rect 5953 6353 5967 6367
rect 5813 6333 5827 6347
rect 5833 6333 5847 6347
rect 5753 6253 5767 6267
rect 5893 6233 5907 6247
rect 5813 6153 5827 6167
rect 5853 6133 5867 6147
rect 5773 6113 5787 6127
rect 5813 6113 5827 6127
rect 5833 6093 5847 6107
rect 5873 6113 5887 6127
rect 5793 6073 5807 6087
rect 5853 6073 5867 6087
rect 5753 6053 5767 6067
rect 5793 6033 5807 6047
rect 5713 5953 5727 5967
rect 5733 5953 5747 5967
rect 5693 5933 5707 5947
rect 5713 5933 5727 5947
rect 5773 5933 5787 5947
rect 5693 5893 5707 5907
rect 5753 5913 5767 5927
rect 5653 5873 5667 5887
rect 5693 5873 5707 5887
rect 5753 5873 5767 5887
rect 5573 5853 5587 5867
rect 5633 5853 5647 5867
rect 5533 5793 5547 5807
rect 5533 5773 5547 5787
rect 5513 5653 5527 5667
rect 5453 5633 5467 5647
rect 5493 5633 5507 5647
rect 5513 5613 5527 5627
rect 5573 5693 5587 5707
rect 5613 5793 5627 5807
rect 5553 5673 5567 5687
rect 5593 5673 5607 5687
rect 5593 5653 5607 5667
rect 5473 5593 5487 5607
rect 5493 5593 5507 5607
rect 5533 5593 5547 5607
rect 5453 5553 5467 5567
rect 5433 5473 5447 5487
rect 5413 5453 5427 5467
rect 5473 5533 5487 5547
rect 5333 5433 5347 5447
rect 5473 5413 5487 5427
rect 5373 5393 5387 5407
rect 5333 5353 5347 5367
rect 5333 5273 5347 5287
rect 5313 5253 5327 5267
rect 5393 5353 5407 5367
rect 5373 5253 5387 5267
rect 5353 5233 5367 5247
rect 5373 5193 5387 5207
rect 5333 5173 5347 5187
rect 5333 5153 5347 5167
rect 5373 5153 5387 5167
rect 5353 5113 5367 5127
rect 5373 5013 5387 5027
rect 5593 5613 5607 5627
rect 5573 5493 5587 5507
rect 5573 5453 5587 5467
rect 5533 5413 5547 5427
rect 5553 5393 5567 5407
rect 5473 5353 5487 5367
rect 5493 5353 5507 5367
rect 5653 5693 5667 5707
rect 5633 5673 5647 5687
rect 5833 5953 5847 5967
rect 6093 6433 6107 6447
rect 6133 6433 6147 6447
rect 5993 6373 6007 6387
rect 6033 6373 6047 6387
rect 6073 6353 6087 6367
rect 5973 6313 5987 6327
rect 5953 6153 5967 6167
rect 5973 6133 5987 6147
rect 5993 6113 6007 6127
rect 5973 6093 5987 6107
rect 5933 6073 5947 6087
rect 5933 6053 5947 6067
rect 5913 5973 5927 5987
rect 5873 5933 5887 5947
rect 5933 5933 5947 5947
rect 5973 5933 5987 5947
rect 5873 5913 5887 5927
rect 5893 5913 5907 5927
rect 5953 5893 5967 5907
rect 5773 5833 5787 5847
rect 5793 5833 5807 5847
rect 5833 5833 5847 5847
rect 5693 5653 5707 5667
rect 5753 5653 5767 5667
rect 5653 5593 5667 5607
rect 5633 5573 5647 5587
rect 5633 5533 5647 5547
rect 5653 5533 5667 5547
rect 5653 5513 5667 5527
rect 5693 5613 5707 5627
rect 5713 5613 5727 5627
rect 5733 5633 5747 5647
rect 5773 5633 5787 5647
rect 5773 5593 5787 5607
rect 5753 5573 5767 5587
rect 5713 5533 5727 5547
rect 5733 5533 5747 5547
rect 5693 5513 5707 5527
rect 5673 5493 5687 5507
rect 5673 5473 5687 5487
rect 5613 5453 5627 5467
rect 5653 5453 5667 5467
rect 5633 5413 5647 5427
rect 5673 5413 5687 5427
rect 5893 5833 5907 5847
rect 5853 5813 5867 5827
rect 6113 6333 6127 6347
rect 6093 6313 6107 6327
rect 6053 6153 6067 6167
rect 6253 6453 6267 6467
rect 6293 6453 6307 6467
rect 6353 6453 6367 6467
rect 6213 6433 6227 6447
rect 6233 6433 6247 6447
rect 6153 6373 6167 6387
rect 6353 6413 6367 6427
rect 6273 6373 6287 6387
rect 6333 6373 6347 6387
rect 6213 6353 6227 6367
rect 6233 6353 6247 6367
rect 6133 6273 6147 6287
rect 6173 6273 6187 6287
rect 6133 6233 6147 6247
rect 6133 6153 6147 6167
rect 6173 6153 6187 6167
rect 6193 6153 6207 6167
rect 6153 6133 6167 6147
rect 6173 6113 6187 6127
rect 6033 6073 6047 6087
rect 6073 6073 6087 6087
rect 6513 6433 6527 6447
rect 6533 6433 6547 6447
rect 6593 6433 6607 6447
rect 6693 6433 6707 6447
rect 6413 6413 6427 6427
rect 6373 6373 6387 6387
rect 6393 6353 6407 6367
rect 6313 6333 6327 6347
rect 6573 6413 6587 6427
rect 6433 6373 6447 6387
rect 6413 6333 6427 6347
rect 6473 6373 6487 6387
rect 6493 6353 6507 6367
rect 6433 6233 6447 6247
rect 6313 6173 6327 6187
rect 6233 6153 6247 6167
rect 6273 6153 6287 6167
rect 6253 6133 6267 6147
rect 6233 6113 6247 6127
rect 6253 6113 6267 6127
rect 6293 6133 6307 6147
rect 6153 6073 6167 6087
rect 6173 6073 6187 6087
rect 6153 6033 6167 6047
rect 6093 6013 6107 6027
rect 6033 5933 6047 5947
rect 6073 5933 6087 5947
rect 6133 5933 6147 5947
rect 6153 5933 6167 5947
rect 6173 5933 6187 5947
rect 6013 5913 6027 5927
rect 5973 5853 5987 5867
rect 5913 5813 5927 5827
rect 5973 5733 5987 5747
rect 5933 5713 5947 5727
rect 5893 5693 5907 5707
rect 5933 5693 5947 5707
rect 5953 5673 5967 5687
rect 5953 5653 5967 5667
rect 5873 5613 5887 5627
rect 5893 5633 5907 5647
rect 5933 5633 5947 5647
rect 5853 5593 5867 5607
rect 5873 5593 5887 5607
rect 6053 5893 6067 5907
rect 6093 5913 6107 5927
rect 6153 5893 6167 5907
rect 6093 5873 6107 5887
rect 6113 5873 6127 5887
rect 6093 5833 6107 5847
rect 6113 5753 6127 5767
rect 6013 5693 6027 5707
rect 6173 5693 6187 5707
rect 5993 5653 6007 5667
rect 6093 5673 6107 5687
rect 6053 5633 6067 5647
rect 6073 5613 6087 5627
rect 5953 5593 5967 5607
rect 5833 5573 5847 5587
rect 5793 5553 5807 5567
rect 5913 5573 5927 5587
rect 5793 5533 5807 5547
rect 5773 5493 5787 5507
rect 5793 5493 5807 5507
rect 5773 5473 5787 5487
rect 5753 5453 5767 5467
rect 5573 5373 5587 5387
rect 5653 5373 5667 5387
rect 5733 5373 5747 5387
rect 5553 5353 5567 5367
rect 5593 5353 5607 5367
rect 5513 5333 5527 5347
rect 5433 5313 5447 5327
rect 5473 5313 5487 5327
rect 5533 5313 5547 5327
rect 5513 5253 5527 5267
rect 5533 5253 5547 5267
rect 5513 5213 5527 5227
rect 5573 5233 5587 5247
rect 5433 5173 5447 5187
rect 5473 5173 5487 5187
rect 5533 5173 5547 5187
rect 5513 5153 5527 5167
rect 5413 5013 5427 5027
rect 5393 4993 5407 5007
rect 5333 4973 5347 4987
rect 5313 4953 5327 4967
rect 5353 4953 5367 4967
rect 5393 4953 5407 4967
rect 5473 5133 5487 5147
rect 5493 5133 5507 5147
rect 5453 4973 5467 4987
rect 5473 4973 5487 4987
rect 5573 5133 5587 5147
rect 5553 5093 5567 5107
rect 5553 5013 5567 5027
rect 5573 5013 5587 5027
rect 5553 4973 5567 4987
rect 5413 4933 5427 4947
rect 5433 4933 5447 4947
rect 5533 4953 5547 4967
rect 5353 4913 5367 4927
rect 5273 4853 5287 4867
rect 5293 4853 5307 4867
rect 5293 4793 5307 4807
rect 5253 4753 5267 4767
rect 5273 4753 5287 4767
rect 5253 4713 5267 4727
rect 5293 4713 5307 4727
rect 5333 4713 5347 4727
rect 5193 4693 5207 4707
rect 5233 4693 5247 4707
rect 4953 4513 4967 4527
rect 4973 4513 4987 4527
rect 5073 4653 5087 4667
rect 5033 4593 5047 4607
rect 5033 4573 5047 4587
rect 4993 4473 5007 4487
rect 5213 4673 5227 4687
rect 5233 4673 5247 4687
rect 5153 4633 5167 4647
rect 5233 4633 5247 4647
rect 5193 4613 5207 4627
rect 5413 4873 5427 4887
rect 5373 4813 5387 4827
rect 5453 4853 5467 4867
rect 5433 4833 5447 4847
rect 5413 4793 5427 4807
rect 5393 4713 5407 4727
rect 5273 4653 5287 4667
rect 5293 4673 5307 4687
rect 5393 4673 5407 4687
rect 5413 4693 5427 4707
rect 5373 4653 5387 4667
rect 5393 4653 5407 4667
rect 5433 4653 5447 4667
rect 5053 4553 5067 4567
rect 5093 4553 5107 4567
rect 4953 4453 4967 4467
rect 4993 4453 5007 4467
rect 4913 4273 4927 4287
rect 4853 4253 4867 4267
rect 4873 4253 4887 4267
rect 4973 4393 4987 4407
rect 5153 4533 5167 4547
rect 5133 4493 5147 4507
rect 5173 4493 5187 4507
rect 5093 4473 5107 4487
rect 5073 4453 5087 4467
rect 5153 4473 5167 4487
rect 5153 4453 5167 4467
rect 5093 4433 5107 4447
rect 4993 4353 5007 4367
rect 4953 4313 4967 4327
rect 4813 4233 4827 4247
rect 4833 4233 4847 4247
rect 4893 4213 4907 4227
rect 4993 4293 5007 4307
rect 4973 4273 4987 4287
rect 5053 4393 5067 4407
rect 4993 4253 5007 4267
rect 5013 4253 5027 4267
rect 5133 4433 5147 4447
rect 5093 4373 5107 4387
rect 5113 4373 5127 4387
rect 5133 4353 5147 4367
rect 5193 4453 5207 4467
rect 5193 4373 5207 4387
rect 5213 4353 5227 4367
rect 5133 4333 5147 4347
rect 5173 4333 5187 4347
rect 5093 4253 5107 4267
rect 5113 4253 5127 4267
rect 5053 4233 5067 4247
rect 5273 4593 5287 4607
rect 5333 4633 5347 4647
rect 5353 4613 5367 4627
rect 5333 4533 5347 4547
rect 5333 4513 5347 4527
rect 5433 4633 5447 4647
rect 5513 4913 5527 4927
rect 5493 4893 5507 4907
rect 5473 4813 5487 4827
rect 5613 5193 5627 5207
rect 5633 5173 5647 5187
rect 5633 5113 5647 5127
rect 5613 5093 5627 5107
rect 5593 4973 5607 4987
rect 5573 4953 5587 4967
rect 5733 5333 5747 5347
rect 5893 5493 5907 5507
rect 5933 5453 5947 5467
rect 5813 5433 5827 5447
rect 5833 5413 5847 5427
rect 5893 5433 5907 5447
rect 5913 5433 5927 5447
rect 5773 5393 5787 5407
rect 5753 5313 5767 5327
rect 5753 5213 5767 5227
rect 5733 5193 5747 5207
rect 5693 5173 5707 5187
rect 5693 5153 5707 5167
rect 5733 5173 5747 5187
rect 5673 5133 5687 5147
rect 5693 5113 5707 5127
rect 5693 5093 5707 5107
rect 5653 4973 5667 4987
rect 5633 4953 5647 4967
rect 5813 5353 5827 5367
rect 5793 5293 5807 5307
rect 5773 5173 5787 5187
rect 5813 5273 5827 5287
rect 5853 5273 5867 5287
rect 5833 5213 5847 5227
rect 5913 5393 5927 5407
rect 5993 5593 6007 5607
rect 6013 5593 6027 5607
rect 5993 5573 6007 5587
rect 5993 5513 6007 5527
rect 6013 5513 6027 5527
rect 6053 5593 6067 5607
rect 6053 5553 6067 5567
rect 6053 5533 6067 5547
rect 6033 5493 6047 5507
rect 5993 5453 6007 5467
rect 6113 5573 6127 5587
rect 6093 5513 6107 5527
rect 6073 5473 6087 5487
rect 6153 5613 6167 5627
rect 6173 5613 6187 5627
rect 6133 5553 6147 5567
rect 6133 5513 6147 5527
rect 6173 5513 6187 5527
rect 6153 5473 6167 5487
rect 6093 5453 6107 5467
rect 6133 5453 6147 5467
rect 6053 5433 6067 5447
rect 6073 5433 6087 5447
rect 6013 5393 6027 5407
rect 6053 5393 6067 5407
rect 5893 5353 5907 5367
rect 5933 5373 5947 5387
rect 5913 5333 5927 5347
rect 5993 5373 6007 5387
rect 5933 5293 5947 5307
rect 5953 5293 5967 5307
rect 5893 5253 5907 5267
rect 6013 5353 6027 5367
rect 5873 5233 5887 5247
rect 5893 5233 5907 5247
rect 5933 5233 5947 5247
rect 5973 5233 5987 5247
rect 5993 5233 6007 5247
rect 5873 5193 5887 5207
rect 5833 5153 5847 5167
rect 5993 5193 6007 5207
rect 6173 5453 6187 5467
rect 6093 5373 6107 5387
rect 6133 5393 6147 5407
rect 6113 5313 6127 5327
rect 6033 5293 6047 5307
rect 6073 5293 6087 5307
rect 6113 5293 6127 5307
rect 5913 5153 5927 5167
rect 5973 5173 5987 5187
rect 5993 5153 6007 5167
rect 5853 5133 5867 5147
rect 5873 5133 5887 5147
rect 5953 5133 5967 5147
rect 6013 5133 6027 5147
rect 5773 5093 5787 5107
rect 5813 5093 5827 5107
rect 5733 5073 5747 5087
rect 5753 5073 5767 5087
rect 5833 5073 5847 5087
rect 5713 4993 5727 5007
rect 5713 4973 5727 4987
rect 5633 4933 5647 4947
rect 5653 4913 5667 4927
rect 5573 4893 5587 4907
rect 5613 4893 5627 4907
rect 5633 4893 5647 4907
rect 5573 4873 5587 4887
rect 5613 4873 5627 4887
rect 5553 4833 5567 4847
rect 5593 4853 5607 4867
rect 5593 4773 5607 4787
rect 5573 4753 5587 4767
rect 5473 4733 5487 4747
rect 5513 4713 5527 4727
rect 5513 4693 5527 4707
rect 5553 4693 5567 4707
rect 5553 4673 5567 4687
rect 5593 4693 5607 4707
rect 5473 4653 5487 4667
rect 5433 4613 5447 4627
rect 5453 4613 5467 4627
rect 5253 4473 5267 4487
rect 5313 4493 5327 4507
rect 5353 4493 5367 4507
rect 5273 4453 5287 4467
rect 5353 4453 5367 4467
rect 5293 4433 5307 4447
rect 5413 4573 5427 4587
rect 5393 4533 5407 4547
rect 5413 4513 5427 4527
rect 5373 4433 5387 4447
rect 5273 4393 5287 4407
rect 5193 4233 5207 4247
rect 5233 4233 5247 4247
rect 4973 4213 4987 4227
rect 5033 4213 5047 4227
rect 4933 4173 4947 4187
rect 4973 4193 4987 4207
rect 4993 4193 5007 4207
rect 5053 4193 5067 4207
rect 5013 4173 5027 4187
rect 4973 4153 4987 4167
rect 5113 4213 5127 4227
rect 5133 4213 5147 4227
rect 5133 4193 5147 4207
rect 5193 4193 5207 4207
rect 5213 4173 5227 4187
rect 5113 4153 5127 4167
rect 5153 4153 5167 4167
rect 5093 4133 5107 4147
rect 4933 4113 4947 4127
rect 5173 4113 5187 4127
rect 4913 4053 4927 4067
rect 4853 3993 4867 4007
rect 4893 3993 4907 4007
rect 4773 3953 4787 3967
rect 4813 3973 4827 3987
rect 4793 3933 4807 3947
rect 4873 3973 4887 3987
rect 4913 3953 4927 3967
rect 4853 3873 4867 3887
rect 5033 3993 5047 4007
rect 4913 3833 4927 3847
rect 4753 3753 4767 3767
rect 4893 3753 4907 3767
rect 4953 3773 4967 3787
rect 4833 3693 4847 3707
rect 4653 3513 4667 3527
rect 4733 3533 4747 3547
rect 4713 3473 4727 3487
rect 5193 3993 5207 4007
rect 5153 3973 5167 3987
rect 5153 3773 5167 3787
rect 5093 3753 5107 3767
rect 5353 4413 5367 4427
rect 5333 4393 5347 4407
rect 5293 4193 5307 4207
rect 5273 4133 5287 4147
rect 5373 4373 5387 4387
rect 5353 4233 5367 4247
rect 5413 4433 5427 4447
rect 5413 4293 5427 4307
rect 5393 4213 5407 4227
rect 5353 4173 5367 4187
rect 5333 4153 5347 4167
rect 5253 4113 5267 4127
rect 5253 4093 5267 4107
rect 5293 4113 5307 4127
rect 5273 4053 5287 4067
rect 5353 4093 5367 4107
rect 5293 4013 5307 4027
rect 5293 3993 5307 4007
rect 5313 3993 5327 4007
rect 5273 3973 5287 3987
rect 5333 3953 5347 3967
rect 5233 3853 5247 3867
rect 5253 3853 5267 3867
rect 5273 3853 5287 3867
rect 5213 3793 5227 3807
rect 5253 3793 5267 3807
rect 5453 4533 5467 4547
rect 5453 4493 5467 4507
rect 5533 4633 5547 4647
rect 5493 4593 5507 4607
rect 5553 4573 5567 4587
rect 5593 4653 5607 4667
rect 5493 4533 5507 4547
rect 5473 4473 5487 4487
rect 5573 4553 5587 4567
rect 5573 4513 5587 4527
rect 5533 4493 5547 4507
rect 5593 4473 5607 4487
rect 5453 4433 5467 4447
rect 5513 4453 5527 4467
rect 5533 4453 5547 4467
rect 5513 4433 5527 4447
rect 5553 4433 5567 4447
rect 5653 4753 5667 4767
rect 5633 4713 5647 4727
rect 5713 4873 5727 4887
rect 5713 4793 5727 4807
rect 5693 4773 5707 4787
rect 5833 5033 5847 5047
rect 5793 4973 5807 4987
rect 5753 4953 5767 4967
rect 5793 4933 5807 4947
rect 5813 4933 5827 4947
rect 5753 4913 5767 4927
rect 5773 4893 5787 4907
rect 5753 4873 5767 4887
rect 5753 4833 5767 4847
rect 5773 4833 5787 4847
rect 5913 5113 5927 5127
rect 5933 5113 5947 5127
rect 5893 5073 5907 5087
rect 5853 5013 5867 5027
rect 5873 5013 5887 5027
rect 5853 4993 5867 5007
rect 5873 4973 5887 4987
rect 5873 4933 5887 4947
rect 5913 4993 5927 5007
rect 5913 4973 5927 4987
rect 5913 4933 5927 4947
rect 5813 4893 5827 4907
rect 5833 4893 5847 4907
rect 5873 4893 5887 4907
rect 5813 4813 5827 4827
rect 5793 4793 5807 4807
rect 5733 4753 5747 4767
rect 5753 4753 5767 4767
rect 5713 4733 5727 4747
rect 5673 4713 5687 4727
rect 5773 4713 5787 4727
rect 5693 4693 5707 4707
rect 5733 4693 5747 4707
rect 5733 4673 5747 4687
rect 5633 4633 5647 4647
rect 5653 4613 5667 4627
rect 5713 4653 5727 4667
rect 5713 4633 5727 4647
rect 5693 4613 5707 4627
rect 5673 4573 5687 4587
rect 5673 4533 5687 4547
rect 5653 4513 5667 4527
rect 5693 4453 5707 4467
rect 5453 4373 5467 4387
rect 5493 4413 5507 4427
rect 5533 4413 5547 4427
rect 5513 4353 5527 4367
rect 5493 4333 5507 4347
rect 5473 4293 5487 4307
rect 5473 4253 5487 4267
rect 5433 4193 5447 4207
rect 5413 4153 5427 4167
rect 5473 4173 5487 4187
rect 5453 4093 5467 4107
rect 5413 4053 5427 4067
rect 5593 4373 5607 4387
rect 5553 4333 5567 4347
rect 5573 4253 5587 4267
rect 5573 4213 5587 4227
rect 5633 4353 5647 4367
rect 5693 4393 5707 4407
rect 5653 4313 5667 4327
rect 5733 4613 5747 4627
rect 5773 4653 5787 4667
rect 5753 4573 5767 4587
rect 5793 4573 5807 4587
rect 5773 4513 5787 4527
rect 5733 4493 5747 4507
rect 5713 4333 5727 4347
rect 5753 4433 5767 4447
rect 5773 4453 5787 4467
rect 5793 4413 5807 4427
rect 5753 4373 5767 4387
rect 5733 4253 5747 4267
rect 5673 4233 5687 4247
rect 5693 4233 5707 4247
rect 5793 4333 5807 4347
rect 5793 4273 5807 4287
rect 5573 4193 5587 4207
rect 5613 4193 5627 4207
rect 5553 4173 5567 4187
rect 5513 4053 5527 4067
rect 5533 4053 5547 4067
rect 5493 4013 5507 4027
rect 5473 3973 5487 3987
rect 5493 3993 5507 4007
rect 5533 4013 5547 4027
rect 5793 4233 5807 4247
rect 5753 4213 5767 4227
rect 5793 4213 5807 4227
rect 5713 4173 5727 4187
rect 5733 4173 5747 4187
rect 5633 4153 5647 4167
rect 5593 4113 5607 4127
rect 5593 4013 5607 4027
rect 5553 3973 5567 3987
rect 5573 3953 5587 3967
rect 5493 3913 5507 3927
rect 5533 3913 5547 3927
rect 5433 3853 5447 3867
rect 5393 3773 5407 3787
rect 5373 3753 5387 3767
rect 5053 3713 5067 3727
rect 5033 3693 5047 3707
rect 5133 3713 5147 3727
rect 5153 3673 5167 3687
rect 4993 3593 5007 3607
rect 5093 3593 5107 3607
rect 4913 3533 4927 3547
rect 4893 3513 4907 3527
rect 4953 3513 4967 3527
rect 4753 3373 4767 3387
rect 4773 3373 4787 3387
rect 4713 3353 4727 3367
rect 4553 3313 4567 3327
rect 4713 3313 4727 3327
rect 4553 3273 4567 3287
rect 4593 3273 4607 3287
rect 4673 3273 4687 3287
rect 4413 3213 4427 3227
rect 4473 3233 4487 3247
rect 4533 3213 4547 3227
rect 4573 3213 4587 3227
rect 4433 3193 4447 3207
rect 4473 3193 4487 3207
rect 4493 3193 4507 3207
rect 4393 3133 4407 3147
rect 4433 3133 4447 3147
rect 4273 3113 4287 3127
rect 4253 3093 4267 3107
rect 4293 3093 4307 3107
rect 4413 3093 4427 3107
rect 4273 3053 4287 3067
rect 4293 3053 4307 3067
rect 4193 2993 4207 3007
rect 4213 3013 4227 3027
rect 4233 3013 4247 3027
rect 4233 2993 4247 3007
rect 4273 2973 4287 2987
rect 4173 2893 4187 2907
rect 4353 3033 4367 3047
rect 4333 2993 4347 3007
rect 4413 2993 4427 3007
rect 4173 2853 4187 2867
rect 4173 2793 4187 2807
rect 4133 2773 4147 2787
rect 4113 2713 4127 2727
rect 4093 2653 4107 2667
rect 4253 2773 4267 2787
rect 4313 2773 4327 2787
rect 4153 2733 4167 2747
rect 4213 2753 4227 2767
rect 4493 3133 4507 3147
rect 4613 3193 4627 3207
rect 4633 3193 4647 3207
rect 4493 3093 4507 3107
rect 4513 3093 4527 3107
rect 4593 3093 4607 3107
rect 4473 3073 4487 3087
rect 4493 3053 4507 3067
rect 4633 3093 4647 3107
rect 4573 3073 4587 3087
rect 4613 3073 4627 3087
rect 4613 3033 4627 3047
rect 4553 2973 4567 2987
rect 4533 2953 4547 2967
rect 4513 2913 4527 2927
rect 4493 2893 4507 2907
rect 4413 2813 4427 2827
rect 4433 2813 4447 2827
rect 4353 2773 4367 2787
rect 4333 2753 4347 2767
rect 4393 2753 4407 2767
rect 4413 2753 4427 2767
rect 4293 2733 4307 2747
rect 4353 2733 4367 2747
rect 4173 2713 4187 2727
rect 4213 2713 4227 2727
rect 4253 2713 4267 2727
rect 4053 2633 4067 2647
rect 4133 2633 4147 2647
rect 3993 2573 4007 2587
rect 4013 2573 4027 2587
rect 4033 2573 4047 2587
rect 3893 2553 3907 2567
rect 3793 2533 3807 2547
rect 3793 2513 3807 2527
rect 3873 2533 3887 2547
rect 4073 2593 4087 2607
rect 4013 2533 4027 2547
rect 4033 2533 4047 2547
rect 3853 2513 3867 2527
rect 3893 2513 3907 2527
rect 3993 2513 4007 2527
rect 3793 2493 3807 2507
rect 3673 2473 3687 2487
rect 3713 2473 3727 2487
rect 3773 2473 3787 2487
rect 3813 2473 3827 2487
rect 3593 2373 3607 2387
rect 3633 2313 3647 2327
rect 3653 2273 3667 2287
rect 3633 2213 3647 2227
rect 3573 2193 3587 2207
rect 3633 2193 3647 2207
rect 3573 2073 3587 2087
rect 3553 1953 3567 1967
rect 3513 1913 3527 1927
rect 3353 1893 3367 1907
rect 3393 1893 3407 1907
rect 3453 1893 3467 1907
rect 3573 1893 3587 1907
rect 3573 1873 3587 1887
rect 3513 1853 3527 1867
rect 3353 1833 3367 1847
rect 3393 1833 3407 1847
rect 3433 1813 3447 1827
rect 3513 1813 3527 1827
rect 3373 1753 3387 1767
rect 3333 1733 3347 1747
rect 3313 1713 3327 1727
rect 3293 1693 3307 1707
rect 3213 1613 3227 1627
rect 2973 1413 2987 1427
rect 2953 1393 2967 1407
rect 2953 1373 2967 1387
rect 2933 1333 2947 1347
rect 3133 1393 3147 1407
rect 3113 1353 3127 1367
rect 2973 1333 2987 1347
rect 2993 1333 3007 1347
rect 3073 1333 3087 1347
rect 2953 1313 2967 1327
rect 3013 1293 3027 1307
rect 3033 1313 3047 1327
rect 2953 1273 2967 1287
rect 3033 1273 3047 1287
rect 2973 1233 2987 1247
rect 2933 1213 2947 1227
rect 2873 1153 2887 1167
rect 2873 1133 2887 1147
rect 2913 1153 2927 1167
rect 2793 953 2807 967
rect 2793 833 2807 847
rect 2773 713 2787 727
rect 2733 693 2747 707
rect 2773 693 2787 707
rect 2713 613 2727 627
rect 2753 613 2767 627
rect 2773 633 2787 647
rect 2733 493 2747 507
rect 2673 313 2687 327
rect 2613 293 2627 307
rect 2653 293 2667 307
rect 2713 353 2727 367
rect 2833 973 2847 987
rect 2813 793 2827 807
rect 2853 933 2867 947
rect 2933 1053 2947 1067
rect 2933 853 2947 867
rect 2993 1113 3007 1127
rect 2993 1033 3007 1047
rect 3053 1233 3067 1247
rect 3053 1113 3067 1127
rect 3033 1033 3047 1047
rect 3093 1313 3107 1327
rect 3093 1133 3107 1147
rect 3233 1553 3247 1567
rect 3313 1633 3327 1647
rect 3373 1633 3387 1647
rect 3293 1553 3307 1567
rect 3393 1613 3407 1627
rect 3333 1553 3347 1567
rect 3353 1573 3367 1587
rect 3493 1773 3507 1787
rect 3473 1753 3487 1767
rect 3513 1753 3527 1767
rect 3653 2133 3667 2147
rect 3613 2093 3627 2107
rect 3773 2413 3787 2427
rect 3953 2493 3967 2507
rect 3833 2393 3847 2407
rect 3853 2393 3867 2407
rect 3893 2393 3907 2407
rect 3773 2293 3787 2307
rect 3793 2293 3807 2307
rect 3753 2253 3767 2267
rect 3833 2293 3847 2307
rect 3933 2333 3947 2347
rect 3893 2293 3907 2307
rect 3813 2253 3827 2267
rect 3713 2193 3727 2207
rect 3773 2193 3787 2207
rect 3773 2173 3787 2187
rect 3693 2153 3707 2167
rect 3713 2133 3727 2147
rect 3673 2073 3687 2087
rect 3733 2053 3747 2067
rect 3873 2253 3887 2267
rect 3893 2253 3907 2267
rect 3853 2153 3867 2167
rect 3833 2113 3847 2127
rect 3813 2093 3827 2107
rect 3933 2253 3947 2267
rect 3913 2213 3927 2227
rect 3893 2193 3907 2207
rect 3773 2053 3787 2067
rect 3813 2053 3827 2067
rect 3873 2073 3887 2087
rect 3653 2033 3667 2047
rect 3613 1993 3627 2007
rect 3673 2013 3687 2027
rect 3693 1993 3707 2007
rect 3673 1833 3687 1847
rect 3713 1973 3727 1987
rect 3753 2033 3767 2047
rect 3753 1973 3767 1987
rect 3733 1953 3747 1967
rect 3833 1953 3847 1967
rect 3813 1893 3827 1907
rect 3793 1853 3807 1867
rect 3773 1813 3787 1827
rect 3553 1653 3567 1667
rect 3593 1653 3607 1667
rect 3473 1633 3487 1647
rect 3533 1613 3547 1627
rect 3433 1593 3447 1607
rect 3413 1573 3427 1587
rect 3513 1573 3527 1587
rect 3393 1513 3407 1527
rect 3353 1493 3367 1507
rect 3313 1453 3327 1467
rect 3253 1413 3267 1427
rect 3273 1413 3287 1427
rect 3253 1393 3267 1407
rect 3233 1353 3247 1367
rect 3213 1333 3227 1347
rect 3193 1213 3207 1227
rect 3133 1173 3147 1187
rect 3133 1153 3147 1167
rect 3233 1273 3247 1287
rect 3113 1073 3127 1087
rect 2993 993 3007 1007
rect 3073 993 3087 1007
rect 2913 833 2927 847
rect 2933 833 2947 847
rect 2973 833 2987 847
rect 2953 813 2967 827
rect 2813 773 2827 787
rect 2813 693 2827 707
rect 2833 673 2847 687
rect 2813 613 2827 627
rect 3093 953 3107 967
rect 3213 1153 3227 1167
rect 3333 1293 3347 1307
rect 3313 1213 3327 1227
rect 3273 1193 3287 1207
rect 3253 1173 3267 1187
rect 3233 1133 3247 1147
rect 3573 1553 3587 1567
rect 3453 1473 3467 1487
rect 3473 1453 3487 1467
rect 3373 1413 3387 1427
rect 3393 1413 3407 1427
rect 3393 1333 3407 1347
rect 3393 1293 3407 1307
rect 3373 1253 3387 1267
rect 3353 1133 3367 1147
rect 3453 1333 3467 1347
rect 3393 1193 3407 1207
rect 3493 1433 3507 1447
rect 3693 1753 3707 1767
rect 3813 1813 3827 1827
rect 4013 2473 4027 2487
rect 3973 2433 3987 2447
rect 4013 2373 4027 2387
rect 3993 2253 4007 2267
rect 3953 2233 3967 2247
rect 3973 2233 3987 2247
rect 3973 2193 3987 2207
rect 4133 2573 4147 2587
rect 4093 2513 4107 2527
rect 4053 2453 4067 2467
rect 4073 2453 4087 2467
rect 4073 2413 4087 2427
rect 4053 2393 4067 2407
rect 4033 2293 4047 2307
rect 4033 2273 4047 2287
rect 4013 2213 4027 2227
rect 4033 2193 4047 2207
rect 4053 2193 4067 2207
rect 3993 2173 4007 2187
rect 4013 2173 4027 2187
rect 3933 2093 3947 2107
rect 3953 2093 3967 2107
rect 4033 2153 4047 2167
rect 4013 2113 4027 2127
rect 4013 2093 4027 2107
rect 4033 2093 4047 2107
rect 3913 2053 3927 2067
rect 3933 2053 3947 2067
rect 4113 2493 4127 2507
rect 4133 2433 4147 2447
rect 4113 2293 4127 2307
rect 4113 2253 4127 2267
rect 4153 2413 4167 2427
rect 4193 2633 4207 2647
rect 4233 2613 4247 2627
rect 4193 2593 4207 2607
rect 4213 2593 4227 2607
rect 4193 2573 4207 2587
rect 4273 2673 4287 2687
rect 4293 2593 4307 2607
rect 4253 2573 4267 2587
rect 4273 2553 4287 2567
rect 4293 2533 4307 2547
rect 4233 2493 4247 2507
rect 4213 2453 4227 2467
rect 4253 2473 4267 2487
rect 4253 2453 4267 2467
rect 4173 2373 4187 2387
rect 4193 2353 4207 2367
rect 4093 2213 4107 2227
rect 4073 2153 4087 2167
rect 4093 2073 4107 2087
rect 4013 2053 4027 2067
rect 3893 2033 3907 2047
rect 3893 1993 3907 2007
rect 3953 2033 3967 2047
rect 3993 2033 4007 2047
rect 4053 2033 4067 2047
rect 3933 1973 3947 1987
rect 3913 1953 3927 1967
rect 4093 2013 4107 2027
rect 4173 2233 4187 2247
rect 4133 2213 4147 2227
rect 4233 2373 4247 2387
rect 4233 2293 4247 2307
rect 4293 2413 4307 2427
rect 4273 2293 4287 2307
rect 4333 2713 4347 2727
rect 4393 2733 4407 2747
rect 4373 2713 4387 2727
rect 4433 2713 4447 2727
rect 4393 2693 4407 2707
rect 4433 2693 4447 2707
rect 4713 3233 4727 3247
rect 4693 3213 4707 3227
rect 4713 3193 4727 3207
rect 4673 3073 4687 3087
rect 4673 3053 4687 3067
rect 4653 3013 4667 3027
rect 4893 3353 4907 3367
rect 4813 3273 4827 3287
rect 4793 3233 4807 3247
rect 4853 3233 4867 3247
rect 4913 3213 4927 3227
rect 4853 3193 4867 3207
rect 4913 3193 4927 3207
rect 4753 3133 4767 3147
rect 4733 3073 4747 3087
rect 4713 3053 4727 3067
rect 4633 2993 4647 3007
rect 4653 2993 4667 3007
rect 4693 2993 4707 3007
rect 4713 2993 4727 3007
rect 4593 2873 4607 2887
rect 4553 2833 4567 2847
rect 4513 2813 4527 2827
rect 4513 2773 4527 2787
rect 4573 2773 4587 2787
rect 4353 2653 4367 2667
rect 4353 2633 4367 2647
rect 4313 2373 4327 2387
rect 4373 2613 4387 2627
rect 4413 2653 4427 2667
rect 4413 2593 4427 2607
rect 4413 2513 4427 2527
rect 4393 2473 4407 2487
rect 4493 2693 4507 2707
rect 4533 2693 4547 2707
rect 4513 2673 4527 2687
rect 4633 2733 4647 2747
rect 4513 2613 4527 2627
rect 4493 2553 4507 2567
rect 4493 2493 4507 2507
rect 4433 2413 4447 2427
rect 4393 2373 4407 2387
rect 4413 2373 4427 2387
rect 4353 2353 4367 2367
rect 4293 2253 4307 2267
rect 4253 2233 4267 2247
rect 4253 2193 4267 2207
rect 4233 2173 4247 2187
rect 4293 2173 4307 2187
rect 4193 2113 4207 2127
rect 4133 2093 4147 2107
rect 4273 2133 4287 2147
rect 4193 2073 4207 2087
rect 4233 2073 4247 2087
rect 4173 2053 4187 2067
rect 3993 1933 4007 1947
rect 4033 1933 4047 1947
rect 3893 1893 3907 1907
rect 4073 1993 4087 2007
rect 4053 1913 4067 1927
rect 4053 1893 4067 1907
rect 3853 1833 3867 1847
rect 4033 1833 4047 1847
rect 3853 1813 3867 1827
rect 3833 1793 3847 1807
rect 3873 1793 3887 1807
rect 3893 1813 3907 1827
rect 3993 1813 4007 1827
rect 3853 1753 3867 1767
rect 3653 1713 3667 1727
rect 3773 1713 3787 1727
rect 3793 1713 3807 1727
rect 3673 1693 3687 1707
rect 3673 1653 3687 1667
rect 3713 1653 3727 1667
rect 3693 1593 3707 1607
rect 3713 1533 3727 1547
rect 3613 1493 3627 1507
rect 3693 1473 3707 1487
rect 3713 1473 3727 1487
rect 3593 1433 3607 1447
rect 3693 1433 3707 1447
rect 3653 1333 3667 1347
rect 3513 1293 3527 1307
rect 3613 1313 3627 1327
rect 3713 1413 3727 1427
rect 3753 1413 3767 1427
rect 3813 1633 3827 1647
rect 3953 1753 3967 1767
rect 3873 1733 3887 1747
rect 3973 1713 3987 1727
rect 3853 1693 3867 1707
rect 3873 1693 3887 1707
rect 3793 1613 3807 1627
rect 3833 1613 3847 1627
rect 3833 1593 3847 1607
rect 3813 1573 3827 1587
rect 3873 1633 3887 1647
rect 3913 1633 3927 1647
rect 4093 1853 4107 1867
rect 4093 1733 4107 1747
rect 4093 1693 4107 1707
rect 4053 1673 4067 1687
rect 4013 1653 4027 1667
rect 3993 1613 4007 1627
rect 4013 1613 4027 1627
rect 3853 1553 3867 1567
rect 3793 1493 3807 1507
rect 3813 1493 3827 1507
rect 3773 1393 3787 1407
rect 3713 1353 3727 1367
rect 3713 1313 3727 1327
rect 3733 1293 3747 1307
rect 3533 1273 3547 1287
rect 3573 1273 3587 1287
rect 3613 1273 3627 1287
rect 3573 1233 3587 1247
rect 3493 1213 3507 1227
rect 3513 1213 3527 1227
rect 3473 1173 3487 1187
rect 3193 1093 3207 1107
rect 3173 1073 3187 1087
rect 3233 1093 3247 1107
rect 3273 1093 3287 1107
rect 3253 1073 3267 1087
rect 3133 953 3147 967
rect 3113 913 3127 927
rect 3093 873 3107 887
rect 3213 993 3227 1007
rect 3173 953 3187 967
rect 3193 953 3207 967
rect 3033 833 3047 847
rect 2993 793 3007 807
rect 2973 773 2987 787
rect 2913 713 2927 727
rect 2933 693 2947 707
rect 3053 713 3067 727
rect 3053 693 3067 707
rect 2873 653 2887 667
rect 2933 653 2947 667
rect 2953 653 2967 667
rect 3013 653 3027 667
rect 2893 613 2907 627
rect 3153 833 3167 847
rect 3173 793 3187 807
rect 3153 753 3167 767
rect 3113 693 3127 707
rect 3093 673 3107 687
rect 3093 653 3107 667
rect 2933 613 2947 627
rect 2853 593 2867 607
rect 3013 593 3027 607
rect 3413 1093 3427 1107
rect 3433 1113 3447 1127
rect 3493 1113 3507 1127
rect 3293 1073 3307 1087
rect 3313 1073 3327 1087
rect 3333 1073 3347 1087
rect 3373 1053 3387 1067
rect 3313 1033 3327 1047
rect 3273 1013 3287 1027
rect 3313 953 3327 967
rect 3253 833 3267 847
rect 3233 773 3247 787
rect 3173 693 3187 707
rect 3153 633 3167 647
rect 3233 733 3247 747
rect 3193 653 3207 667
rect 2973 533 2987 547
rect 2753 373 2767 387
rect 2733 333 2747 347
rect 2793 373 2807 387
rect 2813 373 2827 387
rect 2933 373 2947 387
rect 2773 333 2787 347
rect 2593 253 2607 267
rect 2593 213 2607 227
rect 2573 193 2587 207
rect 2653 193 2667 207
rect 2553 153 2567 167
rect 2533 133 2547 147
rect 2573 133 2587 147
rect 2613 153 2627 167
rect 2633 133 2647 147
rect 2613 113 2627 127
rect 2413 93 2427 107
rect 2433 93 2447 107
rect 2733 113 2747 127
rect 2793 253 2807 267
rect 2853 313 2867 327
rect 2873 313 2887 327
rect 2933 313 2947 327
rect 3013 553 3027 567
rect 3053 533 3067 547
rect 3033 473 3047 487
rect 2993 373 3007 387
rect 2853 273 2867 287
rect 3013 253 3027 267
rect 2833 233 2847 247
rect 2793 173 2807 187
rect 2893 193 2907 207
rect 2993 193 3007 207
rect 3093 413 3107 427
rect 3053 293 3067 307
rect 3073 273 3087 287
rect 3053 173 3067 187
rect 2953 153 2967 167
rect 2893 113 2907 127
rect 3173 553 3187 567
rect 3253 493 3267 507
rect 3493 1033 3507 1047
rect 3433 1013 3447 1027
rect 3453 1013 3467 1027
rect 3393 953 3407 967
rect 3373 933 3387 947
rect 3393 933 3407 947
rect 3453 913 3467 927
rect 3473 913 3487 927
rect 3333 833 3347 847
rect 3373 813 3387 827
rect 3533 1153 3547 1167
rect 3553 1113 3567 1127
rect 3553 1073 3567 1087
rect 3593 1153 3607 1167
rect 3593 1133 3607 1147
rect 3693 1273 3707 1287
rect 3733 1253 3747 1267
rect 3713 1213 3727 1227
rect 3693 1193 3707 1207
rect 3633 1113 3647 1127
rect 3673 1153 3687 1167
rect 3693 1153 3707 1167
rect 3693 1113 3707 1127
rect 3673 1093 3687 1107
rect 3613 1013 3627 1027
rect 3633 1013 3647 1027
rect 3573 973 3587 987
rect 3553 953 3567 967
rect 3613 913 3627 927
rect 3513 873 3527 887
rect 3533 873 3547 887
rect 3573 873 3587 887
rect 3333 713 3347 727
rect 3353 713 3367 727
rect 3293 693 3307 707
rect 3393 673 3407 687
rect 3333 653 3347 667
rect 3353 653 3367 667
rect 3313 613 3327 627
rect 3553 833 3567 847
rect 3493 773 3507 787
rect 3453 713 3467 727
rect 3413 653 3427 667
rect 3593 813 3607 827
rect 3553 773 3567 787
rect 3533 753 3547 767
rect 3373 613 3387 627
rect 3433 633 3447 647
rect 3493 633 3507 647
rect 3413 613 3427 627
rect 3333 593 3347 607
rect 3393 573 3407 587
rect 3413 473 3427 487
rect 3393 453 3407 467
rect 3193 353 3207 367
rect 3093 233 3107 247
rect 3233 233 3247 247
rect 3113 193 3127 207
rect 3153 193 3167 207
rect 3313 393 3327 407
rect 3273 353 3287 367
rect 3453 593 3467 607
rect 3473 613 3487 627
rect 3593 633 3607 647
rect 3493 593 3507 607
rect 3473 493 3487 507
rect 3433 453 3447 467
rect 3853 1433 3867 1447
rect 4013 1513 4027 1527
rect 3953 1433 3967 1447
rect 3953 1373 3967 1387
rect 3973 1373 3987 1387
rect 3873 1333 3887 1347
rect 3793 1253 3807 1267
rect 3753 1213 3767 1227
rect 3773 1153 3787 1167
rect 3833 1253 3847 1267
rect 3713 993 3727 1007
rect 3653 933 3667 947
rect 3693 913 3707 927
rect 3733 833 3747 847
rect 3653 793 3667 807
rect 3713 793 3727 807
rect 3673 753 3687 767
rect 3813 1153 3827 1167
rect 3813 1113 3827 1127
rect 3773 1053 3787 1067
rect 3793 953 3807 967
rect 3773 853 3787 867
rect 3913 1333 3927 1347
rect 3853 1173 3867 1187
rect 3873 1153 3887 1167
rect 3893 1153 3907 1167
rect 3873 1113 3887 1127
rect 3953 1273 3967 1287
rect 3933 1173 3947 1187
rect 3913 1133 3927 1147
rect 3933 1113 3947 1127
rect 3953 1113 3967 1127
rect 3893 1033 3907 1047
rect 3953 1033 3967 1047
rect 3913 1013 3927 1027
rect 3853 953 3867 967
rect 3913 933 3927 947
rect 3833 853 3847 867
rect 3873 873 3887 887
rect 3953 913 3967 927
rect 3913 813 3927 827
rect 3873 773 3887 787
rect 3773 753 3787 767
rect 3793 753 3807 767
rect 3813 753 3827 767
rect 3753 733 3767 747
rect 3713 653 3727 667
rect 3633 633 3647 647
rect 3653 613 3667 627
rect 3713 633 3727 647
rect 3733 613 3747 627
rect 3773 613 3787 627
rect 3613 533 3627 547
rect 3633 513 3647 527
rect 3573 493 3587 507
rect 3573 413 3587 427
rect 3553 393 3567 407
rect 3633 393 3647 407
rect 3513 373 3527 387
rect 3533 373 3547 387
rect 3753 593 3767 607
rect 3853 713 3867 727
rect 3993 1293 4007 1307
rect 4113 1633 4127 1647
rect 4173 2013 4187 2027
rect 4153 1993 4167 2007
rect 4173 1973 4187 1987
rect 4153 1933 4167 1947
rect 4173 1933 4187 1947
rect 4213 1913 4227 1927
rect 4173 1893 4187 1907
rect 4273 2033 4287 2047
rect 4293 1973 4307 1987
rect 4253 1953 4267 1967
rect 4233 1893 4247 1907
rect 4213 1873 4227 1887
rect 4233 1873 4247 1887
rect 4293 1813 4307 1827
rect 4333 2253 4347 2267
rect 4373 2253 4387 2267
rect 4333 2233 4347 2247
rect 4553 2613 4567 2627
rect 4553 2593 4567 2607
rect 4733 2973 4747 2987
rect 4793 3093 4807 3107
rect 4853 3093 4867 3107
rect 4853 3053 4867 3067
rect 4913 3053 4927 3067
rect 4813 3033 4827 3047
rect 4833 3013 4847 3027
rect 4893 3033 4907 3047
rect 4773 2993 4787 3007
rect 4793 2993 4807 3007
rect 4813 2973 4827 2987
rect 4713 2873 4727 2887
rect 4773 2873 4787 2887
rect 4693 2853 4707 2867
rect 4833 2933 4847 2947
rect 4973 3413 4987 3427
rect 4953 3253 4967 3267
rect 5053 3573 5067 3587
rect 5013 3533 5027 3547
rect 5333 3733 5347 3747
rect 5373 3733 5387 3747
rect 5273 3713 5287 3727
rect 5353 3713 5367 3727
rect 5213 3673 5227 3687
rect 5293 3673 5307 3687
rect 5353 3653 5367 3667
rect 5313 3573 5327 3587
rect 5073 3493 5087 3507
rect 5133 3493 5147 3507
rect 4993 3273 5007 3287
rect 4993 3253 5007 3267
rect 4973 3233 4987 3247
rect 5233 3553 5247 3567
rect 5273 3533 5287 3547
rect 5273 3453 5287 3467
rect 5213 3273 5227 3287
rect 5173 3253 5187 3267
rect 5153 3213 5167 3227
rect 5053 3153 5067 3167
rect 5033 3133 5047 3147
rect 5153 3133 5167 3147
rect 4973 3093 4987 3107
rect 4993 3093 5007 3107
rect 4973 3053 4987 3067
rect 5013 3053 5027 3067
rect 5113 3093 5127 3107
rect 4953 3013 4967 3027
rect 4973 3013 4987 3027
rect 4953 2993 4967 3007
rect 4913 2913 4927 2927
rect 4933 2913 4947 2927
rect 4893 2893 4907 2907
rect 4973 2953 4987 2967
rect 4993 2913 5007 2927
rect 4833 2813 4847 2827
rect 4813 2773 4827 2787
rect 4873 2733 4887 2747
rect 4673 2713 4687 2727
rect 4733 2713 4747 2727
rect 4813 2713 4827 2727
rect 4813 2693 4827 2707
rect 4833 2693 4847 2707
rect 4733 2633 4747 2647
rect 4793 2633 4807 2647
rect 4753 2613 4767 2627
rect 4733 2593 4747 2607
rect 4673 2573 4687 2587
rect 4613 2553 4627 2567
rect 4573 2533 4587 2547
rect 4633 2533 4647 2547
rect 4553 2513 4567 2527
rect 4553 2493 4567 2507
rect 4533 2353 4547 2367
rect 4513 2333 4527 2347
rect 4493 2273 4507 2287
rect 4673 2493 4687 2507
rect 4573 2413 4587 2427
rect 4673 2393 4687 2407
rect 4593 2353 4607 2367
rect 4533 2253 4547 2267
rect 4493 2233 4507 2247
rect 4373 2213 4387 2227
rect 4393 2213 4407 2227
rect 4453 2153 4467 2167
rect 4373 2133 4387 2147
rect 4453 2133 4467 2147
rect 4333 2093 4347 2107
rect 4333 2073 4347 2087
rect 4373 2073 4387 2087
rect 4553 2193 4567 2207
rect 4533 2153 4547 2167
rect 4533 2113 4547 2127
rect 4433 2093 4447 2107
rect 4413 2073 4427 2087
rect 4653 2273 4667 2287
rect 4593 2233 4607 2247
rect 4593 2193 4607 2207
rect 4573 2133 4587 2147
rect 4773 2513 4787 2527
rect 4813 2473 4827 2487
rect 4753 2373 4767 2387
rect 4713 2333 4727 2347
rect 4733 2333 4747 2347
rect 4773 2353 4787 2367
rect 4753 2253 4767 2267
rect 4713 2213 4727 2227
rect 4633 2133 4647 2147
rect 4673 2133 4687 2147
rect 4813 2253 4827 2267
rect 4773 2193 4787 2207
rect 4813 2193 4827 2207
rect 4753 2173 4767 2187
rect 4713 2113 4727 2127
rect 4613 2093 4627 2107
rect 4653 2093 4667 2107
rect 4453 2053 4467 2067
rect 4433 2013 4447 2027
rect 4433 1993 4447 2007
rect 4433 1953 4447 1967
rect 4393 1933 4407 1947
rect 4333 1913 4347 1927
rect 4353 1853 4367 1867
rect 4333 1833 4347 1847
rect 4173 1793 4187 1807
rect 4313 1793 4327 1807
rect 4273 1773 4287 1787
rect 4293 1773 4307 1787
rect 4153 1753 4167 1767
rect 4173 1733 4187 1747
rect 4193 1693 4207 1707
rect 4153 1673 4167 1687
rect 4173 1673 4187 1687
rect 4253 1713 4267 1727
rect 4253 1693 4267 1707
rect 4053 1473 4067 1487
rect 4093 1473 4107 1487
rect 4013 1233 4027 1247
rect 4073 1393 4087 1407
rect 4053 1193 4067 1207
rect 4053 1153 4067 1167
rect 4233 1593 4247 1607
rect 4253 1573 4267 1587
rect 4193 1493 4207 1507
rect 4173 1433 4187 1447
rect 4253 1433 4267 1447
rect 4293 1733 4307 1747
rect 4293 1633 4307 1647
rect 4673 2073 4687 2087
rect 4653 2053 4667 2067
rect 4693 2053 4707 2067
rect 4533 2033 4547 2047
rect 4573 2033 4587 2047
rect 4613 2033 4627 2047
rect 4473 1933 4487 1947
rect 4473 1833 4487 1847
rect 4353 1753 4367 1767
rect 4433 1773 4447 1787
rect 4473 1773 4487 1787
rect 4453 1753 4467 1767
rect 4393 1733 4407 1747
rect 4373 1713 4387 1727
rect 4453 1693 4467 1707
rect 4393 1653 4407 1667
rect 4353 1613 4367 1627
rect 4333 1553 4347 1567
rect 4373 1533 4387 1547
rect 4313 1513 4327 1527
rect 4413 1633 4427 1647
rect 4333 1473 4347 1487
rect 4393 1473 4407 1487
rect 4413 1473 4427 1487
rect 4153 1373 4167 1387
rect 4093 1293 4107 1307
rect 4093 1173 4107 1187
rect 4153 1213 4167 1227
rect 4153 1173 4167 1187
rect 4233 1413 4247 1427
rect 4233 1333 4247 1347
rect 4193 1273 4207 1287
rect 4233 1213 4247 1227
rect 4153 1153 4167 1167
rect 4173 1153 4187 1167
rect 3993 1133 4007 1147
rect 4033 1133 4047 1147
rect 4073 1133 4087 1147
rect 4113 1133 4127 1147
rect 4193 1133 4207 1147
rect 3973 893 3987 907
rect 4053 1113 4067 1127
rect 4073 1093 4087 1107
rect 4113 1093 4127 1107
rect 4153 1113 4167 1127
rect 4173 1093 4187 1107
rect 4233 1113 4247 1127
rect 4113 1033 4127 1047
rect 4033 1013 4047 1027
rect 4033 993 4047 1007
rect 3953 773 3967 787
rect 4013 853 4027 867
rect 4013 813 4027 827
rect 4053 953 4067 967
rect 4173 953 4187 967
rect 4133 913 4147 927
rect 4213 913 4227 927
rect 4313 1353 4327 1367
rect 4293 1253 4307 1267
rect 4533 1933 4547 1947
rect 4633 1933 4647 1947
rect 4573 1833 4587 1847
rect 4513 1773 4527 1787
rect 4693 1933 4707 1947
rect 4853 2673 4867 2687
rect 4933 2813 4947 2827
rect 4913 2793 4927 2807
rect 4933 2773 4947 2787
rect 4973 2733 4987 2747
rect 4913 2713 4927 2727
rect 4953 2713 4967 2727
rect 4913 2693 4927 2707
rect 4893 2673 4907 2687
rect 4973 2673 4987 2687
rect 4913 2653 4927 2667
rect 4873 2633 4887 2647
rect 4853 2513 4867 2527
rect 4893 2593 4907 2607
rect 4893 2353 4907 2367
rect 4873 2273 4887 2287
rect 4933 2553 4947 2567
rect 4953 2553 4967 2567
rect 4953 2433 4967 2447
rect 4973 2433 4987 2447
rect 5033 2993 5047 3007
rect 5013 2833 5027 2847
rect 5053 2893 5067 2907
rect 5093 2853 5107 2867
rect 5033 2773 5047 2787
rect 5053 2773 5067 2787
rect 5113 2773 5127 2787
rect 5213 3173 5227 3187
rect 5253 3233 5267 3247
rect 5193 3053 5207 3067
rect 5473 3713 5487 3727
rect 5433 3493 5447 3507
rect 5373 3413 5387 3427
rect 5293 3353 5307 3367
rect 5273 3213 5287 3227
rect 5153 2993 5167 3007
rect 5313 3313 5327 3327
rect 5553 3873 5567 3887
rect 5693 4113 5707 4127
rect 5693 4093 5707 4107
rect 5633 3953 5647 3967
rect 5633 3913 5647 3927
rect 5673 3993 5687 4007
rect 5673 3953 5687 3967
rect 5613 3853 5627 3867
rect 5513 3753 5527 3767
rect 5593 3753 5607 3767
rect 5513 3713 5527 3727
rect 5533 3693 5547 3707
rect 5513 3533 5527 3547
rect 5573 3493 5587 3507
rect 5553 3473 5567 3487
rect 5533 3353 5547 3367
rect 5473 3293 5487 3307
rect 5493 3293 5507 3307
rect 5413 3253 5427 3267
rect 5473 3253 5487 3267
rect 5493 3253 5507 3267
rect 5353 3233 5367 3247
rect 5393 3233 5407 3247
rect 5333 3193 5347 3207
rect 5373 3193 5387 3207
rect 5293 3153 5307 3167
rect 5333 3153 5347 3167
rect 5373 3153 5387 3167
rect 5373 3113 5387 3127
rect 5313 3093 5327 3107
rect 5273 3033 5287 3047
rect 5253 3013 5267 3027
rect 5153 2973 5167 2987
rect 5173 2973 5187 2987
rect 5153 2813 5167 2827
rect 5233 2913 5247 2927
rect 5213 2833 5227 2847
rect 5273 2993 5287 3007
rect 5233 2793 5247 2807
rect 5253 2793 5267 2807
rect 5233 2773 5247 2787
rect 5013 2733 5027 2747
rect 5033 2753 5047 2767
rect 5053 2733 5067 2747
rect 5093 2733 5107 2747
rect 5133 2753 5147 2767
rect 5153 2753 5167 2767
rect 5033 2713 5047 2727
rect 5073 2713 5087 2727
rect 5173 2713 5187 2727
rect 5033 2653 5047 2667
rect 5053 2613 5067 2627
rect 5033 2573 5047 2587
rect 4933 2333 4947 2347
rect 4993 2373 5007 2387
rect 5033 2433 5047 2447
rect 5033 2413 5047 2427
rect 5013 2293 5027 2307
rect 4873 2193 4887 2207
rect 4873 2133 4887 2147
rect 4833 2113 4847 2127
rect 4733 2053 4747 2067
rect 4793 2073 4807 2087
rect 4753 2033 4767 2047
rect 4753 2013 4767 2027
rect 4713 1873 4727 1887
rect 4693 1853 4707 1867
rect 4653 1833 4667 1847
rect 4613 1793 4627 1807
rect 4673 1773 4687 1787
rect 4513 1753 4527 1767
rect 4533 1753 4547 1767
rect 4533 1733 4547 1747
rect 4493 1693 4507 1707
rect 4473 1653 4487 1667
rect 4513 1653 4527 1667
rect 4513 1613 4527 1627
rect 4593 1753 4607 1767
rect 4573 1713 4587 1727
rect 4553 1653 4567 1667
rect 4713 1833 4727 1847
rect 4833 2073 4847 2087
rect 4973 2213 4987 2227
rect 4973 2173 4987 2187
rect 5013 2213 5027 2227
rect 4993 2153 5007 2167
rect 4893 2093 4907 2107
rect 4953 2093 4967 2107
rect 4853 2053 4867 2067
rect 4893 2073 4907 2087
rect 4973 2073 4987 2087
rect 4813 1993 4827 2007
rect 4893 2033 4907 2047
rect 4873 1933 4887 1947
rect 4853 1893 4867 1907
rect 4873 1893 4887 1907
rect 4873 1853 4887 1867
rect 4813 1833 4827 1847
rect 4713 1793 4727 1807
rect 4733 1793 4747 1807
rect 4753 1793 4767 1807
rect 4693 1733 4707 1747
rect 4733 1733 4747 1747
rect 4593 1673 4607 1687
rect 4633 1673 4647 1687
rect 4593 1653 4607 1667
rect 4713 1653 4727 1667
rect 4533 1593 4547 1607
rect 4473 1533 4487 1547
rect 4493 1533 4507 1547
rect 4713 1613 4727 1627
rect 4653 1593 4667 1607
rect 4693 1573 4707 1587
rect 4553 1493 4567 1507
rect 4453 1413 4467 1427
rect 4493 1413 4507 1427
rect 4453 1353 4467 1367
rect 4333 1333 4347 1347
rect 4413 1333 4427 1347
rect 4433 1333 4447 1347
rect 4353 1313 4367 1327
rect 4333 1293 4347 1307
rect 4393 1293 4407 1307
rect 4413 1313 4427 1327
rect 4513 1313 4527 1327
rect 4333 1273 4347 1287
rect 4353 1273 4367 1287
rect 4293 1213 4307 1227
rect 4313 1213 4327 1227
rect 4273 1133 4287 1147
rect 4293 1133 4307 1147
rect 4433 1273 4447 1287
rect 4433 1253 4447 1267
rect 4353 1133 4367 1147
rect 4393 1133 4407 1147
rect 4533 1293 4547 1307
rect 4513 1273 4527 1287
rect 4493 1233 4507 1247
rect 4513 1233 4527 1247
rect 4473 1213 4487 1227
rect 4533 1133 4547 1147
rect 4393 1113 4407 1127
rect 4373 1093 4387 1107
rect 4453 1093 4467 1107
rect 4493 1093 4507 1107
rect 4313 1033 4327 1047
rect 4353 1033 4367 1047
rect 4333 973 4347 987
rect 4453 1073 4467 1087
rect 4453 973 4467 987
rect 4373 953 4387 967
rect 4413 953 4427 967
rect 4313 913 4327 927
rect 4333 913 4347 927
rect 4253 893 4267 907
rect 4353 893 4367 907
rect 4253 873 4267 887
rect 4093 833 4107 847
rect 4073 813 4087 827
rect 4033 793 4047 807
rect 4053 753 4067 767
rect 4073 753 4087 767
rect 3933 733 3947 747
rect 3993 733 4007 747
rect 3973 713 3987 727
rect 3893 693 3907 707
rect 3913 673 3927 687
rect 3893 653 3907 667
rect 3793 593 3807 607
rect 3873 613 3887 627
rect 3673 553 3687 567
rect 3753 553 3767 567
rect 3833 553 3847 567
rect 3713 513 3727 527
rect 3733 513 3747 527
rect 3713 473 3727 487
rect 3673 393 3687 407
rect 3753 413 3767 427
rect 3733 373 3747 387
rect 3293 253 3307 267
rect 3453 333 3467 347
rect 3493 353 3507 367
rect 3413 313 3427 327
rect 3493 313 3507 327
rect 3533 313 3547 327
rect 3553 313 3567 327
rect 3353 273 3367 287
rect 3393 293 3407 307
rect 3373 253 3387 267
rect 3333 213 3347 227
rect 3133 133 3147 147
rect 2913 93 2927 107
rect 3413 253 3427 267
rect 3413 193 3427 207
rect 3173 93 3187 107
rect 3533 293 3547 307
rect 3533 253 3547 267
rect 3513 233 3527 247
rect 3493 113 3507 127
rect 3653 353 3667 367
rect 3853 453 3867 467
rect 3773 373 3787 387
rect 3793 373 3807 387
rect 3633 333 3647 347
rect 3933 633 3947 647
rect 3933 493 3947 507
rect 3913 393 3927 407
rect 3933 373 3947 387
rect 4013 653 4027 667
rect 4133 813 4147 827
rect 4173 833 4187 847
rect 4253 833 4267 847
rect 4233 813 4247 827
rect 3853 353 3867 367
rect 3873 333 3887 347
rect 3893 333 3907 347
rect 3913 353 3927 367
rect 3953 353 3967 367
rect 3973 353 3987 367
rect 3953 333 3967 347
rect 3733 313 3747 327
rect 3773 313 3787 327
rect 3793 313 3807 327
rect 3593 293 3607 307
rect 3573 213 3587 227
rect 3633 213 3647 227
rect 3613 193 3627 207
rect 3593 173 3607 187
rect 3753 293 3767 307
rect 3653 193 3667 207
rect 3753 173 3767 187
rect 3553 153 3567 167
rect 3593 153 3607 167
rect 3613 153 3627 167
rect 3553 133 3567 147
rect 3613 133 3627 147
rect 3673 153 3687 167
rect 3713 133 3727 147
rect 3733 153 3747 167
rect 3653 113 3667 127
rect 3853 273 3867 287
rect 3893 293 3907 307
rect 4073 513 4087 527
rect 4013 493 4027 507
rect 4173 793 4187 807
rect 4193 793 4207 807
rect 4233 773 4247 787
rect 4193 693 4207 707
rect 4193 593 4207 607
rect 4173 533 4187 547
rect 4153 493 4167 507
rect 4153 473 4167 487
rect 4133 413 4147 427
rect 4033 353 4047 367
rect 4073 313 4087 327
rect 3993 293 4007 307
rect 3953 273 3967 287
rect 3893 253 3907 267
rect 3933 253 3947 267
rect 3793 133 3807 147
rect 3813 113 3827 127
rect 3873 193 3887 207
rect 3933 213 3947 227
rect 3773 73 3787 87
rect 4093 193 4107 207
rect 4093 173 4107 187
rect 4053 133 4067 147
rect 4073 153 4087 167
rect 4193 333 4207 347
rect 4273 813 4287 827
rect 4293 833 4307 847
rect 4333 833 4347 847
rect 4273 793 4287 807
rect 4313 793 4327 807
rect 4333 793 4347 807
rect 4253 693 4267 707
rect 4253 633 4267 647
rect 4233 273 4247 287
rect 4513 1073 4527 1087
rect 4513 993 4527 1007
rect 4513 953 4527 967
rect 4493 933 4507 947
rect 4393 853 4407 867
rect 4393 813 4407 827
rect 4373 733 4387 747
rect 4373 693 4387 707
rect 4333 653 4347 667
rect 4353 653 4367 667
rect 4353 633 4367 647
rect 4293 493 4307 507
rect 4333 453 4347 467
rect 4293 313 4307 327
rect 4273 293 4287 307
rect 4313 253 4327 267
rect 4293 233 4307 247
rect 4173 213 4187 227
rect 4213 213 4227 227
rect 4253 213 4267 227
rect 4173 193 4187 207
rect 4133 153 4147 167
rect 4113 133 4127 147
rect 4153 133 4167 147
rect 4213 153 4227 167
rect 4193 133 4207 147
rect 4013 73 4027 87
rect 4253 133 4267 147
rect 4493 833 4507 847
rect 4473 793 4487 807
rect 4433 753 4447 767
rect 4433 733 4447 747
rect 4453 733 4467 747
rect 4413 713 4427 727
rect 4053 53 4067 67
rect 4333 153 4347 167
rect 4393 393 4407 407
rect 4473 653 4487 667
rect 4453 613 4467 627
rect 4493 613 4507 627
rect 4653 1553 4667 1567
rect 4973 2033 4987 2047
rect 5173 2673 5187 2687
rect 5113 2633 5127 2647
rect 5073 2593 5087 2607
rect 5093 2533 5107 2547
rect 5233 2693 5247 2707
rect 5193 2653 5207 2667
rect 5313 3053 5327 3067
rect 5433 3213 5447 3227
rect 5413 3133 5427 3147
rect 5393 3073 5407 3087
rect 5373 3033 5387 3047
rect 5313 2973 5327 2987
rect 5313 2753 5327 2767
rect 5353 2753 5367 2767
rect 5273 2713 5287 2727
rect 5333 2713 5347 2727
rect 5353 2713 5367 2727
rect 5253 2633 5267 2647
rect 5273 2593 5287 2607
rect 5233 2573 5247 2587
rect 5293 2573 5307 2587
rect 5313 2573 5327 2587
rect 5133 2553 5147 2567
rect 5193 2533 5207 2547
rect 5253 2553 5267 2567
rect 5233 2533 5247 2547
rect 5273 2533 5287 2547
rect 5453 3033 5467 3047
rect 5413 2973 5427 2987
rect 5453 2953 5467 2967
rect 5493 3233 5507 3247
rect 5613 3513 5627 3527
rect 5653 3693 5667 3707
rect 5713 3753 5727 3767
rect 5773 4173 5787 4187
rect 5853 4853 5867 4867
rect 5873 4853 5887 4867
rect 5973 5073 5987 5087
rect 6013 5033 6027 5047
rect 6093 5253 6107 5267
rect 6053 5173 6067 5187
rect 6073 5153 6087 5167
rect 6053 5133 6067 5147
rect 6113 5113 6127 5127
rect 6233 6053 6247 6067
rect 6213 5973 6227 5987
rect 6273 6053 6287 6067
rect 6633 6413 6647 6427
rect 6653 6373 6667 6387
rect 6673 6393 6687 6407
rect 6613 6353 6627 6367
rect 6573 6333 6587 6347
rect 6673 6333 6687 6347
rect 6653 6313 6667 6327
rect 6553 6273 6567 6287
rect 6453 6153 6467 6167
rect 6313 6033 6327 6047
rect 6253 6013 6267 6027
rect 6393 6133 6407 6147
rect 6373 6113 6387 6127
rect 6433 6133 6447 6147
rect 6513 6133 6527 6147
rect 6373 6073 6387 6087
rect 6333 5993 6347 6007
rect 6333 5973 6347 5987
rect 6313 5953 6327 5967
rect 6233 5933 6247 5947
rect 6293 5913 6307 5927
rect 6233 5873 6247 5887
rect 6253 5893 6267 5907
rect 6213 5793 6227 5807
rect 6253 5793 6267 5807
rect 6213 5673 6227 5687
rect 6233 5653 6247 5667
rect 6333 5913 6347 5927
rect 6353 5913 6367 5927
rect 6353 5873 6367 5887
rect 6453 6093 6467 6107
rect 6473 6113 6487 6127
rect 6553 6113 6567 6127
rect 6413 6033 6427 6047
rect 6433 6013 6447 6027
rect 6393 5953 6407 5967
rect 6493 6073 6507 6087
rect 6493 6053 6507 6067
rect 6533 6053 6547 6067
rect 6473 5933 6487 5947
rect 6453 5913 6467 5927
rect 6573 6033 6587 6047
rect 6593 5973 6607 5987
rect 6633 5933 6647 5947
rect 6393 5873 6407 5887
rect 6313 5853 6327 5867
rect 6273 5773 6287 5787
rect 6333 5773 6347 5787
rect 6333 5753 6347 5767
rect 6273 5693 6287 5707
rect 6373 5813 6387 5827
rect 6353 5693 6367 5707
rect 6453 5853 6467 5867
rect 6413 5753 6427 5767
rect 6513 5893 6527 5907
rect 6533 5893 6547 5907
rect 6553 5873 6567 5887
rect 6573 5873 6587 5887
rect 6593 5873 6607 5887
rect 6613 5893 6627 5907
rect 6553 5833 6567 5847
rect 6493 5713 6507 5727
rect 6533 5693 6547 5707
rect 6453 5673 6467 5687
rect 6473 5673 6487 5687
rect 6313 5653 6327 5667
rect 6333 5653 6347 5667
rect 6253 5633 6267 5647
rect 6273 5633 6287 5647
rect 6313 5633 6327 5647
rect 6373 5633 6387 5647
rect 6333 5613 6347 5627
rect 6273 5593 6287 5607
rect 6313 5593 6327 5607
rect 6373 5593 6387 5607
rect 6293 5573 6307 5587
rect 6293 5533 6307 5547
rect 6273 5513 6287 5527
rect 6293 5493 6307 5507
rect 6273 5473 6287 5487
rect 6233 5453 6247 5467
rect 6253 5453 6267 5467
rect 6353 5553 6367 5567
rect 6333 5533 6347 5547
rect 6293 5453 6307 5467
rect 6313 5453 6327 5467
rect 6213 5433 6227 5447
rect 6213 5413 6227 5427
rect 6253 5413 6267 5427
rect 6313 5413 6327 5427
rect 6353 5433 6367 5447
rect 6353 5413 6367 5427
rect 6193 5393 6207 5407
rect 6233 5393 6247 5407
rect 6293 5393 6307 5407
rect 6173 5373 6187 5387
rect 6193 5213 6207 5227
rect 6173 5193 6187 5207
rect 6273 5213 6287 5227
rect 6253 5193 6267 5207
rect 6233 5173 6247 5187
rect 6233 5133 6247 5147
rect 6193 5113 6207 5127
rect 6273 5113 6287 5127
rect 6133 5093 6147 5107
rect 6153 5093 6167 5107
rect 6233 5093 6247 5107
rect 6053 5073 6067 5087
rect 6073 5073 6087 5087
rect 6113 5073 6127 5087
rect 6133 5053 6147 5067
rect 6113 5033 6127 5047
rect 6073 5013 6087 5027
rect 6093 5013 6107 5027
rect 6033 4973 6047 4987
rect 5973 4953 5987 4967
rect 5993 4953 6007 4967
rect 5973 4933 5987 4947
rect 6053 4953 6067 4967
rect 6113 4953 6127 4967
rect 6113 4933 6127 4947
rect 5993 4913 6007 4927
rect 6013 4913 6027 4927
rect 5953 4893 5967 4907
rect 5913 4833 5927 4847
rect 5933 4833 5947 4847
rect 5853 4813 5867 4827
rect 5833 4693 5847 4707
rect 6053 4913 6067 4927
rect 6073 4913 6087 4927
rect 6033 4893 6047 4907
rect 6033 4873 6047 4887
rect 6013 4813 6027 4827
rect 5953 4773 5967 4787
rect 5993 4773 6007 4787
rect 5853 4673 5867 4687
rect 5853 4593 5867 4607
rect 5913 4673 5927 4687
rect 5933 4693 5947 4707
rect 6013 4753 6027 4767
rect 5973 4693 5987 4707
rect 5953 4673 5967 4687
rect 5913 4653 5927 4667
rect 5973 4653 5987 4667
rect 5893 4553 5907 4567
rect 5933 4533 5947 4547
rect 5893 4513 5907 4527
rect 5913 4513 5927 4527
rect 6013 4553 6027 4567
rect 5993 4513 6007 4527
rect 5993 4493 6007 4507
rect 6273 5033 6287 5047
rect 6213 5013 6227 5027
rect 6193 4993 6207 5007
rect 6153 4953 6167 4967
rect 6273 4993 6287 5007
rect 6233 4973 6247 4987
rect 6433 5653 6447 5667
rect 6393 5573 6407 5587
rect 6453 5593 6467 5607
rect 6593 5813 6607 5827
rect 6613 5713 6627 5727
rect 6573 5673 6587 5687
rect 6613 5673 6627 5687
rect 6653 5793 6667 5807
rect 6593 5653 6607 5667
rect 6593 5633 6607 5647
rect 6493 5573 6507 5587
rect 6433 5553 6447 5567
rect 6413 5513 6427 5527
rect 6413 5473 6427 5487
rect 6393 5453 6407 5467
rect 6533 5613 6547 5627
rect 6553 5613 6567 5627
rect 6513 5513 6527 5527
rect 6513 5493 6527 5507
rect 6473 5453 6487 5467
rect 6493 5453 6507 5467
rect 6413 5413 6427 5427
rect 6453 5413 6467 5427
rect 6393 5393 6407 5407
rect 6373 5373 6387 5387
rect 6313 5273 6327 5287
rect 6373 5233 6387 5247
rect 6353 5213 6367 5227
rect 6433 5233 6447 5247
rect 6413 5213 6427 5227
rect 6393 5193 6407 5207
rect 6533 5473 6547 5487
rect 6553 5453 6567 5467
rect 6573 5453 6587 5467
rect 6513 5433 6527 5447
rect 6513 5393 6527 5407
rect 6533 5413 6547 5427
rect 6573 5413 6587 5427
rect 6553 5393 6567 5407
rect 6613 5533 6627 5547
rect 6633 5493 6647 5507
rect 6733 6373 6747 6387
rect 6713 6353 6727 6367
rect 6693 6313 6707 6327
rect 6693 5893 6707 5907
rect 6653 5453 6667 5467
rect 6673 5453 6687 5467
rect 6633 5413 6647 5427
rect 6593 5393 6607 5407
rect 6533 5373 6547 5387
rect 6513 5213 6527 5227
rect 6493 5193 6507 5207
rect 6353 5173 6367 5187
rect 6333 5153 6347 5167
rect 6313 5133 6327 5147
rect 6293 4973 6307 4987
rect 6393 5173 6407 5187
rect 6453 5173 6467 5187
rect 6433 5153 6447 5167
rect 6473 5153 6487 5167
rect 6513 5153 6527 5167
rect 6373 5133 6387 5147
rect 6353 5113 6367 5127
rect 6373 5113 6387 5127
rect 6333 5033 6347 5047
rect 6173 4933 6187 4947
rect 6193 4933 6207 4947
rect 6253 4933 6267 4947
rect 6293 4953 6307 4967
rect 6313 4953 6327 4967
rect 6193 4913 6207 4927
rect 6133 4873 6147 4887
rect 6273 4873 6287 4887
rect 6153 4793 6167 4807
rect 6173 4773 6187 4787
rect 6093 4733 6107 4747
rect 6153 4733 6167 4747
rect 6053 4693 6067 4707
rect 6153 4713 6167 4727
rect 6053 4653 6067 4667
rect 6113 4653 6127 4667
rect 6073 4553 6087 4567
rect 6053 4513 6067 4527
rect 5933 4473 5947 4487
rect 5953 4473 5967 4487
rect 5833 4433 5847 4447
rect 5873 4433 5887 4447
rect 5933 4453 5947 4467
rect 6013 4453 6027 4467
rect 6033 4453 6047 4467
rect 5973 4433 5987 4447
rect 5853 4413 5867 4427
rect 5873 4393 5887 4407
rect 5913 4393 5927 4407
rect 5993 4353 6007 4367
rect 5853 4233 5867 4247
rect 5933 4233 5947 4247
rect 5873 4213 5887 4227
rect 5873 4193 5887 4207
rect 5833 4173 5847 4187
rect 5813 4153 5827 4167
rect 5833 4133 5847 4147
rect 5773 4093 5787 4107
rect 5853 4053 5867 4067
rect 5833 4013 5847 4027
rect 5913 4113 5927 4127
rect 5953 4213 5967 4227
rect 6033 4433 6047 4447
rect 6133 4613 6147 4627
rect 6153 4513 6167 4527
rect 6093 4493 6107 4507
rect 6193 4713 6207 4727
rect 6253 4713 6267 4727
rect 6213 4673 6227 4687
rect 6233 4693 6247 4707
rect 6293 4793 6307 4807
rect 6293 4753 6307 4767
rect 6293 4733 6307 4747
rect 6433 5133 6447 5147
rect 6393 5013 6407 5027
rect 6433 4993 6447 5007
rect 6413 4953 6427 4967
rect 6353 4913 6367 4927
rect 6373 4933 6387 4947
rect 6393 4913 6407 4927
rect 6333 4893 6347 4907
rect 6493 5113 6507 5127
rect 6553 5353 6567 5367
rect 6653 5393 6667 5407
rect 6673 5393 6687 5407
rect 6633 5353 6647 5367
rect 6553 5193 6567 5207
rect 6593 5193 6607 5207
rect 6673 5193 6687 5207
rect 6573 5173 6587 5187
rect 6553 5153 6567 5167
rect 6613 5173 6627 5187
rect 6613 5153 6627 5167
rect 6633 5153 6647 5167
rect 6653 5173 6667 5187
rect 6553 5133 6567 5147
rect 6533 5093 6547 5107
rect 6593 5093 6607 5107
rect 6493 4993 6507 5007
rect 6553 4993 6567 5007
rect 6473 4953 6487 4967
rect 6473 4933 6487 4947
rect 6593 4993 6607 5007
rect 6573 4973 6587 4987
rect 6513 4953 6527 4967
rect 6553 4953 6567 4967
rect 6493 4913 6507 4927
rect 6533 4913 6547 4927
rect 6613 4973 6627 4987
rect 6653 5133 6667 5147
rect 6713 5133 6727 5147
rect 6673 5113 6687 5127
rect 6693 5113 6707 5127
rect 6653 4993 6667 5007
rect 6633 4913 6647 4927
rect 6453 4853 6467 4867
rect 6353 4753 6367 4767
rect 6333 4733 6347 4747
rect 6313 4693 6327 4707
rect 6273 4673 6287 4687
rect 6273 4633 6287 4647
rect 6233 4593 6247 4607
rect 6213 4573 6227 4587
rect 6173 4453 6187 4467
rect 6113 4413 6127 4427
rect 6193 4413 6207 4427
rect 6093 4393 6107 4407
rect 6073 4373 6087 4387
rect 6273 4573 6287 4587
rect 6353 4713 6367 4727
rect 6413 4713 6427 4727
rect 6433 4713 6447 4727
rect 6373 4693 6387 4707
rect 6333 4593 6347 4607
rect 6393 4653 6407 4667
rect 6433 4653 6447 4667
rect 6373 4613 6387 4627
rect 6373 4593 6387 4607
rect 6353 4573 6367 4587
rect 6253 4533 6267 4547
rect 6313 4533 6327 4547
rect 6253 4493 6267 4507
rect 6353 4513 6367 4527
rect 6373 4513 6387 4527
rect 6333 4493 6347 4507
rect 6273 4473 6287 4487
rect 6353 4473 6367 4487
rect 6233 4413 6247 4427
rect 6313 4433 6327 4447
rect 6433 4633 6447 4647
rect 6473 4793 6487 4807
rect 6493 4773 6507 4787
rect 6513 4733 6527 4747
rect 6473 4693 6487 4707
rect 6493 4693 6507 4707
rect 6633 4833 6647 4847
rect 6553 4733 6567 4747
rect 6613 4733 6627 4747
rect 6653 4713 6667 4727
rect 6673 4713 6687 4727
rect 6573 4693 6587 4707
rect 6553 4653 6567 4667
rect 6453 4613 6467 4627
rect 6513 4633 6527 4647
rect 6473 4593 6487 4607
rect 6473 4553 6487 4567
rect 6453 4513 6467 4527
rect 6493 4513 6507 4527
rect 6393 4473 6407 4487
rect 6553 4553 6567 4567
rect 6573 4513 6587 4527
rect 6533 4473 6547 4487
rect 6393 4433 6407 4447
rect 6433 4453 6447 4467
rect 6453 4453 6467 4467
rect 6453 4433 6467 4447
rect 6513 4453 6527 4467
rect 6553 4453 6567 4467
rect 6613 4613 6627 4627
rect 6613 4533 6627 4547
rect 6633 4493 6647 4507
rect 6613 4473 6627 4487
rect 6593 4453 6607 4467
rect 6653 4453 6667 4467
rect 6513 4433 6527 4447
rect 6293 4413 6307 4427
rect 6233 4373 6247 4387
rect 6273 4373 6287 4387
rect 6213 4353 6227 4367
rect 6053 4333 6067 4347
rect 6013 4313 6027 4327
rect 6093 4313 6107 4327
rect 6033 4213 6047 4227
rect 5973 4173 5987 4187
rect 5993 4193 6007 4207
rect 6013 4173 6027 4187
rect 6073 4193 6087 4207
rect 6073 4173 6087 4187
rect 6013 4153 6027 4167
rect 5893 4093 5907 4107
rect 5813 3993 5827 4007
rect 5773 3933 5787 3947
rect 5833 3953 5847 3967
rect 5853 3953 5867 3967
rect 6053 4093 6067 4107
rect 6013 3993 6027 4007
rect 6033 3993 6047 4007
rect 5893 3953 5907 3967
rect 5933 3953 5947 3967
rect 5973 3953 5987 3967
rect 5873 3933 5887 3947
rect 5793 3873 5807 3887
rect 5853 3873 5867 3887
rect 5813 3733 5827 3747
rect 5773 3713 5787 3727
rect 5793 3713 5807 3727
rect 5833 3673 5847 3687
rect 5793 3613 5807 3627
rect 5913 3713 5927 3727
rect 5933 3733 5947 3747
rect 5913 3693 5927 3707
rect 5793 3573 5807 3587
rect 5873 3573 5887 3587
rect 5693 3553 5707 3567
rect 5753 3553 5767 3567
rect 5653 3533 5667 3547
rect 5733 3533 5747 3547
rect 5753 3533 5767 3547
rect 5653 3513 5667 3527
rect 5713 3513 5727 3527
rect 5713 3493 5727 3507
rect 5673 3473 5687 3487
rect 5633 3453 5647 3467
rect 5633 3413 5647 3427
rect 5613 3333 5627 3347
rect 5553 3153 5567 3167
rect 5553 3133 5567 3147
rect 5513 3113 5527 3127
rect 5533 3053 5547 3067
rect 5573 3053 5587 3067
rect 5693 3373 5707 3387
rect 5693 3333 5707 3347
rect 5673 3313 5687 3327
rect 5673 3293 5687 3307
rect 5653 3053 5667 3067
rect 5473 2933 5487 2947
rect 5533 3013 5547 3027
rect 5633 3033 5647 3047
rect 5513 2973 5527 2987
rect 5493 2913 5507 2927
rect 5453 2813 5467 2827
rect 5513 2833 5527 2847
rect 5493 2793 5507 2807
rect 5393 2773 5407 2787
rect 5433 2773 5447 2787
rect 5373 2673 5387 2687
rect 5473 2753 5487 2767
rect 5493 2733 5507 2747
rect 5473 2713 5487 2727
rect 5433 2693 5447 2707
rect 5433 2673 5447 2687
rect 5473 2673 5487 2687
rect 5393 2653 5407 2667
rect 5413 2633 5427 2647
rect 5373 2593 5387 2607
rect 5353 2573 5367 2587
rect 5333 2533 5347 2547
rect 5373 2533 5387 2547
rect 5153 2493 5167 2507
rect 5193 2493 5207 2507
rect 5293 2453 5307 2467
rect 5193 2433 5207 2447
rect 5113 2353 5127 2367
rect 5153 2353 5167 2367
rect 5153 2313 5167 2327
rect 5173 2313 5187 2327
rect 5073 2253 5087 2267
rect 5053 2213 5067 2227
rect 5093 2213 5107 2227
rect 5053 2193 5067 2207
rect 5153 2193 5167 2207
rect 5133 2153 5147 2167
rect 5093 2133 5107 2147
rect 5113 2133 5127 2147
rect 5053 2113 5067 2127
rect 5133 2093 5147 2107
rect 5033 2073 5047 2087
rect 5053 2073 5067 2087
rect 5093 2073 5107 2087
rect 5113 2073 5127 2087
rect 5253 2353 5267 2367
rect 5273 2313 5287 2327
rect 5313 2353 5327 2367
rect 5293 2293 5307 2307
rect 5213 2253 5227 2267
rect 5273 2213 5287 2227
rect 5173 2133 5187 2147
rect 5193 2133 5207 2147
rect 5213 2133 5227 2147
rect 4933 1993 4947 2007
rect 4953 1993 4967 2007
rect 5013 2013 5027 2027
rect 5033 2013 5047 2027
rect 4973 1933 4987 1947
rect 4933 1913 4947 1927
rect 4973 1873 4987 1887
rect 4873 1773 4887 1787
rect 4853 1753 4867 1767
rect 4913 1753 4927 1767
rect 4893 1713 4907 1727
rect 4873 1673 4887 1687
rect 4893 1673 4907 1687
rect 4813 1653 4827 1667
rect 4853 1653 4867 1667
rect 4753 1633 4767 1647
rect 4813 1573 4827 1587
rect 4833 1593 4847 1607
rect 4653 1513 4667 1527
rect 4593 1493 4607 1507
rect 4633 1493 4647 1507
rect 4593 1413 4607 1427
rect 4733 1533 4747 1547
rect 4613 1353 4627 1367
rect 4633 1353 4647 1367
rect 4713 1353 4727 1367
rect 4573 1333 4587 1347
rect 4573 1313 4587 1327
rect 4613 1313 4627 1327
rect 4593 1293 4607 1307
rect 4713 1333 4727 1347
rect 4793 1553 4807 1567
rect 4793 1533 4807 1547
rect 4773 1393 4787 1407
rect 4733 1293 4747 1307
rect 4633 1253 4647 1267
rect 4613 1193 4627 1207
rect 4653 1193 4667 1207
rect 4573 1153 4587 1167
rect 4573 1113 4587 1127
rect 4573 1073 4587 1087
rect 4553 1053 4567 1067
rect 4533 873 4547 887
rect 4613 1133 4627 1147
rect 4633 1113 4647 1127
rect 4673 1113 4687 1127
rect 4673 1033 4687 1047
rect 4653 1013 4667 1027
rect 4653 933 4667 947
rect 4673 933 4687 947
rect 4613 913 4627 927
rect 4673 893 4687 907
rect 4613 873 4627 887
rect 4653 873 4667 887
rect 4573 853 4587 867
rect 4553 833 4567 847
rect 4593 833 4607 847
rect 4653 833 4667 847
rect 4653 813 4667 827
rect 4533 793 4547 807
rect 4613 793 4627 807
rect 4533 773 4547 787
rect 4653 773 4667 787
rect 4653 753 4667 767
rect 4573 693 4587 707
rect 4613 653 4627 667
rect 4533 633 4547 647
rect 4553 613 4567 627
rect 4593 613 4607 627
rect 4493 553 4507 567
rect 4513 553 4527 567
rect 4493 513 4507 527
rect 4473 473 4487 487
rect 4433 373 4447 387
rect 4513 453 4527 467
rect 4553 453 4567 467
rect 4493 433 4507 447
rect 4513 353 4527 367
rect 4493 333 4507 347
rect 4393 293 4407 307
rect 4413 293 4427 307
rect 4453 193 4467 207
rect 4433 113 4447 127
rect 4373 73 4387 87
rect 4573 333 4587 347
rect 4553 313 4567 327
rect 4533 273 4547 287
rect 4573 293 4587 307
rect 4613 313 4627 327
rect 4713 1273 4727 1287
rect 4753 1273 4767 1287
rect 4773 1273 4787 1287
rect 4813 1433 4827 1447
rect 5153 2073 5167 2087
rect 5133 2053 5147 2067
rect 5193 2073 5207 2087
rect 5113 2033 5127 2047
rect 5093 1993 5107 2007
rect 5033 1913 5047 1927
rect 5073 1913 5087 1927
rect 5013 1813 5027 1827
rect 4973 1793 4987 1807
rect 5053 1773 5067 1787
rect 4993 1753 5007 1767
rect 4973 1733 4987 1747
rect 4913 1633 4927 1647
rect 4893 1593 4907 1607
rect 4953 1593 4967 1607
rect 5013 1653 5027 1667
rect 5013 1593 5027 1607
rect 5013 1573 5027 1587
rect 4913 1553 4927 1567
rect 4993 1553 5007 1567
rect 4853 1373 4867 1387
rect 5053 1633 5067 1647
rect 5053 1593 5067 1607
rect 5013 1533 5027 1547
rect 5013 1493 5027 1507
rect 5053 1473 5067 1487
rect 4933 1413 4947 1427
rect 4953 1393 4967 1407
rect 5113 1833 5127 1847
rect 5153 1973 5167 1987
rect 5253 2113 5267 2127
rect 5213 1953 5227 1967
rect 5253 1993 5267 2007
rect 5233 1833 5247 1847
rect 5133 1813 5147 1827
rect 5153 1813 5167 1827
rect 5193 1793 5207 1807
rect 5233 1773 5247 1787
rect 5093 1753 5107 1767
rect 5113 1753 5127 1767
rect 5173 1753 5187 1767
rect 5193 1753 5207 1767
rect 5093 1733 5107 1747
rect 5113 1733 5127 1747
rect 5093 1653 5107 1667
rect 5093 1593 5107 1607
rect 5193 1713 5207 1727
rect 5173 1673 5187 1687
rect 5133 1593 5147 1607
rect 5153 1593 5167 1607
rect 5113 1573 5127 1587
rect 4953 1373 4967 1387
rect 5073 1373 5087 1387
rect 5233 1753 5247 1767
rect 5213 1673 5227 1687
rect 5293 2193 5307 2207
rect 5373 2433 5387 2447
rect 5393 2393 5407 2407
rect 5373 2313 5387 2327
rect 5333 2173 5347 2187
rect 5353 2173 5367 2187
rect 5313 2153 5327 2167
rect 5333 2133 5347 2147
rect 5373 2133 5387 2147
rect 5293 2093 5307 2107
rect 5473 2653 5487 2667
rect 5533 2793 5547 2807
rect 5593 2993 5607 3007
rect 5593 2933 5607 2947
rect 5633 2933 5647 2947
rect 5573 2793 5587 2807
rect 5553 2773 5567 2787
rect 5553 2713 5567 2727
rect 5573 2673 5587 2687
rect 5513 2633 5527 2647
rect 5573 2613 5587 2627
rect 5573 2593 5587 2607
rect 5553 2573 5567 2587
rect 5493 2553 5507 2567
rect 5533 2533 5547 2547
rect 5493 2513 5507 2527
rect 5433 2353 5447 2367
rect 5413 2333 5427 2347
rect 5433 2333 5447 2347
rect 5413 2293 5427 2307
rect 5453 2293 5467 2307
rect 5413 2253 5427 2267
rect 5433 2273 5447 2287
rect 5433 2213 5447 2227
rect 5413 2193 5427 2207
rect 5473 2193 5487 2207
rect 5513 2273 5527 2287
rect 5533 2213 5547 2227
rect 5433 2173 5447 2187
rect 5513 2153 5527 2167
rect 5433 2113 5447 2127
rect 5633 2753 5647 2767
rect 5593 2513 5607 2527
rect 5693 3253 5707 3267
rect 5853 3553 5867 3567
rect 5893 3553 5907 3567
rect 5833 3493 5847 3507
rect 5773 3473 5787 3487
rect 5753 3433 5767 3447
rect 5733 3253 5747 3267
rect 5893 3533 5907 3547
rect 5873 3493 5887 3507
rect 5893 3493 5907 3507
rect 6033 3853 6047 3867
rect 6173 4233 6187 4247
rect 6133 4213 6147 4227
rect 6093 4113 6107 4127
rect 6073 3833 6087 3847
rect 6073 3773 6087 3787
rect 6153 4173 6167 4187
rect 6253 4313 6267 4327
rect 6193 4213 6207 4227
rect 6173 4133 6187 4147
rect 6213 4133 6227 4147
rect 6173 4113 6187 4127
rect 6153 4013 6167 4027
rect 6173 3993 6187 4007
rect 6213 3993 6227 4007
rect 6133 3893 6147 3907
rect 6153 3893 6167 3907
rect 6113 3773 6127 3787
rect 6093 3753 6107 3767
rect 5933 3673 5947 3687
rect 5953 3673 5967 3687
rect 6013 3713 6027 3727
rect 6093 3713 6107 3727
rect 6013 3653 6027 3667
rect 6053 3673 6067 3687
rect 6073 3673 6087 3687
rect 6033 3633 6047 3647
rect 5973 3553 5987 3567
rect 5933 3533 5947 3547
rect 6053 3533 6067 3547
rect 5953 3493 5967 3507
rect 5973 3513 5987 3527
rect 6013 3513 6027 3527
rect 5853 3373 5867 3387
rect 5873 3333 5887 3347
rect 5833 3293 5847 3307
rect 5833 3273 5847 3287
rect 5753 3233 5767 3247
rect 5773 3233 5787 3247
rect 5733 3113 5747 3127
rect 5813 3213 5827 3227
rect 5833 3233 5847 3247
rect 5833 3173 5847 3187
rect 5793 3153 5807 3167
rect 5773 3133 5787 3147
rect 5753 3053 5767 3067
rect 5913 3153 5927 3167
rect 5973 3473 5987 3487
rect 6033 3473 6047 3487
rect 6033 3413 6047 3427
rect 5973 3353 5987 3367
rect 5993 3353 6007 3367
rect 6013 3353 6027 3367
rect 6073 3353 6087 3367
rect 6053 3273 6067 3287
rect 6093 3273 6107 3287
rect 6033 3213 6047 3227
rect 6093 3233 6107 3247
rect 6493 4413 6507 4427
rect 6313 4393 6327 4407
rect 6313 4333 6327 4347
rect 6413 4333 6427 4347
rect 6573 4413 6587 4427
rect 6553 4373 6567 4387
rect 6513 4313 6527 4327
rect 6453 4293 6467 4307
rect 6433 4273 6447 4287
rect 6433 4253 6447 4267
rect 6293 4213 6307 4227
rect 6333 4213 6347 4227
rect 6373 4213 6387 4227
rect 6273 4173 6287 4187
rect 6293 4173 6307 4187
rect 6393 4193 6407 4207
rect 6493 4273 6507 4287
rect 6433 4193 6447 4207
rect 6473 4193 6487 4207
rect 6333 4153 6347 4167
rect 6353 4153 6367 4167
rect 6273 3993 6287 4007
rect 6253 3773 6267 3787
rect 6413 3953 6427 3967
rect 6553 4233 6567 4247
rect 6513 4213 6527 4227
rect 6673 4253 6687 4267
rect 6693 4233 6707 4247
rect 6593 4213 6607 4227
rect 6513 4173 6527 4187
rect 6553 4193 6567 4207
rect 6573 4193 6587 4207
rect 6593 4193 6607 4207
rect 6613 4193 6627 4207
rect 6653 4173 6667 4187
rect 6573 4153 6587 4167
rect 6613 4153 6627 4167
rect 6633 4153 6647 4167
rect 6533 4073 6547 4087
rect 6653 4133 6667 4147
rect 6573 3913 6587 3927
rect 6453 3793 6467 3807
rect 6493 3793 6507 3807
rect 6413 3773 6427 3787
rect 6273 3733 6287 3747
rect 6293 3733 6307 3747
rect 6313 3733 6327 3747
rect 6373 3753 6387 3767
rect 6153 3713 6167 3727
rect 6173 3693 6187 3707
rect 6193 3713 6207 3727
rect 6213 3713 6227 3727
rect 6233 3713 6247 3727
rect 6133 3633 6147 3647
rect 6273 3713 6287 3727
rect 6193 3673 6207 3687
rect 6213 3673 6227 3687
rect 6233 3673 6247 3687
rect 6173 3653 6187 3667
rect 6153 3613 6167 3627
rect 6213 3633 6227 3647
rect 6233 3633 6247 3647
rect 6193 3533 6207 3547
rect 6253 3593 6267 3607
rect 6253 3533 6267 3547
rect 6253 3433 6267 3447
rect 6133 3413 6147 3427
rect 6233 3373 6247 3387
rect 6193 3353 6207 3367
rect 6133 3293 6147 3307
rect 6153 3293 6167 3307
rect 6213 3313 6227 3327
rect 6113 3213 6127 3227
rect 5953 3133 5967 3147
rect 5993 3133 6007 3147
rect 6133 3193 6147 3207
rect 5933 3113 5947 3127
rect 6073 3113 6087 3127
rect 5853 3093 5867 3107
rect 5873 3093 5887 3107
rect 5853 3053 5867 3067
rect 5973 3053 5987 3067
rect 5933 3033 5947 3047
rect 5913 3013 5927 3027
rect 6133 3173 6147 3187
rect 6153 3133 6167 3147
rect 6253 3293 6267 3307
rect 6253 3273 6267 3287
rect 6233 3253 6247 3267
rect 6253 3253 6267 3267
rect 6313 3693 6327 3707
rect 6353 3693 6367 3707
rect 6353 3653 6367 3667
rect 6433 3693 6447 3707
rect 6413 3633 6427 3647
rect 6693 4033 6707 4047
rect 6493 3773 6507 3787
rect 6653 3773 6667 3787
rect 6333 3593 6347 3607
rect 6453 3593 6467 3607
rect 6293 3433 6307 3447
rect 6293 3413 6307 3427
rect 6293 3273 6307 3287
rect 6233 3213 6247 3227
rect 6273 3233 6287 3247
rect 6273 3193 6287 3207
rect 6253 3153 6267 3167
rect 6293 3153 6307 3167
rect 6193 3093 6207 3107
rect 6213 3093 6227 3107
rect 6173 3073 6187 3087
rect 6113 3053 6127 3067
rect 6173 3053 6187 3067
rect 5993 3013 6007 3027
rect 6033 3033 6047 3047
rect 6113 3013 6127 3027
rect 6153 3013 6167 3027
rect 5793 2993 5807 3007
rect 5693 2933 5707 2947
rect 5713 2933 5727 2947
rect 5713 2873 5727 2887
rect 5713 2773 5727 2787
rect 5653 2693 5667 2707
rect 5673 2693 5687 2707
rect 5653 2673 5667 2687
rect 5773 2733 5787 2747
rect 5853 2973 5867 2987
rect 5913 2953 5927 2967
rect 5853 2813 5867 2827
rect 5813 2793 5827 2807
rect 5813 2753 5827 2767
rect 5833 2713 5847 2727
rect 5873 2793 5887 2807
rect 5793 2673 5807 2687
rect 5853 2673 5867 2687
rect 5973 2853 5987 2867
rect 5933 2833 5947 2847
rect 5953 2833 5967 2847
rect 6233 3073 6247 3087
rect 6253 3073 6267 3087
rect 6213 3053 6227 3067
rect 6273 3013 6287 3027
rect 6173 2993 6187 3007
rect 6213 2993 6227 3007
rect 6053 2833 6067 2847
rect 6013 2793 6027 2807
rect 6153 2813 6167 2827
rect 6093 2793 6107 2807
rect 5993 2753 6007 2767
rect 6013 2733 6027 2747
rect 5953 2713 5967 2727
rect 5973 2713 5987 2727
rect 6013 2713 6027 2727
rect 5893 2693 5907 2707
rect 5913 2693 5927 2707
rect 5873 2653 5887 2667
rect 5753 2633 5767 2647
rect 5813 2633 5827 2647
rect 5833 2633 5847 2647
rect 5773 2613 5787 2627
rect 5733 2573 5747 2587
rect 5813 2573 5827 2587
rect 5653 2533 5667 2547
rect 5673 2533 5687 2547
rect 5713 2533 5727 2547
rect 5773 2553 5787 2567
rect 5613 2373 5627 2387
rect 5633 2373 5647 2387
rect 5613 2293 5627 2307
rect 5833 2513 5847 2527
rect 5833 2473 5847 2487
rect 5773 2453 5787 2467
rect 5733 2433 5747 2447
rect 5673 2413 5687 2427
rect 5653 2333 5667 2347
rect 5593 2253 5607 2267
rect 5653 2253 5667 2267
rect 5573 2233 5587 2247
rect 5653 2233 5667 2247
rect 5393 2093 5407 2107
rect 5713 2393 5727 2407
rect 5873 2433 5887 2447
rect 5793 2413 5807 2427
rect 5773 2353 5787 2367
rect 5833 2373 5847 2387
rect 5813 2353 5827 2367
rect 5733 2313 5747 2327
rect 5833 2313 5847 2327
rect 5753 2273 5767 2287
rect 5793 2273 5807 2287
rect 5853 2293 5867 2307
rect 5833 2273 5847 2287
rect 5713 2253 5727 2267
rect 5733 2253 5747 2267
rect 5673 2193 5687 2207
rect 5653 2113 5667 2127
rect 5773 2233 5787 2247
rect 5873 2273 5887 2287
rect 5873 2233 5887 2247
rect 5753 2213 5767 2227
rect 5853 2213 5867 2227
rect 5973 2633 5987 2647
rect 5913 2613 5927 2627
rect 5953 2613 5967 2627
rect 5993 2613 6007 2627
rect 5973 2573 5987 2587
rect 5993 2573 6007 2587
rect 5913 2553 5927 2567
rect 5993 2553 6007 2567
rect 5913 2493 5927 2507
rect 5953 2493 5967 2507
rect 5933 2473 5947 2487
rect 5933 2313 5947 2327
rect 5913 2293 5927 2307
rect 5913 2273 5927 2287
rect 5933 2273 5947 2287
rect 5913 2233 5927 2247
rect 5933 2233 5947 2247
rect 5893 2213 5907 2227
rect 5873 2193 5887 2207
rect 5913 2193 5927 2207
rect 5753 2173 5767 2187
rect 5853 2173 5867 2187
rect 5793 2133 5807 2147
rect 5553 2093 5567 2107
rect 5593 2093 5607 2107
rect 5353 2053 5367 2067
rect 5393 2073 5407 2087
rect 5453 2053 5467 2067
rect 5493 2073 5507 2087
rect 5393 2013 5407 2027
rect 5273 1973 5287 1987
rect 5333 1933 5347 1947
rect 5293 1813 5307 1827
rect 5273 1793 5287 1807
rect 5313 1793 5327 1807
rect 5353 1773 5367 1787
rect 5253 1733 5267 1747
rect 5353 1693 5367 1707
rect 5253 1673 5267 1687
rect 5313 1673 5327 1687
rect 5253 1633 5267 1647
rect 5233 1613 5247 1627
rect 5213 1593 5227 1607
rect 5253 1593 5267 1607
rect 5253 1513 5267 1527
rect 5233 1493 5247 1507
rect 5253 1493 5267 1507
rect 5153 1453 5167 1467
rect 4993 1353 5007 1367
rect 4813 1333 4827 1347
rect 4793 1233 4807 1247
rect 4813 1233 4827 1247
rect 4773 1213 4787 1227
rect 4753 1173 4767 1187
rect 4913 1333 4927 1347
rect 4893 1233 4907 1247
rect 4833 1213 4847 1227
rect 4793 1173 4807 1187
rect 4833 1153 4847 1167
rect 4773 1133 4787 1147
rect 4873 1133 4887 1147
rect 4753 1093 4767 1107
rect 4753 1033 4767 1047
rect 4793 1113 4807 1127
rect 4853 1093 4867 1107
rect 4793 1073 4807 1087
rect 4813 1073 4827 1087
rect 4733 893 4747 907
rect 4713 853 4727 867
rect 4953 1313 4967 1327
rect 4933 1293 4947 1307
rect 4953 1293 4967 1307
rect 4933 1233 4947 1247
rect 4913 1213 4927 1227
rect 4913 1173 4927 1187
rect 4873 1013 4887 1027
rect 4893 1013 4907 1027
rect 4853 993 4867 1007
rect 4813 933 4827 947
rect 4793 893 4807 907
rect 4753 873 4767 887
rect 4753 833 4767 847
rect 4713 813 4727 827
rect 4773 813 4787 827
rect 4833 833 4847 847
rect 4713 793 4727 807
rect 4733 793 4747 807
rect 4753 793 4767 807
rect 4713 733 4727 747
rect 4713 693 4727 707
rect 4973 1213 4987 1227
rect 4953 1133 4967 1147
rect 5193 1453 5207 1467
rect 5113 1333 5127 1347
rect 5153 1333 5167 1347
rect 5173 1333 5187 1347
rect 5033 1313 5047 1327
rect 5073 1313 5087 1327
rect 5093 1293 5107 1307
rect 5033 1273 5047 1287
rect 5033 1233 5047 1247
rect 4993 1173 5007 1187
rect 5093 1253 5107 1267
rect 5013 1153 5027 1167
rect 5053 1153 5067 1167
rect 4993 1133 5007 1147
rect 4953 1033 4967 1047
rect 4913 993 4927 1007
rect 4873 853 4887 867
rect 4893 833 4907 847
rect 5373 1673 5387 1687
rect 5333 1593 5347 1607
rect 5353 1573 5367 1587
rect 5353 1473 5367 1487
rect 5373 1473 5387 1487
rect 5313 1433 5327 1447
rect 5273 1413 5287 1427
rect 5253 1353 5267 1367
rect 5233 1333 5247 1347
rect 5193 1313 5207 1327
rect 5233 1313 5247 1327
rect 5313 1393 5327 1407
rect 5373 1413 5387 1427
rect 5353 1353 5367 1367
rect 5453 2013 5467 2027
rect 5413 1973 5427 1987
rect 5453 1853 5467 1867
rect 5433 1833 5447 1847
rect 5413 1773 5427 1787
rect 5573 2073 5587 2087
rect 5553 2053 5567 2067
rect 5613 2073 5627 2087
rect 5593 2053 5607 2067
rect 5633 2053 5647 2067
rect 5673 2053 5687 2067
rect 5753 2053 5767 2067
rect 5533 2033 5547 2047
rect 5573 2033 5587 2047
rect 5553 1993 5567 2007
rect 5533 1913 5547 1927
rect 5493 1873 5507 1887
rect 5553 1873 5567 1887
rect 5573 1873 5587 1887
rect 5533 1853 5547 1867
rect 5513 1833 5527 1847
rect 5473 1813 5487 1827
rect 5433 1733 5447 1747
rect 5433 1633 5447 1647
rect 5493 1753 5507 1767
rect 5473 1693 5487 1707
rect 5533 1813 5547 1827
rect 5553 1793 5567 1807
rect 5693 2013 5707 2027
rect 5653 1893 5667 1907
rect 5673 1893 5687 1907
rect 5593 1853 5607 1867
rect 5693 1833 5707 1847
rect 5793 2053 5807 2067
rect 5853 2053 5867 2067
rect 5873 2053 5887 2067
rect 5773 1993 5787 2007
rect 5753 1973 5767 1987
rect 5813 1973 5827 1987
rect 5653 1813 5667 1827
rect 5673 1813 5687 1827
rect 5593 1793 5607 1807
rect 5593 1773 5607 1787
rect 5713 1813 5727 1827
rect 5773 1813 5787 1827
rect 5893 1953 5907 1967
rect 5873 1913 5887 1927
rect 5853 1893 5867 1907
rect 6113 2753 6127 2767
rect 6073 2733 6087 2747
rect 6093 2733 6107 2747
rect 6133 2733 6147 2747
rect 6053 2713 6067 2727
rect 6093 2713 6107 2727
rect 6073 2673 6087 2687
rect 6053 2653 6067 2667
rect 6033 2593 6047 2607
rect 6053 2573 6067 2587
rect 6033 2533 6047 2547
rect 6293 2973 6307 2987
rect 6273 2833 6287 2847
rect 6173 2773 6187 2787
rect 6293 2793 6307 2807
rect 6173 2733 6187 2747
rect 6093 2613 6107 2627
rect 6093 2553 6107 2567
rect 6073 2493 6087 2507
rect 5973 2433 5987 2447
rect 6013 2433 6027 2447
rect 6113 2433 6127 2447
rect 5973 2253 5987 2267
rect 6033 2273 6047 2287
rect 6073 2273 6087 2287
rect 5973 2233 5987 2247
rect 5953 2193 5967 2207
rect 5933 2153 5947 2167
rect 5953 2113 5967 2127
rect 5933 2073 5947 2087
rect 5933 2033 5947 2047
rect 5913 1913 5927 1927
rect 5893 1853 5907 1867
rect 5733 1793 5747 1807
rect 5613 1753 5627 1767
rect 5633 1753 5647 1767
rect 5593 1733 5607 1747
rect 5573 1713 5587 1727
rect 5693 1733 5707 1747
rect 5713 1733 5727 1747
rect 5673 1713 5687 1727
rect 5533 1673 5547 1687
rect 5633 1673 5647 1687
rect 5653 1673 5667 1687
rect 5473 1613 5487 1627
rect 5613 1633 5627 1647
rect 5533 1613 5547 1627
rect 5453 1573 5467 1587
rect 5493 1573 5507 1587
rect 5553 1593 5567 1607
rect 5593 1573 5607 1587
rect 5553 1553 5567 1567
rect 5493 1513 5507 1527
rect 5413 1473 5427 1487
rect 5433 1473 5447 1487
rect 5393 1393 5407 1407
rect 5473 1453 5487 1467
rect 5493 1453 5507 1467
rect 5433 1393 5447 1407
rect 5253 1293 5267 1307
rect 5273 1293 5287 1307
rect 5113 1213 5127 1227
rect 5213 1253 5227 1267
rect 5253 1233 5267 1247
rect 5173 1213 5187 1227
rect 5153 1173 5167 1187
rect 5233 1173 5247 1187
rect 5333 1313 5347 1327
rect 5353 1293 5367 1307
rect 5373 1293 5387 1307
rect 5433 1313 5447 1327
rect 5453 1293 5467 1307
rect 5333 1253 5347 1267
rect 5313 1193 5327 1207
rect 5113 1153 5127 1167
rect 5133 1133 5147 1147
rect 5033 1113 5047 1127
rect 5013 1093 5027 1107
rect 5173 1153 5187 1167
rect 5113 1053 5127 1067
rect 5013 1013 5027 1027
rect 4993 953 5007 967
rect 4993 933 5007 947
rect 4973 813 4987 827
rect 4933 773 4947 787
rect 4853 693 4867 707
rect 4693 653 4707 667
rect 4733 653 4747 667
rect 4753 653 4767 667
rect 4833 653 4847 667
rect 4873 653 4887 667
rect 4913 653 4927 667
rect 4673 633 4687 647
rect 4733 613 4747 627
rect 4793 633 4807 647
rect 4813 613 4827 627
rect 4693 593 4707 607
rect 4753 593 4767 607
rect 4853 593 4867 607
rect 4893 593 4907 607
rect 4953 753 4967 767
rect 4973 653 4987 667
rect 4953 613 4967 627
rect 4973 533 4987 547
rect 4873 513 4887 527
rect 4933 513 4947 527
rect 4753 493 4767 507
rect 4753 373 4767 387
rect 4713 353 4727 367
rect 4773 313 4787 327
rect 4693 273 4707 287
rect 4953 393 4967 407
rect 4973 393 4987 407
rect 4933 333 4947 347
rect 4873 273 4887 287
rect 4973 313 4987 327
rect 4633 253 4647 267
rect 4653 253 4667 267
rect 4833 253 4847 267
rect 4593 213 4607 227
rect 4613 193 4627 207
rect 4613 173 4627 187
rect 4593 153 4607 167
rect 4513 93 4527 107
rect 4573 93 4587 107
rect 4813 233 4827 247
rect 4693 173 4707 187
rect 4653 153 4667 167
rect 4713 133 4727 147
rect 4673 113 4687 127
rect 4773 133 4787 147
rect 5213 973 5227 987
rect 5113 933 5127 947
rect 5173 913 5187 927
rect 5093 893 5107 907
rect 5193 853 5207 867
rect 5113 833 5127 847
rect 5153 813 5167 827
rect 5033 773 5047 787
rect 5093 753 5107 767
rect 5153 733 5167 747
rect 5153 713 5167 727
rect 5013 633 5027 647
rect 5053 633 5067 647
rect 5073 633 5087 647
rect 5013 593 5027 607
rect 4993 293 5007 307
rect 5093 613 5107 627
rect 5113 613 5127 627
rect 5053 593 5067 607
rect 5093 593 5107 607
rect 5133 533 5147 547
rect 5033 513 5047 527
rect 5093 513 5107 527
rect 5053 433 5067 447
rect 5153 453 5167 467
rect 5293 1173 5307 1187
rect 5273 1133 5287 1147
rect 5273 1093 5287 1107
rect 5393 1233 5407 1247
rect 5373 1213 5387 1227
rect 5353 1173 5367 1187
rect 5253 1073 5267 1087
rect 5233 933 5247 947
rect 5253 933 5267 947
rect 5293 1073 5307 1087
rect 5273 833 5287 847
rect 5353 1013 5367 1027
rect 5333 913 5347 927
rect 5313 873 5327 887
rect 5293 813 5307 827
rect 5293 633 5307 647
rect 5453 1253 5467 1267
rect 5533 1513 5547 1527
rect 5553 1493 5567 1507
rect 5493 1413 5507 1427
rect 5513 1413 5527 1427
rect 5493 1353 5507 1367
rect 5513 1333 5527 1347
rect 5613 1513 5627 1527
rect 5593 1453 5607 1467
rect 5573 1373 5587 1387
rect 5653 1653 5667 1667
rect 5693 1673 5707 1687
rect 5653 1613 5667 1627
rect 5673 1613 5687 1627
rect 5673 1593 5687 1607
rect 5893 1793 5907 1807
rect 5753 1673 5767 1687
rect 5853 1733 5867 1747
rect 5833 1693 5847 1707
rect 5813 1653 5827 1667
rect 5793 1633 5807 1647
rect 5953 1853 5967 1867
rect 5933 1773 5947 1787
rect 5893 1693 5907 1707
rect 6033 2233 6047 2247
rect 6013 2213 6027 2227
rect 6053 2213 6067 2227
rect 6013 2093 6027 2107
rect 6013 2053 6027 2067
rect 6053 2073 6067 2087
rect 6093 2253 6107 2267
rect 6093 2233 6107 2247
rect 6153 2633 6167 2647
rect 6253 2713 6267 2727
rect 6293 2693 6307 2707
rect 6193 2633 6207 2647
rect 6213 2553 6227 2567
rect 6193 2533 6207 2547
rect 6153 2333 6167 2347
rect 6153 2253 6167 2267
rect 6173 2273 6187 2287
rect 6093 2153 6107 2167
rect 6093 2073 6107 2087
rect 6093 2013 6107 2027
rect 6293 2433 6307 2447
rect 6293 2353 6307 2367
rect 6373 3353 6387 3367
rect 6333 3313 6347 3327
rect 6333 3273 6347 3287
rect 6373 3253 6387 3267
rect 6373 3213 6387 3227
rect 6393 3213 6407 3227
rect 6413 3233 6427 3247
rect 6473 3233 6487 3247
rect 6433 3213 6447 3227
rect 6353 3193 6367 3207
rect 6453 3193 6467 3207
rect 6353 3173 6367 3187
rect 6373 3173 6387 3187
rect 6433 3153 6447 3167
rect 6353 3053 6367 3067
rect 6333 3033 6347 3047
rect 6353 3013 6367 3027
rect 6373 3033 6387 3047
rect 6393 3013 6407 3027
rect 6413 3033 6427 3047
rect 6333 2993 6347 3007
rect 6373 2933 6387 2947
rect 6333 2813 6347 2827
rect 6393 2793 6407 2807
rect 6353 2713 6367 2727
rect 6333 2613 6347 2627
rect 6373 2613 6387 2627
rect 6413 2573 6427 2587
rect 6453 3133 6467 3147
rect 6513 3753 6527 3767
rect 6553 3713 6567 3727
rect 6633 3733 6647 3747
rect 6573 3693 6587 3707
rect 6533 3613 6547 3627
rect 6633 3633 6647 3647
rect 6573 3593 6587 3607
rect 6593 3593 6607 3607
rect 6533 3453 6547 3467
rect 6513 3253 6527 3267
rect 6553 3273 6567 3287
rect 6513 3213 6527 3227
rect 6553 3233 6567 3247
rect 6553 3213 6567 3227
rect 6553 3173 6567 3187
rect 6593 3393 6607 3407
rect 6613 3273 6627 3287
rect 6593 3253 6607 3267
rect 6633 3253 6647 3267
rect 6573 3153 6587 3167
rect 6553 3133 6567 3147
rect 6493 3113 6507 3127
rect 6533 3113 6547 3127
rect 6493 3093 6507 3107
rect 6473 3073 6487 3087
rect 6493 3053 6507 3067
rect 6453 3013 6467 3027
rect 6493 3013 6507 3027
rect 6513 3013 6527 3027
rect 6453 2693 6467 2707
rect 6513 2713 6527 2727
rect 6513 2693 6527 2707
rect 6493 2653 6507 2667
rect 6413 2553 6427 2567
rect 6433 2533 6447 2547
rect 6413 2453 6427 2467
rect 6393 2393 6407 2407
rect 6333 2353 6347 2367
rect 6393 2353 6407 2367
rect 6313 2313 6327 2327
rect 6373 2333 6387 2347
rect 6373 2293 6387 2307
rect 6433 2413 6447 2427
rect 6433 2393 6447 2407
rect 6473 2533 6487 2547
rect 6613 3193 6627 3207
rect 6593 3053 6607 3067
rect 6633 3153 6647 3167
rect 6633 3073 6647 3087
rect 6573 3013 6587 3027
rect 6573 2993 6587 3007
rect 6633 2973 6647 2987
rect 6553 2733 6567 2747
rect 6573 2733 6587 2747
rect 6573 2713 6587 2727
rect 6533 2573 6547 2587
rect 6533 2533 6547 2547
rect 6493 2513 6507 2527
rect 6693 2653 6707 2667
rect 6693 2613 6707 2627
rect 6573 2553 6587 2567
rect 6593 2533 6607 2547
rect 6653 2553 6667 2567
rect 6573 2513 6587 2527
rect 6453 2333 6467 2347
rect 6473 2333 6487 2347
rect 6473 2313 6487 2327
rect 6413 2293 6427 2307
rect 6453 2293 6467 2307
rect 6233 2273 6247 2287
rect 6313 2273 6327 2287
rect 6353 2273 6367 2287
rect 6153 2213 6167 2227
rect 6193 2213 6207 2227
rect 6113 1993 6127 2007
rect 6073 1933 6087 1947
rect 6053 1893 6067 1907
rect 5973 1833 5987 1847
rect 5973 1793 5987 1807
rect 5973 1773 5987 1787
rect 5953 1753 5967 1767
rect 5893 1653 5907 1667
rect 5913 1653 5927 1667
rect 5833 1613 5847 1627
rect 5713 1593 5727 1607
rect 5733 1573 5747 1587
rect 5693 1513 5707 1527
rect 5633 1493 5647 1507
rect 5633 1473 5647 1487
rect 5613 1333 5627 1347
rect 5513 1293 5527 1307
rect 5553 1313 5567 1327
rect 5573 1313 5587 1327
rect 5513 1273 5527 1287
rect 5553 1273 5567 1287
rect 5473 1213 5487 1227
rect 5413 1193 5427 1207
rect 5413 1173 5427 1187
rect 5473 1173 5487 1187
rect 5453 1153 5467 1167
rect 5433 1133 5447 1147
rect 5413 1073 5427 1087
rect 5373 973 5387 987
rect 5413 893 5427 907
rect 5433 893 5447 907
rect 5353 873 5367 887
rect 5393 853 5407 867
rect 5433 833 5447 847
rect 5353 793 5367 807
rect 5413 793 5427 807
rect 5433 773 5447 787
rect 5413 733 5427 747
rect 5353 673 5367 687
rect 5353 633 5367 647
rect 5333 613 5347 627
rect 5273 533 5287 547
rect 5233 513 5247 527
rect 5253 473 5267 487
rect 5233 453 5247 467
rect 5133 413 5147 427
rect 5193 413 5207 427
rect 5173 393 5187 407
rect 5353 433 5367 447
rect 5333 393 5347 407
rect 5233 373 5247 387
rect 5313 373 5327 387
rect 5673 1433 5687 1447
rect 5653 1353 5667 1367
rect 5693 1413 5707 1427
rect 5793 1553 5807 1567
rect 5733 1453 5747 1467
rect 5773 1453 5787 1467
rect 5753 1413 5767 1427
rect 5733 1393 5747 1407
rect 5713 1373 5727 1387
rect 5713 1353 5727 1367
rect 5653 1253 5667 1267
rect 5553 1213 5567 1227
rect 5633 1213 5647 1227
rect 5533 1113 5547 1127
rect 5633 1113 5647 1127
rect 5493 1073 5507 1087
rect 5553 1073 5567 1087
rect 5473 793 5487 807
rect 5633 1033 5647 1047
rect 5613 893 5627 907
rect 5573 853 5587 867
rect 5513 833 5527 847
rect 5573 833 5587 847
rect 5593 813 5607 827
rect 5493 773 5507 787
rect 5453 753 5467 767
rect 5733 1333 5747 1347
rect 5733 1293 5747 1307
rect 5693 1233 5707 1247
rect 5713 1233 5727 1247
rect 5673 1213 5687 1227
rect 5673 1133 5687 1147
rect 5773 1393 5787 1407
rect 5993 1753 6007 1767
rect 6033 1693 6047 1707
rect 6193 2193 6207 2207
rect 6173 2073 6187 2087
rect 6173 1973 6187 1987
rect 6153 1873 6167 1887
rect 6173 1873 6187 1887
rect 6093 1853 6107 1867
rect 6113 1853 6127 1867
rect 6173 1853 6187 1867
rect 6233 2233 6247 2247
rect 6253 2233 6267 2247
rect 6273 2233 6287 2247
rect 6313 2233 6327 2247
rect 6333 2233 6347 2247
rect 6213 2173 6227 2187
rect 6233 2153 6247 2167
rect 6233 2133 6247 2147
rect 6213 2113 6227 2127
rect 6233 2073 6247 2087
rect 6213 1973 6227 1987
rect 6193 1813 6207 1827
rect 6133 1793 6147 1807
rect 6153 1773 6167 1787
rect 6333 2133 6347 2147
rect 6373 2253 6387 2267
rect 6433 2273 6447 2287
rect 6433 2253 6447 2267
rect 6373 2233 6387 2247
rect 6413 2233 6427 2247
rect 6373 2173 6387 2187
rect 6353 2113 6367 2127
rect 6293 2073 6307 2087
rect 6293 2053 6307 2067
rect 6233 1913 6247 1927
rect 6253 1913 6267 1927
rect 6333 1953 6347 1967
rect 6313 1833 6327 1847
rect 6393 2153 6407 2167
rect 6493 2273 6507 2287
rect 6513 2293 6527 2307
rect 6593 2333 6607 2347
rect 6593 2293 6607 2307
rect 6553 2273 6567 2287
rect 6573 2273 6587 2287
rect 6493 2213 6507 2227
rect 6473 2193 6487 2207
rect 6453 2173 6467 2187
rect 6433 2113 6447 2127
rect 6393 2093 6407 2107
rect 6413 2093 6427 2107
rect 6413 1993 6427 2007
rect 6653 2433 6667 2447
rect 6693 2553 6707 2567
rect 6673 2313 6687 2327
rect 6653 2273 6667 2287
rect 6533 2233 6547 2247
rect 6673 2233 6687 2247
rect 6513 2113 6527 2127
rect 6573 2213 6587 2227
rect 6633 2193 6647 2207
rect 6593 2173 6607 2187
rect 6553 2133 6567 2147
rect 6533 2093 6547 2107
rect 6453 2053 6467 2067
rect 6513 2073 6527 2087
rect 6493 2033 6507 2047
rect 6493 1933 6507 1947
rect 6453 1893 6467 1907
rect 6393 1853 6407 1867
rect 6433 1853 6447 1867
rect 6293 1813 6307 1827
rect 6333 1813 6347 1827
rect 6373 1813 6387 1827
rect 6213 1773 6227 1787
rect 6273 1793 6287 1807
rect 6073 1733 6087 1747
rect 6133 1753 6147 1767
rect 6073 1673 6087 1687
rect 6113 1673 6127 1687
rect 5973 1613 5987 1627
rect 6053 1653 6067 1667
rect 5973 1593 5987 1607
rect 5833 1553 5847 1567
rect 5893 1553 5907 1567
rect 5933 1573 5947 1587
rect 5993 1573 6007 1587
rect 6113 1653 6127 1667
rect 6153 1733 6167 1747
rect 6133 1633 6147 1647
rect 6093 1593 6107 1607
rect 6073 1573 6087 1587
rect 5953 1553 5967 1567
rect 5973 1553 5987 1567
rect 5813 1473 5827 1487
rect 5853 1473 5867 1487
rect 5833 1453 5847 1467
rect 5813 1393 5827 1407
rect 5793 1353 5807 1367
rect 5813 1353 5827 1367
rect 5833 1333 5847 1347
rect 5773 1293 5787 1307
rect 5793 1293 5807 1307
rect 5773 1273 5787 1287
rect 5753 1253 5767 1267
rect 5973 1533 5987 1547
rect 5993 1533 6007 1547
rect 5913 1413 5927 1427
rect 5893 1393 5907 1407
rect 6113 1553 6127 1567
rect 6133 1553 6147 1567
rect 6093 1513 6107 1527
rect 6113 1513 6127 1527
rect 6033 1453 6047 1467
rect 5973 1393 5987 1407
rect 6073 1373 6087 1387
rect 5913 1353 5927 1367
rect 5933 1353 5947 1367
rect 5893 1333 5907 1347
rect 5873 1313 5887 1327
rect 5813 1253 5827 1267
rect 5673 1093 5687 1107
rect 5653 993 5667 1007
rect 5653 933 5667 947
rect 5693 1073 5707 1087
rect 5673 913 5687 927
rect 5733 1053 5747 1067
rect 5793 1233 5807 1247
rect 5873 1293 5887 1307
rect 5953 1313 5967 1327
rect 5973 1313 5987 1327
rect 5933 1293 5947 1307
rect 5893 1273 5907 1287
rect 5873 1253 5887 1267
rect 5853 1233 5867 1247
rect 5913 1233 5927 1247
rect 5833 1173 5847 1187
rect 5813 1153 5827 1167
rect 5773 1133 5787 1147
rect 5893 1153 5907 1167
rect 6073 1313 6087 1327
rect 6013 1253 6027 1267
rect 6053 1253 6067 1267
rect 6033 1233 6047 1247
rect 5993 1213 6007 1227
rect 6033 1193 6047 1207
rect 6013 1153 6027 1167
rect 5773 1093 5787 1107
rect 5813 1093 5827 1107
rect 5853 1113 5867 1127
rect 5873 1093 5887 1107
rect 5933 1113 5947 1127
rect 5833 1073 5847 1087
rect 5853 1073 5867 1087
rect 5873 1073 5887 1087
rect 5953 1093 5967 1107
rect 5933 1073 5947 1087
rect 5753 1033 5767 1047
rect 5813 1033 5827 1047
rect 5853 1033 5867 1047
rect 5833 913 5847 927
rect 5653 893 5667 907
rect 5693 893 5707 907
rect 5713 893 5727 907
rect 5973 1073 5987 1087
rect 5993 1093 6007 1107
rect 6113 1433 6127 1447
rect 6113 1353 6127 1367
rect 6113 1333 6127 1347
rect 6233 1753 6247 1767
rect 6253 1753 6267 1767
rect 6193 1713 6207 1727
rect 6233 1693 6247 1707
rect 6213 1673 6227 1687
rect 6173 1633 6187 1647
rect 6233 1653 6247 1667
rect 6253 1653 6267 1667
rect 6193 1573 6207 1587
rect 6233 1573 6247 1587
rect 6293 1753 6307 1767
rect 6313 1753 6327 1767
rect 6313 1733 6327 1747
rect 6373 1773 6387 1787
rect 6333 1713 6347 1727
rect 6433 1813 6447 1827
rect 6593 2093 6607 2107
rect 6653 2113 6667 2127
rect 6613 2053 6627 2067
rect 6553 2033 6567 2047
rect 6533 1853 6547 1867
rect 6493 1813 6507 1827
rect 6533 1793 6547 1807
rect 6573 1993 6587 2007
rect 6653 1993 6667 2007
rect 6573 1973 6587 1987
rect 6653 1953 6667 1967
rect 6573 1853 6587 1867
rect 6513 1773 6527 1787
rect 6553 1773 6567 1787
rect 6413 1753 6427 1767
rect 6513 1753 6527 1767
rect 6393 1693 6407 1707
rect 6453 1693 6467 1707
rect 6433 1653 6447 1667
rect 6293 1633 6307 1647
rect 6333 1633 6347 1647
rect 6353 1633 6367 1647
rect 6393 1633 6407 1647
rect 6293 1593 6307 1607
rect 6233 1553 6247 1567
rect 6273 1553 6287 1567
rect 6313 1553 6327 1567
rect 6293 1533 6307 1547
rect 6193 1513 6207 1527
rect 6153 1413 6167 1427
rect 6173 1373 6187 1387
rect 6253 1413 6267 1427
rect 6193 1333 6207 1347
rect 6113 1293 6127 1307
rect 6153 1293 6167 1307
rect 6253 1313 6267 1327
rect 6173 1273 6187 1287
rect 6193 1273 6207 1287
rect 6113 1233 6127 1247
rect 6093 1193 6107 1207
rect 6153 1193 6167 1207
rect 6113 1173 6127 1187
rect 6133 1173 6147 1187
rect 6073 1133 6087 1147
rect 6113 1133 6127 1147
rect 6033 1113 6047 1127
rect 6093 1113 6107 1127
rect 5953 1053 5967 1067
rect 6073 1053 6087 1067
rect 5653 873 5667 887
rect 5713 873 5727 887
rect 5873 873 5887 887
rect 5693 853 5707 867
rect 5633 813 5647 827
rect 5633 793 5647 807
rect 5613 773 5627 787
rect 5553 713 5567 727
rect 5613 693 5627 707
rect 5433 573 5447 587
rect 5433 553 5447 567
rect 5453 553 5467 567
rect 5473 533 5487 547
rect 5433 433 5447 447
rect 5513 613 5527 627
rect 5533 633 5547 647
rect 5593 633 5607 647
rect 5533 593 5547 607
rect 5493 473 5507 487
rect 5453 413 5467 427
rect 5433 393 5447 407
rect 5353 373 5367 387
rect 5413 373 5427 387
rect 5053 353 5067 367
rect 5053 333 5067 347
rect 5113 333 5127 347
rect 5293 353 5307 367
rect 5153 313 5167 327
rect 5093 293 5107 307
rect 4973 253 4987 267
rect 5013 253 5027 267
rect 4973 173 4987 187
rect 4753 73 4767 87
rect 4853 73 4867 87
rect 5093 193 5107 207
rect 5313 333 5327 347
rect 5353 333 5367 347
rect 5193 213 5207 227
rect 5333 273 5347 287
rect 5253 253 5267 267
rect 5213 173 5227 187
rect 5333 233 5347 247
rect 5113 153 5127 167
rect 5173 153 5187 167
rect 5193 133 5207 147
rect 5213 153 5227 167
rect 5253 153 5267 167
rect 5233 133 5247 147
rect 5133 113 5147 127
rect 5293 133 5307 147
rect 5573 573 5587 587
rect 5693 813 5707 827
rect 5673 773 5687 787
rect 5673 693 5687 707
rect 5933 873 5947 887
rect 5733 813 5747 827
rect 5753 833 5767 847
rect 5793 833 5807 847
rect 5853 853 5867 867
rect 5873 833 5887 847
rect 5773 793 5787 807
rect 5713 713 5727 727
rect 5793 773 5807 787
rect 5913 793 5927 807
rect 6033 1013 6047 1027
rect 5953 833 5967 847
rect 5993 853 6007 867
rect 5873 733 5887 747
rect 5893 733 5907 747
rect 5933 733 5947 747
rect 5853 713 5867 727
rect 5913 713 5927 727
rect 5933 713 5947 727
rect 5853 653 5867 667
rect 5713 613 5727 627
rect 5893 673 5907 687
rect 5693 593 5707 607
rect 5713 593 5727 607
rect 5633 553 5647 567
rect 5613 413 5627 427
rect 5593 353 5607 367
rect 5613 373 5627 387
rect 5513 333 5527 347
rect 5393 313 5407 327
rect 5433 313 5447 327
rect 5473 253 5487 267
rect 5373 213 5387 227
rect 5373 153 5387 167
rect 5453 173 5467 187
rect 5493 153 5507 167
rect 5133 93 5147 107
rect 4573 53 4587 67
rect 4633 53 4647 67
rect 5853 633 5867 647
rect 5913 633 5927 647
rect 5893 613 5907 627
rect 5953 693 5967 707
rect 6113 973 6127 987
rect 6093 953 6107 967
rect 6093 913 6107 927
rect 6073 833 6087 847
rect 6053 793 6067 807
rect 6013 773 6027 787
rect 6053 733 6067 747
rect 6053 693 6067 707
rect 6193 1173 6207 1187
rect 6233 1213 6247 1227
rect 6273 1213 6287 1227
rect 6233 1193 6247 1207
rect 6253 1193 6267 1207
rect 6273 1173 6287 1187
rect 6273 1113 6287 1127
rect 6253 1093 6267 1107
rect 6253 953 6267 967
rect 6153 913 6167 927
rect 6393 1613 6407 1627
rect 6373 1573 6387 1587
rect 6413 1453 6427 1467
rect 6353 1353 6367 1367
rect 6333 1273 6347 1287
rect 6393 1173 6407 1187
rect 6333 1153 6347 1167
rect 6413 1153 6427 1167
rect 6473 1593 6487 1607
rect 6513 1413 6527 1427
rect 6553 1413 6567 1427
rect 6533 1393 6547 1407
rect 6493 1293 6507 1307
rect 6533 1273 6547 1287
rect 6633 1833 6647 1847
rect 6593 1813 6607 1827
rect 6613 1793 6627 1807
rect 6593 1673 6607 1687
rect 6653 1573 6667 1587
rect 6713 2313 6727 2327
rect 6713 2293 6727 2307
rect 6693 2053 6707 2067
rect 6733 2093 6747 2107
rect 6713 1933 6727 1947
rect 6733 1913 6747 1927
rect 6693 1873 6707 1887
rect 6673 1433 6687 1447
rect 6573 1273 6587 1287
rect 6453 1133 6467 1147
rect 6333 1053 6347 1067
rect 6393 1073 6407 1087
rect 6433 1013 6447 1027
rect 6453 1013 6467 1027
rect 6513 1153 6527 1167
rect 6473 993 6487 1007
rect 6473 953 6487 967
rect 6453 873 6467 887
rect 6133 813 6147 827
rect 6253 853 6267 867
rect 6293 853 6307 867
rect 6313 853 6327 867
rect 6233 813 6247 827
rect 6213 773 6227 787
rect 6173 753 6187 767
rect 6233 753 6247 767
rect 6153 713 6167 727
rect 6193 673 6207 687
rect 5973 633 5987 647
rect 5953 613 5967 627
rect 6073 633 6087 647
rect 6113 653 6127 667
rect 6173 653 6187 667
rect 6133 633 6147 647
rect 6093 613 6107 627
rect 6153 613 6167 627
rect 6193 633 6207 647
rect 6213 633 6227 647
rect 6193 613 6207 627
rect 5973 593 5987 607
rect 5933 553 5947 567
rect 5793 473 5807 487
rect 5893 473 5907 487
rect 5893 453 5907 467
rect 5673 413 5687 427
rect 5693 413 5707 427
rect 5733 413 5747 427
rect 5813 413 5827 427
rect 5653 333 5667 347
rect 5713 353 5727 367
rect 5553 153 5567 167
rect 5613 153 5627 167
rect 5693 173 5707 187
rect 5793 353 5807 367
rect 5953 453 5967 467
rect 6033 573 6047 587
rect 6353 853 6367 867
rect 6293 833 6307 847
rect 6333 833 6347 847
rect 6313 813 6327 827
rect 6273 773 6287 787
rect 6313 733 6327 747
rect 6353 733 6367 747
rect 6253 633 6267 647
rect 6333 693 6347 707
rect 6233 593 6247 607
rect 6273 613 6287 627
rect 6313 613 6327 627
rect 6053 553 6067 567
rect 6113 493 6127 507
rect 6113 473 6127 487
rect 6053 433 6067 447
rect 5973 373 5987 387
rect 6033 373 6047 387
rect 5853 353 5867 367
rect 5813 333 5827 347
rect 5873 333 5887 347
rect 5913 333 5927 347
rect 5993 353 6007 367
rect 5973 333 5987 347
rect 5753 273 5767 287
rect 5953 313 5967 327
rect 5933 253 5947 267
rect 5933 233 5947 247
rect 5753 153 5767 167
rect 5653 113 5667 127
rect 5813 193 5827 207
rect 5853 153 5867 167
rect 5933 173 5947 187
rect 6053 353 6067 367
rect 6133 413 6147 427
rect 6253 573 6267 587
rect 6233 393 6247 407
rect 6413 833 6427 847
rect 6453 853 6467 867
rect 6433 793 6447 807
rect 6393 653 6407 667
rect 6393 593 6407 607
rect 6373 573 6387 587
rect 6373 473 6387 487
rect 6273 433 6287 447
rect 6333 433 6347 447
rect 6313 413 6327 427
rect 6293 393 6307 407
rect 6053 313 6067 327
rect 5993 293 6007 307
rect 5973 193 5987 207
rect 5953 153 5967 167
rect 5993 133 6007 147
rect 6093 273 6107 287
rect 6073 253 6087 267
rect 6133 353 6147 367
rect 6153 333 6167 347
rect 6253 353 6267 367
rect 6313 373 6327 387
rect 6453 453 6467 467
rect 6393 373 6407 387
rect 6313 333 6327 347
rect 6333 353 6347 367
rect 6393 333 6407 347
rect 6413 333 6427 347
rect 6233 313 6247 327
rect 6273 313 6287 327
rect 6313 313 6327 327
rect 6133 293 6147 307
rect 6153 253 6167 267
rect 6113 213 6127 227
rect 6213 293 6227 307
rect 6233 293 6247 307
rect 6193 213 6207 227
rect 6173 193 6187 207
rect 6113 133 6127 147
rect 6133 153 6147 167
rect 6173 153 6187 167
rect 6193 133 6207 147
rect 6153 113 6167 127
rect 6273 273 6287 287
rect 6253 253 6267 267
rect 6553 1233 6567 1247
rect 6593 1153 6607 1167
rect 6553 1133 6567 1147
rect 6673 1313 6687 1327
rect 6673 1293 6687 1307
rect 6653 1193 6667 1207
rect 6633 1173 6647 1187
rect 6553 1113 6567 1127
rect 6613 1093 6627 1107
rect 6653 1093 6667 1107
rect 6553 1073 6567 1087
rect 6533 853 6547 867
rect 6533 813 6547 827
rect 6653 1073 6667 1087
rect 6573 973 6587 987
rect 6593 973 6607 987
rect 6653 973 6667 987
rect 6573 793 6587 807
rect 6513 673 6527 687
rect 6533 673 6547 687
rect 6553 673 6567 687
rect 6513 613 6527 627
rect 6513 453 6527 467
rect 6493 333 6507 347
rect 6573 653 6587 667
rect 6573 613 6587 627
rect 6613 893 6627 907
rect 6713 1313 6727 1327
rect 6693 1253 6707 1267
rect 6733 1213 6747 1227
rect 6733 1053 6747 1067
rect 6713 1013 6727 1027
rect 6713 973 6727 987
rect 6673 893 6687 907
rect 6653 853 6667 867
rect 6653 653 6667 667
rect 6593 473 6607 487
rect 6533 373 6547 387
rect 6473 293 6487 307
rect 6313 253 6327 267
rect 6233 193 6247 207
rect 6293 193 6307 207
rect 6393 193 6407 207
rect 6413 193 6427 207
rect 6213 113 6227 127
rect 6253 153 6267 167
rect 6293 153 6307 167
rect 6313 133 6327 147
rect 6613 373 6627 387
rect 6713 233 6727 247
rect 6513 173 6527 187
rect 6553 153 6567 167
rect 6233 93 6247 107
rect 6273 93 6287 107
rect 6053 53 6067 67
rect 2773 33 2787 47
rect 2973 33 2987 47
rect 4313 33 4327 47
<< metal3 >>
rect 4407 6496 4753 6504
rect 4907 6496 5893 6504
rect 4347 6476 5113 6484
rect 5167 6476 5533 6484
rect 5556 6476 6173 6484
rect 3107 6456 3453 6464
rect 4687 6456 4913 6464
rect 5027 6456 5473 6464
rect 5556 6464 5564 6476
rect 5507 6456 5564 6464
rect 5747 6456 5793 6464
rect 6027 6456 6053 6464
rect 6167 6456 6253 6464
rect 6307 6456 6353 6464
rect 747 6436 933 6444
rect 1227 6436 1353 6444
rect 1647 6436 1673 6444
rect 2176 6436 2304 6444
rect 147 6416 153 6424
rect 167 6416 693 6424
rect 707 6416 764 6424
rect 107 6396 293 6404
rect 347 6396 413 6404
rect 447 6396 533 6404
rect 587 6396 613 6404
rect 756 6404 764 6416
rect 856 6416 1004 6424
rect 856 6404 864 6416
rect 756 6396 864 6404
rect 996 6404 1004 6416
rect 1076 6416 1173 6424
rect 1076 6404 1084 6416
rect 1187 6416 1293 6424
rect 1307 6416 1664 6424
rect 996 6396 1084 6404
rect 1416 6396 1553 6404
rect 287 6376 373 6384
rect 627 6376 793 6384
rect 827 6376 873 6384
rect 1047 6376 1193 6384
rect 1316 6384 1324 6393
rect 1207 6376 1324 6384
rect 1416 6384 1424 6396
rect 1656 6404 1664 6416
rect 1696 6416 1793 6424
rect 1696 6404 1704 6416
rect 1656 6396 1704 6404
rect 1847 6396 1973 6404
rect 2007 6396 2153 6404
rect 2176 6387 2184 6436
rect 2296 6424 2304 6436
rect 2327 6436 2493 6444
rect 2907 6436 3113 6444
rect 3187 6436 3253 6444
rect 3407 6436 4093 6444
rect 4447 6436 4553 6444
rect 4567 6436 4793 6444
rect 4947 6436 5153 6444
rect 5227 6436 5333 6444
rect 5367 6436 5493 6444
rect 5587 6436 5753 6444
rect 6047 6436 6093 6444
rect 6147 6436 6213 6444
rect 6247 6436 6513 6444
rect 6527 6436 6533 6444
rect 6607 6436 6693 6444
rect 2296 6416 2433 6424
rect 2727 6416 3193 6424
rect 3247 6416 3373 6424
rect 3507 6416 3533 6424
rect 3607 6416 3713 6424
rect 3767 6416 3973 6424
rect 4707 6416 4733 6424
rect 4767 6416 4953 6424
rect 5627 6416 5653 6424
rect 5667 6416 5693 6424
rect 5947 6416 5973 6424
rect 6367 6416 6413 6424
rect 6587 6416 6633 6424
rect 2207 6396 2233 6404
rect 2276 6387 2284 6413
rect 2367 6396 2413 6404
rect 2467 6396 2473 6404
rect 2487 6396 2573 6404
rect 3007 6396 3033 6404
rect 3216 6404 3224 6413
rect 3067 6396 3164 6404
rect 3216 6396 3264 6404
rect 1387 6376 1424 6384
rect 1507 6376 1593 6384
rect 1667 6376 1753 6384
rect 1767 6376 1913 6384
rect 2016 6376 2053 6384
rect 227 6356 353 6364
rect 367 6356 453 6364
rect 507 6356 513 6364
rect 527 6356 673 6364
rect 867 6356 913 6364
rect 1347 6356 1433 6364
rect 1547 6356 1573 6364
rect 2016 6364 2024 6376
rect 2647 6376 2673 6384
rect 2727 6376 2744 6384
rect 2736 6367 2744 6376
rect 2767 6376 2793 6384
rect 2867 6376 2904 6384
rect 1807 6356 2024 6364
rect 2087 6356 2233 6364
rect 2247 6356 2293 6364
rect 2307 6356 2333 6364
rect 2427 6356 2553 6364
rect 2787 6356 2833 6364
rect 2896 6364 2904 6376
rect 2956 6367 2964 6393
rect 3156 6387 3164 6396
rect 2987 6376 3013 6384
rect 3087 6376 3133 6384
rect 3256 6384 3264 6396
rect 3307 6396 3333 6404
rect 3356 6396 3553 6404
rect 3356 6387 3364 6396
rect 3596 6396 3633 6404
rect 3256 6376 3273 6384
rect 3596 6384 3604 6396
rect 3656 6396 3733 6404
rect 3527 6376 3604 6384
rect 3656 6384 3664 6396
rect 3827 6396 3833 6404
rect 4507 6396 4604 6404
rect 3627 6376 3664 6384
rect 3687 6376 3753 6384
rect 2896 6356 2924 6364
rect 407 6336 413 6344
rect 427 6336 813 6344
rect 2287 6336 2353 6344
rect 2367 6336 2373 6344
rect 2696 6344 2704 6353
rect 2387 6336 2773 6344
rect 2876 6344 2884 6353
rect 2876 6336 2893 6344
rect 2916 6344 2924 6356
rect 3036 6364 3044 6373
rect 3776 6367 3784 6393
rect 3816 6367 3824 6393
rect 4087 6376 4193 6384
rect 4307 6376 4444 6384
rect 3036 6356 3193 6364
rect 3207 6356 3573 6364
rect 3607 6356 3653 6364
rect 2916 6336 3153 6344
rect 3547 6336 3593 6344
rect 3807 6336 3853 6344
rect 4016 6344 4024 6373
rect 4147 6356 4213 6364
rect 4227 6356 4313 6364
rect 4327 6356 4373 6364
rect 4436 6364 4444 6376
rect 4547 6376 4573 6384
rect 4596 6384 4604 6396
rect 4636 6387 4644 6413
rect 4756 6404 4764 6413
rect 4716 6396 4764 6404
rect 4716 6387 4724 6396
rect 4787 6396 4813 6404
rect 5036 6396 5053 6404
rect 4596 6376 4613 6384
rect 4647 6376 4684 6384
rect 4436 6356 4473 6364
rect 4527 6356 4553 6364
rect 4587 6356 4653 6364
rect 4676 6364 4684 6376
rect 4767 6376 4793 6384
rect 4856 6384 4864 6393
rect 4856 6376 4893 6384
rect 5036 6384 5044 6396
rect 5227 6396 5373 6404
rect 5387 6396 5393 6404
rect 5807 6396 5844 6404
rect 4956 6376 5044 6384
rect 4956 6364 4964 6376
rect 5207 6376 5253 6384
rect 5567 6376 5633 6384
rect 5756 6384 5764 6393
rect 5687 6376 5813 6384
rect 4676 6356 4964 6364
rect 5007 6356 5133 6364
rect 4016 6336 4033 6344
rect 4127 6336 4173 6344
rect 4416 6344 4424 6353
rect 5256 6347 5264 6373
rect 5296 6347 5304 6373
rect 5396 6364 5404 6373
rect 5396 6356 5453 6364
rect 5687 6356 5733 6364
rect 5836 6364 5844 6396
rect 5887 6396 6673 6404
rect 5927 6376 5993 6384
rect 6047 6376 6153 6384
rect 6167 6376 6264 6384
rect 5816 6356 5844 6364
rect 4187 6336 4713 6344
rect 4727 6336 5233 6344
rect 5327 6336 5593 6344
rect 5607 6336 5713 6344
rect 5796 6344 5804 6353
rect 5816 6347 5824 6356
rect 5887 6356 5913 6364
rect 5967 6356 6073 6364
rect 6087 6356 6213 6364
rect 6227 6356 6233 6364
rect 6256 6364 6264 6376
rect 6287 6376 6333 6384
rect 6387 6376 6433 6384
rect 6487 6376 6524 6384
rect 6256 6356 6393 6364
rect 6407 6356 6493 6364
rect 5727 6336 5804 6344
rect 5847 6336 6113 6344
rect 6127 6336 6313 6344
rect 6327 6336 6413 6344
rect 6516 6344 6524 6376
rect 6667 6376 6733 6384
rect 6627 6356 6713 6364
rect 6496 6336 6524 6344
rect 2107 6316 2533 6324
rect 2547 6316 2793 6324
rect 3487 6316 3493 6324
rect 3507 6316 3913 6324
rect 3927 6316 4493 6324
rect 4627 6316 4993 6324
rect 5027 6316 5213 6324
rect 5987 6316 6093 6324
rect 6496 6324 6504 6336
rect 6587 6336 6673 6344
rect 6107 6316 6504 6324
rect 6667 6316 6693 6324
rect 507 6296 1073 6304
rect 2267 6296 2633 6304
rect 3127 6296 4073 6304
rect 4607 6296 4973 6304
rect 4987 6296 5033 6304
rect 5107 6296 5293 6304
rect 5307 6296 5353 6304
rect 887 6276 953 6284
rect 2027 6276 2653 6284
rect 2867 6276 2913 6284
rect 2927 6276 3173 6284
rect 3187 6276 3233 6284
rect 3247 6276 3433 6284
rect 3847 6276 4053 6284
rect 4067 6276 4893 6284
rect 5127 6276 5413 6284
rect 5427 6276 5493 6284
rect 6147 6276 6173 6284
rect 6187 6276 6553 6284
rect 2047 6256 2113 6264
rect 3127 6256 3253 6264
rect 3267 6256 3773 6264
rect 3907 6256 3993 6264
rect 4007 6256 4273 6264
rect 4727 6256 5253 6264
rect 5427 6256 5553 6264
rect 5567 6256 5613 6264
rect 5627 6256 5753 6264
rect 1907 6236 1953 6244
rect 5907 6236 6133 6244
rect 6147 6236 6433 6244
rect 4647 6216 4753 6224
rect 3147 6196 3253 6204
rect 3267 6196 3273 6204
rect 3287 6196 4173 6204
rect 4447 6196 4513 6204
rect 4567 6196 5453 6204
rect 327 6176 513 6184
rect 2547 6176 2953 6184
rect 3476 6176 3513 6184
rect 407 6156 444 6164
rect 247 6116 293 6124
rect 376 6124 384 6133
rect 347 6116 384 6124
rect 47 6096 73 6104
rect 167 6096 273 6104
rect 336 6104 344 6113
rect 336 6096 373 6104
rect 416 6104 424 6133
rect 396 6096 424 6104
rect 396 6084 404 6096
rect 327 6076 404 6084
rect 436 6084 444 6156
rect 767 6156 833 6164
rect 1007 6156 1053 6164
rect 1227 6156 1353 6164
rect 1627 6156 1713 6164
rect 2087 6156 2133 6164
rect 2607 6156 2693 6164
rect 2907 6156 3173 6164
rect 496 6136 533 6144
rect 496 6104 504 6136
rect 587 6136 684 6144
rect 527 6116 553 6124
rect 636 6116 653 6124
rect 496 6096 513 6104
rect 616 6104 624 6113
rect 567 6096 624 6104
rect 427 6076 444 6084
rect 467 6076 553 6084
rect 636 6084 644 6116
rect 676 6124 684 6136
rect 1607 6136 1644 6144
rect 676 6116 744 6124
rect 736 6107 744 6116
rect 827 6116 913 6124
rect 967 6116 1013 6124
rect 1107 6116 1144 6124
rect 667 6096 713 6104
rect 816 6104 824 6113
rect 1136 6107 1144 6116
rect 1636 6124 1644 6136
rect 2067 6136 2133 6144
rect 2207 6136 2293 6144
rect 2316 6136 2413 6144
rect 2316 6127 2324 6136
rect 2747 6136 2813 6144
rect 2827 6136 3013 6144
rect 3236 6144 3244 6153
rect 3476 6147 3484 6176
rect 4467 6176 4873 6184
rect 6256 6176 6313 6184
rect 3527 6156 3573 6164
rect 4347 6156 4373 6164
rect 4476 6156 4553 6164
rect 3227 6136 3244 6144
rect 3307 6136 3373 6144
rect 3496 6127 3504 6153
rect 3607 6136 3633 6144
rect 3647 6136 3713 6144
rect 3767 6136 3793 6144
rect 1296 6116 1424 6124
rect 1636 6116 1684 6124
rect 796 6096 824 6104
rect 956 6096 1024 6104
rect 636 6076 693 6084
rect 796 6084 804 6096
rect 956 6084 964 6096
rect 787 6076 804 6084
rect 916 6076 964 6084
rect 1016 6084 1024 6096
rect 1276 6104 1284 6113
rect 1296 6107 1304 6116
rect 1247 6096 1284 6104
rect 1416 6104 1424 6116
rect 1336 6096 1404 6104
rect 1416 6096 1433 6104
rect 1336 6084 1344 6096
rect 1016 6076 1344 6084
rect 127 6056 373 6064
rect 916 6064 924 6076
rect 407 6056 924 6064
rect 947 6056 993 6064
rect 1007 6056 1173 6064
rect 1187 6056 1373 6064
rect 1396 6064 1404 6096
rect 1447 6096 1484 6104
rect 1427 6076 1453 6084
rect 1476 6084 1484 6096
rect 1567 6096 1633 6104
rect 1476 6076 1533 6084
rect 1556 6076 1593 6084
rect 1396 6056 1513 6064
rect 1556 6064 1564 6076
rect 1676 6084 1684 6116
rect 1696 6116 1753 6124
rect 1696 6107 1704 6116
rect 1807 6116 1833 6124
rect 1887 6116 1933 6124
rect 1947 6116 1973 6124
rect 2087 6116 2093 6124
rect 2107 6116 2153 6124
rect 2487 6116 2533 6124
rect 2927 6116 2953 6124
rect 3127 6116 3193 6124
rect 1727 6096 1773 6104
rect 2036 6096 2104 6104
rect 2036 6087 2044 6096
rect 1676 6076 1753 6084
rect 1787 6076 1793 6084
rect 1807 6076 1993 6084
rect 2096 6084 2104 6096
rect 2236 6104 2244 6113
rect 2187 6096 2244 6104
rect 2387 6096 2513 6104
rect 2527 6096 2613 6104
rect 2636 6087 2644 6113
rect 2767 6096 2793 6104
rect 2896 6096 2953 6104
rect 2896 6087 2904 6096
rect 3116 6087 3124 6113
rect 3336 6104 3344 6113
rect 3336 6096 3513 6104
rect 3527 6096 3593 6104
rect 2096 6076 2233 6084
rect 2667 6076 2833 6084
rect 2947 6076 3013 6084
rect 3467 6076 3513 6084
rect 3527 6076 3593 6084
rect 3627 6076 3653 6084
rect 1527 6056 1564 6064
rect 1587 6056 1753 6064
rect 1767 6056 1913 6064
rect 1927 6056 2213 6064
rect 2227 6056 2413 6064
rect 2447 6056 2593 6064
rect 2607 6056 2953 6064
rect 2987 6056 3033 6064
rect 3047 6056 3133 6064
rect 3327 6056 3553 6064
rect 3676 6064 3684 6113
rect 3747 6096 3773 6104
rect 3816 6104 3824 6153
rect 4267 6136 4293 6144
rect 4476 6144 4484 6156
rect 4716 6156 4733 6164
rect 4336 6136 4484 6144
rect 3856 6107 3864 6133
rect 3807 6096 3824 6104
rect 3996 6087 4004 6113
rect 4036 6087 4044 6133
rect 4196 6116 4233 6124
rect 4056 6104 4064 6113
rect 4056 6096 4093 6104
rect 4176 6104 4184 6113
rect 4196 6107 4204 6116
rect 4336 6124 4344 6136
rect 4576 6136 4593 6144
rect 4327 6116 4344 6124
rect 4496 6107 4504 6133
rect 4576 6107 4584 6136
rect 4607 6116 4673 6124
rect 4716 6124 4724 6156
rect 5047 6156 5213 6164
rect 5227 6156 5273 6164
rect 5336 6156 5404 6164
rect 4747 6136 4873 6144
rect 5096 6136 5113 6144
rect 4716 6116 4764 6124
rect 4156 6096 4184 6104
rect 4156 6087 4164 6096
rect 4267 6096 4313 6104
rect 4327 6096 4353 6104
rect 3767 6076 3873 6084
rect 4067 6076 4113 6084
rect 4596 6084 4604 6113
rect 4616 6096 4653 6104
rect 4616 6087 4624 6096
rect 4667 6096 4733 6104
rect 4427 6076 4604 6084
rect 4756 6084 4764 6116
rect 4847 6116 4933 6124
rect 4687 6076 4764 6084
rect 3567 6056 4073 6064
rect 4127 6056 4213 6064
rect 4447 6056 4773 6064
rect 4796 6064 4804 6113
rect 5096 6107 5104 6136
rect 5336 6124 5344 6156
rect 5396 6144 5404 6156
rect 5547 6156 5713 6164
rect 5827 6156 5953 6164
rect 5967 6156 6053 6164
rect 6147 6156 6164 6164
rect 6156 6147 6164 6156
rect 6207 6156 6233 6164
rect 5367 6136 5384 6144
rect 5396 6136 5433 6144
rect 5336 6116 5353 6124
rect 4927 6096 4993 6104
rect 5116 6087 5124 6113
rect 5376 6107 5384 6136
rect 5607 6136 5644 6144
rect 5636 6127 5644 6136
rect 5707 6136 5853 6144
rect 6176 6144 6184 6153
rect 6256 6147 6264 6176
rect 6396 6156 6453 6164
rect 6176 6136 6244 6144
rect 5487 6116 5613 6124
rect 5687 6116 5713 6124
rect 5736 6116 5773 6124
rect 5167 6096 5213 6104
rect 5736 6104 5744 6116
rect 5787 6116 5804 6124
rect 5476 6096 5744 6104
rect 5796 6104 5804 6116
rect 5827 6116 5873 6124
rect 5976 6107 5984 6133
rect 6236 6127 6244 6136
rect 6007 6116 6173 6124
rect 6276 6124 6284 6153
rect 6396 6147 6404 6156
rect 6307 6136 6384 6144
rect 6376 6127 6384 6136
rect 6447 6136 6513 6144
rect 6267 6116 6284 6124
rect 6487 6116 6553 6124
rect 5796 6096 5833 6104
rect 4827 6076 4873 6084
rect 4887 6076 4913 6084
rect 5207 6076 5333 6084
rect 5476 6084 5484 6096
rect 6276 6096 6453 6104
rect 5347 6076 5484 6084
rect 5507 6076 5593 6084
rect 5627 6076 5693 6084
rect 5807 6076 5853 6084
rect 5947 6076 6033 6084
rect 6087 6076 6153 6084
rect 6276 6084 6284 6096
rect 6187 6076 6284 6084
rect 6387 6076 6493 6084
rect 4796 6056 4893 6064
rect 4907 6056 5073 6064
rect 5087 6056 5273 6064
rect 5767 6056 5933 6064
rect 6247 6056 6273 6064
rect 6507 6056 6533 6064
rect 527 6036 613 6044
rect 707 6036 813 6044
rect 907 6036 1153 6044
rect 1367 6036 1473 6044
rect 1487 6036 1673 6044
rect 2087 6036 2113 6044
rect 2207 6036 2273 6044
rect 2727 6036 3073 6044
rect 4007 6036 4093 6044
rect 4107 6036 4173 6044
rect 4707 6036 4753 6044
rect 4767 6036 5173 6044
rect 5667 6036 5793 6044
rect 6167 6036 6313 6044
rect 6427 6036 6573 6044
rect 1667 6016 1693 6024
rect 3407 6016 3533 6024
rect 3547 6016 3553 6024
rect 3567 6016 3693 6024
rect 3707 6016 3833 6024
rect 3947 6016 3993 6024
rect 4147 6016 4433 6024
rect 6107 6016 6253 6024
rect 6267 6016 6433 6024
rect 507 5996 613 6004
rect 627 5996 1193 6004
rect 1236 5996 1253 6004
rect 547 5976 653 5984
rect 767 5976 793 5984
rect 1236 5984 1244 5996
rect 1667 5996 1793 6004
rect 2207 5996 2373 6004
rect 2947 5996 3853 6004
rect 3867 5996 5613 6004
rect 5627 5996 6333 6004
rect 807 5976 1244 5984
rect 1727 5976 1733 5984
rect 1747 5976 1813 5984
rect 1827 5976 1913 5984
rect 1927 5976 2333 5984
rect 3687 5976 3973 5984
rect 4067 5976 4073 5984
rect 4087 5976 4713 5984
rect 4987 5976 5193 5984
rect 5927 5976 6213 5984
rect 6347 5976 6593 5984
rect 407 5956 433 5964
rect 807 5956 893 5964
rect 1007 5956 1153 5964
rect 1167 5956 1233 5964
rect 1756 5956 1773 5964
rect 327 5936 413 5944
rect 527 5936 593 5944
rect 867 5936 1044 5944
rect 527 5916 544 5924
rect 207 5896 333 5904
rect 416 5887 424 5913
rect 536 5907 544 5916
rect 587 5916 633 5924
rect 676 5924 684 5933
rect 656 5916 684 5924
rect 656 5887 664 5916
rect 707 5916 733 5924
rect 776 5924 784 5933
rect 776 5916 804 5924
rect -24 5876 13 5884
rect 67 5876 93 5884
rect 247 5876 293 5884
rect 347 5876 373 5884
rect 467 5876 633 5884
rect 796 5884 804 5916
rect 827 5916 873 5924
rect 987 5916 1013 5924
rect 1036 5907 1044 5936
rect 1067 5916 1073 5924
rect 1127 5916 1213 5924
rect 1367 5916 1473 5924
rect 1647 5916 1673 5924
rect 947 5896 973 5904
rect 1076 5904 1084 5913
rect 1696 5907 1704 5933
rect 1756 5924 1764 5956
rect 1827 5956 2013 5964
rect 2196 5956 2233 5964
rect 2007 5936 2053 5944
rect 2196 5944 2204 5956
rect 2276 5956 2353 5964
rect 2176 5936 2204 5944
rect 1756 5916 1784 5924
rect 1776 5907 1784 5916
rect 1807 5916 1873 5924
rect 1936 5916 1953 5924
rect 1936 5907 1944 5916
rect 2176 5924 2184 5936
rect 1967 5916 2184 5924
rect 2216 5907 2224 5933
rect 2256 5924 2264 5933
rect 2236 5916 2264 5924
rect 2236 5907 2244 5916
rect 1076 5896 1093 5904
rect 1547 5896 1573 5904
rect 1856 5896 1893 5904
rect 796 5876 813 5884
rect 827 5876 913 5884
rect 1507 5876 1553 5884
rect 1607 5876 1833 5884
rect 147 5856 213 5864
rect 227 5856 573 5864
rect 787 5856 873 5864
rect 1067 5856 1093 5864
rect 1547 5856 1813 5864
rect 1856 5864 1864 5896
rect 1967 5896 1993 5904
rect 2007 5896 2073 5904
rect 2127 5896 2164 5904
rect 1887 5876 1913 5884
rect 1947 5876 1973 5884
rect 1987 5876 2093 5884
rect 2156 5884 2164 5896
rect 2276 5904 2284 5956
rect 2987 5956 2993 5964
rect 3007 5956 3373 5964
rect 3616 5956 3853 5964
rect 2467 5936 2513 5944
rect 2527 5936 2553 5944
rect 2567 5936 2613 5944
rect 2627 5936 2713 5944
rect 2787 5936 2873 5944
rect 2887 5936 3093 5944
rect 3127 5936 3393 5944
rect 3427 5936 3493 5944
rect 3616 5944 3624 5956
rect 3907 5956 3953 5964
rect 3967 5956 4453 5964
rect 4707 5956 4753 5964
rect 5027 5956 5053 5964
rect 5207 5956 5373 5964
rect 5687 5956 5713 5964
rect 5747 5956 5833 5964
rect 6327 5956 6393 5964
rect 3596 5936 3624 5944
rect 2296 5907 2304 5933
rect 2327 5916 2353 5924
rect 2587 5916 2624 5924
rect 2616 5907 2624 5916
rect 2827 5916 2893 5924
rect 2927 5916 3013 5924
rect 3087 5916 3153 5924
rect 3187 5916 3273 5924
rect 3327 5916 3333 5924
rect 3347 5916 3453 5924
rect 3476 5916 3573 5924
rect 2267 5896 2284 5904
rect 2316 5896 2333 5904
rect 2316 5884 2324 5896
rect 2507 5896 2593 5904
rect 2687 5896 2733 5904
rect 2807 5896 2824 5904
rect 2156 5876 2324 5884
rect 2447 5876 2473 5884
rect 2707 5876 2713 5884
rect 2727 5876 2753 5884
rect 2816 5884 2824 5896
rect 2907 5896 2944 5904
rect 2816 5876 2853 5884
rect 2936 5884 2944 5896
rect 3036 5904 3044 5913
rect 3007 5896 3044 5904
rect 3187 5896 3253 5904
rect 3307 5896 3353 5904
rect 3476 5904 3484 5916
rect 3596 5907 3604 5936
rect 3687 5936 3744 5944
rect 3627 5916 3653 5924
rect 3667 5916 3713 5924
rect 3736 5907 3744 5936
rect 3967 5936 3984 5944
rect 3867 5916 3953 5924
rect 3976 5907 3984 5936
rect 4167 5936 4184 5944
rect 4016 5924 4024 5933
rect 4016 5916 4153 5924
rect 4176 5924 4184 5936
rect 4207 5936 4224 5944
rect 4216 5924 4224 5936
rect 4476 5936 4553 5944
rect 4176 5916 4204 5924
rect 4216 5916 4253 5924
rect 4196 5907 4204 5916
rect 4387 5916 4424 5924
rect 3407 5896 3484 5904
rect 3647 5896 3693 5904
rect 4027 5896 4073 5904
rect 4096 5896 4113 5904
rect 2936 5876 2953 5884
rect 3136 5884 3144 5893
rect 3107 5876 3144 5884
rect 3487 5876 3613 5884
rect 3716 5884 3724 5893
rect 3696 5876 3773 5884
rect 1856 5856 2393 5864
rect 2567 5856 2633 5864
rect 2647 5856 2653 5864
rect 2796 5864 2804 5873
rect 2896 5864 2904 5873
rect 2667 5856 3053 5864
rect 3096 5864 3104 5873
rect 3087 5856 3104 5864
rect 3156 5864 3164 5873
rect 3156 5856 3173 5864
rect 3547 5856 3653 5864
rect 3696 5864 3704 5876
rect 3687 5856 3704 5864
rect 3876 5864 3884 5893
rect 4096 5884 4104 5896
rect 4287 5896 4353 5904
rect 4367 5896 4393 5904
rect 3947 5876 4104 5884
rect 4116 5876 4133 5884
rect 4116 5867 4124 5876
rect 4147 5876 4173 5884
rect 4236 5884 4244 5893
rect 4187 5876 4244 5884
rect 4416 5884 4424 5916
rect 4396 5876 4424 5884
rect 4436 5884 4444 5913
rect 4476 5907 4484 5936
rect 4636 5936 4744 5944
rect 4636 5924 4644 5936
rect 4507 5916 4644 5924
rect 4736 5924 4744 5936
rect 5067 5936 5084 5944
rect 4916 5924 4924 5933
rect 4667 5916 4704 5924
rect 4736 5916 4924 5924
rect 5036 5924 5044 5933
rect 5036 5916 5064 5924
rect 4696 5904 4704 5916
rect 4756 5907 4764 5916
rect 5056 5907 5064 5916
rect 4696 5896 4733 5904
rect 4827 5896 4853 5904
rect 4867 5896 4973 5904
rect 4987 5896 5033 5904
rect 4436 5876 4453 5884
rect 3876 5856 3953 5864
rect 4256 5864 4264 5873
rect 4256 5856 4273 5864
rect 4396 5864 4404 5876
rect 4787 5876 4893 5884
rect 5076 5884 5084 5936
rect 5247 5936 5364 5944
rect 5107 5916 5133 5924
rect 5356 5924 5364 5936
rect 5467 5936 5493 5944
rect 5507 5936 5633 5944
rect 5727 5936 5773 5944
rect 5887 5936 5933 5944
rect 5987 5936 6033 5944
rect 6087 5936 6133 5944
rect 6187 5936 6233 5944
rect 6487 5936 6633 5944
rect 5356 5916 5513 5924
rect 5527 5916 5573 5924
rect 5616 5916 5653 5924
rect 5176 5896 5213 5904
rect 5176 5887 5184 5896
rect 5336 5904 5344 5913
rect 5236 5896 5344 5904
rect 5236 5887 5244 5896
rect 5407 5896 5553 5904
rect 5616 5904 5624 5916
rect 5696 5924 5704 5933
rect 5696 5916 5724 5924
rect 5567 5896 5624 5904
rect 5647 5896 5693 5904
rect 5047 5876 5084 5884
rect 5107 5876 5113 5884
rect 5127 5876 5153 5884
rect 5267 5876 5333 5884
rect 5367 5876 5473 5884
rect 5667 5876 5693 5884
rect 5716 5884 5724 5916
rect 5767 5916 5873 5924
rect 5887 5916 5893 5924
rect 6016 5904 6024 5913
rect 6016 5896 6053 5904
rect 5716 5876 5753 5884
rect 5956 5884 5964 5893
rect 6096 5887 6104 5913
rect 6156 5907 6164 5933
rect 6236 5916 6293 5924
rect 6236 5887 6244 5916
rect 6367 5916 6453 5924
rect 6467 5916 6484 5924
rect 6336 5904 6344 5913
rect 6476 5904 6484 5916
rect 6336 5896 6364 5904
rect 6476 5896 6513 5904
rect 5767 5876 5964 5884
rect 6127 5876 6233 5884
rect 4367 5856 4404 5864
rect 4427 5856 4853 5864
rect 4996 5864 5004 5873
rect 4907 5856 5073 5864
rect 5327 5856 5453 5864
rect 5507 5856 5573 5864
rect 5647 5856 5973 5864
rect 6256 5864 6264 5893
rect 6356 5887 6364 5896
rect 6627 5896 6693 5904
rect 6536 5884 6544 5893
rect 6407 5876 6544 5884
rect 6256 5856 6313 5864
rect 6327 5856 6384 5864
rect 507 5836 673 5844
rect 987 5836 1453 5844
rect 2047 5836 2373 5844
rect 2407 5836 2593 5844
rect 2967 5836 3033 5844
rect 3207 5836 3293 5844
rect 3647 5836 3844 5844
rect 1907 5816 1953 5824
rect 2247 5816 3813 5824
rect 3836 5824 3844 5836
rect 3947 5836 4293 5844
rect 4707 5836 4733 5844
rect 4747 5836 5033 5844
rect 5127 5836 5433 5844
rect 5447 5836 5773 5844
rect 5807 5836 5833 5844
rect 5907 5836 6093 5844
rect 6376 5844 6384 5856
rect 6536 5864 6544 5876
rect 6567 5876 6573 5884
rect 6587 5876 6593 5884
rect 6467 5856 6544 5864
rect 6376 5836 6553 5844
rect 3836 5816 4053 5824
rect 4196 5816 5273 5824
rect 3187 5796 3433 5804
rect 4196 5804 4204 5816
rect 5527 5816 5853 5824
rect 5867 5816 5913 5824
rect 6387 5816 6593 5824
rect 4027 5796 4204 5804
rect 4227 5796 4393 5804
rect 5167 5796 5233 5804
rect 5247 5796 5533 5804
rect 5627 5796 6213 5804
rect 6267 5796 6653 5804
rect 4167 5776 4253 5784
rect 4267 5776 4353 5784
rect 5547 5776 6273 5784
rect 6287 5776 6333 5784
rect 3987 5756 4093 5764
rect 4107 5756 4373 5764
rect 4667 5756 5313 5764
rect 5447 5756 6113 5764
rect 6347 5756 6413 5764
rect 3947 5736 4373 5744
rect 4387 5736 4453 5744
rect 4547 5736 4653 5744
rect 4867 5736 4973 5744
rect 5287 5736 5973 5744
rect 747 5716 913 5724
rect 2387 5716 2873 5724
rect 4067 5716 4273 5724
rect 4287 5716 4393 5724
rect 4627 5716 4793 5724
rect 4807 5716 4873 5724
rect 4887 5716 5353 5724
rect 5407 5716 5933 5724
rect 6507 5716 6613 5724
rect 687 5696 953 5704
rect 967 5696 1233 5704
rect 2007 5696 2033 5704
rect 2047 5696 2613 5704
rect 2687 5696 2733 5704
rect 2827 5696 2833 5704
rect 2847 5696 2973 5704
rect 2987 5696 3073 5704
rect 4147 5696 4333 5704
rect 4347 5696 4493 5704
rect 4507 5696 4513 5704
rect 4527 5696 4633 5704
rect 4647 5696 4833 5704
rect 4847 5696 4853 5704
rect 5427 5696 5573 5704
rect 5667 5696 5893 5704
rect 5947 5696 6013 5704
rect 6187 5696 6273 5704
rect 6367 5696 6524 5704
rect 616 5676 633 5684
rect -24 5644 -16 5664
rect 476 5656 513 5664
rect 476 5644 484 5656
rect 547 5656 564 5664
rect -24 5636 4 5644
rect -4 5624 4 5636
rect 456 5636 484 5644
rect -24 5604 -16 5624
rect -4 5616 33 5624
rect 267 5616 313 5624
rect 456 5624 464 5636
rect 556 5644 564 5656
rect 556 5636 584 5644
rect 447 5616 464 5624
rect -24 5596 113 5604
rect 496 5604 504 5633
rect 467 5596 504 5604
rect 576 5604 584 5636
rect 596 5627 604 5653
rect 527 5596 584 5604
rect 616 5604 624 5676
rect 656 5676 704 5684
rect 656 5664 664 5676
rect 647 5656 664 5664
rect 676 5644 684 5653
rect 636 5636 684 5644
rect 696 5644 704 5676
rect 1047 5676 1113 5684
rect 1887 5676 1993 5684
rect 2107 5676 2133 5684
rect 2187 5676 2213 5684
rect 2227 5676 2273 5684
rect 2427 5676 2433 5684
rect 2447 5676 4033 5684
rect 4056 5676 4233 5684
rect 696 5636 793 5644
rect 636 5627 644 5636
rect 816 5627 824 5673
rect 1987 5656 2013 5664
rect 2147 5656 2233 5664
rect 2307 5656 2353 5664
rect 2756 5656 2773 5664
rect 1007 5636 1033 5644
rect 1307 5636 1404 5644
rect 887 5616 933 5624
rect 676 5604 684 5613
rect 616 5596 684 5604
rect 747 5596 833 5604
rect 1096 5604 1104 5613
rect 1136 5607 1144 5633
rect 1276 5624 1284 5633
rect 1276 5616 1313 5624
rect 1396 5624 1404 5636
rect 1447 5636 1673 5644
rect 1396 5616 1464 5624
rect 1007 5596 1104 5604
rect 1247 5596 1333 5604
rect 1367 5596 1433 5604
rect 1456 5604 1464 5616
rect 1607 5616 1733 5624
rect 1456 5596 1553 5604
rect 467 5576 693 5584
rect 707 5576 1013 5584
rect 1067 5576 1193 5584
rect 1227 5576 1393 5584
rect 1407 5576 1453 5584
rect 1756 5584 1764 5633
rect 1896 5627 1904 5653
rect 2756 5647 2764 5656
rect 2787 5656 2944 5664
rect 1967 5636 1993 5644
rect 2156 5636 2173 5644
rect 2156 5627 2164 5636
rect 2936 5644 2944 5656
rect 3067 5656 3373 5664
rect 3427 5656 3473 5664
rect 3627 5656 3633 5664
rect 3647 5656 3733 5664
rect 4056 5664 4064 5676
rect 4276 5676 4313 5684
rect 3787 5656 4064 5664
rect 4176 5656 4193 5664
rect 2936 5636 2993 5644
rect 3007 5636 3053 5644
rect 3267 5636 3273 5644
rect 3287 5636 3313 5644
rect 3476 5636 3553 5644
rect 1776 5616 1833 5624
rect 1776 5607 1784 5616
rect 2207 5616 2253 5624
rect 2587 5616 2653 5624
rect 2747 5616 2833 5624
rect 3096 5624 3104 5633
rect 3047 5616 3104 5624
rect 3127 5616 3153 5624
rect 1927 5596 1993 5604
rect 2016 5596 2173 5604
rect 2016 5584 2024 5596
rect 2627 5596 2673 5604
rect 3027 5596 3073 5604
rect 3087 5596 3193 5604
rect 3216 5604 3224 5633
rect 3367 5616 3453 5624
rect 3476 5624 3484 5636
rect 3816 5636 3873 5644
rect 3467 5616 3484 5624
rect 3507 5616 3613 5624
rect 3687 5616 3713 5624
rect 3816 5624 3824 5636
rect 3807 5616 3824 5624
rect 3907 5616 3953 5624
rect 3216 5596 3273 5604
rect 3347 5596 3573 5604
rect 3587 5596 3613 5604
rect 3707 5596 3733 5604
rect 4116 5604 4124 5653
rect 4176 5627 4184 5656
rect 4276 5664 4284 5676
rect 4607 5676 5184 5684
rect 4256 5656 4284 5664
rect 4207 5636 4233 5644
rect 4256 5624 4264 5656
rect 4307 5656 4353 5664
rect 4407 5656 4544 5664
rect 4416 5647 4424 5656
rect 4256 5616 4293 5624
rect 4387 5616 4433 5624
rect 4047 5596 4124 5604
rect 4167 5596 4333 5604
rect 4456 5604 4464 5633
rect 4536 5624 4544 5656
rect 4567 5656 4593 5664
rect 4716 5656 4733 5664
rect 4627 5636 4693 5644
rect 4716 5627 4724 5656
rect 4767 5656 4824 5664
rect 4747 5636 4793 5644
rect 4816 5644 4824 5656
rect 4956 5656 5013 5664
rect 4956 5647 4964 5656
rect 5036 5656 5093 5664
rect 4816 5636 4953 5644
rect 4536 5616 4593 5624
rect 4447 5596 4464 5604
rect 4487 5596 4613 5604
rect 4736 5604 4744 5633
rect 5036 5627 5044 5656
rect 5067 5636 5093 5644
rect 5116 5627 5124 5653
rect 5176 5647 5184 5676
rect 5196 5676 5393 5684
rect 5196 5667 5204 5676
rect 5567 5676 5593 5684
rect 5616 5676 5633 5684
rect 5207 5656 5253 5664
rect 5616 5664 5624 5676
rect 5967 5676 6093 5684
rect 6227 5676 6453 5684
rect 5607 5656 5624 5664
rect 5707 5656 5724 5664
rect 5407 5636 5453 5644
rect 4787 5616 5024 5624
rect 4736 5596 4793 5604
rect 4867 5596 4953 5604
rect 5016 5604 5024 5616
rect 5147 5616 5213 5624
rect 5496 5624 5504 5633
rect 5516 5627 5524 5653
rect 5716 5627 5724 5656
rect 5836 5656 5953 5664
rect 5367 5616 5504 5624
rect 5607 5616 5693 5624
rect 5016 5596 5053 5604
rect 5107 5596 5153 5604
rect 5187 5596 5253 5604
rect 5316 5596 5373 5604
rect 1756 5576 2024 5584
rect 2127 5576 2213 5584
rect 2227 5576 2233 5584
rect 3187 5576 3293 5584
rect 3307 5576 3593 5584
rect 3607 5576 3744 5584
rect 487 5556 1173 5564
rect 1187 5556 1253 5564
rect 1887 5556 2073 5564
rect 3047 5556 3113 5564
rect 3127 5556 3653 5564
rect 3667 5556 3713 5564
rect 3736 5564 3744 5576
rect 3827 5576 4033 5584
rect 4207 5576 4273 5584
rect 4747 5576 4813 5584
rect 4907 5576 4933 5584
rect 4956 5576 4993 5584
rect 3736 5556 4073 5564
rect 4247 5556 4313 5564
rect 4587 5556 4753 5564
rect 4787 5556 4853 5564
rect 4956 5564 4964 5576
rect 5027 5576 5053 5584
rect 5316 5584 5324 5596
rect 5387 5596 5473 5604
rect 5507 5596 5533 5604
rect 5716 5604 5724 5613
rect 5667 5596 5724 5604
rect 5247 5576 5324 5584
rect 5347 5576 5633 5584
rect 5736 5584 5744 5633
rect 5756 5624 5764 5653
rect 5836 5644 5844 5656
rect 6007 5656 6044 5664
rect 5787 5636 5844 5644
rect 5756 5616 5873 5624
rect 5787 5596 5853 5604
rect 5896 5604 5904 5633
rect 5887 5596 5904 5604
rect 5936 5604 5944 5633
rect 5936 5596 5953 5604
rect 5976 5596 5993 5604
rect 5647 5576 5744 5584
rect 5767 5576 5833 5584
rect 5976 5584 5984 5596
rect 6036 5604 6044 5656
rect 6247 5656 6313 5664
rect 6347 5656 6404 5664
rect 6327 5636 6373 5644
rect 6056 5607 6064 5633
rect 6087 5616 6153 5624
rect 6256 5624 6264 5633
rect 6187 5616 6264 5624
rect 6276 5607 6284 5633
rect 6316 5607 6324 5633
rect 6396 5624 6404 5656
rect 6476 5664 6484 5673
rect 6447 5656 6484 5664
rect 6516 5644 6524 5696
rect 6547 5696 6604 5704
rect 6576 5644 6584 5673
rect 6596 5667 6604 5696
rect 6516 5636 6544 5644
rect 6576 5636 6593 5644
rect 6536 5627 6544 5636
rect 6347 5616 6404 5624
rect 6616 5624 6624 5673
rect 6567 5616 6624 5624
rect 6027 5596 6044 5604
rect 6387 5596 6453 5604
rect 5927 5576 5984 5584
rect 6007 5576 6113 5584
rect 6307 5576 6393 5584
rect 6407 5576 6493 5584
rect 4927 5556 4964 5564
rect 5067 5556 5313 5564
rect 5467 5556 5793 5564
rect 5807 5556 6053 5564
rect 6067 5556 6133 5564
rect 6367 5556 6433 5564
rect 447 5536 533 5544
rect 567 5536 593 5544
rect 747 5536 953 5544
rect 987 5536 1093 5544
rect 1107 5536 1113 5544
rect 1827 5536 2473 5544
rect 2547 5536 2593 5544
rect 2967 5536 3033 5544
rect 3367 5536 3413 5544
rect 3687 5536 3793 5544
rect 3947 5536 3993 5544
rect 4007 5536 4433 5544
rect 4527 5536 4633 5544
rect 4787 5536 5233 5544
rect 5267 5536 5393 5544
rect 5487 5536 5633 5544
rect 5667 5536 5713 5544
rect 5747 5536 5793 5544
rect 6067 5536 6293 5544
rect 6347 5536 6613 5544
rect 627 5516 644 5524
rect 507 5496 613 5504
rect 636 5504 644 5516
rect 927 5516 973 5524
rect 987 5516 1073 5524
rect 2227 5516 2253 5524
rect 2267 5516 2493 5524
rect 2507 5516 2633 5524
rect 2647 5516 2753 5524
rect 3027 5516 3913 5524
rect 4227 5516 4273 5524
rect 4567 5516 4933 5524
rect 4947 5516 5073 5524
rect 5087 5516 5213 5524
rect 5287 5516 5353 5524
rect 5407 5516 5653 5524
rect 5707 5516 5993 5524
rect 6027 5516 6093 5524
rect 6147 5516 6173 5524
rect 6287 5516 6413 5524
rect 6427 5516 6513 5524
rect 636 5496 693 5504
rect 2467 5496 2733 5504
rect 2747 5496 2853 5504
rect 2867 5496 5573 5504
rect 5687 5496 5773 5504
rect 5807 5496 5893 5504
rect 6047 5496 6293 5504
rect 6527 5496 6633 5504
rect 347 5476 713 5484
rect 887 5476 913 5484
rect 1087 5476 1153 5484
rect 2007 5476 2273 5484
rect 2367 5476 2404 5484
rect 127 5456 173 5464
rect 187 5456 273 5464
rect 407 5456 513 5464
rect 527 5456 793 5464
rect 1036 5456 1293 5464
rect 167 5436 353 5444
rect 536 5436 593 5444
rect 47 5416 93 5424
rect 287 5416 364 5424
rect 96 5404 104 5413
rect 96 5396 253 5404
rect 356 5404 364 5416
rect 536 5407 544 5436
rect 607 5436 613 5444
rect 636 5436 653 5444
rect 636 5424 644 5436
rect 1036 5444 1044 5456
rect 1307 5456 1313 5464
rect 1667 5456 1693 5464
rect 1747 5456 1773 5464
rect 1787 5456 1833 5464
rect 1907 5456 1984 5464
rect 776 5436 1044 5444
rect 776 5424 784 5436
rect 1067 5436 1144 5444
rect 1136 5427 1144 5436
rect 1167 5436 1353 5444
rect 1547 5436 1713 5444
rect 1807 5436 1853 5444
rect 1927 5436 1953 5444
rect 1976 5444 1984 5456
rect 2087 5456 2153 5464
rect 2327 5456 2373 5464
rect 1976 5436 2033 5444
rect 556 5416 644 5424
rect 736 5416 784 5424
rect 556 5407 564 5416
rect 736 5407 744 5416
rect 847 5416 944 5424
rect 356 5396 413 5404
rect 427 5396 453 5404
rect 836 5404 844 5413
rect 816 5396 844 5404
rect 936 5404 944 5416
rect 1027 5416 1124 5424
rect 936 5396 1033 5404
rect 816 5387 824 5396
rect 1116 5404 1124 5416
rect 1687 5416 1733 5424
rect 1116 5396 1173 5404
rect 307 5376 573 5384
rect 587 5376 593 5384
rect 687 5376 693 5384
rect 707 5376 773 5384
rect 927 5376 1233 5384
rect 327 5356 373 5364
rect 387 5356 413 5364
rect 547 5356 613 5364
rect 787 5356 853 5364
rect 1496 5364 1504 5413
rect 1527 5396 1573 5404
rect 1667 5396 1693 5404
rect 1756 5404 1764 5433
rect 1787 5416 1873 5424
rect 2127 5416 2173 5424
rect 2336 5424 2344 5433
rect 2307 5416 2344 5424
rect 2376 5424 2384 5433
rect 2367 5416 2384 5424
rect 1756 5396 1784 5404
rect 1616 5384 1624 5393
rect 1616 5376 1673 5384
rect 1776 5384 1784 5396
rect 1867 5396 1933 5404
rect 2147 5396 2153 5404
rect 2167 5396 2193 5404
rect 2396 5404 2404 5476
rect 2556 5476 2604 5484
rect 2447 5456 2453 5464
rect 2467 5456 2533 5464
rect 2556 5427 2564 5476
rect 2596 5464 2604 5476
rect 2627 5476 2653 5484
rect 2967 5476 3193 5484
rect 3387 5476 3433 5484
rect 3447 5476 3473 5484
rect 3487 5476 3633 5484
rect 3647 5476 4533 5484
rect 4807 5476 5033 5484
rect 5447 5476 5673 5484
rect 5787 5476 6073 5484
rect 6167 5476 6273 5484
rect 6427 5476 6533 5484
rect 2596 5456 2893 5464
rect 2596 5427 2604 5456
rect 2956 5456 2973 5464
rect 2647 5436 2933 5444
rect 2827 5416 2893 5424
rect 2227 5396 2404 5404
rect 2727 5396 2813 5404
rect 2956 5404 2964 5456
rect 3036 5456 3193 5464
rect 3036 5427 3044 5456
rect 3207 5456 3233 5464
rect 3247 5456 3413 5464
rect 3587 5456 3833 5464
rect 3867 5456 3953 5464
rect 4027 5456 4033 5464
rect 4047 5456 4113 5464
rect 4676 5464 4684 5473
rect 4507 5456 4624 5464
rect 4676 5456 4704 5464
rect 3087 5436 3153 5444
rect 3196 5436 3233 5444
rect 2887 5396 2964 5404
rect 3056 5404 3064 5433
rect 3047 5396 3064 5404
rect 3196 5404 3204 5436
rect 3256 5436 3273 5444
rect 3256 5424 3264 5436
rect 3287 5436 3313 5444
rect 3407 5436 3493 5444
rect 3667 5436 3693 5444
rect 3747 5436 3753 5444
rect 3767 5436 3873 5444
rect 4236 5444 4244 5453
rect 4027 5436 4244 5444
rect 3227 5416 3264 5424
rect 3316 5416 3353 5424
rect 3316 5404 3324 5416
rect 3467 5416 3533 5424
rect 3667 5416 3813 5424
rect 3896 5424 3904 5433
rect 3867 5416 3904 5424
rect 3956 5424 3964 5433
rect 3927 5416 3964 5424
rect 3996 5424 4004 5433
rect 4236 5427 4244 5436
rect 4387 5436 4424 5444
rect 3996 5416 4093 5424
rect 4127 5416 4224 5424
rect 3196 5396 3324 5404
rect 3347 5396 3513 5404
rect 3527 5396 3813 5404
rect 3907 5396 4033 5404
rect 4067 5396 4113 5404
rect 4216 5404 4224 5416
rect 4327 5416 4393 5424
rect 4216 5396 4373 5404
rect 1696 5376 1853 5384
rect 1696 5364 1704 5376
rect 2527 5376 2653 5384
rect 3607 5376 3773 5384
rect 3787 5376 3973 5384
rect 4087 5376 4293 5384
rect 4416 5384 4424 5436
rect 4616 5444 4624 5456
rect 4696 5447 4704 5456
rect 4736 5456 4773 5464
rect 4736 5447 4744 5456
rect 4847 5456 4953 5464
rect 4967 5456 5173 5464
rect 5247 5456 5273 5464
rect 5307 5456 5413 5464
rect 5587 5456 5613 5464
rect 5667 5456 5744 5464
rect 4616 5436 4673 5444
rect 4787 5436 4873 5444
rect 4976 5436 5013 5444
rect 4516 5424 4524 5433
rect 4516 5416 4544 5424
rect 4467 5396 4513 5404
rect 4536 5404 4544 5416
rect 4727 5416 4813 5424
rect 4896 5416 4913 5424
rect 4896 5407 4904 5416
rect 4536 5396 4893 5404
rect 4976 5404 4984 5436
rect 5127 5436 5133 5444
rect 5147 5436 5153 5444
rect 5276 5436 5333 5444
rect 5276 5427 5284 5436
rect 5736 5444 5744 5456
rect 5767 5456 5933 5464
rect 5947 5456 5993 5464
rect 6036 5456 6093 5464
rect 5736 5436 5804 5444
rect 5007 5416 5084 5424
rect 5076 5407 5084 5416
rect 5487 5416 5533 5424
rect 5547 5416 5633 5424
rect 5796 5424 5804 5436
rect 5827 5436 5864 5444
rect 5796 5416 5833 5424
rect 5856 5424 5864 5436
rect 6036 5444 6044 5456
rect 6187 5456 6233 5464
rect 6407 5456 6473 5464
rect 6507 5456 6553 5464
rect 6587 5456 6653 5464
rect 6687 5456 6704 5464
rect 6016 5436 6044 5444
rect 5856 5416 5884 5424
rect 4927 5396 4984 5404
rect 5116 5396 5233 5404
rect 4416 5376 4433 5384
rect 4467 5376 4673 5384
rect 4687 5376 4753 5384
rect 4867 5376 4973 5384
rect 5116 5384 5124 5396
rect 5267 5396 5373 5404
rect 5387 5396 5553 5404
rect 5676 5404 5684 5413
rect 5676 5396 5773 5404
rect 4987 5376 5124 5384
rect 5587 5376 5653 5384
rect 5876 5384 5884 5416
rect 5747 5376 5884 5384
rect 5896 5384 5904 5433
rect 5916 5407 5924 5433
rect 6016 5424 6024 5436
rect 6136 5444 6144 5453
rect 6087 5436 6144 5444
rect 6256 5444 6264 5453
rect 6227 5436 6264 5444
rect 5996 5416 6024 5424
rect 5996 5387 6004 5416
rect 6056 5407 6064 5433
rect 6296 5424 6304 5453
rect 6316 5444 6324 5453
rect 6316 5436 6353 5444
rect 6456 5436 6513 5444
rect 6456 5427 6464 5436
rect 6267 5416 6313 5424
rect 6336 5416 6353 5424
rect 6147 5396 6193 5404
rect 6216 5404 6224 5413
rect 6216 5396 6233 5404
rect 6336 5404 6344 5416
rect 6587 5416 6633 5424
rect 6307 5396 6344 5404
rect 6416 5404 6424 5413
rect 6407 5396 6513 5404
rect 5896 5376 5933 5384
rect 6016 5384 6024 5393
rect 6536 5387 6544 5413
rect 6567 5396 6593 5404
rect 6607 5396 6653 5404
rect 6696 5404 6704 5456
rect 6687 5396 6704 5404
rect 6016 5376 6093 5384
rect 6016 5367 6024 5376
rect 6187 5376 6373 5384
rect 1496 5356 1704 5364
rect 2067 5356 2213 5364
rect 2367 5356 2633 5364
rect 3427 5356 4093 5364
rect 4107 5356 4293 5364
rect 4387 5356 4473 5364
rect 4527 5356 4713 5364
rect 4847 5356 5073 5364
rect 5107 5356 5333 5364
rect 5407 5356 5473 5364
rect 5507 5356 5553 5364
rect 5607 5356 5764 5364
rect 1627 5336 1813 5344
rect 1947 5336 2173 5344
rect 2227 5336 2393 5344
rect 3187 5336 3953 5344
rect 4027 5336 4193 5344
rect 4227 5336 4353 5344
rect 4507 5336 4533 5344
rect 4647 5336 4853 5344
rect 4867 5336 4913 5344
rect 5027 5336 5213 5344
rect 5227 5336 5513 5344
rect 5527 5336 5733 5344
rect 5756 5344 5764 5356
rect 5827 5356 5893 5364
rect 6567 5356 6633 5364
rect 5756 5336 5913 5344
rect 1687 5316 2193 5324
rect 3687 5316 4213 5324
rect 4287 5316 4813 5324
rect 5047 5316 5093 5324
rect 5107 5316 5433 5324
rect 5487 5316 5533 5324
rect 5767 5316 6113 5324
rect 2687 5296 2853 5304
rect 2867 5296 3033 5304
rect 3887 5296 4033 5304
rect 4047 5296 4433 5304
rect 4647 5296 4933 5304
rect 5007 5296 5793 5304
rect 5836 5296 5933 5304
rect 3107 5276 3904 5284
rect 3267 5256 3533 5264
rect 3547 5256 3613 5264
rect 3627 5256 3653 5264
rect 3896 5264 3904 5276
rect 4367 5276 4473 5284
rect 4496 5276 4553 5284
rect 3896 5256 4013 5264
rect 4127 5256 4153 5264
rect 4496 5264 4504 5276
rect 4687 5276 5013 5284
rect 5047 5276 5113 5284
rect 5127 5276 5253 5284
rect 5347 5276 5813 5284
rect 4207 5256 4504 5264
rect 4527 5256 4573 5264
rect 4587 5256 4733 5264
rect 4907 5256 5053 5264
rect 5087 5256 5153 5264
rect 5247 5256 5313 5264
rect 5387 5256 5513 5264
rect 5836 5264 5844 5296
rect 5967 5296 6033 5304
rect 6087 5296 6113 5304
rect 5867 5276 6313 5284
rect 5547 5256 5844 5264
rect 5907 5256 6093 5264
rect 2627 5236 2733 5244
rect 3527 5236 3633 5244
rect 4027 5236 4413 5244
rect 4427 5236 4593 5244
rect 4607 5236 4793 5244
rect 4807 5236 5033 5244
rect 5047 5236 5173 5244
rect 5187 5236 5353 5244
rect 5367 5236 5573 5244
rect 5587 5236 5873 5244
rect 5887 5236 5893 5244
rect 5947 5236 5973 5244
rect 6007 5236 6064 5244
rect 527 5216 573 5224
rect 587 5216 933 5224
rect 2707 5216 2793 5224
rect 3187 5216 3653 5224
rect 3967 5216 4173 5224
rect 387 5196 593 5204
rect 827 5196 873 5204
rect 1527 5196 1564 5204
rect -24 5144 -16 5164
rect 127 5156 313 5164
rect 336 5147 344 5193
rect 376 5176 493 5184
rect 376 5164 384 5176
rect 507 5176 533 5184
rect 807 5176 833 5184
rect 1087 5176 1153 5184
rect 367 5156 384 5164
rect 427 5156 453 5164
rect 567 5156 613 5164
rect 867 5156 933 5164
rect 987 5156 1024 5164
rect 1016 5147 1024 5156
rect 1087 5156 1113 5164
rect -24 5136 33 5144
rect 87 5136 113 5144
rect 456 5136 664 5144
rect 207 5116 353 5124
rect 456 5124 464 5136
rect 367 5116 464 5124
rect 487 5116 513 5124
rect 656 5124 664 5136
rect 687 5136 953 5144
rect 1136 5144 1144 5176
rect 1387 5176 1404 5184
rect 1396 5164 1404 5176
rect 1247 5156 1384 5164
rect 1396 5156 1493 5164
rect 1107 5136 1144 5144
rect 1376 5144 1384 5156
rect 1536 5164 1544 5173
rect 1556 5167 1564 5196
rect 2267 5196 2293 5204
rect 2307 5196 2373 5204
rect 2387 5196 2753 5204
rect 2927 5196 3133 5204
rect 3367 5196 3453 5204
rect 3467 5196 3693 5204
rect 1907 5176 2013 5184
rect 2047 5176 2073 5184
rect 2187 5176 2224 5184
rect 1516 5156 1544 5164
rect 1516 5144 1524 5156
rect 1956 5156 1993 5164
rect 1376 5136 1524 5144
rect 1647 5136 1673 5144
rect 1767 5136 1913 5144
rect 656 5116 713 5124
rect 727 5116 733 5124
rect 1007 5116 1053 5124
rect 1236 5107 1244 5133
rect 1936 5127 1944 5153
rect 1956 5147 1964 5156
rect 2027 5136 2053 5144
rect 2136 5144 2144 5173
rect 2167 5156 2193 5164
rect 2216 5164 2224 5176
rect 2247 5176 2413 5184
rect 2507 5176 2593 5184
rect 2687 5176 2744 5184
rect 2216 5156 2233 5164
rect 2407 5156 2453 5164
rect 2507 5156 2564 5164
rect 2556 5147 2564 5156
rect 2736 5147 2744 5176
rect 3127 5176 3173 5184
rect 3227 5176 3233 5184
rect 3247 5176 3273 5184
rect 3296 5176 3373 5184
rect 2876 5164 2884 5173
rect 2876 5156 2933 5164
rect 2956 5164 2964 5173
rect 2956 5156 3013 5164
rect 2127 5136 2353 5144
rect 2447 5136 2493 5144
rect 2756 5127 2764 5153
rect 2847 5136 2993 5144
rect 3096 5144 3104 5173
rect 3296 5167 3304 5176
rect 3716 5176 3744 5184
rect 3147 5156 3193 5164
rect 3347 5156 3493 5164
rect 3536 5147 3544 5173
rect 3096 5136 3113 5144
rect 3176 5136 3433 5144
rect 1327 5116 1713 5124
rect 1727 5116 1753 5124
rect 2127 5116 2573 5124
rect 2587 5116 2613 5124
rect 2787 5116 2793 5124
rect 2807 5116 2853 5124
rect 3007 5116 3013 5124
rect 3176 5124 3184 5136
rect 3456 5136 3504 5144
rect 3456 5127 3464 5136
rect 3027 5116 3184 5124
rect 3367 5116 3393 5124
rect 3416 5116 3453 5124
rect 247 5096 433 5104
rect 1027 5096 1133 5104
rect 2007 5096 2533 5104
rect 2747 5096 2833 5104
rect 2987 5096 3213 5104
rect 3416 5104 3424 5116
rect 3496 5124 3504 5136
rect 3556 5144 3564 5153
rect 3556 5136 3573 5144
rect 3596 5124 3604 5173
rect 3636 5144 3644 5173
rect 3716 5164 3724 5176
rect 3667 5156 3724 5164
rect 3736 5147 3744 5176
rect 3947 5176 3973 5184
rect 4067 5176 4084 5184
rect 3827 5156 3893 5164
rect 3636 5136 3713 5144
rect 3756 5144 3764 5153
rect 4016 5147 4024 5173
rect 4036 5147 4044 5173
rect 3756 5136 3833 5144
rect 3847 5136 3993 5144
rect 3496 5116 3604 5124
rect 3707 5116 3813 5124
rect 4056 5124 4064 5153
rect 4076 5147 4084 5176
rect 4096 5167 4104 5216
rect 4196 5216 4273 5224
rect 4156 5147 4164 5173
rect 4196 5164 4204 5216
rect 4327 5216 4373 5224
rect 4467 5216 4613 5224
rect 4627 5216 5044 5224
rect 4227 5196 4933 5204
rect 5036 5204 5044 5216
rect 5127 5216 5444 5224
rect 5036 5196 5093 5204
rect 4267 5176 4333 5184
rect 4447 5176 4544 5184
rect 4187 5156 4204 5164
rect 4236 5144 4244 5173
rect 4256 5147 4264 5173
rect 4367 5156 4393 5164
rect 4416 5156 4453 5164
rect 4187 5136 4244 5144
rect 4416 5144 4424 5156
rect 4476 5156 4513 5164
rect 4347 5136 4424 5144
rect 4476 5144 4484 5156
rect 4536 5164 4544 5176
rect 4567 5176 4584 5184
rect 4576 5164 4584 5176
rect 4536 5156 4564 5164
rect 4576 5156 4613 5164
rect 4447 5136 4484 5144
rect 4507 5136 4533 5144
rect 4556 5144 4564 5156
rect 4556 5136 4593 5144
rect 4636 5144 4644 5173
rect 4707 5156 4733 5164
rect 4787 5156 4873 5164
rect 4627 5136 4644 5144
rect 4667 5136 4693 5144
rect 4887 5136 4913 5144
rect 4056 5116 4093 5124
rect 4107 5116 4213 5124
rect 4287 5116 4413 5124
rect 4447 5116 4473 5124
rect 4667 5116 4773 5124
rect 5016 5124 5024 5193
rect 5036 5147 5044 5196
rect 5207 5196 5253 5204
rect 5287 5196 5373 5204
rect 5436 5187 5444 5216
rect 5527 5216 5753 5224
rect 6056 5224 6064 5236
rect 6387 5236 6433 5244
rect 5847 5216 5984 5224
rect 6056 5216 6193 5224
rect 5627 5196 5724 5204
rect 5076 5176 5113 5184
rect 5076 5144 5084 5176
rect 5136 5176 5233 5184
rect 5136 5164 5144 5176
rect 5347 5176 5424 5184
rect 5107 5156 5144 5164
rect 5156 5156 5193 5164
rect 5076 5136 5093 5144
rect 5156 5144 5164 5156
rect 5236 5156 5333 5164
rect 5236 5144 5244 5156
rect 5416 5164 5424 5176
rect 5487 5176 5533 5184
rect 5647 5176 5693 5184
rect 5416 5156 5464 5164
rect 5376 5144 5384 5153
rect 5127 5136 5164 5144
rect 5216 5136 5244 5144
rect 5336 5136 5384 5144
rect 5456 5144 5464 5156
rect 5527 5156 5693 5164
rect 5456 5136 5473 5144
rect 5216 5124 5224 5136
rect 5016 5116 5044 5124
rect 3227 5096 3424 5104
rect 3447 5096 3773 5104
rect 3967 5096 4233 5104
rect 4307 5096 4313 5104
rect 4327 5096 4813 5104
rect 4827 5096 4833 5104
rect 5036 5104 5044 5116
rect 5196 5116 5224 5124
rect 5036 5096 5073 5104
rect 1047 5076 1113 5084
rect 1127 5076 1193 5084
rect 2467 5076 2813 5084
rect 2827 5076 3053 5084
rect 3327 5076 3373 5084
rect 3387 5076 3473 5084
rect 3807 5076 3853 5084
rect 3867 5076 4273 5084
rect 4307 5076 4333 5084
rect 5196 5084 5204 5116
rect 5336 5124 5344 5136
rect 5507 5136 5573 5144
rect 5596 5136 5673 5144
rect 5247 5116 5344 5124
rect 5596 5124 5604 5136
rect 5716 5144 5724 5196
rect 5747 5196 5873 5204
rect 5976 5187 5984 5216
rect 6287 5216 6353 5224
rect 6427 5216 6513 5224
rect 6187 5196 6253 5204
rect 6407 5196 6464 5204
rect 5747 5176 5773 5184
rect 5787 5176 5844 5184
rect 5836 5167 5844 5176
rect 5996 5184 6004 5193
rect 6456 5187 6464 5196
rect 6507 5196 6553 5204
rect 6607 5196 6624 5204
rect 6616 5187 6624 5196
rect 6687 5196 6704 5204
rect 5996 5176 6024 5184
rect 5927 5156 5993 5164
rect 6016 5147 6024 5176
rect 6156 5176 6233 5184
rect 6056 5147 6064 5173
rect 6156 5164 6164 5176
rect 6367 5176 6393 5184
rect 6536 5176 6573 5184
rect 6087 5156 6164 5164
rect 6196 5156 6333 5164
rect 5716 5136 5784 5144
rect 5367 5116 5604 5124
rect 5647 5116 5693 5124
rect 5776 5124 5784 5136
rect 5867 5136 5873 5144
rect 5887 5136 5953 5144
rect 6196 5127 6204 5156
rect 6347 5156 6433 5164
rect 6487 5156 6513 5164
rect 6247 5136 6313 5144
rect 6327 5136 6373 5144
rect 6536 5144 6544 5176
rect 6567 5156 6613 5164
rect 6656 5164 6664 5173
rect 6647 5156 6664 5164
rect 6696 5164 6704 5196
rect 6696 5156 6744 5164
rect 6447 5136 6524 5144
rect 6536 5136 6553 5144
rect 5776 5116 5913 5124
rect 5947 5116 6113 5124
rect 6287 5116 6353 5124
rect 6387 5116 6493 5124
rect 6516 5124 6524 5136
rect 6667 5136 6713 5144
rect 6516 5116 6673 5124
rect 6736 5124 6744 5156
rect 6707 5116 6744 5124
rect 5287 5096 5553 5104
rect 5627 5096 5693 5104
rect 5707 5096 5773 5104
rect 5827 5096 6133 5104
rect 6167 5096 6233 5104
rect 6547 5096 6593 5104
rect 4487 5076 5204 5084
rect 5287 5076 5733 5084
rect 5747 5076 5753 5084
rect 5847 5076 5893 5084
rect 5987 5076 6053 5084
rect 6087 5076 6113 5084
rect 2767 5056 2853 5064
rect 2867 5056 2893 5064
rect 2907 5056 2953 5064
rect 2976 5056 3313 5064
rect 1067 5036 1133 5044
rect 1147 5036 1393 5044
rect 2147 5036 2213 5044
rect 2976 5044 2984 5056
rect 3347 5056 3553 5064
rect 3827 5056 3893 5064
rect 4007 5056 4033 5064
rect 4047 5056 6133 5064
rect 2227 5036 2984 5044
rect 3007 5036 3093 5044
rect 3107 5036 3113 5044
rect 3127 5036 3273 5044
rect 3447 5036 3653 5044
rect 3667 5036 4093 5044
rect 4107 5036 4333 5044
rect 4367 5036 4873 5044
rect 4907 5036 5113 5044
rect 5156 5036 5833 5044
rect 87 5016 893 5024
rect 1207 5016 1253 5024
rect 2047 5016 2333 5024
rect 2687 5016 2953 5024
rect 3207 5016 3933 5024
rect 3947 5016 4253 5024
rect 4287 5016 4404 5024
rect 567 4996 613 5004
rect 647 4996 733 5004
rect 987 4996 1173 5004
rect 1227 4996 1353 5004
rect 1587 4996 1613 5004
rect 1967 4996 2033 5004
rect 2227 4996 2233 5004
rect 2247 4996 2373 5004
rect 2396 4996 2593 5004
rect 576 4976 724 4984
rect -24 4956 33 4964
rect 56 4956 113 4964
rect 56 4944 64 4956
rect 167 4956 273 4964
rect 407 4956 513 4964
rect 576 4964 584 4976
rect 536 4956 584 4964
rect 536 4947 544 4956
rect 627 4956 664 4964
rect -24 4936 64 4944
rect -24 4916 -16 4936
rect 227 4936 504 4944
rect 247 4916 273 4924
rect 496 4924 504 4936
rect 616 4944 624 4953
rect 567 4936 624 4944
rect 656 4927 664 4956
rect 676 4956 693 4964
rect 676 4927 684 4956
rect 716 4964 724 4976
rect 827 4976 1093 4984
rect 1367 4976 1493 4984
rect 1507 4976 1593 4984
rect 1607 4976 1653 4984
rect 1667 4976 1673 4984
rect 1687 4976 1933 4984
rect 2167 4976 2273 4984
rect 2396 4984 2404 4996
rect 2807 4996 2924 5004
rect 2367 4976 2404 4984
rect 2427 4976 2624 4984
rect 716 4956 833 4964
rect 1167 4956 1204 4964
rect 1196 4947 1204 4956
rect 1216 4956 1313 4964
rect 707 4936 733 4944
rect 767 4936 793 4944
rect 816 4936 853 4944
rect 816 4927 824 4936
rect 867 4936 893 4944
rect 967 4936 1184 4944
rect 1176 4927 1184 4936
rect 496 4916 573 4924
rect 587 4916 613 4924
rect 727 4916 804 4924
rect 207 4896 593 4904
rect 607 4896 773 4904
rect 796 4904 804 4916
rect 847 4916 1153 4924
rect 1216 4924 1224 4956
rect 1847 4956 1933 4964
rect 1307 4936 1324 4944
rect 1187 4916 1224 4924
rect 1247 4916 1273 4924
rect 1316 4924 1324 4936
rect 1347 4936 1433 4944
rect 1547 4936 1593 4944
rect 1616 4927 1624 4953
rect 1727 4936 1773 4944
rect 1796 4927 1804 4953
rect 1827 4936 1873 4944
rect 1927 4936 1953 4944
rect 1976 4927 1984 4973
rect 1996 4947 2004 4973
rect 2027 4956 2073 4964
rect 2207 4956 2284 4964
rect 2107 4936 2133 4944
rect 2276 4944 2284 4956
rect 2616 4964 2624 4976
rect 2647 4976 2764 4984
rect 2616 4956 2693 4964
rect 2756 4964 2764 4976
rect 2827 4976 2893 4984
rect 2916 4984 2924 4996
rect 2947 4996 3004 5004
rect 2916 4976 2933 4984
rect 2996 4984 3004 4996
rect 3047 4996 3833 5004
rect 3927 4996 4044 5004
rect 2996 4976 3153 4984
rect 3187 4976 3413 4984
rect 3427 4976 3753 4984
rect 3847 4976 3933 4984
rect 3947 4976 3993 4984
rect 4036 4984 4044 4996
rect 4087 4996 4113 5004
rect 4227 4996 4353 5004
rect 4396 5004 4404 5016
rect 5156 5024 5164 5036
rect 6027 5036 6113 5044
rect 6287 5036 6333 5044
rect 4427 5016 5164 5024
rect 5187 5016 5373 5024
rect 5427 5016 5553 5024
rect 5587 5016 5853 5024
rect 5887 5016 6073 5024
rect 6107 5016 6213 5024
rect 6227 5016 6393 5024
rect 4396 4996 4513 5004
rect 4576 4996 4613 5004
rect 4036 4976 4064 4984
rect 2756 4956 2813 4964
rect 2276 4936 2413 4944
rect 2436 4944 2444 4953
rect 2976 4947 2984 4973
rect 3027 4956 3053 4964
rect 3147 4956 3253 4964
rect 3287 4956 3493 4964
rect 3567 4956 3593 4964
rect 3616 4956 3713 4964
rect 2436 4936 2673 4944
rect 2727 4936 2753 4944
rect 2787 4936 2833 4944
rect 2887 4936 2913 4944
rect 3087 4936 3113 4944
rect 3136 4936 3293 4944
rect 1316 4916 1344 4924
rect 796 4896 833 4904
rect 1227 4896 1313 4904
rect 627 4876 693 4884
rect 767 4876 1233 4884
rect 1336 4884 1344 4916
rect 1907 4916 1944 4924
rect 1427 4896 1593 4904
rect 1747 4896 1913 4904
rect 1936 4904 1944 4916
rect 2267 4916 2293 4924
rect 2627 4916 2773 4924
rect 3136 4924 3144 4936
rect 3307 4936 3353 4944
rect 3407 4936 3433 4944
rect 3616 4944 3624 4956
rect 3816 4956 3913 4964
rect 3816 4947 3824 4956
rect 4016 4964 4024 4973
rect 4056 4964 4064 4976
rect 4167 4976 4193 4984
rect 4576 4984 4584 4996
rect 4627 4996 4893 5004
rect 4947 4996 5013 5004
rect 5036 4996 5093 5004
rect 4207 4976 4584 4984
rect 3967 4956 3984 4964
rect 4016 4956 4044 4964
rect 3547 4936 3624 4944
rect 3667 4936 3693 4944
rect 3867 4936 3953 4944
rect 2907 4916 3144 4924
rect 3187 4916 3193 4924
rect 3207 4916 3233 4924
rect 3247 4916 3273 4924
rect 3347 4916 3653 4924
rect 3736 4924 3744 4933
rect 3727 4916 3744 4924
rect 3827 4916 3893 4924
rect 3976 4924 3984 4956
rect 4036 4947 4044 4956
rect 4056 4956 4184 4964
rect 4056 4947 4064 4956
rect 4176 4944 4184 4956
rect 4176 4936 4233 4944
rect 3976 4916 3993 4924
rect 4076 4924 4084 4933
rect 4256 4927 4264 4953
rect 4296 4944 4304 4953
rect 4296 4936 4324 4944
rect 4067 4916 4084 4924
rect 4127 4916 4173 4924
rect 4187 4916 4193 4924
rect 1936 4896 2493 4904
rect 2927 4896 3013 4904
rect 3647 4896 4113 4904
rect 4147 4896 4213 4904
rect 4276 4904 4284 4933
rect 4316 4927 4324 4936
rect 4356 4927 4364 4976
rect 4727 4976 4753 4984
rect 5036 4984 5044 4996
rect 5207 4996 5393 5004
rect 5407 4996 5713 5004
rect 5867 4996 5913 5004
rect 5927 4996 6193 5004
rect 6287 4996 6433 5004
rect 6507 4996 6553 5004
rect 6607 4996 6653 5004
rect 4807 4976 5044 4984
rect 4387 4956 4424 4964
rect 4416 4944 4424 4956
rect 4447 4956 4464 4964
rect 4407 4936 4433 4944
rect 4456 4944 4464 4956
rect 4507 4956 4593 4964
rect 4676 4956 4813 4964
rect 4456 4936 4473 4944
rect 4496 4927 4504 4953
rect 4567 4936 4593 4944
rect 4267 4896 4284 4904
rect 4616 4904 4624 4953
rect 4676 4947 4684 4956
rect 4776 4927 4784 4956
rect 4907 4956 4973 4964
rect 4836 4944 4844 4953
rect 4816 4936 4844 4944
rect 4816 4927 4824 4936
rect 4747 4916 4764 4924
rect 4367 4896 4713 4904
rect 4756 4887 4764 4916
rect 4876 4924 4884 4953
rect 4876 4916 4973 4924
rect 4996 4907 5004 4976
rect 5067 4976 5133 4984
rect 5147 4976 5173 4984
rect 5227 4976 5333 4984
rect 5376 4976 5453 4984
rect 5027 4956 5064 4964
rect 5056 4927 5064 4956
rect 5216 4956 5253 4964
rect 5096 4927 5104 4953
rect 5216 4927 5224 4956
rect 5267 4956 5273 4964
rect 5327 4956 5353 4964
rect 5376 4944 5384 4976
rect 5567 4976 5593 4984
rect 5667 4976 5713 4984
rect 5807 4976 5873 4984
rect 5927 4976 6033 4984
rect 6247 4976 6293 4984
rect 6587 4976 6613 4984
rect 5476 4964 5484 4973
rect 5407 4956 5484 4964
rect 5496 4956 5533 4964
rect 5376 4936 5413 4944
rect 5496 4944 5504 4956
rect 5616 4956 5633 4964
rect 5447 4936 5504 4944
rect 5147 4916 5173 4924
rect 5267 4916 5353 4924
rect 5576 4924 5584 4953
rect 5616 4924 5624 4956
rect 5767 4956 5804 4964
rect 5796 4947 5804 4956
rect 5816 4956 5973 4964
rect 5816 4947 5824 4956
rect 6016 4956 6053 4964
rect 5647 4936 5684 4944
rect 5527 4916 5584 4924
rect 5596 4916 5624 4924
rect 4847 4896 4993 4904
rect 5047 4896 5093 4904
rect 5127 4896 5273 4904
rect 5287 4896 5493 4904
rect 5507 4896 5573 4904
rect 1287 4876 1344 4884
rect 1467 4876 1553 4884
rect 1567 4876 1953 4884
rect 2547 4876 3853 4884
rect 3867 4876 4413 4884
rect 4647 4876 4733 4884
rect 4927 4876 4953 4884
rect 4987 4876 5033 4884
rect 5067 4876 5224 4884
rect 647 4856 753 4864
rect 767 4856 1673 4864
rect 1687 4856 1973 4864
rect 3667 4856 3973 4864
rect 4087 4856 4473 4864
rect 4587 4856 5153 4864
rect 5216 4864 5224 4876
rect 5247 4876 5413 4884
rect 5596 4884 5604 4916
rect 5676 4924 5684 4936
rect 5927 4936 5973 4944
rect 5676 4916 5753 4924
rect 5627 4896 5633 4904
rect 5656 4904 5664 4913
rect 5876 4907 5884 4933
rect 5996 4927 6004 4953
rect 6016 4927 6024 4956
rect 6096 4956 6113 4964
rect 6096 4944 6104 4956
rect 6167 4956 6293 4964
rect 6327 4956 6413 4964
rect 6487 4956 6513 4964
rect 6536 4956 6553 4964
rect 6056 4936 6104 4944
rect 6056 4927 6064 4936
rect 6127 4936 6173 4944
rect 6207 4936 6253 4944
rect 6387 4936 6473 4944
rect 6536 4944 6544 4956
rect 6487 4936 6544 4944
rect 6087 4916 6193 4924
rect 6207 4916 6353 4924
rect 6476 4916 6493 4924
rect 5656 4896 5773 4904
rect 5827 4896 5833 4904
rect 5967 4896 6033 4904
rect 6047 4896 6333 4904
rect 6396 4904 6404 4913
rect 6476 4904 6484 4916
rect 6547 4916 6633 4924
rect 6396 4896 6484 4904
rect 5587 4876 5604 4884
rect 5627 4876 5713 4884
rect 5767 4876 6033 4884
rect 6147 4876 6273 4884
rect 5216 4856 5273 4864
rect 5307 4856 5453 4864
rect 5607 4856 5853 4864
rect 5887 4856 6453 4864
rect 1907 4836 1993 4844
rect 2507 4836 3813 4844
rect 3867 4836 4313 4844
rect 4347 4836 4653 4844
rect 4727 4836 4833 4844
rect 4856 4836 5113 4844
rect 1947 4816 3833 4824
rect 4267 4816 4633 4824
rect 4856 4824 4864 4836
rect 5207 4836 5433 4844
rect 5567 4836 5753 4844
rect 5787 4836 5913 4844
rect 5947 4836 6633 4844
rect 4707 4816 4864 4824
rect 4887 4816 5013 4824
rect 5056 4816 5073 4824
rect 1007 4796 1253 4804
rect 1827 4796 1853 4804
rect 3747 4796 3833 4804
rect 3887 4796 3933 4804
rect 4007 4796 4353 4804
rect 4407 4796 4753 4804
rect 5056 4804 5064 4816
rect 5087 4816 5373 4824
rect 5387 4816 5473 4824
rect 5487 4816 5813 4824
rect 5867 4816 6013 4824
rect 4847 4796 5064 4804
rect 5107 4796 5293 4804
rect 5427 4796 5713 4804
rect 5807 4796 6153 4804
rect 6307 4796 6473 4804
rect 307 4776 413 4784
rect 1347 4776 1393 4784
rect 3587 4776 3993 4784
rect 4107 4776 5593 4784
rect 5707 4776 5953 4784
rect 6007 4776 6173 4784
rect 6187 4776 6493 4784
rect 1367 4756 1413 4764
rect 1627 4756 2093 4764
rect 3767 4756 3853 4764
rect 4207 4756 4273 4764
rect 4607 4756 4673 4764
rect 4967 4756 4993 4764
rect 5107 4756 5193 4764
rect 5227 4756 5253 4764
rect 5287 4756 5573 4764
rect 5667 4756 5733 4764
rect 5767 4756 6013 4764
rect 6307 4756 6353 4764
rect 747 4736 1553 4744
rect 1567 4736 1693 4744
rect 2247 4736 2433 4744
rect 4167 4736 4293 4744
rect 4387 4736 4613 4744
rect 4827 4736 4973 4744
rect 5007 4736 5053 4744
rect 5076 4736 5424 4744
rect 1307 4716 1344 4724
rect 187 4696 544 4704
rect 236 4676 313 4684
rect 236 4667 244 4676
rect 447 4676 513 4684
rect 536 4684 544 4696
rect 847 4696 913 4704
rect 927 4696 933 4704
rect 1247 4696 1324 4704
rect 1316 4687 1324 4696
rect 536 4676 813 4684
rect 907 4676 1193 4684
rect 1287 4676 1304 4684
rect 336 4647 344 4673
rect 367 4656 373 4664
rect 396 4664 404 4673
rect 396 4656 533 4664
rect 547 4656 613 4664
rect 847 4656 893 4664
rect 1087 4656 1213 4664
rect 1296 4664 1304 4676
rect 1336 4684 1344 4716
rect 1587 4716 1733 4724
rect 1856 4716 1933 4724
rect 1856 4704 1864 4716
rect 2176 4716 2393 4724
rect 2176 4704 2184 4716
rect 2407 4716 2413 4724
rect 2427 4716 2513 4724
rect 3007 4716 4473 4724
rect 4507 4716 4653 4724
rect 4687 4716 4784 4724
rect 1647 4696 1864 4704
rect 1876 4696 2184 4704
rect 1336 4676 1373 4684
rect 1447 4676 1484 4684
rect 1476 4667 1484 4676
rect 1507 4676 1544 4684
rect 1536 4667 1544 4676
rect 1567 4676 1624 4684
rect 1616 4667 1624 4676
rect 1727 4676 1764 4684
rect 1296 4656 1353 4664
rect 1407 4656 1453 4664
rect 1547 4656 1584 4664
rect 347 4636 373 4644
rect 507 4636 513 4644
rect 527 4636 553 4644
rect 667 4636 793 4644
rect 827 4636 1033 4644
rect 1447 4636 1553 4644
rect 1576 4644 1584 4656
rect 1696 4647 1704 4673
rect 1756 4667 1764 4676
rect 1827 4676 1853 4684
rect 1876 4667 1884 4696
rect 2207 4696 2253 4704
rect 2276 4696 2353 4704
rect 1947 4676 2213 4684
rect 1767 4656 1833 4664
rect 2276 4664 2284 4696
rect 2376 4696 2433 4704
rect 2376 4687 2384 4696
rect 3287 4696 3313 4704
rect 3327 4696 3633 4704
rect 3647 4696 3773 4704
rect 4127 4696 4153 4704
rect 4247 4696 4273 4704
rect 4467 4696 4513 4704
rect 4776 4704 4784 4716
rect 4807 4716 4873 4724
rect 5076 4724 5084 4736
rect 4927 4716 5084 4724
rect 5187 4716 5253 4724
rect 5267 4716 5293 4724
rect 5347 4716 5393 4724
rect 5416 4724 5424 4736
rect 5487 4736 5564 4744
rect 5416 4716 5513 4724
rect 5556 4724 5564 4736
rect 5727 4736 6093 4744
rect 6167 4736 6293 4744
rect 6347 4736 6513 4744
rect 6567 4736 6613 4744
rect 5556 4716 5633 4724
rect 5556 4707 5564 4716
rect 5787 4716 6153 4724
rect 6167 4716 6193 4724
rect 6207 4716 6253 4724
rect 6427 4716 6433 4724
rect 6447 4716 6653 4724
rect 6667 4716 6673 4724
rect 4707 4696 4744 4704
rect 4776 4696 4913 4704
rect 2307 4676 2344 4684
rect 2276 4656 2313 4664
rect 2336 4664 2344 4676
rect 2396 4676 2504 4684
rect 2396 4664 2404 4676
rect 2336 4656 2404 4664
rect 2496 4664 2504 4676
rect 2607 4676 2633 4684
rect 2647 4676 2893 4684
rect 3507 4676 3553 4684
rect 3707 4676 3753 4684
rect 3807 4676 3853 4684
rect 4196 4684 4204 4693
rect 4147 4676 4673 4684
rect 2496 4656 2564 4664
rect 1576 4636 1633 4644
rect 1807 4636 1813 4644
rect 1827 4636 2293 4644
rect 2347 4636 2373 4644
rect 2467 4636 2533 4644
rect 2556 4644 2564 4656
rect 2587 4656 2684 4664
rect 2556 4636 2593 4644
rect 2676 4644 2684 4656
rect 2827 4656 2953 4664
rect 3107 4656 3153 4664
rect 3407 4656 3533 4664
rect 3556 4664 3564 4673
rect 3556 4656 3613 4664
rect 3667 4656 3753 4664
rect 4247 4656 4293 4664
rect 4427 4656 4533 4664
rect 4596 4656 4633 4664
rect 2676 4636 2793 4644
rect 3127 4636 3353 4644
rect 3587 4636 3733 4644
rect 4067 4636 4173 4644
rect 4507 4636 4573 4644
rect 287 4616 353 4624
rect 576 4624 584 4633
rect 576 4616 713 4624
rect 827 4616 853 4624
rect 867 4616 1273 4624
rect 1527 4616 1573 4624
rect 1587 4616 1773 4624
rect 2327 4616 2453 4624
rect 3787 4616 3913 4624
rect 4596 4624 4604 4656
rect 4696 4647 4704 4673
rect 4716 4644 4724 4673
rect 4736 4667 4744 4696
rect 4987 4696 5033 4704
rect 5067 4696 5093 4704
rect 5147 4696 5153 4704
rect 5207 4696 5224 4704
rect 4956 4684 4964 4693
rect 4867 4676 4964 4684
rect 5067 4676 5113 4684
rect 4716 4636 4733 4644
rect 4756 4627 4764 4673
rect 4807 4656 4833 4664
rect 4887 4656 4933 4664
rect 5007 4656 5073 4664
rect 5136 4664 5144 4693
rect 5216 4687 5224 4696
rect 5247 4696 5324 4704
rect 5247 4676 5293 4684
rect 5316 4684 5324 4696
rect 5527 4696 5544 4704
rect 5316 4676 5393 4684
rect 5416 4684 5424 4693
rect 5416 4676 5464 4684
rect 5087 4656 5144 4664
rect 5287 4656 5373 4664
rect 5407 4656 5433 4664
rect 5456 4664 5464 4676
rect 5456 4656 5473 4664
rect 5536 4664 5544 4696
rect 5576 4696 5593 4704
rect 5576 4684 5584 4696
rect 5567 4676 5584 4684
rect 5536 4656 5593 4664
rect 5676 4664 5684 4713
rect 5747 4696 5833 4704
rect 5947 4696 5973 4704
rect 6196 4696 6233 4704
rect 5696 4684 5704 4693
rect 5696 4676 5733 4684
rect 5927 4676 5953 4684
rect 5616 4656 5684 4664
rect 4807 4636 5153 4644
rect 5167 4636 5233 4644
rect 5347 4636 5433 4644
rect 5616 4644 5624 4656
rect 5727 4656 5773 4664
rect 5856 4664 5864 4673
rect 6056 4667 6064 4693
rect 6196 4684 6204 4696
rect 6356 4704 6364 4713
rect 6356 4696 6373 4704
rect 6456 4696 6473 4704
rect 6096 4676 6204 4684
rect 5856 4656 5913 4664
rect 5987 4656 6044 4664
rect 5547 4636 5624 4644
rect 5647 4636 5713 4644
rect 6036 4644 6044 4656
rect 6096 4644 6104 4676
rect 6227 4676 6273 4684
rect 6316 4684 6324 4693
rect 6316 4676 6344 4684
rect 6127 4656 6304 4664
rect 6036 4636 6273 4644
rect 6296 4644 6304 4656
rect 6336 4644 6344 4676
rect 6407 4656 6433 4664
rect 6296 4636 6344 4644
rect 6456 4644 6464 4696
rect 6507 4696 6573 4704
rect 6516 4656 6553 4664
rect 6516 4647 6524 4656
rect 6447 4636 6464 4644
rect 4007 4616 4604 4624
rect 4627 4616 4673 4624
rect 4687 4616 4713 4624
rect 5207 4616 5344 4624
rect 307 4596 333 4604
rect 376 4596 953 4604
rect 376 4584 384 4596
rect 1667 4596 2653 4604
rect 3087 4596 4093 4604
rect 4187 4596 4273 4604
rect 4327 4596 4353 4604
rect 4467 4596 4773 4604
rect 4847 4596 5033 4604
rect 5047 4596 5273 4604
rect 5336 4604 5344 4616
rect 5367 4616 5433 4624
rect 5447 4616 5453 4624
rect 5476 4616 5653 4624
rect 5476 4604 5484 4616
rect 5707 4616 5733 4624
rect 6147 4616 6373 4624
rect 6467 4616 6613 4624
rect 5336 4596 5484 4604
rect 5507 4596 5853 4604
rect 6247 4596 6333 4604
rect 6387 4596 6473 4604
rect 267 4576 384 4584
rect 407 4576 773 4584
rect 1127 4576 1153 4584
rect 1367 4576 2293 4584
rect 2307 4576 2353 4584
rect 2387 4576 2433 4584
rect 4567 4576 4853 4584
rect 5047 4576 5413 4584
rect 5567 4576 5664 4584
rect 147 4556 453 4564
rect 1387 4556 1873 4564
rect 3827 4556 3933 4564
rect 3947 4556 4373 4564
rect 4607 4556 5053 4564
rect 5107 4556 5573 4564
rect 5656 4564 5664 4576
rect 5687 4576 5753 4584
rect 5807 4576 6213 4584
rect 6287 4576 6353 4584
rect 5656 4556 5893 4564
rect 6027 4556 6073 4564
rect 6487 4556 6553 4564
rect 347 4536 413 4544
rect 447 4536 493 4544
rect 747 4536 913 4544
rect 2987 4536 3644 4544
rect 87 4516 213 4524
rect 427 4516 733 4524
rect 807 4516 973 4524
rect 1247 4516 1653 4524
rect 1667 4516 1833 4524
rect 2067 4516 2193 4524
rect 2407 4516 2513 4524
rect 2527 4516 2573 4524
rect 3387 4516 3453 4524
rect 3636 4524 3644 4536
rect 3867 4536 4693 4544
rect 4767 4536 4853 4544
rect 4907 4536 5153 4544
rect 5347 4536 5393 4544
rect 5467 4536 5493 4544
rect 5507 4536 5673 4544
rect 5947 4536 6253 4544
rect 6327 4536 6613 4544
rect 3636 4516 3933 4524
rect 4076 4516 4133 4524
rect 67 4496 113 4504
rect 207 4496 353 4504
rect 527 4496 613 4504
rect 907 4496 924 4504
rect 196 4476 273 4484
rect -24 4444 -16 4464
rect 47 4456 73 4464
rect 96 4464 104 4473
rect 196 4467 204 4476
rect 327 4476 344 4484
rect 96 4456 153 4464
rect 167 4456 173 4464
rect 247 4456 313 4464
rect 336 4464 344 4476
rect 336 4456 353 4464
rect 376 4464 384 4493
rect 467 4476 513 4484
rect 696 4476 753 4484
rect 376 4456 413 4464
rect 436 4464 444 4473
rect 436 4456 593 4464
rect 696 4464 704 4476
rect 836 4484 844 4493
rect 767 4476 844 4484
rect 627 4456 704 4464
rect 896 4464 904 4473
rect 916 4467 924 4496
rect 1067 4496 1233 4504
rect 1367 4496 1413 4504
rect 1507 4496 1613 4504
rect 1747 4496 1853 4504
rect 1867 4496 2033 4504
rect 2047 4496 2153 4504
rect 2167 4496 2173 4504
rect 2727 4496 2853 4504
rect 3407 4496 3493 4504
rect 3507 4496 3573 4504
rect 1287 4476 1373 4484
rect 1407 4476 1453 4484
rect 1907 4476 1933 4484
rect 1967 4476 2073 4484
rect 3307 4476 3433 4484
rect 3547 4476 3673 4484
rect 867 4456 904 4464
rect 936 4464 944 4473
rect 936 4456 993 4464
rect 1516 4456 1553 4464
rect 1516 4447 1524 4456
rect 2436 4464 2444 4473
rect 2327 4456 2444 4464
rect 2507 4456 2533 4464
rect 2816 4464 2824 4473
rect 2547 4456 2824 4464
rect 2887 4456 2933 4464
rect 3056 4464 3064 4473
rect 3856 4467 3864 4493
rect 3887 4476 4013 4484
rect 4076 4484 4084 4516
rect 4147 4516 4253 4524
rect 4587 4516 4753 4524
rect 4887 4516 4953 4524
rect 4987 4516 5333 4524
rect 4107 4496 4264 4504
rect 4076 4476 4133 4484
rect 4167 4476 4233 4484
rect 4256 4484 4264 4496
rect 4287 4496 4373 4504
rect 4427 4496 4453 4504
rect 4527 4496 4573 4504
rect 4647 4496 4693 4504
rect 4747 4496 4793 4504
rect 4876 4496 4893 4504
rect 4256 4476 4304 4484
rect 4296 4467 4304 4476
rect 4447 4476 4473 4484
rect 4536 4476 4593 4484
rect 3027 4456 3064 4464
rect 3387 4456 3413 4464
rect 3487 4456 3513 4464
rect 4156 4456 4264 4464
rect -24 4436 13 4444
rect 27 4436 1053 4444
rect 1347 4436 1353 4444
rect 1367 4436 1473 4444
rect 1867 4436 1953 4444
rect 1996 4436 3013 4444
rect 487 4416 713 4424
rect 1467 4416 1573 4424
rect 1996 4424 2004 4436
rect 3456 4444 3464 4453
rect 3447 4436 3464 4444
rect 3767 4436 3833 4444
rect 4156 4444 4164 4456
rect 3947 4436 4164 4444
rect 4256 4444 4264 4456
rect 4256 4436 4273 4444
rect 4336 4444 4344 4473
rect 4396 4447 4404 4473
rect 4536 4467 4544 4476
rect 4627 4476 4684 4484
rect 4676 4464 4684 4476
rect 4876 4484 4884 4496
rect 5147 4496 5173 4504
rect 4787 4476 4884 4484
rect 4896 4476 4993 4484
rect 4896 4464 4904 4476
rect 5167 4476 5184 4484
rect 4607 4456 4644 4464
rect 4676 4456 4724 4464
rect 4307 4436 4344 4444
rect 4556 4444 4564 4453
rect 4507 4436 4564 4444
rect 4636 4444 4644 4456
rect 4716 4447 4724 4456
rect 4876 4456 4904 4464
rect 4916 4456 4953 4464
rect 4636 4436 4664 4444
rect 1587 4416 2004 4424
rect 2707 4416 2773 4424
rect 2787 4416 3253 4424
rect 3267 4416 3273 4424
rect 3287 4416 3353 4424
rect 3367 4416 3593 4424
rect 3607 4416 3733 4424
rect 3747 4416 3953 4424
rect 3967 4416 4033 4424
rect 4047 4416 4413 4424
rect 4427 4416 4633 4424
rect 4656 4424 4664 4436
rect 4876 4444 4884 4456
rect 4767 4436 4884 4444
rect 4916 4444 4924 4456
rect 5007 4456 5073 4464
rect 5096 4447 5104 4473
rect 5176 4464 5184 4476
rect 5176 4456 5193 4464
rect 4907 4436 4924 4444
rect 5156 4444 5164 4453
rect 5147 4436 5164 4444
rect 5256 4444 5264 4473
rect 5276 4467 5284 4516
rect 5427 4516 5573 4524
rect 5667 4516 5773 4524
rect 5907 4516 5913 4524
rect 5927 4516 5993 4524
rect 6167 4516 6353 4524
rect 6387 4516 6453 4524
rect 6507 4516 6573 4524
rect 5327 4496 5344 4504
rect 5336 4484 5344 4496
rect 5367 4496 5453 4504
rect 5547 4496 5704 4504
rect 5336 4476 5364 4484
rect 5356 4467 5364 4476
rect 5456 4476 5473 4484
rect 5456 4464 5464 4476
rect 5696 4484 5704 4496
rect 5747 4496 5993 4504
rect 5696 4476 5933 4484
rect 5396 4456 5464 4464
rect 5476 4456 5513 4464
rect 5256 4436 5293 4444
rect 4656 4416 4833 4424
rect 4867 4416 5353 4424
rect 5376 4424 5384 4433
rect 5367 4416 5384 4424
rect 347 4396 373 4404
rect 647 4396 813 4404
rect 3147 4396 4193 4404
rect 4287 4396 4453 4404
rect 4727 4396 4973 4404
rect 5067 4396 5273 4404
rect 5396 4404 5404 4456
rect 5427 4436 5453 4444
rect 5347 4396 5404 4404
rect 5476 4404 5484 4456
rect 5547 4456 5564 4464
rect 5556 4447 5564 4456
rect 5496 4436 5513 4444
rect 5496 4427 5504 4436
rect 5596 4424 5604 4473
rect 5707 4456 5773 4464
rect 5816 4444 5824 4476
rect 6056 4484 6064 4513
rect 6016 4476 6064 4484
rect 6076 4496 6093 4504
rect 5816 4436 5833 4444
rect 5936 4444 5944 4453
rect 5887 4436 5944 4444
rect 5547 4416 5604 4424
rect 5476 4396 5693 4404
rect 5756 4404 5764 4433
rect 5807 4416 5853 4424
rect 5876 4424 5884 4433
rect 5867 4416 5884 4424
rect 5956 4424 5964 4473
rect 6016 4467 6024 4476
rect 6076 4464 6084 4496
rect 6267 4496 6333 4504
rect 6347 4496 6633 4504
rect 6176 4476 6273 4484
rect 6176 4467 6184 4476
rect 6367 4476 6393 4484
rect 6547 4476 6613 4484
rect 6047 4456 6084 4464
rect 6336 4456 6433 4464
rect 5987 4436 6033 4444
rect 6336 4444 6344 4456
rect 6467 4456 6484 4464
rect 6327 4436 6344 4444
rect 6407 4436 6453 4444
rect 6476 4444 6484 4456
rect 6527 4456 6553 4464
rect 6607 4456 6653 4464
rect 6476 4436 6513 4444
rect 5956 4416 6113 4424
rect 6207 4416 6233 4424
rect 6247 4416 6293 4424
rect 6507 4416 6573 4424
rect 5756 4396 5873 4404
rect 5887 4396 5913 4404
rect 6107 4396 6313 4404
rect 1067 4376 3593 4384
rect 4187 4376 4253 4384
rect 4747 4376 4773 4384
rect 4907 4376 5093 4384
rect 5127 4376 5193 4384
rect 5207 4376 5373 4384
rect 5467 4376 5593 4384
rect 5767 4376 6073 4384
rect 6087 4376 6233 4384
rect 6287 4376 6553 4384
rect 3567 4356 3993 4364
rect 4007 4356 4053 4364
rect 4087 4356 4573 4364
rect 4587 4356 4964 4364
rect 3407 4336 3493 4344
rect 4447 4336 4793 4344
rect 4956 4344 4964 4356
rect 5007 4356 5133 4364
rect 5147 4356 5213 4364
rect 5527 4356 5633 4364
rect 6007 4356 6213 4364
rect 4956 4336 5133 4344
rect 5187 4336 5493 4344
rect 5567 4336 5713 4344
rect 5807 4336 6053 4344
rect 6067 4336 6313 4344
rect 6327 4336 6413 4344
rect 1467 4316 1493 4324
rect 2847 4316 2913 4324
rect 3827 4316 3853 4324
rect 3867 4316 3993 4324
rect 4007 4316 4073 4324
rect 4167 4316 4373 4324
rect 4407 4316 4693 4324
rect 4707 4316 4953 4324
rect 4976 4316 5653 4324
rect 4976 4304 4984 4316
rect 6027 4316 6093 4324
rect 6267 4316 6513 4324
rect 4067 4296 4984 4304
rect 5007 4296 5413 4304
rect 5487 4296 6453 4304
rect 4787 4276 4913 4284
rect 4987 4276 5793 4284
rect 6447 4276 6493 4284
rect 567 4256 593 4264
rect 707 4256 753 4264
rect 1287 4256 1673 4264
rect 1707 4256 1753 4264
rect 2687 4256 2733 4264
rect 3427 4256 3573 4264
rect 4147 4256 4673 4264
rect 4687 4256 4853 4264
rect 4887 4256 4993 4264
rect 5027 4256 5093 4264
rect 5127 4256 5473 4264
rect 5587 4256 5733 4264
rect 5747 4256 6433 4264
rect 6687 4256 6724 4264
rect 136 4236 153 4244
rect 136 4204 144 4236
rect 587 4236 593 4244
rect 607 4236 1073 4244
rect 1567 4236 1613 4244
rect 1667 4236 1773 4244
rect 3816 4236 3913 4244
rect 167 4216 373 4224
rect 447 4216 544 4224
rect -24 4184 -16 4204
rect 136 4196 184 4204
rect 176 4187 184 4196
rect 536 4204 544 4216
rect 587 4216 633 4224
rect 647 4216 793 4224
rect 827 4216 873 4224
rect 1096 4216 1273 4224
rect 287 4196 524 4204
rect 536 4196 553 4204
rect -24 4176 33 4184
rect 267 4176 433 4184
rect 516 4184 524 4196
rect 716 4196 1013 4204
rect 716 4184 724 4196
rect 1096 4204 1104 4216
rect 1327 4216 1353 4224
rect 1487 4216 1633 4224
rect 1687 4216 1713 4224
rect 1827 4216 1873 4224
rect 1887 4216 2093 4224
rect 3447 4216 3464 4224
rect 1067 4196 1104 4204
rect 1127 4196 1364 4204
rect 516 4176 724 4184
rect 736 4176 804 4184
rect 87 4156 273 4164
rect 427 4156 453 4164
rect 736 4164 744 4176
rect 467 4156 744 4164
rect 796 4164 804 4176
rect 867 4176 893 4184
rect 1027 4176 1133 4184
rect 1356 4184 1364 4196
rect 1387 4196 1513 4204
rect 1556 4196 1593 4204
rect 1356 4176 1473 4184
rect 1507 4176 1533 4184
rect 796 4156 893 4164
rect 907 4156 1213 4164
rect 1556 4164 1564 4196
rect 1607 4196 1653 4204
rect 1756 4204 1764 4213
rect 1756 4196 1793 4204
rect 2127 4196 2193 4204
rect 2247 4196 2773 4204
rect 1656 4176 1793 4184
rect 1656 4167 1664 4176
rect 2007 4176 2213 4184
rect 2367 4176 2424 4184
rect 1547 4156 1564 4164
rect 1767 4156 1953 4164
rect 1967 4156 2173 4164
rect 2187 4156 2393 4164
rect 2416 4164 2424 4176
rect 2487 4176 2533 4184
rect 2727 4176 2753 4184
rect 2796 4184 2804 4213
rect 2827 4196 2853 4204
rect 3067 4196 3093 4204
rect 3416 4204 3424 4213
rect 3107 4196 3384 4204
rect 3416 4196 3433 4204
rect 2787 4176 2804 4184
rect 2416 4156 2693 4164
rect 2747 4156 2873 4164
rect 2896 4164 2904 4193
rect 3376 4187 3384 4196
rect 3456 4204 3464 4216
rect 3516 4207 3524 4233
rect 3456 4196 3484 4204
rect 2927 4176 2964 4184
rect 2896 4156 2913 4164
rect 2956 4164 2964 4176
rect 3436 4176 3453 4184
rect 2956 4156 3013 4164
rect 3287 4156 3413 4164
rect 247 4136 373 4144
rect 687 4136 933 4144
rect 1587 4136 1693 4144
rect 1707 4136 2013 4144
rect 2027 4136 2113 4144
rect 2127 4136 2153 4144
rect 2167 4136 2213 4144
rect 2227 4136 2253 4144
rect 2547 4136 2593 4144
rect 3436 4144 3444 4176
rect 3476 4164 3484 4196
rect 3747 4196 3784 4204
rect 3776 4184 3784 4196
rect 3816 4204 3824 4236
rect 4067 4236 4273 4244
rect 4687 4236 4813 4244
rect 4847 4236 5053 4244
rect 5207 4236 5233 4244
rect 5367 4236 5673 4244
rect 5707 4236 5793 4244
rect 5947 4236 6173 4244
rect 6567 4236 6624 4244
rect 4487 4216 4753 4224
rect 4767 4216 4893 4224
rect 4907 4216 4973 4224
rect 5047 4216 5113 4224
rect 5147 4216 5393 4224
rect 5416 4216 5573 4224
rect 3807 4196 3824 4204
rect 4047 4196 4073 4204
rect 4287 4196 4724 4204
rect 3776 4176 3813 4184
rect 3987 4176 4093 4184
rect 3467 4156 3484 4164
rect 3496 4156 4053 4164
rect 3496 4144 3504 4156
rect 4196 4164 4204 4193
rect 4227 4176 4253 4184
rect 4567 4176 4693 4184
rect 4716 4184 4724 4196
rect 5007 4196 5053 4204
rect 5147 4196 5193 4204
rect 5416 4204 5424 4216
rect 5587 4216 5753 4224
rect 5307 4196 5424 4204
rect 5447 4196 5573 4204
rect 5587 4196 5613 4204
rect 5796 4204 5804 4213
rect 5676 4196 5804 4204
rect 5856 4204 5864 4233
rect 5887 4216 5953 4224
rect 6047 4216 6133 4224
rect 6207 4216 6244 4224
rect 5856 4196 5873 4204
rect 4716 4176 4933 4184
rect 4976 4184 4984 4193
rect 4976 4176 5013 4184
rect 5227 4176 5353 4184
rect 5396 4176 5473 4184
rect 4196 4156 4213 4164
rect 4527 4156 4593 4164
rect 4987 4156 5113 4164
rect 5167 4156 5333 4164
rect 5396 4164 5404 4176
rect 5676 4184 5684 4196
rect 5896 4196 5993 4204
rect 5567 4176 5684 4184
rect 5727 4176 5733 4184
rect 5747 4176 5773 4184
rect 5896 4184 5904 4196
rect 6196 4204 6204 4213
rect 6087 4196 6204 4204
rect 6236 4204 6244 4216
rect 6307 4216 6324 4224
rect 6316 4204 6324 4216
rect 6347 4216 6373 4224
rect 6527 4216 6593 4224
rect 6616 4207 6624 4236
rect 6676 4236 6693 4244
rect 6236 4196 6304 4204
rect 6316 4196 6384 4204
rect 6296 4187 6304 4196
rect 5847 4176 5904 4184
rect 5987 4176 6013 4184
rect 6027 4176 6073 4184
rect 6167 4176 6273 4184
rect 6376 4184 6384 4196
rect 6407 4196 6433 4204
rect 6487 4196 6553 4204
rect 6376 4176 6513 4184
rect 6576 4167 6584 4193
rect 6596 4184 6604 4193
rect 6596 4176 6653 4184
rect 5347 4156 5404 4164
rect 5427 4156 5633 4164
rect 5827 4156 6013 4164
rect 6027 4156 6333 4164
rect 6347 4156 6353 4164
rect 6587 4156 6613 4164
rect 6676 4164 6684 4236
rect 6647 4156 6684 4164
rect 3436 4136 3504 4144
rect 3587 4136 3873 4144
rect 3927 4136 4013 4144
rect 4027 4136 4133 4144
rect 4147 4136 4173 4144
rect 4187 4136 5093 4144
rect 5287 4136 5833 4144
rect 6187 4136 6213 4144
rect 6716 4144 6724 4256
rect 6667 4136 6724 4144
rect 367 4116 413 4124
rect 687 4116 773 4124
rect 787 4116 873 4124
rect 1267 4116 1613 4124
rect 1747 4116 2933 4124
rect 2947 4116 3153 4124
rect 3407 4116 3553 4124
rect 3567 4116 3753 4124
rect 4127 4116 4353 4124
rect 4947 4116 5173 4124
rect 5187 4116 5253 4124
rect 5307 4116 5593 4124
rect 5707 4116 5913 4124
rect 6107 4116 6173 4124
rect 727 4096 793 4104
rect 5267 4096 5353 4104
rect 5367 4096 5453 4104
rect 5707 4096 5773 4104
rect 5907 4096 6053 4104
rect 1627 4076 2573 4084
rect 2587 4076 2713 4084
rect 4227 4076 6533 4084
rect 907 4056 1253 4064
rect 2947 4056 2973 4064
rect 3687 4056 3913 4064
rect 3927 4056 3933 4064
rect 4247 4056 4333 4064
rect 4347 4056 4764 4064
rect 176 4036 693 4044
rect 176 4024 184 4036
rect 1087 4036 1313 4044
rect 1327 4036 1364 4044
rect -24 4016 184 4024
rect -24 3996 -16 4016
rect 207 4016 453 4024
rect 567 4016 613 4024
rect 747 4016 1133 4024
rect 1307 4016 1324 4024
rect 87 3996 113 4004
rect 247 3996 433 4004
rect 476 4004 484 4013
rect 476 3996 633 4004
rect 747 3996 773 4004
rect 1127 3996 1133 4004
rect 1147 3996 1244 4004
rect 367 3976 384 3984
rect -24 3956 53 3964
rect 127 3956 333 3964
rect 376 3964 384 3976
rect 427 3976 453 3984
rect 576 3976 633 3984
rect 576 3967 584 3976
rect 1076 3984 1084 3993
rect 1056 3976 1084 3984
rect 376 3956 493 3964
rect 507 3956 533 3964
rect 667 3956 773 3964
rect 787 3956 1013 3964
rect 387 3936 593 3944
rect 1036 3944 1044 3973
rect 1056 3967 1064 3976
rect 1107 3976 1124 3984
rect 1036 3936 1053 3944
rect 1067 3936 1073 3944
rect 467 3916 753 3924
rect 1116 3904 1124 3976
rect 1236 3984 1244 3996
rect 1187 3976 1224 3984
rect 1236 3976 1273 3984
rect 1136 3956 1153 3964
rect 1136 3927 1144 3956
rect 1216 3964 1224 3976
rect 1316 3984 1324 4016
rect 1356 4007 1364 4036
rect 1467 4036 1653 4044
rect 1667 4036 1833 4044
rect 2587 4036 2633 4044
rect 2927 4036 2993 4044
rect 3007 4036 3173 4044
rect 3227 4036 3773 4044
rect 4107 4036 4233 4044
rect 4487 4036 4613 4044
rect 4756 4044 4764 4056
rect 4927 4056 5273 4064
rect 5427 4056 5513 4064
rect 5547 4056 5853 4064
rect 4756 4036 6693 4044
rect 1447 4016 1713 4024
rect 1727 4016 1753 4024
rect 1767 4016 1913 4024
rect 2516 4016 2553 4024
rect 1496 3996 1644 4004
rect 1496 3984 1504 3996
rect 1316 3976 1504 3984
rect 1636 3984 1644 3996
rect 1967 3996 2173 4004
rect 2196 3996 2333 4004
rect 2196 3987 2204 3996
rect 2387 3996 2493 4004
rect 2516 3987 2524 4016
rect 2607 4016 2613 4024
rect 2627 4016 2673 4024
rect 2827 4016 2844 4024
rect 2836 4004 2844 4016
rect 2967 4016 3013 4024
rect 3027 4016 3093 4024
rect 3527 4016 3624 4024
rect 2836 3996 2904 4004
rect 1636 3976 1753 3984
rect 1636 3967 1644 3976
rect 2087 3976 2153 3984
rect 2287 3976 2324 3984
rect 2316 3967 2324 3976
rect 2427 3976 2473 3984
rect 2536 3984 2544 3993
rect 2536 3976 2613 3984
rect 2696 3984 2704 3993
rect 2696 3976 2733 3984
rect 2787 3976 2873 3984
rect 2896 3984 2904 3996
rect 3147 3996 3193 4004
rect 3287 3996 3473 4004
rect 3567 3996 3593 4004
rect 3616 4004 3624 4016
rect 3756 4016 3813 4024
rect 3756 4004 3764 4016
rect 4027 4016 4113 4024
rect 4127 4016 4153 4024
rect 4387 4016 5293 4024
rect 5507 4016 5533 4024
rect 5607 4016 5824 4024
rect 5816 4007 5824 4016
rect 5847 4016 6153 4024
rect 3616 3996 3764 4004
rect 4007 3996 4153 4004
rect 4687 3996 4733 4004
rect 4747 3996 4853 4004
rect 4907 3996 5033 4004
rect 5207 3996 5293 4004
rect 5507 3996 5673 4004
rect 5827 3996 6013 4004
rect 6047 3996 6173 4004
rect 6227 3996 6273 4004
rect 2896 3976 3013 3984
rect 3036 3967 3044 3993
rect 3067 3976 3113 3984
rect 3296 3976 3353 3984
rect 3296 3967 3304 3976
rect 3987 3976 4053 3984
rect 4256 3984 4264 3993
rect 4187 3976 4313 3984
rect 4407 3976 4453 3984
rect 4827 3976 4873 3984
rect 5167 3976 5273 3984
rect 1216 3956 1313 3964
rect 1327 3956 1593 3964
rect 1787 3956 1833 3964
rect 1847 3956 2053 3964
rect 2807 3956 2853 3964
rect 2907 3956 2973 3964
rect 3216 3956 3253 3964
rect 1547 3936 1733 3944
rect 2267 3936 2413 3944
rect 2427 3936 2453 3944
rect 3216 3944 3224 3956
rect 3327 3956 3653 3964
rect 4327 3956 4353 3964
rect 4447 3956 4493 3964
rect 4787 3956 4913 3964
rect 2727 3936 3224 3944
rect 3247 3936 3333 3944
rect 3807 3936 3833 3944
rect 3847 3936 4373 3944
rect 4747 3936 4793 3944
rect 5316 3944 5324 3993
rect 5487 3976 5553 3984
rect 5876 3976 6004 3984
rect 5347 3956 5573 3964
rect 5587 3956 5633 3964
rect 5687 3956 5833 3964
rect 5876 3964 5884 3976
rect 5867 3956 5884 3964
rect 5907 3956 5933 3964
rect 5996 3964 6004 3976
rect 5996 3956 6413 3964
rect 5316 3936 5773 3944
rect 5976 3944 5984 3953
rect 5887 3936 5984 3944
rect 2767 3916 3953 3924
rect 4047 3916 4093 3924
rect 5507 3916 5533 3924
rect 5647 3916 6573 3924
rect 1116 3896 1413 3904
rect 4507 3896 6133 3904
rect 6147 3896 6153 3904
rect 3627 3876 4713 3884
rect 4867 3876 5553 3884
rect 5807 3876 5853 3884
rect 3987 3856 4113 3864
rect 5247 3856 5253 3864
rect 5267 3856 5273 3864
rect 5287 3856 5433 3864
rect 5627 3856 6033 3864
rect 2307 3836 2633 3844
rect 4927 3836 6073 3844
rect 1087 3816 1113 3824
rect 2647 3816 2893 3824
rect 2587 3796 2753 3804
rect 2767 3796 2873 3804
rect 3127 3796 3333 3804
rect 3727 3796 3833 3804
rect 4307 3796 4593 3804
rect 5227 3796 5253 3804
rect 6467 3796 6493 3804
rect 587 3776 653 3784
rect 687 3776 753 3784
rect 767 3776 773 3784
rect 827 3776 853 3784
rect 1847 3776 2293 3784
rect 2307 3776 2393 3784
rect 2807 3776 3173 3784
rect 3467 3776 3533 3784
rect 3707 3776 3953 3784
rect 4967 3776 5153 3784
rect 5167 3776 5393 3784
rect 6087 3776 6113 3784
rect 6267 3776 6413 3784
rect 6507 3776 6653 3784
rect 207 3756 593 3764
rect 607 3756 773 3764
rect 787 3756 1193 3764
rect 1507 3756 1544 3764
rect -24 3724 -16 3744
rect 547 3736 604 3744
rect -24 3716 4 3724
rect -4 3704 4 3716
rect 227 3716 573 3724
rect 596 3724 604 3736
rect 747 3736 1113 3744
rect 1187 3736 1233 3744
rect 1327 3736 1413 3744
rect 1427 3736 1453 3744
rect 596 3716 733 3724
rect 807 3716 1073 3724
rect 1236 3716 1373 3724
rect -24 3684 -16 3704
rect -4 3696 33 3704
rect 167 3696 253 3704
rect 407 3696 513 3704
rect 536 3696 833 3704
rect -24 3676 113 3684
rect 367 3676 473 3684
rect 536 3684 544 3696
rect 867 3696 893 3704
rect 1236 3704 1244 3716
rect 1167 3696 1244 3704
rect 1256 3696 1313 3704
rect 487 3676 544 3684
rect 567 3676 693 3684
rect 836 3684 844 3693
rect 836 3676 933 3684
rect 1256 3684 1264 3696
rect 1347 3696 1353 3704
rect 1516 3704 1524 3733
rect 1536 3727 1544 3756
rect 1927 3756 1973 3764
rect 2156 3756 2373 3764
rect 1907 3736 1933 3744
rect 2107 3736 2133 3744
rect 1976 3716 2044 3724
rect 1376 3696 1524 3704
rect 1227 3676 1264 3684
rect 1376 3684 1384 3696
rect 1747 3696 1773 3704
rect 1816 3696 1833 3704
rect 1816 3687 1824 3696
rect 1976 3704 1984 3716
rect 2036 3707 2044 3716
rect 1907 3696 1984 3704
rect 2067 3696 2133 3704
rect 2156 3687 2164 3756
rect 2387 3756 2613 3764
rect 2847 3756 2913 3764
rect 2987 3756 3093 3764
rect 3287 3756 3313 3764
rect 3387 3756 3673 3764
rect 3687 3756 3793 3764
rect 4487 3756 4533 3764
rect 4607 3756 4753 3764
rect 4767 3756 4893 3764
rect 4907 3756 5093 3764
rect 5107 3756 5373 3764
rect 5387 3756 5513 3764
rect 5527 3756 5593 3764
rect 5607 3756 5713 3764
rect 5727 3756 6093 3764
rect 6107 3756 6373 3764
rect 6387 3756 6513 3764
rect 2596 3736 2673 3744
rect 2256 3716 2293 3724
rect 2256 3704 2264 3716
rect 2527 3716 2573 3724
rect 2207 3696 2264 3704
rect 2396 3687 2404 3713
rect 1307 3676 1384 3684
rect 1407 3676 1533 3684
rect 1847 3676 1873 3684
rect 2227 3676 2273 3684
rect 2307 3676 2353 3684
rect 87 3656 893 3664
rect 927 3656 1253 3664
rect 1587 3656 1673 3664
rect 2416 3664 2424 3713
rect 2596 3707 2604 3736
rect 2787 3736 2813 3744
rect 2907 3736 2964 3744
rect 2956 3727 2964 3736
rect 3047 3736 3064 3744
rect 2627 3716 2773 3724
rect 2976 3716 3013 3724
rect 2767 3696 2893 3704
rect 2976 3704 2984 3716
rect 3056 3707 3064 3736
rect 3147 3736 3233 3744
rect 3247 3736 3313 3744
rect 3087 3716 3113 3724
rect 3187 3716 3233 3724
rect 3336 3724 3344 3753
rect 3747 3736 3804 3744
rect 3336 3716 3353 3724
rect 3447 3716 3493 3724
rect 3547 3716 3753 3724
rect 2967 3696 2984 3704
rect 3167 3696 3213 3704
rect 2807 3676 2853 3684
rect 2867 3676 3113 3684
rect 3247 3676 3293 3684
rect 3307 3676 3313 3684
rect 3796 3684 3804 3736
rect 4087 3736 4173 3744
rect 4476 3736 4493 3744
rect 3887 3716 3933 3724
rect 3967 3716 3993 3724
rect 4127 3716 4413 3724
rect 4476 3724 4484 3736
rect 4727 3736 5333 3744
rect 5347 3736 5373 3744
rect 5947 3736 6273 3744
rect 6307 3736 6313 3744
rect 6327 3736 6633 3744
rect 4436 3716 4484 3724
rect 4107 3696 4233 3704
rect 4367 3696 4373 3704
rect 4436 3704 4444 3716
rect 4556 3724 4564 3733
rect 4527 3716 4564 3724
rect 5067 3716 5133 3724
rect 5287 3716 5353 3724
rect 5487 3716 5513 3724
rect 5656 3716 5773 3724
rect 5656 3707 5664 3716
rect 4387 3696 4444 3704
rect 4847 3696 5033 3704
rect 3787 3676 3913 3684
rect 5167 3676 5213 3684
rect 5536 3684 5544 3693
rect 5307 3676 5544 3684
rect 5796 3684 5804 3713
rect 5816 3704 5824 3733
rect 5856 3716 5913 3724
rect 5856 3704 5864 3716
rect 6107 3716 6153 3724
rect 6287 3716 6553 3724
rect 5816 3696 5864 3704
rect 6016 3704 6024 3713
rect 5927 3696 6024 3704
rect 6196 3704 6204 3713
rect 6187 3696 6204 3704
rect 6216 3687 6224 3713
rect 6236 3687 6244 3713
rect 6327 3696 6353 3704
rect 6447 3696 6573 3704
rect 5796 3676 5833 3684
rect 5947 3676 5953 3684
rect 5967 3676 6053 3684
rect 6087 3676 6193 3684
rect 6207 3676 6213 3684
rect 1887 3656 3053 3664
rect 3207 3656 3253 3664
rect 3307 3656 5353 3664
rect 6027 3656 6173 3664
rect 6187 3656 6353 3664
rect 507 3636 553 3644
rect 707 3636 733 3644
rect 1067 3636 1093 3644
rect 1116 3636 1133 3644
rect 467 3616 633 3624
rect 1116 3624 1124 3636
rect 1507 3636 1593 3644
rect 1687 3636 2073 3644
rect 2627 3636 6033 3644
rect 6047 3636 6133 3644
rect 6147 3636 6213 3644
rect 6227 3636 6233 3644
rect 6427 3636 6633 3644
rect 987 3616 1124 3624
rect 1807 3616 2173 3624
rect 2247 3616 2533 3624
rect 2547 3616 2673 3624
rect 2947 3616 2993 3624
rect 3047 3616 3553 3624
rect 3727 3616 3913 3624
rect 5807 3616 6153 3624
rect 6167 3616 6533 3624
rect 427 3596 453 3604
rect 1487 3596 1913 3604
rect 1927 3596 1993 3604
rect 3367 3596 3393 3604
rect 3727 3596 3893 3604
rect 3907 3596 4053 3604
rect 4067 3596 4453 3604
rect 4467 3596 4993 3604
rect 5007 3596 5093 3604
rect 6267 3596 6333 3604
rect 6467 3596 6573 3604
rect 247 3576 513 3584
rect 567 3576 853 3584
rect 1167 3576 1293 3584
rect 1927 3576 1953 3584
rect 2687 3576 2973 3584
rect 2987 3576 3033 3584
rect 5067 3576 5313 3584
rect 5807 3576 5873 3584
rect 427 3556 733 3564
rect 747 3556 753 3564
rect 967 3556 1033 3564
rect 1127 3556 1173 3564
rect 1347 3556 1373 3564
rect 1947 3556 1973 3564
rect 2067 3556 2093 3564
rect 2567 3556 2813 3564
rect 3667 3556 3953 3564
rect 4007 3556 4013 3564
rect 4027 3556 4033 3564
rect 4307 3556 4373 3564
rect 4387 3556 5233 3564
rect 5636 3556 5693 3564
rect 207 3536 473 3544
rect 807 3536 1024 3544
rect -24 3516 33 3524
rect 87 3516 113 3524
rect 327 3516 413 3524
rect 536 3516 693 3524
rect 536 3507 544 3516
rect 707 3516 713 3524
rect 787 3516 813 3524
rect 827 3516 933 3524
rect 956 3516 973 3524
rect -24 3496 213 3504
rect -24 3476 -16 3496
rect 787 3496 853 3504
rect 956 3504 964 3516
rect 1016 3524 1024 3536
rect 1207 3536 1433 3544
rect 1647 3536 1733 3544
rect 1747 3536 1904 3544
rect 1016 3516 1064 3524
rect 927 3496 964 3504
rect 1056 3504 1064 3516
rect 1187 3516 1233 3524
rect 1447 3516 1513 3524
rect 1527 3516 1553 3524
rect 1627 3516 1673 3524
rect 1827 3516 1853 3524
rect 1896 3524 1904 3536
rect 1956 3536 2144 3544
rect 1956 3524 1964 3536
rect 1896 3516 1964 3524
rect 1976 3516 2073 3524
rect 1056 3496 1133 3504
rect 1347 3496 1733 3504
rect 1976 3504 1984 3516
rect 2136 3524 2144 3536
rect 2376 3536 2433 3544
rect 2376 3527 2384 3536
rect 2507 3536 2553 3544
rect 2567 3536 2633 3544
rect 2767 3536 2853 3544
rect 2887 3536 2973 3544
rect 2987 3536 3024 3544
rect 2136 3516 2184 3524
rect 1907 3496 1984 3504
rect 2007 3496 2133 3504
rect 2176 3504 2184 3516
rect 2267 3516 2293 3524
rect 2847 3516 2913 3524
rect 3016 3524 3024 3536
rect 3047 3536 3093 3544
rect 3147 3536 3153 3544
rect 3167 3536 3233 3544
rect 3247 3536 3273 3544
rect 4367 3536 4613 3544
rect 4656 3536 4733 3544
rect 4656 3527 4664 3536
rect 4927 3536 5013 3544
rect 5287 3536 5513 3544
rect 5636 3544 5644 3556
rect 5767 3556 5853 3564
rect 5907 3556 5973 3564
rect 5596 3536 5644 3544
rect 3016 3516 3044 3524
rect 3036 3507 3044 3516
rect 3087 3516 3193 3524
rect 3247 3516 3493 3524
rect 3587 3516 3613 3524
rect 3747 3516 3773 3524
rect 4116 3516 4153 3524
rect 2176 3496 2433 3504
rect 2707 3496 2793 3504
rect 2807 3496 3013 3504
rect 3067 3496 3153 3504
rect 3267 3496 3313 3504
rect 3347 3496 3644 3504
rect 127 3476 333 3484
rect 356 3464 364 3493
rect 387 3476 593 3484
rect 356 3456 573 3464
rect 587 3456 613 3464
rect 636 3464 644 3493
rect 1007 3476 1513 3484
rect 1827 3476 2093 3484
rect 2107 3476 2213 3484
rect 2227 3476 2353 3484
rect 2767 3476 2913 3484
rect 3107 3476 3133 3484
rect 3636 3484 3644 3496
rect 3687 3496 3973 3504
rect 4116 3504 4124 3516
rect 4356 3516 4373 3524
rect 4356 3507 4364 3516
rect 4696 3516 4884 3524
rect 4007 3496 4124 3504
rect 4147 3496 4273 3504
rect 4376 3496 4393 3504
rect 3636 3476 4333 3484
rect 4376 3484 4384 3496
rect 4696 3504 4704 3516
rect 4627 3496 4704 3504
rect 4876 3504 4884 3516
rect 4907 3516 4953 3524
rect 5596 3524 5604 3536
rect 5667 3536 5733 3544
rect 5747 3536 5753 3544
rect 5776 3536 5844 3544
rect 5056 3516 5304 3524
rect 5056 3504 5064 3516
rect 4876 3496 5064 3504
rect 5087 3496 5133 3504
rect 5296 3504 5304 3516
rect 5556 3516 5604 3524
rect 5296 3496 5433 3504
rect 5556 3487 5564 3516
rect 5627 3516 5653 3524
rect 5776 3524 5784 3536
rect 5727 3516 5784 3524
rect 5836 3524 5844 3536
rect 5907 3536 5933 3544
rect 5956 3536 6053 3544
rect 5956 3524 5964 3536
rect 6207 3536 6253 3544
rect 5836 3516 5964 3524
rect 5587 3496 5713 3504
rect 5847 3496 5873 3504
rect 5907 3496 5953 3504
rect 5976 3487 5984 3513
rect 4356 3476 4384 3484
rect 636 3456 653 3464
rect 687 3456 773 3464
rect 2847 3456 2893 3464
rect 3047 3456 3213 3464
rect 3527 3456 3633 3464
rect 4356 3464 4364 3476
rect 4527 3476 4713 3484
rect 5687 3476 5773 3484
rect 6016 3484 6024 3513
rect 6016 3476 6033 3484
rect 4327 3456 4364 3464
rect 4387 3456 4473 3464
rect 5287 3456 5633 3464
rect 5876 3456 6533 3464
rect 227 3436 1053 3444
rect 2787 3436 2853 3444
rect 2887 3436 3693 3444
rect 5876 3444 5884 3456
rect 5767 3436 5884 3444
rect 6267 3436 6293 3444
rect 2667 3416 3113 3424
rect 3127 3416 3253 3424
rect 3967 3416 4973 3424
rect 5387 3416 5633 3424
rect 6047 3416 6133 3424
rect 6147 3416 6293 3424
rect 6596 3407 6604 3593
rect 2407 3396 3573 3404
rect 3707 3396 4804 3404
rect 3087 3376 3233 3384
rect 3447 3376 3473 3384
rect 4427 3376 4753 3384
rect 4767 3376 4773 3384
rect 4796 3384 4804 3396
rect 4796 3376 5693 3384
rect 5867 3376 6233 3384
rect 3047 3356 4713 3364
rect 4907 3356 5293 3364
rect 5547 3356 5973 3364
rect 6007 3356 6013 3364
rect 6027 3356 6073 3364
rect 6087 3356 6193 3364
rect 6207 3356 6373 3364
rect 2287 3336 2593 3344
rect 2967 3336 5613 3344
rect 5707 3336 5873 3344
rect 627 3316 833 3324
rect 907 3316 1013 3324
rect 1027 3316 1113 3324
rect 1267 3316 2233 3324
rect 3067 3316 4393 3324
rect 4487 3316 4553 3324
rect 4727 3316 5313 3324
rect 5327 3316 5673 3324
rect 6227 3316 6333 3324
rect 427 3296 493 3304
rect 587 3296 633 3304
rect 887 3296 1273 3304
rect 1287 3296 1373 3304
rect 1787 3296 1864 3304
rect 387 3276 593 3284
rect 667 3276 973 3284
rect 316 3256 333 3264
rect -24 3224 -16 3244
rect 316 3244 324 3256
rect 467 3256 633 3264
rect 656 3247 664 3273
rect 727 3256 753 3264
rect 896 3256 913 3264
rect 127 3236 324 3244
rect 367 3236 413 3244
rect 707 3236 764 3244
rect -24 3216 33 3224
rect 87 3216 113 3224
rect 247 3216 433 3224
rect 476 3224 484 3233
rect 456 3216 484 3224
rect 456 3207 464 3216
rect 527 3216 553 3224
rect 596 3224 604 3233
rect 756 3227 764 3236
rect 587 3216 604 3224
rect 647 3216 693 3224
rect 707 3216 733 3224
rect 827 3216 873 3224
rect 896 3207 904 3256
rect 967 3256 1053 3264
rect 1707 3256 1813 3264
rect 916 3236 953 3244
rect 916 3227 924 3236
rect 1247 3236 1293 3244
rect 1607 3236 1733 3244
rect 1836 3244 1844 3273
rect 1856 3267 1864 3296
rect 2867 3296 2913 3304
rect 2927 3296 3153 3304
rect 3607 3296 3953 3304
rect 4247 3296 5473 3304
rect 5507 3296 5673 3304
rect 5847 3296 6133 3304
rect 6167 3296 6253 3304
rect 2747 3276 2873 3284
rect 2907 3276 2933 3284
rect 2947 3276 2973 3284
rect 3027 3276 3193 3284
rect 3427 3276 3773 3284
rect 4567 3276 4593 3284
rect 4687 3276 4813 3284
rect 4827 3276 4993 3284
rect 5227 3276 5833 3284
rect 6067 3276 6093 3284
rect 6136 3276 6253 3284
rect 2207 3256 2233 3264
rect 2927 3256 3033 3264
rect 3567 3256 3693 3264
rect 3707 3256 3713 3264
rect 3867 3256 4584 3264
rect 1836 3236 1853 3244
rect 927 3216 1073 3224
rect 1196 3224 1204 3233
rect 1167 3216 1204 3224
rect 1227 3216 1493 3224
rect 1527 3216 1613 3224
rect 1776 3224 1784 3233
rect 1776 3216 1813 3224
rect 1896 3224 1904 3233
rect 1847 3216 1904 3224
rect 487 3196 553 3204
rect 567 3196 633 3204
rect 947 3196 973 3204
rect 1667 3196 1713 3204
rect 1916 3204 1924 3233
rect 2367 3216 2413 3224
rect 2487 3216 2513 3224
rect 1767 3196 1924 3204
rect 1936 3196 2404 3204
rect 527 3176 593 3184
rect 607 3176 673 3184
rect 1936 3184 1944 3196
rect 807 3176 1944 3184
rect 2327 3176 2373 3184
rect 2396 3184 2404 3196
rect 2447 3196 2493 3204
rect 2536 3204 2544 3233
rect 2556 3227 2564 3253
rect 2876 3227 2884 3253
rect 3007 3236 3053 3244
rect 3076 3244 3084 3253
rect 3076 3236 3093 3244
rect 3187 3236 3293 3244
rect 3407 3236 3464 3244
rect 3456 3227 3464 3236
rect 3516 3236 3573 3244
rect 2807 3216 2833 3224
rect 3047 3216 3073 3224
rect 3127 3216 3213 3224
rect 3227 3216 3353 3224
rect 3516 3224 3524 3236
rect 3616 3236 3713 3244
rect 3507 3216 3524 3224
rect 2536 3196 2553 3204
rect 2907 3196 2964 3204
rect 2396 3176 2933 3184
rect 2956 3184 2964 3196
rect 3267 3196 3453 3204
rect 3487 3196 3513 3204
rect 3616 3204 3624 3236
rect 3836 3244 3844 3253
rect 3736 3236 3844 3244
rect 3736 3224 3744 3236
rect 4067 3236 4093 3244
rect 4187 3236 4473 3244
rect 4416 3227 4424 3236
rect 4576 3244 4584 3256
rect 5007 3256 5173 3264
rect 5427 3256 5473 3264
rect 5507 3256 5693 3264
rect 6136 3264 6144 3276
rect 6307 3276 6333 3284
rect 6567 3276 6613 3284
rect 5747 3256 6144 3264
rect 6156 3256 6233 3264
rect 4576 3236 4684 3244
rect 3656 3216 3744 3224
rect 3656 3207 3664 3216
rect 3907 3216 3933 3224
rect 4127 3216 4253 3224
rect 4476 3216 4533 3224
rect 4476 3207 4484 3216
rect 4587 3216 4644 3224
rect 4636 3207 4644 3216
rect 3616 3196 3633 3204
rect 3687 3196 3693 3204
rect 3707 3196 3753 3204
rect 3947 3196 4013 3204
rect 4087 3196 4433 3204
rect 4507 3196 4613 3204
rect 4676 3204 4684 3236
rect 4696 3236 4713 3244
rect 4696 3227 4704 3236
rect 4807 3236 4853 3244
rect 4956 3244 4964 3253
rect 4936 3236 4964 3244
rect 4896 3216 4913 3224
rect 4676 3196 4713 3204
rect 4896 3204 4904 3216
rect 4867 3196 4904 3204
rect 4936 3204 4944 3236
rect 4987 3236 5253 3244
rect 5367 3236 5393 3244
rect 5436 3236 5493 3244
rect 5436 3227 5444 3236
rect 5787 3236 5833 3244
rect 6156 3244 6164 3256
rect 6267 3256 6324 3264
rect 6107 3236 6164 3244
rect 6316 3244 6324 3256
rect 6387 3256 6513 3264
rect 6316 3236 6404 3244
rect 5167 3216 5273 3224
rect 5756 3224 5764 3233
rect 5456 3216 5564 3224
rect 5756 3216 5813 3224
rect 4927 3196 4944 3204
rect 4996 3196 5333 3204
rect 4996 3184 5004 3196
rect 5456 3204 5464 3216
rect 5387 3196 5464 3204
rect 5556 3204 5564 3216
rect 5876 3216 5944 3224
rect 5876 3204 5884 3216
rect 5556 3196 5884 3204
rect 5936 3204 5944 3216
rect 5976 3216 6024 3224
rect 5976 3204 5984 3216
rect 5936 3196 5984 3204
rect 6016 3204 6024 3216
rect 6047 3216 6113 3224
rect 6276 3224 6284 3233
rect 6396 3227 6404 3236
rect 6427 3236 6473 3244
rect 6496 3236 6553 3244
rect 6247 3216 6284 3224
rect 6336 3216 6373 3224
rect 6016 3196 6133 3204
rect 6336 3204 6344 3216
rect 6496 3224 6504 3236
rect 6447 3216 6504 3224
rect 6527 3216 6553 3224
rect 6287 3196 6344 3204
rect 6367 3196 6453 3204
rect 6596 3204 6604 3253
rect 6596 3196 6613 3204
rect 2956 3176 5004 3184
rect 5227 3176 5833 3184
rect 6147 3176 6353 3184
rect 6387 3176 6553 3184
rect 6636 3167 6644 3253
rect 767 3156 1033 3164
rect 1076 3156 1173 3164
rect 1076 3144 1084 3156
rect 1807 3156 1913 3164
rect 2847 3156 2913 3164
rect 3347 3156 3373 3164
rect 3407 3156 3453 3164
rect 3487 3156 5053 3164
rect 5136 3156 5293 3164
rect 1027 3136 1084 3144
rect 1307 3136 1333 3144
rect 2807 3136 3333 3144
rect 3427 3136 3553 3144
rect 3916 3136 4344 3144
rect 3916 3124 3924 3136
rect 2507 3116 3924 3124
rect 4336 3124 4344 3136
rect 4407 3136 4433 3144
rect 4507 3136 4753 3144
rect 5136 3144 5144 3156
rect 5347 3156 5373 3164
rect 5567 3156 5793 3164
rect 5927 3156 6253 3164
rect 6267 3156 6293 3164
rect 6447 3156 6573 3164
rect 5047 3136 5144 3144
rect 5167 3136 5413 3144
rect 5427 3136 5553 3144
rect 5787 3136 5953 3144
rect 6007 3136 6153 3144
rect 6167 3136 6453 3144
rect 6467 3136 6553 3144
rect 4287 3116 4324 3124
rect 4336 3116 5373 3124
rect 387 3096 733 3104
rect 767 3096 1293 3104
rect 1767 3096 1993 3104
rect 2927 3096 2953 3104
rect 3167 3096 3273 3104
rect 3307 3096 3493 3104
rect 3707 3096 3913 3104
rect 3987 3096 4053 3104
rect 4267 3096 4293 3104
rect 4316 3104 4324 3116
rect 5527 3116 5733 3124
rect 5947 3116 6073 3124
rect 6507 3116 6533 3124
rect 4316 3096 4413 3104
rect 4456 3096 4493 3104
rect 687 3076 773 3084
rect 987 3076 1033 3084
rect 1527 3076 1713 3084
rect 1787 3076 1873 3084
rect 2076 3076 2253 3084
rect 527 3056 673 3064
rect 947 3056 973 3064
rect 1167 3056 1453 3064
rect 1467 3056 1473 3064
rect 1547 3056 1653 3064
rect 1847 3056 1953 3064
rect -24 3036 233 3044
rect -24 2996 -16 3036
rect 587 3036 604 3044
rect 416 3024 424 3033
rect 207 3016 453 3024
rect 556 3024 564 3033
rect 556 3016 573 3024
rect 596 3024 604 3036
rect 647 3036 713 3044
rect 1027 3036 1193 3044
rect 1347 3036 1504 3044
rect 596 3016 673 3024
rect 707 3016 993 3024
rect 1096 3016 1393 3024
rect 507 2996 513 3004
rect 527 2996 553 3004
rect 576 2996 593 3004
rect 576 2964 584 2996
rect 667 2996 793 3004
rect 1096 3004 1104 3016
rect 1496 3024 1504 3036
rect 1616 3036 1693 3044
rect 1616 3024 1624 3036
rect 1716 3036 1793 3044
rect 1496 3016 1624 3024
rect 1716 3024 1724 3036
rect 1647 3016 1724 3024
rect 1747 3016 1773 3024
rect 1836 3024 1844 3033
rect 1836 3016 1884 3024
rect 907 2996 1104 3004
rect 1367 2996 1393 3004
rect 1876 3004 1884 3016
rect 1936 3024 1944 3033
rect 1927 3016 1973 3024
rect 2027 3016 2053 3024
rect 2076 3007 2084 3076
rect 2387 3076 2553 3084
rect 2567 3076 2873 3084
rect 2887 3076 2944 3084
rect 2127 3056 2233 3064
rect 2287 3056 2293 3064
rect 2307 3056 2453 3064
rect 2467 3056 2724 3064
rect 1876 2996 1893 3004
rect 2096 3004 2104 3053
rect 2116 3036 2284 3044
rect 2116 3027 2124 3036
rect 2147 3016 2164 3024
rect 2096 2996 2133 3004
rect 2156 3004 2164 3016
rect 2187 3016 2213 3024
rect 2276 3024 2284 3036
rect 2367 3036 2473 3044
rect 2636 3036 2693 3044
rect 2276 3016 2413 3024
rect 2636 3024 2644 3036
rect 2716 3044 2724 3056
rect 2836 3056 2873 3064
rect 2836 3044 2844 3056
rect 2716 3036 2844 3044
rect 2867 3036 2884 3044
rect 2427 3016 2644 3024
rect 2667 3016 2853 3024
rect 2876 3007 2884 3036
rect 2896 3027 2904 3053
rect 2936 3027 2944 3076
rect 4456 3084 4464 3096
rect 4527 3096 4593 3104
rect 4647 3096 4793 3104
rect 4867 3096 4973 3104
rect 5007 3096 5113 3104
rect 5127 3096 5313 3104
rect 5327 3096 5853 3104
rect 5887 3096 6193 3104
rect 6227 3096 6493 3104
rect 3647 3076 4464 3084
rect 4487 3076 4573 3084
rect 4627 3076 4673 3084
rect 4747 3076 5393 3084
rect 5407 3076 6173 3084
rect 6187 3076 6233 3084
rect 6247 3076 6253 3084
rect 6267 3076 6473 3084
rect 6516 3076 6633 3084
rect 3387 3056 3464 3064
rect 2987 3036 3093 3044
rect 3116 3036 3133 3044
rect 3007 3016 3033 3024
rect 2156 2996 2193 3004
rect 2207 2996 2253 3004
rect 2627 2996 2793 3004
rect 2916 2996 3053 3004
rect 607 2976 673 2984
rect 687 2976 813 2984
rect 867 2976 1073 2984
rect 1347 2976 2213 2984
rect 2916 2984 2924 2996
rect 3076 2987 3084 3013
rect 3116 3007 3124 3036
rect 3167 3036 3244 3044
rect 3236 3027 3244 3036
rect 3267 3036 3353 3044
rect 3367 3036 3433 3044
rect 3456 3027 3464 3056
rect 3547 3056 3633 3064
rect 3787 3056 3884 3064
rect 3607 3036 3853 3044
rect 3147 3016 3193 3024
rect 3876 3024 3884 3056
rect 3907 3056 4273 3064
rect 4036 3047 4044 3056
rect 4307 3056 4493 3064
rect 4507 3056 4673 3064
rect 4687 3056 4713 3064
rect 4867 3056 4913 3064
rect 4987 3056 5004 3064
rect 4127 3036 4353 3044
rect 4776 3036 4813 3044
rect 3827 3016 3973 3024
rect 4227 3016 4233 3024
rect 4616 3024 4624 3033
rect 4256 3016 4344 3024
rect 4616 3016 4653 3024
rect 3287 2996 3333 3004
rect 3607 2996 4073 3004
rect 4167 2996 4193 3004
rect 2787 2976 2924 2984
rect 2947 2976 3013 2984
rect 3107 2976 3153 2984
rect 3167 2976 3313 2984
rect 3576 2984 3584 2993
rect 3547 2976 3584 2984
rect 3627 2976 3773 2984
rect 4216 2984 4224 3013
rect 4256 3004 4264 3016
rect 4336 3007 4344 3016
rect 4776 3007 4784 3036
rect 4907 3036 4984 3044
rect 4976 3027 4984 3036
rect 4847 3016 4953 3024
rect 4996 3024 5004 3056
rect 5027 3056 5193 3064
rect 5327 3056 5424 3064
rect 5287 3036 5373 3044
rect 5416 3044 5424 3056
rect 5547 3056 5573 3064
rect 5616 3056 5653 3064
rect 5416 3036 5453 3044
rect 4996 3016 5253 3024
rect 4247 2996 4264 3004
rect 4427 2996 4633 3004
rect 4667 2996 4693 3004
rect 4727 2996 4764 3004
rect 3827 2976 4273 2984
rect 4567 2976 4733 2984
rect 4756 2984 4764 2996
rect 4807 2996 4844 3004
rect 4756 2976 4813 2984
rect 4836 2984 4844 2996
rect 4996 3004 5004 3016
rect 5376 3024 5384 3033
rect 5376 3016 5533 3024
rect 5616 3024 5624 3056
rect 5767 3056 5804 3064
rect 5796 3044 5804 3056
rect 5867 3056 5973 3064
rect 6187 3056 6213 3064
rect 6396 3056 6493 3064
rect 5647 3036 5744 3044
rect 5796 3036 5933 3044
rect 5547 3016 5624 3024
rect 5736 3024 5744 3036
rect 5947 3036 6033 3044
rect 6116 3027 6124 3053
rect 5736 3016 5764 3024
rect 4967 2996 5004 3004
rect 5047 2996 5153 3004
rect 5287 2996 5593 3004
rect 5756 3004 5764 3016
rect 5927 3016 5993 3024
rect 6167 3016 6273 3024
rect 6336 3024 6344 3033
rect 6356 3027 6364 3053
rect 6287 3016 6344 3024
rect 5756 2996 5793 3004
rect 6187 2996 6213 3004
rect 6376 3004 6384 3033
rect 6396 3027 6404 3056
rect 6516 3044 6524 3076
rect 6496 3036 6524 3044
rect 6416 3024 6424 3033
rect 6496 3027 6504 3036
rect 6416 3016 6453 3024
rect 6527 3016 6573 3024
rect 6347 2996 6384 3004
rect 6596 3004 6604 3053
rect 6587 2996 6604 3004
rect 4836 2976 5153 2984
rect 5187 2976 5313 2984
rect 5427 2976 5484 2984
rect 576 2956 613 2964
rect 707 2956 753 2964
rect 887 2956 953 2964
rect 2087 2956 2144 2964
rect 307 2936 853 2944
rect 2136 2944 2144 2956
rect 2167 2956 2193 2964
rect 3067 2956 3213 2964
rect 3307 2956 3613 2964
rect 3627 2956 3993 2964
rect 4127 2956 4533 2964
rect 4987 2956 5453 2964
rect 5476 2964 5484 2976
rect 5527 2976 5853 2984
rect 6307 2976 6633 2984
rect 5476 2956 5913 2964
rect 2136 2936 2253 2944
rect 3207 2936 3313 2944
rect 3347 2936 3393 2944
rect 3407 2936 3633 2944
rect 3727 2936 4833 2944
rect 5487 2936 5593 2944
rect 5647 2936 5693 2944
rect 5727 2936 6373 2944
rect 1787 2916 3053 2924
rect 4527 2916 4913 2924
rect 4947 2916 4993 2924
rect 5247 2916 5493 2924
rect 2327 2896 3653 2904
rect 4187 2896 4493 2904
rect 4907 2896 5053 2904
rect 2827 2876 3073 2884
rect 3087 2876 3753 2884
rect 4607 2876 4713 2884
rect 4787 2876 5713 2884
rect 2347 2856 2493 2864
rect 2727 2856 2893 2864
rect 2927 2856 3004 2864
rect 1007 2836 2973 2844
rect 2996 2844 3004 2856
rect 3027 2856 3113 2864
rect 3127 2856 3573 2864
rect 3587 2856 4173 2864
rect 4707 2856 4964 2864
rect 2996 2836 3313 2844
rect 3336 2836 3553 2844
rect 627 2816 813 2824
rect 1227 2816 1373 2824
rect 2187 2816 2913 2824
rect 3047 2816 3053 2824
rect 3336 2824 3344 2836
rect 4027 2836 4553 2844
rect 4956 2844 4964 2856
rect 5107 2856 5973 2864
rect 4956 2836 5013 2844
rect 5027 2836 5213 2844
rect 5236 2836 5513 2844
rect 3067 2816 3344 2824
rect 3356 2816 3813 2824
rect 767 2796 793 2804
rect 827 2796 853 2804
rect 867 2796 933 2804
rect 967 2796 1053 2804
rect 1107 2796 1613 2804
rect 1627 2796 1673 2804
rect 2067 2796 2233 2804
rect 2387 2796 2413 2804
rect 3007 2796 3133 2804
rect 3356 2804 3364 2816
rect 4007 2816 4413 2824
rect 4447 2816 4513 2824
rect 4847 2816 4933 2824
rect 5236 2824 5244 2836
rect 5527 2836 5933 2844
rect 5947 2836 5953 2844
rect 6067 2836 6273 2844
rect 5167 2816 5244 2824
rect 5467 2816 5604 2824
rect 3147 2796 3364 2804
rect 3427 2796 3553 2804
rect 3807 2796 3993 2804
rect 4087 2796 4124 2804
rect 567 2776 593 2784
rect 607 2776 893 2784
rect 987 2776 1024 2784
rect 47 2756 104 2764
rect 96 2747 104 2756
rect 456 2756 524 2764
rect 116 2736 233 2744
rect 116 2727 124 2736
rect 456 2744 464 2756
rect 516 2747 524 2756
rect 747 2756 844 2764
rect 836 2747 844 2756
rect 1016 2747 1024 2776
rect 1156 2776 1313 2784
rect 1047 2756 1093 2764
rect 1127 2756 1144 2764
rect 376 2736 464 2744
rect 376 2724 384 2736
rect 847 2736 913 2744
rect 1027 2736 1073 2744
rect 147 2716 384 2724
rect 467 2716 653 2724
rect 1136 2724 1144 2756
rect 1156 2747 1164 2776
rect 1456 2776 1593 2784
rect 1456 2767 1464 2776
rect 1667 2776 1753 2784
rect 1767 2776 1853 2784
rect 1907 2776 1933 2784
rect 2007 2776 2273 2784
rect 2527 2776 2873 2784
rect 2916 2776 2933 2784
rect 1216 2756 1273 2764
rect 1176 2724 1184 2753
rect 1216 2744 1224 2756
rect 1367 2756 1393 2764
rect 1507 2756 1544 2764
rect 1207 2736 1224 2744
rect 1247 2736 1293 2744
rect 1336 2744 1344 2753
rect 1536 2747 1544 2756
rect 1847 2756 1913 2764
rect 2087 2756 2113 2764
rect 2167 2756 2433 2764
rect 2456 2764 2464 2773
rect 2456 2756 2573 2764
rect 2796 2756 2873 2764
rect 1316 2736 1344 2744
rect 1136 2716 1184 2724
rect 1316 2724 1324 2736
rect 1387 2736 1473 2744
rect 1556 2727 1564 2753
rect 1607 2736 1813 2744
rect 1867 2736 1893 2744
rect 2067 2736 2093 2744
rect 2136 2744 2144 2753
rect 2116 2736 2193 2744
rect 1207 2716 1324 2724
rect 1427 2716 1453 2724
rect 1507 2716 1533 2724
rect 1567 2716 1593 2724
rect 1727 2716 1853 2724
rect 2116 2724 2124 2736
rect 2207 2736 2244 2744
rect 2056 2716 2124 2724
rect 2236 2724 2244 2736
rect 2236 2716 2293 2724
rect 167 2696 1133 2704
rect 1147 2696 1713 2704
rect 2056 2704 2064 2716
rect 1727 2696 2064 2704
rect 2087 2696 2133 2704
rect 2307 2696 2533 2704
rect 2547 2696 2733 2704
rect 2747 2696 2753 2704
rect 2796 2704 2804 2756
rect 2896 2747 2904 2773
rect 2916 2767 2924 2776
rect 2967 2776 3073 2784
rect 3087 2776 3253 2784
rect 3807 2776 3853 2784
rect 3876 2776 3973 2784
rect 3327 2756 3364 2764
rect 2827 2736 2844 2744
rect 2836 2724 2844 2736
rect 2867 2736 2884 2744
rect 2876 2727 2884 2736
rect 2927 2736 2953 2744
rect 3016 2736 3213 2744
rect 3016 2727 3024 2736
rect 3296 2744 3304 2753
rect 3356 2747 3364 2756
rect 3427 2756 3453 2764
rect 3876 2764 3884 2776
rect 4027 2776 4064 2784
rect 3856 2756 3884 2764
rect 3896 2756 3933 2764
rect 3267 2736 3284 2744
rect 3296 2736 3324 2744
rect 2836 2716 2853 2724
rect 3276 2724 3284 2736
rect 3316 2727 3324 2736
rect 3587 2736 3664 2744
rect 3276 2716 3293 2724
rect 3367 2716 3573 2724
rect 3656 2724 3664 2736
rect 3836 2744 3844 2753
rect 3747 2736 3844 2744
rect 3656 2716 3673 2724
rect 3727 2716 3833 2724
rect 3856 2724 3864 2756
rect 3896 2747 3904 2756
rect 4007 2756 4044 2764
rect 3956 2744 3964 2753
rect 3927 2736 3964 2744
rect 3847 2716 3864 2724
rect 4036 2724 4044 2756
rect 4007 2716 4044 2724
rect 2796 2696 2893 2704
rect 3207 2696 3373 2704
rect 3407 2696 3433 2704
rect 3467 2696 3513 2704
rect 3567 2696 3613 2704
rect 3667 2696 3733 2704
rect 3767 2696 3913 2704
rect 4056 2704 4064 2776
rect 4076 2727 4084 2753
rect 4096 2744 4104 2773
rect 4116 2764 4124 2796
rect 4187 2796 4304 2804
rect 4147 2776 4253 2784
rect 4116 2756 4213 2764
rect 4096 2736 4153 2744
rect 4216 2727 4224 2753
rect 4296 2747 4304 2796
rect 4927 2796 5233 2804
rect 5267 2796 5493 2804
rect 5547 2796 5573 2804
rect 5596 2804 5604 2816
rect 5796 2816 5853 2824
rect 5796 2804 5804 2816
rect 6167 2816 6333 2824
rect 5596 2796 5804 2804
rect 5827 2796 5873 2804
rect 6027 2796 6093 2804
rect 6307 2796 6393 2804
rect 4327 2776 4353 2784
rect 4527 2776 4573 2784
rect 4976 2776 5033 2784
rect 4347 2756 4393 2764
rect 4816 2764 4824 2773
rect 4936 2764 4944 2773
rect 4427 2756 4524 2764
rect 4367 2736 4393 2744
rect 4516 2744 4524 2756
rect 4776 2756 4824 2764
rect 4916 2756 4944 2764
rect 4516 2736 4633 2744
rect 4776 2744 4784 2756
rect 4647 2736 4704 2744
rect 4127 2716 4173 2724
rect 4267 2716 4333 2724
rect 4347 2716 4373 2724
rect 4447 2716 4673 2724
rect 4696 2724 4704 2736
rect 4756 2736 4784 2744
rect 4696 2716 4733 2724
rect 4756 2724 4764 2736
rect 4916 2744 4924 2756
rect 4976 2747 4984 2776
rect 5127 2776 5233 2784
rect 5407 2776 5433 2784
rect 5567 2776 5713 2784
rect 5727 2776 6173 2784
rect 5056 2764 5064 2773
rect 5047 2756 5064 2764
rect 5367 2756 5473 2764
rect 5647 2756 5813 2764
rect 6007 2756 6084 2764
rect 4887 2736 4924 2744
rect 5036 2736 5053 2744
rect 4747 2716 4764 2724
rect 4827 2716 4913 2724
rect 5016 2724 5024 2733
rect 5036 2727 5044 2736
rect 5136 2744 5144 2753
rect 5107 2736 5144 2744
rect 4967 2716 5024 2724
rect 5156 2724 5164 2753
rect 5087 2716 5164 2724
rect 5187 2716 5273 2724
rect 5316 2724 5324 2753
rect 5356 2727 5364 2753
rect 6076 2747 6084 2756
rect 6127 2756 6164 2764
rect 5476 2736 5493 2744
rect 5476 2727 5484 2736
rect 6027 2736 6044 2744
rect 5316 2716 5333 2724
rect 5776 2724 5784 2733
rect 5567 2716 5833 2724
rect 5847 2716 5953 2724
rect 5987 2716 6013 2724
rect 6036 2724 6044 2736
rect 6107 2736 6133 2744
rect 6036 2716 6053 2724
rect 6156 2724 6164 2756
rect 6187 2736 6553 2744
rect 6567 2736 6573 2744
rect 6107 2716 6164 2724
rect 6267 2716 6353 2724
rect 6527 2716 6573 2724
rect 3967 2696 4064 2704
rect 4216 2696 4393 2704
rect 507 2676 613 2684
rect 1167 2676 2113 2684
rect 2967 2676 3053 2684
rect 3227 2676 3413 2684
rect 4216 2684 4224 2696
rect 4447 2696 4493 2704
rect 4547 2696 4813 2704
rect 4827 2696 4833 2704
rect 4927 2696 5233 2704
rect 5447 2696 5653 2704
rect 5687 2696 5893 2704
rect 5927 2696 6293 2704
rect 6307 2696 6453 2704
rect 6467 2696 6513 2704
rect 3607 2676 4224 2684
rect 4287 2676 4513 2684
rect 4867 2676 4893 2684
rect 4987 2676 5173 2684
rect 5387 2676 5433 2684
rect 5487 2676 5573 2684
rect 5667 2676 5793 2684
rect 5867 2676 6073 2684
rect 1347 2656 1593 2664
rect 1667 2656 2033 2664
rect 2287 2656 2413 2664
rect 2427 2656 3073 2664
rect 3096 2656 3213 2664
rect 67 2636 253 2644
rect 267 2636 973 2644
rect 1587 2636 1633 2644
rect 1647 2636 1793 2644
rect 1807 2636 1833 2644
rect 1947 2636 2173 2644
rect 2387 2636 2753 2644
rect 2807 2636 2873 2644
rect 2907 2636 2973 2644
rect 3096 2644 3104 2656
rect 3247 2656 4093 2664
rect 4107 2656 4353 2664
rect 4367 2656 4404 2664
rect 3007 2636 3104 2644
rect 3196 2636 3373 2644
rect 1547 2616 1613 2624
rect 1687 2616 1993 2624
rect 2047 2616 2773 2624
rect 3196 2624 3204 2636
rect 3396 2636 3813 2644
rect 2827 2616 3204 2624
rect 3396 2624 3404 2636
rect 4067 2636 4133 2644
rect 4207 2636 4353 2644
rect 4396 2644 4404 2656
rect 4427 2656 4913 2664
rect 5047 2656 5193 2664
rect 5407 2656 5473 2664
rect 5887 2656 6053 2664
rect 6507 2656 6693 2664
rect 4396 2636 4464 2644
rect 3227 2616 3404 2624
rect 3427 2616 3473 2624
rect 3707 2616 4104 2624
rect 127 2596 273 2604
rect 647 2596 833 2604
rect 847 2596 953 2604
rect 1007 2596 1233 2604
rect 1387 2596 1493 2604
rect 1907 2596 2173 2604
rect 2187 2596 2293 2604
rect 2347 2596 2484 2604
rect 136 2576 153 2584
rect 136 2544 144 2576
rect 287 2576 433 2584
rect 1047 2576 1133 2584
rect 1527 2576 1553 2584
rect 327 2556 353 2564
rect 487 2556 593 2564
rect 1027 2556 1053 2564
rect 1187 2556 1273 2564
rect 1296 2556 1353 2564
rect 136 2536 164 2544
rect 156 2527 164 2536
rect 667 2536 693 2544
rect 707 2536 784 2544
rect 776 2527 784 2536
rect 1296 2544 1304 2556
rect 1436 2564 1444 2573
rect 1436 2556 1513 2564
rect 807 2536 1304 2544
rect -24 2504 -16 2524
rect 367 2516 673 2524
rect 867 2516 993 2524
rect 1007 2516 1033 2524
rect 1296 2524 1304 2536
rect 1436 2544 1444 2556
rect 1327 2536 1444 2544
rect 1536 2544 1544 2576
rect 1827 2576 1893 2584
rect 1916 2576 1973 2584
rect 1916 2564 1924 2576
rect 2087 2576 2253 2584
rect 2267 2576 2373 2584
rect 2476 2584 2484 2596
rect 2507 2596 2533 2604
rect 2567 2596 2653 2604
rect 2767 2596 2813 2604
rect 2907 2596 3113 2604
rect 3147 2596 3593 2604
rect 3647 2596 3773 2604
rect 3947 2596 4073 2604
rect 4096 2604 4104 2616
rect 4247 2616 4373 2624
rect 4456 2624 4464 2636
rect 4747 2636 4793 2644
rect 4887 2636 5113 2644
rect 5267 2636 5413 2644
rect 5427 2636 5513 2644
rect 5767 2636 5813 2644
rect 5847 2636 5973 2644
rect 6167 2636 6193 2644
rect 4456 2616 4513 2624
rect 4567 2616 4744 2624
rect 4736 2607 4744 2616
rect 4767 2616 5053 2624
rect 5067 2616 5573 2624
rect 5787 2616 5913 2624
rect 5967 2616 5993 2624
rect 6107 2616 6333 2624
rect 6387 2616 6693 2624
rect 4096 2596 4193 2604
rect 4227 2596 4293 2604
rect 4307 2596 4413 2604
rect 4496 2596 4553 2604
rect 2476 2576 2753 2584
rect 1896 2556 1924 2564
rect 1936 2556 1953 2564
rect 1467 2536 1544 2544
rect 1767 2536 1813 2544
rect 1896 2544 1904 2556
rect 1827 2536 1904 2544
rect 1936 2544 1944 2556
rect 2016 2547 2024 2573
rect 2596 2567 2604 2576
rect 2787 2576 2993 2584
rect 3047 2576 3104 2584
rect 2247 2556 2353 2564
rect 2727 2556 2744 2564
rect 1927 2536 1944 2544
rect 2107 2536 2133 2544
rect 2347 2536 2553 2544
rect 2736 2544 2744 2556
rect 2787 2556 2833 2564
rect 3096 2564 3104 2576
rect 3396 2576 3533 2584
rect 3096 2556 3213 2564
rect 2607 2536 2724 2544
rect 2736 2536 2873 2544
rect 1296 2516 1333 2524
rect 1507 2516 1553 2524
rect 2227 2516 2313 2524
rect 2487 2516 2693 2524
rect 2716 2524 2724 2536
rect 2716 2516 2773 2524
rect 2796 2516 2953 2524
rect -24 2496 293 2504
rect 567 2496 713 2504
rect 1307 2496 1413 2504
rect 1987 2496 2053 2504
rect 2067 2496 2613 2504
rect 2796 2504 2804 2516
rect 2707 2496 2804 2504
rect 2976 2504 2984 2553
rect 3056 2544 3064 2553
rect 3396 2547 3404 2576
rect 3556 2576 3593 2584
rect 3556 2564 3564 2576
rect 3687 2576 3993 2584
rect 4147 2576 4193 2584
rect 4267 2576 4344 2584
rect 3467 2556 3564 2564
rect 3587 2556 3613 2564
rect 3687 2556 3813 2564
rect 4016 2564 4024 2573
rect 3907 2556 4024 2564
rect 4016 2547 4024 2556
rect 4036 2547 4044 2573
rect 4336 2564 4344 2576
rect 4496 2567 4504 2596
rect 4907 2596 5073 2604
rect 5287 2596 5373 2604
rect 5587 2596 6033 2604
rect 4656 2576 4673 2584
rect 4287 2556 4324 2564
rect 4336 2556 4464 2564
rect 3056 2536 3093 2544
rect 3447 2536 3493 2544
rect 3567 2536 3633 2544
rect 3656 2536 3673 2544
rect 3087 2516 3533 2524
rect 3656 2524 3664 2536
rect 3707 2536 3793 2544
rect 4056 2536 4293 2544
rect 3567 2516 3664 2524
rect 3687 2516 3713 2524
rect 3807 2516 3853 2524
rect 3876 2524 3884 2533
rect 3876 2516 3893 2524
rect 4056 2524 4064 2536
rect 4316 2544 4324 2556
rect 4456 2544 4464 2556
rect 4656 2564 4664 2576
rect 4936 2576 5033 2584
rect 4936 2567 4944 2576
rect 5116 2576 5224 2584
rect 4636 2556 4664 2564
rect 4316 2536 4444 2544
rect 4456 2536 4573 2544
rect 4007 2516 4064 2524
rect 4107 2516 4413 2524
rect 4436 2524 4444 2536
rect 4436 2516 4553 2524
rect 4616 2524 4624 2553
rect 4636 2547 4644 2556
rect 5116 2564 5124 2576
rect 4967 2556 5124 2564
rect 5216 2564 5224 2576
rect 5247 2576 5293 2584
rect 5327 2576 5353 2584
rect 5367 2576 5384 2584
rect 5216 2556 5253 2564
rect 5136 2544 5144 2553
rect 5376 2547 5384 2576
rect 5567 2576 5733 2584
rect 6007 2576 6044 2584
rect 5507 2556 5773 2564
rect 5107 2536 5144 2544
rect 5207 2536 5233 2544
rect 5287 2536 5333 2544
rect 5547 2536 5653 2544
rect 5687 2536 5713 2544
rect 5816 2544 5824 2573
rect 5916 2544 5924 2553
rect 5976 2544 5984 2573
rect 6036 2564 6044 2576
rect 6067 2576 6104 2584
rect 6096 2567 6104 2576
rect 6427 2576 6444 2584
rect 6036 2556 6084 2564
rect 5816 2536 5844 2544
rect 5916 2536 5984 2544
rect 5996 2544 6004 2553
rect 5996 2536 6033 2544
rect 5836 2527 5844 2536
rect 6076 2544 6084 2556
rect 6176 2556 6213 2564
rect 6176 2544 6184 2556
rect 6076 2536 6184 2544
rect 6416 2544 6424 2553
rect 6436 2547 6444 2576
rect 6536 2564 6544 2573
rect 6516 2556 6573 2564
rect 6207 2536 6424 2544
rect 6516 2544 6524 2556
rect 6667 2556 6693 2564
rect 6487 2536 6524 2544
rect 6547 2536 6593 2544
rect 4567 2516 4624 2524
rect 4787 2516 4853 2524
rect 5507 2516 5593 2524
rect 6507 2516 6573 2524
rect 2967 2496 2984 2504
rect 3467 2496 3493 2504
rect 3527 2496 3793 2504
rect 3967 2496 4113 2504
rect 4247 2496 4493 2504
rect 4567 2496 4673 2504
rect 5167 2496 5193 2504
rect 5356 2496 5913 2504
rect 1467 2476 1933 2484
rect 2287 2476 2704 2484
rect 987 2456 2673 2464
rect 2696 2464 2704 2476
rect 2847 2476 3113 2484
rect 3127 2476 3233 2484
rect 3387 2476 3453 2484
rect 3487 2476 3673 2484
rect 3727 2476 3773 2484
rect 3827 2476 4004 2484
rect 2696 2456 2793 2464
rect 2807 2456 2933 2464
rect 3996 2464 4004 2476
rect 4027 2476 4253 2484
rect 4407 2476 4804 2484
rect 2947 2456 3424 2464
rect 3996 2456 4053 2464
rect 1747 2436 2253 2444
rect 2267 2436 2313 2444
rect 2367 2436 2553 2444
rect 2627 2436 3033 2444
rect 3107 2436 3173 2444
rect 3416 2444 3424 2456
rect 4087 2456 4213 2464
rect 4796 2464 4804 2476
rect 5356 2484 5364 2496
rect 5967 2496 6073 2504
rect 4827 2476 5364 2484
rect 5847 2476 5933 2484
rect 4267 2456 4564 2464
rect 4796 2456 5293 2464
rect 3416 2436 3973 2444
rect 4556 2444 4564 2456
rect 5787 2456 6413 2464
rect 4147 2436 4324 2444
rect 4556 2436 4953 2444
rect 1447 2416 2373 2424
rect 2467 2416 2573 2424
rect 2627 2416 2713 2424
rect 2736 2416 2893 2424
rect 1647 2396 1913 2404
rect 2227 2396 2593 2404
rect 2736 2404 2744 2416
rect 2907 2416 3333 2424
rect 3407 2416 3473 2424
rect 3507 2416 3604 2424
rect 2707 2396 2744 2404
rect 2987 2396 3573 2404
rect 3596 2404 3604 2416
rect 3787 2416 4073 2424
rect 4167 2416 4293 2424
rect 4316 2424 4324 2436
rect 4987 2436 5033 2444
rect 5047 2436 5064 2444
rect 4316 2416 4433 2424
rect 4587 2416 5033 2424
rect 5056 2424 5064 2436
rect 5207 2436 5373 2444
rect 5747 2436 5873 2444
rect 5887 2436 5973 2444
rect 6027 2436 6113 2444
rect 6307 2436 6653 2444
rect 5056 2416 5673 2424
rect 5807 2416 6433 2424
rect 3596 2396 3833 2404
rect 3867 2396 3893 2404
rect 4067 2396 4673 2404
rect 5407 2396 5713 2404
rect 6407 2396 6433 2404
rect 1187 2376 1253 2384
rect 1907 2376 2233 2384
rect 2276 2376 2653 2384
rect 2276 2364 2284 2376
rect 3007 2376 3153 2384
rect 3187 2376 3293 2384
rect 3307 2376 3553 2384
rect 3607 2376 4013 2384
rect 4187 2376 4233 2384
rect 4327 2376 4393 2384
rect 4427 2376 4753 2384
rect 5007 2376 5613 2384
rect 5647 2376 5833 2384
rect 2067 2356 2284 2364
rect 2307 2356 2864 2364
rect 387 2336 613 2344
rect 767 2336 784 2344
rect 307 2296 373 2304
rect 427 2296 513 2304
rect 776 2304 784 2336
rect 1047 2336 2533 2344
rect 2567 2336 2833 2344
rect 2856 2344 2864 2356
rect 2887 2356 3133 2364
rect 4207 2356 4353 2364
rect 4547 2356 4593 2364
rect 4787 2356 4893 2364
rect 5127 2356 5153 2364
rect 5167 2356 5253 2364
rect 5327 2356 5433 2364
rect 5787 2356 5813 2364
rect 5836 2356 6293 2364
rect 2856 2336 2873 2344
rect 2947 2336 3213 2344
rect 3236 2336 3473 2344
rect 1547 2316 1613 2324
rect 1627 2316 1653 2324
rect 2407 2316 2544 2324
rect 536 2296 644 2304
rect 96 2276 233 2284
rect 96 2267 104 2276
rect 536 2284 544 2296
rect 427 2276 484 2284
rect 476 2267 484 2276
rect 496 2276 544 2284
rect 556 2276 613 2284
rect 216 2227 224 2253
rect 496 2247 504 2276
rect 527 2256 533 2264
rect 556 2264 564 2276
rect 636 2284 644 2296
rect 696 2296 784 2304
rect 696 2284 704 2296
rect 776 2287 784 2296
rect 807 2296 864 2304
rect 636 2276 704 2284
rect 547 2256 564 2264
rect 747 2256 813 2264
rect 827 2256 833 2264
rect 247 2236 473 2244
rect 527 2236 653 2244
rect 727 2236 813 2244
rect 856 2244 864 2296
rect 1327 2296 1564 2304
rect 1007 2276 1164 2284
rect 1156 2264 1164 2276
rect 1487 2276 1524 2284
rect 1516 2267 1524 2276
rect 1556 2267 1564 2296
rect 1667 2296 1713 2304
rect 1727 2296 2413 2304
rect 2456 2296 2513 2304
rect 1156 2256 1284 2264
rect 827 2236 864 2244
rect 1276 2244 1284 2256
rect 1276 2236 1333 2244
rect 1447 2236 1493 2244
rect 1576 2244 1584 2273
rect 1636 2264 1644 2293
rect 1707 2276 1973 2284
rect 2087 2276 2273 2284
rect 2287 2276 2353 2284
rect 1636 2256 1673 2264
rect 1747 2256 1793 2264
rect 1887 2256 1984 2264
rect 1576 2236 1773 2244
rect 1867 2236 1913 2244
rect 1976 2244 1984 2256
rect 2036 2264 2044 2273
rect 2007 2256 2044 2264
rect 2056 2244 2064 2273
rect 2167 2256 2233 2264
rect 2336 2256 2373 2264
rect 1976 2236 2173 2244
rect 2336 2244 2344 2256
rect 2187 2236 2344 2244
rect 2367 2236 2393 2244
rect 2416 2244 2424 2273
rect 2436 2267 2444 2293
rect 2456 2287 2464 2296
rect 2536 2264 2544 2316
rect 2556 2316 2573 2324
rect 2556 2307 2564 2316
rect 2667 2316 2764 2324
rect 2667 2296 2693 2304
rect 2756 2304 2764 2316
rect 3236 2324 3244 2336
rect 3567 2336 3933 2344
rect 3947 2336 4513 2344
rect 4727 2336 4733 2344
rect 4747 2336 4933 2344
rect 4947 2336 5413 2344
rect 5447 2336 5653 2344
rect 5836 2344 5844 2356
rect 6347 2356 6393 2364
rect 5667 2336 5844 2344
rect 5856 2336 6153 2344
rect 2787 2316 3244 2324
rect 3327 2316 3633 2324
rect 4996 2316 5153 2324
rect 2756 2296 2804 2304
rect 2636 2284 2644 2293
rect 2567 2276 2644 2284
rect 2796 2284 2804 2296
rect 2907 2296 2973 2304
rect 3027 2296 3044 2304
rect 2687 2276 2764 2284
rect 2796 2276 2864 2284
rect 2756 2267 2764 2276
rect 2856 2267 2864 2276
rect 2876 2276 2924 2284
rect 2467 2256 2544 2264
rect 2567 2256 2693 2264
rect 2416 2236 2613 2244
rect 2667 2236 2693 2244
rect 2876 2244 2884 2276
rect 2916 2264 2924 2276
rect 2947 2276 3024 2284
rect 3016 2267 3024 2276
rect 2916 2256 3004 2264
rect 2816 2236 2884 2244
rect 2896 2244 2904 2253
rect 2896 2236 2933 2244
rect 247 2216 553 2224
rect 567 2216 753 2224
rect 767 2216 973 2224
rect 1547 2216 1793 2224
rect 1807 2216 1953 2224
rect 2287 2216 2693 2224
rect 2816 2224 2824 2236
rect 2996 2244 3004 2256
rect 3036 2244 3044 2296
rect 3367 2296 3524 2304
rect 3076 2284 3084 2293
rect 3076 2276 3173 2284
rect 3207 2276 3253 2284
rect 3316 2276 3373 2284
rect 3316 2267 3324 2276
rect 3396 2276 3473 2284
rect 3167 2256 3233 2264
rect 3396 2264 3404 2276
rect 3516 2284 3524 2296
rect 3547 2296 3773 2304
rect 3847 2296 3893 2304
rect 4016 2296 4033 2304
rect 3516 2276 3653 2284
rect 3796 2284 3804 2293
rect 3667 2276 3804 2284
rect 3367 2256 3404 2264
rect 3427 2256 3493 2264
rect 3827 2256 3873 2264
rect 3887 2256 3893 2264
rect 3947 2256 3993 2264
rect 4016 2264 4024 2296
rect 4127 2296 4224 2304
rect 4047 2276 4084 2284
rect 4076 2264 4084 2276
rect 4016 2256 4064 2264
rect 4076 2256 4113 2264
rect 2996 2236 3044 2244
rect 3056 2236 3413 2244
rect 2747 2216 2824 2224
rect 2847 2216 2953 2224
rect 3056 2224 3064 2236
rect 3756 2244 3764 2253
rect 3467 2236 3953 2244
rect 3967 2236 3973 2244
rect 4056 2244 4064 2256
rect 4216 2264 4224 2296
rect 4247 2296 4273 2304
rect 4996 2304 5004 2316
rect 5187 2316 5204 2324
rect 4796 2296 5004 2304
rect 4416 2276 4493 2284
rect 4216 2256 4293 2264
rect 4347 2256 4364 2264
rect 4056 2236 4173 2244
rect 4267 2236 4333 2244
rect 4356 2244 4364 2256
rect 4416 2264 4424 2276
rect 4667 2276 4724 2284
rect 4387 2256 4424 2264
rect 4716 2264 4724 2276
rect 4547 2256 4684 2264
rect 4716 2256 4753 2264
rect 4356 2236 4493 2244
rect 4507 2236 4593 2244
rect 4676 2244 4684 2256
rect 4796 2244 4804 2296
rect 5027 2296 5064 2304
rect 4816 2276 4873 2284
rect 4816 2267 4824 2276
rect 5056 2284 5064 2296
rect 5196 2284 5204 2316
rect 5287 2316 5373 2324
rect 5716 2316 5733 2324
rect 5307 2296 5324 2304
rect 5316 2284 5324 2296
rect 5427 2296 5453 2304
rect 5716 2304 5724 2316
rect 5836 2304 5844 2313
rect 5856 2307 5864 2336
rect 6387 2336 6453 2344
rect 6487 2336 6593 2344
rect 5876 2316 5933 2324
rect 5627 2296 5664 2304
rect 5056 2276 5084 2284
rect 5196 2276 5224 2284
rect 5316 2276 5424 2284
rect 5076 2267 5084 2276
rect 5216 2267 5224 2276
rect 5416 2267 5424 2276
rect 5527 2276 5604 2284
rect 5436 2264 5444 2273
rect 5596 2267 5604 2276
rect 5656 2267 5664 2296
rect 5696 2296 5724 2304
rect 5736 2296 5844 2304
rect 5436 2256 5524 2264
rect 4676 2236 4804 2244
rect 5516 2244 5524 2256
rect 5516 2236 5573 2244
rect 5696 2244 5704 2296
rect 5736 2284 5744 2296
rect 5876 2287 5884 2316
rect 5947 2316 6313 2324
rect 6327 2316 6473 2324
rect 6687 2316 6713 2324
rect 5927 2296 5984 2304
rect 5716 2276 5744 2284
rect 5716 2267 5724 2276
rect 5767 2276 5793 2284
rect 5807 2276 5833 2284
rect 5896 2276 5913 2284
rect 5896 2264 5904 2276
rect 5747 2256 5904 2264
rect 5936 2247 5944 2273
rect 5976 2267 5984 2296
rect 6467 2296 6513 2304
rect 6607 2296 6713 2304
rect 6087 2276 6173 2284
rect 6376 2284 6384 2293
rect 6367 2276 6384 2284
rect 6036 2264 6044 2273
rect 6016 2256 6044 2264
rect 6076 2256 6093 2264
rect 5667 2236 5704 2244
rect 5787 2236 5804 2244
rect 3047 2216 3064 2224
rect 3287 2216 3633 2224
rect 3927 2216 4013 2224
rect 4027 2216 4093 2224
rect 4147 2216 4373 2224
rect 4407 2216 4704 2224
rect 1607 2196 1653 2204
rect 1707 2196 1833 2204
rect 2347 2196 2513 2204
rect 2787 2196 3113 2204
rect 3207 2196 3573 2204
rect 3647 2196 3713 2204
rect 3787 2196 3893 2204
rect 3987 2196 4033 2204
rect 4067 2196 4253 2204
rect 4376 2196 4553 2204
rect 67 2176 173 2184
rect 607 2176 693 2184
rect 707 2176 853 2184
rect 867 2176 1153 2184
rect 1287 2176 1693 2184
rect 1767 2176 1804 2184
rect 587 2156 713 2164
rect 1527 2156 1773 2164
rect 1796 2164 1804 2176
rect 1847 2176 2153 2184
rect 2407 2176 2473 2184
rect 2887 2176 3164 2184
rect 1796 2156 1913 2164
rect 1947 2156 2053 2164
rect 2247 2156 2433 2164
rect 2527 2156 2653 2164
rect 2667 2156 3093 2164
rect 3107 2156 3133 2164
rect 3156 2164 3164 2176
rect 3187 2176 3353 2184
rect 3636 2176 3764 2184
rect 3156 2156 3373 2164
rect 3507 2156 3533 2164
rect 3636 2164 3644 2176
rect 3547 2156 3644 2164
rect 3756 2164 3764 2176
rect 3787 2176 3993 2184
rect 4027 2176 4233 2184
rect 4376 2184 4384 2196
rect 4696 2204 4704 2216
rect 4727 2216 4973 2224
rect 5027 2216 5053 2224
rect 5107 2216 5273 2224
rect 5447 2216 5533 2224
rect 5547 2216 5753 2224
rect 5796 2224 5804 2236
rect 5887 2236 5913 2244
rect 6016 2244 6024 2256
rect 5987 2236 6024 2244
rect 6076 2244 6084 2256
rect 6136 2256 6153 2264
rect 6047 2236 6084 2244
rect 6136 2244 6144 2256
rect 6236 2247 6244 2273
rect 6316 2264 6324 2273
rect 6316 2256 6373 2264
rect 6416 2264 6424 2293
rect 6447 2276 6493 2284
rect 6667 2276 6684 2284
rect 6416 2256 6433 2264
rect 6556 2264 6564 2273
rect 6516 2256 6564 2264
rect 6107 2236 6144 2244
rect 6267 2236 6273 2244
rect 6287 2236 6313 2244
rect 6347 2236 6373 2244
rect 6516 2244 6524 2256
rect 6427 2236 6524 2244
rect 6576 2244 6584 2273
rect 6676 2247 6684 2276
rect 6547 2236 6584 2244
rect 5796 2216 5853 2224
rect 5907 2216 6013 2224
rect 6067 2216 6153 2224
rect 6167 2216 6193 2224
rect 6456 2216 6493 2224
rect 4607 2196 4684 2204
rect 4696 2196 4773 2204
rect 4307 2176 4384 2184
rect 4676 2184 4684 2196
rect 4787 2196 4813 2204
rect 4887 2196 5053 2204
rect 5167 2196 5293 2204
rect 5427 2196 5473 2204
rect 5687 2196 5873 2204
rect 5927 2196 5953 2204
rect 6456 2204 6464 2216
rect 6507 2216 6573 2224
rect 6207 2196 6464 2204
rect 6487 2196 6633 2204
rect 4676 2176 4753 2184
rect 4987 2176 5333 2184
rect 5367 2176 5433 2184
rect 5767 2176 5853 2184
rect 6227 2176 6373 2184
rect 6387 2176 6453 2184
rect 6476 2176 6593 2184
rect 3707 2156 3744 2164
rect 3756 2156 3853 2164
rect 287 2136 313 2144
rect 407 2136 493 2144
rect 587 2136 733 2144
rect 1367 2136 1933 2144
rect 1967 2136 2293 2144
rect 2307 2136 2373 2144
rect 2467 2136 2524 2144
rect 227 2116 473 2124
rect 487 2116 833 2124
rect 1127 2116 1493 2124
rect 1507 2116 1633 2124
rect 1927 2116 2213 2124
rect 2516 2124 2524 2136
rect 2547 2136 2613 2144
rect 2627 2136 2713 2144
rect 2727 2136 2993 2144
rect 3127 2136 3184 2144
rect 2516 2116 2564 2124
rect 87 2096 133 2104
rect 187 2096 213 2104
rect 327 2096 373 2104
rect 576 2096 593 2104
rect 76 2076 164 2084
rect 76 2064 84 2076
rect 67 2056 84 2064
rect 156 2064 164 2076
rect 187 2076 244 2084
rect 156 2056 184 2064
rect 87 2036 153 2044
rect 176 2044 184 2056
rect 236 2047 244 2076
rect 367 2076 493 2084
rect 367 2056 453 2064
rect 436 2047 444 2056
rect 176 2036 193 2044
rect 347 2036 393 2044
rect 527 2036 533 2044
rect 576 2044 584 2096
rect 767 2096 853 2104
rect 1396 2096 1453 2104
rect 627 2076 633 2084
rect 827 2076 864 2084
rect 616 2064 624 2073
rect 856 2067 864 2076
rect 887 2076 913 2084
rect 967 2076 1013 2084
rect 1027 2076 1033 2084
rect 1056 2067 1064 2093
rect 1396 2084 1404 2096
rect 1567 2096 1613 2104
rect 1736 2096 1813 2104
rect 1356 2076 1404 2084
rect 607 2056 624 2064
rect 667 2056 733 2064
rect 787 2056 813 2064
rect 1196 2064 1204 2073
rect 1356 2067 1364 2076
rect 1507 2076 1573 2084
rect 1736 2084 1744 2096
rect 1976 2096 2133 2104
rect 1727 2076 1744 2084
rect 1827 2076 1853 2084
rect 1976 2084 1984 2096
rect 2556 2104 2564 2116
rect 2587 2116 2633 2124
rect 2647 2116 2813 2124
rect 2827 2116 2913 2124
rect 3176 2124 3184 2136
rect 3227 2136 3293 2144
rect 3347 2136 3393 2144
rect 3416 2136 3653 2144
rect 3416 2124 3424 2136
rect 3667 2136 3713 2144
rect 3736 2144 3744 2156
rect 3867 2156 4033 2164
rect 4087 2156 4453 2164
rect 4467 2156 4533 2164
rect 5007 2156 5133 2164
rect 5147 2156 5313 2164
rect 5527 2156 5933 2164
rect 6107 2156 6233 2164
rect 6476 2164 6484 2176
rect 6407 2156 6484 2164
rect 3736 2136 4273 2144
rect 4387 2136 4453 2144
rect 4467 2136 4573 2144
rect 4587 2136 4633 2144
rect 4687 2136 4873 2144
rect 5036 2136 5093 2144
rect 2987 2116 3024 2124
rect 3176 2116 3424 2124
rect 3436 2116 3504 2124
rect 2556 2096 2724 2104
rect 1956 2076 1984 2084
rect 1196 2056 1264 2064
rect 576 2036 613 2044
rect 807 2036 833 2044
rect 927 2036 973 2044
rect 1187 2036 1233 2044
rect 1256 2044 1264 2056
rect 1456 2044 1464 2073
rect 1487 2056 1513 2064
rect 1567 2056 1633 2064
rect 1647 2056 1653 2064
rect 1716 2047 1724 2073
rect 1747 2056 1873 2064
rect 1256 2036 1464 2044
rect 1956 2044 1964 2076
rect 2007 2076 2113 2084
rect 2387 2076 2493 2084
rect 2716 2084 2724 2096
rect 2767 2096 2853 2104
rect 3016 2104 3024 2116
rect 2947 2096 3004 2104
rect 3016 2096 3124 2104
rect 2667 2076 2704 2084
rect 2716 2076 2744 2084
rect 2276 2064 2284 2073
rect 2276 2056 2344 2064
rect 1956 2036 1993 2044
rect 2287 2036 2313 2044
rect 107 2016 193 2024
rect 207 2016 2093 2024
rect 2336 2024 2344 2056
rect 2596 2064 2604 2073
rect 2596 2056 2673 2064
rect 2416 2044 2424 2053
rect 2416 2036 2433 2044
rect 2547 2036 2593 2044
rect 2696 2044 2704 2076
rect 2647 2036 2704 2044
rect 2127 2016 2673 2024
rect 2736 2024 2744 2076
rect 2756 2064 2764 2073
rect 2756 2056 2833 2064
rect 2876 2044 2884 2073
rect 2976 2064 2984 2073
rect 2927 2056 2984 2064
rect 2996 2044 3004 2096
rect 3116 2087 3124 2096
rect 3027 2076 3104 2084
rect 3096 2064 3104 2076
rect 3136 2084 3144 2093
rect 3136 2076 3164 2084
rect 3156 2067 3164 2076
rect 3256 2076 3353 2084
rect 3096 2056 3133 2064
rect 3256 2064 3264 2076
rect 3436 2084 3444 2116
rect 3436 2076 3453 2084
rect 3496 2084 3504 2116
rect 3547 2116 3833 2124
rect 4027 2116 4193 2124
rect 4547 2116 4713 2124
rect 5036 2124 5044 2136
rect 5127 2136 5173 2144
rect 5207 2136 5213 2144
rect 5227 2136 5333 2144
rect 5387 2136 5793 2144
rect 6247 2136 6324 2144
rect 4847 2116 5044 2124
rect 5067 2116 5253 2124
rect 5447 2116 5653 2124
rect 5667 2116 5684 2124
rect 3627 2096 3813 2104
rect 3967 2096 4013 2104
rect 4047 2096 4133 2104
rect 4347 2096 4433 2104
rect 4627 2096 4653 2104
rect 4816 2096 4893 2104
rect 3496 2076 3573 2084
rect 3587 2076 3673 2084
rect 3236 2056 3264 2064
rect 3236 2047 3244 2056
rect 3327 2056 3393 2064
rect 3496 2056 3733 2064
rect 2876 2036 3004 2044
rect 3067 2036 3173 2044
rect 3496 2044 3504 2056
rect 3787 2056 3813 2064
rect 3876 2064 3884 2073
rect 3936 2067 3944 2093
rect 4207 2076 4233 2084
rect 4387 2076 4413 2084
rect 3876 2056 3913 2064
rect 4096 2064 4104 2073
rect 4096 2056 4173 2064
rect 4336 2064 4344 2073
rect 4336 2056 4453 2064
rect 4676 2064 4684 2073
rect 4667 2056 4684 2064
rect 4707 2056 4733 2064
rect 4796 2064 4804 2073
rect 4756 2056 4804 2064
rect 3487 2036 3504 2044
rect 3667 2036 3753 2044
rect 3907 2036 3953 2044
rect 4016 2044 4024 2053
rect 4756 2047 4764 2056
rect 4007 2036 4024 2044
rect 4287 2036 4533 2044
rect 4587 2036 4613 2044
rect 2736 2016 2953 2024
rect 3007 2016 3113 2024
rect 3447 2016 3673 2024
rect 67 1996 113 2004
rect 187 1996 353 2004
rect 407 1996 893 2004
rect 907 1996 933 2004
rect 947 1996 993 2004
rect 1267 1996 1573 2004
rect 2087 1996 2293 2004
rect 2407 1996 2593 2004
rect 2647 1996 3033 2004
rect 3347 1996 3613 2004
rect 3707 1996 3893 2004
rect 87 1976 293 1984
rect 787 1976 1113 1984
rect 1187 1976 1353 1984
rect 1367 1976 1673 1984
rect 1887 1976 1993 1984
rect 2007 1976 2013 1984
rect 2247 1976 2733 1984
rect 2796 1976 2873 1984
rect 387 1956 493 1964
rect 507 1956 593 1964
rect 987 1956 1053 1964
rect 1067 1956 1093 1964
rect 1107 1956 1413 1964
rect 1447 1956 1473 1964
rect 1487 1956 1633 1964
rect 1647 1956 1793 1964
rect 2087 1956 2393 1964
rect 2507 1956 2553 1964
rect 2796 1964 2804 1976
rect 3407 1976 3713 1984
rect 3767 1976 3933 1984
rect 4056 1984 4064 2033
rect 4107 2016 4173 2024
rect 4447 2016 4753 2024
rect 4816 2024 4824 2096
rect 5307 2096 5384 2104
rect 4847 2076 4893 2084
rect 4836 2064 4844 2073
rect 4836 2056 4853 2064
rect 4956 2064 4964 2093
rect 5067 2076 5093 2084
rect 5107 2076 5113 2084
rect 4896 2056 4964 2064
rect 4896 2047 4904 2056
rect 4976 2047 4984 2073
rect 5036 2064 5044 2073
rect 5136 2067 5144 2093
rect 5376 2084 5384 2096
rect 5407 2096 5424 2104
rect 5376 2076 5393 2084
rect 5036 2056 5104 2064
rect 5096 2044 5104 2056
rect 5096 2036 5113 2044
rect 5156 2044 5164 2073
rect 5196 2044 5204 2073
rect 5416 2064 5424 2096
rect 5567 2096 5593 2104
rect 5507 2076 5573 2084
rect 5627 2076 5664 2084
rect 5367 2056 5424 2064
rect 5467 2056 5553 2064
rect 5607 2056 5633 2064
rect 5156 2036 5533 2044
rect 5656 2044 5664 2076
rect 5676 2067 5684 2116
rect 5967 2116 6213 2124
rect 6316 2124 6324 2136
rect 6347 2136 6553 2144
rect 6316 2116 6353 2124
rect 6376 2116 6433 2124
rect 6376 2104 6384 2116
rect 6456 2116 6504 2124
rect 6027 2096 6384 2104
rect 6456 2104 6464 2116
rect 6427 2096 6464 2104
rect 6496 2104 6504 2116
rect 6527 2116 6653 2124
rect 6496 2096 6533 2104
rect 6556 2096 6593 2104
rect 5856 2076 5933 2084
rect 5856 2067 5864 2076
rect 6067 2076 6093 2084
rect 6247 2076 6293 2084
rect 6396 2084 6404 2093
rect 6396 2076 6464 2084
rect 5767 2056 5793 2064
rect 5887 2056 6013 2064
rect 6176 2064 6184 2073
rect 6456 2067 6464 2076
rect 6527 2076 6544 2084
rect 6176 2056 6293 2064
rect 5587 2036 5664 2044
rect 5676 2036 5933 2044
rect 4816 2016 5013 2024
rect 5047 2016 5393 2024
rect 5676 2024 5684 2036
rect 5976 2036 6493 2044
rect 5467 2016 5684 2024
rect 5976 2024 5984 2036
rect 5707 2016 5984 2024
rect 6536 2024 6544 2076
rect 6556 2047 6564 2096
rect 6696 2096 6733 2104
rect 6696 2084 6704 2096
rect 6596 2076 6704 2084
rect 6596 2044 6604 2076
rect 6627 2056 6693 2064
rect 6576 2036 6604 2044
rect 6576 2024 6584 2036
rect 6107 2016 6144 2024
rect 6536 2016 6584 2024
rect 4087 1996 4124 2004
rect 3996 1976 4064 1984
rect 4116 1984 4124 1996
rect 4167 1996 4433 2004
rect 4116 1976 4173 1984
rect 2687 1956 2804 1964
rect 2827 1956 3093 1964
rect 3127 1956 3553 1964
rect 3747 1956 3833 1964
rect 3996 1964 4004 1976
rect 4256 1967 4264 1996
rect 4827 1996 4933 2004
rect 4967 1996 5093 2004
rect 5116 1996 5253 2004
rect 5116 1984 5124 1996
rect 5267 1996 5553 2004
rect 5787 1996 6113 2004
rect 6136 2004 6144 2016
rect 6136 1996 6413 2004
rect 6587 1996 6653 2004
rect 4307 1976 5124 1984
rect 5167 1976 5273 1984
rect 5427 1976 5753 1984
rect 5827 1976 6173 1984
rect 6227 1976 6573 1984
rect 3927 1956 4004 1964
rect 4447 1956 5213 1964
rect 5907 1956 6333 1964
rect 6347 1956 6653 1964
rect 627 1936 1013 1944
rect 1987 1936 2093 1944
rect 2367 1936 2573 1944
rect 2867 1936 3033 1944
rect 3047 1936 3313 1944
rect 4007 1936 4033 1944
rect 4047 1936 4153 1944
rect 4187 1936 4393 1944
rect 4487 1936 4533 1944
rect 4547 1936 4633 1944
rect 4647 1936 4693 1944
rect 4707 1936 4873 1944
rect 4987 1936 5333 1944
rect 5516 1936 6073 1944
rect 887 1916 1173 1924
rect 1367 1916 1433 1924
rect 2347 1916 2373 1924
rect 2427 1916 2473 1924
rect 2587 1916 2693 1924
rect 2847 1916 3193 1924
rect 3527 1916 4053 1924
rect 4227 1916 4333 1924
rect 4947 1916 5033 1924
rect 5516 1924 5524 1936
rect 6507 1936 6713 1944
rect 5087 1916 5524 1924
rect 5547 1916 5873 1924
rect 5927 1916 6233 1924
rect 6267 1916 6733 1924
rect 167 1896 393 1904
rect 407 1896 833 1904
rect 1027 1896 1393 1904
rect 1527 1896 2013 1904
rect 2147 1896 2793 1904
rect 2807 1896 2893 1904
rect 2907 1896 3353 1904
rect 3407 1896 3453 1904
rect 3587 1896 3813 1904
rect 3907 1896 4044 1904
rect 867 1876 1153 1884
rect 1207 1876 1453 1884
rect 1627 1876 1873 1884
rect 1927 1876 1953 1884
rect 2116 1884 2124 1893
rect 2116 1876 2133 1884
rect 2167 1876 2393 1884
rect 2467 1876 2653 1884
rect 2747 1876 2833 1884
rect 2987 1876 3073 1884
rect 3167 1876 3233 1884
rect 3307 1876 3573 1884
rect 4036 1884 4044 1896
rect 4067 1896 4173 1904
rect 4247 1896 4853 1904
rect 4887 1896 5653 1904
rect 5687 1896 5853 1904
rect 6067 1896 6453 1904
rect 4036 1876 4213 1884
rect 4247 1876 4713 1884
rect 4756 1876 4973 1884
rect 496 1856 753 1864
rect 496 1844 504 1856
rect 847 1856 1213 1864
rect 1327 1856 1733 1864
rect 1967 1856 2213 1864
rect 2447 1856 2533 1864
rect 2787 1856 3513 1864
rect 3807 1856 4093 1864
rect 4107 1856 4353 1864
rect 4756 1864 4764 1876
rect 5036 1876 5493 1884
rect 4707 1856 4764 1864
rect 5036 1864 5044 1876
rect 5516 1876 5553 1884
rect 4887 1856 5044 1864
rect 5096 1856 5453 1864
rect 107 1836 504 1844
rect 647 1836 744 1844
rect 416 1816 493 1824
rect 416 1784 424 1816
rect 607 1816 713 1824
rect 736 1824 744 1836
rect 807 1836 1193 1844
rect 736 1816 893 1824
rect 947 1816 993 1824
rect 1116 1824 1124 1836
rect 1056 1816 1124 1824
rect 447 1796 653 1804
rect 1016 1804 1024 1813
rect 967 1796 1024 1804
rect 227 1776 344 1784
rect 416 1776 453 1784
rect 336 1767 344 1776
rect 496 1776 564 1784
rect 207 1756 313 1764
rect 496 1764 504 1776
rect 467 1756 504 1764
rect 556 1764 564 1776
rect 1056 1784 1064 1816
rect 1156 1824 1164 1836
rect 1247 1836 1273 1844
rect 1367 1836 1384 1844
rect 1376 1827 1384 1836
rect 1827 1836 2293 1844
rect 2327 1836 2773 1844
rect 2887 1836 3053 1844
rect 3296 1836 3353 1844
rect 1156 1816 1204 1824
rect 1047 1776 1064 1784
rect 1136 1767 1144 1813
rect 1196 1807 1204 1816
rect 1216 1816 1253 1824
rect 1216 1784 1224 1816
rect 1307 1816 1333 1824
rect 1396 1804 1404 1833
rect 2027 1816 2493 1824
rect 2727 1816 2804 1824
rect 1387 1796 1404 1804
rect 1927 1796 2084 1804
rect 1187 1776 1224 1784
rect 1416 1776 1453 1784
rect 1416 1767 1424 1776
rect 556 1756 733 1764
rect 927 1756 1113 1764
rect 1507 1756 1633 1764
rect 1816 1744 1824 1773
rect 1836 1764 1844 1793
rect 1867 1776 2013 1784
rect 2076 1784 2084 1796
rect 2107 1796 2424 1804
rect 2076 1776 2293 1784
rect 2387 1776 2404 1784
rect 1836 1756 1913 1764
rect 1987 1756 2373 1764
rect 887 1736 1824 1744
rect 1867 1736 2133 1744
rect 2147 1736 2173 1744
rect 2396 1744 2404 1776
rect 2416 1764 2424 1796
rect 2796 1804 2804 1816
rect 2847 1816 3133 1824
rect 2467 1796 2524 1804
rect 2796 1796 2853 1804
rect 2436 1784 2444 1793
rect 2436 1776 2493 1784
rect 2416 1756 2433 1764
rect 2516 1764 2524 1796
rect 2876 1804 2884 1816
rect 3296 1824 3304 1836
rect 3367 1836 3393 1844
rect 3687 1836 3853 1844
rect 3867 1836 4033 1844
rect 4316 1836 4333 1844
rect 3187 1816 3304 1824
rect 2876 1796 3024 1804
rect 2607 1776 2813 1784
rect 2907 1776 2953 1784
rect 2976 1776 2993 1784
rect 2976 1767 2984 1776
rect 3016 1784 3024 1796
rect 3047 1796 3173 1804
rect 3016 1776 3053 1784
rect 3196 1784 3204 1816
rect 3447 1816 3513 1824
rect 3827 1816 3853 1824
rect 4007 1816 4293 1824
rect 3316 1804 3324 1813
rect 3287 1796 3324 1804
rect 3176 1776 3204 1784
rect 3176 1767 3184 1776
rect 3776 1784 3784 1813
rect 3847 1796 3873 1804
rect 3896 1784 3904 1813
rect 4316 1807 4324 1836
rect 4487 1836 4573 1844
rect 4616 1836 4653 1844
rect 4616 1824 4624 1836
rect 4667 1836 4713 1844
rect 5096 1844 5104 1856
rect 5516 1864 5524 1876
rect 5587 1876 6153 1884
rect 6187 1876 6693 1884
rect 5496 1856 5524 1864
rect 4827 1836 5104 1844
rect 5127 1836 5233 1844
rect 5247 1836 5324 1844
rect 4396 1816 4624 1824
rect 4187 1796 4224 1804
rect 3507 1776 3544 1784
rect 3776 1776 3904 1784
rect 4216 1784 4224 1796
rect 4216 1776 4273 1784
rect 2456 1756 2524 1764
rect 2227 1736 2404 1744
rect 2456 1744 2464 1756
rect 2547 1756 2633 1764
rect 2707 1756 2793 1764
rect 2807 1756 2953 1764
rect 3207 1756 3253 1764
rect 3327 1756 3373 1764
rect 3487 1756 3513 1764
rect 3536 1764 3544 1776
rect 3536 1756 3693 1764
rect 3707 1756 3853 1764
rect 3896 1764 3904 1776
rect 4396 1784 4404 1816
rect 4516 1787 4524 1816
rect 5027 1816 5133 1824
rect 5167 1816 5293 1824
rect 5316 1807 5324 1836
rect 5496 1844 5504 1856
rect 5547 1856 5593 1864
rect 5607 1856 5893 1864
rect 5967 1856 6093 1864
rect 6127 1856 6173 1864
rect 6407 1856 6433 1864
rect 6547 1856 6573 1864
rect 5447 1836 5504 1844
rect 5527 1836 5693 1844
rect 5856 1836 5964 1844
rect 5596 1816 5653 1824
rect 4576 1796 4613 1804
rect 4307 1776 4404 1784
rect 4447 1776 4473 1784
rect 4576 1784 4584 1796
rect 4696 1796 4713 1804
rect 4556 1776 4584 1784
rect 3896 1756 3953 1764
rect 4167 1756 4353 1764
rect 4367 1756 4424 1764
rect 2427 1736 2464 1744
rect 2607 1736 2673 1744
rect 2727 1736 2893 1744
rect 3147 1736 3333 1744
rect 3887 1736 4084 1744
rect 387 1716 593 1724
rect 767 1716 1553 1724
rect 1687 1716 2073 1724
rect 2307 1716 2533 1724
rect 2567 1716 2733 1724
rect 2787 1716 3013 1724
rect 3087 1716 3213 1724
rect 3327 1716 3653 1724
rect 3787 1716 3793 1724
rect 3807 1716 3973 1724
rect 4076 1724 4084 1736
rect 4107 1736 4173 1744
rect 4236 1736 4293 1744
rect 4236 1724 4244 1736
rect 4356 1736 4393 1744
rect 4076 1716 4244 1724
rect 4356 1724 4364 1736
rect 4416 1744 4424 1756
rect 4467 1756 4513 1764
rect 4556 1764 4564 1776
rect 4696 1784 4704 1796
rect 4767 1796 4973 1804
rect 5116 1796 5193 1804
rect 4687 1776 4704 1784
rect 4736 1784 4744 1793
rect 4736 1776 4873 1784
rect 5116 1784 5124 1796
rect 5216 1796 5273 1804
rect 5067 1776 5124 1784
rect 4547 1756 4564 1764
rect 4607 1756 4853 1764
rect 4867 1756 4913 1764
rect 5007 1756 5093 1764
rect 5127 1756 5173 1764
rect 5216 1764 5224 1796
rect 5476 1804 5484 1813
rect 5396 1796 5484 1804
rect 5247 1776 5353 1784
rect 5207 1756 5224 1764
rect 5396 1764 5404 1796
rect 5536 1784 5544 1813
rect 5596 1807 5604 1816
rect 5687 1816 5704 1824
rect 5567 1796 5584 1804
rect 5427 1776 5544 1784
rect 5576 1784 5584 1796
rect 5696 1804 5704 1816
rect 5727 1816 5773 1824
rect 5696 1796 5733 1804
rect 5576 1776 5593 1784
rect 5856 1784 5864 1836
rect 5956 1824 5964 1836
rect 5987 1836 6224 1844
rect 5956 1816 6193 1824
rect 5907 1796 5973 1804
rect 5987 1796 6133 1804
rect 6216 1804 6224 1836
rect 6327 1836 6633 1844
rect 6307 1816 6333 1824
rect 6447 1816 6493 1824
rect 6516 1816 6593 1824
rect 6216 1796 6244 1804
rect 5636 1776 5864 1784
rect 5636 1767 5644 1776
rect 5947 1776 5973 1784
rect 6136 1767 6144 1793
rect 6167 1776 6213 1784
rect 6236 1767 6244 1796
rect 6376 1804 6384 1813
rect 6516 1804 6524 1816
rect 6356 1796 6384 1804
rect 6496 1796 6524 1804
rect 5247 1756 5493 1764
rect 5516 1756 5613 1764
rect 4416 1736 4533 1744
rect 4707 1736 4733 1744
rect 4987 1736 5093 1744
rect 5127 1736 5253 1744
rect 5516 1744 5524 1756
rect 5967 1756 5993 1764
rect 6276 1764 6284 1793
rect 6356 1784 6364 1796
rect 6296 1776 6364 1784
rect 6296 1767 6304 1776
rect 6496 1784 6504 1796
rect 6547 1796 6613 1804
rect 6387 1776 6504 1784
rect 6267 1756 6284 1764
rect 6327 1756 6413 1764
rect 6496 1764 6504 1776
rect 6527 1776 6553 1784
rect 6496 1756 6513 1764
rect 5447 1736 5524 1744
rect 5607 1736 5693 1744
rect 5707 1736 5713 1744
rect 5867 1736 6073 1744
rect 6167 1736 6313 1744
rect 4267 1716 4364 1724
rect 4387 1716 4573 1724
rect 4587 1716 4893 1724
rect 5207 1716 5573 1724
rect 5587 1716 5604 1724
rect 507 1696 953 1704
rect 1307 1696 1393 1704
rect 1707 1696 1813 1704
rect 1907 1696 1953 1704
rect 2287 1696 2613 1704
rect 2787 1696 2873 1704
rect 2987 1696 3033 1704
rect 3147 1696 3293 1704
rect 3687 1696 3853 1704
rect 3887 1696 4093 1704
rect 4207 1696 4253 1704
rect 4467 1696 4493 1704
rect 4507 1696 5344 1704
rect 607 1676 1273 1684
rect 1387 1676 1493 1684
rect 1527 1676 2813 1684
rect 3047 1676 3113 1684
rect 3167 1676 4053 1684
rect 4136 1676 4153 1684
rect 367 1656 573 1664
rect 1187 1656 1353 1664
rect 1487 1656 2013 1664
rect 2367 1656 2513 1664
rect 2587 1656 2633 1664
rect 2667 1656 3093 1664
rect 3116 1656 3553 1664
rect 727 1636 1133 1644
rect 1147 1636 1193 1644
rect 1267 1636 1324 1644
rect 27 1616 53 1624
rect 107 1616 193 1624
rect 496 1607 504 1633
rect 587 1616 1053 1624
rect 1107 1616 1213 1624
rect 1227 1616 1264 1624
rect -24 1596 33 1604
rect 47 1596 64 1604
rect 56 1584 64 1596
rect 87 1596 173 1604
rect 1076 1587 1084 1613
rect 1147 1596 1213 1604
rect 56 1576 93 1584
rect 127 1576 153 1584
rect 567 1576 593 1584
rect 647 1576 684 1584
rect 167 1556 393 1564
rect 407 1556 453 1564
rect 676 1564 684 1576
rect 676 1556 773 1564
rect 1096 1564 1104 1593
rect 1127 1576 1233 1584
rect 1256 1567 1264 1616
rect 1316 1584 1324 1636
rect 1467 1636 1533 1644
rect 1607 1636 1753 1644
rect 1847 1636 2233 1644
rect 2287 1636 2313 1644
rect 2387 1636 2473 1644
rect 2687 1636 2913 1644
rect 2927 1636 3033 1644
rect 3116 1644 3124 1656
rect 3607 1656 3673 1664
rect 3727 1656 4013 1664
rect 3067 1636 3124 1644
rect 3327 1636 3373 1644
rect 3387 1636 3473 1644
rect 3827 1636 3873 1644
rect 3927 1636 4113 1644
rect 1456 1616 1533 1624
rect 1316 1576 1353 1584
rect 1416 1567 1424 1593
rect 1456 1584 1464 1616
rect 1767 1616 1853 1624
rect 1876 1616 1964 1624
rect 1616 1604 1624 1613
rect 1496 1596 1624 1604
rect 1447 1576 1464 1584
rect 1476 1567 1484 1593
rect 1496 1587 1504 1596
rect 1727 1596 1773 1604
rect 1876 1604 1884 1616
rect 1787 1596 1884 1604
rect 1956 1604 1964 1616
rect 2207 1616 2353 1624
rect 2407 1616 2453 1624
rect 2467 1616 2553 1624
rect 2656 1616 2693 1624
rect 1956 1596 2013 1604
rect 2027 1596 2084 1604
rect 1527 1576 1553 1584
rect 1647 1576 1873 1584
rect 2076 1584 2084 1596
rect 2156 1596 2213 1604
rect 2076 1576 2093 1584
rect 2156 1584 2164 1596
rect 2236 1596 2413 1604
rect 2236 1587 2244 1596
rect 2656 1604 2664 1616
rect 2747 1616 2853 1624
rect 2867 1616 3213 1624
rect 3407 1616 3533 1624
rect 3807 1616 3824 1624
rect 2567 1596 2664 1604
rect 2576 1587 2584 1596
rect 2687 1596 2773 1604
rect 3447 1596 3524 1604
rect 3516 1587 3524 1596
rect 3816 1604 3824 1616
rect 3847 1616 3993 1624
rect 4136 1624 4144 1676
rect 4187 1676 4593 1684
rect 4647 1676 4873 1684
rect 4907 1676 4984 1684
rect 4407 1656 4473 1664
rect 4527 1656 4553 1664
rect 4607 1656 4713 1664
rect 4827 1656 4853 1664
rect 4976 1664 4984 1676
rect 5076 1676 5173 1684
rect 4976 1656 5013 1664
rect 4307 1636 4413 1644
rect 4427 1636 4753 1644
rect 4927 1636 5053 1644
rect 4027 1616 4144 1624
rect 4336 1616 4353 1624
rect 3816 1596 3833 1604
rect 4336 1604 4344 1616
rect 5076 1624 5084 1676
rect 5227 1676 5253 1684
rect 5336 1684 5344 1696
rect 5367 1696 5473 1704
rect 5596 1704 5604 1716
rect 5687 1716 5864 1724
rect 5596 1696 5833 1704
rect 5856 1704 5864 1716
rect 6207 1716 6333 1724
rect 5856 1696 5893 1704
rect 6047 1696 6233 1704
rect 6407 1696 6453 1704
rect 5327 1676 5373 1684
rect 5547 1676 5633 1684
rect 5667 1676 5693 1684
rect 5767 1676 6073 1684
rect 6127 1676 6204 1684
rect 5107 1656 5644 1664
rect 4727 1616 5084 1624
rect 5116 1636 5253 1644
rect 4247 1596 4344 1604
rect 2116 1576 2164 1584
rect 1067 1556 1104 1564
rect 1287 1556 1313 1564
rect 2116 1564 2124 1576
rect 3367 1576 3413 1584
rect 3696 1584 3704 1593
rect 3696 1576 3813 1584
rect 4516 1584 4524 1613
rect 5016 1607 5024 1616
rect 4616 1596 4653 1604
rect 4267 1576 4524 1584
rect 4536 1584 4544 1593
rect 4616 1584 4624 1596
rect 4736 1596 4833 1604
rect 4536 1576 4624 1584
rect 4736 1584 4744 1596
rect 4967 1596 5004 1604
rect 4707 1576 4744 1584
rect 4896 1584 4904 1593
rect 4827 1576 4904 1584
rect 4996 1584 5004 1596
rect 5067 1596 5093 1604
rect 5116 1604 5124 1636
rect 5447 1636 5613 1644
rect 5636 1644 5644 1656
rect 5667 1656 5813 1664
rect 5907 1656 5913 1664
rect 5927 1656 6053 1664
rect 6196 1664 6204 1676
rect 6227 1676 6593 1684
rect 6127 1656 6164 1664
rect 6196 1656 6233 1664
rect 5636 1636 5793 1644
rect 6116 1636 6133 1644
rect 5247 1616 5473 1624
rect 5487 1616 5533 1624
rect 5616 1616 5653 1624
rect 5116 1596 5133 1604
rect 5167 1596 5213 1604
rect 5227 1596 5253 1604
rect 5347 1596 5524 1604
rect 4996 1576 5013 1584
rect 5127 1576 5353 1584
rect 5467 1576 5493 1584
rect 5516 1584 5524 1596
rect 5616 1604 5624 1616
rect 5687 1616 5704 1624
rect 5567 1596 5624 1604
rect 5516 1576 5544 1584
rect 1967 1556 2124 1564
rect 2807 1556 2824 1564
rect 616 1544 624 1553
rect 616 1536 913 1544
rect 1167 1536 1353 1544
rect 1507 1536 1733 1544
rect 2007 1536 2153 1544
rect 2167 1536 2473 1544
rect 2527 1536 2793 1544
rect 2816 1544 2824 1556
rect 3067 1556 3224 1564
rect 2816 1536 2953 1544
rect 3216 1544 3224 1556
rect 3247 1556 3293 1564
rect 3347 1556 3573 1564
rect 3867 1556 4333 1564
rect 4667 1556 4793 1564
rect 4927 1556 4993 1564
rect 3216 1536 3713 1544
rect 4387 1536 4473 1544
rect 4507 1536 4733 1544
rect 4807 1536 5013 1544
rect 5536 1544 5544 1576
rect 5576 1576 5593 1584
rect 5576 1564 5584 1576
rect 5567 1556 5584 1564
rect 5676 1564 5684 1593
rect 5696 1584 5704 1616
rect 5847 1616 5973 1624
rect 5727 1596 5824 1604
rect 5696 1576 5733 1584
rect 5816 1584 5824 1596
rect 5987 1596 6093 1604
rect 6116 1604 6124 1636
rect 6156 1644 6164 1656
rect 6267 1656 6433 1664
rect 6156 1636 6173 1644
rect 6307 1636 6333 1644
rect 6367 1636 6393 1644
rect 6407 1616 6484 1624
rect 6476 1607 6484 1616
rect 6116 1596 6224 1604
rect 5816 1576 5844 1584
rect 5836 1567 5844 1576
rect 5947 1576 5993 1584
rect 6087 1576 6193 1584
rect 6216 1584 6224 1596
rect 6276 1596 6293 1604
rect 6216 1576 6233 1584
rect 6276 1584 6284 1596
rect 6256 1576 6284 1584
rect 5676 1556 5793 1564
rect 5907 1556 5953 1564
rect 5987 1556 6113 1564
rect 6147 1556 6233 1564
rect 5536 1536 5973 1544
rect 6256 1544 6264 1576
rect 6387 1576 6653 1584
rect 6287 1556 6313 1564
rect 6007 1536 6293 1544
rect 447 1516 653 1524
rect 1007 1516 1413 1524
rect 1427 1516 1593 1524
rect 1607 1516 1693 1524
rect 1887 1516 2273 1524
rect 2307 1516 2853 1524
rect 3407 1516 4013 1524
rect 4327 1516 4653 1524
rect 5267 1516 5493 1524
rect 5547 1516 5613 1524
rect 5707 1516 6093 1524
rect 6127 1516 6193 1524
rect 947 1496 1313 1504
rect 1587 1496 1673 1504
rect 2907 1496 3353 1504
rect 3627 1496 3793 1504
rect 3827 1496 4193 1504
rect 4207 1496 4553 1504
rect 4607 1496 4633 1504
rect 4647 1496 5013 1504
rect 5036 1496 5233 1504
rect 1407 1476 1973 1484
rect 1996 1476 2573 1484
rect 1187 1456 1213 1464
rect 1996 1464 2004 1476
rect 3027 1476 3424 1484
rect 1627 1456 2004 1464
rect 2067 1456 2213 1464
rect 2347 1456 3313 1464
rect 3416 1464 3424 1476
rect 3467 1476 3693 1484
rect 3727 1476 4044 1484
rect 3416 1456 3473 1464
rect 4036 1464 4044 1476
rect 4067 1476 4093 1484
rect 4347 1476 4393 1484
rect 5036 1484 5044 1496
rect 5267 1496 5553 1504
rect 5567 1496 5633 1504
rect 4427 1476 5044 1484
rect 5067 1476 5353 1484
rect 5387 1476 5413 1484
rect 5447 1476 5633 1484
rect 5827 1476 5853 1484
rect 4036 1456 5153 1464
rect 5207 1456 5473 1464
rect 5507 1456 5593 1464
rect 5607 1456 5733 1464
rect 5787 1456 5833 1464
rect 6047 1456 6413 1464
rect 1447 1436 1753 1444
rect 2247 1436 2313 1444
rect 2367 1436 3053 1444
rect 3507 1436 3593 1444
rect 3707 1436 3853 1444
rect 3967 1436 4173 1444
rect 4196 1436 4253 1444
rect 1087 1416 1373 1424
rect 1387 1416 1473 1424
rect 1487 1416 1733 1424
rect 1787 1416 2173 1424
rect 2187 1416 2293 1424
rect 2467 1416 2653 1424
rect 2767 1416 2853 1424
rect 2987 1416 3253 1424
rect 3287 1416 3373 1424
rect 3407 1416 3713 1424
rect 4196 1424 4204 1436
rect 4267 1436 4813 1444
rect 5327 1436 5673 1444
rect 6127 1436 6673 1444
rect 3767 1416 4204 1424
rect 4247 1416 4453 1424
rect 4507 1416 4593 1424
rect 4947 1416 5273 1424
rect 5387 1416 5493 1424
rect 5527 1416 5693 1424
rect 5767 1416 5913 1424
rect 6167 1416 6253 1424
rect 6527 1416 6553 1424
rect 807 1396 1413 1404
rect 1767 1396 2233 1404
rect 2267 1396 2613 1404
rect 2967 1396 3133 1404
rect 3267 1396 3773 1404
rect 3787 1396 4073 1404
rect 4087 1396 4773 1404
rect 4787 1396 4953 1404
rect 5327 1396 5393 1404
rect 5447 1396 5733 1404
rect 5747 1396 5773 1404
rect 5827 1396 5893 1404
rect 5987 1396 6533 1404
rect 287 1376 1333 1384
rect 1347 1376 1573 1384
rect 1687 1376 1713 1384
rect 1727 1376 1993 1384
rect 2007 1376 2073 1384
rect 2247 1376 2293 1384
rect 2967 1376 3953 1384
rect 3987 1376 4153 1384
rect 4296 1376 4853 1384
rect 207 1356 233 1364
rect 267 1356 293 1364
rect 307 1356 533 1364
rect 547 1356 873 1364
rect 927 1356 973 1364
rect 1016 1356 1253 1364
rect 1016 1347 1024 1356
rect 1567 1356 1633 1364
rect 1667 1356 1753 1364
rect 1947 1356 2053 1364
rect 2067 1356 2113 1364
rect 2167 1356 2193 1364
rect 2227 1356 2384 1364
rect 27 1336 53 1344
rect 187 1336 413 1344
rect 787 1336 933 1344
rect 1627 1336 1833 1344
rect 2187 1336 2273 1344
rect 516 1324 524 1333
rect 467 1316 524 1324
rect 547 1316 573 1324
rect 627 1316 733 1324
rect 967 1316 1144 1324
rect 156 1296 213 1304
rect 27 1276 73 1284
rect 87 1276 113 1284
rect 156 1284 164 1296
rect 287 1296 313 1304
rect 396 1287 404 1313
rect 616 1304 624 1313
rect 1136 1307 1144 1316
rect 1327 1316 1433 1324
rect 1756 1316 1773 1324
rect 1756 1307 1764 1316
rect 427 1296 624 1304
rect 647 1296 753 1304
rect 907 1296 973 1304
rect 987 1296 993 1304
rect 1187 1296 1253 1304
rect 1707 1296 1733 1304
rect 1876 1304 1884 1333
rect 1907 1316 1953 1324
rect 1976 1324 1984 1333
rect 1976 1316 2004 1324
rect 1876 1296 1973 1304
rect 1996 1287 2004 1316
rect 2087 1316 2104 1324
rect 2096 1307 2104 1316
rect 2167 1316 2213 1324
rect 2296 1304 2304 1333
rect 2376 1324 2384 1356
rect 2507 1356 2633 1364
rect 2407 1336 2593 1344
rect 2616 1344 2624 1356
rect 2727 1356 3113 1364
rect 3247 1356 3704 1364
rect 2616 1336 2933 1344
rect 3007 1336 3073 1344
rect 3227 1336 3393 1344
rect 3467 1336 3564 1344
rect 2376 1316 2424 1324
rect 2416 1307 2424 1316
rect 2447 1316 2544 1324
rect 2536 1307 2544 1316
rect 2747 1316 2953 1324
rect 2976 1324 2984 1333
rect 2976 1316 3004 1324
rect 2296 1296 2353 1304
rect 2556 1296 2713 1304
rect 2556 1287 2564 1296
rect 147 1276 164 1284
rect 327 1276 353 1284
rect 487 1276 793 1284
rect 876 1276 1033 1284
rect 376 1264 384 1273
rect 876 1267 884 1276
rect 1607 1276 1633 1284
rect 1787 1276 1833 1284
rect 2027 1276 2393 1284
rect 2456 1276 2473 1284
rect 307 1256 384 1264
rect 607 1256 633 1264
rect 747 1256 773 1264
rect 1647 1256 1833 1264
rect 1947 1256 2033 1264
rect 2047 1256 2293 1264
rect 2456 1264 2464 1276
rect 2727 1276 2773 1284
rect 2827 1276 2953 1284
rect 2996 1284 3004 1316
rect 3047 1316 3093 1324
rect 3027 1296 3333 1304
rect 3407 1296 3513 1304
rect 3556 1304 3564 1336
rect 3696 1344 3704 1356
rect 4296 1364 4304 1376
rect 4867 1376 4944 1384
rect 3727 1356 4304 1364
rect 4327 1356 4453 1364
rect 4556 1356 4613 1364
rect 3667 1336 3684 1344
rect 3696 1336 3873 1344
rect 3676 1324 3684 1336
rect 3927 1336 4233 1344
rect 4347 1336 4413 1344
rect 4447 1336 4544 1344
rect 3627 1316 3664 1324
rect 3676 1316 3713 1324
rect 3656 1304 3664 1316
rect 4367 1316 4413 1324
rect 3556 1296 3604 1304
rect 3656 1296 3733 1304
rect 2996 1276 3033 1284
rect 3247 1276 3404 1284
rect 2327 1256 2464 1264
rect 2487 1256 3373 1264
rect 3396 1264 3404 1276
rect 3547 1276 3573 1284
rect 3596 1284 3604 1296
rect 4007 1296 4093 1304
rect 4347 1296 4393 1304
rect 4516 1287 4524 1313
rect 4536 1307 4544 1336
rect 4556 1324 4564 1356
rect 4647 1356 4713 1364
rect 4587 1336 4604 1344
rect 4556 1316 4573 1324
rect 4596 1307 4604 1336
rect 4656 1336 4713 1344
rect 4656 1324 4664 1336
rect 4827 1336 4913 1344
rect 4936 1344 4944 1376
rect 4967 1376 5073 1384
rect 5087 1376 5573 1384
rect 5727 1376 5844 1384
rect 5007 1356 5253 1364
rect 5367 1356 5493 1364
rect 5507 1356 5653 1364
rect 5727 1356 5793 1364
rect 5836 1364 5844 1376
rect 6087 1376 6173 1384
rect 5836 1356 5864 1364
rect 4936 1336 4984 1344
rect 4627 1316 4664 1324
rect 4936 1316 4953 1324
rect 4936 1307 4944 1316
rect 4747 1296 4804 1304
rect 3596 1276 3613 1284
rect 3707 1276 3953 1284
rect 3967 1276 4193 1284
rect 4207 1276 4333 1284
rect 4367 1276 4433 1284
rect 4727 1276 4753 1284
rect 4767 1276 4773 1284
rect 4796 1284 4804 1296
rect 4976 1304 4984 1336
rect 5056 1336 5113 1344
rect 5056 1324 5064 1336
rect 5127 1336 5153 1344
rect 5187 1336 5224 1344
rect 5047 1316 5064 1324
rect 5136 1316 5193 1324
rect 4967 1296 4984 1304
rect 4796 1276 5033 1284
rect 3396 1256 3733 1264
rect 3807 1256 3833 1264
rect 4307 1256 4433 1264
rect 5076 1264 5084 1313
rect 5136 1304 5144 1316
rect 5107 1296 5144 1304
rect 5216 1304 5224 1336
rect 5247 1336 5513 1344
rect 5536 1336 5613 1344
rect 5247 1316 5333 1324
rect 5447 1316 5484 1324
rect 5216 1296 5253 1304
rect 5287 1296 5353 1304
rect 5367 1296 5373 1304
rect 5476 1304 5484 1316
rect 5476 1296 5504 1304
rect 5456 1284 5464 1293
rect 5496 1284 5504 1296
rect 5536 1304 5544 1336
rect 5816 1344 5824 1353
rect 5747 1336 5804 1344
rect 5816 1336 5833 1344
rect 5527 1296 5544 1304
rect 5556 1287 5564 1313
rect 5256 1276 5484 1284
rect 5496 1276 5513 1284
rect 4647 1256 5093 1264
rect 5256 1264 5264 1276
rect 5227 1256 5264 1264
rect 5347 1256 5453 1264
rect 5476 1264 5484 1276
rect 5576 1284 5584 1313
rect 5796 1307 5804 1336
rect 5747 1296 5773 1304
rect 5856 1304 5864 1356
rect 5876 1356 5913 1364
rect 5876 1327 5884 1356
rect 5947 1356 6113 1364
rect 6136 1356 6353 1364
rect 5907 1336 5944 1344
rect 5936 1307 5944 1336
rect 5967 1316 5973 1324
rect 5987 1316 6064 1324
rect 5856 1296 5873 1304
rect 6056 1304 6064 1316
rect 6116 1324 6124 1333
rect 6087 1316 6124 1324
rect 6056 1296 6113 1304
rect 6136 1304 6144 1356
rect 6176 1336 6193 1344
rect 6136 1296 6153 1304
rect 6176 1287 6184 1336
rect 6216 1316 6253 1324
rect 5576 1276 5773 1284
rect 5907 1276 6164 1284
rect 5476 1256 5653 1264
rect 5767 1256 5813 1264
rect 5887 1256 6013 1264
rect 6027 1256 6053 1264
rect 6156 1264 6164 1276
rect 6216 1284 6224 1316
rect 6687 1316 6713 1324
rect 6507 1296 6673 1304
rect 6207 1276 6224 1284
rect 6347 1276 6533 1284
rect 6547 1276 6573 1284
rect 6067 1256 6144 1264
rect 6156 1256 6693 1264
rect 207 1236 333 1244
rect 447 1236 653 1244
rect 1467 1236 1533 1244
rect 1547 1236 1793 1244
rect 1827 1236 2053 1244
rect 2387 1236 2553 1244
rect 2587 1236 2804 1244
rect 1567 1216 1773 1224
rect 1787 1216 2433 1224
rect 2447 1216 2773 1224
rect 2796 1224 2804 1236
rect 2827 1236 2853 1244
rect 2987 1236 3053 1244
rect 3076 1236 3573 1244
rect 2796 1216 2904 1224
rect 1767 1196 1813 1204
rect 1967 1196 2033 1204
rect 2187 1196 2253 1204
rect 2267 1196 2333 1204
rect 2496 1196 2533 1204
rect 627 1176 813 1184
rect 2496 1184 2504 1196
rect 2747 1196 2853 1204
rect 2127 1176 2504 1184
rect 2527 1176 2553 1184
rect 2787 1176 2873 1184
rect 307 1156 373 1164
rect 407 1156 713 1164
rect 767 1156 813 1164
rect 927 1156 1004 1164
rect 127 1136 184 1144
rect 107 1116 153 1124
rect 176 1124 184 1136
rect 316 1136 413 1144
rect 316 1124 324 1136
rect 427 1136 473 1144
rect 807 1136 973 1144
rect 176 1116 324 1124
rect 347 1116 373 1124
rect 776 1116 833 1124
rect 456 1104 464 1113
rect 247 1096 464 1104
rect 667 1096 693 1104
rect 776 1104 784 1116
rect 867 1116 953 1124
rect 707 1096 784 1104
rect 996 1104 1004 1156
rect 1567 1156 1873 1164
rect 1927 1156 1953 1164
rect 2107 1156 2753 1164
rect 2847 1156 2873 1164
rect 1807 1136 1893 1144
rect 1976 1136 2033 1144
rect 1687 1116 1933 1124
rect 1976 1124 1984 1136
rect 2067 1136 2093 1144
rect 2167 1136 2213 1144
rect 2327 1136 2393 1144
rect 2447 1136 2464 1144
rect 1956 1116 1984 1124
rect 987 1096 1004 1104
rect 1307 1096 1333 1104
rect 1447 1096 1573 1104
rect 1887 1096 1933 1104
rect 1956 1104 1964 1116
rect 2116 1124 2124 1133
rect 2067 1116 2124 1124
rect 2276 1116 2293 1124
rect 1947 1096 1964 1104
rect 587 1076 604 1084
rect 596 1024 604 1076
rect 796 1084 804 1093
rect 767 1076 804 1084
rect 847 1056 893 1064
rect 916 1064 924 1093
rect 947 1076 953 1084
rect 967 1076 993 1084
rect 1187 1076 1433 1084
rect 1836 1084 1844 1093
rect 1836 1076 1913 1084
rect 2256 1084 2264 1113
rect 2276 1104 2284 1116
rect 2456 1124 2464 1136
rect 2487 1136 2593 1144
rect 2516 1127 2524 1136
rect 2896 1144 2904 1216
rect 3076 1224 3084 1236
rect 3616 1236 3864 1244
rect 2947 1216 3084 1224
rect 3207 1216 3313 1224
rect 3507 1216 3513 1224
rect 3616 1224 3624 1236
rect 3527 1216 3624 1224
rect 3727 1216 3753 1224
rect 3856 1224 3864 1236
rect 4027 1236 4493 1244
rect 4527 1236 4793 1244
rect 4827 1236 4893 1244
rect 4947 1236 5024 1244
rect 3856 1216 4153 1224
rect 4247 1216 4293 1224
rect 4327 1216 4473 1224
rect 4596 1216 4773 1224
rect 3287 1196 3393 1204
rect 3407 1196 3693 1204
rect 4596 1204 4604 1216
rect 4787 1216 4833 1224
rect 4927 1216 4973 1224
rect 5016 1224 5024 1236
rect 5047 1236 5253 1244
rect 5407 1236 5693 1244
rect 5727 1236 5793 1244
rect 5867 1236 5913 1244
rect 6047 1236 6113 1244
rect 6136 1244 6144 1256
rect 6136 1236 6553 1244
rect 5016 1216 5113 1224
rect 5187 1216 5373 1224
rect 5396 1216 5473 1224
rect 4067 1196 4604 1204
rect 4627 1196 4653 1204
rect 5396 1204 5404 1216
rect 5567 1216 5633 1224
rect 5687 1216 5993 1224
rect 6007 1216 6233 1224
rect 6287 1216 6733 1224
rect 5327 1196 5404 1204
rect 5427 1196 6033 1204
rect 6107 1196 6153 1204
rect 6167 1196 6233 1204
rect 6267 1196 6653 1204
rect 3147 1176 3244 1184
rect 2927 1156 2984 1164
rect 2887 1136 2904 1144
rect 2976 1144 2984 1156
rect 3147 1156 3213 1164
rect 3236 1164 3244 1176
rect 3267 1176 3473 1184
rect 3867 1176 3933 1184
rect 3947 1176 4093 1184
rect 4167 1176 4753 1184
rect 4807 1176 4913 1184
rect 4927 1176 4993 1184
rect 5167 1176 5204 1184
rect 3236 1156 3533 1164
rect 3607 1156 3673 1164
rect 3707 1156 3773 1164
rect 3827 1156 3873 1164
rect 3907 1156 4053 1164
rect 4167 1156 4173 1164
rect 4187 1156 4244 1164
rect 2976 1136 3084 1144
rect 2456 1116 2473 1124
rect 2556 1116 2613 1124
rect 2276 1096 2344 1104
rect 2256 1076 2313 1084
rect 2336 1084 2344 1096
rect 2556 1104 2564 1116
rect 2816 1124 2824 1133
rect 2687 1116 2824 1124
rect 2527 1096 2564 1104
rect 2587 1096 2633 1104
rect 2656 1087 2664 1113
rect 2696 1104 2704 1116
rect 3007 1116 3053 1124
rect 3076 1124 3084 1136
rect 3107 1136 3233 1144
rect 3367 1136 3593 1144
rect 3607 1136 3913 1144
rect 4007 1136 4033 1144
rect 4127 1136 4193 1144
rect 4236 1144 4244 1156
rect 4587 1156 4833 1164
rect 5027 1156 5053 1164
rect 5127 1156 5173 1164
rect 5196 1164 5204 1176
rect 5247 1176 5293 1184
rect 5367 1176 5413 1184
rect 5487 1176 5833 1184
rect 5996 1176 6113 1184
rect 5196 1156 5453 1164
rect 5556 1156 5644 1164
rect 4236 1136 4273 1144
rect 4307 1136 4353 1144
rect 4407 1136 4504 1144
rect 3076 1116 3204 1124
rect 3196 1107 3204 1116
rect 3216 1116 3433 1124
rect 2696 1096 2793 1104
rect 2336 1076 2573 1084
rect 2676 1084 2684 1093
rect 2676 1076 2733 1084
rect 2787 1076 3113 1084
rect 3216 1084 3224 1116
rect 3647 1116 3693 1124
rect 3827 1116 3873 1124
rect 3896 1116 3933 1124
rect 3247 1096 3273 1104
rect 3316 1096 3413 1104
rect 3316 1087 3324 1096
rect 3187 1076 3224 1084
rect 3267 1076 3293 1084
rect 3496 1084 3504 1113
rect 3556 1087 3564 1113
rect 3896 1104 3904 1116
rect 3967 1116 4053 1124
rect 4076 1107 4084 1133
rect 4247 1116 4393 1124
rect 3687 1096 3904 1104
rect 4156 1104 4164 1113
rect 4496 1107 4504 1136
rect 4547 1136 4613 1144
rect 4756 1136 4773 1144
rect 4587 1116 4633 1124
rect 4127 1096 4164 1104
rect 4187 1096 4373 1104
rect 4467 1096 4484 1104
rect 3347 1076 3504 1084
rect 3616 1076 4453 1084
rect 916 1056 933 1064
rect 1507 1056 1793 1064
rect 1807 1056 2193 1064
rect 2207 1056 2753 1064
rect 2827 1056 2933 1064
rect 3616 1064 3624 1076
rect 4476 1084 4484 1096
rect 4476 1076 4513 1084
rect 4676 1084 4684 1113
rect 4756 1107 4764 1136
rect 4887 1136 4953 1144
rect 5007 1136 5133 1144
rect 5287 1136 5324 1144
rect 4856 1116 5033 1124
rect 4796 1087 4804 1113
rect 4856 1107 4864 1116
rect 4896 1096 5013 1104
rect 4587 1076 4684 1084
rect 4896 1084 4904 1096
rect 5316 1104 5324 1136
rect 5287 1096 5324 1104
rect 5336 1136 5433 1144
rect 4827 1076 5253 1084
rect 5336 1084 5344 1136
rect 5556 1144 5564 1156
rect 5476 1136 5564 1144
rect 5636 1144 5644 1156
rect 5736 1156 5813 1164
rect 5636 1136 5673 1144
rect 5307 1076 5344 1084
rect 5476 1084 5484 1136
rect 5536 1127 5544 1136
rect 5736 1124 5744 1156
rect 5996 1164 6004 1176
rect 6147 1176 6193 1184
rect 6216 1176 6273 1184
rect 5907 1156 6004 1164
rect 6216 1164 6224 1176
rect 6407 1176 6633 1184
rect 6027 1156 6224 1164
rect 6347 1156 6413 1164
rect 6527 1156 6593 1164
rect 5787 1136 6073 1144
rect 6127 1136 6453 1144
rect 6567 1136 6624 1144
rect 5647 1116 5684 1124
rect 5736 1116 5824 1124
rect 5676 1107 5684 1116
rect 5816 1107 5824 1116
rect 5836 1116 5853 1124
rect 5716 1096 5773 1104
rect 5427 1076 5484 1084
rect 5507 1076 5553 1084
rect 5716 1084 5724 1096
rect 5836 1087 5844 1116
rect 5896 1116 5933 1124
rect 5856 1096 5873 1104
rect 5856 1087 5864 1096
rect 5707 1076 5724 1084
rect 5896 1084 5904 1116
rect 6047 1116 6084 1124
rect 5967 1096 5993 1104
rect 5887 1076 5904 1084
rect 5947 1076 5973 1084
rect 6076 1067 6084 1116
rect 6616 1124 6624 1136
rect 6567 1116 6604 1124
rect 6616 1116 6684 1124
rect 6096 1084 6104 1113
rect 6276 1104 6284 1113
rect 6267 1096 6284 1104
rect 6096 1076 6393 1084
rect 6596 1084 6604 1116
rect 6627 1096 6653 1104
rect 6567 1076 6604 1084
rect 6676 1084 6684 1116
rect 6667 1076 6684 1084
rect 3387 1056 3624 1064
rect 3787 1056 4384 1064
rect 1887 1036 2273 1044
rect 2287 1036 2613 1044
rect 2847 1036 2993 1044
rect 3047 1036 3313 1044
rect 3507 1036 3893 1044
rect 3967 1036 4113 1044
rect 4327 1036 4353 1044
rect 4376 1044 4384 1056
rect 4567 1056 5113 1064
rect 5747 1056 5953 1064
rect 6347 1056 6733 1064
rect 4376 1036 4673 1044
rect 4767 1036 4953 1044
rect 5647 1036 5753 1044
rect 5827 1036 5853 1044
rect 596 1016 613 1024
rect 787 1016 833 1024
rect 1627 1016 2433 1024
rect 2467 1016 2653 1024
rect 2747 1016 3273 1024
rect 3316 1016 3433 1024
rect 2027 996 2513 1004
rect 3007 996 3073 1004
rect 3316 1004 3324 1016
rect 3467 1016 3613 1024
rect 3627 1016 3633 1024
rect 3927 1016 4033 1024
rect 4667 1016 4873 1024
rect 4907 1016 5013 1024
rect 5367 1016 6033 1024
rect 6047 1016 6433 1024
rect 6467 1016 6713 1024
rect 3227 996 3324 1004
rect 3496 996 3713 1004
rect 1707 976 1893 984
rect 1907 976 2013 984
rect 2047 976 2153 984
rect 2247 976 2533 984
rect 3496 984 3504 996
rect 3727 996 4033 1004
rect 4047 996 4513 1004
rect 4867 996 4913 1004
rect 5667 996 6473 1004
rect 2847 976 3504 984
rect 3587 976 4333 984
rect 4467 976 5213 984
rect 5387 976 6113 984
rect 6127 976 6573 984
rect 6587 976 6593 984
rect 6667 976 6713 984
rect 2187 956 2373 964
rect 2447 956 2713 964
rect 2807 956 3093 964
rect 3147 956 3173 964
rect 3207 956 3313 964
rect 3327 956 3393 964
rect 3407 956 3553 964
rect 3567 956 3793 964
rect 3807 956 3853 964
rect 3867 956 4053 964
rect 4187 956 4373 964
rect 4427 956 4513 964
rect 4527 956 4993 964
rect 5007 956 6093 964
rect 6267 956 6473 964
rect 767 936 813 944
rect 1847 936 1873 944
rect 1887 936 1913 944
rect 2276 936 2853 944
rect 687 916 953 924
rect 987 916 1193 924
rect 2276 924 2284 936
rect 2867 936 3373 944
rect 3407 936 3653 944
rect 3927 936 4493 944
rect 4507 936 4653 944
rect 4687 936 4813 944
rect 5007 936 5113 944
rect 5136 936 5233 944
rect 1347 916 2284 924
rect 2307 916 2413 924
rect 2487 916 2533 924
rect 2547 916 2753 924
rect 3127 916 3453 924
rect 3487 916 3613 924
rect 3627 916 3693 924
rect 3967 916 4133 924
rect 4227 916 4313 924
rect 4347 916 4613 924
rect 5136 924 5144 936
rect 5267 936 5653 944
rect 4627 916 5144 924
rect 5187 916 5333 924
rect 5687 916 5833 924
rect 6107 916 6153 924
rect 127 896 433 904
rect 807 896 893 904
rect 1047 896 1233 904
rect 1247 896 1273 904
rect 2347 896 2493 904
rect 2567 896 3973 904
rect 4267 896 4353 904
rect 4416 896 4673 904
rect 147 876 313 884
rect 467 876 493 884
rect 547 876 713 884
rect 727 876 1033 884
rect 2127 876 2593 884
rect 2627 876 3084 884
rect 187 856 204 864
rect 36 827 44 853
rect 196 844 204 856
rect 627 856 653 864
rect 707 856 753 864
rect 887 856 933 864
rect 947 856 1093 864
rect 1367 856 1453 864
rect 1767 856 1873 864
rect 2267 856 2373 864
rect 2427 856 2624 864
rect 196 836 213 844
rect 576 836 593 844
rect 276 816 333 824
rect 276 804 284 816
rect 476 824 484 833
rect 576 827 584 836
rect 356 816 493 824
rect 236 796 284 804
rect 236 784 244 796
rect 356 804 364 816
rect 527 816 544 824
rect 307 796 364 804
rect 227 776 244 784
rect 536 784 544 816
rect 656 824 664 853
rect 836 844 844 853
rect 816 836 844 844
rect 896 836 1073 844
rect 627 816 664 824
rect 747 816 773 824
rect 816 824 824 836
rect 807 816 824 824
rect 896 824 904 836
rect 1267 836 1324 844
rect 887 816 904 824
rect 927 816 953 824
rect 1007 816 1053 824
rect 1147 816 1173 824
rect 1316 824 1324 836
rect 1987 836 2033 844
rect 2396 844 2404 853
rect 2616 847 2624 856
rect 3076 864 3084 876
rect 3107 876 3513 884
rect 3547 876 3573 884
rect 3887 876 4253 884
rect 4416 884 4424 896
rect 4747 896 4793 904
rect 5107 896 5413 904
rect 5447 896 5613 904
rect 5667 896 5693 904
rect 5727 896 6613 904
rect 6627 896 6673 904
rect 4376 876 4424 884
rect 2947 856 3064 864
rect 3076 856 3773 864
rect 2387 836 2404 844
rect 2516 836 2533 844
rect 1316 816 1333 824
rect 1587 816 1633 824
rect 1967 816 1993 824
rect 2356 824 2364 833
rect 2356 816 2393 824
rect 587 796 1233 804
rect 1427 796 1473 804
rect 1696 804 1704 813
rect 1696 796 1733 804
rect 1747 796 1813 804
rect 2107 796 2333 804
rect 2407 796 2433 804
rect 2456 804 2464 833
rect 2516 827 2524 836
rect 2667 836 2793 844
rect 2947 836 2973 844
rect 2987 836 3033 844
rect 2587 816 2633 824
rect 2916 824 2924 833
rect 2916 816 2953 824
rect 3056 824 3064 856
rect 3847 856 4013 864
rect 4376 864 4384 876
rect 4547 876 4613 884
rect 4667 876 4684 884
rect 4236 856 4384 864
rect 3167 836 3253 844
rect 3347 836 3553 844
rect 3596 836 3733 844
rect 3596 827 3604 836
rect 4107 836 4173 844
rect 4236 844 4244 856
rect 4216 836 4244 844
rect 3056 816 3373 824
rect 3616 816 3913 824
rect 2456 796 2533 804
rect 2567 796 2813 804
rect 3007 796 3173 804
rect 3616 804 3624 816
rect 4027 816 4073 824
rect 4216 824 4224 836
rect 4267 836 4293 844
rect 4147 816 4224 824
rect 4247 816 4273 824
rect 4316 824 4324 856
rect 4456 856 4573 864
rect 4396 844 4404 853
rect 4456 844 4464 856
rect 4347 836 4404 844
rect 4436 836 4464 844
rect 4316 816 4393 824
rect 3196 796 3624 804
rect 487 776 753 784
rect 1027 776 1593 784
rect 1607 776 1833 784
rect 1847 776 2073 784
rect 2087 776 2193 784
rect 2207 776 2213 784
rect 2227 776 2313 784
rect 2327 776 2373 784
rect 2387 776 2533 784
rect 2647 776 2673 784
rect 2827 776 2973 784
rect 3196 784 3204 796
rect 3667 796 3713 804
rect 4047 796 4173 804
rect 4187 796 4193 804
rect 4287 796 4313 804
rect 4436 804 4444 836
rect 4507 836 4553 844
rect 4607 836 4653 844
rect 4676 824 4684 876
rect 4767 876 5184 884
rect 4727 856 4873 864
rect 4767 836 4804 844
rect 4667 816 4684 824
rect 4727 816 4773 824
rect 4347 796 4444 804
rect 4487 796 4524 804
rect 2987 776 3204 784
rect 3247 776 3493 784
rect 3567 776 3873 784
rect 3967 776 4233 784
rect 467 756 513 764
rect 527 756 573 764
rect 687 756 833 764
rect 1107 756 1133 764
rect 1887 756 2093 764
rect 2487 756 2573 764
rect 2667 756 2733 764
rect 2767 756 3153 764
rect 3216 756 3533 764
rect 407 736 553 744
rect 567 736 693 744
rect 707 736 953 744
rect 3216 744 3224 756
rect 3687 756 3773 764
rect 3787 756 3793 764
rect 3827 756 4053 764
rect 4087 756 4433 764
rect 4516 764 4524 796
rect 4547 796 4613 804
rect 4627 796 4713 804
rect 4727 796 4733 804
rect 4796 804 4804 836
rect 4847 836 4893 844
rect 5016 836 5113 844
rect 5016 824 5024 836
rect 4987 816 5024 824
rect 5176 824 5184 876
rect 5327 876 5353 884
rect 5667 876 5713 884
rect 5727 876 5873 884
rect 5947 876 6453 884
rect 5207 856 5393 864
rect 5407 856 5573 864
rect 5836 856 5853 864
rect 5287 836 5433 844
rect 5527 836 5573 844
rect 5696 827 5704 853
rect 5836 844 5844 856
rect 6007 856 6244 864
rect 5807 836 5844 844
rect 5887 836 5953 844
rect 6236 844 6244 856
rect 6267 856 6293 864
rect 6327 856 6353 864
rect 6467 856 6533 864
rect 6547 856 6653 864
rect 6087 836 6224 844
rect 6236 836 6293 844
rect 5167 816 5184 824
rect 5307 816 5584 824
rect 4767 796 4804 804
rect 5367 796 5413 804
rect 5427 796 5473 804
rect 5576 804 5584 816
rect 5607 816 5633 824
rect 5756 824 5764 833
rect 5756 816 5784 824
rect 5576 796 5633 804
rect 4547 776 4653 784
rect 4947 776 5033 784
rect 5447 776 5493 784
rect 5627 776 5673 784
rect 5736 784 5744 813
rect 5776 807 5784 816
rect 6036 816 6133 824
rect 6036 804 6044 816
rect 6216 824 6224 836
rect 6347 836 6413 844
rect 6216 816 6233 824
rect 6327 816 6533 824
rect 5927 796 6044 804
rect 6067 796 6433 804
rect 6447 796 6573 804
rect 5736 776 5764 784
rect 4447 756 4524 764
rect 4667 756 4953 764
rect 4967 756 5093 764
rect 5756 764 5764 776
rect 5807 776 6013 784
rect 6227 776 6273 784
rect 5467 756 5764 764
rect 6187 756 6233 764
rect 1867 736 3224 744
rect 3247 736 3484 744
rect 2527 716 2773 724
rect 2927 716 3053 724
rect 3067 716 3333 724
rect 3367 716 3453 724
rect 3476 724 3484 736
rect 3767 736 3933 744
rect 3947 736 3993 744
rect 4387 736 4433 744
rect 4467 736 4713 744
rect 5167 736 5413 744
rect 5427 736 5873 744
rect 5907 736 5933 744
rect 5947 736 6053 744
rect 6327 736 6353 744
rect 3476 716 3853 724
rect 3867 716 3973 724
rect 3987 716 4413 724
rect 4427 716 5153 724
rect 5567 716 5713 724
rect 5867 716 5913 724
rect 5947 716 6153 724
rect 107 696 253 704
rect 1567 696 2513 704
rect 2587 696 2733 704
rect 2787 696 2813 704
rect 2947 696 3053 704
rect 3127 696 3173 704
rect 3307 696 3893 704
rect 4207 696 4253 704
rect 4387 696 4573 704
rect 4727 696 4853 704
rect 5627 696 5673 704
rect 5876 696 5953 704
rect -4 676 13 684
rect -4 644 4 676
rect 207 676 233 684
rect 867 676 913 684
rect 1487 676 1693 684
rect 2507 676 2673 684
rect 2687 676 2833 684
rect 3107 676 3393 684
rect 3927 676 5353 684
rect 5876 684 5884 696
rect 6067 696 6333 704
rect 5367 676 5884 684
rect 5907 676 6193 684
rect 6527 676 6533 684
rect 6547 676 6553 684
rect 27 656 53 664
rect 327 656 373 664
rect 467 656 533 664
rect 716 656 753 664
rect -4 636 24 644
rect 16 627 24 636
rect 67 636 113 644
rect 116 616 133 624
rect 116 607 124 616
rect 47 596 73 604
rect 176 604 184 653
rect 256 627 264 653
rect 307 636 333 644
rect 716 644 724 656
rect 887 656 1353 664
rect 356 636 724 644
rect 356 627 364 636
rect 847 636 973 644
rect 996 627 1004 656
rect 1387 656 1553 664
rect 2156 664 2164 673
rect 2156 656 2633 664
rect 2716 656 2873 664
rect 1287 636 1313 644
rect 1487 636 1793 644
rect 2467 636 2493 644
rect 2716 627 2724 656
rect 3027 656 3093 664
rect 3107 656 3193 664
rect 3207 656 3333 664
rect 3347 656 3353 664
rect 3367 656 3413 664
rect 3727 656 3764 664
rect 2787 636 2904 644
rect 2896 627 2904 636
rect 2936 627 2944 653
rect 2956 644 2964 653
rect 2956 636 3004 644
rect 467 616 544 624
rect 147 596 184 604
rect 207 596 233 604
rect 247 596 353 604
rect 416 587 424 613
rect 536 607 544 616
rect 567 616 584 624
rect 576 604 584 616
rect 607 616 633 624
rect 687 616 713 624
rect 727 616 733 624
rect 2767 616 2813 624
rect 2996 624 3004 636
rect 3167 636 3433 644
rect 3607 636 3624 644
rect 2996 616 3024 624
rect 3016 607 3024 616
rect 3327 616 3373 624
rect 3427 616 3473 624
rect 3496 607 3504 633
rect 3616 624 3624 636
rect 3647 636 3664 644
rect 3656 627 3664 636
rect 3616 616 3644 624
rect 576 596 593 604
rect 636 596 653 604
rect 287 556 413 564
rect 436 564 444 593
rect 636 587 644 596
rect 787 596 853 604
rect 867 596 893 604
rect 1687 596 2013 604
rect 2107 596 2253 604
rect 2327 596 2393 604
rect 2407 596 2853 604
rect 3347 596 3453 604
rect 3636 604 3644 616
rect 3716 604 3724 633
rect 3756 624 3764 656
rect 3907 656 3944 664
rect 3936 647 3944 656
rect 4027 656 4333 664
rect 4367 656 4473 664
rect 4627 656 4693 664
rect 4747 656 4753 664
rect 4767 656 4833 664
rect 4887 656 4913 664
rect 5867 656 6113 664
rect 6187 656 6393 664
rect 6587 656 6653 664
rect 4267 636 4353 644
rect 4547 636 4584 644
rect 3747 616 3764 624
rect 3887 616 4453 624
rect 4507 616 4553 624
rect 3636 596 3724 604
rect 3776 604 3784 613
rect 3767 596 3784 604
rect 3807 596 4193 604
rect 4576 604 4584 636
rect 4636 636 4673 644
rect 4636 624 4644 636
rect 4736 636 4793 644
rect 4736 627 4744 636
rect 4816 636 4904 644
rect 4816 627 4824 636
rect 4607 616 4644 624
rect 4896 624 4904 636
rect 4896 616 4953 624
rect 4976 624 4984 653
rect 5027 636 5053 644
rect 5096 636 5144 644
rect 5076 624 5084 633
rect 5096 627 5104 636
rect 4976 616 5084 624
rect 4576 596 4693 604
rect 4767 596 4853 604
rect 4907 596 5013 604
rect 5027 596 5053 604
rect 5076 604 5084 616
rect 5136 624 5144 636
rect 5307 636 5353 644
rect 5547 636 5584 644
rect 5136 616 5333 624
rect 5347 616 5513 624
rect 5076 596 5093 604
rect 5116 604 5124 613
rect 5107 596 5124 604
rect 5576 604 5584 636
rect 5796 636 5853 644
rect 5547 596 5584 604
rect 5596 604 5604 633
rect 5796 624 5804 636
rect 5927 636 5973 644
rect 6087 636 6133 644
rect 6156 636 6193 644
rect 5727 616 5804 624
rect 5916 624 5924 633
rect 6156 627 6164 636
rect 6227 636 6253 644
rect 5907 616 5924 624
rect 6056 616 6093 624
rect 5596 596 5693 604
rect 5707 596 5713 604
rect 567 576 613 584
rect 807 576 833 584
rect 1547 576 3384 584
rect 436 556 573 564
rect 587 556 933 564
rect 3027 556 3173 564
rect 3376 564 3384 576
rect 3407 576 4244 584
rect 3376 556 3673 564
rect 3767 556 3833 564
rect 4236 564 4244 576
rect 5447 576 5573 584
rect 5956 584 5964 613
rect 6056 604 6064 616
rect 6207 616 6273 624
rect 6327 616 6513 624
rect 6536 616 6573 624
rect 5987 596 6064 604
rect 6536 604 6544 616
rect 6407 596 6544 604
rect 5956 576 6033 584
rect 6236 584 6244 593
rect 6047 576 6244 584
rect 6267 576 6373 584
rect 4236 556 4493 564
rect 4527 556 5433 564
rect 5467 556 5633 564
rect 5647 556 5933 564
rect 5947 556 6053 564
rect 327 536 553 544
rect 647 536 913 544
rect 2987 536 3053 544
rect 3627 536 4173 544
rect 4476 536 4973 544
rect 407 516 473 524
rect 2247 516 2293 524
rect 3647 516 3713 524
rect 3747 516 4073 524
rect 4476 524 4484 536
rect 5147 536 5273 544
rect 5287 536 5473 544
rect 4087 516 4484 524
rect 4507 516 4873 524
rect 4947 516 5033 524
rect 5107 516 5233 524
rect 2747 496 3253 504
rect 3487 496 3573 504
rect 3947 496 4013 504
rect 4167 496 4293 504
rect 4767 496 6113 504
rect 2507 476 2553 484
rect 2567 476 3033 484
rect 3427 476 3713 484
rect 3727 476 4153 484
rect 4167 476 4473 484
rect 4487 476 5253 484
rect 5267 476 5493 484
rect 5507 476 5793 484
rect 5807 476 5893 484
rect 6127 476 6373 484
rect 6387 476 6593 484
rect 67 456 393 464
rect 1707 456 3393 464
rect 3447 456 3853 464
rect 4347 456 4513 464
rect 4527 456 4553 464
rect 5167 456 5233 464
rect 5907 456 5953 464
rect 6467 456 6513 464
rect 3076 436 4493 444
rect 467 416 513 424
rect 3076 424 3084 436
rect 5067 436 5353 444
rect 5447 436 6053 444
rect 6287 436 6333 444
rect 1767 416 3084 424
rect 3107 416 3484 424
rect 687 396 753 404
rect 1407 396 1453 404
rect 1907 396 2133 404
rect 2207 396 2264 404
rect 267 376 513 384
rect 576 376 853 384
rect 467 356 493 364
rect 576 364 584 376
rect 1567 376 1613 384
rect 2147 376 2173 384
rect 547 356 584 364
rect 696 356 764 364
rect 696 347 704 356
rect 16 336 153 344
rect 16 327 24 336
rect 756 344 764 356
rect 796 356 833 364
rect 796 344 804 356
rect 847 356 853 364
rect 756 336 804 344
rect 1227 336 1273 344
rect 1287 336 1293 344
rect 127 316 373 324
rect 387 316 473 324
rect 787 316 1133 324
rect 587 296 633 304
rect 687 296 733 304
rect 1436 304 1444 373
rect 1476 347 1484 373
rect 2027 356 2073 364
rect 2096 347 2104 373
rect 2216 364 2224 373
rect 2207 356 2224 364
rect 1647 336 1673 344
rect 2176 344 2184 353
rect 2176 336 2213 344
rect 1507 316 1553 324
rect 1627 316 1653 324
rect 2236 324 2244 353
rect 2256 344 2264 396
rect 3327 396 3464 404
rect 2407 376 2753 384
rect 2767 376 2793 384
rect 2827 376 2933 384
rect 2976 376 2993 384
rect 2287 356 2333 364
rect 2976 364 2984 376
rect 2727 356 2984 364
rect 3207 356 3273 364
rect 3456 364 3464 396
rect 3436 356 3464 364
rect 2256 336 2293 344
rect 2447 336 2513 344
rect 2747 336 2773 344
rect 3436 344 3444 356
rect 3416 336 3444 344
rect 3416 327 3424 336
rect 3476 344 3484 416
rect 3587 416 3753 424
rect 3767 416 4133 424
rect 4147 416 5133 424
rect 5207 416 5453 424
rect 5627 416 5673 424
rect 5707 416 5733 424
rect 5747 416 5813 424
rect 6147 416 6313 424
rect 3567 396 3633 404
rect 3687 396 3913 404
rect 4407 396 4953 404
rect 4987 396 5173 404
rect 5347 396 5433 404
rect 6247 396 6293 404
rect 3527 376 3533 384
rect 3547 376 3733 384
rect 3807 376 3904 384
rect 3507 356 3544 364
rect 3467 336 3484 344
rect 3536 344 3544 356
rect 3536 336 3564 344
rect 3556 327 3564 336
rect 3656 344 3664 353
rect 3647 336 3664 344
rect 3776 344 3784 373
rect 3867 356 3884 364
rect 3876 347 3884 356
rect 3896 347 3904 376
rect 3947 376 3964 384
rect 3956 367 3964 376
rect 4447 376 4753 384
rect 4516 367 4524 376
rect 5247 376 5304 384
rect 5296 367 5304 376
rect 5427 376 5564 384
rect 3927 356 3944 364
rect 3776 336 3804 344
rect 3796 327 3804 336
rect 3936 344 3944 356
rect 3987 356 4033 364
rect 4676 356 4713 364
rect 3936 336 3953 344
rect 4176 336 4193 344
rect 2236 316 2353 324
rect 2367 316 2433 324
rect 2687 316 2853 324
rect 2887 316 2933 324
rect 3507 316 3533 324
rect 3747 316 3773 324
rect 4176 324 4184 336
rect 4507 336 4573 344
rect 4676 344 4684 356
rect 5067 356 5104 364
rect 4636 336 4684 344
rect 4836 336 4933 344
rect 4087 316 4184 324
rect 4307 316 4553 324
rect 4636 324 4644 336
rect 4627 316 4644 324
rect 4836 324 4844 336
rect 5096 344 5104 356
rect 5316 347 5324 373
rect 5356 347 5364 373
rect 5556 364 5564 376
rect 5627 376 5724 384
rect 5716 367 5724 376
rect 5987 376 6004 384
rect 5996 367 6004 376
rect 6016 376 6033 384
rect 5556 356 5593 364
rect 5807 356 5853 364
rect 5096 336 5113 344
rect 5527 336 5653 344
rect 5827 336 5873 344
rect 5927 336 5973 344
rect 6016 344 6024 376
rect 6547 376 6613 384
rect 6067 356 6133 364
rect 5996 336 6024 344
rect 4787 316 4844 324
rect 5056 324 5064 333
rect 4987 316 5064 324
rect 5076 316 5153 324
rect 1407 296 1444 304
rect 2047 296 2313 304
rect 2347 296 2613 304
rect 2667 296 3053 304
rect 3067 296 3393 304
rect 3407 296 3533 304
rect 3607 296 3753 304
rect 3907 296 3993 304
rect 4007 296 4273 304
rect 4287 296 4393 304
rect 4407 296 4413 304
rect 4587 296 4993 304
rect 5076 304 5084 316
rect 5407 316 5433 324
rect 5996 324 6004 336
rect 6256 344 6264 353
rect 6316 347 6324 373
rect 6256 336 6284 344
rect 5967 316 6004 324
rect 6156 324 6164 333
rect 6276 327 6284 336
rect 6067 316 6233 324
rect 6336 324 6344 353
rect 6396 347 6404 373
rect 6427 336 6493 344
rect 6327 316 6344 324
rect 5007 296 5084 304
rect 5107 296 5993 304
rect 6147 296 6213 304
rect 6247 296 6473 304
rect 1127 276 1713 284
rect 1727 276 1753 284
rect 1787 276 2253 284
rect 2867 276 3073 284
rect 3087 276 3353 284
rect 3867 276 3953 284
rect 4247 276 4524 284
rect 2307 256 2453 264
rect 2607 256 2793 264
rect 3027 256 3293 264
rect 3387 256 3413 264
rect 3547 256 3893 264
rect 3947 256 4313 264
rect 4516 264 4524 276
rect 4547 276 4693 284
rect 4887 276 5324 284
rect 4516 256 4633 264
rect 4667 256 4833 264
rect 4847 256 4973 264
rect 5027 256 5253 264
rect 5316 264 5324 276
rect 5347 276 5753 284
rect 5767 276 6093 284
rect 6107 276 6273 284
rect 5316 256 5473 264
rect 5487 256 5933 264
rect 6087 256 6153 264
rect 6267 256 6313 264
rect 1227 236 1533 244
rect 2207 236 2373 244
rect 2847 236 3093 244
rect 3247 236 3513 244
rect 3527 236 4293 244
rect 4307 236 4813 244
rect 4827 236 5333 244
rect 5947 236 6713 244
rect 827 216 873 224
rect 887 216 1133 224
rect 1147 216 1153 224
rect 1167 216 1213 224
rect 1347 216 1593 224
rect 1607 216 2053 224
rect 2067 216 2093 224
rect 2107 216 2353 224
rect 2367 216 2513 224
rect 2527 216 2593 224
rect 3347 216 3573 224
rect 3647 216 3933 224
rect 4187 216 4213 224
rect 4267 216 4593 224
rect 4607 216 5193 224
rect 5207 216 5373 224
rect 6127 216 6193 224
rect 567 196 573 204
rect 587 196 653 204
rect 727 196 973 204
rect 1267 196 1433 204
rect 1447 196 1693 204
rect 1707 196 1753 204
rect 1767 196 1833 204
rect 1847 196 1913 204
rect 2587 196 2653 204
rect 2667 196 2893 204
rect 2907 196 2993 204
rect 3036 196 3113 204
rect 127 176 353 184
rect 367 176 833 184
rect 847 176 1173 184
rect 1187 176 1353 184
rect 1467 176 1513 184
rect 1567 176 1793 184
rect 1987 176 2224 184
rect 167 156 273 164
rect 576 156 613 164
rect 576 124 584 156
rect 667 156 713 164
rect 727 156 753 164
rect 767 156 953 164
rect 1187 156 1313 164
rect 1607 156 1653 164
rect 1947 156 2013 164
rect 2067 156 2193 164
rect 2216 164 2224 176
rect 2247 176 2644 184
rect 2216 156 2313 164
rect 2327 156 2333 164
rect 2567 156 2613 164
rect 2636 164 2644 176
rect 2736 176 2793 184
rect 2736 164 2744 176
rect 3036 184 3044 196
rect 3167 196 3413 204
rect 3627 196 3653 204
rect 3887 196 4093 204
rect 4187 196 4453 204
rect 4627 196 5093 204
rect 5827 196 5973 204
rect 6187 196 6233 204
rect 6307 196 6393 204
rect 6407 196 6413 204
rect 3016 176 3044 184
rect 2636 156 2744 164
rect 3016 164 3024 176
rect 3067 176 3084 184
rect 2967 156 3024 164
rect 3076 164 3084 176
rect 3607 176 3664 184
rect 3076 156 3104 164
rect 1107 136 1153 144
rect 1207 136 1493 144
rect 1536 127 1544 153
rect 1567 136 1633 144
rect 1687 136 1733 144
rect 1756 136 1873 144
rect 576 116 593 124
rect 647 116 853 124
rect 1756 124 1764 136
rect 1967 136 2033 144
rect 2356 127 2364 153
rect 2387 136 2413 144
rect 2487 136 2533 144
rect 2587 136 2633 144
rect 3096 144 3104 156
rect 3567 156 3593 164
rect 3627 156 3644 164
rect 3096 136 3133 144
rect 3567 136 3613 144
rect 1627 116 1764 124
rect 2027 116 2073 124
rect 2627 116 2733 124
rect 2907 116 3493 124
rect 3636 124 3644 156
rect 3656 144 3664 176
rect 3767 176 4093 184
rect 4107 176 4613 184
rect 4707 176 4973 184
rect 5196 176 5213 184
rect 3687 156 3733 164
rect 4087 156 4133 164
rect 4227 156 4333 164
rect 4607 156 4653 164
rect 5127 156 5173 164
rect 5196 147 5204 176
rect 5236 176 5444 184
rect 5236 164 5244 176
rect 5227 156 5244 164
rect 5267 156 5373 164
rect 5436 164 5444 176
rect 5467 176 5693 184
rect 5707 176 5933 184
rect 5947 176 6513 184
rect 5436 156 5493 164
rect 5567 156 5613 164
rect 5767 156 5853 164
rect 5967 156 6133 164
rect 6187 156 6253 164
rect 6307 156 6364 164
rect 3656 136 3704 144
rect 3636 116 3653 124
rect 3696 124 3704 136
rect 3727 136 3793 144
rect 3807 136 4053 144
rect 4127 136 4153 144
rect 4207 136 4253 144
rect 4727 136 4773 144
rect 5247 136 5293 144
rect 6007 136 6113 144
rect 6207 136 6313 144
rect 6356 144 6364 156
rect 6516 156 6553 164
rect 6516 144 6524 156
rect 6356 136 6524 144
rect 3696 116 3813 124
rect 4447 116 4673 124
rect 5147 116 5653 124
rect 6167 116 6213 124
rect 1007 96 1593 104
rect 2127 96 2413 104
rect 2447 96 2913 104
rect 2927 96 3173 104
rect 3187 96 4513 104
rect 4587 96 5133 104
rect 6247 96 6273 104
rect 2347 76 3773 84
rect 3787 76 4013 84
rect 4387 76 4753 84
rect 4767 76 4853 84
rect 4067 56 4573 64
rect 4647 56 6053 64
rect 2787 36 2973 44
rect 2987 36 4313 44
rect 1007 16 1033 24
<< m1p >>
rect 4 6482 6716 6498
rect 4 6242 6736 6258
rect 4 6002 6676 6018
rect 4 5762 6736 5778
rect 4 5522 6696 5538
rect 4 5282 6736 5298
rect 4 5042 6736 5058
rect 4 4802 6736 4818
rect 4 4562 6696 4578
rect 4 4322 6736 4338
rect 4 4082 6736 4098
rect 4 3842 6736 3858
rect 4 3602 6716 3618
rect 4 3362 6736 3378
rect 4 3122 6736 3138
rect 4 2882 6736 2898
rect 4 2642 6696 2658
rect 4 2402 6736 2418
rect 4 2162 6716 2178
rect 4 1922 6736 1938
rect 4 1682 6696 1698
rect 4 1442 6736 1458
rect 4 1202 6716 1218
rect 4 962 6736 978
rect 4 722 6696 738
rect 4 482 6736 498
rect 4 242 6656 258
rect 4 2 6736 18
<< m2p >>
rect 833 6413 847 6427
rect 1053 6413 1067 6427
rect 1673 6413 1687 6427
rect 2273 6413 2287 6427
rect 2433 6413 2447 6427
rect 2493 6413 2507 6427
rect 3153 6413 3167 6427
rect 3213 6413 3227 6427
rect 3253 6413 3267 6427
rect 3493 6413 3507 6427
rect 3593 6413 3607 6427
rect 3933 6413 3947 6427
rect 4553 6413 4567 6427
rect 4633 6413 4647 6427
rect 4733 6413 4747 6427
rect 5433 6413 5447 6427
rect 5573 6413 5587 6427
rect 5653 6413 5667 6427
rect 5693 6413 5707 6427
rect 5933 6413 5947 6427
rect 6013 6413 6027 6427
rect 6093 6413 6107 6427
rect 6293 6413 6307 6427
rect 6533 6413 6547 6427
rect 93 6393 107 6407
rect 133 6393 147 6407
rect 213 6393 227 6407
rect 293 6393 307 6407
rect 333 6393 347 6407
rect 613 6393 627 6407
rect 693 6393 707 6407
rect 733 6393 747 6407
rect 893 6393 907 6407
rect 933 6393 947 6407
rect 973 6393 987 6407
rect 1093 6393 1107 6407
rect 1173 6393 1187 6407
rect 1213 6393 1227 6407
rect 1313 6393 1327 6407
rect 1353 6393 1367 6407
rect 1393 6393 1407 6407
rect 1473 6393 1487 6407
rect 1513 6393 1527 6407
rect 1553 6393 1567 6407
rect 1613 6393 1627 6407
rect 1713 6393 1727 6407
rect 1793 6393 1807 6407
rect 1833 6393 1847 6407
rect 1933 6393 1947 6407
rect 1973 6393 1987 6407
rect 2153 6393 2167 6407
rect 2193 6393 2207 6407
rect 2233 6393 2247 6407
rect 2413 6393 2427 6407
rect 2453 6393 2467 6407
rect 2473 6393 2487 6407
rect 2513 6393 2527 6407
rect 2953 6393 2967 6407
rect 2993 6393 3007 6407
rect 3053 6393 3067 6407
rect 3093 6393 3107 6407
rect 3293 6393 3307 6407
rect 3333 6393 3347 6407
rect 3373 6393 3387 6407
rect 3453 6393 3467 6407
rect 3553 6393 3567 6407
rect 3773 6393 3787 6407
rect 3813 6393 3827 6407
rect 3833 6393 3847 6407
rect 3873 6393 3887 6407
rect 4093 6393 4107 6407
rect 4153 6393 4167 6407
rect 4673 6393 4687 6407
rect 4773 6393 4787 6407
rect 4813 6393 4827 6407
rect 4853 6393 4867 6407
rect 4953 6393 4967 6407
rect 4993 6393 5007 6407
rect 5013 6393 5027 6407
rect 5053 6393 5067 6407
rect 5473 6393 5487 6407
rect 5533 6393 5547 6407
rect 5733 6393 5747 6407
rect 5893 6393 5907 6407
rect 6053 6393 6067 6407
rect 6173 6393 6187 6407
rect 6213 6393 6227 6407
rect 6253 6393 6267 6407
rect 6593 6393 6607 6407
rect 6633 6393 6647 6407
rect 6673 6393 6687 6407
rect 273 6373 287 6387
rect 313 6373 327 6387
rect 373 6373 387 6387
rect 473 6373 487 6387
rect 533 6373 547 6387
rect 853 6373 867 6387
rect 913 6373 927 6387
rect 953 6373 967 6387
rect 1033 6373 1047 6387
rect 1333 6373 1347 6387
rect 1373 6373 1387 6387
rect 1453 6373 1467 6387
rect 1493 6373 1507 6387
rect 1653 6373 1667 6387
rect 1953 6373 1967 6387
rect 1993 6373 2007 6387
rect 2053 6373 2067 6387
rect 2133 6373 2147 6387
rect 2173 6373 2187 6387
rect 2253 6373 2267 6387
rect 2293 6373 2307 6387
rect 2353 6373 2367 6387
rect 2573 6373 2587 6387
rect 2673 6373 2687 6387
rect 2713 6373 2727 6387
rect 2753 6373 2767 6387
rect 2853 6373 2867 6387
rect 2893 6373 2907 6387
rect 2933 6373 2947 6387
rect 2973 6373 2987 6387
rect 3033 6373 3047 6387
rect 3073 6373 3087 6387
rect 3133 6373 3147 6387
rect 3193 6373 3207 6387
rect 3233 6373 3247 6387
rect 3273 6373 3287 6387
rect 3353 6373 3367 6387
rect 3393 6373 3407 6387
rect 3473 6373 3487 6387
rect 3513 6373 3527 6387
rect 3573 6373 3587 6387
rect 3613 6373 3627 6387
rect 3633 6373 3647 6387
rect 3673 6373 3687 6387
rect 3753 6373 3767 6387
rect 3793 6373 3807 6387
rect 3853 6373 3867 6387
rect 3893 6373 3907 6387
rect 3953 6373 3967 6387
rect 4013 6373 4027 6387
rect 4193 6373 4207 6387
rect 4293 6373 4307 6387
rect 4333 6373 4347 6387
rect 4393 6373 4407 6387
rect 4433 6373 4447 6387
rect 4493 6373 4507 6387
rect 4533 6373 4547 6387
rect 4573 6373 4587 6387
rect 4613 6373 4627 6387
rect 4653 6373 4667 6387
rect 4713 6373 4727 6387
rect 4753 6373 4767 6387
rect 4833 6373 4847 6387
rect 4873 6373 4887 6387
rect 4933 6373 4947 6387
rect 4973 6373 4987 6387
rect 5033 6373 5047 6387
rect 5073 6373 5087 6387
rect 5153 6373 5167 6387
rect 5193 6373 5207 6387
rect 5253 6373 5267 6387
rect 5293 6373 5307 6387
rect 5353 6373 5367 6387
rect 5393 6373 5407 6387
rect 5413 6373 5427 6387
rect 5453 6373 5467 6387
rect 5553 6373 5567 6387
rect 5593 6373 5607 6387
rect 5633 6373 5647 6387
rect 5673 6373 5687 6387
rect 5713 6373 5727 6387
rect 5773 6373 5787 6387
rect 5813 6373 5827 6387
rect 5913 6373 5927 6387
rect 5953 6373 5967 6387
rect 5993 6373 6007 6387
rect 6073 6373 6087 6387
rect 6113 6373 6127 6387
rect 6153 6373 6167 6387
rect 6193 6373 6207 6387
rect 6273 6373 6287 6387
rect 6313 6373 6327 6387
rect 6333 6373 6347 6387
rect 6373 6373 6387 6387
rect 6473 6373 6487 6387
rect 6513 6373 6527 6387
rect 6553 6373 6567 6387
rect 6613 6373 6627 6387
rect 6653 6373 6667 6387
rect 353 6353 367 6367
rect 393 6353 407 6367
rect 453 6353 467 6367
rect 493 6353 507 6367
rect 513 6353 527 6367
rect 553 6353 567 6367
rect 1573 6353 1587 6367
rect 2033 6353 2047 6367
rect 2073 6353 2087 6367
rect 2333 6353 2347 6367
rect 2373 6353 2387 6367
rect 2553 6353 2567 6367
rect 2593 6353 2607 6367
rect 2653 6353 2667 6367
rect 2693 6353 2707 6367
rect 2733 6353 2747 6367
rect 2773 6353 2787 6367
rect 2833 6353 2847 6367
rect 2873 6353 2887 6367
rect 3653 6353 3667 6367
rect 3693 6353 3707 6367
rect 3993 6353 4007 6367
rect 4033 6353 4047 6367
rect 4113 6353 4127 6367
rect 4173 6353 4187 6367
rect 4213 6353 4227 6367
rect 4273 6353 4287 6367
rect 4313 6353 4327 6367
rect 4373 6353 4387 6367
rect 4413 6353 4427 6367
rect 4473 6353 4487 6367
rect 4513 6353 4527 6367
rect 5133 6353 5147 6367
rect 5173 6353 5187 6367
rect 5233 6353 5247 6367
rect 5273 6353 5287 6367
rect 5333 6353 5347 6367
rect 5373 6353 5387 6367
rect 5793 6353 5807 6367
rect 5833 6353 5847 6367
rect 6353 6353 6367 6367
rect 6393 6353 6407 6367
rect 6453 6353 6467 6367
rect 6493 6353 6507 6367
rect 373 6133 387 6147
rect 413 6133 427 6147
rect 533 6133 547 6147
rect 573 6133 587 6147
rect 2413 6133 2427 6147
rect 2453 6133 2467 6147
rect 2693 6133 2707 6147
rect 2733 6133 2747 6147
rect 2973 6133 2987 6147
rect 3013 6133 3027 6147
rect 3173 6133 3187 6147
rect 3213 6133 3227 6147
rect 3433 6133 3447 6147
rect 3473 6133 3487 6147
rect 3533 6133 3547 6147
rect 3573 6133 3587 6147
rect 3793 6133 3807 6147
rect 3833 6133 3847 6147
rect 3853 6133 3867 6147
rect 3893 6133 3907 6147
rect 4293 6133 4307 6147
rect 4333 6133 4347 6147
rect 4393 6133 4407 6147
rect 4673 6133 4687 6147
rect 4713 6133 4727 6147
rect 4873 6133 4887 6147
rect 4913 6133 4927 6147
rect 4973 6133 4987 6147
rect 5013 6133 5027 6147
rect 5173 6133 5187 6147
rect 5213 6133 5227 6147
rect 5273 6133 5287 6147
rect 5553 6133 5567 6147
rect 5593 6133 5607 6147
rect 5653 6133 5667 6147
rect 5693 6133 5707 6147
rect 5853 6133 5867 6147
rect 5893 6133 5907 6147
rect 6153 6133 6167 6147
rect 6193 6133 6207 6147
rect 6253 6133 6267 6147
rect 6293 6133 6307 6147
rect 6353 6133 6367 6147
rect 6393 6133 6407 6147
rect 293 6113 307 6127
rect 333 6113 347 6127
rect 393 6113 407 6127
rect 553 6113 567 6127
rect 613 6113 627 6127
rect 653 6113 667 6127
rect 713 6113 727 6127
rect 753 6113 767 6127
rect 913 6113 927 6127
rect 953 6113 967 6127
rect 1033 6113 1047 6127
rect 1093 6113 1107 6127
rect 1233 6113 1247 6127
rect 1273 6113 1287 6127
rect 1333 6113 1347 6127
rect 1393 6113 1407 6127
rect 1613 6113 1627 6127
rect 1833 6113 1847 6127
rect 1873 6113 1887 6127
rect 1933 6113 1947 6127
rect 2013 6113 2027 6127
rect 2053 6113 2067 6127
rect 2093 6113 2107 6127
rect 2153 6113 2167 6127
rect 2193 6113 2207 6127
rect 2253 6113 2267 6127
rect 2313 6113 2327 6127
rect 2353 6113 2367 6127
rect 2433 6113 2447 6127
rect 2473 6113 2487 6127
rect 2533 6113 2547 6127
rect 2573 6113 2587 6127
rect 2713 6113 2727 6127
rect 2753 6113 2767 6127
rect 2813 6113 2827 6127
rect 2853 6113 2867 6127
rect 2913 6113 2927 6127
rect 2953 6113 2967 6127
rect 2993 6113 3007 6127
rect 3093 6113 3107 6127
rect 3133 6113 3147 6127
rect 3193 6113 3207 6127
rect 3233 6113 3247 6127
rect 3293 6113 3307 6127
rect 3333 6113 3347 6127
rect 3373 6113 3387 6127
rect 3453 6113 3467 6127
rect 3493 6113 3507 6127
rect 3513 6113 3527 6127
rect 3553 6113 3567 6127
rect 3633 6113 3647 6127
rect 3673 6113 3687 6127
rect 3713 6113 3727 6127
rect 3813 6113 3827 6127
rect 3873 6113 3887 6127
rect 3953 6113 3967 6127
rect 3993 6113 4007 6127
rect 4053 6113 4067 6127
rect 4093 6113 4107 6127
rect 4233 6113 4247 6127
rect 4313 6113 4327 6127
rect 4473 6113 4487 6127
rect 4513 6113 4527 6127
rect 4593 6113 4607 6127
rect 4633 6113 4647 6127
rect 4653 6113 4667 6127
rect 4693 6113 4707 6127
rect 4793 6113 4807 6127
rect 4833 6113 4847 6127
rect 4893 6113 4907 6127
rect 4933 6113 4947 6127
rect 4953 6113 4967 6127
rect 4993 6113 5007 6127
rect 5073 6113 5087 6127
rect 5113 6113 5127 6127
rect 5193 6113 5207 6127
rect 5353 6113 5367 6127
rect 5393 6113 5407 6127
rect 5473 6113 5487 6127
rect 5513 6113 5527 6127
rect 5573 6113 5587 6127
rect 5613 6113 5627 6127
rect 5633 6113 5647 6127
rect 5673 6113 5687 6127
rect 5773 6113 5787 6127
rect 5813 6113 5827 6127
rect 5833 6113 5847 6127
rect 5873 6113 5887 6127
rect 5953 6113 5967 6127
rect 5993 6113 6007 6127
rect 6053 6113 6067 6127
rect 6093 6113 6107 6127
rect 6133 6113 6147 6127
rect 6173 6113 6187 6127
rect 6233 6113 6247 6127
rect 6273 6113 6287 6127
rect 6373 6113 6387 6127
rect 6413 6113 6427 6127
rect 6473 6113 6487 6127
rect 6513 6113 6527 6127
rect 6553 6113 6567 6127
rect 6613 6113 6627 6127
rect 33 6093 47 6107
rect 113 6093 127 6107
rect 153 6093 167 6107
rect 273 6093 287 6107
rect 433 6093 447 6107
rect 473 6093 487 6107
rect 593 6093 607 6107
rect 633 6093 647 6107
rect 733 6093 747 6107
rect 773 6093 787 6107
rect 793 6093 807 6107
rect 833 6093 847 6107
rect 893 6093 907 6107
rect 993 6093 1007 6107
rect 1133 6093 1147 6107
rect 1173 6093 1187 6107
rect 1253 6093 1267 6107
rect 1293 6093 1307 6107
rect 1433 6093 1447 6107
rect 1473 6093 1487 6107
rect 1513 6093 1527 6107
rect 1553 6093 1567 6107
rect 1653 6093 1667 6107
rect 1693 6093 1707 6107
rect 1733 6093 1747 6107
rect 1773 6093 1787 6107
rect 1813 6093 1827 6107
rect 1853 6093 1867 6107
rect 1993 6093 2007 6107
rect 2173 6093 2187 6107
rect 2213 6093 2227 6107
rect 2333 6093 2347 6107
rect 2373 6093 2387 6107
rect 2513 6093 2527 6107
rect 2613 6093 2627 6107
rect 2653 6093 2667 6107
rect 2793 6093 2807 6107
rect 2833 6093 2847 6107
rect 2873 6093 2887 6107
rect 3073 6093 3087 6107
rect 3273 6093 3287 6107
rect 3733 6093 3747 6107
rect 3973 6093 3987 6107
rect 4013 6093 4027 6107
rect 4033 6093 4047 6107
rect 4073 6093 4087 6107
rect 4153 6093 4167 6107
rect 4193 6093 4207 6107
rect 4353 6093 4367 6107
rect 4413 6093 4427 6107
rect 4493 6093 4507 6107
rect 4533 6093 4547 6107
rect 4573 6093 4587 6107
rect 4773 6093 4787 6107
rect 5093 6093 5107 6107
rect 5133 6093 5147 6107
rect 5233 6093 5247 6107
rect 5293 6093 5307 6107
rect 5333 6093 5347 6107
rect 5373 6093 5387 6107
rect 5453 6093 5467 6107
rect 5753 6093 5767 6107
rect 5933 6093 5947 6107
rect 5973 6093 5987 6107
rect 6033 6093 6047 6107
rect 6073 6093 6087 6107
rect 6453 6093 6467 6107
rect 313 6073 327 6087
rect 453 6073 467 6087
rect 813 6073 827 6087
rect 933 6073 947 6087
rect 973 6073 987 6087
rect 1113 6073 1127 6087
rect 1153 6073 1167 6087
rect 1353 6073 1367 6087
rect 1413 6073 1427 6087
rect 1453 6073 1467 6087
rect 1533 6073 1547 6087
rect 1593 6073 1607 6087
rect 1673 6073 1687 6087
rect 1753 6073 1767 6087
rect 1913 6073 1927 6087
rect 2033 6073 2047 6087
rect 2073 6073 2087 6087
rect 2233 6073 2247 6087
rect 2553 6073 2567 6087
rect 2633 6073 2647 6087
rect 2933 6073 2947 6087
rect 3113 6073 3127 6087
rect 3313 6073 3327 6087
rect 3393 6073 3407 6087
rect 3613 6073 3627 6087
rect 3693 6073 3707 6087
rect 4173 6073 4187 6087
rect 4213 6073 4227 6087
rect 4613 6073 4627 6087
rect 4813 6073 4827 6087
rect 5493 6073 5507 6087
rect 5793 6073 5807 6087
rect 6493 6073 6507 6087
rect 6533 6073 6547 6087
rect 6593 6073 6607 6087
rect 313 5933 327 5947
rect 433 5933 447 5947
rect 533 5933 547 5947
rect 593 5933 607 5947
rect 793 5933 807 5947
rect 833 5933 847 5947
rect 1093 5933 1107 5947
rect 1193 5933 1207 5947
rect 1773 5933 1787 5947
rect 1913 5933 1927 5947
rect 2233 5933 2247 5947
rect 2613 5933 2627 5947
rect 3493 5933 3507 5947
rect 3753 5933 3767 5947
rect 3993 5933 4007 5947
rect 4193 5933 4207 5947
rect 4553 5933 4567 5947
rect 4753 5933 4767 5947
rect 4913 5933 4927 5947
rect 5053 5933 5067 5947
rect 5533 5933 5547 5947
rect 5713 5933 5727 5947
rect 33 5913 47 5927
rect 73 5913 87 5927
rect 273 5913 287 5927
rect 513 5913 527 5927
rect 553 5913 567 5927
rect 573 5913 587 5927
rect 613 5913 627 5927
rect 653 5913 667 5927
rect 693 5913 707 5927
rect 813 5913 827 5927
rect 853 5913 867 5927
rect 1013 5913 1027 5927
rect 1053 5913 1067 5927
rect 1073 5913 1087 5927
rect 1113 5913 1127 5927
rect 1233 5913 1247 5927
rect 1313 5913 1327 5927
rect 1353 5913 1367 5927
rect 1673 5913 1687 5927
rect 1713 5913 1727 5927
rect 1753 5913 1767 5927
rect 1793 5913 1807 5927
rect 2013 5913 2027 5927
rect 2053 5913 2067 5927
rect 2193 5913 2207 5927
rect 2273 5913 2287 5927
rect 2313 5913 2327 5927
rect 2573 5913 2587 5927
rect 3273 5913 3287 5927
rect 3313 5913 3327 5927
rect 3333 5913 3347 5927
rect 3373 5913 3387 5927
rect 3453 5913 3467 5927
rect 3573 5913 3587 5927
rect 3613 5913 3627 5927
rect 3793 5913 3807 5927
rect 3953 5913 3967 5927
rect 4153 5913 4167 5927
rect 4453 5913 4467 5927
rect 4493 5913 4507 5927
rect 4533 5913 4547 5927
rect 4573 5913 4587 5927
rect 4593 5913 4607 5927
rect 4653 5913 4667 5927
rect 4713 5913 4727 5927
rect 5093 5913 5107 5927
rect 5133 5913 5147 5927
rect 5173 5913 5187 5927
rect 5233 5913 5247 5927
rect 5273 5913 5287 5927
rect 5333 5913 5347 5927
rect 5373 5913 5387 5927
rect 5413 5913 5427 5927
rect 5753 5913 5767 5927
rect 5833 5913 5847 5927
rect 5873 5913 5887 5927
rect 5893 5913 5907 5927
rect 5933 5913 5947 5927
rect 6033 5913 6047 5927
rect 6073 5913 6087 5927
rect 6093 5913 6107 5927
rect 6133 5913 6147 5927
rect 6173 5913 6187 5927
rect 6293 5913 6307 5927
rect 6353 5913 6367 5927
rect 6393 5913 6407 5927
rect 6433 5913 6447 5927
rect 113 5893 127 5907
rect 193 5893 207 5907
rect 293 5893 307 5907
rect 333 5893 347 5907
rect 393 5893 407 5907
rect 453 5893 467 5907
rect 673 5893 687 5907
rect 713 5893 727 5907
rect 773 5893 787 5907
rect 933 5893 947 5907
rect 993 5893 1007 5907
rect 1033 5893 1047 5907
rect 1173 5893 1187 5907
rect 1473 5893 1487 5907
rect 1573 5893 1587 5907
rect 1613 5893 1627 5907
rect 1653 5893 1667 5907
rect 1693 5893 1707 5907
rect 1853 5893 1867 5907
rect 1893 5893 1907 5907
rect 1933 5893 1947 5907
rect 1993 5893 2007 5907
rect 2033 5893 2047 5907
rect 2073 5893 2087 5907
rect 2113 5893 2127 5907
rect 2213 5893 2227 5907
rect 2253 5893 2267 5907
rect 2293 5893 2307 5907
rect 2333 5893 2347 5907
rect 2413 5893 2427 5907
rect 2493 5893 2507 5907
rect 2533 5893 2547 5907
rect 2593 5893 2607 5907
rect 2633 5893 2647 5907
rect 2673 5893 2687 5907
rect 2773 5893 2787 5907
rect 2813 5893 2827 5907
rect 2873 5893 2887 5907
rect 2913 5893 2927 5907
rect 2973 5893 2987 5907
rect 3013 5893 3027 5907
rect 3073 5893 3087 5907
rect 3113 5893 3127 5907
rect 3133 5893 3147 5907
rect 3173 5893 3187 5907
rect 3253 5893 3267 5907
rect 3293 5893 3307 5907
rect 3353 5893 3367 5907
rect 3393 5893 3407 5907
rect 3473 5893 3487 5907
rect 3513 5893 3527 5907
rect 3553 5893 3567 5907
rect 3593 5893 3607 5907
rect 3673 5893 3687 5907
rect 3713 5893 3727 5907
rect 3733 5893 3747 5907
rect 3773 5893 3787 5907
rect 3873 5893 3887 5907
rect 3913 5893 3927 5907
rect 3973 5893 3987 5907
rect 4013 5893 4027 5907
rect 4073 5893 4087 5907
rect 4113 5893 4127 5907
rect 4173 5893 4187 5907
rect 4213 5893 4227 5907
rect 4233 5893 4247 5907
rect 4273 5893 4287 5907
rect 4353 5893 4367 5907
rect 4433 5893 4447 5907
rect 4473 5893 4487 5907
rect 4733 5893 4747 5907
rect 4773 5893 4787 5907
rect 4813 5893 4827 5907
rect 4893 5893 4907 5907
rect 4973 5893 4987 5907
rect 5013 5893 5027 5907
rect 5033 5893 5047 5907
rect 5073 5893 5087 5907
rect 5153 5893 5167 5907
rect 5193 5893 5207 5907
rect 5253 5893 5267 5907
rect 5293 5893 5307 5907
rect 5353 5893 5367 5907
rect 5393 5893 5407 5907
rect 5493 5893 5507 5907
rect 5553 5893 5567 5907
rect 5633 5893 5647 5907
rect 5673 5893 5687 5907
rect 5693 5893 5707 5907
rect 5733 5893 5747 5907
rect 5813 5893 5827 5907
rect 5853 5893 5867 5907
rect 5913 5893 5927 5907
rect 5953 5893 5967 5907
rect 6013 5893 6027 5907
rect 6053 5893 6067 5907
rect 6113 5893 6127 5907
rect 6153 5893 6167 5907
rect 6253 5893 6267 5907
rect 6413 5893 6427 5907
rect 6453 5893 6467 5907
rect 6493 5893 6507 5907
rect 6533 5893 6547 5907
rect 6613 5893 6627 5907
rect 93 5873 107 5887
rect 133 5873 147 5887
rect 173 5873 187 5887
rect 213 5873 227 5887
rect 373 5873 387 5887
rect 413 5873 427 5887
rect 913 5873 927 5887
rect 953 5873 967 5887
rect 1453 5873 1467 5887
rect 1493 5873 1507 5887
rect 1553 5873 1567 5887
rect 1593 5873 1607 5887
rect 1833 5873 1847 5887
rect 1873 5873 1887 5887
rect 2093 5873 2107 5887
rect 2133 5873 2147 5887
rect 2393 5873 2407 5887
rect 2433 5873 2447 5887
rect 2473 5873 2487 5887
rect 2513 5873 2527 5887
rect 2653 5873 2667 5887
rect 2693 5873 2707 5887
rect 2753 5873 2767 5887
rect 2793 5873 2807 5887
rect 2853 5873 2867 5887
rect 2893 5873 2907 5887
rect 2953 5873 2967 5887
rect 2993 5873 3007 5887
rect 3053 5873 3067 5887
rect 3093 5873 3107 5887
rect 3153 5873 3167 5887
rect 3193 5873 3207 5887
rect 3653 5873 3667 5887
rect 3693 5873 3707 5887
rect 3853 5873 3867 5887
rect 3893 5873 3907 5887
rect 4053 5873 4067 5887
rect 4093 5873 4107 5887
rect 4253 5873 4267 5887
rect 4293 5873 4307 5887
rect 4333 5873 4347 5887
rect 4373 5873 4387 5887
rect 4633 5873 4647 5887
rect 4793 5873 4807 5887
rect 4833 5873 4847 5887
rect 4953 5873 4967 5887
rect 4993 5873 5007 5887
rect 5473 5873 5487 5887
rect 5513 5873 5527 5887
rect 5613 5873 5627 5887
rect 5653 5873 5667 5887
rect 6233 5873 6247 5887
rect 6273 5873 6287 5887
rect 6333 5873 6347 5887
rect 6513 5873 6527 5887
rect 6553 5873 6567 5887
rect 6593 5873 6607 5887
rect 6633 5873 6647 5887
rect 593 5653 607 5667
rect 633 5653 647 5667
rect 713 5653 727 5667
rect 773 5653 787 5667
rect 813 5653 827 5667
rect 853 5653 867 5667
rect 893 5653 907 5667
rect 1933 5653 1947 5667
rect 1973 5653 1987 5667
rect 2233 5653 2247 5667
rect 2273 5653 2287 5667
rect 2513 5653 2527 5667
rect 2553 5653 2567 5667
rect 2593 5653 2607 5667
rect 2633 5653 2647 5667
rect 2693 5653 2707 5667
rect 2733 5653 2747 5667
rect 2773 5653 2787 5667
rect 2813 5653 2827 5667
rect 2973 5653 2987 5667
rect 3013 5653 3027 5667
rect 3333 5653 3347 5667
rect 3373 5653 3387 5667
rect 3433 5653 3447 5667
rect 3473 5653 3487 5667
rect 3533 5653 3547 5667
rect 3573 5653 3587 5667
rect 4253 5653 4267 5667
rect 4293 5653 4307 5667
rect 4533 5653 4547 5667
rect 4593 5653 4607 5667
rect 4633 5653 4647 5667
rect 4893 5653 4907 5667
rect 4933 5653 4947 5667
rect 5193 5653 5207 5667
rect 5233 5653 5247 5667
rect 5273 5653 5287 5667
rect 5313 5653 5327 5667
rect 5373 5653 5387 5667
rect 5413 5653 5427 5667
rect 5553 5653 5567 5667
rect 5593 5653 5607 5667
rect 5653 5653 5667 5667
rect 5693 5653 5707 5667
rect 6133 5653 6147 5667
rect 6173 5653 6187 5667
rect 6393 5653 6407 5667
rect 6433 5653 6447 5667
rect 6493 5653 6507 5667
rect 6533 5653 6547 5667
rect 6593 5653 6607 5667
rect 6633 5653 6647 5667
rect 493 5633 507 5647
rect 533 5633 547 5647
rect 613 5633 627 5647
rect 793 5633 807 5647
rect 873 5633 887 5647
rect 1033 5633 1047 5647
rect 1133 5633 1147 5647
rect 1273 5633 1287 5647
rect 1413 5633 1427 5647
rect 1713 5633 1727 5647
rect 1753 5633 1767 5647
rect 1833 5633 1847 5647
rect 1873 5633 1887 5647
rect 1953 5633 1967 5647
rect 2013 5633 2027 5647
rect 2093 5633 2107 5647
rect 2133 5633 2147 5647
rect 2253 5633 2267 5647
rect 2353 5633 2367 5647
rect 2413 5633 2427 5647
rect 2533 5633 2547 5647
rect 2613 5633 2627 5647
rect 2653 5633 2667 5647
rect 2713 5633 2727 5647
rect 2753 5633 2767 5647
rect 2793 5633 2807 5647
rect 2873 5633 2887 5647
rect 2913 5633 2927 5647
rect 2993 5633 3007 5647
rect 3033 5633 3047 5647
rect 3053 5633 3067 5647
rect 3093 5633 3107 5647
rect 3173 5633 3187 5647
rect 3213 5633 3227 5647
rect 3273 5633 3287 5647
rect 3313 5633 3327 5647
rect 3353 5633 3367 5647
rect 3453 5633 3467 5647
rect 3493 5633 3507 5647
rect 3553 5633 3567 5647
rect 3593 5633 3607 5647
rect 3633 5633 3647 5647
rect 3693 5633 3707 5647
rect 3733 5633 3747 5647
rect 3873 5633 3887 5647
rect 3913 5633 3927 5647
rect 3973 5633 3987 5647
rect 4053 5633 4067 5647
rect 4093 5633 4107 5647
rect 4153 5633 4167 5647
rect 4193 5633 4207 5647
rect 4273 5633 4287 5647
rect 4313 5633 4327 5647
rect 4353 5633 4367 5647
rect 4413 5633 4427 5647
rect 4453 5633 4467 5647
rect 4613 5633 4627 5647
rect 4693 5633 4707 5647
rect 4733 5633 4747 5647
rect 4793 5633 4807 5647
rect 4833 5633 4847 5647
rect 4913 5633 4927 5647
rect 4953 5633 4967 5647
rect 4973 5633 4987 5647
rect 5013 5633 5027 5647
rect 5093 5633 5107 5647
rect 5133 5633 5147 5647
rect 5173 5633 5187 5647
rect 5213 5633 5227 5647
rect 5293 5633 5307 5647
rect 5353 5633 5367 5647
rect 5393 5633 5407 5647
rect 5453 5633 5467 5647
rect 5493 5633 5507 5647
rect 5573 5633 5587 5647
rect 5673 5633 5687 5647
rect 5733 5633 5747 5647
rect 5773 5633 5787 5647
rect 5853 5633 5867 5647
rect 5893 5633 5907 5647
rect 5953 5633 5967 5647
rect 6013 5633 6027 5647
rect 6053 5633 6067 5647
rect 6113 5633 6127 5647
rect 6153 5633 6167 5647
rect 6233 5633 6247 5647
rect 6273 5633 6287 5647
rect 6313 5633 6327 5647
rect 6373 5633 6387 5647
rect 6413 5633 6427 5647
rect 6473 5633 6487 5647
rect 6513 5633 6527 5647
rect 6573 5633 6587 5647
rect 6613 5633 6627 5647
rect 33 5613 47 5627
rect 73 5613 87 5627
rect 113 5613 127 5627
rect 153 5613 167 5627
rect 193 5613 207 5627
rect 273 5613 287 5627
rect 313 5613 327 5627
rect 433 5613 447 5627
rect 473 5613 487 5627
rect 553 5613 567 5627
rect 673 5613 687 5627
rect 733 5613 747 5627
rect 933 5613 947 5627
rect 973 5613 987 5627
rect 1093 5613 1107 5627
rect 1173 5613 1187 5627
rect 1213 5613 1227 5627
rect 1313 5613 1327 5627
rect 1353 5613 1367 5627
rect 1473 5613 1487 5627
rect 1553 5613 1567 5627
rect 1593 5613 1607 5627
rect 1693 5613 1707 5627
rect 1733 5613 1747 5627
rect 1773 5613 1787 5627
rect 1853 5613 1867 5627
rect 1893 5613 1907 5627
rect 2073 5613 2087 5627
rect 2153 5613 2167 5627
rect 2193 5613 2207 5627
rect 2393 5613 2407 5627
rect 2453 5613 2467 5627
rect 2853 5613 2867 5627
rect 2893 5613 2907 5627
rect 3113 5613 3127 5627
rect 3193 5613 3207 5627
rect 3233 5613 3247 5627
rect 3713 5613 3727 5627
rect 3753 5613 3767 5627
rect 3793 5613 3807 5627
rect 3833 5613 3847 5627
rect 3853 5613 3867 5627
rect 3893 5613 3907 5627
rect 4033 5613 4047 5627
rect 4073 5613 4087 5627
rect 4113 5613 4127 5627
rect 4173 5613 4187 5627
rect 4213 5613 4227 5627
rect 4433 5613 4447 5627
rect 4473 5613 4487 5627
rect 4513 5613 4527 5627
rect 4573 5613 4587 5627
rect 4713 5613 4727 5627
rect 4753 5613 4767 5627
rect 4773 5613 4787 5627
rect 4813 5613 4827 5627
rect 5033 5613 5047 5627
rect 5073 5613 5087 5627
rect 5113 5613 5127 5627
rect 5513 5613 5527 5627
rect 5713 5613 5727 5627
rect 5753 5613 5767 5627
rect 5793 5613 5807 5627
rect 5873 5613 5887 5627
rect 5913 5613 5927 5627
rect 5993 5613 6007 5627
rect 6033 5613 6047 5627
rect 6073 5613 6087 5627
rect 6333 5613 6347 5627
rect 453 5593 467 5607
rect 513 5593 527 5607
rect 953 5593 967 5607
rect 1013 5593 1027 5607
rect 1073 5593 1087 5607
rect 1193 5593 1207 5607
rect 1253 5593 1267 5607
rect 1333 5593 1347 5607
rect 1393 5593 1407 5607
rect 1993 5593 2007 5607
rect 2113 5593 2127 5607
rect 2173 5593 2187 5607
rect 3073 5593 3087 5607
rect 3293 5593 3307 5607
rect 3653 5593 3667 5607
rect 3813 5593 3827 5607
rect 3993 5593 4007 5607
rect 4333 5593 4347 5607
rect 4993 5593 5007 5607
rect 5473 5593 5487 5607
rect 5933 5593 5947 5607
rect 6253 5593 6267 5607
rect 6293 5593 6307 5607
rect 393 5453 407 5467
rect 633 5453 647 5467
rect 713 5453 727 5467
rect 933 5453 947 5467
rect 1013 5453 1027 5467
rect 1693 5453 1707 5467
rect 2213 5453 2227 5467
rect 2353 5453 2367 5467
rect 2453 5453 2467 5467
rect 2533 5453 2547 5467
rect 2973 5453 2987 5467
rect 3413 5453 3427 5467
rect 3473 5453 3487 5467
rect 3713 5453 3727 5467
rect 3913 5453 3927 5467
rect 4233 5453 4247 5467
rect 6113 5453 6127 5467
rect 6653 5453 6667 5467
rect 33 5433 47 5447
rect 113 5433 127 5447
rect 153 5433 167 5447
rect 353 5433 367 5447
rect 533 5433 547 5447
rect 593 5433 607 5447
rect 613 5433 627 5447
rect 653 5433 667 5447
rect 693 5433 707 5447
rect 733 5433 747 5447
rect 1053 5433 1067 5447
rect 1113 5433 1127 5447
rect 1153 5433 1167 5447
rect 1193 5433 1207 5447
rect 1233 5433 1247 5447
rect 1313 5433 1327 5447
rect 1353 5433 1367 5447
rect 1753 5433 1767 5447
rect 1793 5433 1807 5447
rect 1833 5433 1847 5447
rect 1893 5433 1907 5447
rect 2033 5433 2047 5447
rect 2073 5433 2087 5447
rect 2273 5433 2287 5447
rect 2313 5433 2327 5447
rect 2333 5433 2347 5447
rect 2373 5433 2387 5447
rect 2493 5433 2507 5447
rect 2573 5433 2587 5447
rect 2613 5433 2627 5447
rect 2953 5433 2967 5447
rect 2993 5433 3007 5447
rect 3013 5433 3027 5447
rect 3053 5433 3067 5447
rect 3193 5433 3207 5447
rect 3233 5433 3247 5447
rect 3313 5433 3327 5447
rect 3373 5433 3387 5447
rect 3393 5433 3407 5447
rect 3433 5433 3447 5447
rect 3493 5433 3507 5447
rect 3573 5433 3587 5447
rect 3613 5433 3627 5447
rect 3693 5433 3707 5447
rect 3733 5433 3747 5447
rect 3753 5433 3767 5447
rect 3793 5433 3807 5447
rect 3833 5433 3847 5447
rect 3893 5433 3907 5447
rect 3933 5433 3947 5447
rect 3953 5433 3967 5447
rect 3993 5433 4007 5447
rect 4333 5433 4347 5447
rect 4373 5433 4387 5447
rect 4593 5433 4607 5447
rect 4633 5433 4647 5447
rect 4693 5433 4707 5447
rect 4733 5433 4747 5447
rect 4773 5433 4787 5447
rect 4833 5433 4847 5447
rect 4893 5433 4907 5447
rect 4933 5433 4947 5447
rect 5053 5433 5067 5447
rect 5113 5433 5127 5447
rect 5213 5433 5227 5447
rect 5253 5433 5267 5447
rect 5333 5433 5347 5447
rect 5393 5433 5407 5447
rect 5413 5433 5427 5447
rect 5453 5433 5467 5447
rect 5713 5433 5727 5447
rect 5773 5433 5787 5447
rect 5813 5433 5827 5447
rect 5853 5433 5867 5447
rect 5893 5433 5907 5447
rect 6153 5433 6167 5447
rect 6233 5433 6247 5447
rect 6273 5433 6287 5447
rect 6293 5433 6307 5447
rect 6333 5433 6347 5447
rect 6433 5433 6447 5447
rect 6473 5433 6487 5447
rect 6613 5433 6627 5447
rect 273 5413 287 5427
rect 373 5413 387 5427
rect 413 5413 427 5427
rect 473 5413 487 5427
rect 793 5413 807 5427
rect 873 5413 887 5427
rect 953 5413 967 5427
rect 993 5413 1007 5427
rect 1033 5413 1047 5427
rect 1133 5413 1147 5427
rect 1173 5413 1187 5427
rect 1493 5413 1507 5427
rect 1533 5413 1547 5427
rect 1593 5413 1607 5427
rect 1633 5413 1647 5427
rect 1673 5413 1687 5427
rect 1733 5413 1747 5427
rect 1773 5413 1787 5427
rect 1953 5413 1967 5427
rect 2013 5413 2027 5427
rect 2053 5413 2067 5427
rect 2113 5413 2127 5427
rect 2193 5413 2207 5427
rect 2253 5413 2267 5427
rect 2293 5413 2307 5427
rect 2433 5413 2447 5427
rect 2513 5413 2527 5427
rect 2553 5413 2567 5427
rect 2593 5413 2607 5427
rect 2633 5413 2647 5427
rect 2693 5413 2707 5427
rect 2793 5413 2807 5427
rect 2833 5413 2847 5427
rect 2893 5413 2907 5427
rect 3033 5413 3047 5427
rect 3073 5413 3087 5427
rect 3153 5413 3167 5427
rect 3213 5413 3227 5427
rect 3253 5413 3267 5427
rect 3533 5413 3547 5427
rect 3593 5413 3607 5427
rect 3633 5413 3647 5427
rect 3773 5413 3787 5427
rect 3813 5413 3827 5427
rect 3973 5413 3987 5427
rect 4013 5413 4027 5427
rect 4093 5413 4107 5427
rect 4133 5413 4147 5427
rect 4193 5413 4207 5427
rect 4253 5413 4267 5427
rect 4313 5413 4327 5427
rect 4353 5413 4367 5427
rect 4433 5413 4447 5427
rect 4493 5413 4507 5427
rect 4573 5413 4587 5427
rect 4613 5413 4627 5427
rect 4673 5413 4687 5427
rect 4713 5413 4727 5427
rect 4873 5413 4887 5427
rect 4913 5413 4927 5427
rect 4993 5413 5007 5427
rect 5153 5413 5167 5427
rect 5233 5413 5247 5427
rect 5273 5413 5287 5427
rect 5433 5413 5447 5427
rect 5473 5413 5487 5427
rect 5533 5413 5547 5427
rect 5593 5413 5607 5427
rect 5633 5413 5647 5427
rect 5833 5413 5847 5427
rect 5873 5413 5887 5427
rect 5933 5413 5947 5427
rect 5993 5413 6007 5427
rect 6033 5413 6047 5427
rect 6093 5413 6107 5427
rect 6133 5413 6147 5427
rect 6213 5413 6227 5427
rect 6253 5413 6267 5427
rect 6313 5413 6327 5427
rect 6353 5413 6367 5427
rect 6413 5413 6427 5427
rect 6453 5413 6467 5427
rect 6533 5413 6547 5427
rect 6573 5413 6587 5427
rect 6633 5413 6647 5427
rect 6673 5413 6687 5427
rect 253 5393 267 5407
rect 293 5393 307 5407
rect 453 5393 467 5407
rect 493 5393 507 5407
rect 553 5393 567 5407
rect 773 5393 787 5407
rect 813 5393 827 5407
rect 853 5393 867 5407
rect 893 5393 907 5407
rect 1473 5393 1487 5407
rect 1513 5393 1527 5407
rect 1573 5393 1587 5407
rect 1613 5393 1627 5407
rect 1853 5393 1867 5407
rect 1933 5393 1947 5407
rect 1973 5393 1987 5407
rect 2093 5393 2107 5407
rect 2133 5393 2147 5407
rect 2673 5393 2687 5407
rect 2713 5393 2727 5407
rect 2773 5393 2787 5407
rect 2813 5393 2827 5407
rect 2873 5393 2887 5407
rect 2913 5393 2927 5407
rect 3133 5393 3147 5407
rect 3173 5393 3187 5407
rect 3333 5393 3347 5407
rect 4073 5393 4087 5407
rect 4113 5393 4127 5407
rect 4173 5393 4187 5407
rect 4213 5393 4227 5407
rect 4413 5393 4427 5407
rect 4453 5393 4467 5407
rect 4473 5393 4487 5407
rect 4513 5393 4527 5407
rect 4793 5393 4807 5407
rect 4973 5393 4987 5407
rect 5013 5393 5027 5407
rect 5073 5393 5087 5407
rect 5133 5393 5147 5407
rect 5173 5393 5187 5407
rect 5353 5393 5367 5407
rect 5513 5393 5527 5407
rect 5553 5393 5567 5407
rect 5613 5393 5627 5407
rect 5653 5393 5667 5407
rect 5733 5393 5747 5407
rect 5913 5393 5927 5407
rect 5953 5393 5967 5407
rect 6013 5393 6027 5407
rect 6053 5393 6067 5407
rect 6513 5393 6527 5407
rect 6553 5393 6567 5407
rect 333 5173 347 5187
rect 373 5173 387 5187
rect 533 5173 547 5187
rect 573 5173 587 5187
rect 833 5173 847 5187
rect 873 5173 887 5187
rect 1153 5173 1167 5187
rect 1473 5173 1487 5187
rect 1513 5173 1527 5187
rect 1533 5173 1547 5187
rect 1573 5173 1587 5187
rect 2073 5173 2087 5187
rect 2133 5173 2147 5187
rect 2173 5173 2187 5187
rect 2333 5173 2347 5187
rect 2373 5173 2387 5187
rect 2413 5173 2427 5187
rect 2453 5173 2467 5187
rect 2673 5173 2687 5187
rect 2833 5173 2847 5187
rect 2873 5173 2887 5187
rect 2913 5173 2927 5187
rect 2953 5173 2967 5187
rect 3113 5173 3127 5187
rect 3173 5173 3187 5187
rect 3213 5173 3227 5187
rect 3273 5173 3287 5187
rect 3313 5173 3327 5187
rect 3873 5173 3887 5187
rect 3913 5173 3927 5187
rect 3973 5173 3987 5187
rect 4013 5173 4027 5187
rect 4153 5173 4167 5187
rect 4193 5173 4207 5187
rect 4253 5173 4267 5187
rect 4333 5173 4347 5187
rect 4373 5173 4387 5187
rect 4593 5173 4607 5187
rect 4633 5173 4647 5187
rect 4673 5173 4687 5187
rect 4713 5173 4727 5187
rect 4833 5173 4847 5187
rect 4873 5173 4887 5187
rect 5073 5173 5087 5187
rect 5113 5173 5127 5187
rect 5233 5173 5247 5187
rect 5273 5173 5287 5187
rect 5433 5173 5447 5187
rect 5473 5173 5487 5187
rect 5533 5173 5547 5187
rect 5573 5173 5587 5187
rect 5693 5173 5707 5187
rect 5733 5173 5747 5187
rect 5893 5173 5907 5187
rect 5933 5173 5947 5187
rect 5973 5173 5987 5187
rect 6013 5173 6027 5187
rect 6053 5173 6067 5187
rect 6093 5173 6107 5187
rect 6313 5173 6327 5187
rect 6353 5173 6367 5187
rect 6413 5173 6427 5187
rect 6453 5173 6467 5187
rect 6573 5173 6587 5187
rect 6613 5173 6627 5187
rect 6653 5173 6667 5187
rect 6693 5173 6707 5187
rect 353 5153 367 5167
rect 453 5153 467 5167
rect 493 5153 507 5167
rect 553 5153 567 5167
rect 853 5153 867 5167
rect 933 5153 947 5167
rect 973 5153 987 5167
rect 1033 5153 1047 5167
rect 1073 5153 1087 5167
rect 1493 5153 1507 5167
rect 1553 5153 1567 5167
rect 1893 5153 1907 5167
rect 1933 5153 1947 5167
rect 1993 5153 2007 5167
rect 2153 5153 2167 5167
rect 2233 5153 2247 5167
rect 2353 5153 2367 5167
rect 2433 5153 2447 5167
rect 2473 5153 2487 5167
rect 2593 5153 2607 5167
rect 2853 5153 2867 5167
rect 2933 5153 2947 5167
rect 3033 5153 3047 5167
rect 3193 5153 3207 5167
rect 3293 5153 3307 5167
rect 3333 5153 3347 5167
rect 3373 5153 3387 5167
rect 3453 5153 3467 5167
rect 3493 5153 3507 5167
rect 3613 5153 3627 5167
rect 3653 5153 3667 5167
rect 3713 5153 3727 5167
rect 3753 5153 3767 5167
rect 3893 5153 3907 5167
rect 3993 5153 4007 5167
rect 4053 5153 4067 5167
rect 4093 5153 4107 5167
rect 4173 5153 4187 5167
rect 4353 5153 4367 5167
rect 4413 5153 4427 5167
rect 4453 5153 4467 5167
rect 4513 5153 4527 5167
rect 4553 5153 4567 5167
rect 4613 5153 4627 5167
rect 4693 5153 4707 5167
rect 4773 5153 4787 5167
rect 4853 5153 4867 5167
rect 4893 5153 4907 5167
rect 4933 5153 4947 5167
rect 4973 5153 4987 5167
rect 5013 5153 5027 5167
rect 5093 5153 5107 5167
rect 5153 5153 5167 5167
rect 5193 5153 5207 5167
rect 5253 5153 5267 5167
rect 5333 5153 5347 5167
rect 5373 5153 5387 5167
rect 5413 5153 5427 5167
rect 5453 5153 5467 5167
rect 5513 5153 5527 5167
rect 5553 5153 5567 5167
rect 5633 5153 5647 5167
rect 5673 5153 5687 5167
rect 5713 5153 5727 5167
rect 5793 5153 5807 5167
rect 5833 5153 5847 5167
rect 5913 5153 5927 5167
rect 5953 5153 5967 5167
rect 5993 5153 6007 5167
rect 6073 5153 6087 5167
rect 6173 5153 6187 5167
rect 6213 5153 6227 5167
rect 6253 5153 6267 5167
rect 6333 5153 6347 5167
rect 6373 5153 6387 5167
rect 6433 5153 6447 5167
rect 6473 5153 6487 5167
rect 6513 5153 6527 5167
rect 6593 5153 6607 5167
rect 6633 5153 6647 5167
rect 6673 5153 6687 5167
rect 33 5133 47 5147
rect 73 5133 87 5147
rect 113 5133 127 5147
rect 193 5133 207 5147
rect 233 5133 247 5147
rect 433 5133 447 5147
rect 673 5133 687 5147
rect 713 5133 727 5147
rect 793 5133 807 5147
rect 953 5133 967 5147
rect 993 5133 1007 5147
rect 1053 5133 1067 5147
rect 1093 5133 1107 5147
rect 1133 5133 1147 5147
rect 1193 5133 1207 5147
rect 1233 5133 1247 5147
rect 1313 5133 1327 5147
rect 1353 5133 1367 5147
rect 1633 5133 1647 5147
rect 1713 5133 1727 5147
rect 1753 5133 1767 5147
rect 1873 5133 1887 5147
rect 1913 5133 1927 5147
rect 1953 5133 1967 5147
rect 2053 5133 2067 5147
rect 2113 5133 2127 5147
rect 2273 5133 2287 5147
rect 2513 5133 2527 5147
rect 2553 5133 2567 5147
rect 2653 5133 2667 5147
rect 2713 5133 2727 5147
rect 2733 5133 2747 5147
rect 2773 5133 2787 5147
rect 2993 5133 3007 5147
rect 3093 5133 3107 5147
rect 3153 5133 3167 5147
rect 3433 5133 3447 5147
rect 3533 5133 3547 5147
rect 3573 5133 3587 5147
rect 3593 5133 3607 5147
rect 3633 5133 3647 5147
rect 3733 5133 3747 5147
rect 3773 5133 3787 5147
rect 3793 5133 3807 5147
rect 3833 5133 3847 5147
rect 4033 5133 4047 5147
rect 4073 5133 4087 5147
rect 4233 5133 4247 5147
rect 4293 5133 4307 5147
rect 4433 5133 4447 5147
rect 4473 5133 4487 5147
rect 4533 5133 4547 5147
rect 4573 5133 4587 5147
rect 4913 5133 4927 5147
rect 4953 5133 4967 5147
rect 5033 5133 5047 5147
rect 5313 5133 5327 5147
rect 5353 5133 5367 5147
rect 5773 5133 5787 5147
rect 5813 5133 5827 5147
rect 6153 5133 6167 5147
rect 473 5113 487 5127
rect 1973 5113 1987 5127
rect 2293 5113 2307 5127
rect 2533 5113 2547 5127
rect 2573 5113 2587 5127
rect 2753 5113 2767 5127
rect 2973 5113 2987 5127
rect 3393 5113 3407 5127
rect 3473 5113 3487 5127
rect 3553 5113 3567 5127
rect 3813 5113 3827 5127
rect 4753 5113 4767 5127
rect 5613 5113 5627 5127
rect 6193 5113 6207 5127
rect 6273 5113 6287 5127
rect 6493 5113 6507 5127
rect 553 4973 567 4987
rect 1213 4973 1227 4987
rect 2233 4973 2247 4987
rect 2333 4973 2347 4987
rect 2453 4973 2467 4987
rect 2793 4973 2807 4987
rect 3153 4973 3167 4987
rect 3833 4973 3847 4987
rect 4033 4973 4047 4987
rect 5793 4973 5807 4987
rect 6653 4973 6667 4987
rect 33 4953 47 4967
rect 73 4953 87 4967
rect 113 4953 127 4967
rect 153 4953 167 4967
rect 273 4953 287 4967
rect 353 4953 367 4967
rect 393 4953 407 4967
rect 513 4953 527 4967
rect 853 4953 867 4967
rect 933 4953 947 4967
rect 973 4953 987 4967
rect 1093 4953 1107 4967
rect 1133 4953 1147 4967
rect 1173 4953 1187 4967
rect 1353 4953 1367 4967
rect 1393 4953 1407 4967
rect 1613 4953 1627 4967
rect 1653 4953 1667 4967
rect 1793 4953 1807 4967
rect 1833 4953 1847 4967
rect 1973 4953 1987 4967
rect 2013 4953 2027 4967
rect 2073 4953 2087 4967
rect 2113 4953 2127 4967
rect 2153 4953 2167 4967
rect 2213 4953 2227 4967
rect 2313 4953 2327 4967
rect 2353 4953 2367 4967
rect 2433 4953 2447 4967
rect 2593 4953 2607 4967
rect 2633 4953 2647 4967
rect 2693 4953 2707 4967
rect 2733 4953 2747 4967
rect 2813 4953 2827 4967
rect 2853 4953 2867 4967
rect 2953 4953 2967 4967
rect 2993 4953 3007 4967
rect 3053 4953 3067 4967
rect 3093 4953 3107 4967
rect 3133 4953 3147 4967
rect 3173 4953 3187 4967
rect 3213 4953 3227 4967
rect 3373 4953 3387 4967
rect 3413 4953 3427 4967
rect 3513 4953 3527 4967
rect 3553 4953 3567 4967
rect 3633 4953 3647 4967
rect 3673 4953 3687 4967
rect 3713 4953 3727 4967
rect 3793 4953 3807 4967
rect 3993 4953 4007 4967
rect 4093 4953 4107 4967
rect 4153 4953 4167 4967
rect 4213 4953 4227 4967
rect 4313 4953 4327 4967
rect 4373 4953 4387 4967
rect 4453 4953 4467 4967
rect 4493 4953 4507 4967
rect 4613 4953 4627 4967
rect 4653 4953 4667 4967
rect 4813 4953 4827 4967
rect 4873 4953 4887 4967
rect 5053 4953 5067 4967
rect 5113 4953 5127 4967
rect 5253 4953 5267 4967
rect 5313 4953 5327 4967
rect 5333 4953 5347 4967
rect 5393 4953 5407 4967
rect 5453 4953 5467 4967
rect 5493 4953 5507 4967
rect 5533 4953 5547 4967
rect 5753 4953 5767 4967
rect 6013 4953 6027 4967
rect 6053 4953 6067 4967
rect 6093 4953 6107 4967
rect 6233 4953 6247 4967
rect 6273 4953 6287 4967
rect 213 4933 227 4947
rect 533 4933 547 4947
rect 573 4933 587 4947
rect 633 4933 647 4947
rect 693 4933 707 4947
rect 793 4933 807 4947
rect 1193 4933 1207 4947
rect 1233 4933 1247 4947
rect 1293 4933 1307 4947
rect 1433 4933 1447 4947
rect 1533 4933 1547 4947
rect 1593 4933 1607 4947
rect 1633 4933 1647 4947
rect 1713 4933 1727 4947
rect 1773 4933 1787 4947
rect 1813 4933 1827 4947
rect 1873 4933 1887 4947
rect 1953 4933 1967 4947
rect 1993 4933 2007 4947
rect 2053 4933 2067 4947
rect 2093 4933 2107 4947
rect 2253 4933 2267 4947
rect 2393 4933 2407 4947
rect 2513 4933 2527 4947
rect 2573 4933 2587 4947
rect 2613 4933 2627 4947
rect 2673 4933 2687 4947
rect 2713 4933 2727 4947
rect 2773 4933 2787 4947
rect 2833 4933 2847 4947
rect 2873 4933 2887 4947
rect 2933 4933 2947 4947
rect 2973 4933 2987 4947
rect 3033 4933 3047 4947
rect 3073 4933 3087 4947
rect 3233 4933 3247 4947
rect 3293 4933 3307 4947
rect 3353 4933 3367 4947
rect 3393 4933 3407 4947
rect 3693 4933 3707 4947
rect 3733 4933 3747 4947
rect 3813 4933 3827 4947
rect 3853 4933 3867 4947
rect 3913 4933 3927 4947
rect 3953 4933 3967 4947
rect 4013 4933 4027 4947
rect 4053 4933 4067 4947
rect 4113 4933 4127 4947
rect 4273 4933 4287 4947
rect 4433 4933 4447 4947
rect 4473 4933 4487 4947
rect 4513 4933 4527 4947
rect 4553 4933 4567 4947
rect 4633 4933 4647 4947
rect 4673 4933 4687 4947
rect 4753 4933 4767 4947
rect 4933 4933 4947 4947
rect 4993 4933 5007 4947
rect 5193 4933 5207 4947
rect 5473 4933 5487 4947
rect 5513 4933 5527 4947
rect 5593 4933 5607 4947
rect 5633 4933 5647 4947
rect 5673 4933 5687 4947
rect 5773 4933 5787 4947
rect 5813 4933 5827 4947
rect 5873 4933 5887 4947
rect 5913 4933 5927 4947
rect 5973 4933 5987 4947
rect 6033 4933 6047 4947
rect 6073 4933 6087 4947
rect 6173 4933 6187 4947
rect 6213 4933 6227 4947
rect 6253 4933 6267 4947
rect 6293 4933 6307 4947
rect 6373 4933 6387 4947
rect 6413 4933 6427 4947
rect 6473 4933 6487 4947
rect 6513 4933 6527 4947
rect 6553 4933 6567 4947
rect 6633 4933 6647 4947
rect 193 4913 207 4927
rect 233 4913 247 4927
rect 613 4913 627 4927
rect 653 4913 667 4927
rect 673 4913 687 4927
rect 713 4913 727 4927
rect 773 4913 787 4927
rect 813 4913 827 4927
rect 1273 4913 1287 4927
rect 1313 4913 1327 4927
rect 1413 4913 1427 4927
rect 1453 4913 1467 4927
rect 1513 4913 1527 4927
rect 1553 4913 1567 4927
rect 1693 4913 1707 4927
rect 1733 4913 1747 4927
rect 1853 4913 1867 4927
rect 1893 4913 1907 4927
rect 2173 4913 2187 4927
rect 2493 4913 2507 4927
rect 2533 4913 2547 4927
rect 3273 4913 3287 4927
rect 3313 4913 3327 4927
rect 3893 4913 3907 4927
rect 3933 4913 3947 4927
rect 4173 4913 4187 4927
rect 4253 4913 4267 4927
rect 4293 4913 4307 4927
rect 4353 4913 4367 4927
rect 4533 4913 4547 4927
rect 4573 4913 4587 4927
rect 4733 4913 4747 4927
rect 4773 4913 4787 4927
rect 4833 4913 4847 4927
rect 4913 4913 4927 4927
rect 4953 4913 4967 4927
rect 4973 4913 4987 4927
rect 5013 4913 5027 4927
rect 5093 4913 5107 4927
rect 5173 4913 5187 4927
rect 5213 4913 5227 4927
rect 5273 4913 5287 4927
rect 5373 4913 5387 4927
rect 5573 4913 5587 4927
rect 5613 4913 5627 4927
rect 5653 4913 5667 4927
rect 5693 4913 5707 4927
rect 5853 4913 5867 4927
rect 5893 4913 5907 4927
rect 5953 4913 5967 4927
rect 5993 4913 6007 4927
rect 6153 4913 6167 4927
rect 6193 4913 6207 4927
rect 6353 4913 6367 4927
rect 6393 4913 6407 4927
rect 6453 4913 6467 4927
rect 6493 4913 6507 4927
rect 6533 4913 6547 4927
rect 6573 4913 6587 4927
rect 633 4693 647 4707
rect 873 4693 887 4707
rect 913 4693 927 4707
rect 1293 4693 1307 4707
rect 1333 4693 1347 4707
rect 1353 4693 1367 4707
rect 1393 4693 1407 4707
rect 2193 4693 2207 4707
rect 2233 4693 2247 4707
rect 2353 4693 2367 4707
rect 2393 4693 2407 4707
rect 3673 4693 3687 4707
rect 3713 4693 3727 4707
rect 4153 4693 4167 4707
rect 4193 4693 4207 4707
rect 4473 4693 4487 4707
rect 4513 4693 4527 4707
rect 4913 4693 4927 4707
rect 4953 4693 4967 4707
rect 4993 4693 5007 4707
rect 5033 4693 5047 4707
rect 5093 4693 5107 4707
rect 5133 4693 5147 4707
rect 5373 4693 5387 4707
rect 5413 4693 5427 4707
rect 5473 4693 5487 4707
rect 5513 4693 5527 4707
rect 5553 4693 5567 4707
rect 5593 4693 5607 4707
rect 5653 4693 5667 4707
rect 5693 4693 5707 4707
rect 5733 4693 5747 4707
rect 5773 4693 5787 4707
rect 5893 4693 5907 4707
rect 5933 4693 5947 4707
rect 6013 4693 6027 4707
rect 6193 4693 6207 4707
rect 6233 4693 6247 4707
rect 6373 4693 6387 4707
rect 6413 4693 6427 4707
rect 6493 4693 6507 4707
rect 6573 4693 6587 4707
rect 6613 4693 6627 4707
rect 33 4673 47 4687
rect 173 4673 187 4687
rect 313 4673 327 4687
rect 393 4673 407 4687
rect 433 4673 447 4687
rect 473 4673 487 4687
rect 893 4673 907 4687
rect 1193 4673 1207 4687
rect 1233 4673 1247 4687
rect 1313 4673 1327 4687
rect 1373 4673 1387 4687
rect 1453 4673 1467 4687
rect 1493 4673 1507 4687
rect 1713 4673 1727 4687
rect 1853 4673 1867 4687
rect 1893 4673 1907 4687
rect 2213 4673 2227 4687
rect 2273 4673 2287 4687
rect 2373 4673 2387 4687
rect 2513 4673 2527 4687
rect 2553 4673 2567 4687
rect 2633 4673 2647 4687
rect 2933 4673 2947 4687
rect 2973 4673 2987 4687
rect 3513 4673 3527 4687
rect 3553 4673 3567 4687
rect 3633 4673 3647 4687
rect 3693 4673 3707 4687
rect 3753 4673 3767 4687
rect 3793 4673 3807 4687
rect 4113 4673 4127 4687
rect 4173 4673 4187 4687
rect 4493 4673 4507 4687
rect 4533 4673 4547 4687
rect 4573 4673 4587 4687
rect 4613 4673 4627 4687
rect 4693 4673 4707 4687
rect 4753 4673 4767 4687
rect 4793 4673 4807 4687
rect 4933 4673 4947 4687
rect 5013 4673 5027 4687
rect 5113 4673 5127 4687
rect 5173 4673 5187 4687
rect 5213 4673 5227 4687
rect 5293 4673 5307 4687
rect 5333 4673 5347 4687
rect 5393 4673 5407 4687
rect 5493 4673 5507 4687
rect 5533 4673 5547 4687
rect 5573 4673 5587 4687
rect 5673 4673 5687 4687
rect 5713 4673 5727 4687
rect 5753 4673 5767 4687
rect 5833 4673 5847 4687
rect 5873 4673 5887 4687
rect 5913 4673 5927 4687
rect 6093 4673 6107 4687
rect 6133 4673 6147 4687
rect 6213 4673 6227 4687
rect 6253 4673 6267 4687
rect 6293 4673 6307 4687
rect 6353 4673 6367 4687
rect 6393 4673 6407 4687
rect 6593 4673 6607 4687
rect 6633 4673 6647 4687
rect 233 4653 247 4667
rect 273 4653 287 4667
rect 373 4653 387 4667
rect 533 4653 547 4667
rect 573 4653 587 4667
rect 613 4653 627 4667
rect 673 4653 687 4667
rect 693 4653 707 4667
rect 733 4653 747 4667
rect 793 4653 807 4667
rect 833 4653 847 4667
rect 953 4653 967 4667
rect 1033 4653 1047 4667
rect 1073 4653 1087 4667
rect 1213 4653 1227 4667
rect 1253 4653 1267 4667
rect 1473 4653 1487 4667
rect 1513 4653 1527 4667
rect 1533 4653 1547 4667
rect 1573 4653 1587 4667
rect 1613 4653 1627 4667
rect 1653 4653 1667 4667
rect 1753 4653 1767 4667
rect 1793 4653 1807 4667
rect 1833 4653 1847 4667
rect 1873 4653 1887 4667
rect 1953 4653 1967 4667
rect 2033 4653 2047 4667
rect 2073 4653 2087 4667
rect 2313 4653 2327 4667
rect 2433 4653 2447 4667
rect 2473 4653 2487 4667
rect 2573 4653 2587 4667
rect 2693 4653 2707 4667
rect 2773 4653 2787 4667
rect 2813 4653 2827 4667
rect 2913 4653 2927 4667
rect 2953 4653 2967 4667
rect 3033 4653 3047 4667
rect 3113 4653 3127 4667
rect 3153 4653 3167 4667
rect 3273 4653 3287 4667
rect 3353 4653 3367 4667
rect 3393 4653 3407 4667
rect 3533 4653 3547 4667
rect 3573 4653 3587 4667
rect 3613 4653 3627 4667
rect 3773 4653 3787 4667
rect 3813 4653 3827 4667
rect 3913 4653 3927 4667
rect 3953 4653 3967 4667
rect 4033 4653 4047 4667
rect 4093 4653 4107 4667
rect 4233 4653 4247 4667
rect 4313 4653 4327 4667
rect 4353 4653 4367 4667
rect 4633 4653 4647 4667
rect 4733 4653 4747 4667
rect 4773 4653 4787 4667
rect 4833 4653 4847 4667
rect 4873 4653 4887 4667
rect 5153 4653 5167 4667
rect 5193 4653 5207 4667
rect 5273 4653 5287 4667
rect 5313 4653 5327 4667
rect 5353 4653 5367 4667
rect 5993 4653 6007 4667
rect 6053 4653 6067 4667
rect 6073 4653 6087 4667
rect 6113 4653 6127 4667
rect 6313 4653 6327 4667
rect 6473 4653 6487 4667
rect 6533 4653 6547 4667
rect 253 4633 267 4647
rect 333 4633 347 4647
rect 413 4633 427 4647
rect 493 4633 507 4647
rect 553 4633 567 4647
rect 713 4633 727 4647
rect 1553 4633 1567 4647
rect 1633 4633 1647 4647
rect 1693 4633 1707 4647
rect 1773 4633 1787 4647
rect 2333 4633 2347 4647
rect 2453 4633 2467 4647
rect 2533 4633 2547 4647
rect 2653 4633 2667 4647
rect 4553 4633 4567 4647
rect 4713 4633 4727 4647
rect 4853 4633 4867 4647
rect 5853 4633 5867 4647
rect 6273 4633 6287 4647
rect 53 4493 67 4507
rect 113 4493 127 4507
rect 193 4493 207 4507
rect 353 4493 367 4507
rect 493 4493 507 4507
rect 613 4493 627 4507
rect 733 4493 747 4507
rect 773 4493 787 4507
rect 833 4493 847 4507
rect 913 4493 927 4507
rect 973 4493 987 4507
rect 1353 4493 1367 4507
rect 1413 4493 1427 4507
rect 2293 4493 2307 4507
rect 2373 4493 2387 4507
rect 2453 4493 2467 4507
rect 2513 4493 2527 4507
rect 3033 4493 3047 4507
rect 4413 4493 4427 4507
rect 4513 4493 4527 4507
rect 4693 4493 4707 4507
rect 4893 4493 4907 4507
rect 5273 4493 5287 4507
rect 5393 4493 5407 4507
rect 6013 4493 6027 4507
rect 6113 4493 6127 4507
rect 6633 4493 6647 4507
rect 93 4473 107 4487
rect 133 4473 147 4487
rect 213 4473 227 4487
rect 253 4473 267 4487
rect 333 4473 347 4487
rect 373 4473 387 4487
rect 393 4473 407 4487
rect 433 4473 447 4487
rect 513 4473 527 4487
rect 653 4473 667 4487
rect 753 4473 767 4487
rect 793 4473 807 4487
rect 893 4473 907 4487
rect 933 4473 947 4487
rect 1233 4473 1247 4487
rect 1273 4473 1287 4487
rect 1393 4473 1407 4487
rect 1433 4473 1447 4487
rect 1653 4473 1667 4487
rect 1693 4473 1707 4487
rect 1813 4473 1827 4487
rect 1853 4473 1867 4487
rect 1933 4473 1947 4487
rect 2073 4473 2087 4487
rect 2153 4473 2167 4487
rect 2193 4473 2207 4487
rect 2353 4473 2367 4487
rect 2393 4473 2407 4487
rect 2433 4473 2447 4487
rect 2473 4473 2487 4487
rect 2593 4473 2607 4487
rect 2673 4473 2687 4487
rect 2713 4473 2727 4487
rect 2813 4473 2827 4487
rect 2853 4473 2867 4487
rect 3053 4473 3067 4487
rect 3093 4473 3107 4487
rect 3173 4473 3187 4487
rect 3253 4473 3267 4487
rect 3293 4473 3307 4487
rect 3393 4473 3407 4487
rect 3433 4473 3447 4487
rect 3533 4473 3547 4487
rect 3573 4473 3587 4487
rect 3673 4473 3687 4487
rect 3713 4473 3727 4487
rect 3793 4473 3807 4487
rect 3833 4473 3847 4487
rect 3873 4473 3887 4487
rect 4013 4473 4027 4487
rect 4053 4473 4067 4487
rect 4133 4473 4147 4487
rect 4273 4473 4287 4487
rect 4313 4473 4327 4487
rect 4393 4473 4407 4487
rect 4433 4473 4447 4487
rect 4473 4473 4487 4487
rect 4713 4473 4727 4487
rect 4753 4473 4767 4487
rect 4873 4473 4887 4487
rect 5093 4473 5107 4487
rect 5133 4473 5147 4487
rect 5253 4473 5267 4487
rect 5293 4473 5307 4487
rect 5333 4473 5347 4487
rect 5633 4473 5647 4487
rect 5673 4473 5687 4487
rect 5953 4473 5967 4487
rect 5993 4473 6007 4487
rect 6273 4473 6287 4487
rect 6313 4473 6327 4487
rect 6533 4473 6547 4487
rect 6573 4473 6587 4487
rect 33 4453 47 4467
rect 173 4453 187 4467
rect 233 4453 247 4467
rect 273 4453 287 4467
rect 413 4453 427 4467
rect 453 4453 467 4467
rect 553 4453 567 4467
rect 593 4453 607 4467
rect 633 4453 647 4467
rect 713 4453 727 4467
rect 853 4453 867 4467
rect 993 4453 1007 4467
rect 1053 4453 1067 4467
rect 1193 4453 1207 4467
rect 1333 4453 1347 4467
rect 1493 4453 1507 4467
rect 1553 4453 1567 4467
rect 1993 4453 2007 4467
rect 2313 4453 2327 4467
rect 2533 4453 2547 4467
rect 2833 4453 2847 4467
rect 2873 4453 2887 4467
rect 2933 4453 2947 4467
rect 3013 4453 3027 4467
rect 3073 4453 3087 4467
rect 3113 4453 3127 4467
rect 3413 4453 3427 4467
rect 3453 4453 3467 4467
rect 3513 4453 3527 4467
rect 3553 4453 3567 4467
rect 3853 4453 3867 4467
rect 3893 4453 3907 4467
rect 4213 4453 4227 4467
rect 4253 4453 4267 4467
rect 4293 4453 4307 4467
rect 4333 4453 4347 4467
rect 4493 4453 4507 4467
rect 4533 4453 4547 4467
rect 4553 4453 4567 4467
rect 4593 4453 4607 4467
rect 4673 4453 4687 4467
rect 4733 4453 4747 4467
rect 4773 4453 4787 4467
rect 4833 4453 4847 4467
rect 4953 4453 4967 4467
rect 5033 4453 5047 4467
rect 5073 4453 5087 4467
rect 5113 4453 5127 4467
rect 5153 4453 5167 4467
rect 5213 4453 5227 4467
rect 5313 4453 5327 4467
rect 5353 4453 5367 4467
rect 5413 4453 5427 4467
rect 5493 4453 5507 4467
rect 5533 4453 5547 4467
rect 5573 4453 5587 4467
rect 5653 4453 5667 4467
rect 5693 4453 5707 4467
rect 5773 4453 5787 4467
rect 5853 4453 5867 4467
rect 5893 4453 5907 4467
rect 5933 4453 5947 4467
rect 5973 4453 5987 4467
rect 6033 4453 6047 4467
rect 6093 4453 6107 4467
rect 6133 4453 6147 4467
rect 6173 4453 6187 4467
rect 6253 4453 6267 4467
rect 6293 4453 6307 4467
rect 6333 4453 6347 4467
rect 6373 4453 6387 4467
rect 6433 4453 6447 4467
rect 6473 4453 6487 4467
rect 6553 4453 6567 4467
rect 6593 4453 6607 4467
rect 6653 4453 6667 4467
rect 1473 4433 1487 4447
rect 1513 4433 1527 4447
rect 1533 4433 1547 4447
rect 1573 4433 1587 4447
rect 1973 4433 1987 4447
rect 2013 4433 2027 4447
rect 2913 4433 2927 4447
rect 2953 4433 2967 4447
rect 4193 4433 4207 4447
rect 4233 4433 4247 4447
rect 4573 4433 4587 4447
rect 4613 4433 4627 4447
rect 4933 4433 4947 4447
rect 4973 4433 4987 4447
rect 5013 4433 5027 4447
rect 5053 4433 5067 4447
rect 5473 4433 5487 4447
rect 5513 4433 5527 4447
rect 5553 4433 5567 4447
rect 5593 4433 5607 4447
rect 5753 4433 5767 4447
rect 5793 4433 5807 4447
rect 5833 4433 5847 4447
rect 5873 4433 5887 4447
rect 6153 4433 6167 4447
rect 6193 4433 6207 4447
rect 6353 4433 6367 4447
rect 6393 4433 6407 4447
rect 6453 4433 6467 4447
rect 6493 4433 6507 4447
rect 533 4213 547 4227
rect 573 4213 587 4227
rect 1033 4213 1047 4227
rect 1073 4213 1087 4227
rect 1353 4213 1367 4227
rect 1393 4213 1407 4227
rect 1713 4213 1727 4227
rect 1753 4213 1767 4227
rect 1773 4213 1787 4227
rect 1813 4213 1827 4227
rect 2093 4213 2107 4227
rect 2133 4213 2147 4227
rect 2753 4213 2767 4227
rect 2793 4213 2807 4227
rect 3493 4213 3507 4227
rect 3533 4213 3547 4227
rect 3773 4213 3787 4227
rect 3813 4213 3827 4227
rect 3853 4213 3867 4227
rect 3893 4213 3907 4227
rect 3953 4213 3967 4227
rect 3993 4213 4007 4227
rect 5033 4213 5047 4227
rect 5073 4213 5087 4227
rect 5513 4213 5527 4227
rect 5553 4213 5567 4227
rect 5793 4213 5807 4227
rect 5873 4213 5887 4227
rect 5913 4213 5927 4227
rect 6193 4213 6207 4227
rect 6233 4213 6247 4227
rect 6313 4213 6327 4227
rect 6373 4213 6387 4227
rect 6413 4213 6427 4227
rect 6633 4213 6647 4227
rect 6673 4213 6687 4227
rect 113 4193 127 4207
rect 153 4193 167 4207
rect 213 4193 227 4207
rect 253 4193 267 4207
rect 553 4193 567 4207
rect 653 4193 667 4207
rect 693 4193 707 4207
rect 753 4193 767 4207
rect 1053 4193 1067 4207
rect 1373 4193 1387 4207
rect 1453 4193 1467 4207
rect 1513 4193 1527 4207
rect 1553 4193 1567 4207
rect 1633 4193 1647 4207
rect 1673 4193 1687 4207
rect 1733 4193 1747 4207
rect 1793 4193 1807 4207
rect 2113 4193 2127 4207
rect 2193 4193 2207 4207
rect 2233 4193 2247 4207
rect 2613 4193 2627 4207
rect 2673 4193 2687 4207
rect 2713 4193 2727 4207
rect 2773 4193 2787 4207
rect 2853 4193 2867 4207
rect 2893 4193 2907 4207
rect 2953 4193 2967 4207
rect 3093 4193 3107 4207
rect 3393 4193 3407 4207
rect 3433 4193 3447 4207
rect 3513 4193 3527 4207
rect 3593 4193 3607 4207
rect 3733 4193 3747 4207
rect 3793 4193 3807 4207
rect 3873 4193 3887 4207
rect 3973 4193 3987 4207
rect 4033 4193 4047 4207
rect 4093 4193 4107 4207
rect 4133 4193 4147 4207
rect 4193 4193 4207 4207
rect 4233 4193 4247 4207
rect 4533 4193 4547 4207
rect 4573 4193 4587 4207
rect 4893 4193 4907 4207
rect 4953 4193 4967 4207
rect 4993 4193 5007 4207
rect 5013 4193 5027 4207
rect 5053 4193 5067 4207
rect 5133 4193 5147 4207
rect 5193 4193 5207 4207
rect 5233 4193 5247 4207
rect 5533 4193 5547 4207
rect 5613 4193 5627 4207
rect 5673 4193 5687 4207
rect 5713 4193 5727 4207
rect 5853 4193 5867 4207
rect 5893 4193 5907 4207
rect 5993 4193 6007 4207
rect 6033 4193 6047 4207
rect 6073 4193 6087 4207
rect 6213 4193 6227 4207
rect 6393 4193 6407 4207
rect 6473 4193 6487 4207
rect 6553 4193 6567 4207
rect 6593 4193 6607 4207
rect 6613 4193 6627 4207
rect 6653 4193 6667 4207
rect 33 4173 47 4187
rect 73 4173 87 4187
rect 133 4173 147 4187
rect 173 4173 187 4187
rect 193 4173 207 4187
rect 233 4173 247 4187
rect 373 4173 387 4187
rect 413 4173 427 4187
rect 493 4173 507 4187
rect 633 4173 647 4187
rect 673 4173 687 4187
rect 713 4173 727 4187
rect 813 4173 827 4187
rect 893 4173 907 4187
rect 933 4173 947 4187
rect 1133 4173 1147 4187
rect 1213 4173 1227 4187
rect 1253 4173 1267 4187
rect 1533 4173 1547 4187
rect 1573 4173 1587 4187
rect 1613 4173 1627 4187
rect 1873 4173 1887 4187
rect 1953 4173 1967 4187
rect 1993 4173 2007 4187
rect 2213 4173 2227 4187
rect 2253 4173 2267 4187
rect 2353 4173 2367 4187
rect 2393 4173 2407 4187
rect 2473 4173 2487 4187
rect 2533 4173 2547 4187
rect 2573 4173 2587 4187
rect 2653 4173 2667 4187
rect 2693 4173 2707 4187
rect 2873 4173 2887 4187
rect 2913 4173 2927 4187
rect 2993 4173 3007 4187
rect 3033 4173 3047 4187
rect 3153 4173 3167 4187
rect 3233 4173 3247 4187
rect 3273 4173 3287 4187
rect 3373 4173 3387 4187
rect 3413 4173 3427 4187
rect 3453 4173 3467 4187
rect 4113 4173 4127 4187
rect 4153 4173 4167 4187
rect 4173 4173 4187 4187
rect 4213 4173 4227 4187
rect 4353 4173 4367 4187
rect 4393 4173 4407 4187
rect 4473 4173 4487 4187
rect 4553 4173 4567 4187
rect 4593 4173 4607 4187
rect 4693 4173 4707 4187
rect 4733 4173 4747 4187
rect 4813 4173 4827 4187
rect 4873 4173 4887 4187
rect 4933 4173 4947 4187
rect 5173 4173 5187 4187
rect 5213 4173 5227 4187
rect 5353 4173 5367 4187
rect 5393 4173 5407 4187
rect 5473 4173 5487 4187
rect 5653 4173 5667 4187
rect 5693 4173 5707 4187
rect 5773 4173 5787 4187
rect 5833 4173 5847 4187
rect 5973 4173 5987 4187
rect 6013 4173 6027 4187
rect 6053 4173 6067 4187
rect 6113 4173 6127 4187
rect 6153 4173 6167 4187
rect 6293 4173 6307 4187
rect 6353 4173 6367 4187
rect 6533 4173 6547 4187
rect 773 4153 787 4167
rect 1433 4153 1447 4167
rect 1653 4153 1667 4167
rect 2553 4153 2567 4167
rect 2593 4153 2607 4167
rect 2933 4153 2947 4167
rect 3013 4153 3027 4167
rect 3113 4153 3127 4167
rect 4013 4153 4027 4167
rect 4973 4153 4987 4167
rect 5153 4153 5167 4167
rect 5593 4153 5607 4167
rect 6453 4153 6467 4167
rect 6573 4153 6587 4167
rect 473 4013 487 4027
rect 1293 4013 1307 4027
rect 2433 4013 2447 4027
rect 2573 4013 2587 4027
rect 2673 4013 2687 4027
rect 2713 4013 2727 4027
rect 2813 4013 2827 4027
rect 2933 4013 2947 4027
rect 3093 4013 3107 4027
rect 3173 4013 3187 4027
rect 3673 4013 3687 4027
rect 4233 4013 4247 4027
rect 4333 4013 4347 4027
rect 5593 4013 5607 4027
rect 5853 4013 5867 4027
rect 33 3993 47 4007
rect 73 3993 87 4007
rect 113 3993 127 4007
rect 193 3993 207 4007
rect 233 3993 247 4007
rect 433 3993 447 4007
rect 693 3993 707 4007
rect 733 3993 747 4007
rect 773 3993 787 4007
rect 853 3993 867 4007
rect 893 3993 907 4007
rect 1253 3993 1267 4007
rect 1353 3993 1367 4007
rect 1433 3993 1447 4007
rect 1473 3993 1487 4007
rect 1653 3993 1667 4007
rect 1693 3993 1707 4007
rect 1833 3993 1847 4007
rect 1913 3993 1927 4007
rect 1953 3993 1967 4007
rect 2173 3993 2187 4007
rect 2213 3993 2227 4007
rect 2493 3993 2507 4007
rect 2533 3993 2547 4007
rect 2553 3993 2567 4007
rect 2593 3993 2607 4007
rect 2653 3993 2667 4007
rect 2693 3993 2707 4007
rect 2913 3993 2927 4007
rect 2953 3993 2967 4007
rect 2993 3993 3007 4007
rect 3033 3993 3047 4007
rect 3153 3993 3167 4007
rect 3193 3993 3207 4007
rect 3473 3993 3487 4007
rect 3513 3993 3527 4007
rect 3593 3993 3607 4007
rect 3773 3993 3787 4007
rect 3813 3993 3827 4007
rect 3893 3993 3907 4007
rect 4153 3993 4167 4007
rect 4193 3993 4207 4007
rect 4213 3993 4227 4007
rect 4253 3993 4267 4007
rect 4473 3993 4487 4007
rect 4513 3993 4527 4007
rect 4613 3993 4627 4007
rect 4653 3993 4667 4007
rect 4733 3993 4747 4007
rect 4893 3993 4907 4007
rect 4933 3993 4947 4007
rect 5033 3993 5047 4007
rect 5073 3993 5087 4007
rect 5153 3993 5167 4007
rect 5313 3993 5327 4007
rect 5353 3993 5367 4007
rect 5453 3993 5467 4007
rect 5493 3993 5507 4007
rect 5693 3993 5707 4007
rect 5733 3993 5747 4007
rect 5813 3993 5827 4007
rect 6033 3993 6047 4007
rect 6113 3993 6127 4007
rect 6153 3993 6167 4007
rect 6273 3993 6287 4007
rect 6353 3993 6367 4007
rect 6393 3993 6407 4007
rect 6513 3993 6527 4007
rect 6593 3993 6607 4007
rect 6633 3993 6647 4007
rect 353 3973 367 3987
rect 453 3973 467 3987
rect 493 3973 507 3987
rect 553 3973 567 3987
rect 633 3973 647 3987
rect 1033 3973 1047 3987
rect 1093 3973 1107 3987
rect 1173 3973 1187 3987
rect 1273 3973 1287 3987
rect 1313 3973 1327 3987
rect 1613 3973 1627 3987
rect 1753 3973 1767 3987
rect 2073 3973 2087 3987
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 2273 3973 2287 3987
rect 2333 3973 2347 3987
rect 2413 3973 2427 3987
rect 2473 3973 2487 3987
rect 2513 3973 2527 3987
rect 2733 3973 2747 3987
rect 2793 3973 2807 3987
rect 2873 3973 2887 3987
rect 3013 3973 3027 3987
rect 3053 3973 3067 3987
rect 3113 3973 3127 3987
rect 3273 3973 3287 3987
rect 3353 3973 3367 3987
rect 3653 3973 3667 3987
rect 3973 3973 3987 3987
rect 4013 3973 4027 3987
rect 4053 3973 4067 3987
rect 4133 3973 4147 3987
rect 4173 3973 4187 3987
rect 4313 3973 4327 3987
rect 4393 3973 4407 3987
rect 4453 3973 4467 3987
rect 4493 3973 4507 3987
rect 4813 3973 4827 3987
rect 4873 3973 4887 3987
rect 4913 3973 4927 3987
rect 5233 3973 5247 3987
rect 5293 3973 5307 3987
rect 5333 3973 5347 3987
rect 5413 3973 5427 3987
rect 5473 3973 5487 3987
rect 5513 3973 5527 3987
rect 5573 3973 5587 3987
rect 5873 3973 5887 3987
rect 5953 3973 5967 3987
rect 5993 3973 6007 3987
rect 333 3953 347 3967
rect 373 3953 387 3967
rect 533 3953 547 3967
rect 573 3953 587 3967
rect 613 3953 627 3967
rect 653 3953 667 3967
rect 1013 3953 1027 3967
rect 1053 3953 1067 3967
rect 1073 3953 1087 3967
rect 1113 3953 1127 3967
rect 1153 3953 1167 3967
rect 1193 3953 1207 3967
rect 1593 3953 1607 3967
rect 1633 3953 1647 3967
rect 1733 3953 1747 3967
rect 1773 3953 1787 3967
rect 2053 3953 2067 3967
rect 2093 3953 2107 3967
rect 2253 3953 2267 3967
rect 2293 3953 2307 3967
rect 2313 3953 2327 3967
rect 2353 3953 2367 3967
rect 2853 3953 2867 3967
rect 2893 3953 2907 3967
rect 3253 3953 3267 3967
rect 3293 3953 3307 3967
rect 3333 3953 3347 3967
rect 3373 3953 3387 3967
rect 3953 3953 3967 3967
rect 3993 3953 4007 3967
rect 4033 3953 4047 3967
rect 4073 3953 4087 3967
rect 4373 3953 4387 3967
rect 4413 3953 4427 3967
rect 4793 3953 4807 3967
rect 4833 3953 4847 3967
rect 5213 3953 5227 3967
rect 5253 3953 5267 3967
rect 5393 3953 5407 3967
rect 5433 3953 5447 3967
rect 5933 3953 5947 3967
rect 5973 3953 5987 3967
rect 193 3733 207 3747
rect 233 3733 247 3747
rect 613 3733 627 3747
rect 653 3733 667 3747
rect 673 3733 687 3747
rect 713 3733 727 3747
rect 773 3733 787 3747
rect 813 3733 827 3747
rect 1193 3733 1207 3747
rect 1233 3733 1247 3747
rect 1453 3733 1467 3747
rect 1493 3733 1507 3747
rect 1513 3733 1527 3747
rect 1553 3733 1567 3747
rect 1933 3733 1947 3747
rect 1973 3733 1987 3747
rect 2673 3733 2687 3747
rect 2713 3733 2727 3747
rect 2833 3733 2847 3747
rect 2873 3733 2887 3747
rect 3333 3733 3347 3747
rect 3373 3733 3387 3747
rect 3413 3733 3427 3747
rect 3453 3733 3467 3747
rect 3733 3733 3747 3747
rect 3773 3733 3787 3747
rect 3973 3733 3987 3747
rect 4013 3733 4027 3747
rect 4393 3733 4407 3747
rect 4433 3733 4447 3747
rect 4493 3733 4507 3747
rect 4533 3733 4547 3747
rect 5113 3733 5127 3747
rect 5153 3733 5167 3747
rect 5193 3733 5207 3747
rect 5233 3733 5247 3747
rect 5813 3733 5827 3747
rect 5853 3733 5867 3747
rect 5893 3733 5907 3747
rect 5933 3733 5947 3747
rect 6633 3733 6647 3747
rect 6673 3733 6687 3747
rect 213 3713 227 3727
rect 533 3713 547 3727
rect 573 3713 587 3727
rect 633 3713 647 3727
rect 693 3713 707 3727
rect 793 3713 807 3727
rect 1073 3713 1087 3727
rect 1113 3713 1127 3727
rect 1213 3713 1227 3727
rect 1373 3713 1387 3727
rect 1413 3713 1427 3727
rect 1473 3713 1487 3727
rect 1533 3713 1547 3727
rect 1953 3713 1967 3727
rect 2093 3713 2107 3727
rect 2153 3713 2167 3727
rect 2193 3713 2207 3727
rect 2253 3713 2267 3727
rect 2293 3713 2307 3727
rect 2373 3713 2387 3727
rect 2413 3713 2427 3727
rect 2453 3713 2467 3727
rect 2513 3713 2527 3727
rect 2573 3713 2587 3727
rect 2613 3713 2627 3727
rect 2653 3713 2667 3727
rect 2693 3713 2707 3727
rect 2773 3713 2787 3727
rect 2853 3713 2867 3727
rect 2913 3713 2927 3727
rect 2953 3713 2967 3727
rect 3013 3713 3027 3727
rect 3053 3713 3067 3727
rect 3093 3713 3107 3727
rect 3133 3713 3147 3727
rect 3233 3713 3247 3727
rect 3273 3713 3287 3727
rect 3353 3713 3367 3727
rect 3433 3713 3447 3727
rect 3753 3713 3767 3727
rect 3833 3713 3847 3727
rect 3873 3713 3887 3727
rect 3933 3713 3947 3727
rect 3993 3713 4007 3727
rect 4073 3713 4087 3727
rect 4113 3713 4127 3727
rect 4413 3713 4427 3727
rect 4513 3713 4527 3727
rect 4573 3713 4587 3727
rect 4713 3713 4727 3727
rect 5013 3713 5027 3727
rect 5053 3713 5067 3727
rect 5133 3713 5147 3727
rect 5213 3713 5227 3727
rect 5273 3713 5287 3727
rect 5333 3713 5347 3727
rect 5473 3713 5487 3727
rect 5773 3713 5787 3727
rect 5833 3713 5847 3727
rect 5913 3713 5927 3727
rect 5993 3713 6007 3727
rect 6193 3713 6207 3727
rect 6233 3713 6247 3727
rect 6553 3713 6567 3727
rect 6593 3713 6607 3727
rect 6653 3713 6667 3727
rect 33 3693 47 3707
rect 73 3693 87 3707
rect 113 3693 127 3707
rect 153 3693 167 3707
rect 273 3693 287 3707
rect 353 3693 367 3707
rect 393 3693 407 3707
rect 513 3693 527 3707
rect 853 3693 867 3707
rect 933 3693 947 3707
rect 973 3693 987 3707
rect 1133 3693 1147 3707
rect 1253 3693 1267 3707
rect 1293 3693 1307 3707
rect 1353 3693 1367 3707
rect 1593 3693 1607 3707
rect 1633 3693 1647 3707
rect 1693 3693 1707 3707
rect 1773 3693 1787 3707
rect 1813 3693 1827 3707
rect 1993 3693 2007 3707
rect 2033 3693 2047 3707
rect 2133 3693 2147 3707
rect 2173 3693 2187 3707
rect 2273 3693 2287 3707
rect 2313 3693 2327 3707
rect 2353 3693 2367 3707
rect 2553 3693 2567 3707
rect 2593 3693 2607 3707
rect 2893 3693 2907 3707
rect 2933 3693 2947 3707
rect 2993 3693 3007 3707
rect 3033 3693 3047 3707
rect 3153 3693 3167 3707
rect 3213 3693 3227 3707
rect 3253 3693 3267 3707
rect 3293 3693 3307 3707
rect 3553 3693 3567 3707
rect 3593 3693 3607 3707
rect 3673 3693 3687 3707
rect 3813 3693 3827 3707
rect 3853 3693 3867 3707
rect 3893 3693 3907 3707
rect 4053 3693 4067 3707
rect 4093 3693 4107 3707
rect 4233 3693 4247 3707
rect 4273 3693 4287 3707
rect 4353 3693 4367 3707
rect 4833 3693 4847 3707
rect 4873 3693 4887 3707
rect 4953 3693 4967 3707
rect 4993 3693 5007 3707
rect 5033 3693 5047 3707
rect 5533 3693 5547 3707
rect 5613 3693 5627 3707
rect 5653 3693 5667 3707
rect 6033 3693 6047 3707
rect 6073 3693 6087 3707
rect 6133 3693 6147 3707
rect 6173 3693 6187 3707
rect 6253 3693 6267 3707
rect 6313 3693 6327 3707
rect 6393 3693 6407 3707
rect 6433 3693 6447 3707
rect 6533 3693 6547 3707
rect 6573 3693 6587 3707
rect 553 3673 567 3687
rect 1093 3673 1107 3687
rect 1393 3673 1407 3687
rect 1613 3673 1627 3687
rect 2013 3673 2027 3687
rect 2073 3673 2087 3687
rect 2393 3673 2407 3687
rect 2433 3673 2447 3687
rect 2533 3673 2547 3687
rect 2793 3673 2807 3687
rect 3113 3673 3127 3687
rect 3913 3673 3927 3687
rect 5293 3673 5307 3687
rect 5793 3673 5807 3687
rect 6013 3673 6027 3687
rect 6053 3673 6067 3687
rect 6153 3673 6167 3687
rect 6213 3673 6227 3687
rect 553 3533 567 3547
rect 1033 3533 1047 3547
rect 1493 3533 1507 3547
rect 1913 3533 1927 3547
rect 2053 3533 2067 3547
rect 2153 3533 2167 3547
rect 2313 3533 2327 3547
rect 2613 3533 2627 3547
rect 2813 3533 2827 3547
rect 3033 3533 3047 3547
rect 3333 3533 3347 3547
rect 3993 3533 4007 3547
rect 4293 3533 4307 3547
rect 4353 3533 4367 3547
rect 4733 3533 4747 3547
rect 5153 3533 5167 3547
rect 5893 3533 5907 3547
rect 6153 3533 6167 3547
rect 6393 3533 6407 3547
rect 33 3513 47 3527
rect 73 3513 87 3527
rect 113 3513 127 3527
rect 193 3513 207 3527
rect 233 3513 247 3527
rect 413 3513 427 3527
rect 453 3513 467 3527
rect 513 3513 527 3527
rect 693 3513 707 3527
rect 733 3513 747 3527
rect 753 3513 767 3527
rect 793 3513 807 3527
rect 933 3513 947 3527
rect 973 3513 987 3527
rect 1073 3513 1087 3527
rect 1113 3513 1127 3527
rect 1153 3513 1167 3527
rect 1193 3513 1207 3527
rect 1233 3513 1247 3527
rect 1313 3513 1327 3527
rect 1353 3513 1367 3527
rect 1473 3513 1487 3527
rect 1513 3513 1527 3527
rect 1553 3513 1567 3527
rect 1633 3513 1647 3527
rect 1673 3513 1687 3527
rect 1793 3513 1807 3527
rect 1853 3513 1867 3527
rect 1973 3513 1987 3527
rect 2013 3513 2027 3527
rect 2033 3513 2047 3527
rect 2073 3513 2087 3527
rect 2193 3513 2207 3527
rect 2253 3513 2267 3527
rect 2293 3513 2307 3527
rect 2333 3513 2347 3527
rect 2373 3513 2387 3527
rect 2453 3513 2467 3527
rect 2493 3513 2507 3527
rect 2593 3513 2607 3527
rect 2633 3513 2647 3527
rect 2673 3513 2687 3527
rect 2713 3513 2727 3527
rect 2913 3513 2927 3527
rect 2953 3513 2967 3527
rect 3073 3513 3087 3527
rect 3133 3513 3147 3527
rect 3193 3513 3207 3527
rect 3233 3513 3247 3527
rect 3273 3513 3287 3527
rect 3373 3513 3387 3527
rect 3453 3513 3467 3527
rect 3493 3513 3507 3527
rect 3613 3513 3627 3527
rect 3653 3513 3667 3527
rect 3693 3513 3707 3527
rect 3733 3513 3747 3527
rect 3813 3513 3827 3527
rect 3853 3513 3867 3527
rect 4033 3513 4047 3527
rect 4113 3513 4127 3527
rect 4153 3513 4167 3527
rect 4533 3513 4547 3527
rect 4573 3513 4587 3527
rect 4653 3513 4667 3527
rect 4773 3513 4787 3527
rect 4853 3513 4867 3527
rect 4893 3513 4907 3527
rect 5013 3513 5027 3527
rect 5053 3513 5067 3527
rect 5093 3513 5107 3527
rect 5193 3513 5207 3527
rect 5273 3513 5287 3527
rect 5313 3513 5327 3527
rect 5433 3513 5447 3527
rect 5513 3513 5527 3527
rect 5553 3513 5567 3527
rect 5653 3513 5667 3527
rect 5693 3513 5707 3527
rect 5753 3513 5767 3527
rect 5793 3513 5807 3527
rect 5933 3513 5947 3527
rect 5973 3513 5987 3527
rect 6013 3513 6027 3527
rect 6193 3513 6207 3527
rect 6253 3513 6267 3527
rect 6433 3513 6447 3527
rect 6513 3513 6527 3527
rect 6553 3513 6567 3527
rect 353 3493 367 3507
rect 533 3493 547 3507
rect 573 3493 587 3507
rect 633 3493 647 3507
rect 853 3493 867 3507
rect 1013 3493 1027 3507
rect 1893 3493 1907 3507
rect 1953 3493 1967 3507
rect 1993 3493 2007 3507
rect 2133 3493 2147 3507
rect 2693 3493 2707 3507
rect 2733 3493 2747 3507
rect 2793 3493 2807 3507
rect 2873 3493 2887 3507
rect 2933 3493 2947 3507
rect 2973 3493 2987 3507
rect 3013 3493 3027 3507
rect 3053 3493 3067 3507
rect 3113 3493 3127 3507
rect 3213 3493 3227 3507
rect 3253 3493 3267 3507
rect 3313 3493 3327 3507
rect 3633 3493 3647 3507
rect 3673 3493 3687 3507
rect 3973 3493 3987 3507
rect 4273 3493 4287 3507
rect 4333 3493 4347 3507
rect 4393 3493 4407 3507
rect 4713 3493 4727 3507
rect 5033 3493 5047 3507
rect 5073 3493 5087 3507
rect 5133 3493 5147 3507
rect 5673 3493 5687 3507
rect 5713 3493 5727 3507
rect 5773 3493 5787 3507
rect 5813 3493 5827 3507
rect 5873 3493 5887 3507
rect 5953 3493 5967 3507
rect 5993 3493 6007 3507
rect 6053 3493 6067 3507
rect 6133 3493 6147 3507
rect 6233 3493 6247 3507
rect 6293 3493 6307 3507
rect 6373 3493 6387 3507
rect 333 3473 347 3487
rect 373 3473 387 3487
rect 613 3473 627 3487
rect 653 3473 667 3487
rect 833 3473 847 3487
rect 873 3473 887 3487
rect 1813 3473 1827 3487
rect 2213 3473 2227 3487
rect 2853 3473 2867 3487
rect 2893 3473 2907 3487
rect 4373 3473 4387 3487
rect 4413 3473 4427 3487
rect 6033 3473 6047 3487
rect 6073 3473 6087 3487
rect 333 3253 347 3267
rect 373 3253 387 3267
rect 533 3253 547 3267
rect 573 3253 587 3267
rect 673 3253 687 3267
rect 713 3253 727 3267
rect 753 3253 767 3267
rect 793 3253 807 3267
rect 1273 3253 1287 3267
rect 1313 3253 1327 3267
rect 1633 3253 1647 3267
rect 1813 3253 1827 3267
rect 1853 3253 1867 3267
rect 2233 3253 2247 3267
rect 2273 3253 2287 3267
rect 2873 3253 2887 3267
rect 2913 3253 2927 3267
rect 2973 3253 2987 3267
rect 3013 3253 3027 3267
rect 3153 3253 3167 3267
rect 3193 3253 3207 3267
rect 6153 3253 6167 3267
rect 6193 3253 6207 3267
rect 6333 3253 6347 3267
rect 6373 3253 6387 3267
rect 353 3233 367 3247
rect 453 3233 467 3247
rect 493 3233 507 3247
rect 553 3233 567 3247
rect 613 3233 627 3247
rect 653 3233 667 3247
rect 693 3233 707 3247
rect 773 3233 787 3247
rect 853 3233 867 3247
rect 893 3233 907 3247
rect 953 3233 967 3247
rect 1093 3233 1107 3247
rect 1133 3233 1147 3247
rect 1193 3233 1207 3247
rect 1233 3233 1247 3247
rect 1293 3233 1307 3247
rect 1733 3233 1747 3247
rect 1773 3233 1787 3247
rect 1833 3233 1847 3247
rect 1873 3233 1887 3247
rect 1893 3233 1907 3247
rect 1933 3233 1947 3247
rect 2253 3233 2267 3247
rect 2493 3233 2507 3247
rect 2533 3233 2547 3247
rect 2593 3233 2607 3247
rect 2893 3233 2907 3247
rect 2993 3233 3007 3247
rect 3053 3233 3067 3247
rect 3093 3233 3107 3247
rect 3173 3233 3187 3247
rect 3233 3233 3247 3247
rect 3293 3233 3307 3247
rect 3333 3233 3347 3247
rect 3393 3233 3407 3247
rect 3553 3233 3567 3247
rect 3593 3233 3607 3247
rect 3953 3233 3967 3247
rect 3993 3233 4007 3247
rect 4093 3233 4107 3247
rect 4133 3233 4147 3247
rect 4513 3233 4527 3247
rect 4553 3233 4567 3247
rect 4793 3233 4807 3247
rect 4853 3233 4867 3247
rect 4893 3233 4907 3247
rect 4953 3233 4967 3247
rect 4993 3233 5007 3247
rect 5313 3233 5327 3247
rect 5353 3233 5367 3247
rect 5413 3233 5427 3247
rect 5493 3233 5507 3247
rect 5793 3233 5807 3247
rect 5833 3233 5847 3247
rect 5893 3233 5907 3247
rect 5973 3233 5987 3247
rect 6013 3233 6027 3247
rect 6053 3233 6067 3247
rect 6093 3233 6107 3247
rect 6173 3233 6187 3247
rect 6253 3233 6267 3247
rect 6293 3233 6307 3247
rect 6353 3233 6367 3247
rect 6413 3233 6427 3247
rect 6453 3233 6467 3247
rect 33 3213 47 3227
rect 73 3213 87 3227
rect 113 3213 127 3227
rect 193 3213 207 3227
rect 233 3213 247 3227
rect 433 3213 447 3227
rect 873 3213 887 3227
rect 913 3213 927 3227
rect 993 3213 1007 3227
rect 1033 3213 1047 3227
rect 1073 3213 1087 3227
rect 1113 3213 1127 3227
rect 1173 3213 1187 3227
rect 1213 3213 1227 3227
rect 1373 3213 1387 3227
rect 1453 3213 1467 3227
rect 1493 3213 1507 3227
rect 1613 3213 1627 3227
rect 1673 3213 1687 3227
rect 1713 3213 1727 3227
rect 1953 3213 1967 3227
rect 2073 3213 2087 3227
rect 2113 3213 2127 3227
rect 2193 3213 2207 3227
rect 2313 3213 2327 3227
rect 2353 3213 2367 3227
rect 2413 3213 2427 3227
rect 2453 3213 2467 3227
rect 2513 3213 2527 3227
rect 2553 3213 2567 3227
rect 2713 3213 2727 3227
rect 2753 3213 2767 3227
rect 2833 3213 2847 3227
rect 3073 3213 3087 3227
rect 3113 3213 3127 3227
rect 3313 3213 3327 3227
rect 3353 3213 3367 3227
rect 3453 3213 3467 3227
rect 3493 3213 3507 3227
rect 3533 3213 3547 3227
rect 3633 3213 3647 3227
rect 3673 3213 3687 3227
rect 3713 3213 3727 3227
rect 3793 3213 3807 3227
rect 3833 3213 3847 3227
rect 3933 3213 3947 3227
rect 3973 3213 3987 3227
rect 4013 3213 4027 3227
rect 4073 3213 4087 3227
rect 4113 3213 4127 3227
rect 4153 3213 4167 3227
rect 4253 3213 4267 3227
rect 4293 3213 4307 3227
rect 4373 3213 4387 3227
rect 4413 3213 4427 3227
rect 4453 3213 4467 3227
rect 4493 3213 4507 3227
rect 4533 3213 4547 3227
rect 4573 3213 4587 3227
rect 4613 3213 4627 3227
rect 4653 3213 4667 3227
rect 4693 3213 4707 3227
rect 4733 3213 4747 3227
rect 4833 3213 4847 3227
rect 4873 3213 4887 3227
rect 4913 3213 4927 3227
rect 5013 3213 5027 3227
rect 5073 3213 5087 3227
rect 5153 3213 5167 3227
rect 5193 3213 5207 3227
rect 5373 3213 5387 3227
rect 5433 3213 5447 3227
rect 5613 3213 5627 3227
rect 5653 3213 5667 3227
rect 5733 3213 5747 3227
rect 5813 3213 5827 3227
rect 5853 3213 5867 3227
rect 5953 3213 5967 3227
rect 6033 3213 6047 3227
rect 6073 3213 6087 3227
rect 6233 3213 6247 3227
rect 6393 3213 6407 3227
rect 6433 3213 6447 3227
rect 6513 3213 6527 3227
rect 6593 3213 6607 3227
rect 6633 3213 6647 3227
rect 473 3193 487 3207
rect 593 3193 607 3207
rect 933 3193 947 3207
rect 1013 3193 1027 3207
rect 1753 3193 1767 3207
rect 1913 3193 1927 3207
rect 2333 3193 2347 3207
rect 2433 3193 2447 3207
rect 2573 3193 2587 3207
rect 3253 3193 3267 3207
rect 3373 3193 3387 3207
rect 3473 3193 3487 3207
rect 3573 3193 3587 3207
rect 3653 3193 3667 3207
rect 4433 3193 4447 3207
rect 4633 3193 4647 3207
rect 4713 3193 4727 3207
rect 4773 3193 4787 3207
rect 4973 3193 4987 3207
rect 5333 3193 5347 3207
rect 5513 3193 5527 3207
rect 5913 3193 5927 3207
rect 5993 3193 6007 3207
rect 6273 3193 6287 3207
rect 973 3053 987 3067
rect 1653 3053 1667 3067
rect 1813 3053 1827 3067
rect 2113 3053 2127 3067
rect 2273 3053 2287 3067
rect 2633 3053 2647 3067
rect 2713 3053 2727 3067
rect 2813 3053 2827 3067
rect 4673 3053 4687 3067
rect 4973 3053 4987 3067
rect 5113 3053 5127 3067
rect 5193 3053 5207 3067
rect 5533 3053 5547 3067
rect 5893 3053 5907 3067
rect 6133 3053 6147 3067
rect 6213 3053 6227 3067
rect 6253 3053 6267 3067
rect 6473 3053 6487 3067
rect 6493 3053 6507 3067
rect 233 3033 247 3047
rect 273 3033 287 3047
rect 373 3033 387 3047
rect 413 3033 427 3047
rect 493 3033 507 3047
rect 733 3033 747 3047
rect 773 3033 787 3047
rect 1013 3033 1027 3047
rect 1073 3033 1087 3047
rect 1153 3033 1167 3047
rect 1193 3033 1207 3047
rect 1393 3033 1407 3047
rect 1473 3033 1487 3047
rect 1513 3033 1527 3047
rect 1713 3033 1727 3047
rect 1753 3033 1767 3047
rect 1793 3033 1807 3047
rect 1833 3033 1847 3047
rect 1873 3033 1887 3047
rect 1933 3033 1947 3047
rect 1953 3033 1967 3047
rect 1993 3033 2007 3047
rect 2073 3033 2087 3047
rect 2293 3033 2307 3047
rect 2353 3033 2367 3047
rect 2473 3033 2487 3047
rect 2513 3033 2527 3047
rect 2593 3033 2607 3047
rect 2693 3033 2707 3047
rect 2733 3033 2747 3047
rect 2873 3033 2887 3047
rect 2913 3033 2927 3047
rect 2953 3033 2967 3047
rect 3213 3033 3227 3047
rect 3253 3033 3267 3047
rect 3433 3033 3447 3047
rect 3473 3033 3487 3047
rect 3533 3033 3547 3047
rect 3593 3033 3607 3047
rect 3653 3033 3667 3047
rect 3693 3033 3707 3047
rect 3733 3033 3747 3047
rect 3913 3033 3927 3047
rect 3953 3033 3967 3047
rect 4033 3033 4047 3047
rect 4073 3033 4087 3047
rect 4113 3033 4127 3047
rect 4353 3033 4367 3047
rect 4393 3033 4407 3047
rect 4473 3033 4487 3047
rect 4533 3033 4547 3047
rect 4573 3033 4587 3047
rect 4613 3033 4627 3047
rect 4713 3033 4727 3047
rect 4773 3033 4787 3047
rect 4813 3033 4827 3047
rect 4853 3033 4867 3047
rect 4893 3033 4907 3047
rect 4993 3033 5007 3047
rect 5033 3033 5047 3047
rect 5073 3033 5087 3047
rect 5173 3033 5187 3047
rect 5213 3033 5227 3047
rect 5333 3033 5347 3047
rect 5373 3033 5387 3047
rect 5453 3033 5467 3047
rect 5513 3033 5527 3047
rect 5553 3033 5567 3047
rect 5573 3033 5587 3047
rect 5613 3033 5627 3047
rect 5793 3033 5807 3047
rect 5833 3033 5847 3047
rect 5873 3033 5887 3047
rect 5973 3033 5987 3047
rect 6033 3033 6047 3047
rect 6093 3033 6107 3047
rect 6193 3033 6207 3047
rect 6233 3033 6247 3047
rect 6333 3033 6347 3047
rect 6373 3033 6387 3047
rect 6413 3033 6427 3047
rect 6553 3033 6567 3047
rect 6593 3033 6607 3047
rect 33 3013 47 3027
rect 173 3013 187 3027
rect 573 3013 587 3027
rect 633 3013 647 3027
rect 713 3013 727 3027
rect 753 3013 767 3027
rect 833 3013 847 3027
rect 913 3013 927 3027
rect 953 3013 967 3027
rect 993 3013 1007 3027
rect 1333 3013 1347 3027
rect 1633 3013 1647 3027
rect 1693 3013 1707 3027
rect 1733 3013 1747 3027
rect 1973 3013 1987 3027
rect 2013 3013 2027 3027
rect 2093 3013 2107 3027
rect 2133 3013 2147 3027
rect 2173 3013 2187 3027
rect 2253 3013 2267 3027
rect 2653 3013 2667 3027
rect 2793 3013 2807 3027
rect 2853 3013 2867 3027
rect 2893 3013 2907 3027
rect 2933 3013 2947 3027
rect 3033 3013 3047 3027
rect 3073 3013 3087 3027
rect 3133 3013 3147 3027
rect 3193 3013 3207 3027
rect 3233 3013 3247 3027
rect 3293 3013 3307 3027
rect 3373 3013 3387 3027
rect 3453 3013 3467 3027
rect 3493 3013 3507 3027
rect 3673 3013 3687 3027
rect 3713 3013 3727 3027
rect 3773 3013 3787 3027
rect 3813 3013 3827 3027
rect 4093 3013 4107 3027
rect 4133 3013 4147 3027
rect 4213 3013 4227 3027
rect 4253 3013 4267 3027
rect 4553 3013 4567 3027
rect 4593 3013 4607 3027
rect 4653 3013 4667 3027
rect 4733 3013 4747 3027
rect 4793 3013 4807 3027
rect 4833 3013 4847 3027
rect 4873 3013 4887 3027
rect 4953 3013 4967 3027
rect 5013 3013 5027 3027
rect 5053 3013 5067 3027
rect 5133 3013 5147 3027
rect 5593 3013 5607 3027
rect 5633 3013 5647 3027
rect 5713 3013 5727 3027
rect 5753 3013 5767 3027
rect 5813 3013 5827 3027
rect 5853 3013 5867 3027
rect 5913 3013 5927 3027
rect 5953 3013 5967 3027
rect 6013 3013 6027 3027
rect 6113 3013 6127 3027
rect 6153 3013 6167 3027
rect 6273 3013 6287 3027
rect 6353 3013 6367 3027
rect 6393 3013 6407 3027
rect 6453 3013 6467 3027
rect 6513 3013 6527 3027
rect 6573 3013 6587 3027
rect 6613 3013 6627 3027
rect 553 2993 567 3007
rect 593 2993 607 3007
rect 613 2993 627 3007
rect 653 2993 667 3007
rect 813 2993 827 3007
rect 853 2993 867 3007
rect 893 2993 907 3007
rect 933 2993 947 3007
rect 1313 2993 1327 3007
rect 1353 2993 1367 3007
rect 1893 2993 1907 3007
rect 2153 2993 2167 3007
rect 2193 2993 2207 3007
rect 2333 2993 2347 3007
rect 3013 2993 3027 3007
rect 3053 2993 3067 3007
rect 3113 2993 3127 3007
rect 3153 2993 3167 3007
rect 3273 2993 3287 3007
rect 3313 2993 3327 3007
rect 3353 2993 3367 3007
rect 3393 2993 3407 3007
rect 3573 2993 3587 3007
rect 4193 2993 4207 3007
rect 4233 2993 4247 3007
rect 5693 2993 5707 3007
rect 5733 2993 5747 3007
rect 933 2773 947 2787
rect 973 2773 987 2787
rect 1013 2773 1027 2787
rect 1053 2773 1067 2787
rect 1613 2773 1627 2787
rect 1653 2773 1667 2787
rect 2413 2773 2427 2787
rect 2453 2773 2467 2787
rect 4353 2773 4367 2787
rect 4393 2773 4407 2787
rect 6213 2773 6227 2787
rect 6393 2773 6407 2787
rect 33 2753 47 2767
rect 413 2753 427 2767
rect 853 2753 867 2767
rect 893 2753 907 2767
rect 953 2753 967 2767
rect 1033 2753 1047 2767
rect 1113 2753 1127 2767
rect 1173 2753 1187 2767
rect 1213 2753 1227 2767
rect 1313 2753 1327 2767
rect 1353 2753 1367 2767
rect 1393 2753 1407 2767
rect 1453 2753 1467 2767
rect 1493 2753 1507 2767
rect 1633 2753 1647 2767
rect 1793 2753 1807 2767
rect 1833 2753 1847 2767
rect 1933 2753 1947 2767
rect 1993 2753 2007 2767
rect 2033 2753 2047 2767
rect 2113 2753 2127 2767
rect 2153 2753 2167 2767
rect 2433 2753 2447 2767
rect 2513 2753 2527 2767
rect 2573 2753 2587 2767
rect 2873 2753 2887 2767
rect 2913 2753 2927 2767
rect 2993 2753 3007 2767
rect 3033 2753 3047 2767
rect 3313 2753 3327 2767
rect 3373 2753 3387 2767
rect 3413 2753 3427 2767
rect 3493 2753 3507 2767
rect 3533 2753 3547 2767
rect 3613 2753 3627 2767
rect 3653 2753 3667 2767
rect 3713 2753 3727 2767
rect 3753 2753 3767 2767
rect 3833 2753 3847 2767
rect 3873 2753 3887 2767
rect 3933 2753 3947 2767
rect 4173 2753 4187 2767
rect 4213 2753 4227 2767
rect 4253 2753 4267 2767
rect 4293 2753 4307 2767
rect 4373 2753 4387 2767
rect 4413 2753 4427 2767
rect 4693 2753 4707 2767
rect 4833 2753 4847 2767
rect 4873 2753 4887 2767
rect 5033 2753 5047 2767
rect 5073 2753 5087 2767
rect 5113 2753 5127 2767
rect 5153 2753 5167 2767
rect 5313 2753 5327 2767
rect 5353 2753 5367 2767
rect 5433 2753 5447 2767
rect 5473 2753 5487 2767
rect 5533 2753 5547 2767
rect 5813 2753 5827 2767
rect 5873 2753 5887 2767
rect 5933 2753 5947 2767
rect 5993 2753 6007 2767
rect 6053 2753 6067 2767
rect 6113 2753 6127 2767
rect 6293 2753 6307 2767
rect 6333 2753 6347 2767
rect 93 2733 107 2747
rect 133 2733 147 2747
rect 233 2733 247 2747
rect 273 2733 287 2747
rect 353 2733 367 2747
rect 473 2733 487 2747
rect 513 2733 527 2747
rect 613 2733 627 2747
rect 653 2733 667 2747
rect 733 2733 747 2747
rect 793 2733 807 2747
rect 833 2733 847 2747
rect 1153 2733 1167 2747
rect 1193 2733 1207 2747
rect 1233 2733 1247 2747
rect 1293 2733 1307 2747
rect 1473 2733 1487 2747
rect 1513 2733 1527 2747
rect 1533 2733 1547 2747
rect 1573 2733 1587 2747
rect 1693 2733 1707 2747
rect 1733 2733 1747 2747
rect 1813 2733 1827 2747
rect 1853 2733 1867 2747
rect 1893 2733 1907 2747
rect 1973 2733 1987 2747
rect 2013 2733 2027 2747
rect 2093 2733 2107 2747
rect 2253 2733 2267 2747
rect 2293 2733 2307 2747
rect 2373 2733 2387 2747
rect 2693 2733 2707 2747
rect 2733 2733 2747 2747
rect 2813 2733 2827 2747
rect 2853 2733 2867 2747
rect 2893 2733 2907 2747
rect 2973 2733 2987 2747
rect 3073 2733 3087 2747
rect 3153 2733 3167 2747
rect 3193 2733 3207 2747
rect 3353 2733 3367 2747
rect 3393 2733 3407 2747
rect 3433 2733 3447 2747
rect 3473 2733 3487 2747
rect 3513 2733 3527 2747
rect 3593 2733 3607 2747
rect 3633 2733 3647 2747
rect 3673 2733 3687 2747
rect 3693 2733 3707 2747
rect 3733 2733 3747 2747
rect 3813 2733 3827 2747
rect 3853 2733 3867 2747
rect 3893 2733 3907 2747
rect 3973 2733 3987 2747
rect 4013 2733 4027 2747
rect 4053 2733 4067 2747
rect 4093 2733 4107 2747
rect 4153 2733 4167 2747
rect 4233 2733 4247 2747
rect 4273 2733 4287 2747
rect 4513 2733 4527 2747
rect 4553 2733 4567 2747
rect 4633 2733 4647 2747
rect 4733 2733 4747 2747
rect 4773 2733 4787 2747
rect 4813 2733 4827 2747
rect 4853 2733 4867 2747
rect 4933 2733 4947 2747
rect 4973 2733 4987 2747
rect 5013 2733 5027 2747
rect 5053 2733 5067 2747
rect 5093 2733 5107 2747
rect 5173 2733 5187 2747
rect 5213 2733 5227 2747
rect 5253 2733 5267 2747
rect 5293 2733 5307 2747
rect 5333 2733 5347 2747
rect 5413 2733 5427 2747
rect 5453 2733 5467 2747
rect 5493 2733 5507 2747
rect 5653 2733 5667 2747
rect 5693 2733 5707 2747
rect 5773 2733 5787 2747
rect 5833 2733 5847 2747
rect 5893 2733 5907 2747
rect 5953 2733 5967 2747
rect 6013 2733 6027 2747
rect 6073 2733 6087 2747
rect 6133 2733 6147 2747
rect 6193 2733 6207 2747
rect 6253 2733 6267 2747
rect 6353 2733 6367 2747
rect 6413 2733 6427 2747
rect 6473 2733 6487 2747
rect 6553 2733 6567 2747
rect 6593 2733 6607 2747
rect 13 2713 27 2727
rect 113 2713 127 2727
rect 393 2713 407 2727
rect 493 2713 507 2727
rect 1093 2713 1107 2727
rect 1333 2713 1347 2727
rect 1413 2713 1427 2727
rect 1553 2713 1567 2727
rect 1713 2713 1727 2727
rect 1873 2713 1887 2727
rect 2133 2713 2147 2727
rect 2493 2713 2507 2727
rect 2593 2713 2607 2727
rect 3013 2713 3027 2727
rect 3293 2713 3307 2727
rect 3953 2713 3967 2727
rect 3993 2713 4007 2727
rect 4073 2713 4087 2727
rect 4193 2713 4207 2727
rect 4673 2713 4687 2727
rect 4753 2713 4767 2727
rect 4953 2713 4967 2727
rect 5133 2713 5147 2727
rect 5553 2713 5567 2727
rect 633 2573 647 2587
rect 1373 2573 1387 2587
rect 1433 2573 1447 2587
rect 1833 2573 1847 2587
rect 1893 2573 1907 2587
rect 2093 2573 2107 2587
rect 2793 2573 2807 2587
rect 3113 2573 3127 2587
rect 3393 2573 3407 2587
rect 3533 2573 3547 2587
rect 4013 2573 4027 2587
rect 4133 2573 4147 2587
rect 4573 2573 4587 2587
rect 5073 2573 5087 2587
rect 5373 2573 5387 2587
rect 5473 2573 5487 2587
rect 5753 2573 5767 2587
rect 6053 2573 6067 2587
rect 6513 2573 6527 2587
rect 33 2553 47 2567
rect 113 2553 127 2567
rect 153 2553 167 2567
rect 273 2553 287 2567
rect 313 2553 327 2567
rect 353 2553 367 2567
rect 433 2553 447 2567
rect 473 2553 487 2567
rect 593 2553 607 2567
rect 1053 2553 1067 2567
rect 1133 2553 1147 2567
rect 1173 2553 1187 2567
rect 1353 2553 1367 2567
rect 1393 2553 1407 2567
rect 1533 2553 1547 2567
rect 1573 2553 1587 2567
rect 1673 2553 1687 2567
rect 1713 2553 1727 2567
rect 1793 2553 1807 2567
rect 1953 2553 1967 2567
rect 1993 2553 2007 2567
rect 2033 2553 2047 2567
rect 2073 2553 2087 2567
rect 2113 2553 2127 2567
rect 2173 2553 2187 2567
rect 2233 2553 2247 2567
rect 2293 2553 2307 2567
rect 2353 2553 2367 2567
rect 2473 2553 2487 2567
rect 2513 2553 2527 2567
rect 2593 2553 2607 2567
rect 2653 2553 2667 2567
rect 2713 2553 2727 2567
rect 2773 2553 2787 2567
rect 2813 2553 2827 2567
rect 2853 2553 2867 2567
rect 2913 2553 2927 2567
rect 2973 2553 2987 2567
rect 3013 2553 3027 2567
rect 3053 2553 3067 2567
rect 3213 2553 3227 2567
rect 3253 2553 3267 2567
rect 3333 2553 3347 2567
rect 3373 2553 3387 2567
rect 3413 2553 3427 2567
rect 3893 2553 3907 2567
rect 3933 2553 3947 2567
rect 4053 2553 4067 2567
rect 4113 2553 4127 2567
rect 4153 2553 4167 2567
rect 4193 2553 4207 2567
rect 4233 2553 4247 2567
rect 4273 2553 4287 2567
rect 4373 2553 4387 2567
rect 4413 2553 4427 2567
rect 4493 2553 4507 2567
rect 4613 2553 4627 2567
rect 4653 2553 4667 2567
rect 4693 2553 4707 2567
rect 4733 2553 4747 2567
rect 4793 2553 4807 2567
rect 4853 2553 4867 2567
rect 4933 2553 4947 2567
rect 4973 2553 4987 2567
rect 5133 2553 5147 2567
rect 5173 2553 5187 2567
rect 5213 2553 5227 2567
rect 5253 2553 5267 2567
rect 5293 2553 5307 2567
rect 5353 2553 5367 2567
rect 5393 2553 5407 2567
rect 5453 2553 5467 2567
rect 5493 2553 5507 2567
rect 5733 2553 5747 2567
rect 5773 2553 5787 2567
rect 5793 2553 5807 2567
rect 5833 2553 5847 2567
rect 5913 2553 5927 2567
rect 5953 2553 5967 2567
rect 5993 2553 6007 2567
rect 6093 2553 6107 2567
rect 6173 2553 6187 2567
rect 6213 2553 6227 2567
rect 6333 2553 6347 2567
rect 6373 2553 6387 2567
rect 6413 2553 6427 2567
rect 6573 2553 6587 2567
rect 6613 2553 6627 2567
rect 6653 2553 6667 2567
rect 613 2533 627 2547
rect 653 2533 667 2547
rect 693 2533 707 2547
rect 793 2533 807 2547
rect 853 2533 867 2547
rect 993 2533 1007 2547
rect 1313 2533 1327 2547
rect 1453 2533 1467 2547
rect 1513 2533 1527 2547
rect 1553 2533 1567 2547
rect 1853 2533 1867 2547
rect 1913 2533 1927 2547
rect 1973 2533 1987 2547
rect 2013 2533 2027 2547
rect 2153 2533 2167 2547
rect 2213 2533 2227 2547
rect 2273 2533 2287 2547
rect 2333 2533 2347 2547
rect 2633 2533 2647 2547
rect 2693 2533 2707 2547
rect 2873 2533 2887 2547
rect 2933 2533 2947 2547
rect 2993 2533 3007 2547
rect 3033 2533 3047 2547
rect 3093 2533 3107 2547
rect 3493 2533 3507 2547
rect 3553 2533 3567 2547
rect 3593 2533 3607 2547
rect 3633 2533 3647 2547
rect 3693 2533 3707 2547
rect 3733 2533 3747 2547
rect 3833 2533 3847 2547
rect 3873 2533 3887 2547
rect 3913 2533 3927 2547
rect 3953 2533 3967 2547
rect 3993 2533 4007 2547
rect 4033 2533 4047 2547
rect 4213 2533 4227 2547
rect 4253 2533 4267 2547
rect 4553 2533 4567 2547
rect 4633 2533 4647 2547
rect 4673 2533 4687 2547
rect 4713 2533 4727 2547
rect 4773 2533 4787 2547
rect 5093 2533 5107 2547
rect 5153 2533 5167 2547
rect 5193 2533 5207 2547
rect 5273 2533 5287 2547
rect 5313 2533 5327 2547
rect 5533 2533 5547 2547
rect 5673 2533 5687 2547
rect 5813 2533 5827 2547
rect 5853 2533 5867 2547
rect 5933 2533 5947 2547
rect 5973 2533 5987 2547
rect 6033 2533 6047 2547
rect 6353 2533 6367 2547
rect 6393 2533 6407 2547
rect 6433 2533 6447 2547
rect 6473 2533 6487 2547
rect 6533 2533 6547 2547
rect 6593 2533 6607 2547
rect 6633 2533 6647 2547
rect 673 2513 687 2527
rect 713 2513 727 2527
rect 773 2513 787 2527
rect 813 2513 827 2527
rect 1293 2513 1307 2527
rect 1333 2513 1347 2527
rect 3473 2513 3487 2527
rect 3513 2513 3527 2527
rect 3613 2513 3627 2527
rect 3653 2513 3667 2527
rect 3713 2513 3727 2527
rect 3753 2513 3767 2527
rect 3813 2513 3827 2527
rect 3853 2513 3867 2527
rect 673 2293 687 2307
rect 753 2293 767 2307
rect 793 2293 807 2307
rect 833 2293 847 2307
rect 873 2293 887 2307
rect 2513 2293 2527 2307
rect 2553 2293 2567 2307
rect 3793 2293 3807 2307
rect 3833 2293 3847 2307
rect 3893 2293 3907 2307
rect 3933 2293 3947 2307
rect 5713 2293 5727 2307
rect 5753 2293 5767 2307
rect 5813 2293 5827 2307
rect 5853 2293 5867 2307
rect 6473 2293 6487 2307
rect 6513 2293 6527 2307
rect 373 2273 387 2287
rect 413 2273 427 2287
rect 553 2273 567 2287
rect 593 2273 607 2287
rect 733 2273 747 2287
rect 773 2273 787 2287
rect 853 2273 867 2287
rect 1173 2273 1187 2287
rect 1473 2273 1487 2287
rect 1533 2273 1547 2287
rect 1573 2273 1587 2287
rect 1653 2273 1667 2287
rect 1693 2273 1707 2287
rect 1933 2273 1947 2287
rect 1973 2273 1987 2287
rect 2033 2273 2047 2287
rect 2413 2273 2427 2287
rect 2453 2273 2467 2287
rect 2533 2273 2547 2287
rect 2573 2273 2587 2287
rect 2633 2273 2647 2287
rect 2673 2273 2687 2287
rect 2713 2273 2727 2287
rect 2753 2273 2767 2287
rect 3133 2273 3147 2287
rect 3173 2273 3187 2287
rect 3253 2273 3267 2287
rect 3293 2273 3307 2287
rect 3433 2273 3447 2287
rect 3813 2273 3827 2287
rect 3873 2273 3887 2287
rect 3913 2273 3927 2287
rect 3973 2273 3987 2287
rect 4033 2273 4047 2287
rect 4093 2273 4107 2287
rect 4153 2273 4167 2287
rect 4213 2273 4227 2287
rect 4273 2273 4287 2287
rect 4493 2273 4507 2287
rect 4553 2273 4567 2287
rect 4653 2273 4667 2287
rect 4713 2273 4727 2287
rect 4733 2273 4747 2287
rect 4793 2273 4807 2287
rect 4933 2273 4947 2287
rect 4993 2273 5007 2287
rect 5093 2273 5107 2287
rect 5133 2273 5147 2287
rect 5173 2273 5187 2287
rect 5233 2273 5247 2287
rect 5273 2273 5287 2287
rect 5373 2273 5387 2287
rect 5433 2273 5447 2287
rect 5453 2273 5467 2287
rect 5513 2273 5527 2287
rect 5573 2273 5587 2287
rect 5633 2273 5647 2287
rect 5733 2273 5747 2287
rect 5773 2273 5787 2287
rect 5833 2273 5847 2287
rect 5873 2273 5887 2287
rect 5913 2273 5927 2287
rect 5993 2273 6007 2287
rect 6033 2273 6047 2287
rect 6113 2273 6127 2287
rect 6173 2273 6187 2287
rect 6233 2273 6247 2287
rect 6293 2273 6307 2287
rect 6333 2273 6347 2287
rect 6393 2273 6407 2287
rect 6433 2273 6447 2287
rect 6493 2273 6507 2287
rect 6553 2273 6567 2287
rect 6593 2273 6607 2287
rect 6673 2273 6687 2287
rect 93 2253 107 2267
rect 133 2253 147 2267
rect 213 2253 227 2267
rect 273 2253 287 2267
rect 313 2253 327 2267
rect 353 2253 367 2267
rect 473 2253 487 2267
rect 513 2253 527 2267
rect 533 2253 547 2267
rect 573 2253 587 2267
rect 653 2253 667 2267
rect 713 2253 727 2267
rect 933 2253 947 2267
rect 1013 2253 1027 2267
rect 1053 2253 1067 2267
rect 1293 2253 1307 2267
rect 1333 2253 1347 2267
rect 1413 2253 1427 2267
rect 1513 2253 1527 2267
rect 1553 2253 1567 2267
rect 1593 2253 1607 2267
rect 1633 2253 1647 2267
rect 1673 2253 1687 2267
rect 1753 2253 1767 2267
rect 1793 2253 1807 2267
rect 1833 2253 1847 2267
rect 1873 2253 1887 2267
rect 1913 2253 1927 2267
rect 1953 2253 1967 2267
rect 1993 2253 2007 2267
rect 2153 2253 2167 2267
rect 2193 2253 2207 2267
rect 2273 2253 2287 2267
rect 2333 2253 2347 2267
rect 2373 2253 2387 2267
rect 2393 2253 2407 2267
rect 2433 2253 2447 2267
rect 2613 2253 2627 2267
rect 2693 2253 2707 2267
rect 2733 2253 2747 2267
rect 2813 2253 2827 2267
rect 2853 2253 2867 2267
rect 2893 2253 2907 2267
rect 2973 2253 2987 2267
rect 3013 2253 3027 2267
rect 3113 2253 3127 2267
rect 3153 2253 3167 2267
rect 3233 2253 3247 2267
rect 3273 2253 3287 2267
rect 3313 2253 3327 2267
rect 3353 2253 3367 2267
rect 3393 2253 3407 2267
rect 3493 2253 3507 2267
rect 3533 2253 3547 2267
rect 3633 2253 3647 2267
rect 3673 2253 3687 2267
rect 3753 2253 3767 2267
rect 3993 2253 4007 2267
rect 4053 2253 4067 2267
rect 4113 2253 4127 2267
rect 4173 2253 4187 2267
rect 4233 2253 4247 2267
rect 4293 2253 4307 2267
rect 4333 2253 4347 2267
rect 4373 2253 4387 2267
rect 4433 2253 4447 2267
rect 4473 2253 4487 2267
rect 4513 2253 4527 2267
rect 4573 2253 4587 2267
rect 4633 2253 4647 2267
rect 4693 2253 4707 2267
rect 4753 2253 4767 2267
rect 4813 2253 4827 2267
rect 4853 2253 4867 2267
rect 4893 2253 4907 2267
rect 4953 2253 4967 2267
rect 5013 2253 5027 2267
rect 5073 2253 5087 2267
rect 5213 2253 5227 2267
rect 5253 2253 5267 2267
rect 5293 2253 5307 2267
rect 5353 2253 5367 2267
rect 5413 2253 5427 2267
rect 5473 2253 5487 2267
rect 5533 2253 5547 2267
rect 5593 2253 5607 2267
rect 5653 2253 5667 2267
rect 5973 2253 5987 2267
rect 6013 2253 6027 2267
rect 6053 2253 6067 2267
rect 6093 2253 6107 2267
rect 6153 2253 6167 2267
rect 6213 2253 6227 2267
rect 6273 2253 6287 2267
rect 6373 2253 6387 2267
rect 6413 2253 6427 2267
rect 6613 2253 6627 2267
rect 433 2233 447 2247
rect 493 2233 507 2247
rect 1153 2233 1167 2247
rect 1493 2233 1507 2247
rect 1773 2233 1787 2247
rect 1853 2233 1867 2247
rect 2053 2233 2067 2247
rect 2353 2233 2367 2247
rect 2653 2233 2667 2247
rect 2833 2233 2847 2247
rect 3373 2233 3387 2247
rect 3453 2233 3467 2247
rect 3513 2233 3527 2247
rect 4453 2233 4467 2247
rect 4873 2233 4887 2247
rect 5113 2233 5127 2247
rect 5153 2233 5167 2247
rect 5933 2233 5947 2247
rect 6313 2233 6327 2247
rect 6573 2233 6587 2247
rect 6653 2233 6667 2247
rect 53 2093 67 2107
rect 593 2093 607 2107
rect 853 2093 867 2107
rect 1353 2093 1367 2107
rect 1773 2093 1787 2107
rect 2513 2093 2527 2107
rect 2913 2093 2927 2107
rect 3153 2093 3167 2107
rect 3193 2093 3207 2107
rect 3393 2093 3407 2107
rect 3733 2093 3747 2107
rect 3933 2093 3947 2107
rect 4173 2093 4187 2107
rect 4453 2093 4467 2107
rect 4653 2093 4667 2107
rect 4853 2093 4867 2107
rect 5133 2093 5147 2107
rect 5173 2093 5187 2107
rect 5553 2093 5567 2107
rect 5753 2093 5767 2107
rect 6473 2093 6487 2107
rect 33 2073 47 2087
rect 73 2073 87 2087
rect 573 2073 587 2087
rect 613 2073 627 2087
rect 633 2073 647 2087
rect 673 2073 687 2087
rect 833 2073 847 2087
rect 873 2073 887 2087
rect 1013 2073 1027 2087
rect 1073 2073 1087 2087
rect 1193 2073 1207 2087
rect 1233 2073 1247 2087
rect 1313 2073 1327 2087
rect 1413 2073 1427 2087
rect 1453 2073 1467 2087
rect 1493 2073 1507 2087
rect 1573 2073 1587 2087
rect 1613 2073 1627 2087
rect 1673 2073 1687 2087
rect 1713 2073 1727 2087
rect 1753 2073 1767 2087
rect 1793 2073 1807 2087
rect 1853 2073 1867 2087
rect 1893 2073 1907 2087
rect 1933 2073 1947 2087
rect 1993 2073 2007 2087
rect 2053 2073 2067 2087
rect 2113 2073 2127 2087
rect 2233 2073 2247 2087
rect 2273 2073 2287 2087
rect 2353 2073 2367 2087
rect 2433 2073 2447 2087
rect 2473 2073 2487 2087
rect 2493 2073 2507 2087
rect 2533 2073 2547 2087
rect 2693 2073 2707 2087
rect 2753 2073 2767 2087
rect 2813 2073 2827 2087
rect 2873 2073 2887 2087
rect 2973 2073 2987 2087
rect 3013 2073 3027 2087
rect 3053 2073 3067 2087
rect 3113 2073 3127 2087
rect 3253 2073 3267 2087
rect 3293 2073 3307 2087
rect 3333 2073 3347 2087
rect 3373 2073 3387 2087
rect 3413 2073 3427 2087
rect 3533 2073 3547 2087
rect 3573 2073 3587 2087
rect 3653 2073 3667 2087
rect 3713 2073 3727 2087
rect 3753 2073 3767 2087
rect 3793 2073 3807 2087
rect 3833 2073 3847 2087
rect 3873 2073 3887 2087
rect 3953 2073 3967 2087
rect 3993 2073 4007 2087
rect 4153 2073 4167 2087
rect 4193 2073 4207 2087
rect 4293 2073 4307 2087
rect 4333 2073 4347 2087
rect 4413 2073 4427 2087
rect 4513 2073 4527 2087
rect 4553 2073 4567 2087
rect 4593 2073 4607 2087
rect 4633 2073 4647 2087
rect 4673 2073 4687 2087
rect 4753 2073 4767 2087
rect 4793 2073 4807 2087
rect 4833 2073 4847 2087
rect 4873 2073 4887 2087
rect 4893 2073 4907 2087
rect 4933 2073 4947 2087
rect 4973 2073 4987 2087
rect 5113 2073 5127 2087
rect 5153 2073 5167 2087
rect 5193 2073 5207 2087
rect 5293 2073 5307 2087
rect 5333 2073 5347 2087
rect 5373 2073 5387 2087
rect 5393 2073 5407 2087
rect 5433 2073 5447 2087
rect 5473 2073 5487 2087
rect 5533 2073 5547 2087
rect 5573 2073 5587 2087
rect 5613 2073 5627 2087
rect 5653 2073 5667 2087
rect 5693 2073 5707 2087
rect 5873 2073 5887 2087
rect 5953 2073 5967 2087
rect 5993 2073 6007 2087
rect 6173 2073 6187 2087
rect 6213 2073 6227 2087
rect 6293 2073 6307 2087
rect 6353 2073 6367 2087
rect 6413 2073 6427 2087
rect 6513 2073 6527 2087
rect 6553 2073 6567 2087
rect 6593 2073 6607 2087
rect 133 2053 147 2067
rect 213 2053 227 2067
rect 253 2053 267 2067
rect 313 2053 327 2067
rect 353 2053 367 2067
rect 413 2053 427 2067
rect 453 2053 467 2067
rect 493 2053 507 2067
rect 653 2053 667 2067
rect 693 2053 707 2067
rect 733 2053 747 2067
rect 773 2053 787 2067
rect 953 2053 967 2067
rect 993 2053 1007 2067
rect 1053 2053 1067 2067
rect 1373 2053 1387 2067
rect 1433 2053 1447 2067
rect 1473 2053 1487 2067
rect 1553 2053 1567 2067
rect 1593 2053 1607 2067
rect 1653 2053 1667 2067
rect 1693 2053 1707 2067
rect 1833 2053 1847 2067
rect 1873 2053 1887 2067
rect 1953 2053 1967 2067
rect 2013 2053 2027 2067
rect 2073 2053 2087 2067
rect 2133 2053 2147 2067
rect 2413 2053 2427 2067
rect 2453 2053 2467 2067
rect 2613 2053 2627 2067
rect 2653 2053 2667 2067
rect 2673 2053 2687 2067
rect 2733 2053 2747 2067
rect 2833 2053 2847 2067
rect 2893 2053 2907 2067
rect 2933 2053 2947 2067
rect 2993 2053 3007 2067
rect 3033 2053 3047 2067
rect 3133 2053 3147 2067
rect 3173 2053 3187 2067
rect 3213 2053 3227 2067
rect 3273 2053 3287 2067
rect 3313 2053 3327 2067
rect 3813 2053 3827 2067
rect 3853 2053 3867 2067
rect 3913 2053 3927 2067
rect 3973 2053 3987 2067
rect 4013 2053 4027 2067
rect 4073 2053 4087 2067
rect 4473 2053 4487 2067
rect 4533 2053 4547 2067
rect 4573 2053 4587 2067
rect 4733 2053 4747 2067
rect 4773 2053 4787 2067
rect 4913 2053 4927 2067
rect 4953 2053 4967 2067
rect 5053 2053 5067 2067
rect 5233 2053 5247 2067
rect 5313 2053 5327 2067
rect 5353 2053 5367 2067
rect 5413 2053 5427 2067
rect 5453 2053 5467 2067
rect 5633 2053 5647 2067
rect 5673 2053 5687 2067
rect 5733 2053 5747 2067
rect 5793 2053 5807 2067
rect 6333 2053 6347 2067
rect 6393 2053 6407 2067
rect 6453 2053 6467 2067
rect 6493 2053 6507 2067
rect 6573 2053 6587 2067
rect 6613 2053 6627 2067
rect 113 2033 127 2047
rect 153 2033 167 2047
rect 193 2033 207 2047
rect 233 2033 247 2047
rect 293 2033 307 2047
rect 333 2033 347 2047
rect 393 2033 407 2047
rect 433 2033 447 2047
rect 473 2033 487 2047
rect 513 2033 527 2047
rect 753 2033 767 2047
rect 793 2033 807 2047
rect 933 2033 947 2047
rect 973 2033 987 2047
rect 2593 2033 2607 2047
rect 2633 2033 2647 2047
rect 4053 2033 4067 2047
rect 4093 2033 4107 2047
rect 5033 2033 5047 2047
rect 5073 2033 5087 2047
rect 5773 2033 5787 2047
rect 5813 2033 5827 2047
rect 893 1813 907 1827
rect 933 1813 947 1827
rect 1013 1813 1027 1827
rect 1253 1813 1267 1827
rect 1293 1813 1307 1827
rect 1333 1813 1347 1827
rect 1373 1813 1387 1827
rect 2833 1813 2847 1827
rect 2873 1813 2887 1827
rect 3393 1813 3407 1827
rect 3433 1813 3447 1827
rect 3533 1813 3547 1827
rect 3573 1813 3587 1827
rect 3733 1813 3747 1827
rect 3773 1813 3787 1827
rect 3853 1813 3867 1827
rect 3893 1813 3907 1827
rect 5293 1813 5307 1827
rect 5333 1813 5347 1827
rect 5673 1813 5687 1827
rect 5713 1813 5727 1827
rect 6593 1813 6607 1827
rect 6633 1813 6647 1827
rect 33 1793 47 1807
rect 493 1793 507 1807
rect 553 1793 567 1807
rect 593 1793 607 1807
rect 913 1793 927 1807
rect 953 1793 967 1807
rect 1093 1793 1107 1807
rect 1153 1793 1167 1807
rect 1193 1793 1207 1807
rect 1273 1793 1287 1807
rect 1353 1793 1367 1807
rect 1393 1793 1407 1807
rect 1433 1793 1447 1807
rect 1733 1793 1747 1807
rect 1793 1793 1807 1807
rect 1833 1793 1847 1807
rect 1993 1793 2007 1807
rect 2033 1793 2047 1807
rect 2353 1793 2367 1807
rect 2393 1793 2407 1807
rect 2453 1793 2467 1807
rect 2813 1793 2827 1807
rect 2853 1793 2867 1807
rect 2933 1793 2947 1807
rect 2973 1793 2987 1807
rect 3133 1793 3147 1807
rect 3173 1793 3187 1807
rect 3233 1793 3247 1807
rect 3273 1793 3287 1807
rect 3413 1793 3427 1807
rect 3553 1793 3567 1807
rect 3633 1793 3647 1807
rect 3673 1793 3687 1807
rect 3753 1793 3767 1807
rect 3813 1793 3827 1807
rect 3873 1793 3887 1807
rect 4033 1793 4047 1807
rect 4073 1793 4087 1807
rect 4233 1793 4247 1807
rect 4273 1793 4287 1807
rect 4313 1793 4327 1807
rect 4353 1793 4367 1807
rect 4413 1793 4427 1807
rect 4453 1793 4467 1807
rect 4613 1793 4627 1807
rect 4653 1793 4667 1807
rect 4713 1793 4727 1807
rect 4993 1793 5007 1807
rect 5033 1793 5047 1807
rect 5193 1793 5207 1807
rect 5233 1793 5247 1807
rect 5273 1793 5287 1807
rect 5313 1793 5327 1807
rect 5473 1793 5487 1807
rect 5553 1793 5567 1807
rect 5593 1793 5607 1807
rect 5633 1793 5647 1807
rect 5693 1793 5707 1807
rect 5793 1793 5807 1807
rect 5833 1793 5847 1807
rect 5973 1793 5987 1807
rect 6013 1793 6027 1807
rect 6093 1793 6107 1807
rect 6133 1793 6147 1807
rect 6173 1793 6187 1807
rect 6233 1793 6247 1807
rect 6293 1793 6307 1807
rect 6353 1793 6367 1807
rect 6433 1793 6447 1807
rect 6493 1793 6507 1807
rect 6533 1793 6547 1807
rect 6613 1793 6627 1807
rect 93 1773 107 1787
rect 173 1773 187 1787
rect 213 1773 227 1787
rect 313 1773 327 1787
rect 353 1773 367 1787
rect 413 1773 427 1787
rect 453 1773 467 1787
rect 573 1773 587 1787
rect 613 1773 627 1787
rect 653 1773 667 1787
rect 733 1773 747 1787
rect 773 1773 787 1787
rect 973 1773 987 1787
rect 1033 1773 1047 1787
rect 1133 1773 1147 1787
rect 1173 1773 1187 1787
rect 1553 1773 1567 1787
rect 1593 1773 1607 1787
rect 1673 1773 1687 1787
rect 1773 1773 1787 1787
rect 1813 1773 1827 1787
rect 1853 1773 1867 1787
rect 1893 1773 1907 1787
rect 1933 1773 1947 1787
rect 1973 1773 1987 1787
rect 2013 1773 2027 1787
rect 2093 1773 2107 1787
rect 2173 1773 2187 1787
rect 2213 1773 2227 1787
rect 2333 1773 2347 1787
rect 2373 1773 2387 1787
rect 2413 1773 2427 1787
rect 2493 1773 2507 1787
rect 2533 1773 2547 1787
rect 2593 1773 2607 1787
rect 2673 1773 2687 1787
rect 2713 1773 2727 1787
rect 2953 1773 2967 1787
rect 2993 1773 3007 1787
rect 3013 1773 3027 1787
rect 3053 1773 3067 1787
rect 3113 1773 3127 1787
rect 3213 1773 3227 1787
rect 3313 1773 3327 1787
rect 3353 1773 3367 1787
rect 3453 1773 3467 1787
rect 3493 1773 3507 1787
rect 3613 1773 3627 1787
rect 3653 1773 3667 1787
rect 3933 1773 3947 1787
rect 3973 1773 3987 1787
rect 4013 1773 4027 1787
rect 4053 1773 4067 1787
rect 4093 1773 4107 1787
rect 4153 1773 4167 1787
rect 4193 1773 4207 1787
rect 4213 1773 4227 1787
rect 4253 1773 4267 1787
rect 4393 1773 4407 1787
rect 4433 1773 4447 1787
rect 4513 1773 4527 1787
rect 4553 1773 4567 1787
rect 4593 1773 4607 1787
rect 4633 1773 4647 1787
rect 4673 1773 4687 1787
rect 4773 1773 4787 1787
rect 4853 1773 4867 1787
rect 4893 1773 4907 1787
rect 5053 1773 5067 1787
rect 5093 1773 5107 1787
rect 5133 1773 5147 1787
rect 5173 1773 5187 1787
rect 5213 1773 5227 1787
rect 5373 1773 5387 1787
rect 5413 1773 5427 1787
rect 5533 1773 5547 1787
rect 5613 1773 5627 1787
rect 5653 1773 5667 1787
rect 5773 1773 5787 1787
rect 5813 1773 5827 1787
rect 5853 1773 5867 1787
rect 5873 1773 5887 1787
rect 5913 1773 5927 1787
rect 5993 1773 6007 1787
rect 6033 1773 6047 1787
rect 6073 1773 6087 1787
rect 6113 1773 6127 1787
rect 6153 1773 6167 1787
rect 6193 1773 6207 1787
rect 6253 1773 6267 1787
rect 6313 1773 6327 1787
rect 6373 1773 6387 1787
rect 6473 1773 6487 1787
rect 6513 1773 6527 1787
rect 53 1753 67 1767
rect 333 1753 347 1767
rect 433 1753 447 1767
rect 513 1753 527 1767
rect 1073 1753 1087 1767
rect 1413 1753 1427 1767
rect 1713 1753 1727 1767
rect 1913 1753 1927 1767
rect 2433 1753 2447 1767
rect 2513 1753 2527 1767
rect 3033 1753 3047 1767
rect 3153 1753 3167 1767
rect 3253 1753 3267 1767
rect 3473 1753 3487 1767
rect 3833 1753 3847 1767
rect 3953 1753 3967 1767
rect 4173 1753 4187 1767
rect 4533 1753 4547 1767
rect 4733 1753 4747 1767
rect 5013 1753 5027 1767
rect 5113 1753 5127 1767
rect 5493 1753 5507 1767
rect 6413 1753 6427 1767
rect 53 1613 67 1627
rect 573 1613 587 1627
rect 713 1613 727 1627
rect 1073 1613 1087 1627
rect 1353 1613 1367 1627
rect 2113 1613 2127 1627
rect 2313 1613 2327 1627
rect 2573 1613 2587 1627
rect 3753 1613 3767 1627
rect 3813 1613 3827 1627
rect 4013 1613 4027 1627
rect 5853 1613 5867 1627
rect 6113 1613 6127 1627
rect 6393 1613 6407 1627
rect 33 1593 47 1607
rect 73 1593 87 1607
rect 373 1593 387 1607
rect 413 1593 427 1607
rect 493 1593 507 1607
rect 753 1593 767 1607
rect 873 1593 887 1607
rect 913 1593 927 1607
rect 993 1593 1007 1607
rect 1093 1593 1107 1607
rect 1133 1593 1147 1607
rect 1173 1593 1187 1607
rect 1253 1593 1267 1607
rect 1293 1593 1307 1607
rect 1333 1593 1347 1607
rect 1373 1593 1387 1607
rect 1413 1593 1427 1607
rect 1473 1593 1487 1607
rect 1533 1593 1547 1607
rect 1593 1593 1607 1607
rect 1653 1593 1667 1607
rect 1713 1593 1727 1607
rect 1773 1593 1787 1607
rect 1853 1593 1867 1607
rect 1893 1593 1907 1607
rect 2013 1593 2027 1607
rect 2073 1593 2087 1607
rect 2173 1593 2187 1607
rect 2213 1593 2227 1607
rect 2253 1593 2267 1607
rect 2293 1593 2307 1607
rect 2333 1593 2347 1607
rect 2413 1593 2427 1607
rect 2453 1593 2467 1607
rect 2493 1593 2507 1607
rect 2533 1593 2547 1607
rect 2553 1593 2567 1607
rect 2593 1593 2607 1607
rect 2813 1593 2827 1607
rect 2873 1593 2887 1607
rect 3033 1593 3047 1607
rect 3153 1593 3167 1607
rect 3193 1593 3207 1607
rect 3273 1593 3287 1607
rect 3433 1593 3447 1607
rect 3473 1593 3487 1607
rect 3493 1593 3507 1607
rect 3533 1593 3547 1607
rect 3573 1593 3587 1607
rect 3653 1593 3667 1607
rect 3693 1593 3707 1607
rect 3793 1593 3807 1607
rect 3833 1593 3847 1607
rect 3873 1593 3887 1607
rect 3913 1593 3927 1607
rect 3953 1593 3967 1607
rect 4113 1593 4127 1607
rect 4153 1593 4167 1607
rect 4233 1593 4247 1607
rect 4293 1593 4307 1607
rect 4353 1593 4367 1607
rect 4413 1593 4427 1607
rect 4473 1593 4487 1607
rect 4533 1593 4547 1607
rect 4593 1593 4607 1607
rect 4653 1593 4667 1607
rect 4713 1593 4727 1607
rect 4773 1593 4787 1607
rect 4833 1593 4847 1607
rect 4893 1593 4907 1607
rect 4953 1593 4967 1607
rect 5013 1593 5027 1607
rect 5093 1593 5107 1607
rect 5133 1593 5147 1607
rect 5253 1593 5267 1607
rect 5333 1593 5347 1607
rect 5373 1593 5387 1607
rect 5473 1593 5487 1607
rect 5513 1593 5527 1607
rect 5553 1593 5567 1607
rect 5613 1593 5627 1607
rect 5673 1593 5687 1607
rect 5753 1593 5767 1607
rect 5793 1593 5807 1607
rect 5833 1593 5847 1607
rect 5873 1593 5887 1607
rect 6013 1593 6027 1607
rect 6053 1593 6067 1607
rect 6093 1593 6107 1607
rect 6133 1593 6147 1607
rect 6173 1593 6187 1607
rect 6213 1593 6227 1607
rect 6253 1593 6267 1607
rect 6293 1593 6307 1607
rect 6353 1593 6367 1607
rect 6473 1593 6487 1607
rect 6553 1593 6567 1607
rect 6593 1593 6607 1607
rect 113 1573 127 1587
rect 253 1573 267 1587
rect 553 1573 567 1587
rect 593 1573 607 1587
rect 633 1573 647 1587
rect 693 1573 707 1587
rect 733 1573 747 1587
rect 1053 1573 1067 1587
rect 1113 1573 1127 1587
rect 1153 1573 1167 1587
rect 1233 1573 1247 1587
rect 1273 1573 1287 1587
rect 1433 1573 1447 1587
rect 1493 1573 1507 1587
rect 1553 1573 1567 1587
rect 1613 1573 1627 1587
rect 1673 1573 1687 1587
rect 1733 1573 1747 1587
rect 1993 1573 2007 1587
rect 2053 1573 2067 1587
rect 2133 1573 2147 1587
rect 2193 1573 2207 1587
rect 2233 1573 2247 1587
rect 2393 1573 2407 1587
rect 2433 1573 2447 1587
rect 2673 1573 2687 1587
rect 2733 1573 2747 1587
rect 2833 1573 2847 1587
rect 2893 1573 2907 1587
rect 2953 1573 2967 1587
rect 2993 1573 3007 1587
rect 3053 1573 3067 1587
rect 3353 1573 3367 1587
rect 3413 1573 3427 1587
rect 3453 1573 3467 1587
rect 3513 1573 3527 1587
rect 3553 1573 3567 1587
rect 3633 1573 3647 1587
rect 3673 1573 3687 1587
rect 3733 1573 3747 1587
rect 3893 1573 3907 1587
rect 3933 1573 3947 1587
rect 3993 1573 4007 1587
rect 4313 1573 4327 1587
rect 4373 1573 4387 1587
rect 4433 1573 4447 1587
rect 4493 1573 4507 1587
rect 4513 1573 4527 1587
rect 4573 1573 4587 1587
rect 4633 1573 4647 1587
rect 4693 1573 4707 1587
rect 4753 1573 4767 1587
rect 4813 1573 4827 1587
rect 4873 1573 4887 1587
rect 4933 1573 4947 1587
rect 5493 1573 5507 1587
rect 5533 1573 5547 1587
rect 5593 1573 5607 1587
rect 5653 1573 5667 1587
rect 5733 1573 5747 1587
rect 5773 1573 5787 1587
rect 5933 1573 5947 1587
rect 5993 1573 6007 1587
rect 6033 1573 6047 1587
rect 6193 1573 6207 1587
rect 6233 1573 6247 1587
rect 6313 1573 6327 1587
rect 6373 1573 6387 1587
rect 6413 1573 6427 1587
rect 613 1553 627 1567
rect 653 1553 667 1567
rect 2653 1553 2667 1567
rect 2693 1553 2707 1567
rect 2713 1553 2727 1567
rect 2753 1553 2767 1567
rect 2933 1553 2947 1567
rect 2973 1553 2987 1567
rect 3333 1553 3347 1567
rect 3373 1553 3387 1567
rect 5913 1553 5927 1567
rect 5953 1553 5967 1567
rect 53 1333 67 1347
rect 513 1333 527 1347
rect 553 1333 567 1347
rect 933 1333 947 1347
rect 973 1333 987 1347
rect 1013 1333 1027 1347
rect 1053 1333 1067 1347
rect 2193 1333 2207 1347
rect 2233 1333 2247 1347
rect 4853 1333 4867 1347
rect 4893 1333 4907 1347
rect 4933 1333 4947 1347
rect 4973 1333 4987 1347
rect 5313 1333 5327 1347
rect 5353 1333 5367 1347
rect 5793 1333 5807 1347
rect 5833 1333 5847 1347
rect 213 1313 227 1327
rect 253 1313 267 1327
rect 393 1313 407 1327
rect 453 1313 467 1327
rect 533 1313 547 1327
rect 573 1313 587 1327
rect 613 1313 627 1327
rect 953 1313 967 1327
rect 993 1313 1007 1327
rect 1033 1313 1047 1327
rect 1433 1313 1447 1327
rect 1573 1313 1587 1327
rect 1653 1313 1667 1327
rect 1713 1313 1727 1327
rect 1853 1313 1867 1327
rect 1893 1313 1907 1327
rect 1953 1313 1967 1327
rect 1993 1313 2007 1327
rect 2053 1313 2067 1327
rect 2113 1313 2127 1327
rect 2153 1313 2167 1327
rect 2213 1313 2227 1327
rect 2273 1313 2287 1327
rect 2333 1313 2347 1327
rect 2433 1313 2447 1327
rect 2493 1313 2507 1327
rect 2553 1313 2567 1327
rect 2593 1313 2607 1327
rect 2653 1313 2667 1327
rect 2693 1313 2707 1327
rect 2793 1313 2807 1327
rect 2833 1313 2847 1327
rect 2993 1313 3007 1327
rect 3033 1313 3047 1327
rect 3093 1313 3107 1327
rect 3173 1313 3187 1327
rect 3233 1313 3247 1327
rect 3613 1313 3627 1327
rect 3653 1313 3667 1327
rect 3713 1313 3727 1327
rect 3753 1313 3767 1327
rect 3813 1313 3827 1327
rect 4353 1313 4367 1327
rect 4413 1313 4427 1327
rect 4453 1313 4467 1327
rect 4513 1313 4527 1327
rect 4573 1313 4587 1327
rect 4673 1313 4687 1327
rect 4713 1313 4727 1327
rect 4873 1313 4887 1327
rect 4953 1313 4967 1327
rect 5033 1313 5047 1327
rect 5073 1313 5087 1327
rect 5153 1313 5167 1327
rect 5193 1313 5207 1327
rect 5233 1313 5247 1327
rect 5333 1313 5347 1327
rect 5393 1313 5407 1327
rect 5433 1313 5447 1327
rect 5533 1313 5547 1327
rect 5573 1313 5587 1327
rect 5593 1313 5607 1327
rect 5653 1313 5667 1327
rect 5713 1313 5727 1327
rect 5813 1313 5827 1327
rect 5873 1313 5887 1327
rect 5913 1313 5927 1327
rect 5973 1313 5987 1327
rect 6033 1313 6047 1327
rect 6073 1313 6087 1327
rect 6133 1313 6147 1327
rect 6173 1313 6187 1327
rect 13 1293 27 1307
rect 73 1293 87 1307
rect 113 1293 127 1307
rect 153 1293 167 1307
rect 233 1293 247 1307
rect 273 1293 287 1307
rect 313 1293 327 1307
rect 353 1293 367 1307
rect 633 1293 647 1307
rect 753 1293 767 1307
rect 793 1293 807 1307
rect 873 1293 887 1307
rect 1093 1293 1107 1307
rect 1133 1293 1147 1307
rect 1253 1293 1267 1307
rect 1293 1293 1307 1307
rect 1373 1293 1387 1307
rect 1633 1293 1647 1307
rect 1693 1293 1707 1307
rect 1753 1293 1767 1307
rect 1793 1293 1807 1307
rect 1833 1293 1847 1307
rect 1873 1293 1887 1307
rect 1913 1293 1927 1307
rect 1973 1293 1987 1307
rect 2013 1293 2027 1307
rect 2093 1293 2107 1307
rect 2133 1293 2147 1307
rect 2293 1293 2307 1307
rect 2353 1293 2367 1307
rect 2413 1293 2427 1307
rect 2473 1293 2487 1307
rect 2533 1293 2547 1307
rect 2573 1293 2587 1307
rect 2613 1293 2627 1307
rect 2633 1293 2647 1307
rect 2673 1293 2687 1307
rect 2713 1293 2727 1307
rect 2773 1293 2787 1307
rect 2813 1293 2827 1307
rect 2853 1293 2867 1307
rect 2873 1293 2887 1307
rect 2913 1293 2927 1307
rect 2973 1293 2987 1307
rect 3013 1293 3027 1307
rect 3053 1293 3067 1307
rect 3153 1293 3167 1307
rect 3213 1293 3227 1307
rect 3333 1293 3347 1307
rect 3373 1293 3387 1307
rect 3453 1293 3467 1307
rect 3513 1293 3527 1307
rect 3553 1293 3567 1307
rect 3593 1293 3607 1307
rect 3633 1293 3647 1307
rect 3673 1293 3687 1307
rect 3733 1293 3747 1307
rect 3773 1293 3787 1307
rect 3873 1293 3887 1307
rect 3953 1293 3967 1307
rect 3993 1293 4007 1307
rect 4113 1293 4127 1307
rect 4193 1293 4207 1307
rect 4233 1293 4247 1307
rect 4393 1293 4407 1307
rect 4433 1293 4447 1307
rect 4473 1293 4487 1307
rect 4533 1293 4547 1307
rect 4593 1293 4607 1307
rect 4653 1293 4667 1307
rect 4693 1293 4707 1307
rect 4733 1293 4747 1307
rect 4773 1293 4787 1307
rect 4813 1293 4827 1307
rect 5013 1293 5027 1307
rect 5053 1293 5067 1307
rect 5093 1293 5107 1307
rect 5133 1293 5147 1307
rect 5173 1293 5187 1307
rect 5213 1293 5227 1307
rect 5253 1293 5267 1307
rect 5373 1293 5387 1307
rect 5413 1293 5427 1307
rect 5453 1293 5467 1307
rect 5513 1293 5527 1307
rect 5613 1293 5627 1307
rect 5673 1293 5687 1307
rect 5733 1293 5747 1307
rect 5893 1293 5907 1307
rect 5933 1293 5947 1307
rect 6013 1293 6027 1307
rect 6053 1293 6067 1307
rect 6113 1293 6127 1307
rect 6153 1293 6167 1307
rect 6193 1293 6207 1307
rect 6253 1293 6267 1307
rect 6333 1293 6347 1307
rect 6373 1293 6387 1307
rect 6493 1293 6507 1307
rect 6573 1293 6587 1307
rect 6613 1293 6627 1307
rect 133 1273 147 1287
rect 333 1273 347 1287
rect 373 1273 387 1287
rect 433 1273 447 1287
rect 593 1273 607 1287
rect 1113 1273 1127 1287
rect 1773 1273 1787 1287
rect 2033 1273 2047 1287
rect 3113 1273 3127 1287
rect 3533 1273 3547 1287
rect 3833 1273 3847 1287
rect 4373 1273 4387 1287
rect 5553 1273 5567 1287
rect 5993 1273 6007 1287
rect 293 1133 307 1147
rect 553 1133 567 1147
rect 733 1133 747 1147
rect 973 1133 987 1147
rect 1753 1133 1767 1147
rect 2153 1133 2167 1147
rect 2593 1133 2607 1147
rect 2793 1133 2807 1147
rect 4093 1133 4107 1147
rect 4293 1133 4307 1147
rect 4513 1133 4527 1147
rect 4953 1133 4967 1147
rect 5133 1133 5147 1147
rect 5193 1133 5207 1147
rect 5273 1133 5287 1147
rect 5433 1133 5447 1147
rect 5513 1133 5527 1147
rect 5593 1133 5607 1147
rect 5673 1133 5687 1147
rect 5813 1133 5827 1147
rect 6193 1133 6207 1147
rect 6253 1133 6267 1147
rect 33 1113 47 1127
rect 113 1113 127 1127
rect 153 1113 167 1127
rect 333 1113 347 1127
rect 413 1113 427 1127
rect 453 1113 467 1127
rect 713 1113 727 1127
rect 753 1113 767 1127
rect 1113 1113 1127 1127
rect 1153 1113 1167 1127
rect 1233 1113 1247 1127
rect 1553 1113 1567 1127
rect 1593 1113 1607 1127
rect 1673 1113 1687 1127
rect 1733 1113 1747 1127
rect 1773 1113 1787 1127
rect 1813 1113 1827 1127
rect 1853 1113 1867 1127
rect 1893 1113 1907 1127
rect 1953 1113 1967 1127
rect 1993 1113 2007 1127
rect 2053 1113 2067 1127
rect 2093 1113 2107 1127
rect 2133 1113 2147 1127
rect 2173 1113 2187 1127
rect 2213 1113 2227 1127
rect 2253 1113 2267 1127
rect 2293 1113 2307 1127
rect 2393 1113 2407 1127
rect 2433 1113 2447 1127
rect 2513 1113 2527 1127
rect 2613 1113 2627 1127
rect 2653 1113 2667 1127
rect 2733 1113 2747 1127
rect 2773 1113 2787 1127
rect 2873 1113 2887 1127
rect 2913 1113 2927 1127
rect 2953 1113 2967 1127
rect 3053 1113 3067 1127
rect 3093 1113 3107 1127
rect 3173 1113 3187 1127
rect 3313 1113 3327 1127
rect 3373 1113 3387 1127
rect 3433 1113 3447 1127
rect 3493 1113 3507 1127
rect 3553 1113 3567 1127
rect 3593 1113 3607 1127
rect 3693 1113 3707 1127
rect 3733 1113 3747 1127
rect 3813 1113 3827 1127
rect 3873 1113 3887 1127
rect 3933 1113 3947 1127
rect 3993 1113 4007 1127
rect 4053 1113 4067 1127
rect 4153 1113 4167 1127
rect 4193 1113 4207 1127
rect 4233 1113 4247 1127
rect 4273 1113 4287 1127
rect 4313 1113 4327 1127
rect 4393 1113 4407 1127
rect 4433 1113 4447 1127
rect 4473 1113 4487 1127
rect 4633 1113 4647 1127
rect 4673 1113 4687 1127
rect 4753 1113 4767 1127
rect 4793 1113 4807 1127
rect 4833 1113 4847 1127
rect 4873 1113 4887 1127
rect 4933 1113 4947 1127
rect 4973 1113 4987 1127
rect 5033 1113 5047 1127
rect 5073 1113 5087 1127
rect 5113 1113 5127 1127
rect 5153 1113 5167 1127
rect 5173 1113 5187 1127
rect 5213 1113 5227 1127
rect 5253 1113 5267 1127
rect 5293 1113 5307 1127
rect 5353 1113 5367 1127
rect 5393 1113 5407 1127
rect 5413 1113 5427 1127
rect 5453 1113 5467 1127
rect 5493 1113 5507 1127
rect 5533 1113 5547 1127
rect 5633 1113 5647 1127
rect 5693 1113 5707 1127
rect 5793 1113 5807 1127
rect 5833 1113 5847 1127
rect 5853 1113 5867 1127
rect 5893 1113 5907 1127
rect 6053 1113 6067 1127
rect 6093 1113 6107 1127
rect 6173 1113 6187 1127
rect 6213 1113 6227 1127
rect 6233 1113 6247 1127
rect 6273 1113 6287 1127
rect 6333 1113 6347 1127
rect 6413 1113 6427 1127
rect 6453 1113 6467 1127
rect 6553 1113 6567 1127
rect 6593 1113 6607 1127
rect 6633 1113 6647 1127
rect 273 1093 287 1107
rect 573 1093 587 1107
rect 613 1093 627 1107
rect 653 1093 667 1107
rect 793 1093 807 1107
rect 833 1093 847 1107
rect 913 1093 927 1107
rect 993 1093 1007 1107
rect 1293 1093 1307 1107
rect 1433 1093 1447 1107
rect 1833 1093 1847 1107
rect 1873 1093 1887 1107
rect 1933 1093 1947 1107
rect 1973 1093 1987 1107
rect 2033 1093 2047 1107
rect 2073 1093 2087 1107
rect 2233 1093 2247 1107
rect 2273 1093 2287 1107
rect 2573 1093 2587 1107
rect 2633 1093 2647 1107
rect 2673 1093 2687 1107
rect 2813 1093 2827 1107
rect 2893 1093 2907 1107
rect 2933 1093 2947 1107
rect 3233 1093 3247 1107
rect 3333 1093 3347 1107
rect 3393 1093 3407 1107
rect 3413 1093 3427 1107
rect 3473 1093 3487 1107
rect 3853 1093 3867 1107
rect 3913 1093 3927 1107
rect 4013 1093 4027 1107
rect 4073 1093 4087 1107
rect 4113 1093 4127 1107
rect 4173 1093 4187 1107
rect 4213 1093 4227 1107
rect 4373 1093 4387 1107
rect 4413 1093 4427 1107
rect 4493 1093 4507 1107
rect 4533 1093 4547 1107
rect 4813 1093 4827 1107
rect 4853 1093 4867 1107
rect 5013 1093 5027 1107
rect 5053 1093 5067 1107
rect 5573 1093 5587 1107
rect 5613 1093 5627 1107
rect 5733 1093 5747 1107
rect 5873 1093 5887 1107
rect 5913 1093 5927 1107
rect 5993 1093 6007 1107
rect 6033 1093 6047 1107
rect 6073 1093 6087 1107
rect 6113 1093 6127 1107
rect 6573 1093 6587 1107
rect 6613 1093 6627 1107
rect 633 1073 647 1087
rect 673 1073 687 1087
rect 813 1073 827 1087
rect 853 1073 867 1087
rect 893 1073 907 1087
rect 933 1073 947 1087
rect 3213 1073 3227 1087
rect 3253 1073 3267 1087
rect 5973 1073 5987 1087
rect 6013 1073 6027 1087
rect 133 853 147 867
rect 173 853 187 867
rect 653 853 667 867
rect 693 853 707 867
rect 753 853 767 867
rect 793 853 807 867
rect 2013 853 2027 867
rect 2053 853 2067 867
rect 3433 853 3447 867
rect 3473 853 3487 867
rect 4393 853 4407 867
rect 4433 853 4447 867
rect 4633 853 4647 867
rect 4673 853 4687 867
rect 4873 853 4887 867
rect 4913 853 4927 867
rect 5653 853 5667 867
rect 5693 853 5707 867
rect 5853 853 5867 867
rect 5893 853 5907 867
rect 6393 853 6407 867
rect 6433 853 6447 867
rect 73 833 87 847
rect 153 833 167 847
rect 453 833 467 847
rect 673 833 687 847
rect 733 833 747 847
rect 773 833 787 847
rect 853 833 867 847
rect 893 833 907 847
rect 973 833 987 847
rect 1013 833 1027 847
rect 1073 833 1087 847
rect 1113 833 1127 847
rect 1193 833 1207 847
rect 1253 833 1267 847
rect 1353 833 1367 847
rect 1393 833 1407 847
rect 1453 833 1467 847
rect 1753 833 1767 847
rect 1793 833 1807 847
rect 1853 833 1867 847
rect 1933 833 1947 847
rect 1973 833 1987 847
rect 2033 833 2047 847
rect 2353 833 2367 847
rect 2413 833 2427 847
rect 2453 833 2467 847
rect 2613 833 2627 847
rect 2653 833 2667 847
rect 2713 833 2727 847
rect 2853 833 2867 847
rect 2893 833 2907 847
rect 2933 833 2947 847
rect 3033 833 3047 847
rect 3073 833 3087 847
rect 3133 833 3147 847
rect 3193 833 3207 847
rect 3253 833 3267 847
rect 3313 833 3327 847
rect 3353 833 3367 847
rect 3393 833 3407 847
rect 3453 833 3467 847
rect 3513 833 3527 847
rect 3573 833 3587 847
rect 3653 833 3667 847
rect 3733 833 3747 847
rect 3793 833 3807 847
rect 4053 833 4067 847
rect 4113 833 4127 847
rect 4173 833 4187 847
rect 4213 833 4227 847
rect 4293 833 4307 847
rect 4333 833 4347 847
rect 4413 833 4427 847
rect 4453 833 4467 847
rect 4493 833 4507 847
rect 4553 833 4567 847
rect 4593 833 4607 847
rect 4653 833 4667 847
rect 4733 833 4747 847
rect 4793 833 4807 847
rect 4833 833 4847 847
rect 4893 833 4907 847
rect 4953 833 4967 847
rect 5013 833 5027 847
rect 5113 833 5127 847
rect 5173 833 5187 847
rect 5213 833 5227 847
rect 5353 833 5367 847
rect 5393 833 5407 847
rect 5433 833 5447 847
rect 5513 833 5527 847
rect 5573 833 5587 847
rect 5613 833 5627 847
rect 5673 833 5687 847
rect 5753 833 5767 847
rect 5793 833 5807 847
rect 5873 833 5887 847
rect 5913 833 5927 847
rect 6193 833 6207 847
rect 6233 833 6247 847
rect 6293 833 6307 847
rect 6333 833 6347 847
rect 6413 833 6427 847
rect 33 813 47 827
rect 213 813 227 827
rect 293 813 307 827
rect 333 813 347 827
rect 513 813 527 827
rect 553 813 567 827
rect 573 813 587 827
rect 613 813 627 827
rect 833 813 847 827
rect 873 813 887 827
rect 913 813 927 827
rect 953 813 967 827
rect 993 813 1007 827
rect 1053 813 1067 827
rect 1093 813 1107 827
rect 1233 813 1247 827
rect 1293 813 1307 827
rect 1333 813 1347 827
rect 1373 813 1387 827
rect 1573 813 1587 827
rect 1613 813 1627 827
rect 1693 813 1707 827
rect 1813 813 1827 827
rect 1873 813 1887 827
rect 1913 813 1927 827
rect 1953 813 1967 827
rect 2113 813 2127 827
rect 2193 813 2207 827
rect 2233 813 2247 827
rect 2393 813 2407 827
rect 2433 813 2447 827
rect 2473 813 2487 827
rect 2513 813 2527 827
rect 2553 813 2567 827
rect 2633 813 2647 827
rect 2673 813 2687 827
rect 2953 813 2967 827
rect 3013 813 3027 827
rect 3113 813 3127 827
rect 3173 813 3187 827
rect 3233 813 3247 827
rect 3293 813 3307 827
rect 3373 813 3387 827
rect 3413 813 3427 827
rect 3533 813 3547 827
rect 3593 813 3607 827
rect 3713 813 3727 827
rect 3773 813 3787 827
rect 3893 813 3907 827
rect 3933 813 3947 827
rect 4013 813 4027 827
rect 4073 813 4087 827
rect 4133 813 4147 827
rect 4233 813 4247 827
rect 4273 813 4287 827
rect 4313 813 4327 827
rect 4533 813 4547 827
rect 4573 813 4587 827
rect 4773 813 4787 827
rect 4813 813 4827 827
rect 4973 813 4987 827
rect 5033 813 5047 827
rect 5093 813 5107 827
rect 5153 813 5167 827
rect 5453 813 5467 827
rect 5553 813 5567 827
rect 5593 813 5607 827
rect 5733 813 5747 827
rect 5773 813 5787 827
rect 6013 813 6027 827
rect 6053 813 6067 827
rect 6133 813 6147 827
rect 6173 813 6187 827
rect 6213 813 6227 827
rect 6273 813 6287 827
rect 6313 813 6327 827
rect 6533 813 6547 827
rect 6573 813 6587 827
rect 6653 813 6667 827
rect 13 793 27 807
rect 473 793 487 807
rect 533 793 547 807
rect 593 793 607 807
rect 1473 793 1487 807
rect 1733 793 1747 807
rect 2333 793 2347 807
rect 2533 793 2547 807
rect 2913 793 2927 807
rect 3053 793 3067 807
rect 3673 793 3687 807
rect 4193 793 4207 807
rect 4473 793 4487 807
rect 4753 793 4767 807
rect 5413 793 5427 807
rect 5533 793 5547 807
rect 13 653 27 667
rect 173 653 187 667
rect 253 653 267 667
rect 373 653 387 667
rect 693 653 707 667
rect 753 653 767 667
rect 853 653 867 667
rect 2833 653 2847 667
rect 2913 653 2927 667
rect 2953 653 2967 667
rect 3293 653 3307 667
rect 3553 653 3567 667
rect 3653 653 3667 667
rect 4193 653 4207 667
rect 4473 653 4487 667
rect 4713 653 4727 667
rect 4973 653 4987 667
rect 5673 653 5687 667
rect 5753 653 5767 667
rect 5833 653 5847 667
rect 5893 653 5907 667
rect 5993 653 6007 667
rect 6553 653 6567 667
rect 6613 653 6627 667
rect 213 633 227 647
rect 333 633 347 647
rect 833 633 847 647
rect 873 633 887 647
rect 973 633 987 647
rect 1033 633 1047 647
rect 1153 633 1167 647
rect 1193 633 1207 647
rect 1273 633 1287 647
rect 1313 633 1327 647
rect 1353 633 1367 647
rect 1553 633 1567 647
rect 1593 633 1607 647
rect 1673 633 1687 647
rect 1793 633 1807 647
rect 1833 633 1847 647
rect 1913 633 1927 647
rect 2033 633 2047 647
rect 2073 633 2087 647
rect 2153 633 2167 647
rect 2273 633 2287 647
rect 2313 633 2327 647
rect 2393 633 2407 647
rect 2453 633 2467 647
rect 2533 633 2547 647
rect 2573 633 2587 647
rect 2693 633 2707 647
rect 2733 633 2747 647
rect 2773 633 2787 647
rect 2873 633 2887 647
rect 3013 633 3027 647
rect 3053 633 3067 647
rect 3353 633 3367 647
rect 3393 633 3407 647
rect 3593 633 3607 647
rect 3633 633 3647 647
rect 3673 633 3687 647
rect 3713 633 3727 647
rect 3753 633 3767 647
rect 3933 633 3947 647
rect 4013 633 4027 647
rect 4053 633 4067 647
rect 4173 633 4187 647
rect 4213 633 4227 647
rect 4253 633 4267 647
rect 4333 633 4347 647
rect 4373 633 4387 647
rect 4533 633 4547 647
rect 4573 633 4587 647
rect 4613 633 4627 647
rect 4673 633 4687 647
rect 4793 633 4807 647
rect 4833 633 4847 647
rect 5013 633 5027 647
rect 5073 633 5087 647
rect 5233 633 5247 647
rect 5313 633 5327 647
rect 5353 633 5367 647
rect 5473 633 5487 647
rect 5533 633 5547 647
rect 5593 633 5607 647
rect 5653 633 5667 647
rect 5693 633 5707 647
rect 5733 633 5747 647
rect 5773 633 5787 647
rect 5813 633 5827 647
rect 5853 633 5867 647
rect 5873 633 5887 647
rect 5913 633 5927 647
rect 5973 633 5987 647
rect 6013 633 6027 647
rect 6033 633 6047 647
rect 6073 633 6087 647
rect 6133 633 6147 647
rect 6173 633 6187 647
rect 6393 633 6407 647
rect 6433 633 6447 647
rect 6513 633 6527 647
rect 33 613 47 627
rect 93 613 107 627
rect 153 613 167 627
rect 193 613 207 627
rect 273 613 287 627
rect 353 613 367 627
rect 393 613 407 627
rect 413 613 427 627
rect 453 613 467 627
rect 553 613 567 627
rect 633 613 647 627
rect 673 613 687 627
rect 713 613 727 627
rect 773 613 787 627
rect 933 613 947 627
rect 993 613 1007 627
rect 1413 613 1427 627
rect 2713 613 2727 627
rect 2753 613 2767 627
rect 2813 613 2827 627
rect 2893 613 2907 627
rect 2933 613 2947 627
rect 2973 613 2987 627
rect 3033 613 3047 627
rect 3073 613 3087 627
rect 3133 613 3147 627
rect 3193 613 3207 627
rect 3233 613 3247 627
rect 3313 613 3327 627
rect 3373 613 3387 627
rect 3413 613 3427 627
rect 3473 613 3487 627
rect 3533 613 3547 627
rect 3573 613 3587 627
rect 3733 613 3747 627
rect 3773 613 3787 627
rect 3853 613 3867 627
rect 3893 613 3907 627
rect 4493 613 4507 627
rect 4553 613 4567 627
rect 4593 613 4607 627
rect 4693 613 4707 627
rect 4733 613 4747 627
rect 4773 613 4787 627
rect 4813 613 4827 627
rect 4873 613 4887 627
rect 4953 613 4967 627
rect 5033 613 5047 627
rect 5093 613 5107 627
rect 5113 613 5127 627
rect 5153 613 5167 627
rect 5453 613 5467 627
rect 5513 613 5527 627
rect 5573 613 5587 627
rect 6053 613 6067 627
rect 6093 613 6107 627
rect 6153 613 6167 627
rect 6193 613 6207 627
rect 6273 613 6287 627
rect 6573 613 6587 627
rect 6633 613 6647 627
rect 73 593 87 607
rect 113 593 127 607
rect 433 593 447 607
rect 473 593 487 607
rect 533 593 547 607
rect 573 593 587 607
rect 613 593 627 607
rect 653 593 667 607
rect 1393 593 1407 607
rect 1433 593 1447 607
rect 3113 593 3127 607
rect 3153 593 3167 607
rect 3213 593 3227 607
rect 3253 593 3267 607
rect 3453 593 3467 607
rect 3493 593 3507 607
rect 3833 593 3847 607
rect 3873 593 3887 607
rect 4853 593 4867 607
rect 4893 593 4907 607
rect 5133 593 5147 607
rect 5173 593 5187 607
rect 6253 593 6267 607
rect 6293 593 6307 607
rect 513 373 527 387
rect 553 373 567 387
rect 753 373 767 387
rect 793 373 807 387
rect 3173 373 3187 387
rect 3213 373 3227 387
rect 4013 373 4027 387
rect 4053 373 4067 387
rect 5573 373 5587 387
rect 5613 373 5627 387
rect 5773 373 5787 387
rect 5813 373 5827 387
rect 493 353 507 367
rect 533 353 547 367
rect 773 353 787 367
rect 853 353 867 367
rect 1393 353 1407 367
rect 1453 353 1467 367
rect 1493 353 1507 367
rect 1553 353 1567 367
rect 1613 353 1627 367
rect 1653 353 1667 367
rect 1953 353 1967 367
rect 2013 353 2027 367
rect 2073 353 2087 367
rect 2113 353 2127 367
rect 2173 353 2187 367
rect 2233 353 2247 367
rect 2273 353 2287 367
rect 2353 353 2367 367
rect 2393 353 2407 367
rect 2773 353 2787 367
rect 2813 353 2827 367
rect 3193 353 3207 367
rect 3273 353 3287 367
rect 3313 353 3327 367
rect 3473 353 3487 367
rect 3513 353 3527 367
rect 3553 353 3567 367
rect 3593 353 3607 367
rect 3713 353 3727 367
rect 3753 353 3767 367
rect 3913 353 3927 367
rect 3953 353 3967 367
rect 4033 353 4047 367
rect 4073 353 4087 367
rect 4513 353 4527 367
rect 4553 353 4567 367
rect 4713 353 4727 367
rect 4753 353 4767 367
rect 4813 353 4827 367
rect 5133 353 5147 367
rect 5173 353 5187 367
rect 5293 353 5307 367
rect 5333 353 5347 367
rect 5453 353 5467 367
rect 5493 353 5507 367
rect 5553 353 5567 367
rect 5593 353 5607 367
rect 5673 353 5687 367
rect 5713 353 5727 367
rect 5793 353 5807 367
rect 5853 353 5867 367
rect 5893 353 5907 367
rect 5953 353 5967 367
rect 5993 353 6007 367
rect 6053 353 6067 367
rect 6093 353 6107 367
rect 6333 353 6347 367
rect 6373 353 6387 367
rect 33 333 47 347
rect 113 333 127 347
rect 153 333 167 347
rect 333 333 347 347
rect 373 333 387 347
rect 453 333 467 347
rect 593 333 607 347
rect 633 333 647 347
rect 693 333 707 347
rect 733 333 747 347
rect 973 333 987 347
rect 1013 333 1027 347
rect 1093 333 1107 347
rect 1153 333 1167 347
rect 1193 333 1207 347
rect 1213 333 1227 347
rect 1253 333 1267 347
rect 1293 333 1307 347
rect 1333 333 1347 347
rect 1433 333 1447 347
rect 1473 333 1487 347
rect 1593 333 1607 347
rect 1633 333 1647 347
rect 1773 333 1787 347
rect 1813 333 1827 347
rect 1893 333 1907 347
rect 2053 333 2067 347
rect 2093 333 2107 347
rect 2213 333 2227 347
rect 2253 333 2267 347
rect 2293 333 2307 347
rect 2373 333 2387 347
rect 2413 333 2427 347
rect 2433 333 2447 347
rect 2473 333 2487 347
rect 2593 333 2607 347
rect 2633 333 2647 347
rect 2713 333 2727 347
rect 2793 333 2807 347
rect 2833 333 2847 347
rect 2853 333 2867 347
rect 2893 333 2907 347
rect 3013 333 3027 347
rect 3053 333 3067 347
rect 3133 333 3147 347
rect 3293 333 3307 347
rect 3333 333 3347 347
rect 3353 333 3367 347
rect 3393 333 3407 347
rect 3453 333 3467 347
rect 3533 333 3547 347
rect 3573 333 3587 347
rect 3633 333 3647 347
rect 3673 333 3687 347
rect 3773 333 3787 347
rect 3833 333 3847 347
rect 3873 333 3887 347
rect 3893 333 3907 347
rect 3933 333 3947 347
rect 4093 333 4107 347
rect 4133 333 4147 347
rect 4193 333 4207 347
rect 4273 333 4287 347
rect 4313 333 4327 347
rect 4413 333 4427 347
rect 4453 333 4467 347
rect 4533 333 4547 347
rect 4573 333 4587 347
rect 4593 333 4607 347
rect 4633 333 4647 347
rect 4693 333 4707 347
rect 4733 333 4747 347
rect 4773 333 4787 347
rect 4933 333 4947 347
rect 4973 333 4987 347
rect 5053 333 5067 347
rect 5113 333 5127 347
rect 5193 333 5207 347
rect 5233 333 5247 347
rect 5313 333 5327 347
rect 5353 333 5367 347
rect 5373 333 5387 347
rect 5413 333 5427 347
rect 5513 333 5527 347
rect 5653 333 5667 347
rect 5693 333 5707 347
rect 5873 333 5887 347
rect 5913 333 5927 347
rect 5933 333 5947 347
rect 5973 333 5987 347
rect 6033 333 6047 347
rect 6073 333 6087 347
rect 6153 333 6167 347
rect 6193 333 6207 347
rect 6233 333 6247 347
rect 6273 333 6287 347
rect 6313 333 6327 347
rect 6353 333 6367 347
rect 6393 333 6407 347
rect 6493 333 6507 347
rect 6533 333 6547 347
rect 6613 333 6627 347
rect 613 313 627 327
rect 713 313 727 327
rect 873 313 887 327
rect 1413 313 1427 327
rect 1573 313 1587 327
rect 1973 313 1987 327
rect 2033 313 2047 327
rect 2153 313 2167 327
rect 2453 313 2467 327
rect 2873 313 2887 327
rect 3373 313 3387 327
rect 3493 313 3507 327
rect 3653 313 3667 327
rect 3733 313 3747 327
rect 3853 313 3867 327
rect 4113 313 4127 327
rect 4433 313 4447 327
rect 4613 313 4627 327
rect 4833 313 4847 327
rect 5153 313 5167 327
rect 5213 313 5227 327
rect 5393 313 5407 327
rect 5473 313 5487 327
rect 6173 313 6187 327
rect 6253 313 6267 327
rect 1513 173 1527 187
rect 1713 173 1727 187
rect 2653 173 2667 187
rect 3053 173 3067 187
rect 3253 173 3267 187
rect 6393 173 6407 187
rect 33 153 47 167
rect 113 153 127 167
rect 153 153 167 167
rect 273 153 287 167
rect 353 153 367 167
rect 393 153 407 167
rect 513 153 527 167
rect 553 153 567 167
rect 573 153 587 167
rect 613 153 627 167
rect 673 153 687 167
rect 713 153 727 167
rect 753 153 767 167
rect 833 153 847 167
rect 873 153 887 167
rect 973 153 987 167
rect 1013 153 1027 167
rect 1173 153 1187 167
rect 1213 153 1227 167
rect 1313 153 1327 167
rect 1353 153 1367 167
rect 1433 153 1447 167
rect 1653 153 1667 167
rect 1693 153 1707 167
rect 2053 153 2067 167
rect 2093 153 2107 167
rect 2193 153 2207 167
rect 2233 153 2247 167
rect 2313 153 2327 167
rect 2553 153 2567 167
rect 2593 153 2607 167
rect 2753 153 2767 167
rect 2793 153 2807 167
rect 2873 153 2887 167
rect 2953 153 2967 167
rect 2993 153 3007 167
rect 3033 153 3047 167
rect 3073 153 3087 167
rect 3113 153 3127 167
rect 3153 153 3167 167
rect 3193 153 3207 167
rect 3293 153 3307 167
rect 3373 153 3387 167
rect 3413 153 3427 167
rect 3633 153 3647 167
rect 3673 153 3687 167
rect 3693 153 3707 167
rect 3733 153 3747 167
rect 3813 153 3827 167
rect 3893 153 3907 167
rect 3933 153 3947 167
rect 4033 153 4047 167
rect 4073 153 4087 167
rect 4133 153 4147 167
rect 4173 153 4187 167
rect 4333 153 4347 167
rect 4413 153 4427 167
rect 4453 153 4467 167
rect 4553 153 4567 167
rect 4593 153 4607 167
rect 4653 153 4667 167
rect 4693 153 4707 167
rect 4853 153 4867 167
rect 4933 153 4947 167
rect 4973 153 4987 167
rect 5113 153 5127 167
rect 5153 153 5167 167
rect 5173 153 5187 167
rect 5213 153 5227 167
rect 5373 153 5387 167
rect 5453 153 5467 167
rect 5493 153 5507 167
rect 5613 153 5627 167
rect 5693 153 5707 167
rect 5733 153 5747 167
rect 5853 153 5867 167
rect 5933 153 5947 167
rect 5973 153 5987 167
rect 6093 153 6107 167
rect 6133 153 6147 167
rect 6173 153 6187 167
rect 6253 153 6267 167
rect 6293 153 6307 167
rect 6333 153 6347 167
rect 6433 153 6447 167
rect 6513 153 6527 167
rect 6553 153 6567 167
rect 1093 133 1107 147
rect 1153 133 1167 147
rect 1193 133 1207 147
rect 1493 133 1507 147
rect 1553 133 1567 147
rect 1633 133 1647 147
rect 1673 133 1687 147
rect 1733 133 1747 147
rect 1793 133 1807 147
rect 1873 133 1887 147
rect 1953 133 1967 147
rect 2033 133 2047 147
rect 2073 133 2087 147
rect 2373 133 2387 147
rect 2473 133 2487 147
rect 2533 133 2547 147
rect 2573 133 2587 147
rect 2633 133 2647 147
rect 2933 133 2947 147
rect 2973 133 2987 147
rect 3133 133 3147 147
rect 3173 133 3187 147
rect 3233 133 3247 147
rect 3553 133 3567 147
rect 3613 133 3627 147
rect 3653 133 3667 147
rect 3713 133 3727 147
rect 3753 133 3767 147
rect 4053 133 4067 147
rect 4093 133 4107 147
rect 4153 133 4167 147
rect 4193 133 4207 147
rect 4253 133 4267 147
rect 4573 133 4587 147
rect 4613 133 4627 147
rect 4673 133 4687 147
rect 4713 133 4727 147
rect 4773 133 4787 147
rect 5093 133 5107 147
rect 5133 133 5147 147
rect 5193 133 5207 147
rect 5233 133 5247 147
rect 5293 133 5307 147
rect 6113 133 6127 147
rect 6153 133 6167 147
rect 6193 133 6207 147
rect 6273 133 6287 147
rect 6313 133 6327 147
rect 6373 133 6387 147
rect 1073 113 1087 127
rect 1113 113 1127 127
rect 1533 113 1547 127
rect 1573 113 1587 127
rect 1773 113 1787 127
rect 1813 113 1827 127
rect 1853 113 1867 127
rect 1893 113 1907 127
rect 1933 113 1947 127
rect 1973 113 1987 127
rect 2353 113 2367 127
rect 2393 113 2407 127
rect 2453 113 2467 127
rect 2493 113 2507 127
rect 3533 113 3547 127
rect 3573 113 3587 127
rect 4233 113 4247 127
rect 4273 113 4287 127
rect 4753 113 4767 127
rect 4793 113 4807 127
rect 5273 113 5287 127
rect 5313 113 5327 127
<< labels >>
flabel metal1 s 6742 2 6802 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s -24 4456 -16 4464 7 FreeSans 16 0 0 0 ap_clk
port 2 nsew
flabel metal2 s 517 -23 523 -17 7 FreeSans 16 270 0 0 ap_done
port 3 nsew
flabel metal2 s 997 -23 1003 -17 7 FreeSans 16 270 0 0 ap_idle
port 4 nsew
flabel metal2 s 597 -23 603 -17 7 FreeSans 16 270 0 0 ap_ready
port 5 nsew
flabel metal3 s -24 1596 -16 1604 7 FreeSans 16 0 0 0 ap_rst
port 6 nsew
flabel metal2 s 737 -23 743 -17 7 FreeSans 16 270 0 0 ap_start
port 7 nsew
flabel metal2 s 1877 -23 1883 -17 7 FreeSans 16 270 0 0 x[7]
port 8 nsew
flabel metal2 s 2457 -23 2463 -17 7 FreeSans 16 270 0 0 x[6]
port 9 nsew
flabel metal2 s 1797 -23 1803 -17 7 FreeSans 16 270 0 0 x[5]
port 10 nsew
flabel metal2 s 1957 -23 1963 -17 7 FreeSans 16 270 0 0 x[4]
port 11 nsew
flabel metal2 s 2377 -23 2383 -17 7 FreeSans 16 270 0 0 x[3]
port 12 nsew
flabel metal2 s 1077 -23 1083 -17 7 FreeSans 16 270 0 0 x[2]
port 13 nsew
flabel metal2 s 1417 -23 1423 -17 7 FreeSans 16 270 0 0 x[1]
port 14 nsew
flabel metal2 s 1557 -23 1563 -17 7 FreeSans 16 270 0 0 x[0]
port 15 nsew
flabel metal3 s -24 3236 -16 3244 7 FreeSans 16 0 0 0 y[15]
port 16 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 y[14]
port 17 nsew
flabel metal3 s -24 3696 -16 3704 7 FreeSans 16 0 0 0 y[13]
port 18 nsew
flabel metal3 s -24 3956 -16 3964 7 FreeSans 16 0 0 0 y[12]
port 19 nsew
flabel metal3 s -24 5156 -16 5164 7 FreeSans 16 0 0 0 y[11]
port 20 nsew
flabel metal3 s -24 5616 -16 5624 7 FreeSans 16 0 0 0 y[10]
port 21 nsew
flabel metal3 s -24 5876 -16 5884 7 FreeSans 16 0 0 0 y[9]
port 22 nsew
flabel metal3 s -24 5656 -16 5664 7 FreeSans 16 0 0 0 y[8]
port 23 nsew
flabel metal3 s -24 2516 -16 2524 7 FreeSans 16 0 0 0 y[7]
port 24 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 y[6]
port 25 nsew
flabel metal3 s -24 3476 -16 3484 7 FreeSans 16 0 0 0 y[5]
port 26 nsew
flabel metal3 s -24 3996 -16 4004 7 FreeSans 16 0 0 0 y[4]
port 27 nsew
flabel metal3 s -24 4196 -16 4204 7 FreeSans 16 0 0 0 y[3]
port 28 nsew
flabel metal3 s -24 4956 -16 4964 7 FreeSans 16 0 0 0 y[2]
port 29 nsew
flabel metal3 s -24 4916 -16 4924 7 FreeSans 16 0 0 0 y[1]
port 30 nsew
flabel metal3 s -24 3736 -16 3744 7 FreeSans 16 0 0 0 y[0]
port 31 nsew
flabel metal2 s 677 -23 683 -17 7 FreeSans 16 270 0 0 y_ap_vld
port 32 nsew
rlabel metal1 4 242 256 258 0 _1607_.gnd
rlabel metal1 4 2 256 18 0 _1607_.vdd
rlabel metal2 153 153 167 167 0 _1607_.D
rlabel metal2 113 153 127 167 0 _1607_.CLK
rlabel metal2 33 153 47 167 0 _1607_.Q
rlabel metal1 244 242 496 258 0 _1606_.gnd
rlabel metal1 244 2 496 18 0 _1606_.vdd
rlabel metal2 393 153 407 167 0 _1606_.D
rlabel metal2 353 153 367 167 0 _1606_.CLK
rlabel metal2 273 153 287 167 0 _1606_.Q
rlabel metal1 4 242 256 258 0 _1605_.gnd
rlabel metal1 4 482 256 498 0 _1605_.vdd
rlabel metal2 153 333 167 347 0 _1605_.D
rlabel metal2 113 333 127 347 0 _1605_.CLK
rlabel metal2 33 333 47 347 0 _1605_.Q
rlabel metal1 244 242 496 258 0 _1484_.gnd
rlabel metal1 244 482 496 498 0 _1484_.vdd
rlabel metal2 333 333 347 347 0 _1484_.D
rlabel metal2 373 333 387 347 0 _1484_.CLK
rlabel metal2 453 333 467 347 0 _1484_.Q
rlabel metal1 484 242 576 258 0 _3028_.gnd
rlabel metal1 484 2 576 18 0 _3028_.vdd
rlabel metal2 553 153 567 167 0 _3028_.A
rlabel metal2 513 153 527 167 0 _3028_.Y
rlabel metal1 484 242 596 258 0 _1473_.gnd
rlabel metal1 484 482 596 498 0 _1473_.vdd
rlabel metal2 493 353 507 367 0 _1473_.A
rlabel metal2 513 373 527 387 0 _1473_.B
rlabel metal2 533 353 547 367 0 _1473_.C
rlabel metal2 553 373 567 387 0 _1473_.Y
rlabel metal1 644 242 736 258 0 _3047_.gnd
rlabel metal1 644 2 736 18 0 _3047_.vdd
rlabel metal2 713 153 727 167 0 _3047_.A
rlabel metal2 673 153 687 167 0 _3047_.Y
rlabel metal1 564 242 656 258 0 _3030_.gnd
rlabel metal1 564 2 656 18 0 _3030_.vdd
rlabel metal2 573 153 587 167 0 _3030_.A
rlabel metal2 613 153 627 167 0 _3030_.Y
rlabel metal1 724 242 976 258 0 _1485_.gnd
rlabel metal1 724 2 976 18 0 _1485_.vdd
rlabel metal2 873 153 887 167 0 _1485_.D
rlabel metal2 833 153 847 167 0 _1485_.CLK
rlabel metal2 753 153 767 167 0 _1485_.Q
rlabel metal1 584 242 676 258 0 _1474_.gnd
rlabel metal1 584 482 676 498 0 _1474_.vdd
rlabel metal2 633 333 647 347 0 _1474_.B
rlabel metal2 593 333 607 347 0 _1474_.A
rlabel metal2 613 313 627 327 0 _1474_.Y
rlabel metal1 664 242 756 258 0 _1414_.gnd
rlabel metal1 664 482 756 498 0 _1414_.vdd
rlabel metal2 693 333 707 347 0 _1414_.B
rlabel metal2 733 333 747 347 0 _1414_.A
rlabel metal2 713 313 727 327 0 _1414_.Y
rlabel metal1 744 242 836 258 0 _1452_.gnd
rlabel metal1 744 482 836 498 0 _1452_.vdd
rlabel metal2 753 373 767 387 0 _1452_.A
rlabel metal2 793 373 807 387 0 _1452_.B
rlabel metal2 773 353 787 367 0 _1452_.Y
rlabel metal1 964 242 1056 258 0 _3029_.gnd
rlabel metal1 964 2 1056 18 0 _3029_.vdd
rlabel metal2 973 153 987 167 0 _3029_.A
rlabel metal2 1013 153 1027 167 0 _3029_.Y
rlabel metal1 884 242 1136 258 0 _1488_.gnd
rlabel metal1 884 482 1136 498 0 _1488_.vdd
rlabel metal2 973 333 987 347 0 _1488_.D
rlabel metal2 1013 333 1027 347 0 _1488_.CLK
rlabel metal2 1093 333 1107 347 0 _1488_.Q
rlabel metal1 824 242 896 258 0 _1413_.gnd
rlabel metal1 824 482 896 498 0 _1413_.vdd
rlabel metal2 873 313 887 327 0 _1413_.A
rlabel metal2 853 353 867 367 0 _1413_.Y
rlabel metal1 1044 242 1136 258 0 _1425_.gnd
rlabel metal1 1044 2 1136 18 0 _1425_.vdd
rlabel metal2 1113 113 1127 127 0 _1425_.A
rlabel metal2 1073 113 1087 127 0 _1425_.B
rlabel metal2 1093 133 1107 147 0 _1425_.Y
rlabel metal1 1204 242 1296 258 0 BUFX2_insert41.gnd
rlabel metal1 1204 482 1296 498 0 BUFX2_insert41.vdd
rlabel metal2 1213 333 1227 347 0 BUFX2_insert41.A
rlabel metal2 1253 333 1267 347 0 BUFX2_insert41.Y
rlabel metal1 1124 242 1216 258 0 BUFX2_insert39.gnd
rlabel metal1 1124 482 1216 498 0 BUFX2_insert39.vdd
rlabel metal2 1193 333 1207 347 0 BUFX2_insert39.A
rlabel metal2 1153 333 1167 347 0 BUFX2_insert39.Y
rlabel metal1 1284 242 1376 258 0 BUFX2_insert38.gnd
rlabel metal1 1284 482 1376 498 0 BUFX2_insert38.vdd
rlabel metal2 1293 333 1307 347 0 BUFX2_insert38.A
rlabel metal2 1333 333 1347 347 0 BUFX2_insert38.Y
rlabel metal1 1224 242 1476 258 0 _1490_.gnd
rlabel metal1 1224 2 1476 18 0 _1490_.vdd
rlabel metal2 1313 153 1327 167 0 _1490_.D
rlabel metal2 1353 153 1367 167 0 _1490_.CLK
rlabel metal2 1433 153 1447 167 0 _1490_.Q
rlabel metal1 1124 242 1236 258 0 _1426_.gnd
rlabel metal1 1124 2 1236 18 0 _1426_.vdd
rlabel metal2 1213 153 1227 167 0 _1426_.A
rlabel metal2 1193 133 1207 147 0 _1426_.B
rlabel metal2 1153 133 1167 147 0 _1426_.C
rlabel metal2 1173 153 1187 167 0 _1426_.Y
rlabel metal1 1584 242 1696 258 0 _1441_.gnd
rlabel metal1 1584 482 1696 498 0 _1441_.vdd
rlabel metal2 1593 333 1607 347 0 _1441_.A
rlabel metal2 1613 353 1627 367 0 _1441_.B
rlabel metal2 1653 353 1667 367 0 _1441_.C
rlabel metal2 1633 333 1647 347 0 _1441_.Y
rlabel metal1 1424 242 1536 258 0 _1435_.gnd
rlabel metal1 1424 482 1536 498 0 _1435_.vdd
rlabel metal2 1433 333 1447 347 0 _1435_.A
rlabel metal2 1453 353 1467 367 0 _1435_.B
rlabel metal2 1493 353 1507 367 0 _1435_.C
rlabel metal2 1473 333 1487 347 0 _1435_.Y
rlabel metal1 1604 242 1716 258 0 _1420_.gnd
rlabel metal1 1604 2 1716 18 0 _1420_.vdd
rlabel metal2 1693 153 1707 167 0 _1420_.A
rlabel metal2 1673 133 1687 147 0 _1420_.B
rlabel metal2 1633 133 1647 147 0 _1420_.C
rlabel metal2 1653 153 1667 167 0 _1420_.Y
rlabel metal1 1524 242 1596 258 0 _1439_.gnd
rlabel metal1 1524 482 1596 498 0 _1439_.vdd
rlabel metal2 1573 313 1587 327 0 _1439_.A
rlabel metal2 1553 353 1567 367 0 _1439_.Y
rlabel metal1 1364 242 1436 258 0 _1433_.gnd
rlabel metal1 1364 482 1436 498 0 _1433_.vdd
rlabel metal2 1413 313 1427 327 0 _1433_.A
rlabel metal2 1393 353 1407 367 0 _1433_.Y
rlabel metal1 1464 242 1536 258 0 _1424_.gnd
rlabel metal1 1464 2 1536 18 0 _1424_.vdd
rlabel metal2 1513 173 1527 187 0 _1424_.A
rlabel metal2 1493 133 1507 147 0 _1424_.Y
rlabel metal1 1524 242 1616 258 0 _1419_.gnd
rlabel metal1 1524 2 1616 18 0 _1419_.vdd
rlabel metal2 1533 113 1547 127 0 _1419_.A
rlabel metal2 1573 113 1587 127 0 _1419_.B
rlabel metal2 1553 133 1567 147 0 _1419_.Y
rlabel metal1 1684 242 1936 258 0 _3025_.gnd
rlabel metal1 1684 482 1936 498 0 _3025_.vdd
rlabel metal2 1773 333 1787 347 0 _3025_.D
rlabel metal2 1813 333 1827 347 0 _3025_.CLK
rlabel metal2 1893 333 1907 347 0 _3025_.Q
rlabel metal1 1704 242 1776 258 0 _1418_.gnd
rlabel metal1 1704 2 1776 18 0 _1418_.vdd
rlabel metal2 1713 173 1727 187 0 _1418_.A
rlabel metal2 1733 133 1747 147 0 _1418_.Y
rlabel metal1 1844 242 1936 258 0 _1440_.gnd
rlabel metal1 1844 2 1936 18 0 _1440_.vdd
rlabel metal2 1853 113 1867 127 0 _1440_.A
rlabel metal2 1893 113 1907 127 0 _1440_.B
rlabel metal2 1873 133 1887 147 0 _1440_.Y
rlabel metal1 1764 242 1856 258 0 _1434_.gnd
rlabel metal1 1764 2 1856 18 0 _1434_.vdd
rlabel metal2 1773 113 1787 127 0 _1434_.A
rlabel metal2 1813 113 1827 127 0 _1434_.B
rlabel metal2 1793 133 1807 147 0 _1434_.Y
rlabel metal1 2104 242 2356 258 0 _1492_.gnd
rlabel metal1 2104 2 2356 18 0 _1492_.vdd
rlabel metal2 2193 153 2207 167 0 _1492_.D
rlabel metal2 2233 153 2247 167 0 _1492_.CLK
rlabel metal2 2313 153 2327 167 0 _1492_.Q
rlabel metal1 2004 242 2116 258 0 _1432_.gnd
rlabel metal1 2004 2 2116 18 0 _1432_.vdd
rlabel metal2 2093 153 2107 167 0 _1432_.A
rlabel metal2 2073 133 2087 147 0 _1432_.B
rlabel metal2 2033 133 2047 147 0 _1432_.C
rlabel metal2 2053 153 2067 167 0 _1432_.Y
rlabel metal1 2044 242 2156 258 0 _1429_.gnd
rlabel metal1 2044 482 2156 498 0 _1429_.vdd
rlabel metal2 2053 333 2067 347 0 _1429_.A
rlabel metal2 2073 353 2087 367 0 _1429_.B
rlabel metal2 2113 353 2127 367 0 _1429_.C
rlabel metal2 2093 333 2107 347 0 _1429_.Y
rlabel metal1 1924 242 1996 258 0 _1430_.gnd
rlabel metal1 1924 482 1996 498 0 _1430_.vdd
rlabel metal2 1973 313 1987 327 0 _1430_.A
rlabel metal2 1953 353 1967 367 0 _1430_.Y
rlabel metal1 1984 242 2056 258 0 _1427_.gnd
rlabel metal1 1984 482 2056 498 0 _1427_.vdd
rlabel metal2 2033 313 2047 327 0 _1427_.A
rlabel metal2 2013 353 2027 367 0 _1427_.Y
rlabel metal1 1924 242 2016 258 0 _1431_.gnd
rlabel metal1 1924 2 2016 18 0 _1431_.vdd
rlabel metal2 1933 113 1947 127 0 _1431_.A
rlabel metal2 1973 113 1987 127 0 _1431_.B
rlabel metal2 1953 133 1967 147 0 _1431_.Y
rlabel metal1 2204 242 2336 258 0 _2939_.gnd
rlabel metal1 2204 482 2336 498 0 _2939_.vdd
rlabel metal2 2213 333 2227 347 0 _2939_.A
rlabel metal2 2233 353 2247 367 0 _2939_.B
rlabel metal2 2293 333 2307 347 0 _2939_.C
rlabel metal2 2253 333 2267 347 0 _2939_.Y
rlabel metal2 2273 353 2287 367 0 _2939_.D
rlabel metal1 2324 242 2436 258 0 _2938_.gnd
rlabel metal1 2324 482 2436 498 0 _2938_.vdd
rlabel metal2 2413 333 2427 347 0 _2938_.A
rlabel metal2 2393 353 2407 367 0 _2938_.B
rlabel metal2 2353 353 2367 367 0 _2938_.C
rlabel metal2 2373 333 2387 347 0 _2938_.Y
rlabel metal1 2144 242 2216 258 0 _2936_.gnd
rlabel metal1 2144 482 2216 498 0 _2936_.vdd
rlabel metal2 2153 313 2167 327 0 _2936_.A
rlabel metal2 2173 353 2187 367 0 _2936_.Y
rlabel metal1 2344 242 2436 258 0 _1428_.gnd
rlabel metal1 2344 2 2436 18 0 _1428_.vdd
rlabel metal2 2353 113 2367 127 0 _1428_.A
rlabel metal2 2393 113 2407 127 0 _1428_.B
rlabel metal2 2373 133 2387 147 0 _1428_.Y
rlabel metal1 2504 242 2756 258 0 _3002_.gnd
rlabel metal1 2504 482 2756 498 0 _3002_.vdd
rlabel metal2 2593 333 2607 347 0 _3002_.D
rlabel metal2 2633 333 2647 347 0 _3002_.CLK
rlabel metal2 2713 333 2727 347 0 _3002_.Q
rlabel metal1 2664 242 2916 258 0 _1494_.gnd
rlabel metal1 2664 2 2916 18 0 _1494_.vdd
rlabel metal2 2753 153 2767 167 0 _1494_.D
rlabel metal2 2793 153 2807 167 0 _1494_.CLK
rlabel metal2 2873 153 2887 167 0 _1494_.Q
rlabel metal1 2504 242 2616 258 0 _1438_.gnd
rlabel metal1 2504 2 2616 18 0 _1438_.vdd
rlabel metal2 2593 153 2607 167 0 _1438_.A
rlabel metal2 2573 133 2587 147 0 _1438_.B
rlabel metal2 2533 133 2547 147 0 _1438_.C
rlabel metal2 2553 153 2567 167 0 _1438_.Y
rlabel metal1 2424 242 2516 258 0 _2937_.gnd
rlabel metal1 2424 482 2516 498 0 _2937_.vdd
rlabel metal2 2473 333 2487 347 0 _2937_.B
rlabel metal2 2433 333 2447 347 0 _2937_.A
rlabel metal2 2453 313 2467 327 0 _2937_.Y
rlabel metal1 2604 242 2676 258 0 _1436_.gnd
rlabel metal1 2604 2 2676 18 0 _1436_.vdd
rlabel metal2 2653 173 2667 187 0 _1436_.A
rlabel metal2 2633 133 2647 147 0 _1436_.Y
rlabel metal1 2424 242 2516 258 0 _1437_.gnd
rlabel metal1 2424 2 2516 18 0 _1437_.vdd
rlabel metal2 2493 113 2507 127 0 _1437_.A
rlabel metal2 2453 113 2467 127 0 _1437_.B
rlabel metal2 2473 133 2487 147 0 _1437_.Y
rlabel metal1 2924 242 3176 258 0 _2994_.gnd
rlabel metal1 2924 482 3176 498 0 _2994_.vdd
rlabel metal2 3013 333 3027 347 0 _2994_.D
rlabel metal2 3053 333 3067 347 0 _2994_.CLK
rlabel metal2 3133 333 3147 347 0 _2994_.Q
rlabel metal1 2904 242 3016 258 0 _2942_.gnd
rlabel metal1 2904 2 3016 18 0 _2942_.vdd
rlabel metal2 2993 153 3007 167 0 _2942_.A
rlabel metal2 2973 133 2987 147 0 _2942_.B
rlabel metal2 2933 133 2947 147 0 _2942_.C
rlabel metal2 2953 153 2967 167 0 _2942_.Y
rlabel metal1 2744 242 2856 258 0 _2836_.gnd
rlabel metal1 2744 482 2856 498 0 _2836_.vdd
rlabel metal2 2833 333 2847 347 0 _2836_.A
rlabel metal2 2813 353 2827 367 0 _2836_.B
rlabel metal2 2773 353 2787 367 0 _2836_.C
rlabel metal2 2793 333 2807 347 0 _2836_.Y
rlabel metal1 2844 242 2936 258 0 _2834_.gnd
rlabel metal1 2844 482 2936 498 0 _2834_.vdd
rlabel metal2 2893 333 2907 347 0 _2834_.B
rlabel metal2 2853 333 2867 347 0 _2834_.A
rlabel metal2 2873 313 2887 327 0 _2834_.Y
rlabel metal1 3084 242 3216 258 0 _2943_.gnd
rlabel metal1 3084 2 3216 18 0 _2943_.vdd
rlabel metal2 3193 153 3207 167 0 _2943_.A
rlabel metal2 3173 133 3187 147 0 _2943_.B
rlabel metal2 3113 153 3127 167 0 _2943_.C
rlabel metal2 3153 153 3167 167 0 _2943_.Y
rlabel metal2 3133 133 3147 147 0 _2943_.D
rlabel metal1 3004 242 3096 258 0 _2941_.gnd
rlabel metal1 3004 2 3096 18 0 _2941_.vdd
rlabel metal2 3033 153 3047 167 0 _2941_.B
rlabel metal2 3073 153 3087 167 0 _2941_.A
rlabel metal2 3053 173 3067 187 0 _2941_.Y
rlabel metal1 3204 242 3276 258 0 _2940_.gnd
rlabel metal1 3204 2 3276 18 0 _2940_.vdd
rlabel metal2 3253 173 3267 187 0 _2940_.A
rlabel metal2 3233 133 3247 147 0 _2940_.Y
rlabel metal1 3164 242 3256 258 0 _2797_.gnd
rlabel metal1 3164 482 3256 498 0 _2797_.vdd
rlabel metal2 3173 373 3187 387 0 _2797_.A
rlabel metal2 3213 373 3227 387 0 _2797_.B
rlabel metal2 3193 353 3207 367 0 _2797_.Y
rlabel metal1 3264 242 3516 258 0 _3026_.gnd
rlabel metal1 3264 2 3516 18 0 _3026_.vdd
rlabel metal2 3413 153 3427 167 0 _3026_.D
rlabel metal2 3373 153 3387 167 0 _3026_.CLK
rlabel metal2 3293 153 3307 167 0 _3026_.Q
rlabel metal1 3244 242 3356 258 0 _2800_.gnd
rlabel metal1 3244 482 3356 498 0 _2800_.vdd
rlabel metal2 3333 333 3347 347 0 _2800_.A
rlabel metal2 3313 353 3327 367 0 _2800_.B
rlabel metal2 3273 353 3287 367 0 _2800_.C
rlabel metal2 3293 333 3307 347 0 _2800_.Y
rlabel metal1 3344 242 3436 258 0 _2798_.gnd
rlabel metal1 3344 482 3436 498 0 _2798_.vdd
rlabel metal2 3393 333 3407 347 0 _2798_.B
rlabel metal2 3353 333 3367 347 0 _2798_.A
rlabel metal2 3373 313 3387 327 0 _2798_.Y
rlabel metal1 3424 242 3536 258 0 _2835_.gnd
rlabel metal1 3424 482 3536 498 0 _2835_.vdd
rlabel metal2 3513 353 3527 367 0 _2835_.A
rlabel metal2 3493 313 3507 327 0 _2835_.B
rlabel metal2 3473 353 3487 367 0 _2835_.C
rlabel metal2 3453 333 3467 347 0 _2835_.Y
rlabel metal1 3524 242 3636 258 0 _2799_.gnd
rlabel metal1 3524 482 3636 498 0 _2799_.vdd
rlabel metal2 3533 333 3547 347 0 _2799_.A
rlabel metal2 3553 353 3567 367 0 _2799_.B
rlabel metal2 3593 353 3607 367 0 _2799_.C
rlabel metal2 3573 333 3587 347 0 _2799_.Y
rlabel metal1 3584 242 3696 258 0 _2796_.gnd
rlabel metal1 3584 2 3696 18 0 _2796_.vdd
rlabel metal2 3673 153 3687 167 0 _2796_.A
rlabel metal2 3653 133 3667 147 0 _2796_.B
rlabel metal2 3613 133 3627 147 0 _2796_.C
rlabel metal2 3633 153 3647 167 0 _2796_.Y
rlabel metal1 3684 242 3796 258 0 _2795_.gnd
rlabel metal1 3684 2 3796 18 0 _2795_.vdd
rlabel metal2 3693 153 3707 167 0 _2795_.A
rlabel metal2 3713 133 3727 147 0 _2795_.B
rlabel metal2 3753 133 3767 147 0 _2795_.C
rlabel metal2 3733 153 3747 167 0 _2795_.Y
rlabel metal1 3624 242 3716 258 0 _2794_.gnd
rlabel metal1 3624 482 3716 498 0 _2794_.vdd
rlabel metal2 3673 333 3687 347 0 _2794_.B
rlabel metal2 3633 333 3647 347 0 _2794_.A
rlabel metal2 3653 313 3667 327 0 _2794_.Y
rlabel metal1 3504 242 3596 258 0 _2793_.gnd
rlabel metal1 3504 2 3596 18 0 _2793_.vdd
rlabel metal2 3573 113 3587 127 0 _2793_.A
rlabel metal2 3533 113 3547 127 0 _2793_.B
rlabel metal2 3553 133 3567 147 0 _2793_.Y
rlabel metal1 3704 242 3816 258 0 _2827_.gnd
rlabel metal1 3704 482 3816 498 0 _2827_.vdd
rlabel metal2 3713 353 3727 367 0 _2827_.A
rlabel metal2 3733 313 3747 327 0 _2827_.B
rlabel metal2 3753 353 3767 367 0 _2827_.C
rlabel metal2 3773 333 3787 347 0 _2827_.Y
rlabel metal1 3784 242 4036 258 0 _2993_.gnd
rlabel metal1 3784 2 4036 18 0 _2993_.vdd
rlabel metal2 3933 153 3947 167 0 _2993_.D
rlabel metal2 3893 153 3907 167 0 _2993_.CLK
rlabel metal2 3813 153 3827 167 0 _2993_.Q
rlabel metal1 3884 242 3996 258 0 _2828_.gnd
rlabel metal1 3884 482 3996 498 0 _2828_.vdd
rlabel metal2 3893 333 3907 347 0 _2828_.A
rlabel metal2 3913 353 3927 367 0 _2828_.B
rlabel metal2 3953 353 3967 367 0 _2828_.C
rlabel metal2 3933 333 3947 347 0 _2828_.Y
rlabel metal1 3804 242 3896 258 0 _2826_.gnd
rlabel metal1 3804 482 3896 498 0 _2826_.vdd
rlabel metal2 3833 333 3847 347 0 _2826_.B
rlabel metal2 3873 333 3887 347 0 _2826_.A
rlabel metal2 3853 313 3867 327 0 _2826_.Y
rlabel metal1 3984 242 4096 258 0 _2825_.gnd
rlabel metal1 3984 482 4096 498 0 _2825_.vdd
rlabel metal2 4073 353 4087 367 0 _2825_.A
rlabel metal2 4053 373 4067 387 0 _2825_.B
rlabel metal2 4033 353 4047 367 0 _2825_.C
rlabel metal2 4013 373 4027 387 0 _2825_.Y
rlabel metal1 4164 242 4416 258 0 _3000_.gnd
rlabel metal1 4164 482 4416 498 0 _3000_.vdd
rlabel metal2 4313 333 4327 347 0 _3000_.D
rlabel metal2 4273 333 4287 347 0 _3000_.CLK
rlabel metal2 4193 333 4207 347 0 _3000_.Q
rlabel metal1 4124 242 4236 258 0 _2792_.gnd
rlabel metal1 4124 2 4236 18 0 _2792_.vdd
rlabel metal2 4133 153 4147 167 0 _2792_.A
rlabel metal2 4153 133 4167 147 0 _2792_.B
rlabel metal2 4193 133 4207 147 0 _2792_.C
rlabel metal2 4173 153 4187 167 0 _2792_.Y
rlabel metal1 4024 242 4136 258 0 _2791_.gnd
rlabel metal1 4024 2 4136 18 0 _2791_.vdd
rlabel metal2 4033 153 4047 167 0 _2791_.A
rlabel metal2 4053 133 4067 147 0 _2791_.B
rlabel metal2 4093 133 4107 147 0 _2791_.C
rlabel metal2 4073 153 4087 167 0 _2791_.Y
rlabel metal1 4084 242 4176 258 0 _2790_.gnd
rlabel metal1 4084 482 4176 498 0 _2790_.vdd
rlabel metal2 4133 333 4147 347 0 _2790_.B
rlabel metal2 4093 333 4107 347 0 _2790_.A
rlabel metal2 4113 313 4127 327 0 _2790_.Y
rlabel metal1 4224 242 4316 258 0 _2789_.gnd
rlabel metal1 4224 2 4316 18 0 _2789_.vdd
rlabel metal2 4233 113 4247 127 0 _2789_.A
rlabel metal2 4273 113 4287 127 0 _2789_.B
rlabel metal2 4253 133 4267 147 0 _2789_.Y
rlabel metal1 4304 242 4556 258 0 _2992_.gnd
rlabel metal1 4304 2 4556 18 0 _2992_.vdd
rlabel metal2 4453 153 4467 167 0 _2992_.D
rlabel metal2 4413 153 4427 167 0 _2992_.CLK
rlabel metal2 4333 153 4347 167 0 _2992_.Q
rlabel metal1 4484 242 4596 258 0 _2918_.gnd
rlabel metal1 4484 482 4596 498 0 _2918_.vdd
rlabel metal2 4573 333 4587 347 0 _2918_.A
rlabel metal2 4553 353 4567 367 0 _2918_.B
rlabel metal2 4513 353 4527 367 0 _2918_.C
rlabel metal2 4533 333 4547 347 0 _2918_.Y
rlabel metal1 4404 242 4496 258 0 _2786_.gnd
rlabel metal1 4404 482 4496 498 0 _2786_.vdd
rlabel metal2 4453 333 4467 347 0 _2786_.B
rlabel metal2 4413 333 4427 347 0 _2786_.A
rlabel metal2 4433 313 4447 327 0 _2786_.Y
rlabel metal1 4664 242 4796 258 0 _2919_.gnd
rlabel metal1 4664 482 4796 498 0 _2919_.vdd
rlabel metal2 4773 333 4787 347 0 _2919_.A
rlabel metal2 4753 353 4767 367 0 _2919_.B
rlabel metal2 4693 333 4707 347 0 _2919_.C
rlabel metal2 4733 333 4747 347 0 _2919_.Y
rlabel metal2 4713 353 4727 367 0 _2919_.D
rlabel metal1 4644 242 4756 258 0 _2788_.gnd
rlabel metal1 4644 2 4756 18 0 _2788_.vdd
rlabel metal2 4653 153 4667 167 0 _2788_.A
rlabel metal2 4673 133 4687 147 0 _2788_.B
rlabel metal2 4713 133 4727 147 0 _2788_.C
rlabel metal2 4693 153 4707 167 0 _2788_.Y
rlabel metal1 4544 242 4656 258 0 _2787_.gnd
rlabel metal1 4544 2 4656 18 0 _2787_.vdd
rlabel metal2 4553 153 4567 167 0 _2787_.A
rlabel metal2 4573 133 4587 147 0 _2787_.B
rlabel metal2 4613 133 4627 147 0 _2787_.C
rlabel metal2 4593 153 4607 167 0 _2787_.Y
rlabel metal1 4584 242 4676 258 0 _2916_.gnd
rlabel metal1 4584 482 4676 498 0 _2916_.vdd
rlabel metal2 4633 333 4647 347 0 _2916_.B
rlabel metal2 4593 333 4607 347 0 _2916_.A
rlabel metal2 4613 313 4627 327 0 _2916_.Y
rlabel metal1 4784 242 4856 258 0 _2913_.gnd
rlabel metal1 4784 482 4856 498 0 _2913_.vdd
rlabel metal2 4833 313 4847 327 0 _2913_.A
rlabel metal2 4813 353 4827 367 0 _2913_.Y
rlabel metal1 4744 242 4836 258 0 _2785_.gnd
rlabel metal1 4744 2 4836 18 0 _2785_.vdd
rlabel metal2 4753 113 4767 127 0 _2785_.A
rlabel metal2 4793 113 4807 127 0 _2785_.B
rlabel metal2 4773 133 4787 147 0 _2785_.Y
rlabel metal1 4844 242 5096 258 0 _3020_.gnd
rlabel metal1 4844 482 5096 498 0 _3020_.vdd
rlabel metal2 4933 333 4947 347 0 _3020_.D
rlabel metal2 4973 333 4987 347 0 _3020_.CLK
rlabel metal2 5053 333 5067 347 0 _3020_.Q
rlabel metal1 4824 242 5076 258 0 _2991_.gnd
rlabel metal1 4824 2 5076 18 0 _2991_.vdd
rlabel metal2 4973 153 4987 167 0 _2991_.D
rlabel metal2 4933 153 4947 167 0 _2991_.CLK
rlabel metal2 4853 153 4867 167 0 _2991_.Q
rlabel metal1 5064 242 5176 258 0 _2775_.gnd
rlabel metal1 5064 2 5176 18 0 _2775_.vdd
rlabel metal2 5153 153 5167 167 0 _2775_.A
rlabel metal2 5133 133 5147 147 0 _2775_.B
rlabel metal2 5093 133 5107 147 0 _2775_.C
rlabel metal2 5113 153 5127 167 0 _2775_.Y
rlabel metal1 5264 242 5376 258 0 _2812_.gnd
rlabel metal1 5264 482 5376 498 0 _2812_.vdd
rlabel metal2 5353 333 5367 347 0 _2812_.A
rlabel metal2 5333 353 5347 367 0 _2812_.B
rlabel metal2 5293 353 5307 367 0 _2812_.C
rlabel metal2 5313 333 5327 347 0 _2812_.Y
rlabel metal1 5164 242 5276 258 0 _2776_.gnd
rlabel metal1 5164 2 5276 18 0 _2776_.vdd
rlabel metal2 5173 153 5187 167 0 _2776_.A
rlabel metal2 5193 133 5207 147 0 _2776_.B
rlabel metal2 5233 133 5247 147 0 _2776_.C
rlabel metal2 5213 153 5227 167 0 _2776_.Y
rlabel metal1 5184 242 5276 258 0 _2774_.gnd
rlabel metal1 5184 482 5276 498 0 _2774_.vdd
rlabel metal2 5233 333 5247 347 0 _2774_.B
rlabel metal2 5193 333 5207 347 0 _2774_.A
rlabel metal2 5213 313 5227 327 0 _2774_.Y
rlabel metal1 5264 242 5356 258 0 _2771_.gnd
rlabel metal1 5264 2 5356 18 0 _2771_.vdd
rlabel metal2 5273 113 5287 127 0 _2771_.A
rlabel metal2 5313 113 5327 127 0 _2771_.B
rlabel metal2 5293 133 5307 147 0 _2771_.Y
rlabel metal1 5084 242 5196 258 0 _2811_.gnd
rlabel metal1 5084 482 5196 498 0 _2811_.vdd
rlabel metal2 5173 353 5187 367 0 _2811_.A
rlabel metal2 5153 313 5167 327 0 _2811_.B
rlabel metal2 5133 353 5147 367 0 _2811_.C
rlabel metal2 5113 333 5127 347 0 _2811_.Y
rlabel metal1 5584 242 5836 258 0 _2997_.gnd
rlabel metal1 5584 2 5836 18 0 _2997_.vdd
rlabel metal2 5733 153 5747 167 0 _2997_.D
rlabel metal2 5693 153 5707 167 0 _2997_.CLK
rlabel metal2 5613 153 5627 167 0 _2997_.Q
rlabel metal1 5344 242 5596 258 0 _2988_.gnd
rlabel metal1 5344 2 5596 18 0 _2988_.vdd
rlabel metal2 5493 153 5507 167 0 _2988_.D
rlabel metal2 5453 153 5467 167 0 _2988_.CLK
rlabel metal2 5373 153 5387 167 0 _2988_.Q
rlabel metal1 5364 242 5456 258 0 _2808_.gnd
rlabel metal1 5364 482 5456 498 0 _2808_.vdd
rlabel metal2 5413 333 5427 347 0 _2808_.B
rlabel metal2 5373 333 5387 347 0 _2808_.A
rlabel metal2 5393 313 5407 327 0 _2808_.Y
rlabel metal1 5444 242 5556 258 0 _2815_.gnd
rlabel metal1 5444 482 5556 498 0 _2815_.vdd
rlabel metal2 5453 353 5467 367 0 _2815_.A
rlabel metal2 5473 313 5487 327 0 _2815_.B
rlabel metal2 5493 353 5507 367 0 _2815_.C
rlabel metal2 5513 333 5527 347 0 _2815_.Y
rlabel metal1 5544 242 5656 258 0 _2813_.gnd
rlabel metal1 5544 482 5656 498 0 _2813_.vdd
rlabel metal2 5553 353 5567 367 0 _2813_.A
rlabel metal2 5573 373 5587 387 0 _2813_.B
rlabel metal2 5593 353 5607 367 0 _2813_.C
rlabel metal2 5613 373 5627 387 0 _2813_.Y
rlabel metal1 5824 242 6076 258 0 _2989_.gnd
rlabel metal1 5824 2 6076 18 0 _2989_.vdd
rlabel metal2 5973 153 5987 167 0 _2989_.D
rlabel metal2 5933 153 5947 167 0 _2989_.CLK
rlabel metal2 5853 153 5867 167 0 _2989_.Q
rlabel metal1 5644 242 5756 258 0 _2816_.gnd
rlabel metal1 5644 482 5756 498 0 _2816_.vdd
rlabel metal2 5653 333 5667 347 0 _2816_.A
rlabel metal2 5673 353 5687 367 0 _2816_.B
rlabel metal2 5713 353 5727 367 0 _2816_.C
rlabel metal2 5693 333 5707 347 0 _2816_.Y
rlabel metal1 5824 242 5936 258 0 _2780_.gnd
rlabel metal1 5824 482 5936 498 0 _2780_.vdd
rlabel metal2 5913 333 5927 347 0 _2780_.A
rlabel metal2 5893 353 5907 367 0 _2780_.B
rlabel metal2 5853 353 5867 367 0 _2780_.C
rlabel metal2 5873 333 5887 347 0 _2780_.Y
rlabel metal1 5744 242 5836 258 0 _2777_.gnd
rlabel metal1 5744 482 5836 498 0 _2777_.vdd
rlabel metal2 5813 373 5827 387 0 _2777_.A
rlabel metal2 5773 373 5787 387 0 _2777_.B
rlabel metal2 5793 353 5807 367 0 _2777_.Y
rlabel metal1 6024 242 6136 258 0 _2946_.gnd
rlabel metal1 6024 482 6136 498 0 _2946_.vdd
rlabel metal2 6033 333 6047 347 0 _2946_.A
rlabel metal2 6053 353 6067 367 0 _2946_.B
rlabel metal2 6093 353 6107 367 0 _2946_.C
rlabel metal2 6073 333 6087 347 0 _2946_.Y
rlabel metal1 6124 242 6236 258 0 _2926_.gnd
rlabel metal1 6124 2 6236 18 0 _2926_.vdd
rlabel metal2 6133 153 6147 167 0 _2926_.A
rlabel metal2 6153 133 6167 147 0 _2926_.B
rlabel metal2 6193 133 6207 147 0 _2926_.C
rlabel metal2 6173 153 6187 167 0 _2926_.Y
rlabel metal1 5924 242 6036 258 0 _2779_.gnd
rlabel metal1 5924 482 6036 498 0 _2779_.vdd
rlabel metal2 5933 333 5947 347 0 _2779_.A
rlabel metal2 5953 353 5967 367 0 _2779_.B
rlabel metal2 5993 353 6007 367 0 _2779_.C
rlabel metal2 5973 333 5987 347 0 _2779_.Y
rlabel metal1 6124 242 6216 258 0 _2925_.gnd
rlabel metal1 6124 482 6216 498 0 _2925_.vdd
rlabel metal2 6153 333 6167 347 0 _2925_.B
rlabel metal2 6193 333 6207 347 0 _2925_.A
rlabel metal2 6173 313 6187 327 0 _2925_.Y
rlabel metal1 6064 242 6136 258 0 _2770_.gnd
rlabel metal1 6064 2 6136 18 0 _2770_.vdd
rlabel metal2 6113 133 6127 147 0 _2770_.A
rlabel metal2 6093 153 6107 167 0 _2770_.Y
rlabel metal1 6404 242 6656 258 0 _3027_.gnd
rlabel metal1 6404 482 6656 498 0 _3027_.vdd
rlabel metal2 6493 333 6507 347 0 _3027_.D
rlabel metal2 6533 333 6547 347 0 _3027_.CLK
rlabel metal2 6613 333 6627 347 0 _3027_.Q
rlabel metal1 6404 242 6656 258 0 _3022_.gnd
rlabel metal1 6404 2 6656 18 0 _3022_.vdd
rlabel metal2 6553 153 6567 167 0 _3022_.D
rlabel metal2 6513 153 6527 167 0 _3022_.CLK
rlabel metal2 6433 153 6447 167 0 _3022_.Q
rlabel metal1 6284 242 6416 258 0 _2947_.gnd
rlabel metal1 6284 482 6416 498 0 _2947_.vdd
rlabel metal2 6393 333 6407 347 0 _2947_.A
rlabel metal2 6373 353 6387 367 0 _2947_.B
rlabel metal2 6313 333 6327 347 0 _2947_.C
rlabel metal2 6353 333 6367 347 0 _2947_.Y
rlabel metal2 6333 353 6347 367 0 _2947_.D
rlabel metal1 6224 242 6356 258 0 _2927_.gnd
rlabel metal1 6224 2 6356 18 0 _2927_.vdd
rlabel metal2 6333 153 6347 167 0 _2927_.A
rlabel metal2 6313 133 6327 147 0 _2927_.B
rlabel metal2 6253 153 6267 167 0 _2927_.C
rlabel metal2 6293 153 6307 167 0 _2927_.Y
rlabel metal2 6273 133 6287 147 0 _2927_.D
rlabel metal1 6204 242 6296 258 0 _2945_.gnd
rlabel metal1 6204 482 6296 498 0 _2945_.vdd
rlabel metal2 6233 333 6247 347 0 _2945_.B
rlabel metal2 6273 333 6287 347 0 _2945_.A
rlabel metal2 6253 313 6267 327 0 _2945_.Y
rlabel metal1 6344 242 6416 258 0 _2924_.gnd
rlabel metal1 6344 2 6416 18 0 _2924_.vdd
rlabel metal2 6393 173 6407 187 0 _2924_.A
rlabel metal2 6373 133 6387 147 0 _2924_.Y
rlabel nsubstratencontact 6676 488 6676 488 0 FILL100050x3750.vdd
rlabel metal1 6664 242 6696 258 0 FILL100050x3750.gnd
rlabel nsubstratencontact 6684 12 6684 12 0 FILL100050x150.vdd
rlabel metal1 6664 242 6696 258 0 FILL100050x150.gnd
rlabel nsubstratencontact 6656 488 6656 488 0 FILL99750x3750.vdd
rlabel metal1 6644 242 6676 258 0 FILL99750x3750.gnd
rlabel nsubstratencontact 6664 12 6664 12 0 FILL99750x150.vdd
rlabel metal1 6644 242 6676 258 0 FILL99750x150.gnd
rlabel nsubstratencontact 6716 488 6716 488 0 FILL100650x3750.vdd
rlabel metal1 6704 242 6736 258 0 FILL100650x3750.gnd
rlabel nsubstratencontact 6724 12 6724 12 0 FILL100650x150.vdd
rlabel metal1 6704 242 6736 258 0 FILL100650x150.gnd
rlabel nsubstratencontact 6696 488 6696 488 0 FILL100350x3750.vdd
rlabel metal1 6684 242 6716 258 0 FILL100350x3750.gnd
rlabel nsubstratencontact 6704 12 6704 12 0 FILL100350x150.vdd
rlabel metal1 6684 242 6716 258 0 FILL100350x150.gnd
rlabel metal1 4 722 76 738 0 _1654_.gnd
rlabel metal1 4 482 76 498 0 _1654_.vdd
rlabel metal2 13 653 27 667 0 _1654_.A
rlabel metal2 33 613 47 627 0 _1654_.Y
rlabel metal1 244 722 316 738 0 _1467_.gnd
rlabel metal1 244 482 316 498 0 _1467_.vdd
rlabel metal2 253 653 267 667 0 _1467_.A
rlabel metal2 273 613 287 627 0 _1467_.Y
rlabel metal1 64 722 156 738 0 _1657_.gnd
rlabel metal1 64 482 156 498 0 _1657_.vdd
rlabel metal2 73 593 87 607 0 _1657_.A
rlabel metal2 113 593 127 607 0 _1657_.B
rlabel metal2 93 613 107 627 0 _1657_.Y
rlabel metal1 144 722 256 738 0 _1660_.gnd
rlabel metal1 144 482 256 498 0 _1660_.vdd
rlabel metal2 153 613 167 627 0 _1660_.A
rlabel metal2 173 653 187 667 0 _1660_.B
rlabel metal2 193 613 207 627 0 _1660_.C
rlabel metal2 213 633 227 647 0 _1660_.Y
rlabel metal1 504 722 596 738 0 _1472_.gnd
rlabel metal1 504 482 596 498 0 _1472_.vdd
rlabel metal2 573 593 587 607 0 _1472_.A
rlabel metal2 533 593 547 607 0 _1472_.B
rlabel metal2 553 613 567 627 0 _1472_.Y
rlabel metal1 304 722 416 738 0 _1471_.gnd
rlabel metal1 304 482 416 498 0 _1471_.vdd
rlabel metal2 393 613 407 627 0 _1471_.A
rlabel metal2 373 653 387 667 0 _1471_.B
rlabel metal2 353 613 367 627 0 _1471_.C
rlabel metal2 333 633 347 647 0 _1471_.Y
rlabel metal1 404 722 516 738 0 _1470_.gnd
rlabel metal1 404 482 516 498 0 _1470_.vdd
rlabel metal2 413 613 427 627 0 _1470_.A
rlabel metal2 433 593 447 607 0 _1470_.B
rlabel metal2 453 613 467 627 0 _1470_.C
rlabel metal2 473 593 487 607 0 _1470_.Y
rlabel metal1 684 722 756 738 0 _1446_.gnd
rlabel metal1 684 482 756 498 0 _1446_.vdd
rlabel metal2 693 653 707 667 0 _1446_.A
rlabel metal2 713 613 727 627 0 _1446_.Y
rlabel metal1 744 722 816 738 0 _1442_.gnd
rlabel metal1 744 482 816 498 0 _1442_.vdd
rlabel metal2 753 653 767 667 0 _1442_.A
rlabel metal2 773 613 787 627 0 _1442_.Y
rlabel metal1 584 722 696 738 0 _1466_.gnd
rlabel metal1 584 482 696 498 0 _1466_.vdd
rlabel metal2 673 613 687 627 0 _1466_.A
rlabel metal2 653 593 667 607 0 _1466_.B
rlabel metal2 633 613 647 627 0 _1466_.C
rlabel metal2 613 593 627 607 0 _1466_.Y
rlabel metal1 1064 722 1316 738 0 _1481_.gnd
rlabel metal1 1064 482 1316 498 0 _1481_.vdd
rlabel metal2 1153 633 1167 647 0 _1481_.D
rlabel metal2 1193 633 1207 647 0 _1481_.CLK
rlabel metal2 1273 633 1287 647 0 _1481_.Q
rlabel metal1 804 722 896 738 0 _1464_.gnd
rlabel metal1 804 482 896 498 0 _1464_.vdd
rlabel metal2 833 633 847 647 0 _1464_.B
rlabel metal2 873 633 887 647 0 _1464_.A
rlabel metal2 853 653 867 667 0 _1464_.Y
rlabel metal1 884 482 1076 498 0 _1469_.vdd
rlabel metal2 1033 633 1047 647 0 _1469_.A
rlabel metal2 993 613 1007 627 0 _1469_.B
rlabel metal2 973 633 987 647 0 _1469_.C
rlabel metal2 933 613 947 627 0 _1469_.Y
rlabel metal1 884 722 1076 738 0 _1469_.gnd
rlabel metal1 1304 722 1396 738 0 BUFX2_insert40.gnd
rlabel metal1 1304 482 1396 498 0 BUFX2_insert40.vdd
rlabel metal2 1313 633 1327 647 0 BUFX2_insert40.A
rlabel metal2 1353 633 1367 647 0 BUFX2_insert40.Y
rlabel metal1 1464 722 1716 738 0 _1489_.gnd
rlabel metal1 1464 482 1716 498 0 _1489_.vdd
rlabel metal2 1553 633 1567 647 0 _1489_.D
rlabel metal2 1593 633 1607 647 0 _1489_.CLK
rlabel metal2 1673 633 1687 647 0 _1489_.Q
rlabel metal1 1384 722 1476 738 0 _1422_.gnd
rlabel metal1 1384 482 1476 498 0 _1422_.vdd
rlabel metal2 1393 593 1407 607 0 _1422_.A
rlabel metal2 1433 593 1447 607 0 _1422_.B
rlabel metal2 1413 613 1427 627 0 _1422_.Y
rlabel metal1 1704 722 1956 738 0 _1493_.gnd
rlabel metal1 1704 482 1956 498 0 _1493_.vdd
rlabel metal2 1793 633 1807 647 0 _1493_.D
rlabel metal2 1833 633 1847 647 0 _1493_.CLK
rlabel metal2 1913 633 1927 647 0 _1493_.Q
rlabel metal1 1944 722 2196 738 0 _1495_.gnd
rlabel metal1 1944 482 2196 498 0 _1495_.vdd
rlabel metal2 2033 633 2047 647 0 _1495_.D
rlabel metal2 2073 633 2087 647 0 _1495_.CLK
rlabel metal2 2153 633 2167 647 0 _1495_.Q
rlabel metal1 2184 722 2436 738 0 _1491_.gnd
rlabel metal1 2184 482 2436 498 0 _1491_.vdd
rlabel metal2 2273 633 2287 647 0 _1491_.D
rlabel metal2 2313 633 2327 647 0 _1491_.CLK
rlabel metal2 2393 633 2407 647 0 _1491_.Q
rlabel metal1 2424 722 2676 738 0 _2986_.gnd
rlabel metal1 2424 482 2676 498 0 _2986_.vdd
rlabel metal2 2573 633 2587 647 0 _2986_.D
rlabel metal2 2533 633 2547 647 0 _2986_.CLK
rlabel metal2 2453 633 2467 647 0 _2986_.Q
rlabel metal1 2664 722 2796 738 0 _2755_.gnd
rlabel metal1 2664 482 2796 498 0 _2755_.vdd
rlabel metal2 2773 633 2787 647 0 _2755_.A
rlabel metal2 2753 613 2767 627 0 _2755_.B
rlabel metal2 2693 633 2707 647 0 _2755_.C
rlabel metal2 2713 613 2727 627 0 _2755_.D
rlabel metal2 2733 633 2747 647 0 _2755_.Y
rlabel metal1 2784 722 2856 738 0 _2744_.gnd
rlabel metal1 2784 482 2856 498 0 _2744_.vdd
rlabel metal2 2833 653 2847 667 0 _2744_.A
rlabel metal2 2813 613 2827 627 0 _2744_.Y
rlabel metal1 2844 722 2956 738 0 _2748_.gnd
rlabel metal1 2844 482 2956 498 0 _2748_.vdd
rlabel metal2 2933 613 2947 627 0 _2748_.A
rlabel metal2 2913 653 2927 667 0 _2748_.B
rlabel metal2 2893 613 2907 627 0 _2748_.C
rlabel metal2 2873 633 2887 647 0 _2748_.Y
rlabel metal1 3004 722 3116 738 0 _2747_.gnd
rlabel metal1 3004 482 3116 498 0 _2747_.vdd
rlabel metal2 3013 633 3027 647 0 _2747_.A
rlabel metal2 3033 613 3047 627 0 _2747_.B
rlabel metal2 3073 613 3087 627 0 _2747_.C
rlabel metal2 3053 633 3067 647 0 _2747_.Y
rlabel metal1 2944 722 3016 738 0 _2745_.gnd
rlabel metal1 2944 482 3016 498 0 _2745_.vdd
rlabel metal2 2953 653 2967 667 0 _2745_.A
rlabel metal2 2973 613 2987 627 0 _2745_.Y
rlabel metal1 3104 722 3196 738 0 _2746_.gnd
rlabel metal1 3104 482 3196 498 0 _2746_.vdd
rlabel metal2 3113 593 3127 607 0 _2746_.A
rlabel metal2 3153 593 3167 607 0 _2746_.B
rlabel metal2 3133 613 3147 627 0 _2746_.Y
rlabel metal1 3184 722 3296 738 0 _2833_.gnd
rlabel metal1 3184 482 3296 498 0 _2833_.vdd
rlabel metal2 3193 613 3207 627 0 _2833_.A
rlabel metal2 3213 593 3227 607 0 _2833_.B
rlabel metal2 3233 613 3247 627 0 _2833_.C
rlabel metal2 3253 593 3267 607 0 _2833_.Y
rlabel metal1 3344 722 3456 738 0 _2735_.gnd
rlabel metal1 3344 482 3456 498 0 _2735_.vdd
rlabel metal2 3353 633 3367 647 0 _2735_.A
rlabel metal2 3373 613 3387 627 0 _2735_.B
rlabel metal2 3413 613 3427 627 0 _2735_.C
rlabel metal2 3393 633 3407 647 0 _2735_.Y
rlabel metal1 3284 722 3356 738 0 _2733_.gnd
rlabel metal1 3284 482 3356 498 0 _2733_.vdd
rlabel metal2 3293 653 3307 667 0 _2733_.A
rlabel metal2 3313 613 3327 627 0 _2733_.Y
rlabel metal1 3444 722 3536 738 0 _2734_.gnd
rlabel metal1 3444 482 3536 498 0 _2734_.vdd
rlabel metal2 3453 593 3467 607 0 _2734_.A
rlabel metal2 3493 593 3507 607 0 _2734_.B
rlabel metal2 3473 613 3487 627 0 _2734_.Y
rlabel metal1 3704 722 3816 738 0 _2832_.gnd
rlabel metal1 3704 482 3816 498 0 _2832_.vdd
rlabel metal2 3713 633 3727 647 0 _2832_.A
rlabel metal2 3733 613 3747 627 0 _2832_.B
rlabel metal2 3773 613 3787 627 0 _2832_.C
rlabel metal2 3753 633 3767 647 0 _2832_.Y
rlabel metal1 3624 722 3716 738 0 _2830_.gnd
rlabel metal1 3624 482 3716 498 0 _2830_.vdd
rlabel metal2 3673 633 3687 647 0 _2830_.B
rlabel metal2 3633 633 3647 647 0 _2830_.A
rlabel metal2 3653 653 3667 667 0 _2830_.Y
rlabel metal1 3524 722 3636 738 0 _2831_.gnd
rlabel metal1 3524 482 3636 498 0 _2831_.vdd
rlabel metal2 3533 613 3547 627 0 _2831_.A
rlabel metal2 3553 653 3567 667 0 _2831_.B
rlabel metal2 3573 613 3587 627 0 _2831_.C
rlabel metal2 3593 633 3607 647 0 _2831_.Y
rlabel metal1 3904 722 4156 738 0 _3001_.gnd
rlabel metal1 3904 482 4156 498 0 _3001_.vdd
rlabel metal2 4053 633 4067 647 0 _3001_.D
rlabel metal2 4013 633 4027 647 0 _3001_.CLK
rlabel metal2 3933 633 3947 647 0 _3001_.Q
rlabel metal1 3804 722 3916 738 0 _2829_.gnd
rlabel metal1 3804 482 3916 498 0 _2829_.vdd
rlabel metal2 3893 613 3907 627 0 _2829_.A
rlabel metal2 3873 593 3887 607 0 _2829_.B
rlabel metal2 3853 613 3867 627 0 _2829_.C
rlabel metal2 3833 593 3847 607 0 _2829_.Y
rlabel metal1 4224 722 4476 738 0 _2980_.gnd
rlabel metal1 4224 482 4476 498 0 _2980_.vdd
rlabel metal2 4373 633 4387 647 0 _2980_.D
rlabel metal2 4333 633 4347 647 0 _2980_.CLK
rlabel metal2 4253 633 4267 647 0 _2980_.Q
rlabel metal1 4144 722 4236 738 0 _2822_.gnd
rlabel metal1 4144 482 4236 498 0 _2822_.vdd
rlabel metal2 4173 633 4187 647 0 _2822_.B
rlabel metal2 4213 633 4227 647 0 _2822_.A
rlabel metal2 4193 653 4207 667 0 _2822_.Y
rlabel metal1 4464 722 4536 738 0 _2669_.gnd
rlabel metal1 4464 482 4536 498 0 _2669_.vdd
rlabel metal2 4473 653 4487 667 0 _2669_.A
rlabel metal2 4493 613 4507 627 0 _2669_.Y
rlabel metal1 4524 722 4656 738 0 _2683_.gnd
rlabel metal1 4524 482 4656 498 0 _2683_.vdd
rlabel metal2 4533 633 4547 647 0 _2683_.A
rlabel metal2 4553 613 4567 627 0 _2683_.B
rlabel metal2 4613 633 4627 647 0 _2683_.C
rlabel metal2 4593 613 4607 627 0 _2683_.D
rlabel metal2 4573 633 4587 647 0 _2683_.Y
rlabel metal1 4744 722 4856 738 0 _2672_.gnd
rlabel metal1 4744 482 4856 498 0 _2672_.vdd
rlabel metal2 4833 633 4847 647 0 _2672_.A
rlabel metal2 4813 613 4827 627 0 _2672_.B
rlabel metal2 4773 613 4787 627 0 _2672_.C
rlabel metal2 4793 633 4807 647 0 _2672_.Y
rlabel metal1 4644 722 4756 738 0 _2675_.gnd
rlabel metal1 4644 482 4756 498 0 _2675_.vdd
rlabel metal2 4733 613 4747 627 0 _2675_.A
rlabel metal2 4713 653 4727 667 0 _2675_.B
rlabel metal2 4693 613 4707 627 0 _2675_.C
rlabel metal2 4673 633 4687 647 0 _2675_.Y
rlabel metal1 4924 722 4996 738 0 _2670_.gnd
rlabel metal1 4924 482 4996 498 0 _2670_.vdd
rlabel metal2 4973 653 4987 667 0 _2670_.A
rlabel metal2 4953 613 4967 627 0 _2670_.Y
rlabel metal1 4844 722 4936 738 0 _2671_.gnd
rlabel metal1 4844 482 4936 498 0 _2671_.vdd
rlabel metal2 4853 593 4867 607 0 _2671_.A
rlabel metal2 4893 593 4907 607 0 _2671_.B
rlabel metal2 4873 613 4887 627 0 _2671_.Y
rlabel metal1 4984 722 5116 738 0 _2591_.gnd
rlabel metal1 4985 482 5116 498 0 _2591_.vdd
rlabel metal2 5093 613 5107 627 0 _2591_.S
rlabel metal2 5073 633 5087 647 0 _2591_.B
rlabel metal2 5033 613 5047 627 0 _2591_.Y
rlabel metal2 5013 633 5027 647 0 _2591_.A
rlabel metal1 5204 722 5456 738 0 _2996_.gnd
rlabel metal1 5204 482 5456 498 0 _2996_.vdd
rlabel metal2 5353 633 5367 647 0 _2996_.D
rlabel metal2 5313 633 5327 647 0 _2996_.CLK
rlabel metal2 5233 633 5247 647 0 _2996_.Q
rlabel metal1 5104 722 5216 738 0 _2807_.gnd
rlabel metal1 5104 482 5216 498 0 _2807_.vdd
rlabel metal2 5113 613 5127 627 0 _2807_.A
rlabel metal2 5133 593 5147 607 0 _2807_.B
rlabel metal2 5153 613 5167 627 0 _2807_.C
rlabel metal2 5173 593 5187 607 0 _2807_.Y
rlabel metal1 5444 722 5516 738 0 _2773_.gnd
rlabel metal1 5444 482 5516 498 0 _2773_.vdd
rlabel metal2 5453 613 5467 627 0 _2773_.A
rlabel metal2 5473 633 5487 647 0 _2773_.Y
rlabel metal1 5504 722 5636 738 0 _2596_.gnd
rlabel metal1 5504 482 5635 498 0 _2596_.vdd
rlabel metal2 5513 613 5527 627 0 _2596_.S
rlabel metal2 5533 633 5547 647 0 _2596_.B
rlabel metal2 5573 613 5587 627 0 _2596_.Y
rlabel metal2 5593 633 5607 647 0 _2596_.A
rlabel metal1 5704 722 5796 738 0 _2818_.gnd
rlabel metal1 5704 482 5796 498 0 _2818_.vdd
rlabel metal2 5733 633 5747 647 0 _2818_.B
rlabel metal2 5773 633 5787 647 0 _2818_.A
rlabel metal2 5753 653 5767 667 0 _2818_.Y
rlabel metal1 5624 722 5716 738 0 _2814_.gnd
rlabel metal1 5624 482 5716 498 0 _2814_.vdd
rlabel metal2 5653 633 5667 647 0 _2814_.B
rlabel metal2 5693 633 5707 647 0 _2814_.A
rlabel metal2 5673 653 5687 667 0 _2814_.Y
rlabel metal1 5864 722 5956 738 0 _2802_.gnd
rlabel metal1 5864 482 5956 498 0 _2802_.vdd
rlabel metal2 5913 633 5927 647 0 _2802_.B
rlabel metal2 5873 633 5887 647 0 _2802_.A
rlabel metal2 5893 653 5907 667 0 _2802_.Y
rlabel metal1 5784 722 5876 738 0 _2778_.gnd
rlabel metal1 5784 482 5876 498 0 _2778_.vdd
rlabel metal2 5813 633 5827 647 0 _2778_.B
rlabel metal2 5853 633 5867 647 0 _2778_.A
rlabel metal2 5833 653 5847 667 0 _2778_.Y
rlabel metal1 6124 722 6236 738 0 _2804_.gnd
rlabel metal1 6124 482 6236 498 0 _2804_.vdd
rlabel metal2 6133 633 6147 647 0 _2804_.A
rlabel metal2 6153 613 6167 627 0 _2804_.B
rlabel metal2 6193 613 6207 627 0 _2804_.C
rlabel metal2 6173 633 6187 647 0 _2804_.Y
rlabel metal1 6024 722 6136 738 0 _2803_.gnd
rlabel metal1 6024 482 6136 498 0 _2803_.vdd
rlabel metal2 6033 633 6047 647 0 _2803_.A
rlabel metal2 6053 613 6067 627 0 _2803_.B
rlabel metal2 6093 613 6107 627 0 _2803_.C
rlabel metal2 6073 633 6087 647 0 _2803_.Y
rlabel metal1 5944 722 6036 738 0 _2782_.gnd
rlabel metal1 5944 482 6036 498 0 _2782_.vdd
rlabel metal2 5973 633 5987 647 0 _2782_.B
rlabel metal2 6013 633 6027 647 0 _2782_.A
rlabel metal2 5993 653 6007 667 0 _2782_.Y
rlabel metal1 6304 722 6556 738 0 _2995_.gnd
rlabel metal1 6304 482 6556 498 0 _2995_.vdd
rlabel metal2 6393 633 6407 647 0 _2995_.D
rlabel metal2 6433 633 6447 647 0 _2995_.CLK
rlabel metal2 6513 633 6527 647 0 _2995_.Q
rlabel metal1 6224 722 6316 738 0 _2801_.gnd
rlabel metal1 6224 482 6316 498 0 _2801_.vdd
rlabel metal2 6293 593 6307 607 0 _2801_.A
rlabel metal2 6253 593 6267 607 0 _2801_.B
rlabel metal2 6273 613 6287 627 0 _2801_.Y
rlabel nsubstratencontact 6684 492 6684 492 0 FILL100050x7350.vdd
rlabel metal1 6664 722 6696 738 0 FILL100050x7350.gnd
rlabel metal1 6544 722 6616 738 0 _2944_.gnd
rlabel metal1 6544 482 6616 498 0 _2944_.vdd
rlabel metal2 6553 653 6567 667 0 _2944_.A
rlabel metal2 6573 613 6587 627 0 _2944_.Y
rlabel metal1 6604 722 6676 738 0 _2920_.gnd
rlabel metal1 6604 482 6676 498 0 _2920_.vdd
rlabel metal2 6613 653 6627 667 0 _2920_.A
rlabel metal2 6633 613 6647 627 0 _2920_.Y
rlabel nsubstratencontact 6724 492 6724 492 0 FILL100650x7350.vdd
rlabel metal1 6704 722 6736 738 0 FILL100650x7350.gnd
rlabel nsubstratencontact 6704 492 6704 492 0 FILL100350x7350.vdd
rlabel metal1 6684 722 6716 738 0 FILL100350x7350.gnd
rlabel metal1 184 722 436 738 0 _1663_.gnd
rlabel metal1 184 962 436 978 0 _1663_.vdd
rlabel metal2 333 813 347 827 0 _1663_.D
rlabel metal2 293 813 307 827 0 _1663_.CLK
rlabel metal2 213 813 227 827 0 _1663_.Q
rlabel metal1 104 722 196 738 0 _1656_.gnd
rlabel metal1 104 962 196 978 0 _1656_.vdd
rlabel metal2 173 853 187 867 0 _1656_.A
rlabel metal2 133 853 147 867 0 _1656_.B
rlabel metal2 153 833 167 847 0 _1656_.Y
rlabel metal1 4 722 116 738 0 _1561_.gnd
rlabel metal1 4 962 116 978 0 _1561_.vdd
rlabel metal2 13 793 27 807 0 _1561_.A
rlabel metal2 33 813 47 827 0 _1561_.B
rlabel metal2 73 833 87 847 0 _1561_.Y
rlabel metal1 484 722 576 738 0 _1468_.gnd
rlabel metal1 484 962 576 978 0 _1468_.vdd
rlabel metal2 513 813 527 827 0 _1468_.B
rlabel metal2 553 813 567 827 0 _1468_.A
rlabel metal2 533 793 547 807 0 _1468_.Y
rlabel metal1 424 722 496 738 0 _1444_.gnd
rlabel metal1 424 962 496 978 0 _1444_.vdd
rlabel metal2 473 793 487 807 0 _1444_.A
rlabel metal2 453 833 467 847 0 _1444_.Y
rlabel metal1 564 722 656 738 0 _1465_.gnd
rlabel metal1 564 962 656 978 0 _1465_.vdd
rlabel metal2 613 813 627 827 0 _1465_.B
rlabel metal2 573 813 587 827 0 _1465_.A
rlabel metal2 593 793 607 807 0 _1465_.Y
rlabel metal1 644 722 736 738 0 _1445_.gnd
rlabel metal1 644 962 736 978 0 _1445_.vdd
rlabel metal2 653 853 667 867 0 _1445_.A
rlabel metal2 693 853 707 867 0 _1445_.B
rlabel metal2 673 833 687 847 0 _1445_.Y
rlabel metal1 724 722 836 738 0 _1450_.gnd
rlabel metal1 724 962 836 978 0 _1450_.vdd
rlabel metal2 733 833 747 847 0 _1450_.A
rlabel metal2 753 853 767 867 0 _1450_.B
rlabel metal2 773 833 787 847 0 _1450_.C
rlabel metal2 793 853 807 867 0 _1450_.Y
rlabel metal1 824 722 956 738 0 _1451_.gnd
rlabel metal1 824 962 956 978 0 _1451_.vdd
rlabel metal2 833 813 847 827 0 _1451_.A
rlabel metal2 853 833 867 847 0 _1451_.B
rlabel metal2 913 813 927 827 0 _1451_.C
rlabel metal2 873 813 887 827 0 _1451_.Y
rlabel metal2 893 833 907 847 0 _1451_.D
rlabel metal1 1044 722 1156 738 0 _1455_.gnd
rlabel metal1 1044 962 1156 978 0 _1455_.vdd
rlabel metal2 1053 813 1067 827 0 _1455_.A
rlabel metal2 1073 833 1087 847 0 _1455_.B
rlabel metal2 1113 833 1127 847 0 _1455_.C
rlabel metal2 1093 813 1107 827 0 _1455_.Y
rlabel metal1 944 722 1056 738 0 _1454_.gnd
rlabel metal1 944 962 1056 978 0 _1454_.vdd
rlabel metal2 953 813 967 827 0 _1454_.A
rlabel metal2 973 833 987 847 0 _1454_.B
rlabel metal2 1013 833 1027 847 0 _1454_.C
rlabel metal2 993 813 1007 827 0 _1454_.Y
rlabel metal1 1324 722 1436 738 0 _1423_.gnd
rlabel metal1 1324 962 1436 978 0 _1423_.vdd
rlabel metal2 1333 813 1347 827 0 _1423_.A
rlabel metal2 1353 833 1367 847 0 _1423_.B
rlabel metal2 1393 833 1407 847 0 _1423_.C
rlabel metal2 1373 813 1387 827 0 _1423_.Y
rlabel metal1 1144 962 1336 978 0 _1458_.vdd
rlabel metal2 1293 813 1307 827 0 _1458_.A
rlabel metal2 1253 833 1267 847 0 _1458_.B
rlabel metal2 1233 813 1247 827 0 _1458_.C
rlabel metal2 1193 833 1207 847 0 _1458_.Y
rlabel metal1 1144 722 1336 738 0 _1458_.gnd
rlabel metal1 1484 722 1736 738 0 _2968_.gnd
rlabel metal1 1484 962 1736 978 0 _2968_.vdd
rlabel metal2 1573 813 1587 827 0 _2968_.D
rlabel metal2 1613 813 1627 827 0 _2968_.CLK
rlabel metal2 1693 813 1707 827 0 _2968_.Q
rlabel metal1 1424 722 1496 738 0 _1421_.gnd
rlabel metal1 1424 962 1496 978 0 _1421_.vdd
rlabel metal2 1473 793 1487 807 0 _1421_.A
rlabel metal2 1453 833 1467 847 0 _1421_.Y
rlabel metal1 1724 722 1796 738 0 _2569_.gnd
rlabel metal1 1724 962 1796 978 0 _2569_.vdd
rlabel metal2 1733 793 1747 807 0 _2569_.A
rlabel metal2 1753 833 1767 847 0 _2569_.Y
rlabel metal1 1784 722 1916 738 0 _2630_.gnd
rlabel metal1 1784 962 1915 978 0 _2630_.vdd
rlabel metal2 1793 833 1807 847 0 _2630_.S
rlabel metal2 1813 813 1827 827 0 _2630_.B
rlabel metal2 1853 833 1867 847 0 _2630_.Y
rlabel metal2 1873 813 1887 827 0 _2630_.A
rlabel metal1 2084 722 2336 738 0 _3024_.gnd
rlabel metal1 2084 962 2336 978 0 _3024_.vdd
rlabel metal2 2233 813 2247 827 0 _3024_.D
rlabel metal2 2193 813 2207 827 0 _3024_.CLK
rlabel metal2 2113 813 2127 827 0 _3024_.Q
rlabel metal1 1904 722 2016 738 0 _2729_.gnd
rlabel metal1 1904 962 2016 978 0 _2729_.vdd
rlabel metal2 1913 813 1927 827 0 _2729_.A
rlabel metal2 1933 833 1947 847 0 _2729_.B
rlabel metal2 1973 833 1987 847 0 _2729_.C
rlabel metal2 1953 813 1967 827 0 _2729_.Y
rlabel metal1 2004 722 2096 738 0 _2728_.gnd
rlabel metal1 2004 962 2096 978 0 _2728_.vdd
rlabel metal2 2013 853 2027 867 0 _2728_.A
rlabel metal2 2053 853 2067 867 0 _2728_.B
rlabel metal2 2033 833 2047 847 0 _2728_.Y
rlabel metal1 2384 722 2516 738 0 _2935_.gnd
rlabel metal1 2384 962 2516 978 0 _2935_.vdd
rlabel metal2 2393 813 2407 827 0 _2935_.A
rlabel metal2 2413 833 2427 847 0 _2935_.B
rlabel metal2 2473 813 2487 827 0 _2935_.C
rlabel metal2 2433 813 2447 827 0 _2935_.Y
rlabel metal2 2453 833 2467 847 0 _2935_.D
rlabel metal1 2324 722 2396 738 0 _2932_.gnd
rlabel metal1 2324 962 2396 978 0 _2932_.vdd
rlabel metal2 2333 793 2347 807 0 _2932_.A
rlabel metal2 2353 833 2367 847 0 _2932_.Y
rlabel metal1 2584 722 2696 738 0 _2934_.gnd
rlabel metal1 2584 962 2696 978 0 _2934_.vdd
rlabel metal2 2673 813 2687 827 0 _2934_.A
rlabel metal2 2653 833 2667 847 0 _2934_.B
rlabel metal2 2613 833 2627 847 0 _2934_.C
rlabel metal2 2633 813 2647 827 0 _2934_.Y
rlabel metal1 2504 722 2596 738 0 _2933_.gnd
rlabel metal1 2504 962 2596 978 0 _2933_.vdd
rlabel metal2 2553 813 2567 827 0 _2933_.B
rlabel metal2 2513 813 2527 827 0 _2933_.A
rlabel metal2 2533 793 2547 807 0 _2933_.Y
rlabel metal1 2684 722 2896 738 0 CLKBUF1_insert32.gnd
rlabel metal1 2684 962 2896 978 0 CLKBUF1_insert32.vdd
rlabel metal2 2853 833 2867 847 0 CLKBUF1_insert32.A
rlabel metal2 2713 833 2727 847 0 CLKBUF1_insert32.Y
rlabel metal1 2884 722 2996 738 0 _2724_.gnd
rlabel metal1 2884 962 2996 978 0 _2724_.vdd
rlabel metal2 2893 833 2907 847 0 _2724_.A
rlabel metal2 2913 793 2927 807 0 _2724_.B
rlabel metal2 2933 833 2947 847 0 _2724_.C
rlabel metal2 2953 813 2967 827 0 _2724_.Y
rlabel metal1 2984 722 3096 738 0 _2736_.gnd
rlabel metal1 2984 962 3096 978 0 _2736_.vdd
rlabel metal2 3073 833 3087 847 0 _2736_.A
rlabel metal2 3053 793 3067 807 0 _2736_.B
rlabel metal2 3033 833 3047 847 0 _2736_.C
rlabel metal2 3013 813 3027 827 0 _2736_.Y
rlabel metal1 3084 722 3216 738 0 _2649_.gnd
rlabel metal1 3085 962 3216 978 0 _2649_.vdd
rlabel metal2 3193 833 3207 847 0 _2649_.S
rlabel metal2 3173 813 3187 827 0 _2649_.B
rlabel metal2 3133 833 3147 847 0 _2649_.Y
rlabel metal2 3113 813 3127 827 0 _2649_.A
rlabel metal1 3204 722 3336 738 0 _2639_.gnd
rlabel metal1 3205 962 3336 978 0 _2639_.vdd
rlabel metal2 3313 833 3327 847 0 _2639_.S
rlabel metal2 3293 813 3307 827 0 _2639_.B
rlabel metal2 3253 833 3267 847 0 _2639_.Y
rlabel metal2 3233 813 3247 827 0 _2639_.A
rlabel metal1 3324 722 3436 738 0 _2723_.gnd
rlabel metal1 3324 962 3436 978 0 _2723_.vdd
rlabel metal2 3413 813 3427 827 0 _2723_.A
rlabel metal2 3393 833 3407 847 0 _2723_.B
rlabel metal2 3353 833 3367 847 0 _2723_.C
rlabel metal2 3373 813 3387 827 0 _2723_.Y
rlabel metal1 3424 722 3516 738 0 _2722_.gnd
rlabel metal1 3424 962 3516 978 0 _2722_.vdd
rlabel metal2 3433 853 3447 867 0 _2722_.A
rlabel metal2 3473 853 3487 867 0 _2722_.B
rlabel metal2 3453 833 3467 847 0 _2722_.Y
rlabel metal1 3624 722 3696 738 0 _2721_.gnd
rlabel metal1 3624 962 3696 978 0 _2721_.vdd
rlabel metal2 3673 793 3687 807 0 _2721_.A
rlabel metal2 3653 833 3667 847 0 _2721_.Y
rlabel metal1 3504 722 3636 738 0 _2632_.gnd
rlabel metal1 3504 962 3635 978 0 _2632_.vdd
rlabel metal2 3513 833 3527 847 0 _2632_.S
rlabel metal2 3533 813 3547 827 0 _2632_.B
rlabel metal2 3573 833 3587 847 0 _2632_.Y
rlabel metal2 3593 813 3607 827 0 _2632_.A
rlabel metal1 3684 722 3816 738 0 _2631_.gnd
rlabel metal1 3685 962 3816 978 0 _2631_.vdd
rlabel metal2 3793 833 3807 847 0 _2631_.S
rlabel metal2 3773 813 3787 827 0 _2631_.B
rlabel metal2 3733 833 3747 847 0 _2631_.Y
rlabel metal2 3713 813 3727 827 0 _2631_.A
rlabel metal1 3804 722 4056 738 0 _2999_.gnd
rlabel metal1 3804 962 4056 978 0 _2999_.vdd
rlabel metal2 3893 813 3907 827 0 _2999_.D
rlabel metal2 3933 813 3947 827 0 _2999_.CLK
rlabel metal2 4013 813 4027 827 0 _2999_.Q
rlabel metal1 4264 722 4376 738 0 _2824_.gnd
rlabel metal1 4264 962 4376 978 0 _2824_.vdd
rlabel metal2 4273 813 4287 827 0 _2824_.A
rlabel metal2 4293 833 4307 847 0 _2824_.B
rlabel metal2 4333 833 4347 847 0 _2824_.C
rlabel metal2 4313 813 4327 827 0 _2824_.Y
rlabel metal1 4164 722 4276 738 0 _2823_.gnd
rlabel metal1 4164 962 4276 978 0 _2823_.vdd
rlabel metal2 4173 833 4187 847 0 _2823_.A
rlabel metal2 4193 793 4207 807 0 _2823_.B
rlabel metal2 4213 833 4227 847 0 _2823_.C
rlabel metal2 4233 813 4247 827 0 _2823_.Y
rlabel metal1 4044 722 4176 738 0 _2620_.gnd
rlabel metal1 4044 962 4175 978 0 _2620_.vdd
rlabel metal2 4053 833 4067 847 0 _2620_.S
rlabel metal2 4073 813 4087 827 0 _2620_.B
rlabel metal2 4113 833 4127 847 0 _2620_.Y
rlabel metal2 4133 813 4147 827 0 _2620_.A
rlabel metal1 4524 722 4636 738 0 _2711_.gnd
rlabel metal1 4524 962 4636 978 0 _2711_.vdd
rlabel metal2 4533 813 4547 827 0 _2711_.A
rlabel metal2 4553 833 4567 847 0 _2711_.B
rlabel metal2 4593 833 4607 847 0 _2711_.C
rlabel metal2 4573 813 4587 827 0 _2711_.Y
rlabel metal1 4464 722 4536 738 0 _2709_.gnd
rlabel metal1 4464 962 4536 978 0 _2709_.vdd
rlabel metal2 4473 793 4487 807 0 _2709_.A
rlabel metal2 4493 833 4507 847 0 _2709_.Y
rlabel metal1 4364 722 4476 738 0 _2821_.gnd
rlabel metal1 4364 962 4476 978 0 _2821_.vdd
rlabel metal2 4453 833 4467 847 0 _2821_.A
rlabel metal2 4433 853 4447 867 0 _2821_.B
rlabel metal2 4413 833 4427 847 0 _2821_.C
rlabel metal2 4393 853 4407 867 0 _2821_.Y
rlabel metal1 4764 722 4876 738 0 _2681_.gnd
rlabel metal1 4764 962 4876 978 0 _2681_.vdd
rlabel metal2 4773 813 4787 827 0 _2681_.A
rlabel metal2 4793 833 4807 847 0 _2681_.B
rlabel metal2 4833 833 4847 847 0 _2681_.C
rlabel metal2 4813 813 4827 827 0 _2681_.Y
rlabel metal1 4704 722 4776 738 0 _2546_.gnd
rlabel metal1 4704 962 4776 978 0 _2546_.vdd
rlabel metal2 4753 793 4767 807 0 _2546_.A
rlabel metal2 4733 833 4747 847 0 _2546_.Y
rlabel metal1 4624 722 4716 738 0 _2710_.gnd
rlabel metal1 4624 962 4716 978 0 _2710_.vdd
rlabel metal2 4633 853 4647 867 0 _2710_.A
rlabel metal2 4673 853 4687 867 0 _2710_.B
rlabel metal2 4653 833 4667 847 0 _2710_.Y
rlabel metal1 4864 722 4956 738 0 _2680_.gnd
rlabel metal1 4864 962 4956 978 0 _2680_.vdd
rlabel metal2 4873 853 4887 867 0 _2680_.A
rlabel metal2 4913 853 4927 867 0 _2680_.B
rlabel metal2 4893 833 4907 847 0 _2680_.Y
rlabel metal1 4944 722 5076 738 0 _2592_.gnd
rlabel metal1 4944 962 5075 978 0 _2592_.vdd
rlabel metal2 4953 833 4967 847 0 _2592_.S
rlabel metal2 4973 813 4987 827 0 _2592_.B
rlabel metal2 5013 833 5027 847 0 _2592_.Y
rlabel metal2 5033 813 5047 827 0 _2592_.A
rlabel metal1 5064 722 5196 738 0 _2590_.gnd
rlabel metal1 5065 962 5196 978 0 _2590_.vdd
rlabel metal2 5173 833 5187 847 0 _2590_.S
rlabel metal2 5153 813 5167 827 0 _2590_.B
rlabel metal2 5113 833 5127 847 0 _2590_.Y
rlabel metal2 5093 813 5107 827 0 _2590_.A
rlabel metal1 5184 722 5396 738 0 CLKBUF1_insert30.gnd
rlabel metal1 5184 962 5396 978 0 CLKBUF1_insert30.vdd
rlabel metal2 5213 833 5227 847 0 CLKBUF1_insert30.A
rlabel metal2 5353 833 5367 847 0 CLKBUF1_insert30.Y
rlabel metal1 5544 722 5656 738 0 _2687_.gnd
rlabel metal1 5544 962 5656 978 0 _2687_.vdd
rlabel metal2 5553 813 5567 827 0 _2687_.A
rlabel metal2 5573 833 5587 847 0 _2687_.B
rlabel metal2 5613 833 5627 847 0 _2687_.C
rlabel metal2 5593 813 5607 827 0 _2687_.Y
rlabel metal1 5484 722 5556 738 0 _2685_.gnd
rlabel metal1 5484 962 5556 978 0 _2685_.vdd
rlabel metal2 5533 793 5547 807 0 _2685_.A
rlabel metal2 5513 833 5527 847 0 _2685_.Y
rlabel metal1 5384 722 5496 738 0 _2819_.gnd
rlabel metal1 5384 962 5496 978 0 _2819_.vdd
rlabel metal2 5393 833 5407 847 0 _2819_.A
rlabel metal2 5413 793 5427 807 0 _2819_.B
rlabel metal2 5433 833 5447 847 0 _2819_.C
rlabel metal2 5453 813 5467 827 0 _2819_.Y
rlabel metal1 5724 722 5836 738 0 _2820_.gnd
rlabel metal1 5724 962 5836 978 0 _2820_.vdd
rlabel metal2 5733 813 5747 827 0 _2820_.A
rlabel metal2 5753 833 5767 847 0 _2820_.B
rlabel metal2 5793 833 5807 847 0 _2820_.C
rlabel metal2 5773 813 5787 827 0 _2820_.Y
rlabel metal1 5644 722 5736 738 0 _2686_.gnd
rlabel metal1 5644 962 5736 978 0 _2686_.vdd
rlabel metal2 5653 853 5667 867 0 _2686_.A
rlabel metal2 5693 853 5707 867 0 _2686_.B
rlabel metal2 5673 833 5687 847 0 _2686_.Y
rlabel metal1 5824 722 5936 738 0 _2817_.gnd
rlabel metal1 5824 962 5936 978 0 _2817_.vdd
rlabel metal2 5913 833 5927 847 0 _2817_.A
rlabel metal2 5893 853 5907 867 0 _2817_.B
rlabel metal2 5873 833 5887 847 0 _2817_.C
rlabel metal2 5853 853 5867 867 0 _2817_.Y
rlabel metal1 5924 722 6176 738 0 _2998_.gnd
rlabel metal1 5924 962 6176 978 0 _2998_.vdd
rlabel metal2 6013 813 6027 827 0 _2998_.D
rlabel metal2 6053 813 6067 827 0 _2998_.CLK
rlabel metal2 6133 813 6147 827 0 _2998_.Q
rlabel metal1 6264 722 6376 738 0 _2784_.gnd
rlabel metal1 6264 962 6376 978 0 _2784_.vdd
rlabel metal2 6273 813 6287 827 0 _2784_.A
rlabel metal2 6293 833 6307 847 0 _2784_.B
rlabel metal2 6333 833 6347 847 0 _2784_.C
rlabel metal2 6313 813 6327 827 0 _2784_.Y
rlabel metal1 6164 722 6276 738 0 _2783_.gnd
rlabel metal1 6164 962 6276 978 0 _2783_.vdd
rlabel metal2 6173 813 6187 827 0 _2783_.A
rlabel metal2 6193 833 6207 847 0 _2783_.B
rlabel metal2 6233 833 6247 847 0 _2783_.C
rlabel metal2 6213 813 6227 827 0 _2783_.Y
rlabel metal1 6364 722 6456 738 0 _2781_.gnd
rlabel metal1 6364 962 6456 978 0 _2781_.vdd
rlabel metal2 6433 853 6447 867 0 _2781_.A
rlabel metal2 6393 853 6407 867 0 _2781_.B
rlabel metal2 6413 833 6427 847 0 _2781_.Y
rlabel metal1 6444 722 6696 738 0 _2990_.gnd
rlabel metal1 6444 962 6696 978 0 _2990_.vdd
rlabel metal2 6533 813 6547 827 0 _2990_.D
rlabel metal2 6573 813 6587 827 0 _2990_.CLK
rlabel metal2 6653 813 6667 827 0 _2990_.Q
rlabel nsubstratencontact 6716 968 6716 968 0 FILL100650x10950.vdd
rlabel metal1 6704 722 6736 738 0 FILL100650x10950.gnd
rlabel nsubstratencontact 6696 968 6696 968 0 FILL100350x10950.vdd
rlabel metal1 6684 722 6716 738 0 FILL100350x10950.gnd
rlabel metal1 4 1202 256 1218 0 _1628_.gnd
rlabel metal1 4 962 256 978 0 _1628_.vdd
rlabel metal2 153 1113 167 1127 0 _1628_.D
rlabel metal2 113 1113 127 1127 0 _1628_.CLK
rlabel metal2 33 1113 47 1127 0 _1628_.Q
rlabel metal1 244 1202 316 1218 0 _1658_.gnd
rlabel metal1 244 962 316 978 0 _1658_.vdd
rlabel metal2 293 1133 307 1147 0 _1658_.A
rlabel metal2 273 1093 287 1107 0 _1658_.Y
rlabel metal1 304 1202 556 1218 0 _1664_.gnd
rlabel metal1 304 962 556 978 0 _1664_.vdd
rlabel metal2 453 1113 467 1127 0 _1664_.D
rlabel metal2 413 1113 427 1127 0 _1664_.CLK
rlabel metal2 333 1113 347 1127 0 _1664_.Q
rlabel metal1 704 1202 796 1218 0 _1457_.gnd
rlabel metal1 704 962 796 978 0 _1457_.vdd
rlabel metal2 753 1113 767 1127 0 _1457_.B
rlabel metal2 713 1113 727 1127 0 _1457_.A
rlabel metal2 733 1133 747 1147 0 _1457_.Y
rlabel metal1 544 1202 616 1218 0 _1443_.gnd
rlabel metal1 544 962 616 978 0 _1443_.vdd
rlabel metal2 553 1133 567 1147 0 _1443_.A
rlabel metal2 573 1093 587 1107 0 _1443_.Y
rlabel metal1 604 1202 716 1218 0 _1453_.gnd
rlabel metal1 604 962 716 978 0 _1453_.vdd
rlabel metal2 613 1093 627 1107 0 _1453_.A
rlabel metal2 633 1073 647 1087 0 _1453_.B
rlabel metal2 653 1093 667 1107 0 _1453_.C
rlabel metal2 673 1073 687 1087 0 _1453_.Y
rlabel metal1 784 1202 896 1218 0 _1447_.gnd
rlabel metal1 784 962 896 978 0 _1447_.vdd
rlabel metal2 793 1093 807 1107 0 _1447_.A
rlabel metal2 813 1073 827 1087 0 _1447_.B
rlabel metal2 833 1093 847 1107 0 _1447_.C
rlabel metal2 853 1073 867 1087 0 _1447_.Y
rlabel metal1 1024 1202 1276 1218 0 _1483_.gnd
rlabel metal1 1024 962 1276 978 0 _1483_.vdd
rlabel metal2 1113 1113 1127 1127 0 _1483_.D
rlabel metal2 1153 1113 1167 1127 0 _1483_.CLK
rlabel metal2 1233 1113 1247 1127 0 _1483_.Q
rlabel metal1 964 1202 1036 1218 0 _1448_.gnd
rlabel metal1 964 962 1036 978 0 _1448_.vdd
rlabel metal2 973 1133 987 1147 0 _1448_.A
rlabel metal2 993 1093 1007 1107 0 _1448_.Y
rlabel metal1 884 1202 976 1218 0 _1449_.gnd
rlabel metal1 884 962 976 978 0 _1449_.vdd
rlabel metal2 893 1073 907 1087 0 _1449_.A
rlabel metal2 933 1073 947 1087 0 _1449_.B
rlabel metal2 913 1093 927 1107 0 _1449_.Y
rlabel metal1 1264 1202 1476 1218 0 CLKBUF1_insert29.gnd
rlabel metal1 1264 962 1476 978 0 CLKBUF1_insert29.vdd
rlabel metal2 1293 1093 1307 1107 0 CLKBUF1_insert29.A
rlabel metal2 1433 1093 1447 1107 0 CLKBUF1_insert29.Y
rlabel metal1 1464 1202 1716 1218 0 _2969_.gnd
rlabel metal1 1464 962 1716 978 0 _2969_.vdd
rlabel metal2 1553 1113 1567 1127 0 _2969_.D
rlabel metal2 1593 1113 1607 1127 0 _2969_.CLK
rlabel metal2 1673 1113 1687 1127 0 _2969_.Q
rlabel metal1 1784 1202 1916 1218 0 _2572_.gnd
rlabel metal1 1784 962 1916 978 0 _2572_.vdd
rlabel metal2 1893 1113 1907 1127 0 _2572_.A
rlabel metal2 1873 1093 1887 1107 0 _2572_.B
rlabel metal2 1813 1113 1827 1127 0 _2572_.C
rlabel metal2 1853 1113 1867 1127 0 _2572_.Y
rlabel metal2 1833 1093 1847 1107 0 _2572_.D
rlabel metal1 1704 1202 1796 1218 0 _2570_.gnd
rlabel metal1 1704 962 1796 978 0 _2570_.vdd
rlabel metal2 1733 1113 1747 1127 0 _2570_.B
rlabel metal2 1773 1113 1787 1127 0 _2570_.A
rlabel metal2 1753 1133 1767 1147 0 _2570_.Y
rlabel metal1 2004 1202 2116 1218 0 _2579_.gnd
rlabel metal1 2004 962 2116 978 0 _2579_.vdd
rlabel metal2 2093 1113 2107 1127 0 _2579_.A
rlabel metal2 2073 1093 2087 1107 0 _2579_.B
rlabel metal2 2033 1093 2047 1107 0 _2579_.C
rlabel metal2 2053 1113 2067 1127 0 _2579_.Y
rlabel metal1 1904 1202 2016 1218 0 _2571_.gnd
rlabel metal1 1904 962 2016 978 0 _2571_.vdd
rlabel metal2 1993 1113 2007 1127 0 _2571_.A
rlabel metal2 1973 1093 1987 1107 0 _2571_.B
rlabel metal2 1933 1093 1947 1107 0 _2571_.C
rlabel metal2 1953 1113 1967 1127 0 _2571_.Y
rlabel metal1 2104 1202 2196 1218 0 _2578_.gnd
rlabel metal1 2104 962 2196 978 0 _2578_.vdd
rlabel metal2 2133 1113 2147 1127 0 _2578_.B
rlabel metal2 2173 1113 2187 1127 0 _2578_.A
rlabel metal2 2153 1133 2167 1147 0 _2578_.Y
rlabel metal1 2304 1202 2556 1218 0 _2970_.gnd
rlabel metal1 2304 962 2556 978 0 _2970_.vdd
rlabel metal2 2393 1113 2407 1127 0 _2970_.D
rlabel metal2 2433 1113 2447 1127 0 _2970_.CLK
rlabel metal2 2513 1113 2527 1127 0 _2970_.Q
rlabel metal1 2184 1202 2316 1218 0 _2580_.gnd
rlabel metal1 2184 962 2316 978 0 _2580_.vdd
rlabel metal2 2293 1113 2307 1127 0 _2580_.A
rlabel metal2 2273 1093 2287 1107 0 _2580_.B
rlabel metal2 2213 1113 2227 1127 0 _2580_.C
rlabel metal2 2253 1113 2267 1127 0 _2580_.Y
rlabel metal2 2233 1093 2247 1107 0 _2580_.D
rlabel metal1 2604 1202 2716 1218 0 _2753_.gnd
rlabel metal1 2604 962 2716 978 0 _2753_.vdd
rlabel metal2 2613 1113 2627 1127 0 _2753_.A
rlabel metal2 2633 1093 2647 1107 0 _2753_.B
rlabel metal2 2673 1093 2687 1107 0 _2753_.C
rlabel metal2 2653 1113 2667 1127 0 _2753_.Y
rlabel metal1 2544 1202 2616 1218 0 _2577_.gnd
rlabel metal1 2544 962 2616 978 0 _2577_.vdd
rlabel metal2 2593 1133 2607 1147 0 _2577_.A
rlabel metal2 2573 1093 2587 1107 0 _2577_.Y
rlabel metal1 2704 1202 2796 1218 0 BUFX2_insert6.gnd
rlabel metal1 2704 962 2796 978 0 BUFX2_insert6.vdd
rlabel metal2 2773 1113 2787 1127 0 BUFX2_insert6.A
rlabel metal2 2733 1113 2747 1127 0 BUFX2_insert6.Y
rlabel metal1 2784 1202 2856 1218 0 _2720_.gnd
rlabel metal1 2784 962 2856 978 0 _2720_.vdd
rlabel metal2 2793 1133 2807 1147 0 _2720_.A
rlabel metal2 2813 1093 2827 1107 0 _2720_.Y
rlabel metal1 2844 1202 2976 1218 0 _2731_.gnd
rlabel metal1 2844 962 2976 978 0 _2731_.vdd
rlabel metal2 2953 1113 2967 1127 0 _2731_.A
rlabel metal2 2933 1093 2947 1107 0 _2731_.B
rlabel metal2 2873 1113 2887 1127 0 _2731_.C
rlabel metal2 2893 1093 2907 1107 0 _2731_.D
rlabel metal2 2913 1113 2927 1127 0 _2731_.Y
rlabel metal1 2964 1202 3216 1218 0 _2984_.gnd
rlabel metal1 2964 962 3216 978 0 _2984_.vdd
rlabel metal2 3053 1113 3067 1127 0 _2984_.D
rlabel metal2 3093 1113 3107 1127 0 _2984_.CLK
rlabel metal2 3173 1113 3187 1127 0 _2984_.Q
rlabel metal1 3204 1202 3296 1218 0 _2752_.gnd
rlabel metal1 3204 962 3296 978 0 _2752_.vdd
rlabel metal2 3213 1073 3227 1087 0 _2752_.A
rlabel metal2 3253 1073 3267 1087 0 _2752_.B
rlabel metal2 3233 1093 3247 1107 0 _2752_.Y
rlabel metal1 3404 1202 3536 1218 0 _2651_.gnd
rlabel metal1 3404 962 3535 978 0 _2651_.vdd
rlabel metal2 3413 1093 3427 1107 0 _2651_.S
rlabel metal2 3433 1113 3447 1127 0 _2651_.B
rlabel metal2 3473 1093 3487 1107 0 _2651_.Y
rlabel metal2 3493 1113 3507 1127 0 _2651_.A
rlabel metal1 3284 1202 3416 1218 0 _2650_.gnd
rlabel metal1 3285 962 3416 978 0 _2650_.vdd
rlabel metal2 3393 1093 3407 1107 0 _2650_.S
rlabel metal2 3373 1113 3387 1127 0 _2650_.B
rlabel metal2 3333 1093 3347 1107 0 _2650_.Y
rlabel metal2 3313 1113 3327 1127 0 _2650_.A
rlabel metal1 3524 1202 3616 1218 0 BUFX2_insert9.gnd
rlabel metal1 3524 962 3616 978 0 BUFX2_insert9.vdd
rlabel metal2 3593 1113 3607 1127 0 BUFX2_insert9.A
rlabel metal2 3553 1113 3567 1127 0 BUFX2_insert9.Y
rlabel metal1 3604 1202 3856 1218 0 _2967_.gnd
rlabel metal1 3604 962 3856 978 0 _2967_.vdd
rlabel metal2 3693 1113 3707 1127 0 _2967_.D
rlabel metal2 3733 1113 3747 1127 0 _2967_.CLK
rlabel metal2 3813 1113 3827 1127 0 _2967_.Q
rlabel metal1 3964 1202 4096 1218 0 _2622_.gnd
rlabel metal1 3965 962 4096 978 0 _2622_.vdd
rlabel metal2 4073 1093 4087 1107 0 _2622_.S
rlabel metal2 4053 1113 4067 1127 0 _2622_.B
rlabel metal2 4013 1093 4027 1107 0 _2622_.Y
rlabel metal2 3993 1113 4007 1127 0 _2622_.A
rlabel metal1 3844 1202 3976 1218 0 _2621_.gnd
rlabel metal1 3844 962 3975 978 0 _2621_.vdd
rlabel metal2 3853 1093 3867 1107 0 _2621_.S
rlabel metal2 3873 1113 3887 1127 0 _2621_.B
rlabel metal2 3913 1093 3927 1107 0 _2621_.Y
rlabel metal2 3933 1113 3947 1127 0 _2621_.A
rlabel metal1 4144 1202 4276 1218 0 _2931_.gnd
rlabel metal1 4144 962 4276 978 0 _2931_.vdd
rlabel metal2 4153 1113 4167 1127 0 _2931_.A
rlabel metal2 4173 1093 4187 1107 0 _2931_.B
rlabel metal2 4233 1113 4247 1127 0 _2931_.C
rlabel metal2 4193 1113 4207 1127 0 _2931_.Y
rlabel metal2 4213 1093 4227 1107 0 _2931_.D
rlabel metal1 4264 1202 4356 1218 0 _2929_.gnd
rlabel metal1 4264 962 4356 978 0 _2929_.vdd
rlabel metal2 4313 1113 4327 1127 0 _2929_.B
rlabel metal2 4273 1113 4287 1127 0 _2929_.A
rlabel metal2 4293 1133 4307 1147 0 _2929_.Y
rlabel metal1 4084 1202 4156 1218 0 _2928_.gnd
rlabel metal1 4084 962 4156 978 0 _2928_.vdd
rlabel metal2 4093 1133 4107 1147 0 _2928_.A
rlabel metal2 4113 1093 4127 1107 0 _2928_.Y
rlabel metal1 4344 1202 4456 1218 0 _2930_.gnd
rlabel metal1 4344 962 4456 978 0 _2930_.vdd
rlabel metal2 4433 1113 4447 1127 0 _2930_.A
rlabel metal2 4413 1093 4427 1107 0 _2930_.B
rlabel metal2 4373 1093 4387 1107 0 _2930_.C
rlabel metal2 4393 1113 4407 1127 0 _2930_.Y
rlabel metal1 4444 1202 4556 1218 0 _2712_.gnd
rlabel metal1 4444 962 4556 978 0 _2712_.vdd
rlabel metal2 4533 1093 4547 1107 0 _2712_.A
rlabel metal2 4513 1133 4527 1147 0 _2712_.B
rlabel metal2 4493 1093 4507 1107 0 _2712_.C
rlabel metal2 4473 1113 4487 1127 0 _2712_.Y
rlabel metal1 4544 1202 4796 1218 0 _2964_.gnd
rlabel metal1 4544 962 4796 978 0 _2964_.vdd
rlabel metal2 4633 1113 4647 1127 0 _2964_.D
rlabel metal2 4673 1113 4687 1127 0 _2964_.CLK
rlabel metal2 4753 1113 4767 1127 0 _2964_.Q
rlabel metal1 4784 1202 4916 1218 0 _2556_.gnd
rlabel metal1 4784 962 4916 978 0 _2556_.vdd
rlabel metal2 4793 1113 4807 1127 0 _2556_.A
rlabel metal2 4813 1093 4827 1107 0 _2556_.B
rlabel metal2 4873 1113 4887 1127 0 _2556_.C
rlabel metal2 4833 1113 4847 1127 0 _2556_.Y
rlabel metal2 4853 1093 4867 1107 0 _2556_.D
rlabel metal1 4984 1202 5096 1218 0 _2555_.gnd
rlabel metal1 4984 962 5096 978 0 _2555_.vdd
rlabel metal2 5073 1113 5087 1127 0 _2555_.A
rlabel metal2 5053 1093 5067 1107 0 _2555_.B
rlabel metal2 5013 1093 5027 1107 0 _2555_.C
rlabel metal2 5033 1113 5047 1127 0 _2555_.Y
rlabel metal1 4904 1202 4996 1218 0 _2553_.gnd
rlabel metal1 4904 962 4996 978 0 _2553_.vdd
rlabel metal2 4933 1113 4947 1127 0 _2553_.B
rlabel metal2 4973 1113 4987 1127 0 _2553_.A
rlabel metal2 4953 1133 4967 1147 0 _2553_.Y
rlabel metal1 5324 1202 5416 1218 0 BUFX2_insert5.gnd
rlabel metal1 5324 962 5416 978 0 BUFX2_insert5.vdd
rlabel metal2 5393 1113 5407 1127 0 BUFX2_insert5.A
rlabel metal2 5353 1113 5367 1127 0 BUFX2_insert5.Y
rlabel metal1 5084 1202 5176 1218 0 _2917_.gnd
rlabel metal1 5084 962 5176 978 0 _2917_.vdd
rlabel metal2 5113 1113 5127 1127 0 _2917_.B
rlabel metal2 5153 1113 5167 1127 0 _2917_.A
rlabel metal2 5133 1133 5147 1147 0 _2917_.Y
rlabel metal1 5244 1202 5336 1218 0 _2810_.gnd
rlabel metal1 5244 962 5336 978 0 _2810_.vdd
rlabel metal2 5293 1113 5307 1127 0 _2810_.B
rlabel metal2 5253 1113 5267 1127 0 _2810_.A
rlabel metal2 5273 1133 5287 1147 0 _2810_.Y
rlabel metal1 5164 1202 5256 1218 0 _2554_.gnd
rlabel metal1 5164 962 5256 978 0 _2554_.vdd
rlabel metal2 5213 1113 5227 1127 0 _2554_.B
rlabel metal2 5173 1113 5187 1127 0 _2554_.A
rlabel metal2 5193 1133 5207 1147 0 _2554_.Y
rlabel metal1 5484 1202 5576 1218 0 _2809_.gnd
rlabel metal1 5484 962 5576 978 0 _2809_.vdd
rlabel metal2 5533 1113 5547 1127 0 _2809_.B
rlabel metal2 5493 1113 5507 1127 0 _2809_.A
rlabel metal2 5513 1133 5527 1147 0 _2809_.Y
rlabel metal1 5404 1202 5496 1218 0 _2772_.gnd
rlabel metal1 5404 962 5496 978 0 _2772_.vdd
rlabel metal2 5453 1113 5467 1127 0 _2772_.B
rlabel metal2 5413 1113 5427 1127 0 _2772_.A
rlabel metal2 5433 1133 5447 1147 0 _2772_.Y
rlabel metal1 5564 1202 5676 1218 0 _2839_.gnd
rlabel metal1 5564 962 5676 978 0 _2839_.vdd
rlabel metal2 5573 1093 5587 1107 0 _2839_.A
rlabel metal2 5593 1133 5607 1147 0 _2839_.B
rlabel metal2 5613 1093 5627 1107 0 _2839_.C
rlabel metal2 5633 1113 5647 1127 0 _2839_.Y
rlabel metal1 5844 1202 5956 1218 0 _2840_.gnd
rlabel metal1 5844 962 5956 978 0 _2840_.vdd
rlabel metal2 5853 1113 5867 1127 0 _2840_.A
rlabel metal2 5873 1093 5887 1107 0 _2840_.B
rlabel metal2 5913 1093 5927 1107 0 _2840_.C
rlabel metal2 5893 1113 5907 1127 0 _2840_.Y
rlabel metal1 5764 1202 5856 1218 0 _2838_.gnd
rlabel metal1 5764 962 5856 978 0 _2838_.vdd
rlabel metal2 5793 1113 5807 1127 0 _2838_.B
rlabel metal2 5833 1113 5847 1127 0 _2838_.A
rlabel metal2 5813 1133 5827 1147 0 _2838_.Y
rlabel metal1 5664 1202 5776 1218 0 _2805_.gnd
rlabel metal1 5664 962 5776 978 0 _2805_.vdd
rlabel metal2 5673 1133 5687 1147 0 _2805_.A
rlabel metal2 5693 1113 5707 1127 0 _2805_.B
rlabel metal2 5733 1093 5747 1107 0 _2805_.Y
rlabel metal1 6044 1202 6156 1218 0 _2922_.gnd
rlabel metal1 6044 962 6156 978 0 _2922_.vdd
rlabel metal2 6053 1113 6067 1127 0 _2922_.A
rlabel metal2 6073 1093 6087 1107 0 _2922_.B
rlabel metal2 6113 1093 6127 1107 0 _2922_.C
rlabel metal2 6093 1113 6107 1127 0 _2922_.Y
rlabel metal1 5944 1202 6056 1218 0 _2837_.gnd
rlabel metal1 5944 962 6056 978 0 _2837_.vdd
rlabel metal2 6033 1093 6047 1107 0 _2837_.A
rlabel metal2 6013 1073 6027 1087 0 _2837_.B
rlabel metal2 5993 1093 6007 1107 0 _2837_.C
rlabel metal2 5973 1073 5987 1087 0 _2837_.Y
rlabel metal1 6304 1202 6556 1218 0 _3003_.gnd
rlabel metal1 6304 962 6556 978 0 _3003_.vdd
rlabel metal2 6453 1113 6467 1127 0 _3003_.D
rlabel metal2 6413 1113 6427 1127 0 _3003_.CLK
rlabel metal2 6333 1113 6347 1127 0 _3003_.Q
rlabel metal1 6224 1202 6316 1218 0 _2921_.gnd
rlabel metal1 6224 962 6316 978 0 _2921_.vdd
rlabel metal2 6273 1113 6287 1127 0 _2921_.B
rlabel metal2 6233 1113 6247 1127 0 _2921_.A
rlabel metal2 6253 1133 6267 1147 0 _2921_.Y
rlabel metal1 6144 1202 6236 1218 0 _2558_.gnd
rlabel metal1 6144 962 6236 978 0 _2558_.vdd
rlabel metal2 6173 1113 6187 1127 0 _2558_.B
rlabel metal2 6213 1113 6227 1127 0 _2558_.A
rlabel metal2 6193 1133 6207 1147 0 _2558_.Y
rlabel nsubstratencontact 6684 972 6684 972 0 FILL100050x14550.vdd
rlabel metal1 6664 1202 6696 1218 0 FILL100050x14550.gnd
rlabel metal1 6544 1202 6676 1218 0 _2923_.gnd
rlabel metal1 6544 962 6676 978 0 _2923_.vdd
rlabel metal2 6553 1113 6567 1127 0 _2923_.A
rlabel metal2 6573 1093 6587 1107 0 _2923_.B
rlabel metal2 6633 1113 6647 1127 0 _2923_.C
rlabel metal2 6593 1113 6607 1127 0 _2923_.Y
rlabel metal2 6613 1093 6627 1107 0 _2923_.D
rlabel nsubstratencontact 6724 972 6724 972 0 FILL100650x14550.vdd
rlabel metal1 6704 1202 6736 1218 0 FILL100650x14550.gnd
rlabel nsubstratencontact 6704 972 6704 972 0 FILL100350x14550.vdd
rlabel metal1 6684 1202 6716 1218 0 FILL100350x14550.gnd
rlabel metal1 184 1202 296 1218 0 _1662_.gnd
rlabel metal1 184 1442 296 1458 0 _1662_.vdd
rlabel metal2 273 1293 287 1307 0 _1662_.A
rlabel metal2 253 1313 267 1327 0 _1662_.B
rlabel metal2 213 1313 227 1327 0 _1662_.C
rlabel metal2 233 1293 247 1307 0 _1662_.Y
rlabel metal1 104 1202 196 1218 0 _1661_.gnd
rlabel metal1 104 1442 196 1458 0 _1661_.vdd
rlabel metal2 153 1293 167 1307 0 _1661_.B
rlabel metal2 113 1293 127 1307 0 _1661_.A
rlabel metal2 133 1273 147 1287 0 _1661_.Y
rlabel metal1 4 1202 116 1218 0 _1600_.gnd
rlabel metal1 4 1442 116 1458 0 _1600_.vdd
rlabel metal2 13 1293 27 1307 0 _1600_.A
rlabel metal2 73 1293 87 1307 0 _1600_.Y
rlabel metal2 53 1333 67 1347 0 _1600_.B
rlabel metal1 284 1202 376 1218 0 _1659_.gnd
rlabel metal1 284 1442 376 1458 0 _1659_.vdd
rlabel metal2 313 1293 327 1307 0 _1659_.B
rlabel metal2 353 1293 367 1307 0 _1659_.A
rlabel metal2 333 1273 347 1287 0 _1659_.Y
rlabel metal1 364 1202 436 1218 0 _1655_.gnd
rlabel metal1 364 1442 436 1458 0 _1655_.vdd
rlabel metal2 373 1273 387 1287 0 _1655_.A
rlabel metal2 393 1313 407 1327 0 _1655_.Y
rlabel metal1 424 1202 496 1218 0 _1478_.gnd
rlabel metal1 424 1442 496 1458 0 _1478_.vdd
rlabel metal2 433 1273 447 1287 0 _1478_.A
rlabel metal2 453 1313 467 1327 0 _1478_.Y
rlabel metal1 484 1202 576 1218 0 _1479_.gnd
rlabel metal1 484 1442 576 1458 0 _1479_.vdd
rlabel metal2 553 1333 567 1347 0 _1479_.A
rlabel metal2 513 1333 527 1347 0 _1479_.B
rlabel metal2 533 1313 547 1327 0 _1479_.Y
rlabel metal1 664 1202 916 1218 0 _1487_.gnd
rlabel metal1 664 1442 916 1458 0 _1487_.vdd
rlabel metal2 753 1293 767 1307 0 _1487_.D
rlabel metal2 793 1293 807 1307 0 _1487_.CLK
rlabel metal2 873 1293 887 1307 0 _1487_.Q
rlabel metal1 564 1202 676 1218 0 _1480_.gnd
rlabel metal1 564 1442 676 1458 0 _1480_.vdd
rlabel metal2 573 1313 587 1327 0 _1480_.A
rlabel metal2 593 1273 607 1287 0 _1480_.B
rlabel metal2 613 1313 627 1327 0 _1480_.C
rlabel metal2 633 1293 647 1307 0 _1480_.Y
rlabel metal1 904 1202 996 1218 0 _1461_.gnd
rlabel metal1 904 1442 996 1458 0 _1461_.vdd
rlabel metal2 973 1333 987 1347 0 _1461_.A
rlabel metal2 933 1333 947 1347 0 _1461_.B
rlabel metal2 953 1313 967 1327 0 _1461_.Y
rlabel metal1 984 1202 1096 1218 0 _1462_.gnd
rlabel metal1 984 1442 1096 1458 0 _1462_.vdd
rlabel metal2 993 1313 1007 1327 0 _1462_.A
rlabel metal2 1013 1333 1027 1347 0 _1462_.B
rlabel metal2 1033 1313 1047 1327 0 _1462_.C
rlabel metal2 1053 1333 1067 1347 0 _1462_.Y
rlabel metal1 1164 1202 1416 1218 0 _2952_.gnd
rlabel metal1 1164 1442 1416 1458 0 _2952_.vdd
rlabel metal2 1253 1293 1267 1307 0 _2952_.D
rlabel metal2 1293 1293 1307 1307 0 _2952_.CLK
rlabel metal2 1373 1293 1387 1307 0 _2952_.Q
rlabel metal1 1084 1202 1176 1218 0 _1463_.gnd
rlabel metal1 1084 1442 1176 1458 0 _1463_.vdd
rlabel metal2 1133 1293 1147 1307 0 _1463_.B
rlabel metal2 1093 1293 1107 1307 0 _1463_.A
rlabel metal2 1113 1273 1127 1287 0 _1463_.Y
rlabel metal1 1404 1202 1616 1218 0 CLKBUF1_insert25.gnd
rlabel metal1 1404 1442 1616 1458 0 CLKBUF1_insert25.vdd
rlabel metal2 1573 1313 1587 1327 0 CLKBUF1_insert25.A
rlabel metal2 1433 1313 1447 1327 0 CLKBUF1_insert25.Y
rlabel metal1 1804 1202 1936 1218 0 _2576_.gnd
rlabel metal1 1804 1442 1936 1458 0 _2576_.vdd
rlabel metal2 1913 1293 1927 1307 0 _2576_.A
rlabel metal2 1893 1313 1907 1327 0 _2576_.B
rlabel metal2 1833 1293 1847 1307 0 _2576_.C
rlabel metal2 1873 1293 1887 1307 0 _2576_.Y
rlabel metal2 1853 1313 1867 1327 0 _2576_.D
rlabel metal1 1724 1202 1816 1218 0 _2574_.gnd
rlabel metal1 1724 1442 1816 1458 0 _2574_.vdd
rlabel metal2 1753 1293 1767 1307 0 _2574_.B
rlabel metal2 1793 1293 1807 1307 0 _2574_.A
rlabel metal2 1773 1273 1787 1287 0 _2574_.Y
rlabel metal1 1604 1202 1736 1218 0 _2725_.gnd
rlabel metal1 1605 1442 1736 1458 0 _2725_.vdd
rlabel metal2 1713 1313 1727 1327 0 _2725_.S
rlabel metal2 1693 1293 1707 1307 0 _2725_.B
rlabel metal2 1653 1313 1667 1327 0 _2725_.Y
rlabel metal2 1633 1293 1647 1307 0 _2725_.A
rlabel metal1 2084 1202 2196 1218 0 _2741_.gnd
rlabel metal1 2084 1442 2196 1458 0 _2741_.vdd
rlabel metal2 2093 1293 2107 1307 0 _2741_.A
rlabel metal2 2113 1313 2127 1327 0 _2741_.B
rlabel metal2 2153 1313 2167 1327 0 _2741_.C
rlabel metal2 2133 1293 2147 1307 0 _2741_.Y
rlabel metal1 1924 1202 2036 1218 0 _2575_.gnd
rlabel metal1 1924 1442 2036 1458 0 _2575_.vdd
rlabel metal2 2013 1293 2027 1307 0 _2575_.A
rlabel metal2 1993 1313 2007 1327 0 _2575_.B
rlabel metal2 1953 1313 1967 1327 0 _2575_.C
rlabel metal2 1973 1293 1987 1307 0 _2575_.Y
rlabel metal1 2024 1202 2096 1218 0 _2573_.gnd
rlabel metal1 2024 1442 2096 1458 0 _2573_.vdd
rlabel metal2 2033 1273 2047 1287 0 _2573_.A
rlabel metal2 2053 1313 2067 1327 0 _2573_.Y
rlabel metal1 2184 1202 2276 1218 0 _2740_.gnd
rlabel metal1 2184 1442 2276 1458 0 _2740_.vdd
rlabel metal2 2193 1333 2207 1347 0 _2740_.A
rlabel metal2 2233 1333 2247 1347 0 _2740_.B
rlabel metal2 2213 1313 2227 1327 0 _2740_.Y
rlabel metal1 2384 1202 2516 1218 0 _2727_.gnd
rlabel metal1 2385 1442 2516 1458 0 _2727_.vdd
rlabel metal2 2493 1313 2507 1327 0 _2727_.S
rlabel metal2 2473 1293 2487 1307 0 _2727_.B
rlabel metal2 2433 1313 2447 1327 0 _2727_.Y
rlabel metal2 2413 1293 2427 1307 0 _2727_.A
rlabel metal1 2264 1202 2396 1218 0 _2640_.gnd
rlabel metal1 2264 1442 2395 1458 0 _2640_.vdd
rlabel metal2 2273 1313 2287 1327 0 _2640_.S
rlabel metal2 2293 1293 2307 1307 0 _2640_.B
rlabel metal2 2333 1313 2347 1327 0 _2640_.Y
rlabel metal2 2353 1293 2367 1307 0 _2640_.A
rlabel metal1 2624 1202 2756 1218 0 _2754_.gnd
rlabel metal1 2624 1442 2756 1458 0 _2754_.vdd
rlabel metal2 2633 1293 2647 1307 0 _2754_.A
rlabel metal2 2653 1313 2667 1327 0 _2754_.B
rlabel metal2 2713 1293 2727 1307 0 _2754_.C
rlabel metal2 2693 1313 2707 1327 0 _2754_.D
rlabel metal2 2673 1293 2687 1307 0 _2754_.Y
rlabel metal1 2504 1202 2636 1218 0 _2730_.gnd
rlabel metal1 2504 1442 2636 1458 0 _2730_.vdd
rlabel metal2 2613 1293 2627 1307 0 _2730_.A
rlabel metal2 2593 1313 2607 1327 0 _2730_.B
rlabel metal2 2533 1293 2547 1307 0 _2730_.C
rlabel metal2 2553 1313 2567 1327 0 _2730_.D
rlabel metal2 2573 1293 2587 1307 0 _2730_.Y
rlabel metal1 2864 1202 2956 1218 0 BUFX2_insert12.gnd
rlabel metal1 2864 1442 2956 1458 0 BUFX2_insert12.vdd
rlabel metal2 2873 1293 2887 1307 0 BUFX2_insert12.A
rlabel metal2 2913 1293 2927 1307 0 BUFX2_insert12.Y
rlabel metal1 2744 1202 2876 1218 0 _2742_.gnd
rlabel metal1 2744 1442 2876 1458 0 _2742_.vdd
rlabel metal2 2853 1293 2867 1307 0 _2742_.A
rlabel metal2 2833 1313 2847 1327 0 _2742_.B
rlabel metal2 2773 1293 2787 1307 0 _2742_.C
rlabel metal2 2793 1313 2807 1327 0 _2742_.D
rlabel metal2 2813 1293 2827 1307 0 _2742_.Y
rlabel metal1 3064 1202 3136 1218 0 _2732_.gnd
rlabel metal1 3064 1442 3136 1458 0 _2732_.vdd
rlabel metal2 3113 1273 3127 1287 0 _2732_.A
rlabel metal2 3093 1313 3107 1327 0 _2732_.Y
rlabel metal1 2944 1202 3076 1218 0 _2743_.gnd
rlabel metal1 2944 1442 3076 1458 0 _2743_.vdd
rlabel metal2 3053 1293 3067 1307 0 _2743_.A
rlabel metal2 3033 1313 3047 1327 0 _2743_.B
rlabel metal2 2973 1293 2987 1307 0 _2743_.C
rlabel metal2 2993 1313 3007 1327 0 _2743_.D
rlabel metal2 3013 1293 3027 1307 0 _2743_.Y
rlabel metal1 3124 1202 3256 1218 0 _2641_.gnd
rlabel metal1 3125 1442 3256 1458 0 _2641_.vdd
rlabel metal2 3233 1313 3247 1327 0 _2641_.S
rlabel metal2 3213 1293 3227 1307 0 _2641_.B
rlabel metal2 3173 1313 3187 1327 0 _2641_.Y
rlabel metal2 3153 1293 3167 1307 0 _2641_.A
rlabel metal1 3244 1202 3496 1218 0 _2985_.gnd
rlabel metal1 3244 1442 3496 1458 0 _2985_.vdd
rlabel metal2 3333 1293 3347 1307 0 _2985_.D
rlabel metal2 3373 1293 3387 1307 0 _2985_.CLK
rlabel metal2 3453 1293 3467 1307 0 _2985_.Q
rlabel metal1 3564 1202 3696 1218 0 _2568_.gnd
rlabel metal1 3564 1442 3696 1458 0 _2568_.vdd
rlabel metal2 3673 1293 3687 1307 0 _2568_.A
rlabel metal2 3653 1313 3667 1327 0 _2568_.B
rlabel metal2 3593 1293 3607 1307 0 _2568_.C
rlabel metal2 3633 1293 3647 1307 0 _2568_.Y
rlabel metal2 3613 1313 3627 1327 0 _2568_.D
rlabel metal1 3684 1202 3796 1218 0 _2567_.gnd
rlabel metal1 3684 1442 3796 1458 0 _2567_.vdd
rlabel metal2 3773 1293 3787 1307 0 _2567_.A
rlabel metal2 3753 1313 3767 1327 0 _2567_.B
rlabel metal2 3713 1313 3727 1327 0 _2567_.C
rlabel metal2 3733 1293 3747 1307 0 _2567_.Y
rlabel metal1 3484 1202 3576 1218 0 _2566_.gnd
rlabel metal1 3484 1442 3576 1458 0 _2566_.vdd
rlabel metal2 3513 1293 3527 1307 0 _2566_.B
rlabel metal2 3553 1293 3567 1307 0 _2566_.A
rlabel metal2 3533 1273 3547 1287 0 _2566_.Y
rlabel metal1 3844 1202 4096 1218 0 _3023_.gnd
rlabel metal1 3844 1442 4096 1458 0 _3023_.vdd
rlabel metal2 3993 1293 4007 1307 0 _3023_.D
rlabel metal2 3953 1293 3967 1307 0 _3023_.CLK
rlabel metal2 3873 1293 3887 1307 0 _3023_.Q
rlabel metal1 3784 1202 3856 1218 0 _2565_.gnd
rlabel metal1 3784 1442 3856 1458 0 _2565_.vdd
rlabel metal2 3833 1273 3847 1287 0 _2565_.A
rlabel metal2 3813 1313 3827 1327 0 _2565_.Y
rlabel metal1 4084 1202 4336 1218 0 _2983_.gnd
rlabel metal1 4084 1442 4336 1458 0 _2983_.vdd
rlabel metal2 4233 1293 4247 1307 0 _2983_.D
rlabel metal2 4193 1293 4207 1307 0 _2983_.CLK
rlabel metal2 4113 1293 4127 1307 0 _2983_.Q
rlabel metal1 4324 1202 4396 1218 0 _2708_.gnd
rlabel metal1 4324 1442 4396 1458 0 _2708_.vdd
rlabel metal2 4373 1273 4387 1287 0 _2708_.A
rlabel metal2 4353 1313 4367 1327 0 _2708_.Y
rlabel metal1 4384 1202 4516 1218 0 _2719_.gnd
rlabel metal1 4384 1442 4516 1458 0 _2719_.vdd
rlabel metal2 4393 1293 4407 1307 0 _2719_.A
rlabel metal2 4413 1313 4427 1327 0 _2719_.B
rlabel metal2 4473 1293 4487 1307 0 _2719_.C
rlabel metal2 4453 1313 4467 1327 0 _2719_.D
rlabel metal2 4433 1293 4447 1307 0 _2719_.Y
rlabel metal1 4504 1202 4636 1218 0 _2679_.gnd
rlabel metal1 4504 1442 4635 1458 0 _2679_.vdd
rlabel metal2 4513 1313 4527 1327 0 _2679_.S
rlabel metal2 4533 1293 4547 1307 0 _2679_.B
rlabel metal2 4573 1313 4587 1327 0 _2679_.Y
rlabel metal2 4593 1293 4607 1307 0 _2679_.A
rlabel metal1 4744 1202 4836 1218 0 BUFX2_insert10.gnd
rlabel metal1 4744 1442 4836 1458 0 BUFX2_insert10.vdd
rlabel metal2 4813 1293 4827 1307 0 BUFX2_insert10.A
rlabel metal2 4773 1293 4787 1307 0 BUFX2_insert10.Y
rlabel metal1 4624 1202 4756 1218 0 _2682_.gnd
rlabel metal1 4624 1442 4756 1458 0 _2682_.vdd
rlabel metal2 4733 1293 4747 1307 0 _2682_.A
rlabel metal2 4713 1313 4727 1327 0 _2682_.B
rlabel metal2 4653 1293 4667 1307 0 _2682_.C
rlabel metal2 4673 1313 4687 1327 0 _2682_.D
rlabel metal2 4693 1293 4707 1307 0 _2682_.Y
rlabel metal1 4984 1202 5116 1218 0 _2550_.gnd
rlabel metal1 4984 1442 5116 1458 0 _2550_.vdd
rlabel metal2 5093 1293 5107 1307 0 _2550_.A
rlabel metal2 5073 1313 5087 1327 0 _2550_.B
rlabel metal2 5013 1293 5027 1307 0 _2550_.C
rlabel metal2 5053 1293 5067 1307 0 _2550_.Y
rlabel metal2 5033 1313 5047 1327 0 _2550_.D
rlabel metal1 4824 1202 4916 1218 0 _2768_.gnd
rlabel metal1 4824 1442 4916 1458 0 _2768_.vdd
rlabel metal2 4893 1333 4907 1347 0 _2768_.A
rlabel metal2 4853 1333 4867 1347 0 _2768_.B
rlabel metal2 4873 1313 4887 1327 0 _2768_.Y
rlabel metal1 4904 1202 4996 1218 0 _2549_.gnd
rlabel metal1 4904 1442 4996 1458 0 _2549_.vdd
rlabel metal2 4973 1333 4987 1347 0 _2549_.A
rlabel metal2 4933 1333 4947 1347 0 _2549_.B
rlabel metal2 4953 1313 4967 1327 0 _2549_.Y
rlabel metal1 5104 1202 5236 1218 0 _2914_.gnd
rlabel metal1 5104 1442 5236 1458 0 _2914_.vdd
rlabel metal2 5213 1293 5227 1307 0 _2914_.A
rlabel metal2 5193 1313 5207 1327 0 _2914_.B
rlabel metal2 5133 1293 5147 1307 0 _2914_.C
rlabel metal2 5173 1293 5187 1307 0 _2914_.Y
rlabel metal2 5153 1313 5167 1327 0 _2914_.D
rlabel metal1 5284 1202 5376 1218 0 _2548_.gnd
rlabel metal1 5284 1442 5376 1458 0 _2548_.vdd
rlabel metal2 5353 1333 5367 1347 0 _2548_.A
rlabel metal2 5313 1333 5327 1347 0 _2548_.B
rlabel metal2 5333 1313 5347 1327 0 _2548_.Y
rlabel metal1 5224 1202 5296 1218 0 _2676_.gnd
rlabel metal1 5224 1442 5296 1458 0 _2676_.vdd
rlabel metal2 5233 1313 5247 1327 0 _2676_.A
rlabel metal2 5253 1293 5267 1307 0 _2676_.Y
rlabel metal1 5364 1202 5496 1218 0 _2769_.gnd
rlabel metal1 5364 1442 5496 1458 0 _2769_.vdd
rlabel metal2 5373 1293 5387 1307 0 _2769_.A
rlabel metal2 5393 1313 5407 1327 0 _2769_.B
rlabel metal2 5453 1293 5467 1307 0 _2769_.C
rlabel metal2 5413 1293 5427 1307 0 _2769_.Y
rlabel metal2 5433 1313 5447 1327 0 _2769_.D
rlabel metal1 5484 1202 5596 1218 0 _2688_.gnd
rlabel metal1 5484 1442 5596 1458 0 _2688_.vdd
rlabel metal2 5573 1313 5587 1327 0 _2688_.A
rlabel metal2 5553 1273 5567 1287 0 _2688_.B
rlabel metal2 5533 1313 5547 1327 0 _2688_.C
rlabel metal2 5513 1293 5527 1307 0 _2688_.Y
rlabel metal1 5584 1202 5656 1218 0 _2462_.gnd
rlabel metal1 5584 1442 5656 1458 0 _2462_.vdd
rlabel metal2 5593 1313 5607 1327 0 _2462_.A
rlabel metal2 5613 1293 5627 1307 0 _2462_.Y
rlabel metal1 5844 1202 5956 1218 0 _2693_.gnd
rlabel metal1 5844 1442 5956 1458 0 _2693_.vdd
rlabel metal2 5933 1293 5947 1307 0 _2693_.A
rlabel metal2 5913 1313 5927 1327 0 _2693_.B
rlabel metal2 5873 1313 5887 1327 0 _2693_.C
rlabel metal2 5893 1293 5907 1307 0 _2693_.Y
rlabel metal1 5764 1202 5856 1218 0 _2692_.gnd
rlabel metal1 5764 1442 5856 1458 0 _2692_.vdd
rlabel metal2 5833 1333 5847 1347 0 _2692_.A
rlabel metal2 5793 1333 5807 1347 0 _2692_.B
rlabel metal2 5813 1313 5827 1327 0 _2692_.Y
rlabel metal1 5644 1202 5776 1218 0 _2597_.gnd
rlabel metal1 5644 1442 5775 1458 0 _2597_.vdd
rlabel metal2 5653 1313 5667 1327 0 _2597_.S
rlabel metal2 5673 1293 5687 1307 0 _2597_.B
rlabel metal2 5713 1313 5727 1327 0 _2597_.Y
rlabel metal2 5733 1293 5747 1307 0 _2597_.A
rlabel metal1 6104 1202 6236 1218 0 _2560_.gnd
rlabel metal1 6104 1442 6236 1458 0 _2560_.vdd
rlabel metal2 6113 1293 6127 1307 0 _2560_.A
rlabel metal2 6133 1313 6147 1327 0 _2560_.B
rlabel metal2 6193 1293 6207 1307 0 _2560_.C
rlabel metal2 6153 1293 6167 1307 0 _2560_.Y
rlabel metal2 6173 1313 6187 1327 0 _2560_.D
rlabel metal1 6004 1202 6116 1218 0 _2559_.gnd
rlabel metal1 6004 1442 6116 1458 0 _2559_.vdd
rlabel metal2 6013 1293 6027 1307 0 _2559_.A
rlabel metal2 6033 1313 6047 1327 0 _2559_.B
rlabel metal2 6073 1313 6087 1327 0 _2559_.C
rlabel metal2 6053 1293 6067 1307 0 _2559_.Y
rlabel metal1 5944 1202 6016 1218 0 _2557_.gnd
rlabel metal1 5944 1442 6016 1458 0 _2557_.vdd
rlabel metal2 5993 1273 6007 1287 0 _2557_.A
rlabel metal2 5973 1313 5987 1327 0 _2557_.Y
rlabel metal1 6224 1202 6476 1218 0 _2965_.gnd
rlabel metal1 6224 1442 6476 1458 0 _2965_.vdd
rlabel metal2 6373 1293 6387 1307 0 _2965_.D
rlabel metal2 6333 1293 6347 1307 0 _2965_.CLK
rlabel metal2 6253 1293 6267 1307 0 _2965_.Q
rlabel metal1 6464 1202 6716 1218 0 _3021_.gnd
rlabel metal1 6464 1442 6716 1458 0 _3021_.vdd
rlabel metal2 6613 1293 6627 1307 0 _3021_.D
rlabel metal2 6573 1293 6587 1307 0 _3021_.CLK
rlabel metal2 6493 1293 6507 1307 0 _3021_.Q
rlabel nsubstratencontact 6716 1448 6716 1448 0 FILL100650x18150.vdd
rlabel metal1 6704 1202 6736 1218 0 FILL100650x18150.gnd
rlabel metal1 84 1682 296 1698 0 CLKBUF1_insert31.gnd
rlabel metal1 84 1442 296 1458 0 CLKBUF1_insert31.vdd
rlabel metal2 253 1573 267 1587 0 CLKBUF1_insert31.A
rlabel metal2 113 1573 127 1587 0 CLKBUF1_insert31.Y
rlabel metal1 4 1682 96 1698 0 _1599_.gnd
rlabel metal1 4 1442 96 1458 0 _1599_.vdd
rlabel metal2 33 1593 47 1607 0 _1599_.B
rlabel metal2 73 1593 87 1607 0 _1599_.A
rlabel metal2 53 1613 67 1627 0 _1599_.Y
rlabel metal1 284 1682 536 1698 0 _1604_.gnd
rlabel metal1 284 1442 536 1458 0 _1604_.vdd
rlabel metal2 373 1593 387 1607 0 _1604_.D
rlabel metal2 413 1593 427 1607 0 _1604_.CLK
rlabel metal2 493 1593 507 1607 0 _1604_.Q
rlabel metal1 524 1682 596 1698 0 _1456_.gnd
rlabel metal1 524 1442 596 1458 0 _1456_.vdd
rlabel metal2 573 1613 587 1627 0 _1456_.A
rlabel metal2 553 1573 567 1587 0 _1456_.Y
rlabel metal1 784 1682 1036 1698 0 _2960_.gnd
rlabel metal1 784 1442 1036 1458 0 _2960_.vdd
rlabel metal2 873 1593 887 1607 0 _2960_.D
rlabel metal2 913 1593 927 1607 0 _2960_.CLK
rlabel metal2 993 1593 1007 1607 0 _2960_.Q
rlabel metal1 684 1682 796 1698 0 _1460_.gnd
rlabel metal1 684 1442 796 1458 0 _1460_.vdd
rlabel metal2 693 1573 707 1587 0 _1460_.A
rlabel metal2 713 1613 727 1627 0 _1460_.B
rlabel metal2 733 1573 747 1587 0 _1460_.C
rlabel metal2 753 1593 767 1607 0 _1460_.Y
rlabel metal1 584 1682 696 1698 0 _1459_.gnd
rlabel metal1 584 1442 696 1458 0 _1459_.vdd
rlabel metal2 593 1573 607 1587 0 _1459_.A
rlabel metal2 613 1553 627 1567 0 _1459_.B
rlabel metal2 633 1573 647 1587 0 _1459_.C
rlabel metal2 653 1553 667 1567 0 _1459_.Y
rlabel metal1 1024 1682 1096 1698 0 _2492_.gnd
rlabel metal1 1024 1442 1096 1458 0 _2492_.vdd
rlabel metal2 1073 1613 1087 1627 0 _2492_.A
rlabel metal2 1053 1573 1067 1587 0 _2492_.Y
rlabel metal1 1084 1682 1216 1698 0 _2495_.gnd
rlabel metal1 1084 1442 1216 1458 0 _2495_.vdd
rlabel metal2 1093 1593 1107 1607 0 _2495_.A
rlabel metal2 1113 1573 1127 1587 0 _2495_.B
rlabel metal2 1173 1593 1187 1607 0 _2495_.C
rlabel metal2 1133 1593 1147 1607 0 _2495_.Y
rlabel metal2 1153 1573 1167 1587 0 _2495_.D
rlabel metal1 1204 1682 1316 1698 0 _2494_.gnd
rlabel metal1 1204 1442 1316 1458 0 _2494_.vdd
rlabel metal2 1293 1593 1307 1607 0 _2494_.A
rlabel metal2 1273 1573 1287 1587 0 _2494_.B
rlabel metal2 1233 1573 1247 1587 0 _2494_.C
rlabel metal2 1253 1593 1267 1607 0 _2494_.Y
rlabel metal1 1304 1682 1396 1698 0 _2493_.gnd
rlabel metal1 1304 1442 1396 1458 0 _2493_.vdd
rlabel metal2 1333 1593 1347 1607 0 _2493_.B
rlabel metal2 1373 1593 1387 1607 0 _2493_.A
rlabel metal2 1353 1613 1367 1627 0 _2493_.Y
rlabel metal1 1504 1682 1636 1698 0 _2635_.gnd
rlabel metal1 1505 1442 1636 1458 0 _2635_.vdd
rlabel metal2 1613 1573 1627 1587 0 _2635_.S
rlabel metal2 1593 1593 1607 1607 0 _2635_.B
rlabel metal2 1553 1573 1567 1587 0 _2635_.Y
rlabel metal2 1533 1593 1547 1607 0 _2635_.A
rlabel metal1 1384 1682 1516 1698 0 _2634_.gnd
rlabel metal1 1385 1442 1516 1458 0 _2634_.vdd
rlabel metal2 1493 1573 1507 1587 0 _2634_.S
rlabel metal2 1473 1593 1487 1607 0 _2634_.B
rlabel metal2 1433 1573 1447 1587 0 _2634_.Y
rlabel metal2 1413 1593 1427 1607 0 _2634_.A
rlabel metal1 1744 1682 1996 1698 0 _3008_.gnd
rlabel metal1 1744 1442 1996 1458 0 _3008_.vdd
rlabel metal2 1893 1593 1907 1607 0 _3008_.D
rlabel metal2 1853 1593 1867 1607 0 _3008_.CLK
rlabel metal2 1773 1593 1787 1607 0 _3008_.Q
rlabel metal1 1624 1682 1756 1698 0 _2633_.gnd
rlabel metal1 1625 1442 1756 1458 0 _2633_.vdd
rlabel metal2 1733 1573 1747 1587 0 _2633_.S
rlabel metal2 1713 1593 1727 1607 0 _2633_.B
rlabel metal2 1673 1573 1687 1587 0 _2633_.Y
rlabel metal2 1653 1593 1667 1607 0 _2633_.A
rlabel metal1 2104 1682 2176 1698 0 _2862_.gnd
rlabel metal1 2104 1442 2176 1458 0 _2862_.vdd
rlabel metal2 2113 1613 2127 1627 0 _2862_.A
rlabel metal2 2133 1573 2147 1587 0 _2862_.Y
rlabel metal1 1984 1682 2116 1698 0 _2726_.gnd
rlabel metal1 1984 1442 2115 1458 0 _2726_.vdd
rlabel metal2 1993 1573 2007 1587 0 _2726_.S
rlabel metal2 2013 1593 2027 1607 0 _2726_.B
rlabel metal2 2053 1573 2067 1587 0 _2726_.Y
rlabel metal2 2073 1593 2087 1607 0 _2726_.A
rlabel metal1 2164 1682 2296 1698 0 _2865_.gnd
rlabel metal1 2164 1442 2296 1458 0 _2865_.vdd
rlabel metal2 2173 1593 2187 1607 0 _2865_.A
rlabel metal2 2193 1573 2207 1587 0 _2865_.B
rlabel metal2 2253 1593 2267 1607 0 _2865_.C
rlabel metal2 2213 1593 2227 1607 0 _2865_.Y
rlabel metal2 2233 1573 2247 1587 0 _2865_.D
rlabel metal1 2364 1682 2476 1698 0 _2864_.gnd
rlabel metal1 2364 1442 2476 1458 0 _2864_.vdd
rlabel metal2 2453 1593 2467 1607 0 _2864_.A
rlabel metal2 2433 1573 2447 1587 0 _2864_.B
rlabel metal2 2393 1573 2407 1587 0 _2864_.C
rlabel metal2 2413 1593 2427 1607 0 _2864_.Y
rlabel metal1 2284 1682 2376 1698 0 _2863_.gnd
rlabel metal1 2284 1442 2376 1458 0 _2863_.vdd
rlabel metal2 2333 1593 2347 1607 0 _2863_.B
rlabel metal2 2293 1593 2307 1607 0 _2863_.A
rlabel metal2 2313 1613 2327 1627 0 _2863_.Y
rlabel metal1 2464 1682 2556 1698 0 BUFX2_insert16.gnd
rlabel metal1 2464 1442 2556 1458 0 BUFX2_insert16.vdd
rlabel metal2 2533 1593 2547 1607 0 BUFX2_insert16.A
rlabel metal2 2493 1593 2507 1607 0 BUFX2_insert16.Y
rlabel metal1 2544 1682 2636 1698 0 _2551_.gnd
rlabel metal1 2544 1442 2636 1458 0 _2551_.vdd
rlabel metal2 2593 1593 2607 1607 0 _2551_.B
rlabel metal2 2553 1593 2567 1607 0 _2551_.A
rlabel metal2 2573 1613 2587 1627 0 _2551_.Y
rlabel metal1 2624 1682 2716 1698 0 _2915_.gnd
rlabel metal1 2624 1442 2716 1458 0 _2915_.vdd
rlabel metal2 2693 1553 2707 1567 0 _2915_.A
rlabel metal2 2653 1553 2667 1567 0 _2915_.B
rlabel metal2 2673 1573 2687 1587 0 _2915_.Y
rlabel metal1 2704 1682 2796 1698 0 _2552_.gnd
rlabel metal1 2704 1442 2796 1458 0 _2552_.vdd
rlabel metal2 2713 1553 2727 1567 0 _2552_.A
rlabel metal2 2753 1553 2767 1567 0 _2552_.B
rlabel metal2 2733 1573 2747 1587 0 _2552_.Y
rlabel metal1 2904 1682 3016 1698 0 _2806_.gnd
rlabel metal1 2904 1442 3016 1458 0 _2806_.vdd
rlabel metal2 2993 1573 3007 1587 0 _2806_.A
rlabel metal2 2973 1553 2987 1567 0 _2806_.B
rlabel metal2 2953 1573 2967 1587 0 _2806_.C
rlabel metal2 2933 1553 2947 1567 0 _2806_.Y
rlabel metal1 2784 1682 2916 1698 0 _2636_.gnd
rlabel metal1 2785 1442 2916 1458 0 _2636_.vdd
rlabel metal2 2893 1573 2907 1587 0 _2636_.S
rlabel metal2 2873 1593 2887 1607 0 _2636_.B
rlabel metal2 2833 1573 2847 1587 0 _2636_.Y
rlabel metal2 2813 1593 2827 1607 0 _2636_.A
rlabel metal1 3064 1682 3316 1698 0 _2948_.gnd
rlabel metal1 3064 1442 3316 1458 0 _2948_.vdd
rlabel metal2 3153 1593 3167 1607 0 _2948_.D
rlabel metal2 3193 1593 3207 1607 0 _2948_.CLK
rlabel metal2 3273 1593 3287 1607 0 _2948_.Q
rlabel metal1 3004 1682 3076 1698 0 _2466_.gnd
rlabel metal1 3004 1442 3076 1458 0 _2466_.vdd
rlabel metal2 3053 1573 3067 1587 0 _2466_.A
rlabel metal2 3033 1593 3047 1607 0 _2466_.Y
rlabel metal1 3384 1682 3496 1698 0 _2717_.gnd
rlabel metal1 3384 1442 3496 1458 0 _2717_.vdd
rlabel metal2 3473 1593 3487 1607 0 _2717_.A
rlabel metal2 3453 1573 3467 1587 0 _2717_.B
rlabel metal2 3413 1573 3427 1587 0 _2717_.C
rlabel metal2 3433 1593 3447 1607 0 _2717_.Y
rlabel metal1 3304 1682 3396 1698 0 _2716_.gnd
rlabel metal1 3304 1442 3396 1458 0 _2716_.vdd
rlabel metal2 3373 1553 3387 1567 0 _2716_.A
rlabel metal2 3333 1553 3347 1567 0 _2716_.B
rlabel metal2 3353 1573 3367 1587 0 _2716_.Y
rlabel metal1 3604 1682 3716 1698 0 _2849_.gnd
rlabel metal1 3604 1442 3716 1458 0 _2849_.vdd
rlabel metal2 3693 1593 3707 1607 0 _2849_.A
rlabel metal2 3673 1573 3687 1587 0 _2849_.B
rlabel metal2 3633 1573 3647 1587 0 _2849_.C
rlabel metal2 3653 1593 3667 1607 0 _2849_.Y
rlabel metal1 3704 1682 3776 1698 0 _2461_.gnd
rlabel metal1 3704 1442 3776 1458 0 _2461_.vdd
rlabel metal2 3753 1613 3767 1627 0 _2461_.A
rlabel metal2 3733 1573 3747 1587 0 _2461_.Y
rlabel metal1 3484 1682 3616 1698 0 _2718_.gnd
rlabel metal1 3484 1442 3616 1458 0 _2718_.vdd
rlabel metal2 3493 1593 3507 1607 0 _2718_.A
rlabel metal2 3513 1573 3527 1587 0 _2718_.B
rlabel metal2 3573 1593 3587 1607 0 _2718_.C
rlabel metal2 3553 1573 3567 1587 0 _2718_.D
rlabel metal2 3533 1593 3547 1607 0 _2718_.Y
rlabel metal1 3844 1682 3976 1698 0 _2850_.gnd
rlabel metal1 3844 1442 3976 1458 0 _2850_.vdd
rlabel metal2 3953 1593 3967 1607 0 _2850_.A
rlabel metal2 3933 1573 3947 1587 0 _2850_.B
rlabel metal2 3873 1593 3887 1607 0 _2850_.C
rlabel metal2 3913 1593 3927 1607 0 _2850_.Y
rlabel metal2 3893 1573 3907 1587 0 _2850_.D
rlabel metal1 3764 1682 3856 1698 0 _2847_.gnd
rlabel metal1 3764 1442 3856 1458 0 _2847_.vdd
rlabel metal2 3793 1593 3807 1607 0 _2847_.B
rlabel metal2 3833 1593 3847 1607 0 _2847_.A
rlabel metal2 3813 1613 3827 1627 0 _2847_.Y
rlabel metal1 3964 1682 4036 1698 0 _2841_.gnd
rlabel metal1 3964 1442 4036 1458 0 _2841_.vdd
rlabel metal2 4013 1613 4027 1627 0 _2841_.A
rlabel metal2 3993 1573 4007 1587 0 _2841_.Y
rlabel metal1 4024 1682 4276 1698 0 _3004_.gnd
rlabel metal1 4024 1442 4276 1458 0 _3004_.vdd
rlabel metal2 4113 1593 4127 1607 0 _3004_.D
rlabel metal2 4153 1593 4167 1607 0 _3004_.CLK
rlabel metal2 4233 1593 4247 1607 0 _3004_.Q
rlabel metal1 4264 1682 4396 1698 0 _2587_.gnd
rlabel metal1 4265 1442 4396 1458 0 _2587_.vdd
rlabel metal2 4373 1573 4387 1587 0 _2587_.S
rlabel metal2 4353 1593 4367 1607 0 _2587_.B
rlabel metal2 4313 1573 4327 1587 0 _2587_.Y
rlabel metal2 4293 1593 4307 1607 0 _2587_.A
rlabel metal1 4504 1682 4636 1698 0 _2678_.gnd
rlabel metal1 4504 1442 4635 1458 0 _2678_.vdd
rlabel metal2 4513 1573 4527 1587 0 _2678_.S
rlabel metal2 4533 1593 4547 1607 0 _2678_.B
rlabel metal2 4573 1573 4587 1587 0 _2678_.Y
rlabel metal2 4593 1593 4607 1607 0 _2678_.A
rlabel metal1 4384 1682 4516 1698 0 _2677_.gnd
rlabel metal1 4385 1442 4516 1458 0 _2677_.vdd
rlabel metal2 4493 1573 4507 1587 0 _2677_.S
rlabel metal2 4473 1593 4487 1607 0 _2677_.B
rlabel metal2 4433 1573 4447 1587 0 _2677_.Y
rlabel metal2 4413 1593 4427 1607 0 _2677_.A
rlabel metal1 4744 1682 4876 1698 0 _2589_.gnd
rlabel metal1 4744 1442 4875 1458 0 _2589_.vdd
rlabel metal2 4753 1573 4767 1587 0 _2589_.S
rlabel metal2 4773 1593 4787 1607 0 _2589_.B
rlabel metal2 4813 1573 4827 1587 0 _2589_.Y
rlabel metal2 4833 1593 4847 1607 0 _2589_.A
rlabel metal1 4624 1682 4756 1698 0 _2588_.gnd
rlabel metal1 4624 1442 4755 1458 0 _2588_.vdd
rlabel metal2 4633 1573 4647 1587 0 _2588_.S
rlabel metal2 4653 1593 4667 1607 0 _2588_.B
rlabel metal2 4693 1573 4707 1587 0 _2588_.Y
rlabel metal2 4713 1593 4727 1607 0 _2588_.A
rlabel metal1 4984 1682 5236 1698 0 _3012_.gnd
rlabel metal1 4984 1442 5236 1458 0 _3012_.vdd
rlabel metal2 5133 1593 5147 1607 0 _3012_.D
rlabel metal2 5093 1593 5107 1607 0 _3012_.CLK
rlabel metal2 5013 1593 5027 1607 0 _3012_.Q
rlabel metal1 4864 1682 4996 1698 0 _2593_.gnd
rlabel metal1 4864 1442 4995 1458 0 _2593_.vdd
rlabel metal2 4873 1573 4887 1587 0 _2593_.S
rlabel metal2 4893 1593 4907 1607 0 _2593_.B
rlabel metal2 4933 1573 4947 1587 0 _2593_.Y
rlabel metal2 4953 1593 4967 1607 0 _2593_.A
rlabel metal1 5224 1682 5476 1698 0 _2981_.gnd
rlabel metal1 5224 1442 5476 1458 0 _2981_.vdd
rlabel metal2 5373 1593 5387 1607 0 _2981_.D
rlabel metal2 5333 1593 5347 1607 0 _2981_.CLK
rlabel metal2 5253 1593 5267 1607 0 _2981_.Q
rlabel metal1 5464 1682 5596 1698 0 _2695_.gnd
rlabel metal1 5464 1442 5596 1458 0 _2695_.vdd
rlabel metal2 5473 1593 5487 1607 0 _2695_.A
rlabel metal2 5493 1573 5507 1587 0 _2695_.B
rlabel metal2 5553 1593 5567 1607 0 _2695_.C
rlabel metal2 5533 1573 5547 1587 0 _2695_.D
rlabel metal2 5513 1593 5527 1607 0 _2695_.Y
rlabel metal1 5584 1682 5716 1698 0 _2598_.gnd
rlabel metal1 5584 1442 5715 1458 0 _2598_.vdd
rlabel metal2 5593 1573 5607 1587 0 _2598_.S
rlabel metal2 5613 1593 5627 1607 0 _2598_.B
rlabel metal2 5653 1573 5667 1587 0 _2598_.Y
rlabel metal2 5673 1593 5687 1607 0 _2598_.A
rlabel metal1 5704 1682 5816 1698 0 _2563_.gnd
rlabel metal1 5704 1442 5816 1458 0 _2563_.vdd
rlabel metal2 5793 1593 5807 1607 0 _2563_.A
rlabel metal2 5773 1573 5787 1587 0 _2563_.B
rlabel metal2 5733 1573 5747 1587 0 _2563_.C
rlabel metal2 5753 1593 5767 1607 0 _2563_.Y
rlabel metal1 5804 1682 5896 1698 0 _2582_.gnd
rlabel metal1 5804 1442 5896 1458 0 _2582_.vdd
rlabel metal2 5833 1593 5847 1607 0 _2582_.B
rlabel metal2 5873 1593 5887 1607 0 _2582_.A
rlabel metal2 5853 1613 5867 1627 0 _2582_.Y
rlabel metal1 5964 1682 6076 1698 0 _2705_.gnd
rlabel metal1 5964 1442 6076 1458 0 _2705_.vdd
rlabel metal2 6053 1593 6067 1607 0 _2705_.A
rlabel metal2 6033 1573 6047 1587 0 _2705_.B
rlabel metal2 5993 1573 6007 1587 0 _2705_.C
rlabel metal2 6013 1593 6027 1607 0 _2705_.Y
rlabel metal1 6064 1682 6156 1698 0 _2562_.gnd
rlabel metal1 6064 1442 6156 1458 0 _2562_.vdd
rlabel metal2 6093 1593 6107 1607 0 _2562_.B
rlabel metal2 6133 1593 6147 1607 0 _2562_.A
rlabel metal2 6113 1613 6127 1627 0 _2562_.Y
rlabel metal1 5884 1682 5976 1698 0 _2704_.gnd
rlabel metal1 5884 1442 5976 1458 0 _2704_.vdd
rlabel metal2 5953 1553 5967 1567 0 _2704_.A
rlabel metal2 5913 1553 5927 1567 0 _2704_.B
rlabel metal2 5933 1573 5947 1587 0 _2704_.Y
rlabel metal1 6144 1682 6276 1698 0 _2564_.gnd
rlabel metal1 6144 1442 6276 1458 0 _2564_.vdd
rlabel metal2 6253 1593 6267 1607 0 _2564_.A
rlabel metal2 6233 1573 6247 1587 0 _2564_.B
rlabel metal2 6173 1593 6187 1607 0 _2564_.C
rlabel metal2 6213 1593 6227 1607 0 _2564_.Y
rlabel metal2 6193 1573 6207 1587 0 _2564_.D
rlabel metal1 6384 1682 6456 1698 0 _2561_.gnd
rlabel metal1 6384 1442 6456 1458 0 _2561_.vdd
rlabel metal2 6393 1613 6407 1627 0 _2561_.A
rlabel metal2 6413 1573 6427 1587 0 _2561_.Y
rlabel metal1 6264 1682 6396 1698 0 _2611_.gnd
rlabel metal1 6265 1442 6396 1458 0 _2611_.vdd
rlabel metal2 6373 1573 6387 1587 0 _2611_.S
rlabel metal2 6353 1593 6367 1607 0 _2611_.B
rlabel metal2 6313 1573 6327 1587 0 _2611_.Y
rlabel metal2 6293 1593 6307 1607 0 _2611_.A
rlabel metal1 6444 1682 6696 1698 0 _2966_.gnd
rlabel metal1 6444 1442 6696 1458 0 _2966_.vdd
rlabel metal2 6593 1593 6607 1607 0 _2966_.D
rlabel metal2 6553 1593 6567 1607 0 _2966_.CLK
rlabel metal2 6473 1593 6487 1607 0 _2966_.Q
rlabel nsubstratencontact 6724 1452 6724 1452 0 FILL100650x21750.vdd
rlabel metal1 6704 1682 6736 1698 0 FILL100650x21750.gnd
rlabel nsubstratencontact 6704 1452 6704 1452 0 FILL100350x21750.vdd
rlabel metal1 6684 1682 6716 1698 0 FILL100350x21750.gnd
rlabel metal1 64 1682 316 1698 0 _1626_.gnd
rlabel metal1 64 1922 316 1938 0 _1626_.vdd
rlabel metal2 213 1773 227 1787 0 _1626_.D
rlabel metal2 173 1773 187 1787 0 _1626_.CLK
rlabel metal2 93 1773 107 1787 0 _1626_.Q
rlabel metal1 4 1682 76 1698 0 _1560_.gnd
rlabel metal1 4 1922 76 1938 0 _1560_.vdd
rlabel metal2 53 1753 67 1767 0 _1560_.A
rlabel metal2 33 1793 47 1807 0 _1560_.Y
rlabel metal1 524 1682 636 1698 0 _1596_.gnd
rlabel metal1 524 1922 636 1938 0 _1596_.vdd
rlabel metal2 613 1773 627 1787 0 _1596_.A
rlabel metal2 593 1793 607 1807 0 _1596_.B
rlabel metal2 553 1793 567 1807 0 _1596_.C
rlabel metal2 573 1773 587 1787 0 _1596_.Y
rlabel metal1 304 1682 396 1698 0 _1597_.gnd
rlabel metal1 304 1922 396 1938 0 _1597_.vdd
rlabel metal2 353 1773 367 1787 0 _1597_.B
rlabel metal2 313 1773 327 1787 0 _1597_.A
rlabel metal2 333 1753 347 1767 0 _1597_.Y
rlabel metal1 384 1682 476 1698 0 _1508_.gnd
rlabel metal1 384 1922 476 1938 0 _1508_.vdd
rlabel metal2 413 1773 427 1787 0 _1508_.B
rlabel metal2 453 1773 467 1787 0 _1508_.A
rlabel metal2 433 1753 447 1767 0 _1508_.Y
rlabel metal1 464 1682 536 1698 0 _1507_.gnd
rlabel metal1 464 1922 536 1938 0 _1507_.vdd
rlabel metal2 513 1753 527 1767 0 _1507_.A
rlabel metal2 493 1793 507 1807 0 _1507_.Y
rlabel metal1 624 1682 876 1698 0 _1601_.gnd
rlabel metal1 624 1922 876 1938 0 _1601_.vdd
rlabel metal2 773 1773 787 1787 0 _1601_.D
rlabel metal2 733 1773 747 1787 0 _1601_.CLK
rlabel metal2 653 1773 667 1787 0 _1601_.Q
rlabel metal1 1064 1682 1136 1698 0 _1571_.gnd
rlabel metal1 1064 1922 1136 1938 0 _1571_.vdd
rlabel metal2 1073 1753 1087 1767 0 _1571_.A
rlabel metal2 1093 1793 1107 1807 0 _1571_.Y
rlabel metal1 864 1682 976 1698 0 _1595_.gnd
rlabel metal1 864 1922 976 1938 0 _1595_.vdd
rlabel metal2 953 1793 967 1807 0 _1595_.A
rlabel metal2 933 1813 947 1827 0 _1595_.B
rlabel metal2 913 1793 927 1807 0 _1595_.C
rlabel metal2 893 1813 907 1827 0 _1595_.Y
rlabel metal1 964 1682 1076 1698 0 _1504_.gnd
rlabel metal1 964 1922 1076 1938 0 _1504_.vdd
rlabel metal2 973 1773 987 1787 0 _1504_.A
rlabel metal2 1033 1773 1047 1787 0 _1504_.Y
rlabel metal2 1013 1813 1027 1827 0 _1504_.B
rlabel metal1 1124 1682 1236 1698 0 _1572_.gnd
rlabel metal1 1124 1922 1236 1938 0 _1572_.vdd
rlabel metal2 1133 1773 1147 1787 0 _1572_.A
rlabel metal2 1153 1793 1167 1807 0 _1572_.B
rlabel metal2 1193 1793 1207 1807 0 _1572_.C
rlabel metal2 1173 1773 1187 1787 0 _1572_.Y
rlabel metal1 1224 1682 1316 1698 0 _1575_.gnd
rlabel metal1 1224 1922 1316 1938 0 _1575_.vdd
rlabel metal2 1293 1813 1307 1827 0 _1575_.A
rlabel metal2 1253 1813 1267 1827 0 _1575_.B
rlabel metal2 1273 1793 1287 1807 0 _1575_.Y
rlabel metal1 1304 1682 1416 1698 0 _1574_.gnd
rlabel metal1 1304 1922 1416 1938 0 _1574_.vdd
rlabel metal2 1393 1793 1407 1807 0 _1574_.A
rlabel metal2 1373 1813 1387 1827 0 _1574_.B
rlabel metal2 1353 1793 1367 1807 0 _1574_.C
rlabel metal2 1333 1813 1347 1827 0 _1574_.Y
rlabel metal1 1464 1682 1716 1698 0 _1482_.gnd
rlabel metal1 1464 1922 1716 1938 0 _1482_.vdd
rlabel metal2 1553 1773 1567 1787 0 _1482_.D
rlabel metal2 1593 1773 1607 1787 0 _1482_.CLK
rlabel metal2 1673 1773 1687 1787 0 _1482_.Q
rlabel metal1 1404 1682 1476 1698 0 _1573_.gnd
rlabel metal1 1404 1922 1476 1938 0 _1573_.vdd
rlabel metal2 1413 1753 1427 1767 0 _1573_.A
rlabel metal2 1433 1793 1447 1807 0 _1573_.Y
rlabel metal1 1764 1682 1896 1698 0 _2533_.gnd
rlabel metal1 1764 1922 1896 1938 0 _2533_.vdd
rlabel metal2 1773 1773 1787 1787 0 _2533_.A
rlabel metal2 1793 1793 1807 1807 0 _2533_.B
rlabel metal2 1853 1773 1867 1787 0 _2533_.C
rlabel metal2 1813 1773 1827 1787 0 _2533_.Y
rlabel metal2 1833 1793 1847 1807 0 _2533_.D
rlabel metal1 1704 1682 1776 1698 0 _2530_.gnd
rlabel metal1 1704 1922 1776 1938 0 _2530_.vdd
rlabel metal2 1713 1753 1727 1767 0 _2530_.A
rlabel metal2 1733 1793 1747 1807 0 _2530_.Y
rlabel metal1 2064 1682 2316 1698 0 _2953_.gnd
rlabel metal1 2064 1922 2316 1938 0 _2953_.vdd
rlabel metal2 2213 1773 2227 1787 0 _2953_.D
rlabel metal2 2173 1773 2187 1787 0 _2953_.CLK
rlabel metal2 2093 1773 2107 1787 0 _2953_.Q
rlabel metal1 1964 1682 2076 1698 0 _2532_.gnd
rlabel metal1 1964 1922 2076 1938 0 _2532_.vdd
rlabel metal2 1973 1773 1987 1787 0 _2532_.A
rlabel metal2 1993 1793 2007 1807 0 _2532_.B
rlabel metal2 2033 1793 2047 1807 0 _2532_.C
rlabel metal2 2013 1773 2027 1787 0 _2532_.Y
rlabel metal1 1884 1682 1976 1698 0 _2531_.gnd
rlabel metal1 1884 1922 1976 1938 0 _2531_.vdd
rlabel metal2 1933 1773 1947 1787 0 _2531_.B
rlabel metal2 1893 1773 1907 1787 0 _2531_.A
rlabel metal2 1913 1753 1927 1767 0 _2531_.Y
rlabel metal1 2304 1682 2436 1698 0 _2499_.gnd
rlabel metal1 2304 1922 2436 1938 0 _2499_.vdd
rlabel metal2 2413 1773 2427 1787 0 _2499_.A
rlabel metal2 2393 1793 2407 1807 0 _2499_.B
rlabel metal2 2333 1773 2347 1787 0 _2499_.C
rlabel metal2 2373 1773 2387 1787 0 _2499_.Y
rlabel metal2 2353 1793 2367 1807 0 _2499_.D
rlabel metal1 2564 1682 2816 1698 0 _3016_.gnd
rlabel metal1 2564 1922 2816 1938 0 _3016_.vdd
rlabel metal2 2713 1773 2727 1787 0 _3016_.D
rlabel metal2 2673 1773 2687 1787 0 _3016_.CLK
rlabel metal2 2593 1773 2607 1787 0 _3016_.Q
rlabel metal1 2484 1682 2576 1698 0 _2497_.gnd
rlabel metal1 2484 1922 2576 1938 0 _2497_.vdd
rlabel metal2 2533 1773 2547 1787 0 _2497_.B
rlabel metal2 2493 1773 2507 1787 0 _2497_.A
rlabel metal2 2513 1753 2527 1767 0 _2497_.Y
rlabel metal1 2424 1682 2496 1698 0 _2496_.gnd
rlabel metal1 2424 1922 2496 1938 0 _2496_.vdd
rlabel metal2 2433 1753 2447 1767 0 _2496_.A
rlabel metal2 2453 1793 2467 1807 0 _2496_.Y
rlabel metal1 2904 1682 3016 1698 0 _2900_.gnd
rlabel metal1 2904 1922 3016 1938 0 _2900_.vdd
rlabel metal2 2993 1773 3007 1787 0 _2900_.A
rlabel metal2 2973 1793 2987 1807 0 _2900_.B
rlabel metal2 2933 1793 2947 1807 0 _2900_.C
rlabel metal2 2953 1773 2967 1787 0 _2900_.Y
rlabel metal1 2804 1682 2916 1698 0 _2897_.gnd
rlabel metal1 2804 1922 2916 1938 0 _2897_.vdd
rlabel metal2 2813 1793 2827 1807 0 _2897_.A
rlabel metal2 2833 1813 2847 1827 0 _2897_.B
rlabel metal2 2853 1793 2867 1807 0 _2897_.C
rlabel metal2 2873 1813 2887 1827 0 _2897_.Y
rlabel metal1 3004 1682 3096 1698 0 _2898_.gnd
rlabel metal1 3004 1922 3096 1938 0 _2898_.vdd
rlabel metal2 3053 1773 3067 1787 0 _2898_.B
rlabel metal2 3013 1773 3027 1787 0 _2898_.A
rlabel metal2 3033 1753 3047 1767 0 _2898_.Y
rlabel metal1 3084 1682 3196 1698 0 _2903_.gnd
rlabel metal1 3084 1922 3196 1938 0 _2903_.vdd
rlabel metal2 3173 1793 3187 1807 0 _2903_.A
rlabel metal2 3153 1753 3167 1767 0 _2903_.B
rlabel metal2 3133 1793 3147 1807 0 _2903_.C
rlabel metal2 3113 1773 3127 1787 0 _2903_.Y
rlabel metal1 3184 1682 3296 1698 0 _2899_.gnd
rlabel metal1 3184 1922 3296 1938 0 _2899_.vdd
rlabel metal2 3273 1793 3287 1807 0 _2899_.A
rlabel metal2 3253 1753 3267 1767 0 _2899_.B
rlabel metal2 3233 1793 3247 1807 0 _2899_.C
rlabel metal2 3213 1773 3227 1787 0 _2899_.Y
rlabel metal1 3284 1682 3376 1698 0 BUFX2_insert14.gnd
rlabel metal1 3284 1922 3376 1938 0 BUFX2_insert14.vdd
rlabel metal2 3353 1773 3367 1787 0 BUFX2_insert14.A
rlabel metal2 3313 1773 3327 1787 0 BUFX2_insert14.Y
rlabel metal1 3444 1682 3536 1698 0 _2845_.gnd
rlabel metal1 3444 1922 3536 1938 0 _2845_.vdd
rlabel metal2 3493 1773 3507 1787 0 _2845_.B
rlabel metal2 3453 1773 3467 1787 0 _2845_.A
rlabel metal2 3473 1753 3487 1767 0 _2845_.Y
rlabel metal1 3364 1682 3456 1698 0 _2846_.gnd
rlabel metal1 3364 1922 3456 1938 0 _2846_.vdd
rlabel metal2 3433 1813 3447 1827 0 _2846_.A
rlabel metal2 3393 1813 3407 1827 0 _2846_.B
rlabel metal2 3413 1793 3427 1807 0 _2846_.Y
rlabel metal1 3604 1682 3716 1698 0 _2868_.gnd
rlabel metal1 3604 1922 3716 1938 0 _2868_.vdd
rlabel metal2 3613 1773 3627 1787 0 _2868_.A
rlabel metal2 3633 1793 3647 1807 0 _2868_.B
rlabel metal2 3673 1793 3687 1807 0 _2868_.C
rlabel metal2 3653 1773 3667 1787 0 _2868_.Y
rlabel metal1 3524 1682 3616 1698 0 _2878_.gnd
rlabel metal1 3524 1922 3616 1938 0 _2878_.vdd
rlabel metal2 3533 1813 3547 1827 0 _2878_.A
rlabel metal2 3573 1813 3587 1827 0 _2878_.B
rlabel metal2 3553 1793 3567 1807 0 _2878_.Y
rlabel metal1 3704 1682 3796 1698 0 _2475_.gnd
rlabel metal1 3704 1922 3796 1938 0 _2475_.vdd
rlabel metal2 3773 1813 3787 1827 0 _2475_.A
rlabel metal2 3733 1813 3747 1827 0 _2475_.B
rlabel metal2 3753 1793 3767 1807 0 _2475_.Y
rlabel metal1 4004 1682 4136 1698 0 _2479_.gnd
rlabel metal1 4004 1922 4136 1938 0 _2479_.vdd
rlabel metal2 4013 1773 4027 1787 0 _2479_.A
rlabel metal2 4033 1793 4047 1807 0 _2479_.B
rlabel metal2 4093 1773 4107 1787 0 _2479_.C
rlabel metal2 4053 1773 4067 1787 0 _2479_.Y
rlabel metal2 4073 1793 4087 1807 0 _2479_.D
rlabel metal1 3924 1682 4016 1698 0 _2472_.gnd
rlabel metal1 3924 1922 4016 1938 0 _2472_.vdd
rlabel metal2 3973 1773 3987 1787 0 _2472_.B
rlabel metal2 3933 1773 3947 1787 0 _2472_.A
rlabel metal2 3953 1753 3967 1767 0 _2472_.Y
rlabel metal1 3784 1682 3856 1698 0 _2512_.gnd
rlabel metal1 3784 1922 3856 1938 0 _2512_.vdd
rlabel metal2 3833 1753 3847 1767 0 _2512_.A
rlabel metal2 3813 1793 3827 1807 0 _2512_.Y
rlabel metal1 3844 1682 3936 1698 0 _2513_.gnd
rlabel metal1 3844 1922 3936 1938 0 _2513_.vdd
rlabel metal2 3853 1813 3867 1827 0 _2513_.A
rlabel metal2 3893 1813 3907 1827 0 _2513_.B
rlabel metal2 3873 1793 3887 1807 0 _2513_.Y
rlabel metal1 4204 1682 4316 1698 0 _2478_.gnd
rlabel metal1 4204 1922 4316 1938 0 _2478_.vdd
rlabel metal2 4213 1773 4227 1787 0 _2478_.A
rlabel metal2 4233 1793 4247 1807 0 _2478_.B
rlabel metal2 4273 1793 4287 1807 0 _2478_.C
rlabel metal2 4253 1773 4267 1787 0 _2478_.Y
rlabel metal1 4124 1682 4216 1698 0 _2476_.gnd
rlabel metal1 4124 1922 4216 1938 0 _2476_.vdd
rlabel metal2 4153 1773 4167 1787 0 _2476_.B
rlabel metal2 4193 1773 4207 1787 0 _2476_.A
rlabel metal2 4173 1753 4187 1767 0 _2476_.Y
rlabel metal1 4384 1682 4496 1698 0 _2516_.gnd
rlabel metal1 4384 1922 4496 1938 0 _2516_.vdd
rlabel metal2 4393 1773 4407 1787 0 _2516_.A
rlabel metal2 4413 1793 4427 1807 0 _2516_.B
rlabel metal2 4453 1793 4467 1807 0 _2516_.C
rlabel metal2 4433 1773 4447 1787 0 _2516_.Y
rlabel metal1 4484 1682 4576 1698 0 _2514_.gnd
rlabel metal1 4484 1922 4576 1938 0 _2514_.vdd
rlabel metal2 4513 1773 4527 1787 0 _2514_.B
rlabel metal2 4553 1773 4567 1787 0 _2514_.A
rlabel metal2 4533 1753 4547 1767 0 _2514_.Y
rlabel metal1 4304 1682 4396 1698 0 _2471_.gnd
rlabel metal1 4304 1922 4396 1938 0 _2471_.vdd
rlabel metal2 4313 1793 4327 1807 0 _2471_.A
rlabel metal2 4353 1793 4367 1807 0 _2471_.Y
rlabel metal1 4744 1682 4996 1698 0 _2956_.gnd
rlabel metal1 4744 1922 4996 1938 0 _2956_.vdd
rlabel metal2 4893 1773 4907 1787 0 _2956_.D
rlabel metal2 4853 1773 4867 1787 0 _2956_.CLK
rlabel metal2 4773 1773 4787 1787 0 _2956_.Q
rlabel metal1 4564 1682 4696 1698 0 _2517_.gnd
rlabel metal1 4564 1922 4696 1938 0 _2517_.vdd
rlabel metal2 4673 1773 4687 1787 0 _2517_.A
rlabel metal2 4653 1793 4667 1807 0 _2517_.B
rlabel metal2 4593 1773 4607 1787 0 _2517_.C
rlabel metal2 4633 1773 4647 1787 0 _2517_.Y
rlabel metal2 4613 1793 4627 1807 0 _2517_.D
rlabel metal1 4684 1682 4756 1698 0 _2508_.gnd
rlabel metal1 4684 1922 4756 1938 0 _2508_.vdd
rlabel metal2 4733 1753 4747 1767 0 _2508_.A
rlabel metal2 4713 1793 4727 1807 0 _2508_.Y
rlabel metal1 4984 1682 5096 1698 0 _2883_.gnd
rlabel metal1 4984 1922 5096 1938 0 _2883_.vdd
rlabel metal2 4993 1793 5007 1807 0 _2883_.A
rlabel metal2 5013 1753 5027 1767 0 _2883_.B
rlabel metal2 5033 1793 5047 1807 0 _2883_.C
rlabel metal2 5053 1773 5067 1787 0 _2883_.Y
rlabel metal1 5164 1682 5276 1698 0 _2884_.gnd
rlabel metal1 5164 1922 5276 1938 0 _2884_.vdd
rlabel metal2 5173 1773 5187 1787 0 _2884_.A
rlabel metal2 5193 1793 5207 1807 0 _2884_.B
rlabel metal2 5233 1793 5247 1807 0 _2884_.C
rlabel metal2 5213 1773 5227 1787 0 _2884_.Y
rlabel metal1 5084 1682 5176 1698 0 _2880_.gnd
rlabel metal1 5084 1922 5176 1938 0 _2880_.vdd
rlabel metal2 5133 1773 5147 1787 0 _2880_.B
rlabel metal2 5093 1773 5107 1787 0 _2880_.A
rlabel metal2 5113 1753 5127 1767 0 _2880_.Y
rlabel metal1 5264 1682 5376 1698 0 _2879_.gnd
rlabel metal1 5264 1922 5376 1938 0 _2879_.vdd
rlabel metal2 5273 1793 5287 1807 0 _2879_.A
rlabel metal2 5293 1813 5307 1827 0 _2879_.B
rlabel metal2 5313 1793 5327 1807 0 _2879_.C
rlabel metal2 5333 1813 5347 1827 0 _2879_.Y
rlabel metal1 5364 1682 5456 1698 0 BUFX2_insert8.gnd
rlabel metal1 5364 1922 5456 1938 0 BUFX2_insert8.vdd
rlabel metal2 5373 1773 5387 1787 0 BUFX2_insert8.A
rlabel metal2 5413 1773 5427 1787 0 BUFX2_insert8.Y
rlabel metal1 5564 1682 5676 1698 0 _2520_.gnd
rlabel metal1 5564 1922 5676 1938 0 _2520_.vdd
rlabel metal2 5653 1773 5667 1787 0 _2520_.A
rlabel metal2 5633 1793 5647 1807 0 _2520_.B
rlabel metal2 5593 1793 5607 1807 0 _2520_.C
rlabel metal2 5613 1773 5627 1787 0 _2520_.Y
rlabel metal1 5444 1682 5516 1698 0 _2684_.gnd
rlabel metal1 5444 1922 5516 1938 0 _2684_.vdd
rlabel metal2 5493 1753 5507 1767 0 _2684_.A
rlabel metal2 5473 1793 5487 1807 0 _2684_.Y
rlabel metal1 5504 1682 5576 1698 0 _2674_.gnd
rlabel metal1 5504 1922 5576 1938 0 _2674_.vdd
rlabel metal2 5553 1793 5567 1807 0 _2674_.A
rlabel metal2 5533 1773 5547 1787 0 _2674_.Y
rlabel metal1 5864 1682 5956 1698 0 BUFX2_insert15.gnd
rlabel metal1 5864 1922 5956 1938 0 BUFX2_insert15.vdd
rlabel metal2 5873 1773 5887 1787 0 BUFX2_insert15.A
rlabel metal2 5913 1773 5927 1787 0 BUFX2_insert15.Y
rlabel metal1 5664 1682 5756 1698 0 _2673_.gnd
rlabel metal1 5664 1922 5756 1938 0 _2673_.vdd
rlabel metal2 5673 1813 5687 1827 0 _2673_.A
rlabel metal2 5713 1813 5727 1827 0 _2673_.B
rlabel metal2 5693 1793 5707 1807 0 _2673_.Y
rlabel metal1 5744 1682 5876 1698 0 _2694_.gnd
rlabel metal1 5744 1922 5876 1938 0 _2694_.vdd
rlabel metal2 5853 1773 5867 1787 0 _2694_.A
rlabel metal2 5833 1793 5847 1807 0 _2694_.B
rlabel metal2 5773 1773 5787 1787 0 _2694_.C
rlabel metal2 5793 1793 5807 1807 0 _2694_.D
rlabel metal2 5813 1773 5827 1787 0 _2694_.Y
rlabel metal1 6044 1682 6176 1698 0 _2584_.gnd
rlabel metal1 6044 1922 6176 1938 0 _2584_.vdd
rlabel metal2 6153 1773 6167 1787 0 _2584_.A
rlabel metal2 6133 1793 6147 1807 0 _2584_.B
rlabel metal2 6073 1773 6087 1787 0 _2584_.C
rlabel metal2 6113 1773 6127 1787 0 _2584_.Y
rlabel metal2 6093 1793 6107 1807 0 _2584_.D
rlabel metal1 5944 1682 6056 1698 0 _2583_.gnd
rlabel metal1 5944 1922 6056 1938 0 _2583_.vdd
rlabel metal2 6033 1773 6047 1787 0 _2583_.A
rlabel metal2 6013 1793 6027 1807 0 _2583_.B
rlabel metal2 5973 1793 5987 1807 0 _2583_.C
rlabel metal2 5993 1773 6007 1787 0 _2583_.Y
rlabel metal1 6404 1682 6476 1698 0 _2697_.gnd
rlabel metal1 6404 1922 6476 1938 0 _2697_.vdd
rlabel metal2 6413 1753 6427 1767 0 _2697_.A
rlabel metal2 6433 1793 6447 1807 0 _2697_.Y
rlabel metal1 6164 1682 6296 1698 0 _2612_.gnd
rlabel metal1 6164 1922 6295 1938 0 _2612_.vdd
rlabel metal2 6173 1793 6187 1807 0 _2612_.S
rlabel metal2 6193 1773 6207 1787 0 _2612_.B
rlabel metal2 6233 1793 6247 1807 0 _2612_.Y
rlabel metal2 6253 1773 6267 1787 0 _2612_.A
rlabel metal1 6284 1682 6416 1698 0 _2610_.gnd
rlabel metal1 6284 1922 6415 1938 0 _2610_.vdd
rlabel metal2 6293 1793 6307 1807 0 _2610_.S
rlabel metal2 6313 1773 6327 1787 0 _2610_.B
rlabel metal2 6353 1793 6367 1807 0 _2610_.Y
rlabel metal2 6373 1773 6387 1787 0 _2610_.A
rlabel nsubstratencontact 6676 1928 6676 1928 0 FILL100050x25350.vdd
rlabel metal1 6664 1682 6696 1698 0 FILL100050x25350.gnd
rlabel nsubstratencontact 6656 1928 6656 1928 0 FILL99750x25350.vdd
rlabel metal1 6644 1682 6676 1698 0 FILL99750x25350.gnd
rlabel metal1 6464 1682 6576 1698 0 _2699_.gnd
rlabel metal1 6464 1922 6576 1938 0 _2699_.vdd
rlabel metal2 6473 1773 6487 1787 0 _2699_.A
rlabel metal2 6493 1793 6507 1807 0 _2699_.B
rlabel metal2 6533 1793 6547 1807 0 _2699_.C
rlabel metal2 6513 1773 6527 1787 0 _2699_.Y
rlabel metal1 6564 1682 6656 1698 0 _2698_.gnd
rlabel metal1 6564 1922 6656 1938 0 _2698_.vdd
rlabel metal2 6633 1813 6647 1827 0 _2698_.A
rlabel metal2 6593 1813 6607 1827 0 _2698_.B
rlabel metal2 6613 1793 6627 1807 0 _2698_.Y
rlabel nsubstratencontact 6716 1928 6716 1928 0 FILL100650x25350.vdd
rlabel metal1 6704 1682 6736 1698 0 FILL100650x25350.gnd
rlabel nsubstratencontact 6696 1928 6696 1928 0 FILL100350x25350.vdd
rlabel metal1 6684 1682 6716 1698 0 FILL100350x25350.gnd
rlabel metal1 4 2162 96 2178 0 _1598_.gnd
rlabel metal1 4 1922 96 1938 0 _1598_.vdd
rlabel metal2 33 2073 47 2087 0 _1598_.B
rlabel metal2 73 2073 87 2087 0 _1598_.A
rlabel metal2 53 2093 67 2107 0 _1598_.Y
rlabel metal1 84 2162 176 2178 0 _1564_.gnd
rlabel metal1 84 1922 176 1938 0 _1564_.vdd
rlabel metal2 153 2033 167 2047 0 _1564_.A
rlabel metal2 113 2033 127 2047 0 _1564_.B
rlabel metal2 133 2053 147 2067 0 _1564_.Y
rlabel metal1 164 2162 276 2178 0 _1563_.gnd
rlabel metal1 164 1922 276 1938 0 _1563_.vdd
rlabel metal2 253 2053 267 2067 0 _1563_.A
rlabel metal2 233 2033 247 2047 0 _1563_.B
rlabel metal2 213 2053 227 2067 0 _1563_.C
rlabel metal2 193 2033 207 2047 0 _1563_.Y
rlabel metal1 264 2162 376 2178 0 _1562_.gnd
rlabel metal1 264 1922 376 1938 0 _1562_.vdd
rlabel metal2 353 2053 367 2067 0 _1562_.A
rlabel metal2 333 2033 347 2047 0 _1562_.B
rlabel metal2 313 2053 327 2067 0 _1562_.C
rlabel metal2 293 2033 307 2047 0 _1562_.Y
rlabel metal1 364 2162 456 2178 0 _1503_.gnd
rlabel metal1 364 1922 456 1938 0 _1503_.vdd
rlabel metal2 433 2033 447 2047 0 _1503_.A
rlabel metal2 393 2033 407 2047 0 _1503_.B
rlabel metal2 413 2053 427 2067 0 _1503_.Y
rlabel metal1 444 2162 556 2178 0 _1568_.gnd
rlabel metal1 444 1922 556 1938 0 _1568_.vdd
rlabel metal2 453 2053 467 2067 0 _1568_.A
rlabel metal2 473 2033 487 2047 0 _1568_.B
rlabel metal2 493 2053 507 2067 0 _1568_.C
rlabel metal2 513 2033 527 2047 0 _1568_.Y
rlabel metal1 624 2162 736 2178 0 _1565_.gnd
rlabel metal1 624 1922 736 1938 0 _1565_.vdd
rlabel metal2 633 2073 647 2087 0 _1565_.A
rlabel metal2 653 2053 667 2067 0 _1565_.B
rlabel metal2 693 2053 707 2067 0 _1565_.C
rlabel metal2 673 2073 687 2087 0 _1565_.Y
rlabel metal1 544 2162 636 2178 0 _1569_.gnd
rlabel metal1 544 1922 636 1938 0 _1569_.vdd
rlabel metal2 573 2073 587 2087 0 _1569_.B
rlabel metal2 613 2073 627 2087 0 _1569_.A
rlabel metal2 593 2093 607 2107 0 _1569_.Y
rlabel metal1 724 2162 836 2178 0 _1506_.gnd
rlabel metal1 724 1922 836 1938 0 _1506_.vdd
rlabel metal2 733 2053 747 2067 0 _1506_.A
rlabel metal2 753 2033 767 2047 0 _1506_.B
rlabel metal2 773 2053 787 2067 0 _1506_.C
rlabel metal2 793 2033 807 2047 0 _1506_.Y
rlabel metal1 824 2162 916 2178 0 _1505_.gnd
rlabel metal1 824 1922 916 1938 0 _1505_.vdd
rlabel metal2 873 2073 887 2087 0 _1505_.B
rlabel metal2 833 2073 847 2087 0 _1505_.A
rlabel metal2 853 2093 867 2107 0 _1505_.Y
rlabel metal1 904 2162 996 2178 0 _1501_.gnd
rlabel metal1 904 1922 996 1938 0 _1501_.vdd
rlabel metal2 973 2033 987 2047 0 _1501_.A
rlabel metal2 933 2033 947 2047 0 _1501_.B
rlabel metal2 953 2053 967 2067 0 _1501_.Y
rlabel metal1 984 2162 1116 2178 0 _1570_.gnd
rlabel metal1 984 1922 1115 1938 0 _1570_.vdd
rlabel metal2 993 2053 1007 2067 0 _1570_.S
rlabel metal2 1013 2073 1027 2087 0 _1570_.B
rlabel metal2 1053 2053 1067 2067 0 _1570_.Y
rlabel metal2 1073 2073 1087 2087 0 _1570_.A
rlabel metal1 1104 2162 1356 2178 0 _2961_.gnd
rlabel metal1 1104 1922 1356 1938 0 _2961_.vdd
rlabel metal2 1193 2073 1207 2087 0 _2961_.D
rlabel metal2 1233 2073 1247 2087 0 _2961_.CLK
rlabel metal2 1313 2073 1327 2087 0 _2961_.Q
rlabel metal1 1404 2162 1536 2178 0 _2537_.gnd
rlabel metal1 1404 1922 1536 1938 0 _2537_.vdd
rlabel metal2 1413 2073 1427 2087 0 _2537_.A
rlabel metal2 1433 2053 1447 2067 0 _2537_.B
rlabel metal2 1493 2073 1507 2087 0 _2537_.C
rlabel metal2 1453 2073 1467 2087 0 _2537_.Y
rlabel metal2 1473 2053 1487 2067 0 _2537_.D
rlabel metal1 1524 2162 1636 2178 0 _2536_.gnd
rlabel metal1 1524 1922 1636 1938 0 _2536_.vdd
rlabel metal2 1613 2073 1627 2087 0 _2536_.A
rlabel metal2 1593 2053 1607 2067 0 _2536_.B
rlabel metal2 1553 2053 1567 2067 0 _2536_.C
rlabel metal2 1573 2073 1587 2087 0 _2536_.Y
rlabel metal1 1344 2162 1416 2178 0 _2534_.gnd
rlabel metal1 1344 1922 1416 1938 0 _2534_.vdd
rlabel metal2 1353 2093 1367 2107 0 _2534_.A
rlabel metal2 1373 2053 1387 2067 0 _2534_.Y
rlabel metal1 1624 2162 1736 2178 0 _2540_.gnd
rlabel metal1 1624 1922 1736 1938 0 _2540_.vdd
rlabel metal2 1713 2073 1727 2087 0 _2540_.A
rlabel metal2 1693 2053 1707 2067 0 _2540_.B
rlabel metal2 1653 2053 1667 2067 0 _2540_.C
rlabel metal2 1673 2073 1687 2087 0 _2540_.Y
rlabel metal1 1804 2162 1916 2178 0 _2498_.gnd
rlabel metal1 1804 1922 1916 1938 0 _2498_.vdd
rlabel metal2 1893 2073 1907 2087 0 _2498_.A
rlabel metal2 1873 2053 1887 2067 0 _2498_.B
rlabel metal2 1833 2053 1847 2067 0 _2498_.C
rlabel metal2 1853 2073 1867 2087 0 _2498_.Y
rlabel metal1 1724 2162 1816 2178 0 _2535_.gnd
rlabel metal1 1724 1922 1816 1938 0 _2535_.vdd
rlabel metal2 1753 2073 1767 2087 0 _2535_.B
rlabel metal2 1793 2073 1807 2087 0 _2535_.A
rlabel metal2 1773 2093 1787 2107 0 _2535_.Y
rlabel metal1 2024 2162 2156 2178 0 _2737_.gnd
rlabel metal1 2025 1922 2156 1938 0 _2737_.vdd
rlabel metal2 2133 2053 2147 2067 0 _2737_.S
rlabel metal2 2113 2073 2127 2087 0 _2737_.B
rlabel metal2 2073 2053 2087 2067 0 _2737_.Y
rlabel metal2 2053 2073 2067 2087 0 _2737_.A
rlabel metal1 1904 2162 2036 2178 0 _2643_.gnd
rlabel metal1 1905 1922 2036 1938 0 _2643_.vdd
rlabel metal2 2013 2053 2027 2067 0 _2643_.S
rlabel metal2 1993 2073 2007 2087 0 _2643_.B
rlabel metal2 1953 2053 1967 2067 0 _2643_.Y
rlabel metal2 1933 2073 1947 2087 0 _2643_.A
rlabel metal1 2144 2162 2396 2178 0 _3017_.gnd
rlabel metal1 2144 1922 2396 1938 0 _3017_.vdd
rlabel metal2 2233 2073 2247 2087 0 _3017_.D
rlabel metal2 2273 2073 2287 2087 0 _3017_.CLK
rlabel metal2 2353 2073 2367 2087 0 _3017_.Q
rlabel metal1 2384 2162 2496 2178 0 _2904_.gnd
rlabel metal1 2384 1922 2496 1938 0 _2904_.vdd
rlabel metal2 2473 2073 2487 2087 0 _2904_.A
rlabel metal2 2453 2053 2467 2067 0 _2904_.B
rlabel metal2 2413 2053 2427 2067 0 _2904_.C
rlabel metal2 2433 2073 2447 2087 0 _2904_.Y
rlabel metal1 2484 2162 2576 2178 0 _2902_.gnd
rlabel metal1 2484 1922 2576 1938 0 _2902_.vdd
rlabel metal2 2533 2073 2547 2087 0 _2902_.B
rlabel metal2 2493 2073 2507 2087 0 _2902_.A
rlabel metal2 2513 2093 2527 2107 0 _2902_.Y
rlabel metal1 2564 2162 2676 2178 0 _2901_.gnd
rlabel metal1 2564 1922 2676 1938 0 _2901_.vdd
rlabel metal2 2653 2053 2667 2067 0 _2901_.A
rlabel metal2 2633 2033 2647 2047 0 _2901_.B
rlabel metal2 2613 2053 2627 2067 0 _2901_.C
rlabel metal2 2593 2033 2607 2047 0 _2901_.Y
rlabel metal1 2664 2162 2796 2178 0 _2739_.gnd
rlabel metal1 2664 1922 2795 1938 0 _2739_.vdd
rlabel metal2 2673 2053 2687 2067 0 _2739_.S
rlabel metal2 2693 2073 2707 2087 0 _2739_.B
rlabel metal2 2733 2053 2747 2067 0 _2739_.Y
rlabel metal2 2753 2073 2767 2087 0 _2739_.A
rlabel metal1 2904 2162 2976 2178 0 _2642_.gnd
rlabel metal1 2904 1922 2976 1938 0 _2642_.vdd
rlabel metal2 2913 2093 2927 2107 0 _2642_.A
rlabel metal2 2933 2053 2947 2067 0 _2642_.Y
rlabel metal1 2784 2162 2916 2178 0 _2738_.gnd
rlabel metal1 2785 1922 2916 1938 0 _2738_.vdd
rlabel metal2 2893 2053 2907 2067 0 _2738_.S
rlabel metal2 2873 2073 2887 2087 0 _2738_.B
rlabel metal2 2833 2053 2847 2067 0 _2738_.Y
rlabel metal2 2813 2073 2827 2087 0 _2738_.A
rlabel metal1 2964 2162 3096 2178 0 _2644_.gnd
rlabel metal1 2964 1922 3096 1938 0 _2644_.vdd
rlabel metal2 2973 2073 2987 2087 0 _2644_.A
rlabel metal2 2993 2053 3007 2067 0 _2644_.B
rlabel metal2 3053 2073 3067 2087 0 _2644_.C
rlabel metal2 3013 2073 3027 2087 0 _2644_.Y
rlabel metal2 3033 2053 3047 2067 0 _2644_.D
rlabel metal1 3184 2162 3256 2178 0 _2866_.gnd
rlabel metal1 3184 1922 3256 1938 0 _2866_.vdd
rlabel metal2 3193 2093 3207 2107 0 _2866_.A
rlabel metal2 3213 2053 3227 2067 0 _2866_.Y
rlabel metal1 3084 2162 3196 2178 0 _2645_.gnd
rlabel metal1 3084 1922 3196 1938 0 _2645_.vdd
rlabel metal2 3173 2053 3187 2067 0 _2645_.A
rlabel metal2 3153 2093 3167 2107 0 _2645_.B
rlabel metal2 3133 2053 3147 2067 0 _2645_.C
rlabel metal2 3113 2073 3127 2087 0 _2645_.Y
rlabel metal1 3444 2162 3696 2178 0 _2951_.gnd
rlabel metal1 3444 1922 3696 1938 0 _2951_.vdd
rlabel metal2 3533 2073 3547 2087 0 _2951_.D
rlabel metal2 3573 2073 3587 2087 0 _2951_.CLK
rlabel metal2 3653 2073 3667 2087 0 _2951_.Q
rlabel metal1 3244 2162 3376 2178 0 _2869_.gnd
rlabel metal1 3244 1922 3376 1938 0 _2869_.vdd
rlabel metal2 3253 2073 3267 2087 0 _2869_.A
rlabel metal2 3273 2053 3287 2067 0 _2869_.B
rlabel metal2 3333 2073 3347 2087 0 _2869_.C
rlabel metal2 3293 2073 3307 2087 0 _2869_.Y
rlabel metal2 3313 2053 3327 2067 0 _2869_.D
rlabel metal1 3364 2162 3456 2178 0 _2867_.gnd
rlabel metal1 3364 1922 3456 1938 0 _2867_.vdd
rlabel metal2 3413 2073 3427 2087 0 _2867_.B
rlabel metal2 3373 2073 3387 2087 0 _2867_.A
rlabel metal2 3393 2093 3407 2107 0 _2867_.Y
rlabel metal1 3684 2162 3776 2178 0 _2489_.gnd
rlabel metal1 3684 1922 3776 1938 0 _2489_.vdd
rlabel metal2 3713 2073 3727 2087 0 _2489_.B
rlabel metal2 3753 2073 3767 2087 0 _2489_.A
rlabel metal2 3733 2093 3747 2107 0 _2489_.Y
rlabel metal1 3764 2162 3896 2178 0 _2491_.gnd
rlabel metal1 3764 1922 3896 1938 0 _2491_.vdd
rlabel metal2 3873 2073 3887 2087 0 _2491_.A
rlabel metal2 3853 2053 3867 2067 0 _2491_.B
rlabel metal2 3793 2073 3807 2087 0 _2491_.C
rlabel metal2 3833 2073 3847 2087 0 _2491_.Y
rlabel metal2 3813 2053 3827 2067 0 _2491_.D
rlabel metal1 3944 2162 4056 2178 0 _2490_.gnd
rlabel metal1 3944 1922 4056 1938 0 _2490_.vdd
rlabel metal2 3953 2073 3967 2087 0 _2490_.A
rlabel metal2 3973 2053 3987 2067 0 _2490_.B
rlabel metal2 4013 2053 4027 2067 0 _2490_.C
rlabel metal2 3993 2073 4007 2087 0 _2490_.Y
rlabel metal1 3884 2162 3956 2178 0 _2488_.gnd
rlabel metal1 3884 1922 3956 1938 0 _2488_.vdd
rlabel metal2 3933 2093 3947 2107 0 _2488_.A
rlabel metal2 3913 2053 3927 2067 0 _2488_.Y
rlabel metal1 4204 2162 4456 2178 0 _2958_.gnd
rlabel metal1 4204 1922 4456 1938 0 _2958_.vdd
rlabel metal2 4293 2073 4307 2087 0 _2958_.D
rlabel metal2 4333 2073 4347 2087 0 _2958_.CLK
rlabel metal2 4413 2073 4427 2087 0 _2958_.Q
rlabel metal1 4124 2162 4216 2178 0 _2848_.gnd
rlabel metal1 4124 1922 4216 1938 0 _2848_.vdd
rlabel metal2 4153 2073 4167 2087 0 _2848_.B
rlabel metal2 4193 2073 4207 2087 0 _2848_.A
rlabel metal2 4173 2093 4187 2107 0 _2848_.Y
rlabel metal1 4044 2162 4136 2178 0 _2842_.gnd
rlabel metal1 4044 1922 4136 1938 0 _2842_.vdd
rlabel metal2 4053 2033 4067 2047 0 _2842_.A
rlabel metal2 4093 2033 4107 2047 0 _2842_.B
rlabel metal2 4073 2053 4087 2067 0 _2842_.Y
rlabel metal1 4504 2162 4636 2178 0 _2525_.gnd
rlabel metal1 4504 1922 4636 1938 0 _2525_.vdd
rlabel metal2 4513 2073 4527 2087 0 _2525_.A
rlabel metal2 4533 2053 4547 2067 0 _2525_.B
rlabel metal2 4593 2073 4607 2087 0 _2525_.C
rlabel metal2 4553 2073 4567 2087 0 _2525_.Y
rlabel metal2 4573 2053 4587 2067 0 _2525_.D
rlabel metal1 4444 2162 4516 2178 0 _2522_.gnd
rlabel metal1 4444 1922 4516 1938 0 _2522_.vdd
rlabel metal2 4453 2093 4467 2107 0 _2522_.A
rlabel metal2 4473 2053 4487 2067 0 _2522_.Y
rlabel metal1 4704 2162 4816 2178 0 _2524_.gnd
rlabel metal1 4704 1922 4816 1938 0 _2524_.vdd
rlabel metal2 4793 2073 4807 2087 0 _2524_.A
rlabel metal2 4773 2053 4787 2067 0 _2524_.B
rlabel metal2 4733 2053 4747 2067 0 _2524_.C
rlabel metal2 4753 2073 4767 2087 0 _2524_.Y
rlabel metal1 4804 2162 4896 2178 0 _2882_.gnd
rlabel metal1 4804 1922 4896 1938 0 _2882_.vdd
rlabel metal2 4833 2073 4847 2087 0 _2882_.B
rlabel metal2 4873 2073 4887 2087 0 _2882_.A
rlabel metal2 4853 2093 4867 2107 0 _2882_.Y
rlabel metal1 4624 2162 4716 2178 0 _2523_.gnd
rlabel metal1 4624 1922 4716 1938 0 _2523_.vdd
rlabel metal2 4673 2073 4687 2087 0 _2523_.B
rlabel metal2 4633 2073 4647 2087 0 _2523_.A
rlabel metal2 4653 2093 4667 2107 0 _2523_.Y
rlabel metal1 4884 2162 5016 2178 0 _2844_.gnd
rlabel metal1 4884 1922 5016 1938 0 _2844_.vdd
rlabel metal2 4893 2073 4907 2087 0 _2844_.A
rlabel metal2 4913 2053 4927 2067 0 _2844_.B
rlabel metal2 4973 2073 4987 2087 0 _2844_.C
rlabel metal2 4933 2073 4947 2087 0 _2844_.Y
rlabel metal2 4953 2053 4967 2067 0 _2844_.D
rlabel metal1 5004 2162 5096 2178 0 _2843_.gnd
rlabel metal1 5004 1922 5096 1938 0 _2843_.vdd
rlabel metal2 5073 2033 5087 2047 0 _2843_.A
rlabel metal2 5033 2033 5047 2047 0 _2843_.B
rlabel metal2 5053 2053 5067 2067 0 _2843_.Y
rlabel metal1 5264 2162 5396 2178 0 _2470_.gnd
rlabel metal1 5264 1922 5396 1938 0 _2470_.vdd
rlabel metal2 5373 2073 5387 2087 0 _2470_.A
rlabel metal2 5353 2053 5367 2067 0 _2470_.B
rlabel metal2 5293 2073 5307 2087 0 _2470_.C
rlabel metal2 5333 2073 5347 2087 0 _2470_.Y
rlabel metal2 5313 2053 5327 2067 0 _2470_.D
rlabel metal1 5084 2162 5176 2178 0 _2881_.gnd
rlabel metal1 5084 1922 5176 1938 0 _2881_.vdd
rlabel metal2 5113 2073 5127 2087 0 _2881_.B
rlabel metal2 5153 2073 5167 2087 0 _2881_.A
rlabel metal2 5133 2093 5147 2107 0 _2881_.Y
rlabel metal1 5164 2162 5276 2178 0 _2877_.gnd
rlabel metal1 5164 1922 5276 1938 0 _2877_.vdd
rlabel metal2 5173 2093 5187 2107 0 _2877_.A
rlabel metal2 5193 2073 5207 2087 0 _2877_.B
rlabel metal2 5233 2053 5247 2067 0 _2877_.Y
rlabel metal1 5584 2162 5716 2178 0 _2521_.gnd
rlabel metal1 5584 1922 5716 1938 0 _2521_.vdd
rlabel metal2 5693 2073 5707 2087 0 _2521_.A
rlabel metal2 5673 2053 5687 2067 0 _2521_.B
rlabel metal2 5613 2073 5627 2087 0 _2521_.C
rlabel metal2 5653 2073 5667 2087 0 _2521_.Y
rlabel metal2 5633 2053 5647 2067 0 _2521_.D
rlabel metal1 5384 2162 5516 2178 0 _2511_.gnd
rlabel metal1 5384 1922 5516 1938 0 _2511_.vdd
rlabel metal2 5393 2073 5407 2087 0 _2511_.A
rlabel metal2 5413 2053 5427 2067 0 _2511_.B
rlabel metal2 5473 2073 5487 2087 0 _2511_.C
rlabel metal2 5433 2073 5447 2087 0 _2511_.Y
rlabel metal2 5453 2053 5467 2067 0 _2511_.D
rlabel metal1 5504 2162 5596 2178 0 _2519_.gnd
rlabel metal1 5504 1922 5596 1938 0 _2519_.vdd
rlabel metal2 5533 2073 5547 2087 0 _2519_.B
rlabel metal2 5573 2073 5587 2087 0 _2519_.A
rlabel metal2 5553 2093 5567 2107 0 _2519_.Y
rlabel metal1 5844 2162 6096 2178 0 _2957_.gnd
rlabel metal1 5844 1922 6096 1938 0 _2957_.vdd
rlabel metal2 5993 2073 6007 2087 0 _2957_.D
rlabel metal2 5953 2073 5967 2087 0 _2957_.CLK
rlabel metal2 5873 2073 5887 2087 0 _2957_.Q
rlabel metal1 5704 2162 5776 2178 0 _2518_.gnd
rlabel metal1 5704 1922 5776 1938 0 _2518_.vdd
rlabel metal2 5753 2093 5767 2107 0 _2518_.A
rlabel metal2 5733 2053 5747 2067 0 _2518_.Y
rlabel metal1 5764 2162 5856 2178 0 _2463_.gnd
rlabel metal1 5764 1922 5856 1938 0 _2463_.vdd
rlabel metal2 5773 2033 5787 2047 0 _2463_.A
rlabel metal2 5813 2033 5827 2047 0 _2463_.B
rlabel metal2 5793 2053 5807 2067 0 _2463_.Y
rlabel metal1 6084 2162 6336 2178 0 _2971_.gnd
rlabel metal1 6084 1922 6336 1938 0 _2971_.vdd
rlabel metal2 6173 2073 6187 2087 0 _2971_.D
rlabel metal2 6213 2073 6227 2087 0 _2971_.CLK
rlabel metal2 6293 2073 6307 2087 0 _2971_.Q
rlabel metal1 6324 2162 6456 2178 0 _2660_.gnd
rlabel metal1 6324 1922 6455 1938 0 _2660_.vdd
rlabel metal2 6333 2053 6347 2067 0 _2660_.S
rlabel metal2 6353 2073 6367 2087 0 _2660_.B
rlabel metal2 6393 2053 6407 2067 0 _2660_.Y
rlabel metal2 6413 2073 6427 2087 0 _2660_.A
rlabel nsubstratencontact 6684 1932 6684 1932 0 FILL100050x28950.vdd
rlabel metal1 6664 2162 6696 2178 0 FILL100050x28950.gnd
rlabel nsubstratencontact 6664 1932 6664 1932 0 FILL99750x28950.vdd
rlabel metal1 6644 2162 6676 2178 0 FILL99750x28950.gnd
rlabel metal1 6544 2162 6656 2178 0 _2765_.gnd
rlabel metal1 6544 1922 6656 1938 0 _2765_.vdd
rlabel metal2 6553 2073 6567 2087 0 _2765_.A
rlabel metal2 6573 2053 6587 2067 0 _2765_.B
rlabel metal2 6613 2053 6627 2067 0 _2765_.C
rlabel metal2 6593 2073 6607 2087 0 _2765_.Y
rlabel metal1 6444 2162 6556 2178 0 _2700_.gnd
rlabel metal1 6444 1922 6556 1938 0 _2700_.vdd
rlabel metal2 6453 2053 6467 2067 0 _2700_.A
rlabel metal2 6473 2093 6487 2107 0 _2700_.B
rlabel metal2 6493 2053 6507 2067 0 _2700_.C
rlabel metal2 6513 2073 6527 2087 0 _2700_.Y
rlabel nsubstratencontact 6724 1932 6724 1932 0 FILL100650x28950.vdd
rlabel metal1 6704 2162 6736 2178 0 FILL100650x28950.gnd
rlabel nsubstratencontact 6704 1932 6704 1932 0 FILL100350x28950.vdd
rlabel metal1 6684 2162 6716 2178 0 FILL100350x28950.gnd
rlabel metal1 244 2162 336 2178 0 BUFX2_insert20.gnd
rlabel metal1 244 2402 336 2418 0 BUFX2_insert20.vdd
rlabel metal2 313 2253 327 2267 0 BUFX2_insert20.A
rlabel metal2 273 2253 287 2267 0 BUFX2_insert20.Y
rlabel metal1 4 2162 256 2178 0 _1602_.gnd
rlabel metal1 4 2402 256 2418 0 _1602_.vdd
rlabel metal2 93 2253 107 2267 0 _1602_.D
rlabel metal2 133 2253 147 2267 0 _1602_.CLK
rlabel metal2 213 2253 227 2267 0 _1602_.Q
rlabel metal1 524 2162 636 2178 0 _1594_.gnd
rlabel metal1 524 2402 636 2418 0 _1594_.vdd
rlabel metal2 533 2253 547 2267 0 _1594_.A
rlabel metal2 553 2273 567 2287 0 _1594_.B
rlabel metal2 593 2273 607 2287 0 _1594_.C
rlabel metal2 573 2253 587 2267 0 _1594_.Y
rlabel metal1 444 2162 536 2178 0 _1497_.gnd
rlabel metal1 444 2402 536 2418 0 _1497_.vdd
rlabel metal2 473 2253 487 2267 0 _1497_.B
rlabel metal2 513 2253 527 2267 0 _1497_.A
rlabel metal2 493 2233 507 2247 0 _1497_.Y
rlabel metal1 384 2162 456 2178 0 _1496_.gnd
rlabel metal1 384 2402 456 2418 0 _1496_.vdd
rlabel metal2 433 2233 447 2247 0 _1496_.A
rlabel metal2 413 2273 427 2287 0 _1496_.Y
rlabel metal1 324 2162 396 2178 0 _1498_.gnd
rlabel metal1 324 2402 396 2418 0 _1498_.vdd
rlabel metal2 373 2273 387 2287 0 _1498_.A
rlabel metal2 353 2253 367 2267 0 _1498_.Y
rlabel metal1 724 2162 836 2178 0 _1566_.gnd
rlabel metal1 724 2402 836 2418 0 _1566_.vdd
rlabel metal2 733 2273 747 2287 0 _1566_.A
rlabel metal2 753 2293 767 2307 0 _1566_.B
rlabel metal2 773 2273 787 2287 0 _1566_.C
rlabel metal2 793 2293 807 2307 0 _1566_.Y
rlabel metal1 624 2162 736 2178 0 _1567_.gnd
rlabel metal1 624 2402 736 2418 0 _1567_.vdd
rlabel metal2 713 2253 727 2267 0 _1567_.A
rlabel metal2 653 2253 667 2267 0 _1567_.Y
rlabel metal2 673 2293 687 2307 0 _1567_.B
rlabel metal1 904 2162 1156 2178 0 _1603_.gnd
rlabel metal1 904 2402 1156 2418 0 _1603_.vdd
rlabel metal2 1053 2253 1067 2267 0 _1603_.D
rlabel metal2 1013 2253 1027 2267 0 _1603_.CLK
rlabel metal2 933 2253 947 2267 0 _1603_.Q
rlabel metal1 824 2162 916 2178 0 _1499_.gnd
rlabel metal1 824 2402 916 2418 0 _1499_.vdd
rlabel metal2 833 2293 847 2307 0 _1499_.A
rlabel metal2 873 2293 887 2307 0 _1499_.B
rlabel metal2 853 2273 867 2287 0 _1499_.Y
rlabel metal1 1204 2162 1456 2178 0 _2962_.gnd
rlabel metal1 1204 2402 1456 2418 0 _2962_.vdd
rlabel metal2 1293 2253 1307 2267 0 _2962_.D
rlabel metal2 1333 2253 1347 2267 0 _2962_.CLK
rlabel metal2 1413 2253 1427 2267 0 _2962_.Q
rlabel metal1 1144 2162 1216 2178 0 _1500_.gnd
rlabel metal1 1144 2402 1216 2418 0 _1500_.vdd
rlabel metal2 1153 2233 1167 2247 0 _1500_.A
rlabel metal2 1173 2273 1187 2287 0 _1500_.Y
rlabel metal1 1504 2162 1636 2178 0 _2541_.gnd
rlabel metal1 1504 2402 1636 2418 0 _2541_.vdd
rlabel metal2 1513 2253 1527 2267 0 _2541_.A
rlabel metal2 1533 2273 1547 2287 0 _2541_.B
rlabel metal2 1593 2253 1607 2267 0 _2541_.C
rlabel metal2 1553 2253 1567 2267 0 _2541_.Y
rlabel metal2 1573 2273 1587 2287 0 _2541_.D
rlabel metal1 1444 2162 1516 2178 0 _2538_.gnd
rlabel metal1 1444 2402 1516 2418 0 _2538_.vdd
rlabel metal2 1493 2233 1507 2247 0 _2538_.A
rlabel metal2 1473 2273 1487 2287 0 _2538_.Y
rlabel metal1 1624 2162 1736 2178 0 _2482_.gnd
rlabel metal1 1624 2402 1736 2418 0 _2482_.vdd
rlabel metal2 1633 2253 1647 2267 0 _2482_.A
rlabel metal2 1653 2273 1667 2287 0 _2482_.B
rlabel metal2 1693 2273 1707 2287 0 _2482_.C
rlabel metal2 1673 2253 1687 2267 0 _2482_.Y
rlabel metal1 1724 2162 1816 2178 0 _2539_.gnd
rlabel metal1 1724 2402 1816 2418 0 _2539_.vdd
rlabel metal2 1753 2253 1767 2267 0 _2539_.B
rlabel metal2 1793 2253 1807 2267 0 _2539_.A
rlabel metal2 1773 2233 1787 2247 0 _2539_.Y
rlabel metal1 1804 2162 1896 2178 0 _2481_.gnd
rlabel metal1 1804 2402 1896 2418 0 _2481_.vdd
rlabel metal2 1833 2253 1847 2267 0 _2481_.B
rlabel metal2 1873 2253 1887 2267 0 _2481_.A
rlabel metal2 1853 2233 1867 2247 0 _2481_.Y
rlabel metal1 2064 2162 2316 2178 0 _2949_.gnd
rlabel metal1 2064 2402 2316 2418 0 _2949_.vdd
rlabel metal2 2153 2253 2167 2267 0 _2949_.D
rlabel metal2 2193 2253 2207 2267 0 _2949_.CLK
rlabel metal2 2273 2253 2287 2267 0 _2949_.Q
rlabel metal1 1884 2162 2016 2178 0 _2483_.gnd
rlabel metal1 1884 2402 2016 2418 0 _2483_.vdd
rlabel metal2 1993 2253 2007 2267 0 _2483_.A
rlabel metal2 1973 2273 1987 2287 0 _2483_.B
rlabel metal2 1913 2253 1927 2267 0 _2483_.C
rlabel metal2 1953 2253 1967 2267 0 _2483_.Y
rlabel metal2 1933 2273 1947 2287 0 _2483_.D
rlabel metal1 2004 2162 2076 2178 0 _2480_.gnd
rlabel metal1 2004 2402 2076 2418 0 _2480_.vdd
rlabel metal2 2053 2233 2067 2247 0 _2480_.A
rlabel metal2 2033 2273 2047 2287 0 _2480_.Y
rlabel metal1 2384 2162 2496 2178 0 _2888_.gnd
rlabel metal1 2384 2402 2496 2418 0 _2888_.vdd
rlabel metal2 2393 2253 2407 2267 0 _2888_.A
rlabel metal2 2413 2273 2427 2287 0 _2888_.B
rlabel metal2 2453 2273 2467 2287 0 _2888_.C
rlabel metal2 2433 2253 2447 2267 0 _2888_.Y
rlabel metal1 2304 2162 2396 2178 0 _2886_.gnd
rlabel metal1 2304 2402 2396 2418 0 _2886_.vdd
rlabel metal2 2333 2253 2347 2267 0 _2886_.B
rlabel metal2 2373 2253 2387 2267 0 _2886_.A
rlabel metal2 2353 2233 2367 2247 0 _2886_.Y
rlabel metal1 2584 2162 2696 2178 0 _2887_.gnd
rlabel metal1 2584 2402 2696 2418 0 _2887_.vdd
rlabel metal2 2673 2273 2687 2287 0 _2887_.A
rlabel metal2 2653 2233 2667 2247 0 _2887_.B
rlabel metal2 2633 2273 2647 2287 0 _2887_.C
rlabel metal2 2613 2253 2627 2267 0 _2887_.Y
rlabel metal1 2484 2162 2596 2178 0 _2885_.gnd
rlabel metal1 2484 2402 2596 2418 0 _2885_.vdd
rlabel metal2 2573 2273 2587 2287 0 _2885_.A
rlabel metal2 2553 2293 2567 2307 0 _2885_.B
rlabel metal2 2533 2273 2547 2287 0 _2885_.C
rlabel metal2 2513 2293 2527 2307 0 _2885_.Y
rlabel metal1 2864 2162 3116 2178 0 _3009_.gnd
rlabel metal1 2864 2402 3116 2418 0 _3009_.vdd
rlabel metal2 3013 2253 3027 2267 0 _3009_.D
rlabel metal2 2973 2253 2987 2267 0 _3009_.CLK
rlabel metal2 2893 2253 2907 2267 0 _3009_.Q
rlabel metal1 2684 2162 2796 2178 0 _2853_.gnd
rlabel metal1 2684 2402 2796 2418 0 _2853_.vdd
rlabel metal2 2693 2253 2707 2267 0 _2853_.A
rlabel metal2 2713 2273 2727 2287 0 _2853_.B
rlabel metal2 2753 2273 2767 2287 0 _2853_.C
rlabel metal2 2733 2253 2747 2267 0 _2853_.Y
rlabel metal1 2784 2162 2876 2178 0 _2852_.gnd
rlabel metal1 2784 2402 2876 2418 0 _2852_.vdd
rlabel metal2 2813 2253 2827 2267 0 _2852_.B
rlabel metal2 2853 2253 2867 2267 0 _2852_.A
rlabel metal2 2833 2233 2847 2247 0 _2852_.Y
rlabel metal1 3204 2162 3336 2178 0 _2529_.gnd
rlabel metal1 3204 2402 3336 2418 0 _2529_.vdd
rlabel metal2 3313 2253 3327 2267 0 _2529_.A
rlabel metal2 3293 2273 3307 2287 0 _2529_.B
rlabel metal2 3233 2253 3247 2267 0 _2529_.C
rlabel metal2 3273 2253 3287 2267 0 _2529_.Y
rlabel metal2 3253 2273 3267 2287 0 _2529_.D
rlabel metal1 3104 2162 3216 2178 0 _2528_.gnd
rlabel metal1 3104 2402 3216 2418 0 _2528_.vdd
rlabel metal2 3113 2253 3127 2267 0 _2528_.A
rlabel metal2 3133 2273 3147 2287 0 _2528_.B
rlabel metal2 3173 2273 3187 2287 0 _2528_.C
rlabel metal2 3153 2253 3167 2267 0 _2528_.Y
rlabel metal1 3324 2162 3416 2178 0 _2527_.gnd
rlabel metal1 3324 2402 3416 2418 0 _2527_.vdd
rlabel metal2 3353 2253 3367 2267 0 _2527_.B
rlabel metal2 3393 2253 3407 2267 0 _2527_.A
rlabel metal2 3373 2233 3387 2247 0 _2527_.Y
rlabel metal1 3464 2162 3556 2178 0 _2474_.gnd
rlabel metal1 3464 2402 3556 2418 0 _2474_.vdd
rlabel metal2 3493 2253 3507 2267 0 _2474_.B
rlabel metal2 3533 2253 3547 2267 0 _2474_.A
rlabel metal2 3513 2233 3527 2247 0 _2474_.Y
rlabel metal1 3404 2162 3476 2178 0 _2526_.gnd
rlabel metal1 3404 2402 3476 2418 0 _2526_.vdd
rlabel metal2 3453 2233 3467 2247 0 _2526_.A
rlabel metal2 3433 2273 3447 2287 0 _2526_.Y
rlabel metal1 3544 2162 3796 2178 0 _2959_.gnd
rlabel metal1 3544 2402 3796 2418 0 _2959_.vdd
rlabel metal2 3633 2253 3647 2267 0 _2959_.D
rlabel metal2 3673 2253 3687 2267 0 _2959_.CLK
rlabel metal2 3753 2253 3767 2267 0 _2959_.Q
rlabel metal1 3784 2162 3876 2178 0 _2467_.gnd
rlabel metal1 3784 2402 3876 2418 0 _2467_.vdd
rlabel metal2 3793 2293 3807 2307 0 _2467_.A
rlabel metal2 3833 2293 3847 2307 0 _2467_.B
rlabel metal2 3813 2273 3827 2287 0 _2467_.Y
rlabel metal1 3864 2162 3976 2178 0 _2600_.gnd
rlabel metal1 3864 2402 3976 2418 0 _2600_.vdd
rlabel metal2 3873 2273 3887 2287 0 _2600_.A
rlabel metal2 3893 2293 3907 2307 0 _2600_.B
rlabel metal2 3913 2273 3927 2287 0 _2600_.C
rlabel metal2 3933 2293 3947 2307 0 _2600_.Y
rlabel metal1 3964 2162 4096 2178 0 _2713_.gnd
rlabel metal1 3964 2402 4095 2418 0 _2713_.vdd
rlabel metal2 3973 2273 3987 2287 0 _2713_.S
rlabel metal2 3993 2253 4007 2267 0 _2713_.B
rlabel metal2 4033 2273 4047 2287 0 _2713_.Y
rlabel metal2 4053 2253 4067 2267 0 _2713_.A
rlabel metal1 4084 2162 4216 2178 0 _2715_.gnd
rlabel metal1 4084 2402 4215 2418 0 _2715_.vdd
rlabel metal2 4093 2273 4107 2287 0 _2715_.S
rlabel metal2 4113 2253 4127 2267 0 _2715_.B
rlabel metal2 4153 2273 4167 2287 0 _2715_.Y
rlabel metal2 4173 2253 4187 2267 0 _2715_.A
rlabel metal1 4204 2162 4336 2178 0 _2625_.gnd
rlabel metal1 4204 2402 4335 2418 0 _2625_.vdd
rlabel metal2 4213 2273 4227 2287 0 _2625_.S
rlabel metal2 4233 2253 4247 2267 0 _2625_.B
rlabel metal2 4273 2273 4287 2287 0 _2625_.Y
rlabel metal2 4293 2253 4307 2267 0 _2625_.A
rlabel metal1 4324 2162 4416 2178 0 BUFX2_insert7.gnd
rlabel metal1 4324 2402 4416 2418 0 BUFX2_insert7.vdd
rlabel metal2 4333 2253 4347 2267 0 BUFX2_insert7.A
rlabel metal2 4373 2253 4387 2267 0 BUFX2_insert7.Y
rlabel metal1 4404 2162 4496 2178 0 _2477_.gnd
rlabel metal1 4404 2402 4496 2418 0 _2477_.vdd
rlabel metal2 4433 2253 4447 2267 0 _2477_.B
rlabel metal2 4473 2253 4487 2267 0 _2477_.A
rlabel metal2 4453 2233 4467 2247 0 _2477_.Y
rlabel metal1 4484 2162 4616 2178 0 _2615_.gnd
rlabel metal1 4484 2402 4615 2418 0 _2615_.vdd
rlabel metal2 4493 2273 4507 2287 0 _2615_.S
rlabel metal2 4513 2253 4527 2267 0 _2615_.B
rlabel metal2 4553 2273 4567 2287 0 _2615_.Y
rlabel metal2 4573 2253 4587 2267 0 _2615_.A
rlabel metal1 4724 2162 4856 2178 0 _2703_.gnd
rlabel metal1 4724 2402 4855 2418 0 _2703_.vdd
rlabel metal2 4733 2273 4747 2287 0 _2703_.S
rlabel metal2 4753 2253 4767 2267 0 _2703_.B
rlabel metal2 4793 2273 4807 2287 0 _2703_.Y
rlabel metal2 4813 2253 4827 2267 0 _2703_.A
rlabel metal1 4604 2162 4736 2178 0 _2701_.gnd
rlabel metal1 4605 2402 4736 2418 0 _2701_.vdd
rlabel metal2 4713 2273 4727 2287 0 _2701_.S
rlabel metal2 4693 2253 4707 2267 0 _2701_.B
rlabel metal2 4653 2273 4667 2287 0 _2701_.Y
rlabel metal2 4633 2253 4647 2267 0 _2701_.A
rlabel metal1 4844 2162 4936 2178 0 _2515_.gnd
rlabel metal1 4844 2402 4936 2418 0 _2515_.vdd
rlabel metal2 4893 2253 4907 2267 0 _2515_.B
rlabel metal2 4853 2253 4867 2267 0 _2515_.A
rlabel metal2 4873 2233 4887 2247 0 _2515_.Y
rlabel metal1 5044 2162 5156 2178 0 _2603_.gnd
rlabel metal1 5044 2402 5156 2418 0 _2603_.vdd
rlabel metal2 5133 2273 5147 2287 0 _2603_.A
rlabel metal2 5113 2233 5127 2247 0 _2603_.B
rlabel metal2 5093 2273 5107 2287 0 _2603_.C
rlabel metal2 5073 2253 5087 2267 0 _2603_.Y
rlabel metal1 4924 2162 5056 2178 0 _2690_.gnd
rlabel metal1 4924 2402 5055 2418 0 _2690_.vdd
rlabel metal2 4933 2273 4947 2287 0 _2690_.S
rlabel metal2 4953 2253 4967 2267 0 _2690_.B
rlabel metal2 4993 2273 5007 2287 0 _2690_.Y
rlabel metal2 5013 2253 5027 2267 0 _2690_.A
rlabel metal1 5204 2162 5336 2178 0 _2602_.gnd
rlabel metal1 5204 2402 5336 2418 0 _2602_.vdd
rlabel metal2 5213 2253 5227 2267 0 _2602_.A
rlabel metal2 5233 2273 5247 2287 0 _2602_.B
rlabel metal2 5293 2253 5307 2267 0 _2602_.C
rlabel metal2 5253 2253 5267 2267 0 _2602_.Y
rlabel metal2 5273 2273 5287 2287 0 _2602_.D
rlabel metal1 5144 2162 5216 2178 0 _2599_.gnd
rlabel metal1 5144 2402 5216 2418 0 _2599_.vdd
rlabel metal2 5153 2233 5167 2247 0 _2599_.A
rlabel metal2 5173 2273 5187 2287 0 _2599_.Y
rlabel metal1 5324 2162 5456 2178 0 _2601_.gnd
rlabel metal1 5325 2402 5456 2418 0 _2601_.vdd
rlabel metal2 5433 2273 5447 2287 0 _2601_.S
rlabel metal2 5413 2253 5427 2267 0 _2601_.B
rlabel metal2 5373 2273 5387 2287 0 _2601_.Y
rlabel metal2 5353 2253 5367 2267 0 _2601_.A
rlabel metal1 5564 2162 5696 2178 0 _2691_.gnd
rlabel metal1 5564 2402 5695 2418 0 _2691_.vdd
rlabel metal2 5573 2273 5587 2287 0 _2691_.S
rlabel metal2 5593 2253 5607 2267 0 _2691_.B
rlabel metal2 5633 2273 5647 2287 0 _2691_.Y
rlabel metal2 5653 2253 5667 2267 0 _2691_.A
rlabel metal1 5444 2162 5576 2178 0 _2689_.gnd
rlabel metal1 5444 2402 5575 2418 0 _2689_.vdd
rlabel metal2 5453 2273 5467 2287 0 _2689_.S
rlabel metal2 5473 2253 5487 2267 0 _2689_.B
rlabel metal2 5513 2273 5527 2287 0 _2689_.Y
rlabel metal2 5533 2253 5547 2267 0 _2689_.A
rlabel metal1 5784 2162 5896 2178 0 _2509_.gnd
rlabel metal1 5784 2402 5896 2418 0 _2509_.vdd
rlabel metal2 5873 2273 5887 2287 0 _2509_.A
rlabel metal2 5853 2293 5867 2307 0 _2509_.B
rlabel metal2 5833 2273 5847 2287 0 _2509_.C
rlabel metal2 5813 2293 5827 2307 0 _2509_.Y
rlabel metal1 5684 2162 5796 2178 0 _2465_.gnd
rlabel metal1 5684 2402 5796 2418 0 _2465_.vdd
rlabel metal2 5773 2273 5787 2287 0 _2465_.A
rlabel metal2 5753 2293 5767 2307 0 _2465_.B
rlabel metal2 5733 2273 5747 2287 0 _2465_.C
rlabel metal2 5713 2293 5727 2307 0 _2465_.Y
rlabel metal1 5884 2162 5956 2178 0 _2464_.gnd
rlabel metal1 5884 2402 5956 2418 0 _2464_.vdd
rlabel metal2 5933 2233 5947 2247 0 _2464_.A
rlabel metal2 5913 2273 5927 2287 0 _2464_.Y
rlabel metal1 5944 2162 6076 2178 0 _2706_.gnd
rlabel metal1 5944 2402 6076 2418 0 _2706_.vdd
rlabel metal2 6053 2253 6067 2267 0 _2706_.A
rlabel metal2 6033 2273 6047 2287 0 _2706_.B
rlabel metal2 5973 2253 5987 2267 0 _2706_.C
rlabel metal2 5993 2273 6007 2287 0 _2706_.D
rlabel metal2 6013 2253 6027 2267 0 _2706_.Y
rlabel metal1 6064 2162 6196 2178 0 _2661_.gnd
rlabel metal1 6065 2402 6196 2418 0 _2661_.vdd
rlabel metal2 6173 2273 6187 2287 0 _2661_.S
rlabel metal2 6153 2253 6167 2267 0 _2661_.B
rlabel metal2 6113 2273 6127 2287 0 _2661_.Y
rlabel metal2 6093 2253 6107 2267 0 _2661_.A
rlabel metal1 6364 2162 6476 2178 0 _2759_.gnd
rlabel metal1 6364 2402 6476 2418 0 _2759_.vdd
rlabel metal2 6373 2253 6387 2267 0 _2759_.A
rlabel metal2 6393 2273 6407 2287 0 _2759_.B
rlabel metal2 6433 2273 6447 2287 0 _2759_.C
rlabel metal2 6413 2253 6427 2267 0 _2759_.Y
rlabel metal1 6304 2162 6376 2178 0 _2757_.gnd
rlabel metal1 6304 2402 6376 2418 0 _2757_.vdd
rlabel metal2 6313 2233 6327 2247 0 _2757_.A
rlabel metal2 6333 2273 6347 2287 0 _2757_.Y
rlabel metal1 6184 2162 6316 2178 0 _2659_.gnd
rlabel metal1 6185 2402 6316 2418 0 _2659_.vdd
rlabel metal2 6293 2273 6307 2287 0 _2659_.S
rlabel metal2 6273 2253 6287 2267 0 _2659_.B
rlabel metal2 6233 2273 6247 2287 0 _2659_.Y
rlabel metal2 6213 2253 6227 2267 0 _2659_.A
rlabel metal1 6644 2162 6716 2178 0 _2696_.gnd
rlabel metal1 6644 2402 6716 2418 0 _2696_.vdd
rlabel metal2 6653 2233 6667 2247 0 _2696_.A
rlabel metal2 6673 2273 6687 2287 0 _2696_.Y
rlabel metal1 6464 2162 6556 2178 0 _2758_.gnd
rlabel metal1 6464 2402 6556 2418 0 _2758_.vdd
rlabel metal2 6473 2293 6487 2307 0 _2758_.A
rlabel metal2 6513 2293 6527 2307 0 _2758_.B
rlabel metal2 6493 2273 6507 2287 0 _2758_.Y
rlabel metal1 6544 2162 6656 2178 0 _2760_.gnd
rlabel metal1 6544 2402 6656 2418 0 _2760_.vdd
rlabel metal2 6553 2273 6567 2287 0 _2760_.A
rlabel metal2 6573 2233 6587 2247 0 _2760_.B
rlabel metal2 6593 2273 6607 2287 0 _2760_.C
rlabel metal2 6613 2253 6627 2267 0 _2760_.Y
rlabel nsubstratencontact 6716 2408 6716 2408 0 FILL100650x32550.vdd
rlabel metal1 6704 2162 6736 2178 0 FILL100650x32550.gnd
rlabel metal1 244 2642 336 2658 0 _3044_.gnd
rlabel metal1 244 2402 336 2418 0 _3044_.vdd
rlabel metal2 313 2553 327 2567 0 _3044_.A
rlabel metal2 273 2553 287 2567 0 _3044_.Y
rlabel metal1 4 2642 256 2658 0 _1627_.gnd
rlabel metal1 4 2402 256 2418 0 _1627_.vdd
rlabel metal2 153 2553 167 2567 0 _1627_.D
rlabel metal2 113 2553 127 2567 0 _1627_.CLK
rlabel metal2 33 2553 47 2567 0 _1627_.Q
rlabel metal1 324 2642 576 2658 0 _1615_.gnd
rlabel metal1 324 2402 576 2418 0 _1615_.vdd
rlabel metal2 473 2553 487 2567 0 _1615_.D
rlabel metal2 433 2553 447 2567 0 _1615_.CLK
rlabel metal2 353 2553 367 2567 0 _1615_.Q
rlabel metal1 744 2642 836 2658 0 _1533_.gnd
rlabel metal1 744 2402 836 2418 0 _1533_.vdd
rlabel metal2 813 2513 827 2527 0 _1533_.A
rlabel metal2 773 2513 787 2527 0 _1533_.B
rlabel metal2 793 2533 807 2547 0 _1533_.Y
rlabel metal1 664 2642 756 2658 0 _1531_.gnd
rlabel metal1 664 2402 756 2418 0 _1531_.vdd
rlabel metal2 673 2513 687 2527 0 _1531_.A
rlabel metal2 713 2513 727 2527 0 _1531_.B
rlabel metal2 693 2533 707 2547 0 _1531_.Y
rlabel metal1 564 2642 676 2658 0 _1583_.gnd
rlabel metal1 564 2402 676 2418 0 _1583_.vdd
rlabel metal2 653 2533 667 2547 0 _1583_.A
rlabel metal2 633 2573 647 2587 0 _1583_.B
rlabel metal2 613 2533 627 2547 0 _1583_.C
rlabel metal2 593 2553 607 2567 0 _1583_.Y
rlabel metal1 824 2642 1036 2658 0 CLKBUF1_insert35.gnd
rlabel metal1 824 2402 1036 2418 0 CLKBUF1_insert35.vdd
rlabel metal2 993 2533 1007 2547 0 CLKBUF1_insert35.A
rlabel metal2 853 2533 867 2547 0 CLKBUF1_insert35.Y
rlabel metal1 1024 2642 1276 2658 0 _2387_.gnd
rlabel metal1 1024 2402 1276 2418 0 _2387_.vdd
rlabel metal2 1173 2553 1187 2567 0 _2387_.D
rlabel metal2 1133 2553 1147 2567 0 _2387_.CLK
rlabel metal2 1053 2553 1067 2567 0 _2387_.Q
rlabel metal1 1264 2642 1356 2658 0 _2250_.gnd
rlabel metal1 1264 2402 1356 2418 0 _2250_.vdd
rlabel metal2 1333 2513 1347 2527 0 _2250_.A
rlabel metal2 1293 2513 1307 2527 0 _2250_.B
rlabel metal2 1313 2533 1327 2547 0 _2250_.Y
rlabel metal1 1584 2642 1836 2658 0 _2954_.gnd
rlabel metal1 1584 2402 1836 2418 0 _2954_.vdd
rlabel metal2 1673 2553 1687 2567 0 _2954_.D
rlabel metal2 1713 2553 1727 2567 0 _2954_.CLK
rlabel metal2 1793 2553 1807 2567 0 _2954_.Q
rlabel metal1 1484 2642 1596 2658 0 _2264_.gnd
rlabel metal1 1484 2402 1596 2418 0 _2264_.vdd
rlabel metal2 1573 2553 1587 2567 0 _2264_.A
rlabel metal2 1553 2533 1567 2547 0 _2264_.B
rlabel metal2 1513 2533 1527 2547 0 _2264_.C
rlabel metal2 1533 2553 1547 2567 0 _2264_.Y
rlabel metal1 1344 2642 1436 2658 0 _2252_.gnd
rlabel metal1 1344 2402 1436 2418 0 _2252_.vdd
rlabel metal2 1393 2553 1407 2567 0 _2252_.B
rlabel metal2 1353 2553 1367 2567 0 _2252_.A
rlabel metal2 1373 2573 1387 2587 0 _2252_.Y
rlabel metal1 1424 2642 1496 2658 0 _2251_.gnd
rlabel metal1 1424 2402 1496 2418 0 _2251_.vdd
rlabel metal2 1433 2573 1447 2587 0 _2251_.A
rlabel metal2 1453 2533 1467 2547 0 _2251_.Y
rlabel metal1 1824 2642 1896 2658 0 _2242_.gnd
rlabel metal1 1824 2402 1896 2418 0 _2242_.vdd
rlabel metal2 1833 2573 1847 2587 0 _2242_.A
rlabel metal2 1853 2533 1867 2547 0 _2242_.Y
rlabel metal1 1944 2642 2076 2658 0 _2503_.gnd
rlabel metal1 1944 2402 2076 2418 0 _2503_.vdd
rlabel metal2 1953 2553 1967 2567 0 _2503_.A
rlabel metal2 1973 2533 1987 2547 0 _2503_.B
rlabel metal2 2033 2553 2047 2567 0 _2503_.C
rlabel metal2 1993 2553 2007 2567 0 _2503_.Y
rlabel metal2 2013 2533 2027 2547 0 _2503_.D
rlabel metal1 2064 2642 2156 2658 0 _2501_.gnd
rlabel metal1 2064 2402 2156 2418 0 _2501_.vdd
rlabel metal2 2113 2553 2127 2567 0 _2501_.B
rlabel metal2 2073 2553 2087 2567 0 _2501_.A
rlabel metal2 2093 2573 2107 2587 0 _2501_.Y
rlabel metal1 1884 2642 1956 2658 0 _2500_.gnd
rlabel metal1 1884 2402 1956 2418 0 _2500_.vdd
rlabel metal2 1893 2573 1907 2587 0 _2500_.A
rlabel metal2 1913 2533 1927 2547 0 _2500_.Y
rlabel metal1 2384 2642 2636 2658 0 _3013_.gnd
rlabel metal1 2384 2402 2636 2418 0 _3013_.vdd
rlabel metal2 2473 2553 2487 2567 0 _3013_.D
rlabel metal2 2513 2553 2527 2567 0 _3013_.CLK
rlabel metal2 2593 2553 2607 2567 0 _3013_.Q
rlabel metal1 2264 2642 2396 2658 0 _2749_.gnd
rlabel metal1 2264 2402 2395 2418 0 _2749_.vdd
rlabel metal2 2273 2533 2287 2547 0 _2749_.S
rlabel metal2 2293 2553 2307 2567 0 _2749_.B
rlabel metal2 2333 2533 2347 2547 0 _2749_.Y
rlabel metal2 2353 2553 2367 2567 0 _2749_.A
rlabel metal1 2144 2642 2276 2658 0 _2654_.gnd
rlabel metal1 2144 2402 2275 2418 0 _2654_.vdd
rlabel metal2 2153 2533 2167 2547 0 _2654_.S
rlabel metal2 2173 2553 2187 2567 0 _2654_.B
rlabel metal2 2213 2533 2227 2547 0 _2654_.Y
rlabel metal2 2233 2553 2247 2567 0 _2654_.A
rlabel metal1 2624 2642 2756 2658 0 _2751_.gnd
rlabel metal1 2624 2402 2755 2418 0 _2751_.vdd
rlabel metal2 2633 2533 2647 2547 0 _2751_.S
rlabel metal2 2653 2553 2667 2567 0 _2751_.B
rlabel metal2 2693 2533 2707 2547 0 _2751_.Y
rlabel metal2 2713 2553 2727 2567 0 _2751_.A
rlabel metal1 2744 2642 2836 2658 0 _2906_.gnd
rlabel metal1 2744 2402 2836 2418 0 _2906_.vdd
rlabel metal2 2773 2553 2787 2567 0 _2906_.B
rlabel metal2 2813 2553 2827 2567 0 _2906_.A
rlabel metal2 2793 2573 2807 2587 0 _2906_.Y
rlabel metal1 2824 2642 2956 2658 0 _2750_.gnd
rlabel metal1 2825 2402 2956 2418 0 _2750_.vdd
rlabel metal2 2933 2533 2947 2547 0 _2750_.S
rlabel metal2 2913 2553 2927 2567 0 _2750_.B
rlabel metal2 2873 2533 2887 2547 0 _2750_.Y
rlabel metal2 2853 2553 2867 2567 0 _2750_.A
rlabel metal1 3124 2642 3376 2658 0 _3005_.gnd
rlabel metal1 3124 2402 3376 2418 0 _3005_.vdd
rlabel metal2 3213 2553 3227 2567 0 _3005_.D
rlabel metal2 3253 2553 3267 2567 0 _3005_.CLK
rlabel metal2 3333 2553 3347 2567 0 _3005_.Q
rlabel metal1 2944 2642 3076 2658 0 _2854_.gnd
rlabel metal1 2944 2402 3076 2418 0 _2854_.vdd
rlabel metal2 3053 2553 3067 2567 0 _2854_.A
rlabel metal2 3033 2533 3047 2547 0 _2854_.B
rlabel metal2 2973 2553 2987 2567 0 _2854_.C
rlabel metal2 3013 2553 3027 2567 0 _2854_.Y
rlabel metal2 2993 2533 3007 2547 0 _2854_.D
rlabel metal1 3064 2642 3136 2658 0 _2851_.gnd
rlabel metal1 3064 2402 3136 2418 0 _2851_.vdd
rlabel metal2 3113 2573 3127 2587 0 _2851_.A
rlabel metal2 3093 2533 3107 2547 0 _2851_.Y
rlabel metal1 3364 2642 3456 2658 0 _2870_.gnd
rlabel metal1 3364 2402 3456 2418 0 _2870_.vdd
rlabel metal2 3413 2553 3427 2567 0 _2870_.B
rlabel metal2 3373 2553 3387 2567 0 _2870_.A
rlabel metal2 3393 2573 3407 2587 0 _2870_.Y
rlabel metal1 3444 2642 3536 2658 0 _2473_.gnd
rlabel metal1 3444 2402 3536 2418 0 _2473_.vdd
rlabel metal2 3513 2513 3527 2527 0 _2473_.A
rlabel metal2 3473 2513 3487 2527 0 _2473_.B
rlabel metal2 3493 2533 3507 2547 0 _2473_.Y
rlabel metal1 3524 2642 3596 2658 0 _2468_.gnd
rlabel metal1 3524 2402 3596 2418 0 _2468_.vdd
rlabel metal2 3533 2573 3547 2587 0 _2468_.A
rlabel metal2 3553 2533 3567 2547 0 _2468_.Y
rlabel metal1 3584 2642 3696 2658 0 _2604_.gnd
rlabel metal1 3584 2402 3696 2418 0 _2604_.vdd
rlabel metal2 3593 2533 3607 2547 0 _2604_.A
rlabel metal2 3613 2513 3627 2527 0 _2604_.B
rlabel metal2 3633 2533 3647 2547 0 _2604_.C
rlabel metal2 3653 2513 3667 2527 0 _2604_.Y
rlabel metal1 3684 2642 3796 2658 0 _2469_.gnd
rlabel metal1 3684 2402 3796 2418 0 _2469_.vdd
rlabel metal2 3693 2533 3707 2547 0 _2469_.A
rlabel metal2 3713 2513 3727 2527 0 _2469_.B
rlabel metal2 3733 2533 3747 2547 0 _2469_.C
rlabel metal2 3753 2513 3767 2527 0 _2469_.Y
rlabel metal1 3884 2642 3996 2658 0 _2856_.gnd
rlabel metal1 3884 2402 3996 2418 0 _2856_.vdd
rlabel metal2 3893 2553 3907 2567 0 _2856_.A
rlabel metal2 3913 2533 3927 2547 0 _2856_.B
rlabel metal2 3953 2533 3967 2547 0 _2856_.C
rlabel metal2 3933 2553 3947 2567 0 _2856_.Y
rlabel metal1 3984 2642 4096 2658 0 _2891_.gnd
rlabel metal1 3984 2402 4096 2418 0 _2891_.vdd
rlabel metal2 3993 2533 4007 2547 0 _2891_.A
rlabel metal2 4013 2573 4027 2587 0 _2891_.B
rlabel metal2 4033 2533 4047 2547 0 _2891_.C
rlabel metal2 4053 2553 4067 2567 0 _2891_.Y
rlabel metal1 3784 2642 3896 2658 0 _2510_.gnd
rlabel metal1 3784 2402 3896 2418 0 _2510_.vdd
rlabel metal2 3873 2533 3887 2547 0 _2510_.A
rlabel metal2 3853 2513 3867 2527 0 _2510_.B
rlabel metal2 3833 2533 3847 2547 0 _2510_.C
rlabel metal2 3813 2513 3827 2527 0 _2510_.Y
rlabel metal1 4164 2642 4296 2658 0 _2857_.gnd
rlabel metal1 4164 2402 4296 2418 0 _2857_.vdd
rlabel metal2 4273 2553 4287 2567 0 _2857_.A
rlabel metal2 4253 2533 4267 2547 0 _2857_.B
rlabel metal2 4193 2553 4207 2567 0 _2857_.C
rlabel metal2 4233 2553 4247 2567 0 _2857_.Y
rlabel metal2 4213 2533 4227 2547 0 _2857_.D
rlabel metal1 4084 2642 4176 2658 0 _2855_.gnd
rlabel metal1 4084 2402 4176 2418 0 _2855_.vdd
rlabel metal2 4113 2553 4127 2567 0 _2855_.B
rlabel metal2 4153 2553 4167 2567 0 _2855_.A
rlabel metal2 4133 2573 4147 2587 0 _2855_.Y
rlabel metal1 4284 2642 4536 2658 0 _3006_.gnd
rlabel metal1 4284 2402 4536 2418 0 _3006_.vdd
rlabel metal2 4373 2553 4387 2567 0 _3006_.D
rlabel metal2 4413 2553 4427 2567 0 _3006_.CLK
rlabel metal2 4493 2553 4507 2567 0 _3006_.Q
rlabel metal1 4524 2642 4596 2658 0 _2614_.gnd
rlabel metal1 4524 2402 4596 2418 0 _2614_.vdd
rlabel metal2 4573 2573 4587 2587 0 _2614_.A
rlabel metal2 4553 2533 4567 2547 0 _2614_.Y
rlabel metal1 4584 2642 4716 2658 0 _2616_.gnd
rlabel metal1 4584 2402 4716 2418 0 _2616_.vdd
rlabel metal2 4693 2553 4707 2567 0 _2616_.A
rlabel metal2 4673 2533 4687 2547 0 _2616_.B
rlabel metal2 4613 2553 4627 2567 0 _2616_.C
rlabel metal2 4653 2553 4667 2567 0 _2616_.Y
rlabel metal2 4633 2533 4647 2547 0 _2616_.D
rlabel metal1 4704 2642 4836 2658 0 _2702_.gnd
rlabel metal1 4704 2402 4835 2418 0 _2702_.vdd
rlabel metal2 4713 2533 4727 2547 0 _2702_.S
rlabel metal2 4733 2553 4747 2567 0 _2702_.B
rlabel metal2 4773 2533 4787 2547 0 _2702_.Y
rlabel metal2 4793 2553 4807 2567 0 _2702_.A
rlabel metal1 4824 2642 5076 2658 0 _2950_.gnd
rlabel metal1 4824 2402 5076 2418 0 _2950_.vdd
rlabel metal2 4973 2553 4987 2567 0 _2950_.D
rlabel metal2 4933 2553 4947 2567 0 _2950_.CLK
rlabel metal2 4853 2553 4867 2567 0 _2950_.Q
rlabel metal1 5064 2642 5136 2658 0 _2484_.gnd
rlabel metal1 5064 2402 5136 2418 0 _2484_.vdd
rlabel metal2 5073 2573 5087 2587 0 _2484_.A
rlabel metal2 5093 2533 5107 2547 0 _2484_.Y
rlabel metal1 5124 2642 5256 2658 0 _2487_.gnd
rlabel metal1 5124 2402 5256 2418 0 _2487_.vdd
rlabel metal2 5133 2553 5147 2567 0 _2487_.A
rlabel metal2 5153 2533 5167 2547 0 _2487_.B
rlabel metal2 5213 2553 5227 2567 0 _2487_.C
rlabel metal2 5173 2553 5187 2567 0 _2487_.Y
rlabel metal2 5193 2533 5207 2547 0 _2487_.D
rlabel metal1 5244 2642 5356 2658 0 _2486_.gnd
rlabel metal1 5244 2402 5356 2418 0 _2486_.vdd
rlabel metal2 5253 2553 5267 2567 0 _2486_.A
rlabel metal2 5273 2533 5287 2547 0 _2486_.B
rlabel metal2 5313 2533 5327 2547 0 _2486_.C
rlabel metal2 5293 2553 5307 2567 0 _2486_.Y
rlabel metal1 5504 2642 5716 2658 0 CLKBUF1_insert37.gnd
rlabel metal1 5504 2402 5716 2418 0 CLKBUF1_insert37.vdd
rlabel metal2 5533 2533 5547 2547 0 CLKBUF1_insert37.A
rlabel metal2 5673 2533 5687 2547 0 CLKBUF1_insert37.Y
rlabel metal1 5424 2642 5516 2658 0 _2505_.gnd
rlabel metal1 5424 2402 5516 2418 0 _2505_.vdd
rlabel metal2 5453 2553 5467 2567 0 _2505_.B
rlabel metal2 5493 2553 5507 2567 0 _2505_.A
rlabel metal2 5473 2573 5487 2587 0 _2505_.Y
rlabel metal1 5344 2642 5436 2658 0 _2485_.gnd
rlabel metal1 5344 2402 5436 2418 0 _2485_.vdd
rlabel metal2 5393 2553 5407 2567 0 _2485_.B
rlabel metal2 5353 2553 5367 2567 0 _2485_.A
rlabel metal2 5373 2573 5387 2587 0 _2485_.Y
rlabel metal1 5784 2642 5896 2658 0 _2544_.gnd
rlabel metal1 5784 2402 5896 2418 0 _2544_.vdd
rlabel metal2 5793 2553 5807 2567 0 _2544_.A
rlabel metal2 5813 2533 5827 2547 0 _2544_.B
rlabel metal2 5853 2533 5867 2547 0 _2544_.C
rlabel metal2 5833 2553 5847 2567 0 _2544_.Y
rlabel metal1 5704 2642 5796 2658 0 _2543_.gnd
rlabel metal1 5704 2402 5796 2418 0 _2543_.vdd
rlabel metal2 5733 2553 5747 2567 0 _2543_.B
rlabel metal2 5773 2553 5787 2567 0 _2543_.A
rlabel metal2 5753 2573 5767 2587 0 _2543_.Y
rlabel metal1 6064 2642 6316 2658 0 _2963_.gnd
rlabel metal1 6064 2402 6316 2418 0 _2963_.vdd
rlabel metal2 6213 2553 6227 2567 0 _2963_.D
rlabel metal2 6173 2553 6187 2567 0 _2963_.CLK
rlabel metal2 6093 2553 6107 2567 0 _2963_.Q
rlabel metal1 5884 2642 6016 2658 0 _2545_.gnd
rlabel metal1 5884 2402 6016 2418 0 _2545_.vdd
rlabel metal2 5993 2553 6007 2567 0 _2545_.A
rlabel metal2 5973 2533 5987 2547 0 _2545_.B
rlabel metal2 5913 2553 5927 2567 0 _2545_.C
rlabel metal2 5953 2553 5967 2567 0 _2545_.Y
rlabel metal2 5933 2533 5947 2547 0 _2545_.D
rlabel metal1 6004 2642 6076 2658 0 _2542_.gnd
rlabel metal1 6004 2402 6076 2418 0 _2542_.vdd
rlabel metal2 6053 2573 6067 2587 0 _2542_.A
rlabel metal2 6033 2533 6047 2547 0 _2542_.Y
rlabel metal1 6304 2642 6436 2658 0 _2766_.gnd
rlabel metal1 6304 2402 6436 2418 0 _2766_.vdd
rlabel metal2 6413 2553 6427 2567 0 _2766_.A
rlabel metal2 6393 2533 6407 2547 0 _2766_.B
rlabel metal2 6333 2553 6347 2567 0 _2766_.C
rlabel metal2 6353 2533 6367 2547 0 _2766_.D
rlabel metal2 6373 2553 6387 2567 0 _2766_.Y
rlabel metal1 6504 2642 6576 2658 0 _2756_.gnd
rlabel metal1 6504 2402 6576 2418 0 _2756_.vdd
rlabel metal2 6513 2573 6527 2587 0 _2756_.A
rlabel metal2 6533 2533 6547 2547 0 _2756_.Y
rlabel metal1 6564 2642 6696 2658 0 _2767_.gnd
rlabel metal1 6564 2402 6696 2418 0 _2767_.vdd
rlabel metal2 6573 2553 6587 2567 0 _2767_.A
rlabel metal2 6593 2533 6607 2547 0 _2767_.B
rlabel metal2 6653 2553 6667 2567 0 _2767_.C
rlabel metal2 6633 2533 6647 2547 0 _2767_.D
rlabel metal2 6613 2553 6627 2567 0 _2767_.Y
rlabel metal1 6424 2642 6516 2658 0 _2668_.gnd
rlabel metal1 6424 2402 6516 2418 0 _2668_.vdd
rlabel metal2 6433 2533 6447 2547 0 _2668_.A
rlabel metal2 6473 2533 6487 2547 0 _2668_.Y
rlabel nsubstratencontact 6724 2412 6724 2412 0 FILL100650x36150.vdd
rlabel metal1 6704 2642 6736 2658 0 FILL100650x36150.gnd
rlabel nsubstratencontact 6704 2412 6704 2412 0 FILL100350x36150.vdd
rlabel metal1 6684 2642 6716 2658 0 FILL100350x36150.gnd
rlabel metal1 144 2642 396 2658 0 _1625_.gnd
rlabel metal1 144 2882 396 2898 0 _1625_.vdd
rlabel metal2 233 2733 247 2747 0 _1625_.D
rlabel metal2 273 2733 287 2747 0 _1625_.CLK
rlabel metal2 353 2733 367 2747 0 _1625_.Q
rlabel metal1 64 2642 156 2658 0 _1593_.gnd
rlabel metal1 64 2882 156 2898 0 _1593_.vdd
rlabel metal2 93 2733 107 2747 0 _1593_.B
rlabel metal2 133 2733 147 2747 0 _1593_.A
rlabel metal2 113 2713 127 2727 0 _1593_.Y
rlabel metal1 4 2642 76 2658 0 _1559_.gnd
rlabel metal1 4 2882 76 2898 0 _1559_.vdd
rlabel metal2 13 2713 27 2727 0 _1559_.A
rlabel metal2 33 2753 47 2767 0 _1559_.Y
rlabel metal1 524 2642 776 2658 0 _1624_.gnd
rlabel metal1 524 2882 776 2898 0 _1624_.vdd
rlabel metal2 613 2733 627 2747 0 _1624_.D
rlabel metal2 653 2733 667 2747 0 _1624_.CLK
rlabel metal2 733 2733 747 2747 0 _1624_.Q
rlabel metal1 444 2642 536 2658 0 _1592_.gnd
rlabel metal1 444 2882 536 2898 0 _1592_.vdd
rlabel metal2 473 2733 487 2747 0 _1592_.B
rlabel metal2 513 2733 527 2747 0 _1592_.A
rlabel metal2 493 2713 507 2727 0 _1592_.Y
rlabel metal1 384 2642 456 2658 0 _1558_.gnd
rlabel metal1 384 2882 456 2898 0 _1558_.vdd
rlabel metal2 393 2713 407 2727 0 _1558_.A
rlabel metal2 413 2753 427 2767 0 _1558_.Y
rlabel metal1 764 2642 856 2658 0 BUFX2_insert23.gnd
rlabel metal1 764 2882 856 2898 0 BUFX2_insert23.vdd
rlabel metal2 833 2733 847 2747 0 BUFX2_insert23.A
rlabel metal2 793 2733 807 2747 0 BUFX2_insert23.Y
rlabel metal1 924 2642 1016 2658 0 _1532_.gnd
rlabel metal1 924 2882 1016 2898 0 _1532_.vdd
rlabel metal2 933 2773 947 2787 0 _1532_.A
rlabel metal2 973 2773 987 2787 0 _1532_.B
rlabel metal2 953 2753 967 2767 0 _1532_.Y
rlabel metal1 1004 2642 1096 2658 0 _1530_.gnd
rlabel metal1 1004 2882 1096 2898 0 _1530_.vdd
rlabel metal2 1013 2773 1027 2787 0 _1530_.A
rlabel metal2 1053 2773 1067 2787 0 _1530_.B
rlabel metal2 1033 2753 1047 2767 0 _1530_.Y
rlabel metal1 844 2642 936 2658 0 _1509_.gnd
rlabel metal1 844 2882 936 2898 0 _1509_.vdd
rlabel metal2 853 2753 867 2767 0 _1509_.A
rlabel metal2 893 2753 907 2767 0 _1509_.Y
rlabel metal1 1084 2642 1156 2658 0 _2248_.gnd
rlabel metal1 1084 2882 1156 2898 0 _2248_.vdd
rlabel metal2 1093 2713 1107 2727 0 _2248_.A
rlabel metal2 1113 2753 1127 2767 0 _2248_.Y
rlabel metal1 1264 2642 1376 2658 0 _2256_.gnd
rlabel metal1 1264 2882 1376 2898 0 _2256_.vdd
rlabel metal2 1353 2753 1367 2767 0 _2256_.A
rlabel metal2 1333 2713 1347 2727 0 _2256_.B
rlabel metal2 1313 2753 1327 2767 0 _2256_.C
rlabel metal2 1293 2733 1307 2747 0 _2256_.Y
rlabel metal1 1144 2642 1276 2658 0 _2257_.gnd
rlabel metal1 1144 2882 1276 2898 0 _2257_.vdd
rlabel metal2 1153 2733 1167 2747 0 _2257_.A
rlabel metal2 1173 2753 1187 2767 0 _2257_.B
rlabel metal2 1233 2733 1247 2747 0 _2257_.C
rlabel metal2 1213 2753 1227 2767 0 _2257_.D
rlabel metal2 1193 2733 1207 2747 0 _2257_.Y
rlabel metal1 1424 2642 1536 2658 0 _2253_.gnd
rlabel metal1 1424 2882 1536 2898 0 _2253_.vdd
rlabel metal2 1513 2733 1527 2747 0 _2253_.A
rlabel metal2 1493 2753 1507 2767 0 _2253_.B
rlabel metal2 1453 2753 1467 2767 0 _2253_.C
rlabel metal2 1473 2733 1487 2747 0 _2253_.Y
rlabel metal1 1524 2642 1616 2658 0 _2255_.gnd
rlabel metal1 1524 2882 1616 2898 0 _2255_.vdd
rlabel metal2 1573 2733 1587 2747 0 _2255_.B
rlabel metal2 1533 2733 1547 2747 0 _2255_.A
rlabel metal2 1553 2713 1567 2727 0 _2255_.Y
rlabel metal1 1364 2642 1436 2658 0 _2254_.gnd
rlabel metal1 1364 2882 1436 2898 0 _2254_.vdd
rlabel metal2 1413 2713 1427 2727 0 _2254_.A
rlabel metal2 1393 2753 1407 2767 0 _2254_.Y
rlabel metal1 1604 2642 1696 2658 0 _2241_.gnd
rlabel metal1 1604 2882 1696 2898 0 _2241_.vdd
rlabel metal2 1613 2773 1627 2787 0 _2241_.A
rlabel metal2 1653 2773 1667 2787 0 _2241_.B
rlabel metal2 1633 2753 1647 2767 0 _2241_.Y
rlabel metal1 1764 2642 1876 2658 0 _2249_.gnd
rlabel metal1 1764 2882 1876 2898 0 _2249_.vdd
rlabel metal2 1853 2733 1867 2747 0 _2249_.A
rlabel metal2 1833 2753 1847 2767 0 _2249_.B
rlabel metal2 1793 2753 1807 2767 0 _2249_.C
rlabel metal2 1813 2733 1827 2747 0 _2249_.Y
rlabel metal1 1684 2642 1776 2658 0 _2243_.gnd
rlabel metal1 1684 2882 1776 2898 0 _2243_.vdd
rlabel metal2 1733 2733 1747 2747 0 _2243_.B
rlabel metal2 1693 2733 1707 2747 0 _2243_.A
rlabel metal2 1713 2713 1727 2727 0 _2243_.Y
rlabel metal1 1864 2642 1976 2658 0 _2244_.gnd
rlabel metal1 1864 2882 1976 2898 0 _2244_.vdd
rlabel metal2 1873 2713 1887 2727 0 _2244_.A
rlabel metal2 1893 2733 1907 2747 0 _2244_.B
rlabel metal2 1933 2753 1947 2767 0 _2244_.Y
rlabel metal1 1964 2642 2076 2658 0 _2502_.gnd
rlabel metal1 1964 2882 2076 2898 0 _2502_.vdd
rlabel metal2 1973 2733 1987 2747 0 _2502_.A
rlabel metal2 1993 2753 2007 2767 0 _2502_.B
rlabel metal2 2033 2753 2047 2767 0 _2502_.C
rlabel metal2 2013 2733 2027 2747 0 _2502_.Y
rlabel metal1 2064 2642 2176 2658 0 _1477_.gnd
rlabel metal1 2064 2882 2176 2898 0 _1477_.vdd
rlabel metal2 2153 2753 2167 2767 0 _1477_.A
rlabel metal2 2133 2713 2147 2727 0 _1477_.B
rlabel metal2 2113 2753 2127 2767 0 _1477_.C
rlabel metal2 2093 2733 2107 2747 0 _1477_.Y
rlabel metal1 2164 2642 2416 2658 0 _1486_.gnd
rlabel metal1 2164 2882 2416 2898 0 _1486_.vdd
rlabel metal2 2253 2733 2267 2747 0 _1486_.D
rlabel metal2 2293 2733 2307 2747 0 _1486_.CLK
rlabel metal2 2373 2733 2387 2747 0 _1486_.Q
rlabel metal1 2404 2642 2496 2658 0 _1476_.gnd
rlabel metal1 2404 2882 2496 2898 0 _1476_.vdd
rlabel metal2 2413 2773 2427 2787 0 _1476_.A
rlabel metal2 2453 2773 2467 2787 0 _1476_.B
rlabel metal2 2433 2753 2447 2767 0 _1476_.Y
rlabel metal1 2604 2642 2856 2658 0 _3018_.gnd
rlabel metal1 2604 2882 2856 2898 0 _3018_.vdd
rlabel metal2 2693 2733 2707 2747 0 _3018_.D
rlabel metal2 2733 2733 2747 2747 0 _3018_.CLK
rlabel metal2 2813 2733 2827 2747 0 _3018_.Q
rlabel metal1 2484 2642 2556 2658 0 _1502_.gnd
rlabel metal1 2484 2882 2556 2898 0 _1502_.vdd
rlabel metal2 2493 2713 2507 2727 0 _1502_.A
rlabel metal2 2513 2753 2527 2767 0 _1502_.Y
rlabel metal1 2544 2642 2616 2658 0 _1475_.gnd
rlabel metal1 2544 2882 2616 2898 0 _1475_.vdd
rlabel metal2 2593 2713 2607 2727 0 _1475_.A
rlabel metal2 2573 2753 2587 2767 0 _1475_.Y
rlabel metal1 2844 2642 2956 2658 0 _2908_.gnd
rlabel metal1 2844 2882 2956 2898 0 _2908_.vdd
rlabel metal2 2853 2733 2867 2747 0 _2908_.A
rlabel metal2 2873 2753 2887 2767 0 _2908_.B
rlabel metal2 2913 2753 2927 2767 0 _2908_.C
rlabel metal2 2893 2733 2907 2747 0 _2908_.Y
rlabel metal1 3044 2642 3296 2658 0 _3010_.gnd
rlabel metal1 3044 2882 3296 2898 0 _3010_.vdd
rlabel metal2 3193 2733 3207 2747 0 _3010_.D
rlabel metal2 3153 2733 3167 2747 0 _3010_.CLK
rlabel metal2 3073 2733 3087 2747 0 _3010_.Q
rlabel metal1 2944 2642 3056 2658 0 _2907_.gnd
rlabel metal1 2944 2882 3056 2898 0 _2907_.vdd
rlabel metal2 3033 2753 3047 2767 0 _2907_.A
rlabel metal2 3013 2713 3027 2727 0 _2907_.B
rlabel metal2 2993 2753 3007 2767 0 _2907_.C
rlabel metal2 2973 2733 2987 2747 0 _2907_.Y
rlabel metal1 3344 2642 3476 2658 0 _2872_.gnd
rlabel metal1 3344 2882 3476 2898 0 _2872_.vdd
rlabel metal2 3353 2733 3367 2747 0 _2872_.A
rlabel metal2 3373 2753 3387 2767 0 _2872_.B
rlabel metal2 3433 2733 3447 2747 0 _2872_.C
rlabel metal2 3393 2733 3407 2747 0 _2872_.Y
rlabel metal2 3413 2753 3427 2767 0 _2872_.D
rlabel metal1 3464 2642 3576 2658 0 _2871_.gnd
rlabel metal1 3464 2882 3576 2898 0 _2871_.vdd
rlabel metal2 3473 2733 3487 2747 0 _2871_.A
rlabel metal2 3493 2753 3507 2767 0 _2871_.B
rlabel metal2 3533 2753 3547 2767 0 _2871_.C
rlabel metal2 3513 2733 3527 2747 0 _2871_.Y
rlabel metal1 3284 2642 3356 2658 0 _2653_.gnd
rlabel metal1 3284 2882 3356 2898 0 _2653_.vdd
rlabel metal2 3293 2713 3307 2727 0 _2653_.A
rlabel metal2 3313 2753 3327 2767 0 _2653_.Y
rlabel metal1 3564 2642 3696 2658 0 _2655_.gnd
rlabel metal1 3564 2882 3696 2898 0 _2655_.vdd
rlabel metal2 3673 2733 3687 2747 0 _2655_.A
rlabel metal2 3653 2753 3667 2767 0 _2655_.B
rlabel metal2 3593 2733 3607 2747 0 _2655_.C
rlabel metal2 3633 2733 3647 2747 0 _2655_.Y
rlabel metal2 3613 2753 3627 2767 0 _2655_.D
rlabel metal1 3684 2642 3796 2658 0 _2860_.gnd
rlabel metal1 3684 2882 3796 2898 0 _2860_.vdd
rlabel metal2 3693 2733 3707 2747 0 _2860_.A
rlabel metal2 3713 2753 3727 2767 0 _2860_.B
rlabel metal2 3753 2753 3767 2767 0 _2860_.C
rlabel metal2 3733 2733 3747 2747 0 _2860_.Y
rlabel metal1 3784 2642 3916 2658 0 _2861_.gnd
rlabel metal1 3784 2882 3916 2898 0 _2861_.vdd
rlabel metal2 3893 2733 3907 2747 0 _2861_.A
rlabel metal2 3873 2753 3887 2767 0 _2861_.B
rlabel metal2 3813 2733 3827 2747 0 _2861_.C
rlabel metal2 3853 2733 3867 2747 0 _2861_.Y
rlabel metal2 3833 2753 3847 2767 0 _2861_.D
rlabel metal1 3964 2642 4056 2658 0 _2859_.gnd
rlabel metal1 3964 2882 4056 2898 0 _2859_.vdd
rlabel metal2 4013 2733 4027 2747 0 _2859_.B
rlabel metal2 3973 2733 3987 2747 0 _2859_.A
rlabel metal2 3993 2713 4007 2727 0 _2859_.Y
rlabel metal1 3904 2642 3976 2658 0 _2858_.gnd
rlabel metal1 3904 2882 3976 2898 0 _2858_.vdd
rlabel metal2 3953 2713 3967 2727 0 _2858_.A
rlabel metal2 3933 2753 3947 2767 0 _2858_.Y
rlabel metal1 4224 2642 4336 2658 0 _2892_.gnd
rlabel metal1 4224 2882 4336 2898 0 _2892_.vdd
rlabel metal2 4233 2733 4247 2747 0 _2892_.A
rlabel metal2 4253 2753 4267 2767 0 _2892_.B
rlabel metal2 4293 2753 4307 2767 0 _2892_.C
rlabel metal2 4273 2733 4287 2747 0 _2892_.Y
rlabel metal1 4044 2642 4136 2658 0 _2894_.gnd
rlabel metal1 4044 2882 4136 2898 0 _2894_.vdd
rlabel metal2 4093 2733 4107 2747 0 _2894_.B
rlabel metal2 4053 2733 4067 2747 0 _2894_.A
rlabel metal2 4073 2713 4087 2727 0 _2894_.Y
rlabel metal1 4124 2642 4236 2658 0 _2895_.gnd
rlabel metal1 4124 2882 4236 2898 0 _2895_.vdd
rlabel metal2 4213 2753 4227 2767 0 _2895_.A
rlabel metal2 4193 2713 4207 2727 0 _2895_.B
rlabel metal2 4173 2753 4187 2767 0 _2895_.C
rlabel metal2 4153 2733 4167 2747 0 _2895_.Y
rlabel metal1 4424 2642 4676 2658 0 _3014_.gnd
rlabel metal1 4424 2882 4676 2898 0 _3014_.vdd
rlabel metal2 4513 2733 4527 2747 0 _3014_.D
rlabel metal2 4553 2733 4567 2747 0 _3014_.CLK
rlabel metal2 4633 2733 4647 2747 0 _3014_.Q
rlabel metal1 4324 2642 4436 2658 0 _2889_.gnd
rlabel metal1 4324 2882 4436 2898 0 _2889_.vdd
rlabel metal2 4413 2753 4427 2767 0 _2889_.A
rlabel metal2 4393 2773 4407 2787 0 _2889_.B
rlabel metal2 4373 2753 4387 2767 0 _2889_.C
rlabel metal2 4353 2773 4367 2787 0 _2889_.Y
rlabel metal1 4804 2642 4916 2658 0 _2875_.gnd
rlabel metal1 4804 2882 4916 2898 0 _2875_.vdd
rlabel metal2 4813 2733 4827 2747 0 _2875_.A
rlabel metal2 4833 2753 4847 2767 0 _2875_.B
rlabel metal2 4873 2753 4887 2767 0 _2875_.C
rlabel metal2 4853 2733 4867 2747 0 _2875_.Y
rlabel metal1 4724 2642 4816 2658 0 _2890_.gnd
rlabel metal1 4724 2882 4816 2898 0 _2890_.vdd
rlabel metal2 4773 2733 4787 2747 0 _2890_.B
rlabel metal2 4733 2733 4747 2747 0 _2890_.A
rlabel metal2 4753 2713 4767 2727 0 _2890_.Y
rlabel metal1 4664 2642 4736 2658 0 _2605_.gnd
rlabel metal1 4664 2882 4736 2898 0 _2605_.vdd
rlabel metal2 4673 2713 4687 2727 0 _2605_.A
rlabel metal2 4693 2753 4707 2767 0 _2605_.Y
rlabel metal1 4984 2642 5116 2658 0 _2876_.gnd
rlabel metal1 4984 2882 5116 2898 0 _2876_.vdd
rlabel metal2 5093 2733 5107 2747 0 _2876_.A
rlabel metal2 5073 2753 5087 2767 0 _2876_.B
rlabel metal2 5013 2733 5027 2747 0 _2876_.C
rlabel metal2 5053 2733 5067 2747 0 _2876_.Y
rlabel metal2 5033 2753 5047 2767 0 _2876_.D
rlabel metal1 4904 2642 4996 2658 0 _2874_.gnd
rlabel metal1 4904 2882 4996 2898 0 _2874_.vdd
rlabel metal2 4933 2733 4947 2747 0 _2874_.B
rlabel metal2 4973 2733 4987 2747 0 _2874_.A
rlabel metal2 4953 2713 4967 2727 0 _2874_.Y
rlabel metal1 5204 2642 5296 2658 0 BUFX2_insert11.gnd
rlabel metal1 5204 2882 5296 2898 0 BUFX2_insert11.vdd
rlabel metal2 5213 2733 5227 2747 0 BUFX2_insert11.A
rlabel metal2 5253 2733 5267 2747 0 BUFX2_insert11.Y
rlabel metal1 5284 2642 5396 2658 0 _2506_.gnd
rlabel metal1 5284 2882 5396 2898 0 _2506_.vdd
rlabel metal2 5293 2733 5307 2747 0 _2506_.A
rlabel metal2 5313 2753 5327 2767 0 _2506_.B
rlabel metal2 5353 2753 5367 2767 0 _2506_.C
rlabel metal2 5333 2733 5347 2747 0 _2506_.Y
rlabel metal1 5104 2642 5216 2658 0 _2911_.gnd
rlabel metal1 5104 2882 5216 2898 0 _2911_.vdd
rlabel metal2 5113 2753 5127 2767 0 _2911_.A
rlabel metal2 5133 2713 5147 2727 0 _2911_.B
rlabel metal2 5153 2753 5167 2767 0 _2911_.C
rlabel metal2 5173 2733 5187 2747 0 _2911_.Y
rlabel metal1 5564 2642 5816 2658 0 _2955_.gnd
rlabel metal1 5564 2882 5816 2898 0 _2955_.vdd
rlabel metal2 5653 2733 5667 2747 0 _2955_.D
rlabel metal2 5693 2733 5707 2747 0 _2955_.CLK
rlabel metal2 5773 2733 5787 2747 0 _2955_.Q
rlabel metal1 5384 2642 5516 2658 0 _2507_.gnd
rlabel metal1 5384 2882 5516 2898 0 _2507_.vdd
rlabel metal2 5493 2733 5507 2747 0 _2507_.A
rlabel metal2 5473 2753 5487 2767 0 _2507_.B
rlabel metal2 5413 2733 5427 2747 0 _2507_.C
rlabel metal2 5453 2733 5467 2747 0 _2507_.Y
rlabel metal2 5433 2753 5447 2767 0 _2507_.D
rlabel metal1 5504 2642 5576 2658 0 _2504_.gnd
rlabel metal1 5504 2882 5576 2898 0 _2504_.vdd
rlabel metal2 5553 2713 5567 2727 0 _2504_.A
rlabel metal2 5533 2753 5547 2767 0 _2504_.Y
rlabel metal1 5804 2642 5936 2658 0 _2664_.gnd
rlabel metal1 5804 2882 5935 2898 0 _2664_.vdd
rlabel metal2 5813 2753 5827 2767 0 _2664_.S
rlabel metal2 5833 2733 5847 2747 0 _2664_.B
rlabel metal2 5873 2753 5887 2767 0 _2664_.Y
rlabel metal2 5893 2733 5907 2747 0 _2664_.A
rlabel metal1 6044 2642 6176 2658 0 _2763_.gnd
rlabel metal1 6044 2882 6175 2898 0 _2763_.vdd
rlabel metal2 6053 2753 6067 2767 0 _2763_.S
rlabel metal2 6073 2733 6087 2747 0 _2763_.B
rlabel metal2 6113 2753 6127 2767 0 _2763_.Y
rlabel metal2 6133 2733 6147 2747 0 _2763_.A
rlabel metal1 5924 2642 6056 2658 0 _2761_.gnd
rlabel metal1 5924 2882 6055 2898 0 _2761_.vdd
rlabel metal2 5933 2753 5947 2767 0 _2761_.S
rlabel metal2 5953 2733 5967 2747 0 _2761_.B
rlabel metal2 5993 2753 6007 2767 0 _2761_.Y
rlabel metal2 6013 2733 6027 2747 0 _2761_.A
rlabel metal1 6264 2642 6356 2658 0 _2547_.gnd
rlabel metal1 6264 2882 6356 2898 0 _2547_.vdd
rlabel metal2 6333 2753 6347 2767 0 _2547_.A
rlabel metal2 6293 2753 6307 2767 0 _2547_.Y
rlabel metal1 6344 2642 6456 2658 0 _1417_.gnd
rlabel metal1 6344 2882 6456 2898 0 _1417_.vdd
rlabel metal2 6353 2733 6367 2747 0 _1417_.A
rlabel metal2 6413 2733 6427 2747 0 _1417_.Y
rlabel metal2 6393 2773 6407 2787 0 _1417_.B
rlabel metal1 6164 2642 6276 2658 0 _1415_.gnd
rlabel metal1 6164 2882 6276 2898 0 _1415_.vdd
rlabel metal2 6253 2733 6267 2747 0 _1415_.A
rlabel metal2 6193 2733 6207 2747 0 _1415_.Y
rlabel metal2 6213 2773 6227 2787 0 _1415_.B
rlabel metal1 6444 2642 6696 2658 0 _2987_.gnd
rlabel metal1 6444 2882 6696 2898 0 _2987_.vdd
rlabel metal2 6593 2733 6607 2747 0 _2987_.D
rlabel metal2 6553 2733 6567 2747 0 _2987_.CLK
rlabel metal2 6473 2733 6487 2747 0 _2987_.Q
rlabel nsubstratencontact 6716 2888 6716 2888 0 FILL100650x39750.vdd
rlabel metal1 6704 2642 6736 2658 0 FILL100650x39750.gnd
rlabel nsubstratencontact 6696 2888 6696 2888 0 FILL100350x39750.vdd
rlabel metal1 6684 2642 6716 2658 0 FILL100350x39750.gnd
rlabel metal1 4 3122 216 3138 0 CLKBUF1_insert34.gnd
rlabel metal1 4 2882 216 2898 0 CLKBUF1_insert34.vdd
rlabel metal2 33 3013 47 3027 0 CLKBUF1_insert34.A
rlabel metal2 173 3013 187 3027 0 CLKBUF1_insert34.Y
rlabel metal1 204 3122 296 3138 0 _3043_.gnd
rlabel metal1 204 2882 296 2898 0 _3043_.vdd
rlabel metal2 273 3033 287 3047 0 _3043_.A
rlabel metal2 233 3033 247 3047 0 _3043_.Y
rlabel metal1 4 3122 96 3138 0 _3038_.gnd
rlabel metal1 4 3362 96 3378 0 _3038_.vdd
rlabel metal2 73 3213 87 3227 0 _3038_.A
rlabel metal2 33 3213 47 3227 0 _3038_.Y
rlabel metal1 84 3122 336 3138 0 _1623_.gnd
rlabel metal1 84 3362 336 3378 0 _1623_.vdd
rlabel metal2 233 3213 247 3227 0 _1623_.D
rlabel metal2 193 3213 207 3227 0 _1623_.CLK
rlabel metal2 113 3213 127 3227 0 _1623_.Q
rlabel metal1 284 3122 536 3138 0 _2395_.gnd
rlabel metal1 284 2882 536 2898 0 _2395_.vdd
rlabel metal2 373 3033 387 3047 0 _2395_.D
rlabel metal2 413 3033 427 3047 0 _2395_.CLK
rlabel metal2 493 3033 507 3047 0 _2395_.Q
rlabel metal1 504 3122 596 3138 0 _1557_.gnd
rlabel metal1 504 3362 596 3378 0 _1557_.vdd
rlabel metal2 573 3253 587 3267 0 _1557_.A
rlabel metal2 533 3253 547 3267 0 _1557_.B
rlabel metal2 553 3233 567 3247 0 _1557_.Y
rlabel metal1 524 3122 616 3138 0 _1556_.gnd
rlabel metal1 524 2882 616 2898 0 _1556_.vdd
rlabel metal2 593 2993 607 3007 0 _1556_.A
rlabel metal2 553 2993 567 3007 0 _1556_.B
rlabel metal2 573 3013 587 3027 0 _1556_.Y
rlabel metal1 324 3122 416 3138 0 _1555_.gnd
rlabel metal1 324 3362 416 3378 0 _1555_.vdd
rlabel metal2 333 3253 347 3267 0 _1555_.A
rlabel metal2 373 3253 387 3267 0 _1555_.B
rlabel metal2 353 3233 367 3247 0 _1555_.Y
rlabel metal1 404 3122 516 3138 0 _1591_.gnd
rlabel metal1 404 3362 516 3378 0 _1591_.vdd
rlabel metal2 493 3233 507 3247 0 _1591_.A
rlabel metal2 473 3193 487 3207 0 _1591_.B
rlabel metal2 453 3233 467 3247 0 _1591_.C
rlabel metal2 433 3213 447 3227 0 _1591_.Y
rlabel metal1 684 3122 796 3138 0 _2351_.gnd
rlabel metal1 684 2882 796 2898 0 _2351_.vdd
rlabel metal2 773 3033 787 3047 0 _2351_.A
rlabel metal2 753 3013 767 3027 0 _2351_.B
rlabel metal2 713 3013 727 3027 0 _2351_.C
rlabel metal2 733 3033 747 3047 0 _2351_.Y
rlabel metal1 584 3122 656 3138 0 _2348_.gnd
rlabel metal1 584 3362 656 3378 0 _2348_.vdd
rlabel metal2 593 3193 607 3207 0 _2348_.A
rlabel metal2 613 3233 627 3247 0 _2348_.Y
rlabel metal1 744 3122 836 3138 0 _2350_.gnd
rlabel metal1 744 3362 836 3378 0 _2350_.vdd
rlabel metal2 753 3253 767 3267 0 _2350_.A
rlabel metal2 793 3253 807 3267 0 _2350_.B
rlabel metal2 773 3233 787 3247 0 _2350_.Y
rlabel metal1 604 3122 696 3138 0 _2346_.gnd
rlabel metal1 604 2882 696 2898 0 _2346_.vdd
rlabel metal2 613 2993 627 3007 0 _2346_.A
rlabel metal2 653 2993 667 3007 0 _2346_.B
rlabel metal2 633 3013 647 3027 0 _2346_.Y
rlabel metal1 784 3122 876 3138 0 _1528_.gnd
rlabel metal1 784 2882 876 2898 0 _1528_.vdd
rlabel metal2 853 2993 867 3007 0 _1528_.A
rlabel metal2 813 2993 827 3007 0 _1528_.B
rlabel metal2 833 3013 847 3027 0 _1528_.Y
rlabel metal1 644 3122 756 3138 0 _2347_.gnd
rlabel metal1 644 3362 756 3378 0 _2347_.vdd
rlabel metal2 653 3233 667 3247 0 _2347_.A
rlabel metal2 673 3253 687 3267 0 _2347_.B
rlabel metal2 693 3233 707 3247 0 _2347_.C
rlabel metal2 713 3253 727 3267 0 _2347_.Y
rlabel metal1 1044 3122 1296 3138 0 _1614_.gnd
rlabel metal1 1044 2882 1296 2898 0 _1614_.vdd
rlabel metal2 1193 3033 1207 3047 0 _1614_.D
rlabel metal2 1153 3033 1167 3047 0 _1614_.CLK
rlabel metal2 1073 3033 1087 3047 0 _1614_.Q
rlabel metal1 824 3122 936 3138 0 _2349_.gnd
rlabel metal1 824 3362 936 3378 0 _2349_.vdd
rlabel metal2 913 3213 927 3227 0 _2349_.A
rlabel metal2 893 3233 907 3247 0 _2349_.B
rlabel metal2 853 3233 867 3247 0 _2349_.C
rlabel metal2 873 3213 887 3227 0 _2349_.Y
rlabel metal1 1064 3122 1176 3138 0 _2344_.gnd
rlabel metal1 1064 3362 1176 3378 0 _2344_.vdd
rlabel metal2 1073 3213 1087 3227 0 _2344_.A
rlabel metal2 1093 3233 1107 3247 0 _2344_.B
rlabel metal2 1133 3233 1147 3247 0 _2344_.C
rlabel metal2 1113 3213 1127 3227 0 _2344_.Y
rlabel metal1 984 3122 1076 3138 0 _2341_.gnd
rlabel metal1 984 3362 1076 3378 0 _2341_.vdd
rlabel metal2 1033 3213 1047 3227 0 _2341_.B
rlabel metal2 993 3213 1007 3227 0 _2341_.A
rlabel metal2 1013 3193 1027 3207 0 _2341_.Y
rlabel metal1 924 3122 996 3138 0 _2342_.gnd
rlabel metal1 924 3362 996 3378 0 _2342_.vdd
rlabel metal2 933 3193 947 3207 0 _2342_.A
rlabel metal2 953 3233 967 3247 0 _2342_.Y
rlabel metal1 864 3122 956 3138 0 _1529_.gnd
rlabel metal1 864 2882 956 2898 0 _1529_.vdd
rlabel metal2 933 2993 947 3007 0 _1529_.A
rlabel metal2 893 2993 907 3007 0 _1529_.B
rlabel metal2 913 3013 927 3027 0 _1529_.Y
rlabel metal1 944 3122 1056 3138 0 _1582_.gnd
rlabel metal1 944 2882 1056 2898 0 _1582_.vdd
rlabel metal2 953 3013 967 3027 0 _1582_.A
rlabel metal2 973 3053 987 3067 0 _1582_.B
rlabel metal2 993 3013 1007 3027 0 _1582_.C
rlabel metal2 1013 3033 1027 3047 0 _1582_.Y
rlabel metal1 1164 3122 1276 3138 0 _2345_.gnd
rlabel metal1 1164 3362 1276 3378 0 _2345_.vdd
rlabel metal2 1173 3213 1187 3227 0 _2345_.A
rlabel metal2 1193 3233 1207 3247 0 _2345_.B
rlabel metal2 1233 3233 1247 3247 0 _2345_.C
rlabel metal2 1213 3213 1227 3227 0 _2345_.Y
rlabel metal1 1264 3122 1356 3138 0 _2336_.gnd
rlabel metal1 1264 3362 1356 3378 0 _2336_.vdd
rlabel metal2 1273 3253 1287 3267 0 _2336_.A
rlabel metal2 1313 3253 1327 3267 0 _2336_.B
rlabel metal2 1293 3233 1307 3247 0 _2336_.Y
rlabel metal1 1284 3122 1376 3138 0 _2236_.gnd
rlabel metal1 1284 2882 1376 2898 0 _2236_.vdd
rlabel metal2 1353 2993 1367 3007 0 _2236_.A
rlabel metal2 1313 2993 1327 3007 0 _2236_.B
rlabel metal2 1333 3013 1347 3027 0 _2236_.Y
rlabel metal1 1344 3122 1596 3138 0 _2394_.gnd
rlabel metal1 1344 3362 1596 3378 0 _2394_.vdd
rlabel metal2 1493 3213 1507 3227 0 _2394_.D
rlabel metal2 1453 3213 1467 3227 0 _2394_.CLK
rlabel metal2 1373 3213 1387 3227 0 _2394_.Q
rlabel metal1 1364 3122 1616 3138 0 _2386_.gnd
rlabel metal1 1364 2882 1616 2898 0 _2386_.vdd
rlabel metal2 1513 3033 1527 3047 0 _2386_.D
rlabel metal2 1473 3033 1487 3047 0 _2386_.CLK
rlabel metal2 1393 3033 1407 3047 0 _2386_.Q
rlabel metal1 1604 3122 1676 3138 0 _2265_.gnd
rlabel metal1 1604 2882 1676 2898 0 _2265_.vdd
rlabel metal2 1653 3053 1667 3067 0 _2265_.A
rlabel metal2 1633 3013 1647 3027 0 _2265_.Y
rlabel metal1 1584 3122 1696 3138 0 _2269_.gnd
rlabel metal1 1584 3362 1696 3378 0 _2269_.vdd
rlabel metal2 1673 3213 1687 3227 0 _2269_.A
rlabel metal2 1613 3213 1627 3227 0 _2269_.Y
rlabel metal2 1633 3253 1647 3267 0 _2269_.B
rlabel metal1 1664 3122 1776 3138 0 _2247_.gnd
rlabel metal1 1664 2882 1776 2898 0 _2247_.vdd
rlabel metal2 1753 3033 1767 3047 0 _2247_.A
rlabel metal2 1733 3013 1747 3027 0 _2247_.B
rlabel metal2 1693 3013 1707 3027 0 _2247_.C
rlabel metal2 1713 3033 1727 3047 0 _2247_.Y
rlabel metal1 1764 3122 1856 3138 0 _2266_.gnd
rlabel metal1 1764 2882 1856 2898 0 _2266_.vdd
rlabel metal2 1793 3033 1807 3047 0 _2266_.B
rlabel metal2 1833 3033 1847 3047 0 _2266_.A
rlabel metal2 1813 3053 1827 3067 0 _2266_.Y
rlabel metal1 1684 3122 1796 3138 0 _2267_.gnd
rlabel metal1 1684 3362 1796 3378 0 _2267_.vdd
rlabel metal2 1773 3233 1787 3247 0 _2267_.A
rlabel metal2 1753 3193 1767 3207 0 _2267_.B
rlabel metal2 1733 3233 1747 3247 0 _2267_.C
rlabel metal2 1713 3213 1727 3227 0 _2267_.Y
rlabel metal1 1784 3122 1896 3138 0 _2268_.gnd
rlabel metal1 1784 3362 1896 3378 0 _2268_.vdd
rlabel metal2 1873 3233 1887 3247 0 _2268_.A
rlabel metal2 1853 3253 1867 3267 0 _2268_.B
rlabel metal2 1833 3233 1847 3247 0 _2268_.C
rlabel metal2 1813 3253 1827 3267 0 _2268_.Y
rlabel metal1 1844 3122 1956 3138 0 _2245_.gnd
rlabel metal1 1844 2882 1956 2898 0 _2245_.vdd
rlabel metal2 1933 3033 1947 3047 0 _2245_.A
rlabel metal2 1873 3033 1887 3047 0 _2245_.Y
rlabel metal2 1893 2993 1907 3007 0 _2245_.B
rlabel metal1 1984 3122 2236 3138 0 _2459_.gnd
rlabel metal1 1984 3362 2236 3378 0 _2459_.vdd
rlabel metal2 2073 3213 2087 3227 0 _2459_.D
rlabel metal2 2113 3213 2127 3227 0 _2459_.CLK
rlabel metal2 2193 3213 2207 3227 0 _2459_.Q
rlabel metal1 1944 3122 2056 3138 0 _2246_.gnd
rlabel metal1 1944 2882 2056 2898 0 _2246_.vdd
rlabel metal2 1953 3033 1967 3047 0 _2246_.A
rlabel metal2 1973 3013 1987 3027 0 _2246_.B
rlabel metal2 2013 3013 2027 3027 0 _2246_.C
rlabel metal2 1993 3033 2007 3047 0 _2246_.Y
rlabel metal1 2044 3122 2156 3138 0 _2456_.gnd
rlabel metal1 2044 2882 2156 2898 0 _2456_.vdd
rlabel metal2 2133 3013 2147 3027 0 _2456_.A
rlabel metal2 2113 3053 2127 3067 0 _2456_.B
rlabel metal2 2093 3013 2107 3027 0 _2456_.C
rlabel metal2 2073 3033 2087 3047 0 _2456_.Y
rlabel metal1 1884 3122 1996 3138 0 _2240_.gnd
rlabel metal1 1884 3362 1996 3378 0 _2240_.vdd
rlabel metal2 1893 3233 1907 3247 0 _2240_.A
rlabel metal2 1913 3193 1927 3207 0 _2240_.B
rlabel metal2 1933 3233 1947 3247 0 _2240_.C
rlabel metal2 1953 3213 1967 3227 0 _2240_.Y
rlabel metal1 2384 3122 2636 3138 0 _2445_.gnd
rlabel metal1 2384 2882 2636 2898 0 _2445_.vdd
rlabel metal2 2473 3033 2487 3047 0 _2445_.D
rlabel metal2 2513 3033 2527 3047 0 _2445_.CLK
rlabel metal2 2593 3033 2607 3047 0 _2445_.Q
rlabel metal1 2384 3122 2476 3138 0 _2457_.gnd
rlabel metal1 2384 3362 2476 3378 0 _2457_.vdd
rlabel metal2 2413 3213 2427 3227 0 _2457_.B
rlabel metal2 2453 3213 2467 3227 0 _2457_.A
rlabel metal2 2433 3193 2447 3207 0 _2457_.Y
rlabel metal1 2304 3122 2396 3138 0 _2438_.gnd
rlabel metal1 2304 3362 2396 3378 0 _2438_.vdd
rlabel metal2 2353 3213 2367 3227 0 _2438_.B
rlabel metal2 2313 3213 2327 3227 0 _2438_.A
rlabel metal2 2333 3193 2347 3207 0 _2438_.Y
rlabel metal1 2224 3122 2296 3138 0 _2450_.gnd
rlabel metal1 2224 2882 2296 2898 0 _2450_.vdd
rlabel metal2 2273 3053 2287 3067 0 _2450_.A
rlabel metal2 2253 3013 2267 3027 0 _2450_.Y
rlabel metal1 2144 3122 2236 3138 0 _2453_.gnd
rlabel metal1 2144 2882 2236 2898 0 _2453_.vdd
rlabel metal2 2153 2993 2167 3007 0 _2453_.A
rlabel metal2 2193 2993 2207 3007 0 _2453_.B
rlabel metal2 2173 3013 2187 3027 0 _2453_.Y
rlabel metal1 2224 3122 2316 3138 0 _2452_.gnd
rlabel metal1 2224 3362 2316 3378 0 _2452_.vdd
rlabel metal2 2233 3253 2247 3267 0 _2452_.A
rlabel metal2 2273 3253 2287 3267 0 _2452_.B
rlabel metal2 2253 3233 2267 3247 0 _2452_.Y
rlabel metal1 2284 3122 2396 3138 0 _2439_.gnd
rlabel metal1 2284 2882 2396 2898 0 _2439_.vdd
rlabel metal2 2293 3033 2307 3047 0 _2439_.A
rlabel metal2 2353 3033 2367 3047 0 _2439_.Y
rlabel metal2 2333 2993 2347 3007 0 _2439_.B
rlabel metal1 2624 3122 2876 3138 0 _2444_.gnd
rlabel metal1 2624 3362 2876 3378 0 _2444_.vdd
rlabel metal2 2713 3213 2727 3227 0 _2444_.D
rlabel metal2 2753 3213 2767 3227 0 _2444_.CLK
rlabel metal2 2833 3213 2847 3227 0 _2444_.Q
rlabel metal1 2464 3122 2576 3138 0 _2458_.gnd
rlabel metal1 2464 3362 2576 3378 0 _2458_.vdd
rlabel metal2 2553 3213 2567 3227 0 _2458_.A
rlabel metal2 2533 3233 2547 3247 0 _2458_.B
rlabel metal2 2493 3233 2507 3247 0 _2458_.C
rlabel metal2 2513 3213 2527 3227 0 _2458_.Y
rlabel metal1 2564 3122 2636 3138 0 _2451_.gnd
rlabel metal1 2564 3362 2636 3378 0 _2451_.vdd
rlabel metal2 2573 3193 2587 3207 0 _2451_.A
rlabel metal2 2593 3233 2607 3247 0 _2451_.Y
rlabel metal1 2624 3122 2696 3138 0 _2425_.gnd
rlabel metal1 2624 2882 2696 2898 0 _2425_.vdd
rlabel metal2 2633 3053 2647 3067 0 _2425_.A
rlabel metal2 2653 3013 2667 3027 0 _2425_.Y
rlabel metal1 2824 3122 2936 3138 0 _2426_.gnd
rlabel metal1 2824 2882 2936 2898 0 _2426_.vdd
rlabel metal2 2913 3033 2927 3047 0 _2426_.A
rlabel metal2 2893 3013 2907 3027 0 _2426_.B
rlabel metal2 2853 3013 2867 3027 0 _2426_.C
rlabel metal2 2873 3033 2887 3047 0 _2426_.Y
rlabel metal1 2684 3122 2776 3138 0 _2437_.gnd
rlabel metal1 2684 2882 2776 2898 0 _2437_.vdd
rlabel metal2 2733 3033 2747 3047 0 _2437_.B
rlabel metal2 2693 3033 2707 3047 0 _2437_.A
rlabel metal2 2713 3053 2727 3067 0 _2437_.Y
rlabel metal1 2764 3122 2836 3138 0 _2406_.gnd
rlabel metal1 2764 2882 2836 2898 0 _2406_.vdd
rlabel metal2 2813 3053 2827 3067 0 _2406_.A
rlabel metal2 2793 3013 2807 3027 0 _2406_.Y
rlabel metal1 2864 3122 2956 3138 0 _2405_.gnd
rlabel metal1 2864 3362 2956 3378 0 _2405_.vdd
rlabel metal2 2873 3253 2887 3267 0 _2405_.A
rlabel metal2 2913 3253 2927 3267 0 _2405_.B
rlabel metal2 2893 3233 2907 3247 0 _2405_.Y
rlabel metal1 2924 3122 2996 3138 0 _2401_.gnd
rlabel metal1 2924 2882 2996 2898 0 _2401_.vdd
rlabel metal2 2933 3013 2947 3027 0 _2401_.A
rlabel metal2 2953 3033 2967 3047 0 _2401_.Y
rlabel metal1 3164 3122 3276 3138 0 _1409_.gnd
rlabel metal1 3164 2882 3276 2898 0 _1409_.vdd
rlabel metal2 3253 3033 3267 3047 0 _1409_.A
rlabel metal2 3233 3013 3247 3027 0 _1409_.B
rlabel metal2 3193 3013 3207 3027 0 _1409_.C
rlabel metal2 3213 3033 3227 3047 0 _1409_.Y
rlabel metal1 3024 3122 3136 3138 0 _1406_.gnd
rlabel metal1 3024 3362 3136 3378 0 _1406_.vdd
rlabel metal2 3113 3213 3127 3227 0 _1406_.A
rlabel metal2 3093 3233 3107 3247 0 _1406_.B
rlabel metal2 3053 3233 3067 3247 0 _1406_.C
rlabel metal2 3073 3213 3087 3227 0 _1406_.Y
rlabel metal1 3204 3122 3276 3138 0 _1404_.gnd
rlabel metal1 3204 3362 3276 3378 0 _1404_.vdd
rlabel metal2 3253 3193 3267 3207 0 _1404_.A
rlabel metal2 3233 3233 3247 3247 0 _1404_.Y
rlabel metal1 3124 3122 3216 3138 0 _1411_.gnd
rlabel metal1 3124 3362 3216 3378 0 _1411_.vdd
rlabel metal2 3193 3253 3207 3267 0 _1411_.A
rlabel metal2 3153 3253 3167 3267 0 _1411_.B
rlabel metal2 3173 3233 3187 3247 0 _1411_.Y
rlabel metal1 3084 3122 3176 3138 0 _1408_.gnd
rlabel metal1 3084 2882 3176 2898 0 _1408_.vdd
rlabel metal2 3153 2993 3167 3007 0 _1408_.A
rlabel metal2 3113 2993 3127 3007 0 _1408_.B
rlabel metal2 3133 3013 3147 3027 0 _1408_.Y
rlabel metal1 2944 3122 3036 3138 0 _1405_.gnd
rlabel metal1 2944 3362 3036 3378 0 _1405_.vdd
rlabel metal2 3013 3253 3027 3267 0 _1405_.A
rlabel metal2 2973 3253 2987 3267 0 _1405_.B
rlabel metal2 2993 3233 3007 3247 0 _1405_.Y
rlabel metal1 2984 3122 3096 3138 0 _2905_.gnd
rlabel metal1 2984 2882 3096 2898 0 _2905_.vdd
rlabel metal2 3073 3013 3087 3027 0 _2905_.A
rlabel metal2 3053 2993 3067 3007 0 _2905_.B
rlabel metal2 3033 3013 3047 3027 0 _2905_.C
rlabel metal2 3013 2993 3027 3007 0 _2905_.Y
rlabel metal1 3264 3122 3376 3138 0 _1412_.gnd
rlabel metal1 3264 3362 3376 3378 0 _1412_.vdd
rlabel metal2 3353 3213 3367 3227 0 _1412_.A
rlabel metal2 3333 3233 3347 3247 0 _1412_.B
rlabel metal2 3293 3233 3307 3247 0 _1412_.C
rlabel metal2 3313 3213 3327 3227 0 _1412_.Y
rlabel metal1 3424 3122 3536 3138 0 _1403_.gnd
rlabel metal1 3424 2882 3536 2898 0 _1403_.vdd
rlabel metal2 3433 3033 3447 3047 0 _1403_.A
rlabel metal2 3453 3013 3467 3027 0 _1403_.B
rlabel metal2 3493 3013 3507 3027 0 _1403_.C
rlabel metal2 3473 3033 3487 3047 0 _1403_.Y
rlabel metal1 3424 3122 3516 3138 0 _2424_.gnd
rlabel metal1 3424 3362 3516 3378 0 _2424_.vdd
rlabel metal2 3453 3213 3467 3227 0 _2424_.B
rlabel metal2 3493 3213 3507 3227 0 _2424_.A
rlabel metal2 3473 3193 3487 3207 0 _2424_.Y
rlabel metal1 3364 3122 3436 3138 0 _2423_.gnd
rlabel metal1 3364 3362 3436 3378 0 _2423_.vdd
rlabel metal2 3373 3193 3387 3207 0 _2423_.A
rlabel metal2 3393 3233 3407 3247 0 _2423_.Y
rlabel metal1 3264 3122 3356 3138 0 _1402_.gnd
rlabel metal1 3264 2882 3356 2898 0 _1402_.vdd
rlabel metal2 3273 2993 3287 3007 0 _1402_.A
rlabel metal2 3313 2993 3327 3007 0 _1402_.B
rlabel metal2 3293 3013 3307 3027 0 _1402_.Y
rlabel metal1 3344 3122 3436 3138 0 _1401_.gnd
rlabel metal1 3344 2882 3436 2898 0 _1401_.vdd
rlabel metal2 3353 2993 3367 3007 0 _1401_.A
rlabel metal2 3393 2993 3407 3007 0 _1401_.B
rlabel metal2 3373 3013 3387 3027 0 _1401_.Y
rlabel metal1 3684 3122 3936 3138 0 _2443_.gnd
rlabel metal1 3684 3362 3936 3378 0 _2443_.vdd
rlabel metal2 3833 3213 3847 3227 0 _2443_.D
rlabel metal2 3793 3213 3807 3227 0 _2443_.CLK
rlabel metal2 3713 3213 3727 3227 0 _2443_.Q
rlabel metal1 3604 3122 3696 3138 0 _2656_.gnd
rlabel metal1 3604 3362 3696 3378 0 _2656_.vdd
rlabel metal2 3633 3213 3647 3227 0 _2656_.B
rlabel metal2 3673 3213 3687 3227 0 _2656_.A
rlabel metal2 3653 3193 3667 3207 0 _2656_.Y
rlabel metal1 3504 3122 3616 3138 0 _2646_.gnd
rlabel metal1 3504 3362 3616 3378 0 _2646_.vdd
rlabel metal2 3593 3233 3607 3247 0 _2646_.A
rlabel metal2 3573 3193 3587 3207 0 _2646_.B
rlabel metal2 3553 3233 3567 3247 0 _2646_.C
rlabel metal2 3533 3213 3547 3227 0 _2646_.Y
rlabel metal1 3624 3122 3756 3138 0 _2652_.gnd
rlabel metal1 3624 2882 3756 2898 0 _2652_.vdd
rlabel metal2 3733 3033 3747 3047 0 _2652_.A
rlabel metal2 3713 3013 3727 3027 0 _2652_.B
rlabel metal2 3653 3033 3667 3047 0 _2652_.C
rlabel metal2 3673 3013 3687 3027 0 _2652_.D
rlabel metal2 3693 3033 3707 3047 0 _2652_.Y
rlabel metal1 3524 3122 3636 3138 0 _1416_.gnd
rlabel metal1 3524 2882 3636 2898 0 _1416_.vdd
rlabel metal2 3533 3033 3547 3047 0 _1416_.A
rlabel metal2 3593 3033 3607 3047 0 _1416_.Y
rlabel metal2 3573 2993 3587 3007 0 _1416_.B
rlabel metal1 3824 3122 4076 3138 0 _3007_.gnd
rlabel metal1 3824 2882 4076 2898 0 _3007_.vdd
rlabel metal2 3913 3033 3927 3047 0 _3007_.D
rlabel metal2 3953 3033 3967 3047 0 _3007_.CLK
rlabel metal2 4033 3033 4047 3047 0 _3007_.Q
rlabel metal1 3924 3122 4056 3138 0 _2623_.gnd
rlabel metal1 3924 3362 4056 3378 0 _2623_.vdd
rlabel metal2 3933 3213 3947 3227 0 _2623_.A
rlabel metal2 3953 3233 3967 3247 0 _2623_.B
rlabel metal2 4013 3213 4027 3227 0 _2623_.C
rlabel metal2 3993 3233 4007 3247 0 _2623_.D
rlabel metal2 3973 3213 3987 3227 0 _2623_.Y
rlabel metal1 3744 3122 3836 3138 0 _2585_.gnd
rlabel metal1 3744 2882 3836 2898 0 _2585_.vdd
rlabel metal2 3813 3013 3827 3027 0 _2585_.A
rlabel metal2 3773 3013 3787 3027 0 _2585_.Y
rlabel metal1 4264 3122 4516 3138 0 _3015_.gnd
rlabel metal1 4264 2882 4516 2898 0 _3015_.vdd
rlabel metal2 4353 3033 4367 3047 0 _3015_.D
rlabel metal2 4393 3033 4407 3047 0 _3015_.CLK
rlabel metal2 4473 3033 4487 3047 0 _3015_.Q
rlabel metal1 4164 3122 4416 3138 0 _2975_.gnd
rlabel metal1 4164 3362 4416 3378 0 _2975_.vdd
rlabel metal2 4253 3213 4267 3227 0 _2975_.D
rlabel metal2 4293 3213 4307 3227 0 _2975_.CLK
rlabel metal2 4373 3213 4387 3227 0 _2975_.Q
rlabel metal1 4064 3122 4176 3138 0 _2896_.gnd
rlabel metal1 4064 2882 4176 2898 0 _2896_.vdd
rlabel metal2 4073 3033 4087 3047 0 _2896_.A
rlabel metal2 4093 3013 4107 3027 0 _2896_.B
rlabel metal2 4133 3013 4147 3027 0 _2896_.C
rlabel metal2 4113 3033 4127 3047 0 _2896_.Y
rlabel metal1 4164 3122 4276 3138 0 _2893_.gnd
rlabel metal1 4164 2882 4276 2898 0 _2893_.vdd
rlabel metal2 4253 3013 4267 3027 0 _2893_.A
rlabel metal2 4233 2993 4247 3007 0 _2893_.B
rlabel metal2 4213 3013 4227 3027 0 _2893_.C
rlabel metal2 4193 2993 4207 3007 0 _2893_.Y
rlabel metal1 4044 3122 4176 3138 0 _2628_.gnd
rlabel metal1 4044 3362 4176 3378 0 _2628_.vdd
rlabel metal2 4153 3213 4167 3227 0 _2628_.A
rlabel metal2 4133 3233 4147 3247 0 _2628_.B
rlabel metal2 4073 3213 4087 3227 0 _2628_.C
rlabel metal2 4093 3233 4107 3247 0 _2628_.D
rlabel metal2 4113 3213 4127 3227 0 _2628_.Y
rlabel metal1 4504 3122 4636 3138 0 _2626_.gnd
rlabel metal1 4504 2882 4636 2898 0 _2626_.vdd
rlabel metal2 4613 3033 4627 3047 0 _2626_.A
rlabel metal2 4593 3013 4607 3027 0 _2626_.B
rlabel metal2 4533 3033 4547 3047 0 _2626_.C
rlabel metal2 4573 3033 4587 3047 0 _2626_.Y
rlabel metal2 4553 3013 4567 3027 0 _2626_.D
rlabel metal1 4404 3122 4496 3138 0 _2627_.gnd
rlabel metal1 4404 3362 4496 3378 0 _2627_.vdd
rlabel metal2 4453 3213 4467 3227 0 _2627_.B
rlabel metal2 4413 3213 4427 3227 0 _2627_.A
rlabel metal2 4433 3193 4447 3207 0 _2627_.Y
rlabel metal1 4484 3122 4616 3138 0 _2618_.gnd
rlabel metal1 4484 3362 4616 3378 0 _2618_.vdd
rlabel metal2 4493 3213 4507 3227 0 _2618_.A
rlabel metal2 4513 3233 4527 3247 0 _2618_.B
rlabel metal2 4573 3213 4587 3227 0 _2618_.C
rlabel metal2 4553 3233 4567 3247 0 _2618_.D
rlabel metal2 4533 3213 4547 3227 0 _2618_.Y
rlabel metal1 4604 3122 4696 3138 0 _2617_.gnd
rlabel metal1 4604 3362 4696 3378 0 _2617_.vdd
rlabel metal2 4653 3213 4667 3227 0 _2617_.B
rlabel metal2 4613 3213 4627 3227 0 _2617_.A
rlabel metal2 4633 3193 4647 3207 0 _2617_.Y
rlabel metal1 4684 3122 4776 3138 0 _2411_.gnd
rlabel metal1 4684 3362 4776 3378 0 _2411_.vdd
rlabel metal2 4733 3213 4747 3227 0 _2411_.B
rlabel metal2 4693 3213 4707 3227 0 _2411_.A
rlabel metal2 4713 3193 4727 3207 0 _2411_.Y
rlabel metal1 4764 3122 4836 3138 0 _2658_.gnd
rlabel metal1 4764 3362 4836 3378 0 _2658_.vdd
rlabel metal2 4773 3193 4787 3207 0 _2658_.A
rlabel metal2 4793 3233 4807 3247 0 _2658_.Y
rlabel metal1 4624 3122 4696 3138 0 _2624_.gnd
rlabel metal1 4624 2882 4696 2898 0 _2624_.vdd
rlabel metal2 4673 3053 4687 3067 0 _2624_.A
rlabel metal2 4653 3013 4667 3027 0 _2624_.Y
rlabel metal1 4804 3122 4936 3138 0 _2613_.gnd
rlabel metal1 4804 2882 4936 2898 0 _2613_.vdd
rlabel metal2 4813 3033 4827 3047 0 _2613_.A
rlabel metal2 4833 3013 4847 3027 0 _2613_.B
rlabel metal2 4893 3033 4907 3047 0 _2613_.C
rlabel metal2 4873 3013 4887 3027 0 _2613_.D
rlabel metal2 4853 3033 4867 3047 0 _2613_.Y
rlabel metal1 4684 3122 4816 3138 0 _2714_.gnd
rlabel metal1 4685 2882 4816 2898 0 _2714_.vdd
rlabel metal2 4793 3013 4807 3027 0 _2714_.S
rlabel metal2 4773 3033 4787 3047 0 _2714_.B
rlabel metal2 4733 3013 4747 3027 0 _2714_.Y
rlabel metal2 4713 3033 4727 3047 0 _2714_.A
rlabel metal1 5044 3122 5296 3138 0 _2440_.gnd
rlabel metal1 5044 3362 5296 3378 0 _2440_.vdd
rlabel metal2 5193 3213 5207 3227 0 _2440_.D
rlabel metal2 5153 3213 5167 3227 0 _2440_.CLK
rlabel metal2 5073 3213 5087 3227 0 _2440_.Q
rlabel metal1 4924 3122 4996 3138 0 _2609_.gnd
rlabel metal1 4924 2882 4996 2898 0 _2609_.vdd
rlabel metal2 4973 3053 4987 3067 0 _2609_.A
rlabel metal2 4953 3013 4967 3027 0 _2609_.Y
rlabel metal1 4944 3122 5056 3138 0 _2606_.gnd
rlabel metal1 4944 3362 5056 3378 0 _2606_.vdd
rlabel metal2 4953 3233 4967 3247 0 _2606_.A
rlabel metal2 4973 3193 4987 3207 0 _2606_.B
rlabel metal2 4993 3233 5007 3247 0 _2606_.C
rlabel metal2 5013 3213 5027 3227 0 _2606_.Y
rlabel metal1 4824 3122 4956 3138 0 _2667_.gnd
rlabel metal1 4824 3362 4956 3378 0 _2667_.vdd
rlabel metal2 4833 3213 4847 3227 0 _2667_.A
rlabel metal2 4853 3233 4867 3247 0 _2667_.B
rlabel metal2 4913 3213 4927 3227 0 _2667_.C
rlabel metal2 4893 3233 4907 3247 0 _2667_.D
rlabel metal2 4873 3213 4887 3227 0 _2667_.Y
rlabel metal1 4984 3122 5116 3138 0 _2662_.gnd
rlabel metal1 4984 2882 5116 2898 0 _2662_.vdd
rlabel metal2 4993 3033 5007 3047 0 _2662_.A
rlabel metal2 5013 3013 5027 3027 0 _2662_.B
rlabel metal2 5073 3033 5087 3047 0 _2662_.C
rlabel metal2 5053 3013 5067 3027 0 _2662_.D
rlabel metal2 5033 3033 5047 3047 0 _2662_.Y
rlabel metal1 5244 3122 5496 3138 0 _3011_.gnd
rlabel metal1 5244 2882 5496 2898 0 _3011_.vdd
rlabel metal2 5333 3033 5347 3047 0 _3011_.D
rlabel metal2 5373 3033 5387 3047 0 _3011_.CLK
rlabel metal2 5453 3033 5467 3047 0 _3011_.Q
rlabel metal1 5164 3122 5256 3138 0 _2666_.gnd
rlabel metal1 5164 2882 5256 2898 0 _2666_.vdd
rlabel metal2 5213 3033 5227 3047 0 _2666_.B
rlabel metal2 5173 3033 5187 3047 0 _2666_.A
rlabel metal2 5193 3053 5207 3067 0 _2666_.Y
rlabel metal1 5104 3122 5176 3138 0 _2873_.gnd
rlabel metal1 5104 2882 5176 2898 0 _2873_.vdd
rlabel metal2 5113 3053 5127 3067 0 _2873_.A
rlabel metal2 5133 3013 5147 3027 0 _2873_.Y
rlabel metal1 5284 3122 5356 3138 0 _2404_.gnd
rlabel metal1 5284 3362 5356 3378 0 _2404_.vdd
rlabel metal2 5333 3193 5347 3207 0 _2404_.A
rlabel metal2 5313 3233 5327 3247 0 _2404_.Y
rlabel metal1 5524 3122 5776 3138 0 _3019_.gnd
rlabel metal1 5524 3362 5776 3378 0 _3019_.vdd
rlabel metal2 5613 3213 5627 3227 0 _3019_.D
rlabel metal2 5653 3213 5667 3227 0 _3019_.CLK
rlabel metal2 5733 3213 5747 3227 0 _3019_.Q
rlabel metal1 5564 3122 5676 3138 0 _2912_.gnd
rlabel metal1 5564 2882 5676 2898 0 _2912_.vdd
rlabel metal2 5573 3033 5587 3047 0 _2912_.A
rlabel metal2 5593 3013 5607 3027 0 _2912_.B
rlabel metal2 5633 3013 5647 3027 0 _2912_.C
rlabel metal2 5613 3033 5627 3047 0 _2912_.Y
rlabel metal1 5484 3122 5576 3138 0 _2910_.gnd
rlabel metal1 5484 2882 5576 2898 0 _2910_.vdd
rlabel metal2 5513 3033 5527 3047 0 _2910_.B
rlabel metal2 5553 3033 5567 3047 0 _2910_.A
rlabel metal2 5533 3053 5547 3067 0 _2910_.Y
rlabel metal1 5464 3122 5536 3138 0 _2419_.gnd
rlabel metal1 5464 3362 5536 3378 0 _2419_.vdd
rlabel metal2 5513 3193 5527 3207 0 _2419_.A
rlabel metal2 5493 3233 5507 3247 0 _2419_.Y
rlabel metal1 5344 3122 5476 3138 0 _2420_.gnd
rlabel metal1 5344 3362 5475 3378 0 _2420_.vdd
rlabel metal2 5353 3233 5367 3247 0 _2420_.S
rlabel metal2 5373 3213 5387 3227 0 _2420_.B
rlabel metal2 5413 3233 5427 3247 0 _2420_.Y
rlabel metal2 5433 3213 5447 3227 0 _2420_.A
rlabel metal1 5764 3122 5896 3138 0 _2665_.gnd
rlabel metal1 5764 2882 5896 2898 0 _2665_.vdd
rlabel metal2 5873 3033 5887 3047 0 _2665_.A
rlabel metal2 5853 3013 5867 3027 0 _2665_.B
rlabel metal2 5793 3033 5807 3047 0 _2665_.C
rlabel metal2 5833 3033 5847 3047 0 _2665_.Y
rlabel metal2 5813 3013 5827 3027 0 _2665_.D
rlabel metal1 5764 3122 5876 3138 0 _2435_.gnd
rlabel metal1 5764 3362 5876 3378 0 _2435_.vdd
rlabel metal2 5853 3213 5867 3227 0 _2435_.A
rlabel metal2 5833 3233 5847 3247 0 _2435_.B
rlabel metal2 5793 3233 5807 3247 0 _2435_.C
rlabel metal2 5813 3213 5827 3227 0 _2435_.Y
rlabel metal1 5864 3122 5936 3138 0 _2421_.gnd
rlabel metal1 5864 3362 5936 3378 0 _2421_.vdd
rlabel metal2 5913 3193 5927 3207 0 _2421_.A
rlabel metal2 5893 3233 5907 3247 0 _2421_.Y
rlabel metal1 5664 3122 5776 3138 0 _2909_.gnd
rlabel metal1 5664 2882 5776 2898 0 _2909_.vdd
rlabel metal2 5753 3013 5767 3027 0 _2909_.A
rlabel metal2 5733 2993 5747 3007 0 _2909_.B
rlabel metal2 5713 3013 5727 3027 0 _2909_.C
rlabel metal2 5693 2993 5707 3007 0 _2909_.Y
rlabel metal1 6024 3122 6136 3138 0 _1738_.gnd
rlabel metal1 6024 3362 6136 3378 0 _1738_.vdd
rlabel metal2 6033 3213 6047 3227 0 _1738_.A
rlabel metal2 6053 3233 6067 3247 0 _1738_.B
rlabel metal2 6093 3233 6107 3247 0 _1738_.C
rlabel metal2 6073 3213 6087 3227 0 _1738_.Y
rlabel metal1 5884 3122 5956 3138 0 _2663_.gnd
rlabel metal1 5884 2882 5956 2898 0 _2663_.vdd
rlabel metal2 5893 3053 5907 3067 0 _2663_.A
rlabel metal2 5913 3013 5927 3027 0 _2663_.Y
rlabel metal1 6124 3122 6216 3138 0 _2410_.gnd
rlabel metal1 6124 3362 6216 3378 0 _2410_.vdd
rlabel metal2 6193 3253 6207 3267 0 _2410_.A
rlabel metal2 6153 3253 6167 3267 0 _2410_.B
rlabel metal2 6173 3233 6187 3247 0 _2410_.Y
rlabel metal1 5924 3122 6036 3138 0 _2433_.gnd
rlabel metal1 5924 3362 6036 3378 0 _2433_.vdd
rlabel metal2 6013 3233 6027 3247 0 _2433_.A
rlabel metal2 5993 3193 6007 3207 0 _2433_.B
rlabel metal2 5973 3233 5987 3247 0 _2433_.C
rlabel metal2 5953 3213 5967 3227 0 _2433_.Y
rlabel metal1 6064 3122 6176 3138 0 _2413_.gnd
rlabel metal1 6064 2882 6176 2898 0 _2413_.vdd
rlabel metal2 6153 3013 6167 3027 0 _2413_.A
rlabel metal2 6133 3053 6147 3067 0 _2413_.B
rlabel metal2 6113 3013 6127 3027 0 _2413_.C
rlabel metal2 6093 3033 6107 3047 0 _2413_.Y
rlabel metal1 5944 3122 6076 3138 0 _2762_.gnd
rlabel metal1 5944 2882 6075 2898 0 _2762_.vdd
rlabel metal2 5953 3013 5967 3027 0 _2762_.S
rlabel metal2 5973 3033 5987 3047 0 _2762_.B
rlabel metal2 6013 3013 6027 3027 0 _2762_.Y
rlabel metal2 6033 3033 6047 3047 0 _2762_.A
rlabel metal1 6384 3122 6496 3138 0 _2436_.gnd
rlabel metal1 6384 3362 6496 3378 0 _2436_.vdd
rlabel metal2 6393 3213 6407 3227 0 _2436_.A
rlabel metal2 6413 3233 6427 3247 0 _2436_.B
rlabel metal2 6453 3233 6467 3247 0 _2436_.C
rlabel metal2 6433 3213 6447 3227 0 _2436_.Y
rlabel metal1 6164 3122 6256 3138 0 _2422_.gnd
rlabel metal1 6164 2882 6256 2898 0 _2422_.vdd
rlabel metal2 6193 3033 6207 3047 0 _2422_.B
rlabel metal2 6233 3033 6247 3047 0 _2422_.A
rlabel metal2 6213 3053 6227 3067 0 _2422_.Y
rlabel metal1 6244 3122 6316 3138 0 _2412_.gnd
rlabel metal1 6244 2882 6316 2898 0 _2412_.vdd
rlabel metal2 6253 3053 6267 3067 0 _2412_.A
rlabel metal2 6273 3013 6287 3027 0 _2412_.Y
rlabel metal1 6304 3122 6396 3138 0 _2403_.gnd
rlabel metal1 6304 3362 6396 3378 0 _2403_.vdd
rlabel metal2 6373 3253 6387 3267 0 _2403_.A
rlabel metal2 6333 3253 6347 3267 0 _2403_.B
rlabel metal2 6353 3233 6367 3247 0 _2403_.Y
rlabel metal1 6204 3122 6316 3138 0 _2402_.gnd
rlabel metal1 6204 3362 6316 3378 0 _2402_.vdd
rlabel metal2 6293 3233 6307 3247 0 _2402_.A
rlabel metal2 6273 3193 6287 3207 0 _2402_.B
rlabel metal2 6253 3233 6267 3247 0 _2402_.C
rlabel metal2 6233 3213 6247 3227 0 _2402_.Y
rlabel metal1 6304 3122 6436 3138 0 _2416_.gnd
rlabel metal1 6304 2882 6436 2898 0 _2416_.vdd
rlabel metal2 6413 3033 6427 3047 0 _2416_.A
rlabel metal2 6393 3013 6407 3027 0 _2416_.B
rlabel metal2 6333 3033 6347 3047 0 _2416_.C
rlabel metal2 6353 3013 6367 3027 0 _2416_.D
rlabel metal2 6373 3033 6387 3047 0 _2416_.Y
rlabel nsubstratencontact 6684 2892 6684 2892 0 FILL100050x43350.vdd
rlabel metal1 6664 3122 6696 3138 0 FILL100050x43350.gnd
rlabel nsubstratencontact 6664 2892 6664 2892 0 FILL99750x43350.vdd
rlabel metal1 6644 3122 6676 3138 0 FILL99750x43350.gnd
rlabel metal1 6484 3122 6736 3138 0 _2449_.gnd
rlabel metal1 6484 3362 6736 3378 0 _2449_.vdd
rlabel metal2 6633 3213 6647 3227 0 _2449_.D
rlabel metal2 6593 3213 6607 3227 0 _2449_.CLK
rlabel metal2 6513 3213 6527 3227 0 _2449_.Q
rlabel metal1 6544 3122 6656 3138 0 _2431_.gnd
rlabel metal1 6544 2882 6656 2898 0 _2431_.vdd
rlabel metal2 6553 3033 6567 3047 0 _2431_.A
rlabel metal2 6573 3013 6587 3027 0 _2431_.B
rlabel metal2 6613 3013 6627 3027 0 _2431_.C
rlabel metal2 6593 3033 6607 3047 0 _2431_.Y
rlabel metal1 6484 3122 6556 3138 0 _2430_.gnd
rlabel metal1 6484 2882 6556 2898 0 _2430_.vdd
rlabel metal2 6493 3053 6507 3067 0 _2430_.A
rlabel metal2 6513 3013 6527 3027 0 _2430_.Y
rlabel metal1 6424 3122 6496 3138 0 _2414_.gnd
rlabel metal1 6424 2882 6496 2898 0 _2414_.vdd
rlabel metal2 6473 3053 6487 3067 0 _2414_.A
rlabel metal2 6453 3013 6467 3027 0 _2414_.Y
rlabel nsubstratencontact 6724 2892 6724 2892 0 FILL100650x43350.vdd
rlabel metal1 6704 3122 6736 3138 0 FILL100650x43350.gnd
rlabel nsubstratencontact 6704 2892 6704 2892 0 FILL100350x43350.vdd
rlabel metal1 6684 3122 6716 3138 0 FILL100350x43350.gnd
rlabel metal1 4 3602 96 3618 0 _3037_.gnd
rlabel metal1 4 3362 96 3378 0 _3037_.vdd
rlabel metal2 73 3513 87 3527 0 _3037_.A
rlabel metal2 33 3513 47 3527 0 _3037_.Y
rlabel metal1 84 3602 336 3618 0 _1622_.gnd
rlabel metal1 84 3362 336 3378 0 _1622_.vdd
rlabel metal2 233 3513 247 3527 0 _1622_.D
rlabel metal2 193 3513 207 3527 0 _1622_.CLK
rlabel metal2 113 3513 127 3527 0 _1622_.Q
rlabel metal1 404 3602 496 3618 0 BUFX2_insert18.gnd
rlabel metal1 404 3362 496 3378 0 BUFX2_insert18.vdd
rlabel metal2 413 3513 427 3527 0 BUFX2_insert18.A
rlabel metal2 453 3513 467 3527 0 BUFX2_insert18.Y
rlabel metal1 324 3602 416 3618 0 _1552_.gnd
rlabel metal1 324 3362 416 3378 0 _1552_.vdd
rlabel metal2 333 3473 347 3487 0 _1552_.A
rlabel metal2 373 3473 387 3487 0 _1552_.B
rlabel metal2 353 3493 367 3507 0 _1552_.Y
rlabel metal1 484 3602 596 3618 0 _1590_.gnd
rlabel metal1 484 3362 596 3378 0 _1590_.vdd
rlabel metal2 573 3493 587 3507 0 _1590_.A
rlabel metal2 553 3533 567 3547 0 _1590_.B
rlabel metal2 533 3493 547 3507 0 _1590_.C
rlabel metal2 513 3513 527 3527 0 _1590_.Y
rlabel metal1 744 3602 836 3618 0 BUFX2_insert19.gnd
rlabel metal1 744 3362 836 3378 0 BUFX2_insert19.vdd
rlabel metal2 753 3513 767 3527 0 BUFX2_insert19.A
rlabel metal2 793 3513 807 3527 0 BUFX2_insert19.Y
rlabel metal1 664 3602 756 3618 0 BUFX2_insert17.gnd
rlabel metal1 664 3362 756 3378 0 BUFX2_insert17.vdd
rlabel metal2 733 3513 747 3527 0 BUFX2_insert17.A
rlabel metal2 693 3513 707 3527 0 BUFX2_insert17.Y
rlabel metal1 584 3602 676 3618 0 _1554_.gnd
rlabel metal1 584 3362 676 3378 0 _1554_.vdd
rlabel metal2 653 3473 667 3487 0 _1554_.A
rlabel metal2 613 3473 627 3487 0 _1554_.B
rlabel metal2 633 3493 647 3507 0 _1554_.Y
rlabel metal1 904 3602 996 3618 0 BUFX2_insert24.gnd
rlabel metal1 904 3362 996 3378 0 BUFX2_insert24.vdd
rlabel metal2 973 3513 987 3527 0 BUFX2_insert24.A
rlabel metal2 933 3513 947 3527 0 BUFX2_insert24.Y
rlabel metal1 1044 3602 1136 3618 0 _3042_.gnd
rlabel metal1 1044 3362 1136 3378 0 _3042_.vdd
rlabel metal2 1113 3513 1127 3527 0 _3042_.A
rlabel metal2 1073 3513 1087 3527 0 _3042_.Y
rlabel metal1 984 3602 1056 3618 0 _2343_.gnd
rlabel metal1 984 3362 1056 3378 0 _2343_.vdd
rlabel metal2 1033 3533 1047 3547 0 _2343_.A
rlabel metal2 1013 3493 1027 3507 0 _2343_.Y
rlabel metal1 824 3602 916 3618 0 _1553_.gnd
rlabel metal1 824 3362 916 3378 0 _1553_.vdd
rlabel metal2 833 3473 847 3487 0 _1553_.A
rlabel metal2 873 3473 887 3487 0 _1553_.B
rlabel metal2 853 3493 867 3507 0 _1553_.Y
rlabel metal1 1124 3602 1216 3618 0 BUFX2_insert1.gnd
rlabel metal1 1124 3362 1216 3378 0 BUFX2_insert1.vdd
rlabel metal2 1193 3513 1207 3527 0 BUFX2_insert1.A
rlabel metal2 1153 3513 1167 3527 0 BUFX2_insert1.Y
rlabel metal1 1204 3602 1456 3618 0 _1613_.gnd
rlabel metal1 1204 3362 1456 3378 0 _1613_.vdd
rlabel metal2 1353 3513 1367 3527 0 _1613_.D
rlabel metal2 1313 3513 1327 3527 0 _1613_.CLK
rlabel metal2 1233 3513 1247 3527 0 _1613_.Q
rlabel metal1 1524 3602 1776 3618 0 _2373_.gnd
rlabel metal1 1524 3362 1776 3378 0 _2373_.vdd
rlabel metal2 1673 3513 1687 3527 0 _2373_.D
rlabel metal2 1633 3513 1647 3527 0 _2373_.CLK
rlabel metal2 1553 3513 1567 3527 0 _2373_.Q
rlabel metal1 1444 3602 1536 3618 0 _1917_.gnd
rlabel metal1 1444 3362 1536 3378 0 _1917_.vdd
rlabel metal2 1473 3513 1487 3527 0 _1917_.B
rlabel metal2 1513 3513 1527 3527 0 _1917_.A
rlabel metal2 1493 3533 1507 3547 0 _1917_.Y
rlabel metal1 1864 3602 1936 3618 0 _2229_.gnd
rlabel metal1 1864 3362 1936 3378 0 _2229_.vdd
rlabel metal2 1913 3533 1927 3547 0 _2229_.A
rlabel metal2 1893 3493 1907 3507 0 _2229_.Y
rlabel metal1 1764 3602 1876 3618 0 _2239_.gnd
rlabel metal1 1764 3362 1876 3378 0 _2239_.vdd
rlabel metal2 1853 3513 1867 3527 0 _2239_.A
rlabel metal2 1793 3513 1807 3527 0 _2239_.Y
rlabel metal2 1813 3473 1827 3487 0 _2239_.B
rlabel metal1 1924 3602 2036 3618 0 _2238_.gnd
rlabel metal1 1924 3362 2036 3378 0 _2238_.vdd
rlabel metal2 2013 3513 2027 3527 0 _2238_.A
rlabel metal2 1993 3493 2007 3507 0 _2238_.B
rlabel metal2 1953 3493 1967 3507 0 _2238_.C
rlabel metal2 1973 3513 1987 3527 0 _2238_.Y
rlabel metal1 2024 3602 2116 3618 0 _2231_.gnd
rlabel metal1 2024 3362 2116 3378 0 _2231_.vdd
rlabel metal2 2073 3513 2087 3527 0 _2231_.B
rlabel metal2 2033 3513 2047 3527 0 _2231_.A
rlabel metal2 2053 3533 2067 3547 0 _2231_.Y
rlabel metal1 2104 3602 2176 3618 0 _2237_.gnd
rlabel metal1 2104 3362 2176 3378 0 _2237_.vdd
rlabel metal2 2153 3533 2167 3547 0 _2237_.A
rlabel metal2 2133 3493 2147 3507 0 _2237_.Y
rlabel metal1 2344 3602 2596 3618 0 _2460_.gnd
rlabel metal1 2344 3362 2596 3378 0 _2460_.vdd
rlabel metal2 2493 3513 2507 3527 0 _2460_.D
rlabel metal2 2453 3513 2467 3527 0 _2460_.CLK
rlabel metal2 2373 3513 2387 3527 0 _2460_.Q
rlabel metal1 2264 3602 2356 3618 0 _2232_.gnd
rlabel metal1 2264 3362 2356 3378 0 _2232_.vdd
rlabel metal2 2293 3513 2307 3527 0 _2232_.B
rlabel metal2 2333 3513 2347 3527 0 _2232_.A
rlabel metal2 2313 3533 2327 3547 0 _2232_.Y
rlabel metal1 2164 3602 2276 3618 0 _2233_.gnd
rlabel metal1 2164 3362 2276 3378 0 _2233_.vdd
rlabel metal2 2253 3513 2267 3527 0 _2233_.A
rlabel metal2 2193 3513 2207 3527 0 _2233_.Y
rlabel metal2 2213 3473 2227 3487 0 _2233_.B
rlabel metal1 2664 3602 2776 3618 0 _1635_.gnd
rlabel metal1 2664 3362 2776 3378 0 _1635_.vdd
rlabel metal2 2673 3513 2687 3527 0 _1635_.A
rlabel metal2 2693 3493 2707 3507 0 _1635_.B
rlabel metal2 2733 3493 2747 3507 0 _1635_.C
rlabel metal2 2713 3513 2727 3527 0 _1635_.Y
rlabel metal1 2584 3602 2676 3618 0 _2455_.gnd
rlabel metal1 2584 3362 2676 3378 0 _2455_.vdd
rlabel metal2 2633 3513 2647 3527 0 _2455_.B
rlabel metal2 2593 3513 2607 3527 0 _2455_.A
rlabel metal2 2613 3533 2627 3547 0 _2455_.Y
rlabel metal1 2904 3602 3016 3618 0 _1640_.gnd
rlabel metal1 2904 3362 3016 3378 0 _1640_.vdd
rlabel metal2 2913 3513 2927 3527 0 _1640_.A
rlabel metal2 2933 3493 2947 3507 0 _1640_.B
rlabel metal2 2973 3493 2987 3507 0 _1640_.C
rlabel metal2 2953 3513 2967 3527 0 _1640_.Y
rlabel metal1 2764 3602 2836 3618 0 _1634_.gnd
rlabel metal1 2764 3362 2836 3378 0 _1634_.vdd
rlabel metal2 2813 3533 2827 3547 0 _1634_.A
rlabel metal2 2793 3493 2807 3507 0 _1634_.Y
rlabel metal1 2824 3602 2916 3618 0 _1639_.gnd
rlabel metal1 2824 3362 2916 3378 0 _1639_.vdd
rlabel metal2 2893 3473 2907 3487 0 _1639_.A
rlabel metal2 2853 3473 2867 3487 0 _1639_.B
rlabel metal2 2873 3493 2887 3507 0 _1639_.Y
rlabel metal1 3004 3602 3116 3618 0 _1648_.gnd
rlabel metal1 3004 3362 3116 3378 0 _1648_.vdd
rlabel metal2 3013 3493 3027 3507 0 _1648_.A
rlabel metal2 3033 3533 3047 3547 0 _1648_.B
rlabel metal2 3053 3493 3067 3507 0 _1648_.C
rlabel metal2 3073 3513 3087 3527 0 _1648_.Y
rlabel metal1 3104 3602 3176 3618 0 _1629_.gnd
rlabel metal1 3104 3362 3176 3378 0 _1629_.vdd
rlabel metal2 3113 3493 3127 3507 0 _1629_.A
rlabel metal2 3133 3513 3147 3527 0 _1629_.Y
rlabel metal1 3164 3602 3296 3618 0 _1649_.gnd
rlabel metal1 3164 3362 3296 3378 0 _1649_.vdd
rlabel metal2 3273 3513 3287 3527 0 _1649_.A
rlabel metal2 3253 3493 3267 3507 0 _1649_.B
rlabel metal2 3193 3513 3207 3527 0 _1649_.C
rlabel metal2 3213 3493 3227 3507 0 _1649_.D
rlabel metal2 3233 3513 3247 3527 0 _1649_.Y
rlabel metal1 3344 3602 3596 3618 0 _1653_.gnd
rlabel metal1 3344 3362 3596 3378 0 _1653_.vdd
rlabel metal2 3493 3513 3507 3527 0 _1653_.D
rlabel metal2 3453 3513 3467 3527 0 _1653_.CLK
rlabel metal2 3373 3513 3387 3527 0 _1653_.Q
rlabel metal1 3284 3602 3356 3618 0 _1647_.gnd
rlabel metal1 3284 3362 3356 3378 0 _1647_.vdd
rlabel metal2 3333 3533 3347 3547 0 _1647_.A
rlabel metal2 3313 3493 3327 3507 0 _1647_.Y
rlabel metal1 3704 3602 3956 3618 0 _2978_.gnd
rlabel metal1 3704 3362 3956 3378 0 _2978_.vdd
rlabel metal2 3853 3513 3867 3527 0 _2978_.D
rlabel metal2 3813 3513 3827 3527 0 _2978_.CLK
rlabel metal2 3733 3513 3747 3527 0 _2978_.Q
rlabel metal1 3584 3602 3716 3618 0 _2647_.gnd
rlabel metal1 3584 3362 3716 3378 0 _2647_.vdd
rlabel metal2 3693 3513 3707 3527 0 _2647_.A
rlabel metal2 3673 3493 3687 3507 0 _2647_.B
rlabel metal2 3613 3513 3627 3527 0 _2647_.C
rlabel metal2 3633 3493 3647 3507 0 _2647_.D
rlabel metal2 3653 3513 3667 3527 0 _2647_.Y
rlabel metal1 4004 3602 4256 3618 0 _2977_.gnd
rlabel metal1 4004 3362 4256 3378 0 _2977_.vdd
rlabel metal2 4153 3513 4167 3527 0 _2977_.D
rlabel metal2 4113 3513 4127 3527 0 _2977_.CLK
rlabel metal2 4033 3513 4047 3527 0 _2977_.Q
rlabel metal1 3944 3602 4016 3618 0 _2638_.gnd
rlabel metal1 3944 3362 4016 3378 0 _2638_.vdd
rlabel metal2 3993 3533 4007 3547 0 _2638_.A
rlabel metal2 3973 3493 3987 3507 0 _2638_.Y
rlabel metal1 4244 3602 4316 3618 0 _2619_.gnd
rlabel metal1 4244 3362 4316 3378 0 _2619_.vdd
rlabel metal2 4293 3533 4307 3547 0 _2619_.A
rlabel metal2 4273 3493 4287 3507 0 _2619_.Y
rlabel metal1 4444 3602 4696 3618 0 _2974_.gnd
rlabel metal1 4444 3362 4696 3378 0 _2974_.vdd
rlabel metal2 4533 3513 4547 3527 0 _2974_.D
rlabel metal2 4573 3513 4587 3527 0 _2974_.CLK
rlabel metal2 4653 3513 4667 3527 0 _2974_.Q
rlabel metal1 4304 3602 4376 3618 0 _1410_.gnd
rlabel metal1 4304 3362 4376 3378 0 _1410_.vdd
rlabel metal2 4353 3533 4367 3547 0 _1410_.A
rlabel metal2 4333 3493 4347 3507 0 _1410_.Y
rlabel metal1 4364 3602 4456 3618 0 _1705_.gnd
rlabel metal1 4364 3362 4456 3378 0 _1705_.vdd
rlabel metal2 4373 3473 4387 3487 0 _1705_.A
rlabel metal2 4413 3473 4427 3487 0 _1705_.B
rlabel metal2 4393 3493 4407 3507 0 _1705_.Y
rlabel metal1 4744 3602 4996 3618 0 _2979_.gnd
rlabel metal1 4744 3362 4996 3378 0 _2979_.vdd
rlabel metal2 4893 3513 4907 3527 0 _2979_.D
rlabel metal2 4853 3513 4867 3527 0 _2979_.CLK
rlabel metal2 4773 3513 4787 3527 0 _2979_.Q
rlabel metal1 4684 3602 4756 3618 0 _2608_.gnd
rlabel metal1 4684 3362 4756 3378 0 _2608_.vdd
rlabel metal2 4733 3533 4747 3547 0 _2608_.A
rlabel metal2 4713 3493 4727 3507 0 _2608_.Y
rlabel metal1 4984 3602 5116 3618 0 _2607_.gnd
rlabel metal1 4984 3362 5116 3378 0 _2607_.vdd
rlabel metal2 5093 3513 5107 3527 0 _2607_.A
rlabel metal2 5073 3493 5087 3507 0 _2607_.B
rlabel metal2 5013 3513 5027 3527 0 _2607_.C
rlabel metal2 5033 3493 5047 3507 0 _2607_.D
rlabel metal2 5053 3513 5067 3527 0 _2607_.Y
rlabel metal1 5164 3602 5416 3618 0 _2973_.gnd
rlabel metal1 5164 3362 5416 3378 0 _2973_.vdd
rlabel metal2 5313 3513 5327 3527 0 _2973_.D
rlabel metal2 5273 3513 5287 3527 0 _2973_.CLK
rlabel metal2 5193 3513 5207 3527 0 _2973_.Q
rlabel metal1 5104 3602 5176 3618 0 _2595_.gnd
rlabel metal1 5104 3362 5176 3378 0 _2595_.vdd
rlabel metal2 5153 3533 5167 3547 0 _2595_.A
rlabel metal2 5133 3493 5147 3507 0 _2595_.Y
rlabel metal1 5404 3602 5656 3618 0 _2442_.gnd
rlabel metal1 5404 3362 5656 3378 0 _2442_.vdd
rlabel metal2 5553 3513 5567 3527 0 _2442_.D
rlabel metal2 5513 3513 5527 3527 0 _2442_.CLK
rlabel metal2 5433 3513 5447 3527 0 _2442_.Q
rlabel metal1 5644 3602 5756 3618 0 _2434_.gnd
rlabel metal1 5644 3362 5756 3378 0 _2434_.vdd
rlabel metal2 5653 3513 5667 3527 0 _2434_.A
rlabel metal2 5673 3493 5687 3507 0 _2434_.B
rlabel metal2 5713 3493 5727 3507 0 _2434_.C
rlabel metal2 5693 3513 5707 3527 0 _2434_.Y
rlabel metal1 5744 3602 5856 3618 0 _2428_.gnd
rlabel metal1 5744 3362 5856 3378 0 _2428_.vdd
rlabel metal2 5753 3513 5767 3527 0 _2428_.A
rlabel metal2 5773 3493 5787 3507 0 _2428_.B
rlabel metal2 5813 3493 5827 3507 0 _2428_.C
rlabel metal2 5793 3513 5807 3527 0 _2428_.Y
rlabel metal1 5844 3602 5916 3618 0 _2408_.gnd
rlabel metal1 5844 3362 5916 3378 0 _2408_.vdd
rlabel metal2 5893 3533 5907 3547 0 _2408_.A
rlabel metal2 5873 3493 5887 3507 0 _2408_.Y
rlabel metal1 6104 3602 6176 3618 0 _2398_.gnd
rlabel metal1 6104 3362 6176 3378 0 _2398_.vdd
rlabel metal2 6153 3533 6167 3547 0 _2398_.A
rlabel metal2 6133 3493 6147 3507 0 _2398_.Y
rlabel metal1 6024 3602 6116 3618 0 _2400_.gnd
rlabel metal1 6024 3362 6116 3378 0 _2400_.vdd
rlabel metal2 6033 3473 6047 3487 0 _2400_.A
rlabel metal2 6073 3473 6087 3487 0 _2400_.B
rlabel metal2 6053 3493 6067 3507 0 _2400_.Y
rlabel metal1 5904 3602 6036 3618 0 _2418_.gnd
rlabel metal1 5904 3362 6036 3378 0 _2418_.vdd
rlabel metal2 6013 3513 6027 3527 0 _2418_.A
rlabel metal2 5993 3493 6007 3507 0 _2418_.B
rlabel metal2 5933 3513 5947 3527 0 _2418_.C
rlabel metal2 5953 3493 5967 3507 0 _2418_.D
rlabel metal2 5973 3513 5987 3527 0 _2418_.Y
rlabel metal1 6404 3602 6656 3618 0 _2448_.gnd
rlabel metal1 6404 3362 6656 3378 0 _2448_.vdd
rlabel metal2 6553 3513 6567 3527 0 _2448_.D
rlabel metal2 6513 3513 6527 3527 0 _2448_.CLK
rlabel metal2 6433 3513 6447 3527 0 _2448_.Q
rlabel metal1 6344 3602 6416 3618 0 _2399_.gnd
rlabel metal1 6344 3362 6416 3378 0 _2399_.vdd
rlabel metal2 6393 3533 6407 3547 0 _2399_.A
rlabel metal2 6373 3493 6387 3507 0 _2399_.Y
rlabel metal1 6164 3362 6356 3378 0 _2409_.vdd
rlabel metal2 6193 3513 6207 3527 0 _2409_.A
rlabel metal2 6233 3493 6247 3507 0 _2409_.B
rlabel metal2 6253 3513 6267 3527 0 _2409_.C
rlabel metal2 6293 3493 6307 3507 0 _2409_.Y
rlabel metal1 6164 3602 6356 3618 0 _2409_.gnd
rlabel nsubstratencontact 6684 3372 6684 3372 0 FILL100050x50550.vdd
rlabel metal1 6664 3602 6696 3618 0 FILL100050x50550.gnd
rlabel nsubstratencontact 6664 3372 6664 3372 0 FILL99750x50550.vdd
rlabel metal1 6644 3602 6676 3618 0 FILL99750x50550.gnd
rlabel nsubstratencontact 6724 3372 6724 3372 0 FILL100650x50550.vdd
rlabel metal1 6704 3602 6736 3618 0 FILL100650x50550.gnd
rlabel nsubstratencontact 6704 3372 6704 3372 0 FILL100350x50550.vdd
rlabel metal1 6684 3602 6716 3618 0 FILL100350x50550.gnd
rlabel metal1 84 3602 176 3618 0 _3036_.gnd
rlabel metal1 84 3842 176 3858 0 _3036_.vdd
rlabel metal2 153 3693 167 3707 0 _3036_.A
rlabel metal2 113 3693 127 3707 0 _3036_.Y
rlabel metal1 4 3602 96 3618 0 _3031_.gnd
rlabel metal1 4 3842 96 3858 0 _3031_.vdd
rlabel metal2 73 3693 87 3707 0 _3031_.A
rlabel metal2 33 3693 47 3707 0 _3031_.Y
rlabel metal1 244 3602 496 3618 0 _1621_.gnd
rlabel metal1 244 3842 496 3858 0 _1621_.vdd
rlabel metal2 393 3693 407 3707 0 _1621_.D
rlabel metal2 353 3693 367 3707 0 _1621_.CLK
rlabel metal2 273 3693 287 3707 0 _1621_.Q
rlabel metal1 164 3602 256 3618 0 _1549_.gnd
rlabel metal1 164 3842 256 3858 0 _1549_.vdd
rlabel metal2 233 3733 247 3747 0 _1549_.A
rlabel metal2 193 3733 207 3747 0 _1549_.B
rlabel metal2 213 3713 227 3727 0 _1549_.Y
rlabel metal1 484 3602 596 3618 0 _1589_.gnd
rlabel metal1 484 3842 596 3858 0 _1589_.vdd
rlabel metal2 573 3713 587 3727 0 _1589_.A
rlabel metal2 553 3673 567 3687 0 _1589_.B
rlabel metal2 533 3713 547 3727 0 _1589_.C
rlabel metal2 513 3693 527 3707 0 _1589_.Y
rlabel metal1 584 3602 676 3618 0 _1551_.gnd
rlabel metal1 584 3842 676 3858 0 _1551_.vdd
rlabel metal2 653 3733 667 3747 0 _1551_.A
rlabel metal2 613 3733 627 3747 0 _1551_.B
rlabel metal2 633 3713 647 3727 0 _1551_.Y
rlabel metal1 664 3602 756 3618 0 _1550_.gnd
rlabel metal1 664 3842 756 3858 0 _1550_.vdd
rlabel metal2 673 3733 687 3747 0 _1550_.A
rlabel metal2 713 3733 727 3747 0 _1550_.B
rlabel metal2 693 3713 707 3727 0 _1550_.Y
rlabel metal1 744 3602 836 3618 0 _1510_.gnd
rlabel metal1 744 3842 836 3858 0 _1510_.vdd
rlabel metal2 813 3733 827 3747 0 _1510_.A
rlabel metal2 773 3733 787 3747 0 _1510_.B
rlabel metal2 793 3713 807 3727 0 _1510_.Y
rlabel metal1 824 3602 1076 3618 0 _1608_.gnd
rlabel metal1 824 3842 1076 3858 0 _1608_.vdd
rlabel metal2 973 3693 987 3707 0 _1608_.D
rlabel metal2 933 3693 947 3707 0 _1608_.CLK
rlabel metal2 853 3693 867 3707 0 _1608_.Q
rlabel metal1 1064 3602 1176 3618 0 _1576_.gnd
rlabel metal1 1064 3842 1176 3858 0 _1576_.vdd
rlabel metal2 1073 3713 1087 3727 0 _1576_.A
rlabel metal2 1093 3673 1107 3687 0 _1576_.B
rlabel metal2 1113 3713 1127 3727 0 _1576_.C
rlabel metal2 1133 3693 1147 3707 0 _1576_.Y
rlabel metal1 1244 3602 1336 3618 0 BUFX2_insert22.gnd
rlabel metal1 1244 3842 1336 3858 0 BUFX2_insert22.vdd
rlabel metal2 1253 3693 1267 3707 0 BUFX2_insert22.A
rlabel metal2 1293 3693 1307 3707 0 BUFX2_insert22.Y
rlabel metal1 1164 3602 1256 3618 0 _1525_.gnd
rlabel metal1 1164 3842 1256 3858 0 _1525_.vdd
rlabel metal2 1233 3733 1247 3747 0 _1525_.A
rlabel metal2 1193 3733 1207 3747 0 _1525_.B
rlabel metal2 1213 3713 1227 3727 0 _1525_.Y
rlabel metal1 1324 3602 1436 3618 0 _1581_.gnd
rlabel metal1 1324 3842 1436 3858 0 _1581_.vdd
rlabel metal2 1413 3713 1427 3727 0 _1581_.A
rlabel metal2 1393 3673 1407 3687 0 _1581_.B
rlabel metal2 1373 3713 1387 3727 0 _1581_.C
rlabel metal2 1353 3693 1367 3707 0 _1581_.Y
rlabel metal1 1584 3602 1676 3618 0 _1980_.gnd
rlabel metal1 1584 3842 1676 3858 0 _1980_.vdd
rlabel metal2 1633 3693 1647 3707 0 _1980_.B
rlabel metal2 1593 3693 1607 3707 0 _1980_.A
rlabel metal2 1613 3673 1627 3687 0 _1980_.Y
rlabel metal1 1424 3602 1516 3618 0 _1527_.gnd
rlabel metal1 1424 3842 1516 3858 0 _1527_.vdd
rlabel metal2 1493 3733 1507 3747 0 _1527_.A
rlabel metal2 1453 3733 1467 3747 0 _1527_.B
rlabel metal2 1473 3713 1487 3727 0 _1527_.Y
rlabel metal1 1504 3602 1596 3618 0 _1526_.gnd
rlabel metal1 1504 3842 1596 3858 0 _1526_.vdd
rlabel metal2 1513 3733 1527 3747 0 _1526_.A
rlabel metal2 1553 3733 1567 3747 0 _1526_.B
rlabel metal2 1533 3713 1547 3727 0 _1526_.Y
rlabel metal1 1664 3602 1916 3618 0 _2385_.gnd
rlabel metal1 1664 3842 1916 3858 0 _2385_.vdd
rlabel metal2 1813 3693 1827 3707 0 _2385_.D
rlabel metal2 1773 3693 1787 3707 0 _2385_.CLK
rlabel metal2 1693 3693 1707 3707 0 _2385_.Q
rlabel metal1 2124 3602 2236 3618 0 _2235_.gnd
rlabel metal1 2124 3842 2236 3858 0 _2235_.vdd
rlabel metal2 2133 3693 2147 3707 0 _2235_.A
rlabel metal2 2153 3713 2167 3727 0 _2235_.B
rlabel metal2 2193 3713 2207 3727 0 _2235_.C
rlabel metal2 2173 3693 2187 3707 0 _2235_.Y
rlabel metal1 1984 3602 2076 3618 0 _2230_.gnd
rlabel metal1 1984 3842 2076 3858 0 _2230_.vdd
rlabel metal2 2033 3693 2047 3707 0 _2230_.B
rlabel metal2 1993 3693 2007 3707 0 _2230_.A
rlabel metal2 2013 3673 2027 3687 0 _2230_.Y
rlabel metal1 2064 3602 2136 3618 0 _2226_.gnd
rlabel metal1 2064 3842 2136 3858 0 _2226_.vdd
rlabel metal2 2073 3673 2087 3687 0 _2226_.A
rlabel metal2 2093 3713 2107 3727 0 _2226_.Y
rlabel metal1 1904 3602 1996 3618 0 _2228_.gnd
rlabel metal1 1904 3842 1996 3858 0 _2228_.vdd
rlabel metal2 1973 3733 1987 3747 0 _2228_.A
rlabel metal2 1933 3733 1947 3747 0 _2228_.B
rlabel metal2 1953 3713 1967 3727 0 _2228_.Y
rlabel metal1 2224 3602 2336 3618 0 _2234_.gnd
rlabel metal1 2224 3842 2336 3858 0 _2234_.vdd
rlabel metal2 2313 3693 2327 3707 0 _2234_.A
rlabel metal2 2293 3713 2307 3727 0 _2234_.B
rlabel metal2 2253 3713 2267 3727 0 _2234_.C
rlabel metal2 2273 3693 2287 3707 0 _2234_.Y
rlabel metal1 2324 3602 2436 3618 0 _2227_.gnd
rlabel metal1 2324 3842 2436 3858 0 _2227_.vdd
rlabel metal2 2413 3713 2427 3727 0 _2227_.A
rlabel metal2 2393 3673 2407 3687 0 _2227_.B
rlabel metal2 2373 3713 2387 3727 0 _2227_.C
rlabel metal2 2353 3693 2367 3707 0 _2227_.Y
rlabel metal1 2544 3602 2656 3618 0 _1633_.gnd
rlabel metal1 2544 3842 2656 3858 0 _1633_.vdd
rlabel metal2 2553 3693 2567 3707 0 _1633_.A
rlabel metal2 2573 3713 2587 3727 0 _1633_.B
rlabel metal2 2613 3713 2627 3727 0 _1633_.C
rlabel metal2 2593 3693 2607 3707 0 _1633_.Y
rlabel metal1 2424 3602 2496 3618 0 _2454_.gnd
rlabel metal1 2424 3842 2496 3858 0 _2454_.vdd
rlabel metal2 2433 3673 2447 3687 0 _2454_.A
rlabel metal2 2453 3713 2467 3727 0 _2454_.Y
rlabel metal1 2484 3602 2556 3618 0 _1631_.gnd
rlabel metal1 2484 3842 2556 3858 0 _1631_.vdd
rlabel metal2 2533 3673 2547 3687 0 _1631_.A
rlabel metal2 2513 3713 2527 3727 0 _1631_.Y
rlabel metal1 2644 3602 2756 3618 0 _1636_.gnd
rlabel metal1 2644 3842 2756 3858 0 _1636_.vdd
rlabel metal2 2653 3713 2667 3727 0 _1636_.A
rlabel metal2 2673 3733 2687 3747 0 _1636_.B
rlabel metal2 2693 3713 2707 3727 0 _1636_.C
rlabel metal2 2713 3733 2727 3747 0 _1636_.Y
rlabel metal1 2884 3602 2996 3618 0 _1641_.gnd
rlabel metal1 2884 3842 2996 3858 0 _1641_.vdd
rlabel metal2 2893 3693 2907 3707 0 _1641_.A
rlabel metal2 2913 3713 2927 3727 0 _1641_.B
rlabel metal2 2953 3713 2967 3727 0 _1641_.C
rlabel metal2 2933 3693 2947 3707 0 _1641_.Y
rlabel metal1 2744 3602 2816 3618 0 _1632_.gnd
rlabel metal1 2744 3842 2816 3858 0 _1632_.vdd
rlabel metal2 2793 3673 2807 3687 0 _1632_.A
rlabel metal2 2773 3713 2787 3727 0 _1632_.Y
rlabel metal1 2804 3602 2896 3618 0 _1645_.gnd
rlabel metal1 2804 3842 2896 3858 0 _1645_.vdd
rlabel metal2 2873 3733 2887 3747 0 _1645_.A
rlabel metal2 2833 3733 2847 3747 0 _1645_.B
rlabel metal2 2853 3713 2867 3727 0 _1645_.Y
rlabel metal1 2984 3602 3096 3618 0 _1642_.gnd
rlabel metal1 2984 3842 3096 3858 0 _1642_.vdd
rlabel metal2 2993 3693 3007 3707 0 _1642_.A
rlabel metal2 3013 3713 3027 3727 0 _1642_.B
rlabel metal2 3053 3713 3067 3727 0 _1642_.C
rlabel metal2 3033 3693 3047 3707 0 _1642_.Y
rlabel metal1 3084 3602 3196 3618 0 _1644_.gnd
rlabel metal1 3084 3842 3196 3858 0 _1644_.vdd
rlabel metal2 3093 3713 3107 3727 0 _1644_.A
rlabel metal2 3113 3673 3127 3687 0 _1644_.B
rlabel metal2 3133 3713 3147 3727 0 _1644_.C
rlabel metal2 3153 3693 3167 3707 0 _1644_.Y
rlabel metal1 3184 3602 3316 3618 0 _1646_.gnd
rlabel metal1 3184 3842 3316 3858 0 _1646_.vdd
rlabel metal2 3293 3693 3307 3707 0 _1646_.A
rlabel metal2 3273 3713 3287 3727 0 _1646_.B
rlabel metal2 3213 3693 3227 3707 0 _1646_.C
rlabel metal2 3233 3713 3247 3727 0 _1646_.D
rlabel metal2 3253 3693 3267 3707 0 _1646_.Y
rlabel metal1 3464 3602 3716 3618 0 _1651_.gnd
rlabel metal1 3464 3842 3716 3858 0 _1651_.vdd
rlabel metal2 3553 3693 3567 3707 0 _1651_.D
rlabel metal2 3593 3693 3607 3707 0 _1651_.CLK
rlabel metal2 3673 3693 3687 3707 0 _1651_.Q
rlabel metal1 3384 3602 3476 3618 0 _1675_.gnd
rlabel metal1 3384 3842 3476 3858 0 _1675_.vdd
rlabel metal2 3453 3733 3467 3747 0 _1675_.A
rlabel metal2 3413 3733 3427 3747 0 _1675_.B
rlabel metal2 3433 3713 3447 3727 0 _1675_.Y
rlabel metal1 3304 3602 3396 3618 0 _1638_.gnd
rlabel metal1 3304 3842 3396 3858 0 _1638_.vdd
rlabel metal2 3373 3733 3387 3747 0 _1638_.A
rlabel metal2 3333 3733 3347 3747 0 _1638_.B
rlabel metal2 3353 3713 3367 3727 0 _1638_.Y
rlabel metal1 3704 3602 3796 3618 0 _1702_.gnd
rlabel metal1 3704 3842 3796 3858 0 _1702_.vdd
rlabel metal2 3773 3733 3787 3747 0 _1702_.A
rlabel metal2 3733 3733 3747 3747 0 _1702_.B
rlabel metal2 3753 3713 3767 3727 0 _1702_.Y
rlabel metal1 3904 3602 3976 3618 0 _2648_.gnd
rlabel metal1 3904 3842 3976 3858 0 _2648_.vdd
rlabel metal2 3913 3673 3927 3687 0 _2648_.A
rlabel metal2 3933 3713 3947 3727 0 _2648_.Y
rlabel metal1 3964 3602 4056 3618 0 _1699_.gnd
rlabel metal1 3964 3842 4056 3858 0 _1699_.vdd
rlabel metal2 3973 3733 3987 3747 0 _1699_.A
rlabel metal2 4013 3733 4027 3747 0 _1699_.B
rlabel metal2 3993 3713 4007 3727 0 _1699_.Y
rlabel metal1 3784 3602 3916 3618 0 _2657_.gnd
rlabel metal1 3784 3842 3916 3858 0 _2657_.vdd
rlabel metal2 3893 3693 3907 3707 0 _2657_.A
rlabel metal2 3873 3713 3887 3727 0 _2657_.B
rlabel metal2 3813 3693 3827 3707 0 _2657_.C
rlabel metal2 3833 3713 3847 3727 0 _2657_.D
rlabel metal2 3853 3693 3867 3707 0 _2657_.Y
rlabel metal1 4144 3602 4396 3618 0 _2976_.gnd
rlabel metal1 4144 3842 4396 3858 0 _2976_.vdd
rlabel metal2 4233 3693 4247 3707 0 _2976_.D
rlabel metal2 4273 3693 4287 3707 0 _2976_.CLK
rlabel metal2 4353 3693 4367 3707 0 _2976_.Q
rlabel metal1 4044 3602 4156 3618 0 _2637_.gnd
rlabel metal1 4044 3842 4156 3858 0 _2637_.vdd
rlabel metal2 4053 3693 4067 3707 0 _2637_.A
rlabel metal2 4073 3713 4087 3727 0 _2637_.B
rlabel metal2 4113 3713 4127 3727 0 _2637_.C
rlabel metal2 4093 3693 4107 3707 0 _2637_.Y
rlabel metal1 4384 3602 4476 3618 0 _2629_.gnd
rlabel metal1 4384 3842 4476 3858 0 _2629_.vdd
rlabel metal2 4393 3733 4407 3747 0 _2629_.A
rlabel metal2 4433 3733 4447 3747 0 _2629_.B
rlabel metal2 4413 3713 4427 3727 0 _2629_.Y
rlabel metal1 4464 3602 4556 3618 0 _1696_.gnd
rlabel metal1 4464 3842 4556 3858 0 _1696_.vdd
rlabel metal2 4533 3733 4547 3747 0 _1696_.A
rlabel metal2 4493 3733 4507 3747 0 _1696_.B
rlabel metal2 4513 3713 4527 3727 0 _1696_.Y
rlabel metal1 4544 3602 4756 3618 0 CLKBUF1_insert27.gnd
rlabel metal1 4544 3842 4756 3858 0 CLKBUF1_insert27.vdd
rlabel metal2 4713 3713 4727 3727 0 CLKBUF1_insert27.A
rlabel metal2 4573 3713 4587 3727 0 CLKBUF1_insert27.Y
rlabel metal1 4744 3602 4996 3618 0 _2972_.gnd
rlabel metal1 4744 3842 4996 3858 0 _2972_.vdd
rlabel metal2 4833 3693 4847 3707 0 _2972_.D
rlabel metal2 4873 3693 4887 3707 0 _2972_.CLK
rlabel metal2 4953 3693 4967 3707 0 _2972_.Q
rlabel metal1 4984 3602 5096 3618 0 _2594_.gnd
rlabel metal1 4984 3842 5096 3858 0 _2594_.vdd
rlabel metal2 4993 3693 5007 3707 0 _2594_.A
rlabel metal2 5013 3713 5027 3727 0 _2594_.B
rlabel metal2 5053 3713 5067 3727 0 _2594_.C
rlabel metal2 5033 3693 5047 3707 0 _2594_.Y
rlabel metal1 5304 3602 5516 3618 0 CLKBUF1_insert26.gnd
rlabel metal1 5304 3842 5516 3858 0 CLKBUF1_insert26.vdd
rlabel metal2 5333 3713 5347 3727 0 CLKBUF1_insert26.A
rlabel metal2 5473 3713 5487 3727 0 CLKBUF1_insert26.Y
rlabel metal1 5244 3602 5316 3618 0 _1407_.gnd
rlabel metal1 5244 3842 5316 3858 0 _1407_.vdd
rlabel metal2 5293 3673 5307 3687 0 _1407_.A
rlabel metal2 5273 3713 5287 3727 0 _1407_.Y
rlabel metal1 5084 3602 5176 3618 0 _2586_.gnd
rlabel metal1 5084 3842 5176 3858 0 _2586_.vdd
rlabel metal2 5153 3733 5167 3747 0 _2586_.A
rlabel metal2 5113 3733 5127 3747 0 _2586_.B
rlabel metal2 5133 3713 5147 3727 0 _2586_.Y
rlabel metal1 5164 3602 5256 3618 0 _1687_.gnd
rlabel metal1 5164 3842 5256 3858 0 _1687_.vdd
rlabel metal2 5233 3733 5247 3747 0 _1687_.A
rlabel metal2 5193 3733 5207 3747 0 _1687_.B
rlabel metal2 5213 3713 5227 3727 0 _1687_.Y
rlabel metal1 5504 3602 5756 3618 0 _2441_.gnd
rlabel metal1 5504 3842 5756 3858 0 _2441_.vdd
rlabel metal2 5653 3693 5667 3707 0 _2441_.D
rlabel metal2 5613 3693 5627 3707 0 _2441_.CLK
rlabel metal2 5533 3693 5547 3707 0 _2441_.Q
rlabel metal1 5744 3602 5816 3618 0 _2397_.gnd
rlabel metal1 5744 3842 5816 3858 0 _2397_.vdd
rlabel metal2 5793 3673 5807 3687 0 _2397_.A
rlabel metal2 5773 3713 5787 3727 0 _2397_.Y
rlabel metal1 5804 3602 5896 3618 0 _2429_.gnd
rlabel metal1 5804 3842 5896 3858 0 _2429_.vdd
rlabel metal2 5813 3733 5827 3747 0 _2429_.A
rlabel metal2 5853 3733 5867 3747 0 _2429_.B
rlabel metal2 5833 3713 5847 3727 0 _2429_.Y
rlabel metal1 6024 3602 6116 3618 0 _2407_.gnd
rlabel metal1 6024 3842 6116 3858 0 _2407_.vdd
rlabel metal2 6073 3693 6087 3707 0 _2407_.B
rlabel metal2 6033 3693 6047 3707 0 _2407_.A
rlabel metal2 6053 3673 6067 3687 0 _2407_.Y
rlabel metal1 6104 3602 6196 3618 0 _2396_.gnd
rlabel metal1 6104 3842 6196 3858 0 _2396_.vdd
rlabel metal2 6133 3693 6147 3707 0 _2396_.B
rlabel metal2 6173 3693 6187 3707 0 _2396_.A
rlabel metal2 6153 3673 6167 3687 0 _2396_.Y
rlabel metal1 5964 3602 6036 3618 0 _2417_.gnd
rlabel metal1 5964 3842 6036 3858 0 _2417_.vdd
rlabel metal2 6013 3673 6027 3687 0 _2417_.A
rlabel metal2 5993 3713 6007 3727 0 _2417_.Y
rlabel metal1 5884 3602 5976 3618 0 _2427_.gnd
rlabel metal1 5884 3842 5976 3858 0 _2427_.vdd
rlabel metal2 5893 3733 5907 3747 0 _2427_.A
rlabel metal2 5933 3733 5947 3747 0 _2427_.B
rlabel metal2 5913 3713 5927 3727 0 _2427_.Y
rlabel metal1 6284 3602 6536 3618 0 _2447_.gnd
rlabel metal1 6284 3842 6536 3858 0 _2447_.vdd
rlabel metal2 6433 3693 6447 3707 0 _2447_.D
rlabel metal2 6393 3693 6407 3707 0 _2447_.CLK
rlabel metal2 6313 3693 6327 3707 0 _2447_.Q
rlabel metal1 6184 3602 6296 3618 0 _2415_.gnd
rlabel metal1 6184 3842 6296 3858 0 _2415_.vdd
rlabel metal2 6193 3713 6207 3727 0 _2415_.A
rlabel metal2 6213 3673 6227 3687 0 _2415_.B
rlabel metal2 6233 3713 6247 3727 0 _2415_.C
rlabel metal2 6253 3693 6267 3707 0 _2415_.Y
rlabel metal1 6524 3602 6636 3618 0 _2432_.gnd
rlabel metal1 6524 3842 6636 3858 0 _2432_.vdd
rlabel metal2 6533 3693 6547 3707 0 _2432_.A
rlabel metal2 6553 3713 6567 3727 0 _2432_.B
rlabel metal2 6593 3713 6607 3727 0 _2432_.C
rlabel metal2 6573 3693 6587 3707 0 _2432_.Y
rlabel metal1 6624 3602 6716 3618 0 _2764_.gnd
rlabel metal1 6624 3842 6716 3858 0 _2764_.vdd
rlabel metal2 6633 3733 6647 3747 0 _2764_.A
rlabel metal2 6673 3733 6687 3747 0 _2764_.B
rlabel metal2 6653 3713 6667 3727 0 _2764_.Y
rlabel nsubstratencontact 6716 3848 6716 3848 0 FILL100650x54150.vdd
rlabel metal1 6704 3602 6736 3618 0 FILL100650x54150.gnd
rlabel metal1 4 4082 96 4098 0 _3035_.gnd
rlabel metal1 4 3842 96 3858 0 _3035_.vdd
rlabel metal2 73 3993 87 4007 0 _3035_.A
rlabel metal2 33 3993 47 4007 0 _3035_.Y
rlabel metal1 84 4082 336 4098 0 _1620_.gnd
rlabel metal1 84 3842 336 3858 0 _1620_.vdd
rlabel metal2 233 3993 247 4007 0 _1620_.D
rlabel metal2 193 3993 207 4007 0 _1620_.CLK
rlabel metal2 113 3993 127 4007 0 _1620_.Q
rlabel metal1 504 4082 596 4098 0 _1548_.gnd
rlabel metal1 504 3842 596 3858 0 _1548_.vdd
rlabel metal2 573 3953 587 3967 0 _1548_.A
rlabel metal2 533 3953 547 3967 0 _1548_.B
rlabel metal2 553 3973 567 3987 0 _1548_.Y
rlabel metal1 324 4082 416 4098 0 _1546_.gnd
rlabel metal1 324 3842 416 3858 0 _1546_.vdd
rlabel metal2 333 3953 347 3967 0 _1546_.A
rlabel metal2 373 3953 387 3967 0 _1546_.B
rlabel metal2 353 3973 367 3987 0 _1546_.Y
rlabel metal1 404 4082 516 4098 0 _1588_.gnd
rlabel metal1 404 3842 516 3858 0 _1588_.vdd
rlabel metal2 493 3973 507 3987 0 _1588_.A
rlabel metal2 473 4013 487 4027 0 _1588_.B
rlabel metal2 453 3973 467 3987 0 _1588_.C
rlabel metal2 433 3993 447 4007 0 _1588_.Y
rlabel metal1 664 4082 756 4098 0 _3041_.gnd
rlabel metal1 664 3842 756 3858 0 _3041_.vdd
rlabel metal2 733 3993 747 4007 0 _3041_.A
rlabel metal2 693 3993 707 4007 0 _3041_.Y
rlabel metal1 744 4082 996 4098 0 _1612_.gnd
rlabel metal1 744 3842 996 3858 0 _1612_.vdd
rlabel metal2 893 3993 907 4007 0 _1612_.D
rlabel metal2 853 3993 867 4007 0 _1612_.CLK
rlabel metal2 773 3993 787 4007 0 _1612_.Q
rlabel metal1 584 4082 676 4098 0 _1547_.gnd
rlabel metal1 584 3842 676 3858 0 _1547_.vdd
rlabel metal2 653 3953 667 3967 0 _1547_.A
rlabel metal2 613 3953 627 3967 0 _1547_.B
rlabel metal2 633 3973 647 3987 0 _1547_.Y
rlabel metal1 1064 4082 1156 4098 0 _1512_.gnd
rlabel metal1 1064 3842 1156 3858 0 _1512_.vdd
rlabel metal2 1073 3953 1087 3967 0 _1512_.A
rlabel metal2 1113 3953 1127 3967 0 _1512_.B
rlabel metal2 1093 3973 1107 3987 0 _1512_.Y
rlabel metal1 984 4082 1076 4098 0 _1511_.gnd
rlabel metal1 984 3842 1076 3858 0 _1511_.vdd
rlabel metal2 1053 3953 1067 3967 0 _1511_.A
rlabel metal2 1013 3953 1027 3967 0 _1511_.B
rlabel metal2 1033 3973 1047 3987 0 _1511_.Y
rlabel metal1 1324 4082 1576 4098 0 _2380_.gnd
rlabel metal1 1324 3842 1576 3858 0 _2380_.vdd
rlabel metal2 1473 3993 1487 4007 0 _2380_.D
rlabel metal2 1433 3993 1447 4007 0 _2380_.CLK
rlabel metal2 1353 3993 1367 4007 0 _2380_.Q
rlabel metal1 1144 4082 1236 4098 0 _1522_.gnd
rlabel metal1 1144 3842 1236 3858 0 _1522_.vdd
rlabel metal2 1153 3953 1167 3967 0 _1522_.A
rlabel metal2 1193 3953 1207 3967 0 _1522_.B
rlabel metal2 1173 3973 1187 3987 0 _1522_.Y
rlabel metal1 1224 4082 1336 4098 0 _1580_.gnd
rlabel metal1 1224 3842 1336 3858 0 _1580_.vdd
rlabel metal2 1313 3973 1327 3987 0 _1580_.A
rlabel metal2 1293 4013 1307 4027 0 _1580_.B
rlabel metal2 1273 3973 1287 3987 0 _1580_.C
rlabel metal2 1253 3993 1267 4007 0 _1580_.Y
rlabel metal1 1564 4082 1656 4098 0 _1524_.gnd
rlabel metal1 1564 3842 1656 3858 0 _1524_.vdd
rlabel metal2 1633 3953 1647 3967 0 _1524_.A
rlabel metal2 1593 3953 1607 3967 0 _1524_.B
rlabel metal2 1613 3973 1627 3987 0 _1524_.Y
rlabel metal1 1644 4082 1736 4098 0 BUFX2_insert3.gnd
rlabel metal1 1644 3842 1736 3858 0 BUFX2_insert3.vdd
rlabel metal2 1653 3993 1667 4007 0 BUFX2_insert3.A
rlabel metal2 1693 3993 1707 4007 0 BUFX2_insert3.Y
rlabel metal1 1804 4082 2056 4098 0 _2384_.gnd
rlabel metal1 1804 3842 2056 3858 0 _2384_.vdd
rlabel metal2 1953 3993 1967 4007 0 _2384_.D
rlabel metal2 1913 3993 1927 4007 0 _2384_.CLK
rlabel metal2 1833 3993 1847 4007 0 _2384_.Q
rlabel metal1 1724 4082 1816 4098 0 _1523_.gnd
rlabel metal1 1724 3842 1816 3858 0 _1523_.vdd
rlabel metal2 1733 3953 1747 3967 0 _1523_.A
rlabel metal2 1773 3953 1787 3967 0 _1523_.B
rlabel metal2 1753 3973 1767 3987 0 _1523_.Y
rlabel metal1 2124 4082 2236 4098 0 _2225_.gnd
rlabel metal1 2124 3842 2236 3858 0 _2225_.vdd
rlabel metal2 2213 3993 2227 4007 0 _2225_.A
rlabel metal2 2193 3973 2207 3987 0 _2225_.B
rlabel metal2 2153 3973 2167 3987 0 _2225_.C
rlabel metal2 2173 3993 2187 4007 0 _2225_.Y
rlabel metal1 2044 4082 2136 4098 0 _2214_.gnd
rlabel metal1 2044 3842 2136 3858 0 _2214_.vdd
rlabel metal2 2053 3953 2067 3967 0 _2214_.A
rlabel metal2 2093 3953 2107 3967 0 _2214_.B
rlabel metal2 2073 3973 2087 3987 0 _2214_.Y
rlabel metal1 2384 4082 2456 4098 0 _2220_.gnd
rlabel metal1 2384 3842 2456 3858 0 _2220_.vdd
rlabel metal2 2433 4013 2447 4027 0 _2220_.A
rlabel metal2 2413 3973 2427 3987 0 _2220_.Y
rlabel metal1 2304 4082 2396 4098 0 _2224_.gnd
rlabel metal1 2304 3842 2396 3858 0 _2224_.vdd
rlabel metal2 2313 3953 2327 3967 0 _2224_.A
rlabel metal2 2353 3953 2367 3967 0 _2224_.B
rlabel metal2 2333 3973 2347 3987 0 _2224_.Y
rlabel metal1 2224 4082 2316 4098 0 _2223_.gnd
rlabel metal1 2224 3842 2316 3858 0 _2223_.vdd
rlabel metal2 2293 3953 2307 3967 0 _2223_.A
rlabel metal2 2253 3953 2267 3967 0 _2223_.B
rlabel metal2 2273 3973 2287 3987 0 _2223_.Y
rlabel metal1 2444 4082 2556 4098 0 _2221_.gnd
rlabel metal1 2444 3842 2556 3858 0 _2221_.vdd
rlabel metal2 2533 3993 2547 4007 0 _2221_.A
rlabel metal2 2513 3973 2527 3987 0 _2221_.B
rlabel metal2 2473 3973 2487 3987 0 _2221_.C
rlabel metal2 2493 3993 2507 4007 0 _2221_.Y
rlabel metal1 2544 4082 2636 4098 0 _2222_.gnd
rlabel metal1 2544 3842 2636 3858 0 _2222_.vdd
rlabel metal2 2593 3993 2607 4007 0 _2222_.B
rlabel metal2 2553 3993 2567 4007 0 _2222_.A
rlabel metal2 2573 4013 2587 4027 0 _2222_.Y
rlabel metal1 2624 4082 2716 4098 0 _2216_.gnd
rlabel metal1 2624 3842 2716 3858 0 _2216_.vdd
rlabel metal2 2653 3993 2667 4007 0 _2216_.B
rlabel metal2 2693 3993 2707 4007 0 _2216_.A
rlabel metal2 2673 4013 2687 4027 0 _2216_.Y
rlabel metal1 2904 4082 2996 4098 0 _2208_.gnd
rlabel metal1 2904 3842 2996 3858 0 _2208_.vdd
rlabel metal2 2953 3993 2967 4007 0 _2208_.B
rlabel metal2 2913 3993 2927 4007 0 _2208_.A
rlabel metal2 2933 4013 2947 4027 0 _2208_.Y
rlabel metal1 2704 4082 2776 4098 0 _2215_.gnd
rlabel metal1 2704 3842 2776 3858 0 _2215_.vdd
rlabel metal2 2713 4013 2727 4027 0 _2215_.A
rlabel metal2 2733 3973 2747 3987 0 _2215_.Y
rlabel metal1 2764 4082 2836 4098 0 _2204_.gnd
rlabel metal1 2764 3842 2836 3858 0 _2204_.vdd
rlabel metal2 2813 4013 2827 4027 0 _2204_.A
rlabel metal2 2793 3973 2807 3987 0 _2204_.Y
rlabel metal1 2824 4082 2916 4098 0 _2209_.gnd
rlabel metal1 2824 3842 2916 3858 0 _2209_.vdd
rlabel metal2 2893 3953 2907 3967 0 _2209_.A
rlabel metal2 2853 3953 2867 3967 0 _2209_.B
rlabel metal2 2873 3973 2887 3987 0 _2209_.Y
rlabel metal1 2984 4082 3096 4098 0 _2219_.gnd
rlabel metal1 2984 3842 3096 3858 0 _2219_.vdd
rlabel metal2 2993 3993 3007 4007 0 _2219_.A
rlabel metal2 3013 3973 3027 3987 0 _2219_.B
rlabel metal2 3053 3973 3067 3987 0 _2219_.C
rlabel metal2 3033 3993 3047 4007 0 _2219_.Y
rlabel metal1 3144 4082 3236 4098 0 _2207_.gnd
rlabel metal1 3144 3842 3236 3858 0 _2207_.vdd
rlabel metal2 3193 3993 3207 4007 0 _2207_.B
rlabel metal2 3153 3993 3167 4007 0 _2207_.A
rlabel metal2 3173 4013 3187 4027 0 _2207_.Y
rlabel metal1 3084 4082 3156 4098 0 _2218_.gnd
rlabel metal1 3084 3842 3156 3858 0 _2218_.vdd
rlabel metal2 3093 4013 3107 4027 0 _2218_.A
rlabel metal2 3113 3973 3127 3987 0 _2218_.Y
rlabel metal1 3384 4082 3636 4098 0 _1650_.gnd
rlabel metal1 3384 3842 3636 3858 0 _1650_.vdd
rlabel metal2 3473 3993 3487 4007 0 _1650_.D
rlabel metal2 3513 3993 3527 4007 0 _1650_.CLK
rlabel metal2 3593 3993 3607 4007 0 _1650_.Q
rlabel metal1 3224 4082 3316 4098 0 _1637_.gnd
rlabel metal1 3224 3842 3316 3858 0 _1637_.vdd
rlabel metal2 3293 3953 3307 3967 0 _1637_.A
rlabel metal2 3253 3953 3267 3967 0 _1637_.B
rlabel metal2 3273 3973 3287 3987 0 _1637_.Y
rlabel metal1 3304 4082 3396 4098 0 _1630_.gnd
rlabel metal1 3304 3842 3396 3858 0 _1630_.vdd
rlabel metal2 3373 3953 3387 3967 0 _1630_.A
rlabel metal2 3333 3953 3347 3967 0 _1630_.B
rlabel metal2 3353 3973 3367 3987 0 _1630_.Y
rlabel metal1 3684 4082 3936 4098 0 _1652_.gnd
rlabel metal1 3684 3842 3936 3858 0 _1652_.vdd
rlabel metal2 3773 3993 3787 4007 0 _1652_.D
rlabel metal2 3813 3993 3827 4007 0 _1652_.CLK
rlabel metal2 3893 3993 3907 4007 0 _1652_.Q
rlabel metal1 3624 4082 3696 4098 0 _1643_.gnd
rlabel metal1 3624 3842 3696 3858 0 _1643_.vdd
rlabel metal2 3673 4013 3687 4027 0 _1643_.A
rlabel metal2 3653 3973 3667 3987 0 _1643_.Y
rlabel metal1 3924 4082 4036 4098 0 _1795_.gnd
rlabel metal1 3924 3842 4036 3858 0 _1795_.vdd
rlabel metal2 4013 3973 4027 3987 0 _1795_.A
rlabel metal2 3993 3953 4007 3967 0 _1795_.B
rlabel metal2 3973 3973 3987 3987 0 _1795_.C
rlabel metal2 3953 3953 3967 3967 0 _1795_.Y
rlabel metal1 4104 4082 4216 4098 0 _1791_.gnd
rlabel metal1 4104 3842 4216 3858 0 _1791_.vdd
rlabel metal2 4193 3993 4207 4007 0 _1791_.A
rlabel metal2 4173 3973 4187 3987 0 _1791_.B
rlabel metal2 4133 3973 4147 3987 0 _1791_.C
rlabel metal2 4153 3993 4167 4007 0 _1791_.Y
rlabel metal1 4204 4082 4296 4098 0 _1793_.gnd
rlabel metal1 4204 3842 4296 3858 0 _1793_.vdd
rlabel metal2 4253 3993 4267 4007 0 _1793_.B
rlabel metal2 4213 3993 4227 4007 0 _1793_.A
rlabel metal2 4233 4013 4247 4027 0 _1793_.Y
rlabel metal1 4024 4082 4116 4098 0 _1794_.gnd
rlabel metal1 4024 3842 4116 3858 0 _1794_.vdd
rlabel metal2 4033 3953 4047 3967 0 _1794_.A
rlabel metal2 4073 3953 4087 3967 0 _1794_.B
rlabel metal2 4053 3973 4067 3987 0 _1794_.Y
rlabel metal1 4524 4082 4776 4098 0 _2353_.gnd
rlabel metal1 4524 3842 4776 3858 0 _2353_.vdd
rlabel metal2 4613 3993 4627 4007 0 _2353_.D
rlabel metal2 4653 3993 4667 4007 0 _2353_.CLK
rlabel metal2 4733 3993 4747 4007 0 _2353_.Q
rlabel metal1 4424 4082 4536 4098 0 _1670_.gnd
rlabel metal1 4424 3842 4536 3858 0 _1670_.vdd
rlabel metal2 4513 3993 4527 4007 0 _1670_.A
rlabel metal2 4493 3973 4507 3987 0 _1670_.B
rlabel metal2 4453 3973 4467 3987 0 _1670_.C
rlabel metal2 4473 3993 4487 4007 0 _1670_.Y
rlabel metal1 4284 4082 4356 4098 0 _1790_.gnd
rlabel metal1 4284 3842 4356 3858 0 _1790_.vdd
rlabel metal2 4333 4013 4347 4027 0 _1790_.A
rlabel metal2 4313 3973 4327 3987 0 _1790_.Y
rlabel metal1 4344 4082 4436 4098 0 _1669_.gnd
rlabel metal1 4344 3842 4436 3858 0 _1669_.vdd
rlabel metal2 4413 3953 4427 3967 0 _1669_.A
rlabel metal2 4373 3953 4387 3967 0 _1669_.B
rlabel metal2 4393 3973 4407 3987 0 _1669_.Y
rlabel metal1 4764 4082 4856 4098 0 _1690_.gnd
rlabel metal1 4764 3842 4856 3858 0 _1690_.vdd
rlabel metal2 4833 3953 4847 3967 0 _1690_.A
rlabel metal2 4793 3953 4807 3967 0 _1690_.B
rlabel metal2 4813 3973 4827 3987 0 _1690_.Y
rlabel metal1 4944 4082 5196 4098 0 _2360_.gnd
rlabel metal1 4944 3842 5196 3858 0 _2360_.vdd
rlabel metal2 5033 3993 5047 4007 0 _2360_.D
rlabel metal2 5073 3993 5087 4007 0 _2360_.CLK
rlabel metal2 5153 3993 5167 4007 0 _2360_.Q
rlabel metal1 4844 4082 4956 4098 0 _1691_.gnd
rlabel metal1 4844 3842 4956 3858 0 _1691_.vdd
rlabel metal2 4933 3993 4947 4007 0 _1691_.A
rlabel metal2 4913 3973 4927 3987 0 _1691_.B
rlabel metal2 4873 3973 4887 3987 0 _1691_.C
rlabel metal2 4893 3993 4907 4007 0 _1691_.Y
rlabel metal1 5264 4082 5376 4098 0 _1688_.gnd
rlabel metal1 5264 3842 5376 3858 0 _1688_.vdd
rlabel metal2 5353 3993 5367 4007 0 _1688_.A
rlabel metal2 5333 3973 5347 3987 0 _1688_.B
rlabel metal2 5293 3973 5307 3987 0 _1688_.C
rlabel metal2 5313 3993 5327 4007 0 _1688_.Y
rlabel metal1 5184 4082 5276 4098 0 _1693_.gnd
rlabel metal1 5184 3842 5276 3858 0 _1693_.vdd
rlabel metal2 5253 3953 5267 3967 0 _1693_.A
rlabel metal2 5213 3953 5227 3967 0 _1693_.B
rlabel metal2 5233 3973 5247 3987 0 _1693_.Y
rlabel metal1 5604 4082 5856 4098 0 _2359_.gnd
rlabel metal1 5604 3842 5856 3858 0 _2359_.vdd
rlabel metal2 5693 3993 5707 4007 0 _2359_.D
rlabel metal2 5733 3993 5747 4007 0 _2359_.CLK
rlabel metal2 5813 3993 5827 4007 0 _2359_.Q
rlabel metal1 5444 4082 5556 4098 0 _1685_.gnd
rlabel metal1 5444 3842 5556 3858 0 _1685_.vdd
rlabel metal2 5453 3993 5467 4007 0 _1685_.A
rlabel metal2 5473 3973 5487 3987 0 _1685_.B
rlabel metal2 5513 3973 5527 3987 0 _1685_.C
rlabel metal2 5493 3993 5507 4007 0 _1685_.Y
rlabel metal1 5544 4082 5616 4098 0 _1686_.gnd
rlabel metal1 5544 3842 5616 3858 0 _1686_.vdd
rlabel metal2 5593 4013 5607 4027 0 _1686_.A
rlabel metal2 5573 3973 5587 3987 0 _1686_.Y
rlabel metal1 5364 4082 5456 4098 0 _1684_.gnd
rlabel metal1 5364 3842 5456 3858 0 _1684_.vdd
rlabel metal2 5433 3953 5447 3967 0 _1684_.A
rlabel metal2 5393 3953 5407 3967 0 _1684_.B
rlabel metal2 5413 3973 5427 3987 0 _1684_.Y
rlabel metal1 5844 4082 5916 4098 0 _1734_.gnd
rlabel metal1 5844 3842 5916 3858 0 _1734_.vdd
rlabel metal2 5853 4013 5867 4027 0 _1734_.A
rlabel metal2 5873 3973 5887 3987 0 _1734_.Y
rlabel metal1 6004 4082 6256 4098 0 _2358_.gnd
rlabel metal1 6004 3842 6256 3858 0 _2358_.vdd
rlabel metal2 6153 3993 6167 4007 0 _2358_.D
rlabel metal2 6113 3993 6127 4007 0 _2358_.CLK
rlabel metal2 6033 3993 6047 4007 0 _2358_.Q
rlabel metal1 5904 4082 6016 4098 0 _1739_.gnd
rlabel metal1 5904 3842 6016 3858 0 _1739_.vdd
rlabel metal2 5993 3973 6007 3987 0 _1739_.A
rlabel metal2 5973 3953 5987 3967 0 _1739_.B
rlabel metal2 5953 3973 5967 3987 0 _1739_.C
rlabel metal2 5933 3953 5947 3967 0 _1739_.Y
rlabel metal1 6244 4082 6496 4098 0 _2446_.gnd
rlabel metal1 6244 3842 6496 3858 0 _2446_.vdd
rlabel metal2 6393 3993 6407 4007 0 _2446_.D
rlabel metal2 6353 3993 6367 4007 0 _2446_.CLK
rlabel metal2 6273 3993 6287 4007 0 _2446_.Q
rlabel metal1 6484 4082 6736 4098 0 _2982_.gnd
rlabel metal1 6484 3842 6736 3858 0 _2982_.vdd
rlabel metal2 6633 3993 6647 4007 0 _2982_.D
rlabel metal2 6593 3993 6607 4007 0 _2982_.CLK
rlabel metal2 6513 3993 6527 4007 0 _2982_.Q
rlabel metal1 4 4082 96 4098 0 _3040_.gnd
rlabel metal1 4 4322 96 4338 0 _3040_.vdd
rlabel metal2 73 4173 87 4187 0 _3040_.A
rlabel metal2 33 4173 47 4187 0 _3040_.Y
rlabel metal1 184 4082 296 4098 0 _2325_.gnd
rlabel metal1 184 4322 296 4338 0 _2325_.vdd
rlabel metal2 193 4173 207 4187 0 _2325_.A
rlabel metal2 213 4193 227 4207 0 _2325_.B
rlabel metal2 253 4193 267 4207 0 _2325_.C
rlabel metal2 233 4173 247 4187 0 _2325_.Y
rlabel metal1 84 4082 196 4098 0 _2324_.gnd
rlabel metal1 84 4322 196 4338 0 _2324_.vdd
rlabel metal2 173 4173 187 4187 0 _2324_.A
rlabel metal2 153 4193 167 4207 0 _2324_.B
rlabel metal2 113 4193 127 4207 0 _2324_.C
rlabel metal2 133 4173 147 4187 0 _2324_.Y
rlabel metal1 284 4082 536 4098 0 _2392_.gnd
rlabel metal1 284 4322 536 4338 0 _2392_.vdd
rlabel metal2 373 4173 387 4187 0 _2392_.D
rlabel metal2 413 4173 427 4187 0 _2392_.CLK
rlabel metal2 493 4173 507 4187 0 _2392_.Q
rlabel metal1 524 4082 616 4098 0 _2308_.gnd
rlabel metal1 524 4322 616 4338 0 _2308_.vdd
rlabel metal2 533 4213 547 4227 0 _2308_.A
rlabel metal2 573 4213 587 4227 0 _2308_.B
rlabel metal2 553 4193 567 4207 0 _2308_.Y
rlabel metal1 784 4082 1036 4098 0 _2393_.gnd
rlabel metal1 784 4322 1036 4338 0 _2393_.vdd
rlabel metal2 933 4173 947 4187 0 _2393_.D
rlabel metal2 893 4173 907 4187 0 _2393_.CLK
rlabel metal2 813 4173 827 4187 0 _2393_.Q
rlabel metal1 724 4082 796 4098 0 _2326_.gnd
rlabel metal1 724 4322 796 4338 0 _2326_.vdd
rlabel metal2 773 4153 787 4167 0 _2326_.A
rlabel metal2 753 4193 767 4207 0 _2326_.Y
rlabel metal1 604 4082 736 4098 0 _2335_.gnd
rlabel metal1 604 4322 736 4338 0 _2335_.vdd
rlabel metal2 713 4173 727 4187 0 _2335_.A
rlabel metal2 693 4193 707 4207 0 _2335_.B
rlabel metal2 633 4173 647 4187 0 _2335_.C
rlabel metal2 653 4193 667 4207 0 _2335_.D
rlabel metal2 673 4173 687 4187 0 _2335_.Y
rlabel metal1 1024 4082 1116 4098 0 _1519_.gnd
rlabel metal1 1024 4322 1116 4338 0 _1519_.vdd
rlabel metal2 1033 4213 1047 4227 0 _1519_.A
rlabel metal2 1073 4213 1087 4227 0 _1519_.B
rlabel metal2 1053 4193 1067 4207 0 _1519_.Y
rlabel metal1 1104 4082 1356 4098 0 _1611_.gnd
rlabel metal1 1104 4322 1356 4338 0 _1611_.vdd
rlabel metal2 1253 4173 1267 4187 0 _1611_.D
rlabel metal2 1213 4173 1227 4187 0 _1611_.CLK
rlabel metal2 1133 4173 1147 4187 0 _1611_.Q
rlabel metal1 1484 4082 1596 4098 0 _2183_.gnd
rlabel metal1 1484 4322 1596 4338 0 _2183_.vdd
rlabel metal2 1573 4173 1587 4187 0 _2183_.A
rlabel metal2 1553 4193 1567 4207 0 _2183_.B
rlabel metal2 1513 4193 1527 4207 0 _2183_.C
rlabel metal2 1533 4173 1547 4187 0 _2183_.Y
rlabel metal1 1424 4082 1496 4098 0 _2177_.gnd
rlabel metal1 1424 4322 1496 4338 0 _2177_.vdd
rlabel metal2 1433 4153 1447 4167 0 _2177_.A
rlabel metal2 1453 4193 1467 4207 0 _2177_.Y
rlabel metal1 1344 4082 1436 4098 0 _2182_.gnd
rlabel metal1 1344 4322 1436 4338 0 _2182_.vdd
rlabel metal2 1353 4213 1367 4227 0 _2182_.A
rlabel metal2 1393 4213 1407 4227 0 _2182_.B
rlabel metal2 1373 4193 1387 4207 0 _2182_.Y
rlabel metal1 1584 4082 1696 4098 0 _1579_.gnd
rlabel metal1 1584 4322 1696 4338 0 _1579_.vdd
rlabel metal2 1673 4193 1687 4207 0 _1579_.A
rlabel metal2 1653 4153 1667 4167 0 _1579_.B
rlabel metal2 1633 4193 1647 4207 0 _1579_.C
rlabel metal2 1613 4173 1627 4187 0 _1579_.Y
rlabel metal1 1844 4082 2096 4098 0 _2383_.gnd
rlabel metal1 1844 4322 2096 4338 0 _2383_.vdd
rlabel metal2 1993 4173 2007 4187 0 _2383_.D
rlabel metal2 1953 4173 1967 4187 0 _2383_.CLK
rlabel metal2 1873 4173 1887 4187 0 _2383_.Q
rlabel metal1 1684 4082 1776 4098 0 _1521_.gnd
rlabel metal1 1684 4322 1776 4338 0 _1521_.vdd
rlabel metal2 1753 4213 1767 4227 0 _1521_.A
rlabel metal2 1713 4213 1727 4227 0 _1521_.B
rlabel metal2 1733 4193 1747 4207 0 _1521_.Y
rlabel metal1 1764 4082 1856 4098 0 _1520_.gnd
rlabel metal1 1764 4322 1856 4338 0 _1520_.vdd
rlabel metal2 1773 4213 1787 4227 0 _1520_.A
rlabel metal2 1813 4213 1827 4227 0 _1520_.B
rlabel metal2 1793 4193 1807 4207 0 _1520_.Y
rlabel metal1 2084 4082 2176 4098 0 _2212_.gnd
rlabel metal1 2084 4322 2176 4338 0 _2212_.vdd
rlabel metal2 2093 4213 2107 4227 0 _2212_.A
rlabel metal2 2133 4213 2147 4227 0 _2212_.B
rlabel metal2 2113 4193 2127 4207 0 _2212_.Y
rlabel metal1 2264 4082 2516 4098 0 _2370_.gnd
rlabel metal1 2264 4322 2516 4338 0 _2370_.vdd
rlabel metal2 2353 4173 2367 4187 0 _2370_.D
rlabel metal2 2393 4173 2407 4187 0 _2370_.CLK
rlabel metal2 2473 4173 2487 4187 0 _2370_.Q
rlabel metal1 2164 4082 2276 4098 0 _2213_.gnd
rlabel metal1 2164 4322 2276 4338 0 _2213_.vdd
rlabel metal2 2253 4173 2267 4187 0 _2213_.A
rlabel metal2 2233 4193 2247 4207 0 _2213_.B
rlabel metal2 2193 4193 2207 4207 0 _2213_.C
rlabel metal2 2213 4173 2227 4187 0 _2213_.Y
rlabel metal1 2644 4082 2756 4098 0 _1796_.gnd
rlabel metal1 2644 4322 2756 4338 0 _1796_.vdd
rlabel metal2 2653 4173 2667 4187 0 _1796_.A
rlabel metal2 2673 4193 2687 4207 0 _1796_.B
rlabel metal2 2713 4193 2727 4207 0 _1796_.C
rlabel metal2 2693 4173 2707 4187 0 _1796_.Y
rlabel metal1 2504 4082 2596 4098 0 _2217_.gnd
rlabel metal1 2504 4322 2596 4338 0 _2217_.vdd
rlabel metal2 2533 4173 2547 4187 0 _2217_.B
rlabel metal2 2573 4173 2587 4187 0 _2217_.A
rlabel metal2 2553 4153 2567 4167 0 _2217_.Y
rlabel metal1 2584 4082 2656 4098 0 _1755_.gnd
rlabel metal1 2584 4322 2656 4338 0 _1755_.vdd
rlabel metal2 2593 4153 2607 4167 0 _1755_.A
rlabel metal2 2613 4193 2627 4207 0 _1755_.Y
rlabel metal1 2824 4082 2936 4098 0 _2210_.gnd
rlabel metal1 2824 4322 2936 4338 0 _2210_.vdd
rlabel metal2 2913 4173 2927 4187 0 _2210_.A
rlabel metal2 2893 4193 2907 4207 0 _2210_.B
rlabel metal2 2853 4193 2867 4207 0 _2210_.C
rlabel metal2 2873 4173 2887 4187 0 _2210_.Y
rlabel metal1 2924 4082 2996 4098 0 _2205_.gnd
rlabel metal1 2924 4322 2996 4338 0 _2205_.vdd
rlabel metal2 2933 4153 2947 4167 0 _2205_.A
rlabel metal2 2953 4193 2967 4207 0 _2205_.Y
rlabel metal1 2744 4082 2836 4098 0 _2211_.gnd
rlabel metal1 2744 4322 2836 4338 0 _2211_.vdd
rlabel metal2 2753 4213 2767 4227 0 _2211_.A
rlabel metal2 2793 4213 2807 4227 0 _2211_.B
rlabel metal2 2773 4193 2787 4207 0 _2211_.Y
rlabel metal1 3124 4082 3376 4098 0 _2369_.gnd
rlabel metal1 3124 4322 3376 4338 0 _2369_.vdd
rlabel metal2 3273 4173 3287 4187 0 _2369_.D
rlabel metal2 3233 4173 3247 4187 0 _2369_.CLK
rlabel metal2 3153 4173 3167 4187 0 _2369_.Q
rlabel metal1 2984 4082 3076 4098 0 _2206_.gnd
rlabel metal1 2984 4322 3076 4338 0 _2206_.vdd
rlabel metal2 3033 4173 3047 4187 0 _2206_.B
rlabel metal2 2993 4173 3007 4187 0 _2206_.A
rlabel metal2 3013 4153 3027 4167 0 _2206_.Y
rlabel metal1 3064 4082 3136 4098 0 _1731_.gnd
rlabel metal1 3064 4322 3136 4338 0 _1731_.vdd
rlabel metal2 3113 4153 3127 4167 0 _1731_.A
rlabel metal2 3093 4193 3107 4207 0 _1731_.Y
rlabel metal1 3364 4082 3496 4098 0 _1754_.gnd
rlabel metal1 3364 4322 3496 4338 0 _1754_.vdd
rlabel metal2 3373 4173 3387 4187 0 _1754_.A
rlabel metal2 3393 4193 3407 4207 0 _1754_.B
rlabel metal2 3453 4173 3467 4187 0 _1754_.C
rlabel metal2 3413 4173 3427 4187 0 _1754_.Y
rlabel metal2 3433 4193 3447 4207 0 _1754_.D
rlabel metal1 3564 4082 3776 4098 0 CLKBUF1_insert28.gnd
rlabel metal1 3564 4322 3776 4338 0 CLKBUF1_insert28.vdd
rlabel metal2 3593 4193 3607 4207 0 CLKBUF1_insert28.A
rlabel metal2 3733 4193 3747 4207 0 CLKBUF1_insert28.Y
rlabel metal1 3484 4082 3576 4098 0 _1678_.gnd
rlabel metal1 3484 4322 3576 4338 0 _1678_.vdd
rlabel metal2 3493 4213 3507 4227 0 _1678_.A
rlabel metal2 3533 4213 3547 4227 0 _1678_.B
rlabel metal2 3513 4193 3527 4207 0 _1678_.Y
rlabel metal1 4004 4082 4076 4098 0 _1792_.gnd
rlabel metal1 4004 4322 4076 4338 0 _1792_.vdd
rlabel metal2 4013 4153 4027 4167 0 _1792_.A
rlabel metal2 4033 4193 4047 4207 0 _1792_.Y
rlabel metal1 3844 4082 3936 4098 0 _1753_.gnd
rlabel metal1 3844 4322 3936 4338 0 _1753_.vdd
rlabel metal2 3853 4213 3867 4227 0 _1753_.A
rlabel metal2 3893 4213 3907 4227 0 _1753_.B
rlabel metal2 3873 4193 3887 4207 0 _1753_.Y
rlabel metal1 3924 4082 4016 4098 0 _1672_.gnd
rlabel metal1 3924 4322 4016 4338 0 _1672_.vdd
rlabel metal2 3993 4213 4007 4227 0 _1672_.A
rlabel metal2 3953 4213 3967 4227 0 _1672_.B
rlabel metal2 3973 4193 3987 4207 0 _1672_.Y
rlabel metal1 3764 4082 3856 4098 0 _1666_.gnd
rlabel metal1 3764 4322 3856 4338 0 _1666_.vdd
rlabel metal2 3773 4213 3787 4227 0 _1666_.A
rlabel metal2 3813 4213 3827 4227 0 _1666_.B
rlabel metal2 3793 4193 3807 4207 0 _1666_.Y
rlabel metal1 4264 4082 4516 4098 0 _2354_.gnd
rlabel metal1 4264 4322 4516 4338 0 _2354_.vdd
rlabel metal2 4353 4173 4367 4187 0 _2354_.D
rlabel metal2 4393 4173 4407 4187 0 _2354_.CLK
rlabel metal2 4473 4173 4487 4187 0 _2354_.Q
rlabel metal1 4164 4082 4276 4098 0 _1799_.gnd
rlabel metal1 4164 4322 4276 4338 0 _1799_.vdd
rlabel metal2 4173 4173 4187 4187 0 _1799_.A
rlabel metal2 4193 4193 4207 4207 0 _1799_.B
rlabel metal2 4233 4193 4247 4207 0 _1799_.C
rlabel metal2 4213 4173 4227 4187 0 _1799_.Y
rlabel metal1 4064 4082 4176 4098 0 _1673_.gnd
rlabel metal1 4064 4322 4176 4338 0 _1673_.vdd
rlabel metal2 4153 4173 4167 4187 0 _1673_.A
rlabel metal2 4133 4193 4147 4207 0 _1673_.B
rlabel metal2 4093 4193 4107 4207 0 _1673_.C
rlabel metal2 4113 4173 4127 4187 0 _1673_.Y
rlabel metal1 4504 4082 4616 4098 0 _1697_.gnd
rlabel metal1 4504 4322 4616 4338 0 _1697_.vdd
rlabel metal2 4593 4173 4607 4187 0 _1697_.A
rlabel metal2 4573 4193 4587 4207 0 _1697_.B
rlabel metal2 4533 4193 4547 4207 0 _1697_.C
rlabel metal2 4553 4173 4567 4187 0 _1697_.Y
rlabel metal1 4604 4082 4856 4098 0 _2362_.gnd
rlabel metal1 4604 4322 4856 4338 0 _2362_.vdd
rlabel metal2 4693 4173 4707 4187 0 _2362_.D
rlabel metal2 4733 4173 4747 4187 0 _2362_.CLK
rlabel metal2 4813 4173 4827 4187 0 _2362_.Q
rlabel metal1 4904 4082 5016 4098 0 _1751_.gnd
rlabel metal1 4904 4322 5016 4338 0 _1751_.vdd
rlabel metal2 4993 4193 5007 4207 0 _1751_.A
rlabel metal2 4973 4153 4987 4167 0 _1751_.B
rlabel metal2 4953 4193 4967 4207 0 _1751_.C
rlabel metal2 4933 4173 4947 4187 0 _1751_.Y
rlabel metal1 5004 4082 5116 4098 0 _1752_.gnd
rlabel metal1 5004 4322 5116 4338 0 _1752_.vdd
rlabel metal2 5013 4193 5027 4207 0 _1752_.A
rlabel metal2 5033 4213 5047 4227 0 _1752_.B
rlabel metal2 5053 4193 5067 4207 0 _1752_.C
rlabel metal2 5073 4213 5087 4227 0 _1752_.Y
rlabel metal1 4844 4082 4916 4098 0 _1671_.gnd
rlabel metal1 4844 4322 4916 4338 0 _1671_.vdd
rlabel metal2 4893 4193 4907 4207 0 _1671_.A
rlabel metal2 4873 4173 4887 4187 0 _1671_.Y
rlabel metal1 5264 4082 5516 4098 0 _2361_.gnd
rlabel metal1 5264 4322 5516 4338 0 _2361_.vdd
rlabel metal2 5353 4173 5367 4187 0 _2361_.D
rlabel metal2 5393 4173 5407 4187 0 _2361_.CLK
rlabel metal2 5473 4173 5487 4187 0 _2361_.Q
rlabel metal1 5164 4082 5276 4098 0 _1694_.gnd
rlabel metal1 5164 4322 5276 4338 0 _1694_.vdd
rlabel metal2 5173 4173 5187 4187 0 _1694_.A
rlabel metal2 5193 4193 5207 4207 0 _1694_.B
rlabel metal2 5233 4193 5247 4207 0 _1694_.C
rlabel metal2 5213 4173 5227 4187 0 _1694_.Y
rlabel metal1 5104 4082 5176 4098 0 _1692_.gnd
rlabel metal1 5104 4322 5176 4338 0 _1692_.vdd
rlabel metal2 5153 4153 5167 4167 0 _1692_.A
rlabel metal2 5133 4193 5147 4207 0 _1692_.Y
rlabel metal1 5584 4082 5656 4098 0 _1683_.gnd
rlabel metal1 5584 4322 5656 4338 0 _1683_.vdd
rlabel metal2 5593 4153 5607 4167 0 _1683_.A
rlabel metal2 5613 4193 5627 4207 0 _1683_.Y
rlabel metal1 5504 4082 5596 4098 0 _1733_.gnd
rlabel metal1 5504 4322 5596 4338 0 _1733_.vdd
rlabel metal2 5513 4213 5527 4227 0 _1733_.A
rlabel metal2 5553 4213 5567 4227 0 _1733_.B
rlabel metal2 5533 4193 5547 4207 0 _1733_.Y
rlabel metal1 5644 4082 5756 4098 0 _1740_.gnd
rlabel metal1 5644 4322 5756 4338 0 _1740_.vdd
rlabel metal2 5653 4173 5667 4187 0 _1740_.A
rlabel metal2 5673 4193 5687 4207 0 _1740_.B
rlabel metal2 5713 4193 5727 4207 0 _1740_.C
rlabel metal2 5693 4173 5707 4187 0 _1740_.Y
rlabel metal1 5844 4082 5956 4098 0 _1742_.gnd
rlabel metal1 5844 4322 5956 4338 0 _1742_.vdd
rlabel metal2 5853 4193 5867 4207 0 _1742_.A
rlabel metal2 5873 4213 5887 4227 0 _1742_.B
rlabel metal2 5893 4193 5907 4207 0 _1742_.C
rlabel metal2 5913 4213 5927 4227 0 _1742_.Y
rlabel metal1 5744 4082 5856 4098 0 _1736_.gnd
rlabel metal1 5744 4322 5856 4338 0 _1736_.vdd
rlabel metal2 5833 4173 5847 4187 0 _1736_.A
rlabel metal2 5773 4173 5787 4187 0 _1736_.Y
rlabel metal2 5793 4213 5807 4227 0 _1736_.B
rlabel metal1 6104 4082 6196 4098 0 BUFX2_insert13.gnd
rlabel metal1 6104 4322 6196 4338 0 BUFX2_insert13.vdd
rlabel metal2 6113 4173 6127 4187 0 BUFX2_insert13.A
rlabel metal2 6153 4173 6167 4187 0 BUFX2_insert13.Y
rlabel metal1 6004 4082 6116 4098 0 _1741_.gnd
rlabel metal1 6004 4322 6116 4338 0 _1741_.vdd
rlabel metal2 6013 4173 6027 4187 0 _1741_.A
rlabel metal2 6033 4193 6047 4207 0 _1741_.B
rlabel metal2 6073 4193 6087 4207 0 _1741_.C
rlabel metal2 6053 4173 6067 4187 0 _1741_.Y
rlabel metal1 5944 4082 6016 4098 0 _1689_.gnd
rlabel metal1 5944 4322 6016 4338 0 _1689_.vdd
rlabel metal2 5993 4193 6007 4207 0 _1689_.A
rlabel metal2 5973 4173 5987 4187 0 _1689_.Y
rlabel metal1 6184 4082 6276 4098 0 _1737_.gnd
rlabel metal1 6184 4322 6276 4338 0 _1737_.vdd
rlabel metal2 6193 4213 6207 4227 0 _1737_.A
rlabel metal2 6233 4213 6247 4227 0 _1737_.B
rlabel metal2 6213 4193 6227 4207 0 _1737_.Y
rlabel metal1 6364 4082 6456 4098 0 _1720_.gnd
rlabel metal1 6364 4322 6456 4338 0 _1720_.vdd
rlabel metal2 6373 4213 6387 4227 0 _1720_.A
rlabel metal2 6413 4213 6427 4227 0 _1720_.B
rlabel metal2 6393 4193 6407 4207 0 _1720_.Y
rlabel metal1 6264 4082 6376 4098 0 _1735_.gnd
rlabel metal1 6264 4322 6376 4338 0 _1735_.vdd
rlabel metal2 6353 4173 6367 4187 0 _1735_.A
rlabel metal2 6293 4173 6307 4187 0 _1735_.Y
rlabel metal2 6313 4213 6327 4227 0 _1735_.B
rlabel metal1 6444 4082 6516 4098 0 _1756_.gnd
rlabel metal1 6444 4322 6516 4338 0 _1756_.vdd
rlabel metal2 6453 4153 6467 4167 0 _1756_.A
rlabel metal2 6473 4193 6487 4207 0 _1756_.Y
rlabel metal1 6504 4082 6616 4098 0 _1788_.gnd
rlabel metal1 6504 4322 6616 4338 0 _1788_.vdd
rlabel metal2 6593 4193 6607 4207 0 _1788_.A
rlabel metal2 6573 4153 6587 4167 0 _1788_.B
rlabel metal2 6553 4193 6567 4207 0 _1788_.C
rlabel metal2 6533 4173 6547 4187 0 _1788_.Y
rlabel metal1 6604 4082 6716 4098 0 _1789_.gnd
rlabel metal1 6604 4322 6716 4338 0 _1789_.vdd
rlabel metal2 6613 4193 6627 4207 0 _1789_.A
rlabel metal2 6633 4213 6647 4227 0 _1789_.B
rlabel metal2 6653 4193 6667 4207 0 _1789_.C
rlabel metal2 6673 4213 6687 4227 0 _1789_.Y
rlabel nsubstratencontact 6716 4328 6716 4328 0 FILL100650x61350.vdd
rlabel metal1 6704 4082 6736 4098 0 FILL100650x61350.gnd
rlabel metal1 204 4562 316 4578 0 _2340_.gnd
rlabel metal1 204 4322 316 4338 0 _2340_.vdd
rlabel metal2 213 4473 227 4487 0 _2340_.A
rlabel metal2 233 4453 247 4467 0 _2340_.B
rlabel metal2 273 4453 287 4467 0 _2340_.C
rlabel metal2 253 4473 267 4487 0 _2340_.Y
rlabel metal1 64 4562 156 4578 0 _2338_.gnd
rlabel metal1 64 4322 156 4338 0 _2338_.vdd
rlabel metal2 93 4473 107 4487 0 _2338_.B
rlabel metal2 133 4473 147 4487 0 _2338_.A
rlabel metal2 113 4493 127 4507 0 _2338_.Y
rlabel metal1 4 4562 76 4578 0 _2339_.gnd
rlabel metal1 4 4322 76 4338 0 _2339_.vdd
rlabel metal2 53 4493 67 4507 0 _2339_.A
rlabel metal2 33 4453 47 4467 0 _2339_.Y
rlabel metal1 144 4562 216 4578 0 _2323_.gnd
rlabel metal1 144 4322 216 4338 0 _2323_.vdd
rlabel metal2 193 4493 207 4507 0 _2323_.A
rlabel metal2 173 4453 187 4467 0 _2323_.Y
rlabel metal1 384 4562 496 4578 0 _2328_.gnd
rlabel metal1 384 4322 496 4338 0 _2328_.vdd
rlabel metal2 393 4473 407 4487 0 _2328_.A
rlabel metal2 413 4453 427 4467 0 _2328_.B
rlabel metal2 453 4453 467 4467 0 _2328_.C
rlabel metal2 433 4473 447 4487 0 _2328_.Y
rlabel metal1 304 4562 396 4578 0 _2321_.gnd
rlabel metal1 304 4322 396 4338 0 _2321_.vdd
rlabel metal2 333 4473 347 4487 0 _2321_.B
rlabel metal2 373 4473 387 4487 0 _2321_.A
rlabel metal2 353 4493 367 4507 0 _2321_.Y
rlabel metal1 484 4562 596 4578 0 _2333_.gnd
rlabel metal1 484 4322 596 4338 0 _2333_.vdd
rlabel metal2 493 4493 507 4507 0 _2333_.A
rlabel metal2 513 4473 527 4487 0 _2333_.B
rlabel metal2 553 4453 567 4467 0 _2333_.Y
rlabel metal1 744 4562 836 4578 0 _2320_.gnd
rlabel metal1 744 4322 836 4338 0 _2320_.vdd
rlabel metal2 793 4473 807 4487 0 _2320_.B
rlabel metal2 753 4473 767 4487 0 _2320_.A
rlabel metal2 773 4493 787 4507 0 _2320_.Y
rlabel metal1 684 4562 756 4578 0 _2327_.gnd
rlabel metal1 684 4322 756 4338 0 _2327_.vdd
rlabel metal2 733 4493 747 4507 0 _2327_.A
rlabel metal2 713 4453 727 4467 0 _2327_.Y
rlabel metal1 584 4562 696 4578 0 _2334_.gnd
rlabel metal1 584 4322 696 4338 0 _2334_.vdd
rlabel metal2 593 4453 607 4467 0 _2334_.A
rlabel metal2 613 4493 627 4507 0 _2334_.B
rlabel metal2 633 4453 647 4467 0 _2334_.C
rlabel metal2 653 4473 667 4487 0 _2334_.Y
rlabel metal1 1024 4562 1236 4578 0 CLKBUF1_insert33.gnd
rlabel metal1 1024 4322 1236 4338 0 CLKBUF1_insert33.vdd
rlabel metal2 1053 4453 1067 4467 0 CLKBUF1_insert33.A
rlabel metal2 1193 4453 1207 4467 0 CLKBUF1_insert33.Y
rlabel metal1 884 4562 976 4578 0 _2319_.gnd
rlabel metal1 884 4322 976 4338 0 _2319_.vdd
rlabel metal2 933 4473 947 4487 0 _2319_.B
rlabel metal2 893 4473 907 4487 0 _2319_.A
rlabel metal2 913 4493 927 4507 0 _2319_.Y
rlabel metal1 964 4562 1036 4578 0 _2318_.gnd
rlabel metal1 964 4322 1036 4338 0 _2318_.vdd
rlabel metal2 973 4493 987 4507 0 _2318_.A
rlabel metal2 993 4453 1007 4467 0 _2318_.Y
rlabel metal1 824 4562 896 4578 0 _2317_.gnd
rlabel metal1 824 4322 896 4338 0 _2317_.vdd
rlabel metal2 833 4493 847 4507 0 _2317_.A
rlabel metal2 853 4453 867 4467 0 _2317_.Y
rlabel metal1 1224 4562 1316 4578 0 BUFX2_insert2.gnd
rlabel metal1 1224 4322 1316 4338 0 BUFX2_insert2.vdd
rlabel metal2 1233 4473 1247 4487 0 BUFX2_insert2.A
rlabel metal2 1273 4473 1287 4487 0 BUFX2_insert2.Y
rlabel metal1 1304 4562 1376 4578 0 _2179_.gnd
rlabel metal1 1304 4322 1376 4338 0 _2179_.vdd
rlabel metal2 1353 4493 1367 4507 0 _2179_.A
rlabel metal2 1333 4453 1347 4467 0 _2179_.Y
rlabel metal1 1364 4562 1456 4578 0 _2178_.gnd
rlabel metal1 1364 4322 1456 4338 0 _2178_.vdd
rlabel metal2 1393 4473 1407 4487 0 _2178_.B
rlabel metal2 1433 4473 1447 4487 0 _2178_.A
rlabel metal2 1413 4493 1427 4507 0 _2178_.Y
rlabel metal1 1444 4562 1536 4578 0 _2181_.gnd
rlabel metal1 1444 4322 1536 4338 0 _2181_.vdd
rlabel metal2 1513 4433 1527 4447 0 _2181_.A
rlabel metal2 1473 4433 1487 4447 0 _2181_.B
rlabel metal2 1493 4453 1507 4467 0 _2181_.Y
rlabel metal1 1524 4562 1616 4578 0 _2180_.gnd
rlabel metal1 1524 4322 1616 4338 0 _2180_.vdd
rlabel metal2 1533 4433 1547 4447 0 _2180_.A
rlabel metal2 1573 4433 1587 4447 0 _2180_.B
rlabel metal2 1553 4453 1567 4467 0 _2180_.Y
rlabel metal1 1604 4562 1736 4578 0 _1797_.gnd
rlabel metal1 1604 4322 1736 4338 0 _1797_.vdd
rlabel metal2 1693 4473 1707 4487 0 _1797_.A
rlabel metal2 1653 4473 1667 4487 0 _1797_.Y
rlabel metal1 1724 4562 1976 4578 0 _2371_.gnd
rlabel metal1 1724 4322 1976 4338 0 _2371_.vdd
rlabel metal2 1813 4473 1827 4487 0 _2371_.D
rlabel metal2 1853 4473 1867 4487 0 _2371_.CLK
rlabel metal2 1933 4473 1947 4487 0 _2371_.Q
rlabel metal1 2044 4562 2296 4578 0 _2372_.gnd
rlabel metal1 2044 4322 2296 4338 0 _2372_.vdd
rlabel metal2 2193 4473 2207 4487 0 _2372_.D
rlabel metal2 2153 4473 2167 4487 0 _2372_.CLK
rlabel metal2 2073 4473 2087 4487 0 _2372_.Q
rlabel metal1 1964 4562 2056 4578 0 _1852_.gnd
rlabel metal1 1964 4322 2056 4338 0 _1852_.vdd
rlabel metal2 1973 4433 1987 4447 0 _1852_.A
rlabel metal2 2013 4433 2027 4447 0 _1852_.B
rlabel metal2 1993 4453 2007 4467 0 _1852_.Y
rlabel metal1 2344 4562 2436 4578 0 _2196_.gnd
rlabel metal1 2344 4322 2436 4338 0 _2196_.vdd
rlabel metal2 2393 4473 2407 4487 0 _2196_.B
rlabel metal2 2353 4473 2367 4487 0 _2196_.A
rlabel metal2 2373 4493 2387 4507 0 _2196_.Y
rlabel metal1 2284 4562 2356 4578 0 _2194_.gnd
rlabel metal1 2284 4322 2356 4338 0 _2194_.vdd
rlabel metal2 2293 4493 2307 4507 0 _2194_.A
rlabel metal2 2313 4453 2327 4467 0 _2194_.Y
rlabel metal1 2564 4562 2816 4578 0 _2368_.gnd
rlabel metal1 2564 4322 2816 4338 0 _2368_.vdd
rlabel metal2 2713 4473 2727 4487 0 _2368_.D
rlabel metal2 2673 4473 2687 4487 0 _2368_.CLK
rlabel metal2 2593 4473 2607 4487 0 _2368_.Q
rlabel metal1 2424 4562 2516 4578 0 _2195_.gnd
rlabel metal1 2424 4322 2516 4338 0 _2195_.vdd
rlabel metal2 2473 4473 2487 4487 0 _2195_.B
rlabel metal2 2433 4473 2447 4487 0 _2195_.A
rlabel metal2 2453 4493 2467 4507 0 _2195_.Y
rlabel metal1 2504 4562 2576 4578 0 _1718_.gnd
rlabel metal1 2504 4322 2576 4338 0 _1718_.vdd
rlabel metal2 2513 4493 2527 4507 0 _1718_.A
rlabel metal2 2533 4453 2547 4467 0 _1718_.Y
rlabel metal1 2804 4562 2916 4578 0 _1730_.gnd
rlabel metal1 2804 4322 2916 4338 0 _1730_.vdd
rlabel metal2 2813 4473 2827 4487 0 _1730_.A
rlabel metal2 2833 4453 2847 4467 0 _1730_.B
rlabel metal2 2873 4453 2887 4467 0 _1730_.C
rlabel metal2 2853 4473 2867 4487 0 _1730_.Y
rlabel metal1 2904 4562 2996 4578 0 _1729_.gnd
rlabel metal1 2904 4322 2996 4338 0 _1729_.vdd
rlabel metal2 2913 4433 2927 4447 0 _1729_.A
rlabel metal2 2953 4433 2967 4447 0 _1729_.B
rlabel metal2 2933 4453 2947 4467 0 _1729_.Y
rlabel metal1 3144 4562 3396 4578 0 _2364_.gnd
rlabel metal1 3144 4322 3396 4338 0 _2364_.vdd
rlabel metal2 3293 4473 3307 4487 0 _2364_.D
rlabel metal2 3253 4473 3267 4487 0 _2364_.CLK
rlabel metal2 3173 4473 3187 4487 0 _2364_.Q
rlabel metal1 3044 4562 3156 4578 0 _1709_.gnd
rlabel metal1 3044 4322 3156 4338 0 _1709_.vdd
rlabel metal2 3053 4473 3067 4487 0 _1709_.A
rlabel metal2 3073 4453 3087 4467 0 _1709_.B
rlabel metal2 3113 4453 3127 4467 0 _1709_.C
rlabel metal2 3093 4473 3107 4487 0 _1709_.Y
rlabel metal1 2984 4562 3056 4578 0 _1707_.gnd
rlabel metal1 2984 4322 3056 4338 0 _1707_.vdd
rlabel metal2 3033 4493 3047 4507 0 _1707_.A
rlabel metal2 3013 4453 3027 4467 0 _1707_.Y
rlabel metal1 3384 4562 3496 4578 0 _1703_.gnd
rlabel metal1 3384 4322 3496 4338 0 _1703_.vdd
rlabel metal2 3393 4473 3407 4487 0 _1703_.A
rlabel metal2 3413 4453 3427 4467 0 _1703_.B
rlabel metal2 3453 4453 3467 4467 0 _1703_.C
rlabel metal2 3433 4473 3447 4487 0 _1703_.Y
rlabel metal1 3584 4562 3836 4578 0 _2355_.gnd
rlabel metal1 3584 4322 3836 4338 0 _2355_.vdd
rlabel metal2 3673 4473 3687 4487 0 _2355_.D
rlabel metal2 3713 4473 3727 4487 0 _2355_.CLK
rlabel metal2 3793 4473 3807 4487 0 _2355_.Q
rlabel metal1 3484 4562 3596 4578 0 _1676_.gnd
rlabel metal1 3484 4322 3596 4338 0 _1676_.vdd
rlabel metal2 3573 4473 3587 4487 0 _1676_.A
rlabel metal2 3553 4453 3567 4467 0 _1676_.B
rlabel metal2 3513 4453 3527 4467 0 _1676_.C
rlabel metal2 3533 4473 3547 4487 0 _1676_.Y
rlabel metal1 3924 4562 4176 4578 0 _2352_.gnd
rlabel metal1 3924 4322 4176 4338 0 _2352_.vdd
rlabel metal2 4013 4473 4027 4487 0 _2352_.D
rlabel metal2 4053 4473 4067 4487 0 _2352_.CLK
rlabel metal2 4133 4473 4147 4487 0 _2352_.Q
rlabel metal1 3824 4562 3936 4578 0 _1667_.gnd
rlabel metal1 3824 4322 3936 4338 0 _1667_.vdd
rlabel metal2 3833 4473 3847 4487 0 _1667_.A
rlabel metal2 3853 4453 3867 4467 0 _1667_.B
rlabel metal2 3893 4453 3907 4467 0 _1667_.C
rlabel metal2 3873 4473 3887 4487 0 _1667_.Y
rlabel metal1 4264 4562 4376 4578 0 _1706_.gnd
rlabel metal1 4264 4322 4376 4338 0 _1706_.vdd
rlabel metal2 4273 4473 4287 4487 0 _1706_.A
rlabel metal2 4293 4453 4307 4467 0 _1706_.B
rlabel metal2 4333 4453 4347 4467 0 _1706_.C
rlabel metal2 4313 4473 4327 4487 0 _1706_.Y
rlabel metal1 4164 4562 4276 4578 0 _1708_.gnd
rlabel metal1 4164 4322 4276 4338 0 _1708_.vdd
rlabel metal2 4253 4453 4267 4467 0 _1708_.A
rlabel metal2 4233 4433 4247 4447 0 _1708_.B
rlabel metal2 4213 4453 4227 4467 0 _1708_.C
rlabel metal2 4193 4433 4207 4447 0 _1708_.Y
rlabel metal1 4364 4562 4456 4578 0 _1728_.gnd
rlabel metal1 4364 4322 4456 4338 0 _1728_.vdd
rlabel metal2 4393 4473 4407 4487 0 _1728_.B
rlabel metal2 4433 4473 4447 4487 0 _1728_.A
rlabel metal2 4413 4493 4427 4507 0 _1728_.Y
rlabel metal1 4444 4562 4556 4578 0 _1727_.gnd
rlabel metal1 4444 4322 4556 4338 0 _1727_.vdd
rlabel metal2 4533 4453 4547 4467 0 _1727_.A
rlabel metal2 4513 4493 4527 4507 0 _1727_.B
rlabel metal2 4493 4453 4507 4467 0 _1727_.C
rlabel metal2 4473 4473 4487 4487 0 _1727_.Y
rlabel metal1 4704 4562 4816 4578 0 _1724_.gnd
rlabel metal1 4704 4322 4816 4338 0 _1724_.vdd
rlabel metal2 4713 4473 4727 4487 0 _1724_.A
rlabel metal2 4733 4453 4747 4467 0 _1724_.B
rlabel metal2 4773 4453 4787 4467 0 _1724_.C
rlabel metal2 4753 4473 4767 4487 0 _1724_.Y
rlabel metal1 4644 4562 4716 4578 0 _1726_.gnd
rlabel metal1 4644 4322 4716 4338 0 _1726_.vdd
rlabel metal2 4693 4493 4707 4507 0 _1726_.A
rlabel metal2 4673 4453 4687 4467 0 _1726_.Y
rlabel metal1 4544 4562 4656 4578 0 _1725_.gnd
rlabel metal1 4544 4322 4656 4338 0 _1725_.vdd
rlabel metal2 4553 4453 4567 4467 0 _1725_.A
rlabel metal2 4573 4433 4587 4447 0 _1725_.B
rlabel metal2 4593 4453 4607 4467 0 _1725_.C
rlabel metal2 4613 4433 4627 4447 0 _1725_.Y
rlabel metal1 4804 4562 4916 4578 0 _1723_.gnd
rlabel metal1 4804 4322 4916 4338 0 _1723_.vdd
rlabel metal2 4893 4493 4907 4507 0 _1723_.A
rlabel metal2 4873 4473 4887 4487 0 _1723_.B
rlabel metal2 4833 4453 4847 4467 0 _1723_.Y
rlabel metal1 4904 4562 4996 4578 0 _1722_.gnd
rlabel metal1 4904 4322 4996 4338 0 _1722_.vdd
rlabel metal2 4973 4433 4987 4447 0 _1722_.A
rlabel metal2 4933 4433 4947 4447 0 _1722_.B
rlabel metal2 4953 4453 4967 4467 0 _1722_.Y
rlabel metal1 4984 4562 5096 4578 0 _1748_.gnd
rlabel metal1 4984 4322 5096 4338 0 _1748_.vdd
rlabel metal2 5073 4453 5087 4467 0 _1748_.A
rlabel metal2 5053 4433 5067 4447 0 _1748_.B
rlabel metal2 5033 4453 5047 4467 0 _1748_.C
rlabel metal2 5013 4433 5027 4447 0 _1748_.Y
rlabel metal1 5084 4562 5196 4578 0 _1749_.gnd
rlabel metal1 5084 4322 5196 4338 0 _1749_.vdd
rlabel metal2 5093 4473 5107 4487 0 _1749_.A
rlabel metal2 5113 4453 5127 4467 0 _1749_.B
rlabel metal2 5153 4453 5167 4467 0 _1749_.C
rlabel metal2 5133 4473 5147 4487 0 _1749_.Y
rlabel metal1 5284 4562 5396 4578 0 _1721_.gnd
rlabel metal1 5284 4322 5396 4338 0 _1721_.vdd
rlabel metal2 5293 4473 5307 4487 0 _1721_.A
rlabel metal2 5313 4453 5327 4467 0 _1721_.B
rlabel metal2 5353 4453 5367 4467 0 _1721_.C
rlabel metal2 5333 4473 5347 4487 0 _1721_.Y
rlabel metal1 5184 4562 5296 4578 0 _1732_.gnd
rlabel metal1 5184 4322 5296 4338 0 _1732_.vdd
rlabel metal2 5273 4493 5287 4507 0 _1732_.A
rlabel metal2 5253 4473 5267 4487 0 _1732_.B
rlabel metal2 5213 4453 5227 4467 0 _1732_.Y
rlabel metal1 5384 4562 5456 4578 0 _1695_.gnd
rlabel metal1 5384 4322 5456 4338 0 _1695_.vdd
rlabel metal2 5393 4493 5407 4507 0 _1695_.A
rlabel metal2 5413 4453 5427 4467 0 _1695_.Y
rlabel metal1 5544 4562 5636 4578 0 _1747_.gnd
rlabel metal1 5544 4322 5636 4338 0 _1747_.vdd
rlabel metal2 5553 4433 5567 4447 0 _1747_.A
rlabel metal2 5593 4433 5607 4447 0 _1747_.B
rlabel metal2 5573 4453 5587 4467 0 _1747_.Y
rlabel metal1 5444 4562 5556 4578 0 _1750_.gnd
rlabel metal1 5444 4322 5556 4338 0 _1750_.vdd
rlabel metal2 5533 4453 5547 4467 0 _1750_.A
rlabel metal2 5513 4433 5527 4447 0 _1750_.B
rlabel metal2 5493 4453 5507 4467 0 _1750_.C
rlabel metal2 5473 4433 5487 4447 0 _1750_.Y
rlabel metal1 5624 4562 5736 4578 0 _1744_.gnd
rlabel metal1 5624 4322 5736 4338 0 _1744_.vdd
rlabel metal2 5633 4473 5647 4487 0 _1744_.A
rlabel metal2 5653 4453 5667 4467 0 _1744_.B
rlabel metal2 5693 4453 5707 4467 0 _1744_.C
rlabel metal2 5673 4473 5687 4487 0 _1744_.Y
rlabel metal1 5724 4562 5816 4578 0 _1743_.gnd
rlabel metal1 5724 4322 5816 4338 0 _1743_.vdd
rlabel metal2 5793 4433 5807 4447 0 _1743_.A
rlabel metal2 5753 4433 5767 4447 0 _1743_.B
rlabel metal2 5773 4453 5787 4467 0 _1743_.Y
rlabel metal1 5804 4562 5916 4578 0 _1746_.gnd
rlabel metal1 5804 4322 5916 4338 0 _1746_.vdd
rlabel metal2 5893 4453 5907 4467 0 _1746_.A
rlabel metal2 5873 4433 5887 4447 0 _1746_.B
rlabel metal2 5853 4453 5867 4467 0 _1746_.C
rlabel metal2 5833 4433 5847 4447 0 _1746_.Y
rlabel metal1 5904 4562 6016 4578 0 _1758_.gnd
rlabel metal1 5904 4322 6016 4338 0 _1758_.vdd
rlabel metal2 5993 4473 6007 4487 0 _1758_.A
rlabel metal2 5973 4453 5987 4467 0 _1758_.B
rlabel metal2 5933 4453 5947 4467 0 _1758_.C
rlabel metal2 5953 4473 5967 4487 0 _1758_.Y
rlabel metal1 6064 4562 6136 4578 0 _1784_.gnd
rlabel metal1 6064 4322 6136 4338 0 _1784_.vdd
rlabel metal2 6113 4493 6127 4507 0 _1784_.A
rlabel metal2 6093 4453 6107 4467 0 _1784_.Y
rlabel metal1 6004 4562 6076 4578 0 _1757_.gnd
rlabel metal1 6004 4322 6076 4338 0 _1757_.vdd
rlabel metal2 6013 4493 6027 4507 0 _1757_.A
rlabel metal2 6033 4453 6047 4467 0 _1757_.Y
rlabel metal1 6124 4562 6236 4578 0 _1783_.gnd
rlabel metal1 6124 4322 6236 4338 0 _1783_.vdd
rlabel metal2 6133 4453 6147 4467 0 _1783_.A
rlabel metal2 6153 4433 6167 4447 0 _1783_.B
rlabel metal2 6173 4453 6187 4467 0 _1783_.C
rlabel metal2 6193 4433 6207 4447 0 _1783_.Y
rlabel metal1 6224 4562 6336 4578 0 _1782_.gnd
rlabel metal1 6224 4322 6336 4338 0 _1782_.vdd
rlabel metal2 6313 4473 6327 4487 0 _1782_.A
rlabel metal2 6293 4453 6307 4467 0 _1782_.B
rlabel metal2 6253 4453 6267 4467 0 _1782_.C
rlabel metal2 6273 4473 6287 4487 0 _1782_.Y
rlabel metal1 6324 4562 6436 4578 0 _1786_.gnd
rlabel metal1 6324 4322 6436 4338 0 _1786_.vdd
rlabel metal2 6333 4453 6347 4467 0 _1786_.A
rlabel metal2 6353 4433 6367 4447 0 _1786_.B
rlabel metal2 6373 4453 6387 4467 0 _1786_.C
rlabel metal2 6393 4433 6407 4447 0 _1786_.Y
rlabel metal1 6524 4562 6636 4578 0 _1785_.gnd
rlabel metal1 6524 4322 6636 4338 0 _1785_.vdd
rlabel metal2 6533 4473 6547 4487 0 _1785_.A
rlabel metal2 6553 4453 6567 4467 0 _1785_.B
rlabel metal2 6593 4453 6607 4467 0 _1785_.C
rlabel metal2 6573 4473 6587 4487 0 _1785_.Y
rlabel metal1 6624 4562 6696 4578 0 _1759_.gnd
rlabel metal1 6624 4322 6696 4338 0 _1759_.vdd
rlabel metal2 6633 4493 6647 4507 0 _1759_.A
rlabel metal2 6653 4453 6667 4467 0 _1759_.Y
rlabel metal1 6424 4562 6536 4578 0 _1787_.gnd
rlabel metal1 6424 4322 6536 4338 0 _1787_.vdd
rlabel metal2 6433 4453 6447 4467 0 _1787_.A
rlabel metal2 6453 4433 6467 4447 0 _1787_.B
rlabel metal2 6473 4453 6487 4467 0 _1787_.C
rlabel metal2 6493 4433 6507 4447 0 _1787_.Y
rlabel nsubstratencontact 6724 4332 6724 4332 0 FILL100650x64950.vdd
rlabel metal1 6704 4562 6736 4578 0 FILL100650x64950.gnd
rlabel nsubstratencontact 6704 4332 6704 4332 0 FILL100350x64950.vdd
rlabel metal1 6684 4562 6716 4578 0 FILL100350x64950.gnd
rlabel metal1 4 4562 216 4578 0 CLKBUF1_insert36.gnd
rlabel metal1 4 4802 216 4818 0 CLKBUF1_insert36.vdd
rlabel metal2 33 4673 47 4687 0 CLKBUF1_insert36.A
rlabel metal2 173 4673 187 4687 0 CLKBUF1_insert36.Y
rlabel metal1 204 4562 296 4578 0 _2322_.gnd
rlabel metal1 204 4802 296 4818 0 _2322_.vdd
rlabel metal2 233 4653 247 4667 0 _2322_.B
rlabel metal2 273 4653 287 4667 0 _2322_.A
rlabel metal2 253 4633 267 4647 0 _2322_.Y
rlabel metal1 504 4562 596 4578 0 _2331_.gnd
rlabel metal1 504 4802 596 4818 0 _2331_.vdd
rlabel metal2 533 4653 547 4667 0 _2331_.B
rlabel metal2 573 4653 587 4667 0 _2331_.A
rlabel metal2 553 4633 567 4647 0 _2331_.Y
rlabel metal1 444 4562 516 4578 0 _2332_.gnd
rlabel metal1 444 4802 516 4818 0 _2332_.vdd
rlabel metal2 493 4633 507 4647 0 _2332_.A
rlabel metal2 473 4673 487 4687 0 _2332_.Y
rlabel metal1 284 4562 356 4578 0 _2316_.gnd
rlabel metal1 284 4802 356 4818 0 _2316_.vdd
rlabel metal2 333 4633 347 4647 0 _2316_.A
rlabel metal2 313 4673 327 4687 0 _2316_.Y
rlabel metal1 344 4562 456 4578 0 _2337_.gnd
rlabel metal1 344 4802 456 4818 0 _2337_.vdd
rlabel metal2 433 4673 447 4687 0 _2337_.A
rlabel metal2 413 4633 427 4647 0 _2337_.B
rlabel metal2 393 4673 407 4687 0 _2337_.C
rlabel metal2 373 4653 387 4667 0 _2337_.Y
rlabel metal1 764 4562 856 4578 0 BUFX2_insert21.gnd
rlabel metal1 764 4802 856 4818 0 BUFX2_insert21.vdd
rlabel metal2 833 4653 847 4667 0 BUFX2_insert21.A
rlabel metal2 793 4653 807 4667 0 BUFX2_insert21.Y
rlabel metal1 684 4562 776 4578 0 _2330_.gnd
rlabel metal1 684 4802 776 4818 0 _2330_.vdd
rlabel metal2 733 4653 747 4667 0 _2330_.B
rlabel metal2 693 4653 707 4667 0 _2330_.A
rlabel metal2 713 4633 727 4647 0 _2330_.Y
rlabel metal1 584 4562 696 4578 0 _2329_.gnd
rlabel metal1 584 4802 696 4818 0 _2329_.vdd
rlabel metal2 673 4653 687 4667 0 _2329_.A
rlabel metal2 613 4653 627 4667 0 _2329_.Y
rlabel metal2 633 4693 647 4707 0 _2329_.B
rlabel metal1 924 4562 1176 4578 0 _2381_.gnd
rlabel metal1 924 4802 1176 4818 0 _2381_.vdd
rlabel metal2 1073 4653 1087 4667 0 _2381_.D
rlabel metal2 1033 4653 1047 4667 0 _2381_.CLK
rlabel metal2 953 4653 967 4667 0 _2381_.Q
rlabel metal1 844 4562 936 4578 0 _2191_.gnd
rlabel metal1 844 4802 936 4818 0 _2191_.vdd
rlabel metal2 913 4693 927 4707 0 _2191_.A
rlabel metal2 873 4693 887 4707 0 _2191_.B
rlabel metal2 893 4673 907 4687 0 _2191_.Y
rlabel metal1 1164 4562 1276 4578 0 _2192_.gnd
rlabel metal1 1164 4802 1276 4818 0 _2192_.vdd
rlabel metal2 1253 4653 1267 4667 0 _2192_.A
rlabel metal2 1233 4673 1247 4687 0 _2192_.B
rlabel metal2 1193 4673 1207 4687 0 _2192_.C
rlabel metal2 1213 4653 1227 4667 0 _2192_.Y
rlabel metal1 1264 4562 1356 4578 0 _2190_.gnd
rlabel metal1 1264 4802 1356 4818 0 _2190_.vdd
rlabel metal2 1333 4693 1347 4707 0 _2190_.A
rlabel metal2 1293 4693 1307 4707 0 _2190_.B
rlabel metal2 1313 4673 1327 4687 0 _2190_.Y
rlabel metal1 1424 4562 1536 4578 0 _2189_.gnd
rlabel metal1 1424 4802 1536 4818 0 _2189_.vdd
rlabel metal2 1513 4653 1527 4667 0 _2189_.A
rlabel metal2 1493 4673 1507 4687 0 _2189_.B
rlabel metal2 1453 4673 1467 4687 0 _2189_.C
rlabel metal2 1473 4653 1487 4667 0 _2189_.Y
rlabel metal1 1524 4562 1616 4578 0 _2187_.gnd
rlabel metal1 1524 4802 1616 4818 0 _2187_.vdd
rlabel metal2 1573 4653 1587 4667 0 _2187_.B
rlabel metal2 1533 4653 1547 4667 0 _2187_.A
rlabel metal2 1553 4633 1567 4647 0 _2187_.Y
rlabel metal1 1604 4562 1696 4578 0 _2186_.gnd
rlabel metal1 1604 4802 1696 4818 0 _2186_.vdd
rlabel metal2 1653 4653 1667 4667 0 _2186_.B
rlabel metal2 1613 4653 1627 4667 0 _2186_.A
rlabel metal2 1633 4633 1647 4647 0 _2186_.Y
rlabel metal1 1344 4562 1436 4578 0 _2188_.gnd
rlabel metal1 1344 4802 1436 4818 0 _2188_.vdd
rlabel metal2 1353 4693 1367 4707 0 _2188_.A
rlabel metal2 1393 4693 1407 4707 0 _2188_.B
rlabel metal2 1373 4673 1387 4687 0 _2188_.Y
rlabel metal1 1824 4562 1936 4578 0 _2193_.gnd
rlabel metal1 1824 4802 1936 4818 0 _2193_.vdd
rlabel metal2 1833 4653 1847 4667 0 _2193_.A
rlabel metal2 1853 4673 1867 4687 0 _2193_.B
rlabel metal2 1893 4673 1907 4687 0 _2193_.C
rlabel metal2 1873 4653 1887 4667 0 _2193_.Y
rlabel metal1 1744 4562 1836 4578 0 _2185_.gnd
rlabel metal1 1744 4802 1836 4818 0 _2185_.vdd
rlabel metal2 1793 4653 1807 4667 0 _2185_.B
rlabel metal2 1753 4653 1767 4667 0 _2185_.A
rlabel metal2 1773 4633 1787 4647 0 _2185_.Y
rlabel metal1 1684 4562 1756 4578 0 _2184_.gnd
rlabel metal1 1684 4802 1756 4818 0 _2184_.vdd
rlabel metal2 1693 4633 1707 4647 0 _2184_.A
rlabel metal2 1713 4673 1727 4687 0 _2184_.Y
rlabel metal1 1924 4562 2176 4578 0 _2382_.gnd
rlabel metal1 1924 4802 2176 4818 0 _2382_.vdd
rlabel metal2 2073 4653 2087 4667 0 _2382_.D
rlabel metal2 2033 4653 2047 4667 0 _2382_.CLK
rlabel metal2 1953 4653 1967 4667 0 _2382_.Q
rlabel metal1 2164 4562 2256 4578 0 _2200_.gnd
rlabel metal1 2164 4802 2256 4818 0 _2200_.vdd
rlabel metal2 2233 4693 2247 4707 0 _2200_.A
rlabel metal2 2193 4693 2207 4707 0 _2200_.B
rlabel metal2 2213 4673 2227 4687 0 _2200_.Y
rlabel metal1 2344 4562 2436 4578 0 _2198_.gnd
rlabel metal1 2344 4802 2436 4818 0 _2198_.vdd
rlabel metal2 2353 4693 2367 4707 0 _2198_.A
rlabel metal2 2393 4693 2407 4707 0 _2198_.B
rlabel metal2 2373 4673 2387 4687 0 _2198_.Y
rlabel metal1 2244 4562 2356 4578 0 _2199_.gnd
rlabel metal1 2244 4802 2356 4818 0 _2199_.vdd
rlabel metal2 2333 4633 2347 4647 0 _2199_.A
rlabel metal2 2313 4653 2327 4667 0 _2199_.B
rlabel metal2 2273 4673 2287 4687 0 _2199_.Y
rlabel metal1 2664 4562 2916 4578 0 _2367_.gnd
rlabel metal1 2664 4802 2916 4818 0 _2367_.vdd
rlabel metal2 2813 4653 2827 4667 0 _2367_.D
rlabel metal2 2773 4653 2787 4667 0 _2367_.CLK
rlabel metal2 2693 4653 2707 4667 0 _2367_.Q
rlabel metal1 2424 4562 2516 4578 0 _2197_.gnd
rlabel metal1 2424 4802 2516 4818 0 _2197_.vdd
rlabel metal2 2473 4653 2487 4667 0 _2197_.B
rlabel metal2 2433 4653 2447 4667 0 _2197_.A
rlabel metal2 2453 4633 2467 4647 0 _2197_.Y
rlabel metal1 2604 4562 2676 4578 0 _1710_.gnd
rlabel metal1 2604 4802 2676 4818 0 _1710_.vdd
rlabel metal2 2653 4633 2667 4647 0 _1710_.A
rlabel metal2 2633 4673 2647 4687 0 _1710_.Y
rlabel metal1 2504 4562 2616 4578 0 _2203_.gnd
rlabel metal1 2504 4802 2616 4818 0 _2203_.vdd
rlabel metal2 2513 4673 2527 4687 0 _2203_.A
rlabel metal2 2533 4633 2547 4647 0 _2203_.B
rlabel metal2 2553 4673 2567 4687 0 _2203_.C
rlabel metal2 2573 4653 2587 4667 0 _2203_.Y
rlabel metal1 2904 4562 3016 4578 0 _1717_.gnd
rlabel metal1 2904 4802 3016 4818 0 _1717_.vdd
rlabel metal2 2913 4653 2927 4667 0 _1717_.A
rlabel metal2 2933 4673 2947 4687 0 _1717_.B
rlabel metal2 2973 4673 2987 4687 0 _1717_.C
rlabel metal2 2953 4653 2967 4667 0 _1717_.Y
rlabel metal1 3004 4562 3256 4578 0 _2366_.gnd
rlabel metal1 3004 4802 3256 4818 0 _2366_.vdd
rlabel metal2 3153 4653 3167 4667 0 _2366_.D
rlabel metal2 3113 4653 3127 4667 0 _2366_.CLK
rlabel metal2 3033 4653 3047 4667 0 _2366_.Q
rlabel metal1 3244 4562 3496 4578 0 _2356_.gnd
rlabel metal1 3244 4802 3496 4818 0 _2356_.vdd
rlabel metal2 3393 4653 3407 4667 0 _2356_.D
rlabel metal2 3353 4653 3367 4667 0 _2356_.CLK
rlabel metal2 3273 4653 3287 4667 0 _2356_.Q
rlabel metal1 3724 4562 3836 4578 0 _1682_.gnd
rlabel metal1 3724 4802 3836 4818 0 _1682_.vdd
rlabel metal2 3813 4653 3827 4667 0 _1682_.A
rlabel metal2 3793 4673 3807 4687 0 _1682_.B
rlabel metal2 3753 4673 3767 4687 0 _1682_.C
rlabel metal2 3773 4653 3787 4667 0 _1682_.Y
rlabel metal1 3484 4562 3596 4578 0 _1679_.gnd
rlabel metal1 3484 4802 3596 4818 0 _1679_.vdd
rlabel metal2 3573 4653 3587 4667 0 _1679_.A
rlabel metal2 3553 4673 3567 4687 0 _1679_.B
rlabel metal2 3513 4673 3527 4687 0 _1679_.C
rlabel metal2 3533 4653 3547 4667 0 _1679_.Y
rlabel metal1 3644 4562 3736 4578 0 _1681_.gnd
rlabel metal1 3644 4802 3736 4818 0 _1681_.vdd
rlabel metal2 3713 4693 3727 4707 0 _1681_.A
rlabel metal2 3673 4693 3687 4707 0 _1681_.B
rlabel metal2 3693 4673 3707 4687 0 _1681_.Y
rlabel metal1 3584 4562 3656 4578 0 _1677_.gnd
rlabel metal1 3584 4802 3656 4818 0 _1677_.vdd
rlabel metal2 3633 4673 3647 4687 0 _1677_.A
rlabel metal2 3613 4653 3627 4667 0 _1677_.Y
rlabel metal1 3824 4562 4076 4578 0 _2357_.gnd
rlabel metal1 3824 4802 4076 4818 0 _2357_.vdd
rlabel metal2 3913 4653 3927 4667 0 _2357_.D
rlabel metal2 3953 4653 3967 4667 0 _2357_.CLK
rlabel metal2 4033 4653 4047 4667 0 _2357_.Q
rlabel metal1 4204 4562 4456 4578 0 _2365_.gnd
rlabel metal1 4204 4802 4456 4818 0 _2365_.vdd
rlabel metal2 4353 4653 4367 4667 0 _2365_.D
rlabel metal2 4313 4653 4327 4667 0 _2365_.CLK
rlabel metal2 4233 4653 4247 4667 0 _2365_.Q
rlabel metal1 4124 4562 4216 4578 0 _1927_.gnd
rlabel metal1 4124 4802 4216 4818 0 _1927_.vdd
rlabel metal2 4193 4693 4207 4707 0 _1927_.A
rlabel metal2 4153 4693 4167 4707 0 _1927_.B
rlabel metal2 4173 4673 4187 4687 0 _1927_.Y
rlabel metal1 4064 4562 4136 4578 0 _1704_.gnd
rlabel metal1 4064 4802 4136 4818 0 _1704_.vdd
rlabel metal2 4113 4673 4127 4687 0 _1704_.A
rlabel metal2 4093 4653 4107 4667 0 _1704_.Y
rlabel metal1 4444 4562 4556 4578 0 _1716_.gnd
rlabel metal1 4444 4802 4556 4818 0 _1716_.vdd
rlabel metal2 4533 4673 4547 4687 0 _1716_.A
rlabel metal2 4513 4693 4527 4707 0 _1716_.B
rlabel metal2 4493 4673 4507 4687 0 _1716_.C
rlabel metal2 4473 4693 4487 4707 0 _1716_.Y
rlabel metal1 4724 4562 4836 4578 0 _1715_.gnd
rlabel metal1 4724 4802 4836 4818 0 _1715_.vdd
rlabel metal2 4733 4653 4747 4667 0 _1715_.A
rlabel metal2 4753 4673 4767 4687 0 _1715_.B
rlabel metal2 4793 4673 4807 4687 0 _1715_.C
rlabel metal2 4773 4653 4787 4667 0 _1715_.Y
rlabel metal1 4544 4562 4616 4578 0 _1714_.gnd
rlabel metal1 4544 4802 4616 4818 0 _1714_.vdd
rlabel metal2 4553 4633 4567 4647 0 _1714_.A
rlabel metal2 4573 4673 4587 4687 0 _1714_.Y
rlabel metal1 4664 4562 4736 4578 0 _1665_.gnd
rlabel metal1 4664 4802 4736 4818 0 _1665_.vdd
rlabel metal2 4713 4633 4727 4647 0 _1665_.A
rlabel metal2 4693 4673 4707 4687 0 _1665_.Y
rlabel metal1 4604 4562 4676 4578 0 _1674_.gnd
rlabel metal1 4604 4802 4676 4818 0 _1674_.vdd
rlabel metal2 4613 4673 4627 4687 0 _1674_.A
rlabel metal2 4633 4653 4647 4667 0 _1674_.Y
rlabel metal1 4824 4562 4916 4578 0 _1713_.gnd
rlabel metal1 4824 4802 4916 4818 0 _1713_.vdd
rlabel metal2 4873 4653 4887 4667 0 _1713_.B
rlabel metal2 4833 4653 4847 4667 0 _1713_.A
rlabel metal2 4853 4633 4867 4647 0 _1713_.Y
rlabel metal1 5064 4562 5156 4578 0 _1764_.gnd
rlabel metal1 5064 4802 5156 4818 0 _1764_.vdd
rlabel metal2 5133 4693 5147 4707 0 _1764_.A
rlabel metal2 5093 4693 5107 4707 0 _1764_.B
rlabel metal2 5113 4673 5127 4687 0 _1764_.Y
rlabel metal1 4904 4562 4996 4578 0 _1712_.gnd
rlabel metal1 4904 4802 4996 4818 0 _1712_.vdd
rlabel metal2 4913 4693 4927 4707 0 _1712_.A
rlabel metal2 4953 4693 4967 4707 0 _1712_.B
rlabel metal2 4933 4673 4947 4687 0 _1712_.Y
rlabel metal1 4984 4562 5076 4578 0 _1711_.gnd
rlabel metal1 4984 4802 5076 4818 0 _1711_.vdd
rlabel metal2 4993 4693 5007 4707 0 _1711_.A
rlabel metal2 5033 4693 5047 4707 0 _1711_.B
rlabel metal2 5013 4673 5027 4687 0 _1711_.Y
rlabel metal1 5244 4562 5376 4578 0 _1719_.gnd
rlabel metal1 5244 4802 5376 4818 0 _1719_.vdd
rlabel metal2 5353 4653 5367 4667 0 _1719_.A
rlabel metal2 5333 4673 5347 4687 0 _1719_.B
rlabel metal2 5273 4653 5287 4667 0 _1719_.C
rlabel metal2 5313 4653 5327 4667 0 _1719_.Y
rlabel metal2 5293 4673 5307 4687 0 _1719_.D
rlabel metal1 5144 4562 5256 4578 0 _1765_.gnd
rlabel metal1 5144 4802 5256 4818 0 _1765_.vdd
rlabel metal2 5153 4653 5167 4667 0 _1765_.A
rlabel metal2 5173 4673 5187 4687 0 _1765_.B
rlabel metal2 5213 4673 5227 4687 0 _1765_.C
rlabel metal2 5193 4653 5207 4667 0 _1765_.Y
rlabel metal1 5364 4562 5456 4578 0 _1801_.gnd
rlabel metal1 5364 4802 5456 4818 0 _1801_.vdd
rlabel metal2 5373 4693 5387 4707 0 _1801_.A
rlabel metal2 5413 4693 5427 4707 0 _1801_.B
rlabel metal2 5393 4673 5407 4687 0 _1801_.Y
rlabel metal1 5444 4562 5536 4578 0 _1760_.gnd
rlabel metal1 5444 4802 5536 4818 0 _1760_.vdd
rlabel metal2 5513 4693 5527 4707 0 _1760_.A
rlabel metal2 5473 4693 5487 4707 0 _1760_.B
rlabel metal2 5493 4673 5507 4687 0 _1760_.Y
rlabel metal1 5524 4562 5636 4578 0 _1767_.gnd
rlabel metal1 5524 4802 5636 4818 0 _1767_.vdd
rlabel metal2 5533 4673 5547 4687 0 _1767_.A
rlabel metal2 5553 4693 5567 4707 0 _1767_.B
rlabel metal2 5573 4673 5587 4687 0 _1767_.C
rlabel metal2 5593 4693 5607 4707 0 _1767_.Y
rlabel metal1 5804 4562 5876 4578 0 _1761_.gnd
rlabel metal1 5804 4802 5876 4818 0 _1761_.vdd
rlabel metal2 5853 4633 5867 4647 0 _1761_.A
rlabel metal2 5833 4673 5847 4687 0 _1761_.Y
rlabel metal1 5624 4562 5716 4578 0 _1763_.gnd
rlabel metal1 5624 4802 5716 4818 0 _1763_.vdd
rlabel metal2 5693 4693 5707 4707 0 _1763_.A
rlabel metal2 5653 4693 5667 4707 0 _1763_.B
rlabel metal2 5673 4673 5687 4687 0 _1763_.Y
rlabel metal1 5864 4562 5976 4578 0 _1770_.gnd
rlabel metal1 5864 4802 5976 4818 0 _1770_.vdd
rlabel metal2 5873 4673 5887 4687 0 _1770_.A
rlabel metal2 5893 4693 5907 4707 0 _1770_.B
rlabel metal2 5913 4673 5927 4687 0 _1770_.C
rlabel metal2 5933 4693 5947 4707 0 _1770_.Y
rlabel metal1 5704 4562 5816 4578 0 _1766_.gnd
rlabel metal1 5704 4802 5816 4818 0 _1766_.vdd
rlabel metal2 5713 4673 5727 4687 0 _1766_.A
rlabel metal2 5733 4693 5747 4707 0 _1766_.B
rlabel metal2 5753 4673 5767 4687 0 _1766_.C
rlabel metal2 5773 4693 5787 4707 0 _1766_.Y
rlabel metal1 6064 4562 6176 4578 0 _1802_.gnd
rlabel metal1 6064 4802 6176 4818 0 _1802_.vdd
rlabel metal2 6073 4653 6087 4667 0 _1802_.A
rlabel metal2 6093 4673 6107 4687 0 _1802_.B
rlabel metal2 6133 4673 6147 4687 0 _1802_.C
rlabel metal2 6113 4653 6127 4667 0 _1802_.Y
rlabel metal1 5964 4562 6076 4578 0 _1745_.gnd
rlabel metal1 5964 4802 6076 4818 0 _1745_.vdd
rlabel metal2 6053 4653 6067 4667 0 _1745_.A
rlabel metal2 5993 4653 6007 4667 0 _1745_.Y
rlabel metal2 6013 4693 6027 4707 0 _1745_.B
rlabel metal1 6164 4562 6256 4578 0 _1775_.gnd
rlabel metal1 6164 4802 6256 4818 0 _1775_.vdd
rlabel metal2 6233 4693 6247 4707 0 _1775_.A
rlabel metal2 6193 4693 6207 4707 0 _1775_.B
rlabel metal2 6213 4673 6227 4687 0 _1775_.Y
rlabel metal1 6244 4562 6356 4578 0 _1781_.gnd
rlabel metal1 6244 4802 6356 4818 0 _1781_.vdd
rlabel metal2 6253 4673 6267 4687 0 _1781_.A
rlabel metal2 6273 4633 6287 4647 0 _1781_.B
rlabel metal2 6293 4673 6307 4687 0 _1781_.C
rlabel metal2 6313 4653 6327 4667 0 _1781_.Y
rlabel metal1 6344 4562 6456 4578 0 _1774_.gnd
rlabel metal1 6344 4802 6456 4818 0 _1774_.vdd
rlabel metal2 6353 4673 6367 4687 0 _1774_.A
rlabel metal2 6373 4693 6387 4707 0 _1774_.B
rlabel metal2 6393 4673 6407 4687 0 _1774_.C
rlabel metal2 6413 4693 6427 4707 0 _1774_.Y
rlabel nsubstratencontact 6676 4808 6676 4808 0 FILL100050x68550.vdd
rlabel metal1 6664 4562 6696 4578 0 FILL100050x68550.gnd
rlabel nsubstratencontact 6656 4808 6656 4808 0 FILL99750x68550.vdd
rlabel metal1 6644 4562 6676 4578 0 FILL99750x68550.gnd
rlabel metal1 6544 4562 6656 4578 0 _1779_.gnd
rlabel metal1 6544 4802 6656 4818 0 _1779_.vdd
rlabel metal2 6633 4673 6647 4687 0 _1779_.A
rlabel metal2 6613 4693 6627 4707 0 _1779_.B
rlabel metal2 6593 4673 6607 4687 0 _1779_.C
rlabel metal2 6573 4693 6587 4707 0 _1779_.Y
rlabel metal1 6444 4562 6556 4578 0 _1844_.gnd
rlabel metal1 6444 4802 6556 4818 0 _1844_.vdd
rlabel metal2 6533 4653 6547 4667 0 _1844_.A
rlabel metal2 6473 4653 6487 4667 0 _1844_.Y
rlabel metal2 6493 4693 6507 4707 0 _1844_.B
rlabel nsubstratencontact 6716 4808 6716 4808 0 FILL100650x68550.vdd
rlabel metal1 6704 4562 6736 4578 0 FILL100650x68550.gnd
rlabel nsubstratencontact 6696 4808 6696 4808 0 FILL100350x68550.vdd
rlabel metal1 6684 4562 6716 4578 0 FILL100350x68550.gnd
rlabel metal1 4 5042 96 5058 0 _3039_.gnd
rlabel metal1 4 4802 96 4818 0 _3039_.vdd
rlabel metal2 73 4953 87 4967 0 _3039_.A
rlabel metal2 33 4953 47 4967 0 _3039_.Y
rlabel metal1 84 5042 176 5058 0 _3032_.gnd
rlabel metal1 84 4802 176 4818 0 _3032_.vdd
rlabel metal2 153 4953 167 4967 0 _3032_.A
rlabel metal2 113 4953 127 4967 0 _3032_.Y
rlabel metal1 244 5042 496 5058 0 _1609_.gnd
rlabel metal1 244 4802 496 4818 0 _1609_.vdd
rlabel metal2 393 4953 407 4967 0 _1609_.D
rlabel metal2 353 4953 367 4967 0 _1609_.CLK
rlabel metal2 273 4953 287 4967 0 _1609_.Q
rlabel metal1 164 5042 256 5058 0 _1513_.gnd
rlabel metal1 164 4802 256 4818 0 _1513_.vdd
rlabel metal2 233 4913 247 4927 0 _1513_.A
rlabel metal2 193 4913 207 4927 0 _1513_.B
rlabel metal2 213 4933 227 4947 0 _1513_.Y
rlabel metal1 484 5042 596 5058 0 _1577_.gnd
rlabel metal1 484 4802 596 4818 0 _1577_.vdd
rlabel metal2 573 4933 587 4947 0 _1577_.A
rlabel metal2 553 4973 567 4987 0 _1577_.B
rlabel metal2 533 4933 547 4947 0 _1577_.C
rlabel metal2 513 4953 527 4967 0 _1577_.Y
rlabel metal1 744 5042 836 5058 0 _1516_.gnd
rlabel metal1 744 4802 836 4818 0 _1516_.vdd
rlabel metal2 813 4913 827 4927 0 _1516_.A
rlabel metal2 773 4913 787 4927 0 _1516_.B
rlabel metal2 793 4933 807 4947 0 _1516_.Y
rlabel metal1 584 5042 676 5058 0 _1515_.gnd
rlabel metal1 584 4802 676 4818 0 _1515_.vdd
rlabel metal2 653 4913 667 4927 0 _1515_.A
rlabel metal2 613 4913 627 4927 0 _1515_.B
rlabel metal2 633 4933 647 4947 0 _1515_.Y
rlabel metal1 664 5042 756 5058 0 _1514_.gnd
rlabel metal1 664 4802 756 4818 0 _1514_.vdd
rlabel metal2 673 4913 687 4927 0 _1514_.A
rlabel metal2 713 4913 727 4927 0 _1514_.B
rlabel metal2 693 4933 707 4947 0 _1514_.Y
rlabel metal1 1064 5042 1156 5058 0 BUFX2_insert0.gnd
rlabel metal1 1064 4802 1156 4818 0 BUFX2_insert0.vdd
rlabel metal2 1133 4953 1147 4967 0 BUFX2_insert0.A
rlabel metal2 1093 4953 1107 4967 0 BUFX2_insert0.Y
rlabel metal1 824 5042 1076 5058 0 _1610_.gnd
rlabel metal1 824 4802 1076 4818 0 _1610_.vdd
rlabel metal2 973 4953 987 4967 0 _1610_.D
rlabel metal2 933 4953 947 4967 0 _1610_.CLK
rlabel metal2 853 4953 867 4967 0 _1610_.Q
rlabel metal1 1324 5042 1416 5058 0 BUFX2_insert4.gnd
rlabel metal1 1324 4802 1416 4818 0 BUFX2_insert4.vdd
rlabel metal2 1393 4953 1407 4967 0 BUFX2_insert4.A
rlabel metal2 1353 4953 1367 4967 0 BUFX2_insert4.Y
rlabel metal1 1244 5042 1336 5058 0 _1518_.gnd
rlabel metal1 1244 4802 1336 4818 0 _1518_.vdd
rlabel metal2 1313 4913 1327 4927 0 _1518_.A
rlabel metal2 1273 4913 1287 4927 0 _1518_.B
rlabel metal2 1293 4933 1307 4947 0 _1518_.Y
rlabel metal1 1144 5042 1256 5058 0 _1578_.gnd
rlabel metal1 1144 4802 1256 4818 0 _1578_.vdd
rlabel metal2 1233 4933 1247 4947 0 _1578_.A
rlabel metal2 1213 4973 1227 4987 0 _1578_.B
rlabel metal2 1193 4933 1207 4947 0 _1578_.C
rlabel metal2 1173 4953 1187 4967 0 _1578_.Y
rlabel metal1 1564 5042 1676 5058 0 _2202_.gnd
rlabel metal1 1564 4802 1676 4818 0 _2202_.vdd
rlabel metal2 1653 4953 1667 4967 0 _2202_.A
rlabel metal2 1633 4933 1647 4947 0 _2202_.B
rlabel metal2 1593 4933 1607 4947 0 _2202_.C
rlabel metal2 1613 4953 1627 4967 0 _2202_.Y
rlabel metal1 1484 5042 1576 5058 0 _2201_.gnd
rlabel metal1 1484 4802 1576 4818 0 _2201_.vdd
rlabel metal2 1553 4913 1567 4927 0 _2201_.A
rlabel metal2 1513 4913 1527 4927 0 _2201_.B
rlabel metal2 1533 4933 1547 4947 0 _2201_.Y
rlabel metal1 1404 5042 1496 5058 0 _1517_.gnd
rlabel metal1 1404 4802 1496 4818 0 _1517_.vdd
rlabel metal2 1413 4913 1427 4927 0 _1517_.A
rlabel metal2 1453 4913 1467 4927 0 _1517_.B
rlabel metal2 1433 4933 1447 4947 0 _1517_.Y
rlabel metal1 1744 5042 1856 5058 0 _1851_.gnd
rlabel metal1 1744 4802 1856 4818 0 _1851_.vdd
rlabel metal2 1833 4953 1847 4967 0 _1851_.A
rlabel metal2 1813 4933 1827 4947 0 _1851_.B
rlabel metal2 1773 4933 1787 4947 0 _1851_.C
rlabel metal2 1793 4953 1807 4967 0 _1851_.Y
rlabel metal1 1844 5042 1936 5058 0 _1850_.gnd
rlabel metal1 1844 4802 1936 4818 0 _1850_.vdd
rlabel metal2 1853 4913 1867 4927 0 _1850_.A
rlabel metal2 1893 4913 1907 4927 0 _1850_.B
rlabel metal2 1873 4933 1887 4947 0 _1850_.Y
rlabel metal1 1664 5042 1756 5058 0 _1798_.gnd
rlabel metal1 1664 4802 1756 4818 0 _1798_.vdd
rlabel metal2 1733 4913 1747 4927 0 _1798_.A
rlabel metal2 1693 4913 1707 4927 0 _1798_.B
rlabel metal2 1713 4933 1727 4947 0 _1798_.Y
rlabel metal1 1924 5042 2036 5058 0 _1916_.gnd
rlabel metal1 1924 4802 2036 4818 0 _1916_.vdd
rlabel metal2 2013 4953 2027 4967 0 _1916_.A
rlabel metal2 1993 4933 2007 4947 0 _1916_.B
rlabel metal2 1953 4933 1967 4947 0 _1916_.C
rlabel metal2 1973 4953 1987 4967 0 _1916_.Y
rlabel metal1 2024 5042 2136 5058 0 _1915_.gnd
rlabel metal1 2024 4802 2136 4818 0 _1915_.vdd
rlabel metal2 2113 4953 2127 4967 0 _1915_.A
rlabel metal2 2093 4933 2107 4947 0 _1915_.B
rlabel metal2 2053 4933 2067 4947 0 _1915_.C
rlabel metal2 2073 4953 2087 4967 0 _1915_.Y
rlabel metal1 2124 5042 2236 5058 0 _2158_.gnd
rlabel metal1 2124 4802 2236 4818 0 _2158_.vdd
rlabel metal2 2213 4953 2227 4967 0 _2158_.A
rlabel metal2 2153 4953 2167 4967 0 _2158_.Y
rlabel metal2 2173 4913 2187 4927 0 _2158_.B
rlabel metal1 2284 5042 2376 5058 0 _2174_.gnd
rlabel metal1 2284 4802 2376 4818 0 _2174_.vdd
rlabel metal2 2313 4953 2327 4967 0 _2174_.B
rlabel metal2 2353 4953 2367 4967 0 _2174_.A
rlabel metal2 2333 4973 2347 4987 0 _2174_.Y
rlabel metal1 2224 5042 2296 5058 0 _2172_.gnd
rlabel metal1 2224 4802 2296 4818 0 _2172_.vdd
rlabel metal2 2233 4973 2247 4987 0 _2172_.A
rlabel metal2 2253 4933 2267 4947 0 _2172_.Y
rlabel metal1 2364 5042 2476 5058 0 _2157_.gnd
rlabel metal1 2364 4802 2476 4818 0 _2157_.vdd
rlabel metal2 2453 4973 2467 4987 0 _2157_.A
rlabel metal2 2433 4953 2447 4967 0 _2157_.B
rlabel metal2 2393 4933 2407 4947 0 _2157_.Y
rlabel metal1 2544 5042 2656 5058 0 _2173_.gnd
rlabel metal1 2544 4802 2656 4818 0 _2173_.vdd
rlabel metal2 2633 4953 2647 4967 0 _2173_.A
rlabel metal2 2613 4933 2627 4947 0 _2173_.B
rlabel metal2 2573 4933 2587 4947 0 _2173_.C
rlabel metal2 2593 4953 2607 4967 0 _2173_.Y
rlabel metal1 2644 5042 2756 5058 0 _2156_.gnd
rlabel metal1 2644 4802 2756 4818 0 _2156_.vdd
rlabel metal2 2733 4953 2747 4967 0 _2156_.A
rlabel metal2 2713 4933 2727 4947 0 _2156_.B
rlabel metal2 2673 4933 2687 4947 0 _2156_.C
rlabel metal2 2693 4953 2707 4967 0 _2156_.Y
rlabel metal1 2464 5042 2556 5058 0 _1853_.gnd
rlabel metal1 2464 4802 2556 4818 0 _1853_.vdd
rlabel metal2 2533 4913 2547 4927 0 _1853_.A
rlabel metal2 2493 4913 2507 4927 0 _1853_.B
rlabel metal2 2513 4933 2527 4947 0 _1853_.Y
rlabel metal1 2904 5042 3016 5058 0 _2155_.gnd
rlabel metal1 2904 4802 3016 4818 0 _2155_.vdd
rlabel metal2 2993 4953 3007 4967 0 _2155_.A
rlabel metal2 2973 4933 2987 4947 0 _2155_.B
rlabel metal2 2933 4933 2947 4947 0 _2155_.C
rlabel metal2 2953 4953 2967 4967 0 _2155_.Y
rlabel metal1 2804 5042 2916 5058 0 _2129_.gnd
rlabel metal1 2804 4802 2916 4818 0 _2129_.vdd
rlabel metal2 2813 4953 2827 4967 0 _2129_.A
rlabel metal2 2833 4933 2847 4947 0 _2129_.B
rlabel metal2 2873 4933 2887 4947 0 _2129_.C
rlabel metal2 2853 4953 2867 4967 0 _2129_.Y
rlabel metal1 2744 5042 2816 5058 0 _2127_.gnd
rlabel metal1 2744 4802 2816 4818 0 _2127_.vdd
rlabel metal2 2793 4973 2807 4987 0 _2127_.A
rlabel metal2 2773 4933 2787 4947 0 _2127_.Y
rlabel metal1 3004 5042 3116 5058 0 _2128_.gnd
rlabel metal1 3004 4802 3116 4818 0 _2128_.vdd
rlabel metal2 3093 4953 3107 4967 0 _2128_.A
rlabel metal2 3073 4933 3087 4947 0 _2128_.B
rlabel metal2 3033 4933 3047 4947 0 _2128_.C
rlabel metal2 3053 4953 3067 4967 0 _2128_.Y
rlabel metal1 3104 5042 3196 5058 0 _2126_.gnd
rlabel metal1 3104 4802 3196 4818 0 _2126_.vdd
rlabel metal2 3133 4953 3147 4967 0 _2126_.B
rlabel metal2 3173 4953 3187 4967 0 _2126_.A
rlabel metal2 3153 4973 3167 4987 0 _2126_.Y
rlabel metal1 3184 5042 3256 5058 0 _1701_.gnd
rlabel metal1 3184 4802 3256 4818 0 _1701_.vdd
rlabel metal2 3233 4933 3247 4947 0 _1701_.A
rlabel metal2 3213 4953 3227 4967 0 _1701_.Y
rlabel metal1 3424 5042 3676 5058 0 _2363_.gnd
rlabel metal1 3424 4802 3676 4818 0 _2363_.vdd
rlabel metal2 3513 4953 3527 4967 0 _2363_.D
rlabel metal2 3553 4953 3567 4967 0 _2363_.CLK
rlabel metal2 3633 4953 3647 4967 0 _2363_.Q
rlabel metal1 3324 5042 3436 5058 0 _2098_.gnd
rlabel metal1 3324 4802 3436 4818 0 _2098_.vdd
rlabel metal2 3413 4953 3427 4967 0 _2098_.A
rlabel metal2 3393 4933 3407 4947 0 _2098_.B
rlabel metal2 3353 4933 3367 4947 0 _2098_.C
rlabel metal2 3373 4953 3387 4967 0 _2098_.Y
rlabel metal1 3244 5042 3336 5058 0 _2097_.gnd
rlabel metal1 3244 4802 3336 4818 0 _2097_.vdd
rlabel metal2 3313 4913 3327 4927 0 _2097_.A
rlabel metal2 3273 4913 3287 4927 0 _2097_.B
rlabel metal2 3293 4933 3307 4947 0 _2097_.Y
rlabel metal1 3664 5042 3776 5058 0 _1700_.gnd
rlabel metal1 3664 4802 3776 4818 0 _1700_.vdd
rlabel metal2 3673 4953 3687 4967 0 _1700_.A
rlabel metal2 3693 4933 3707 4947 0 _1700_.B
rlabel metal2 3733 4933 3747 4947 0 _1700_.C
rlabel metal2 3713 4953 3727 4967 0 _1700_.Y
rlabel metal1 3964 5042 4076 5058 0 _1914_.gnd
rlabel metal1 3964 4802 4076 4818 0 _1914_.vdd
rlabel metal2 4053 4933 4067 4947 0 _1914_.A
rlabel metal2 4033 4973 4047 4987 0 _1914_.B
rlabel metal2 4013 4933 4027 4947 0 _1914_.C
rlabel metal2 3993 4953 4007 4967 0 _1914_.Y
rlabel metal1 3764 5042 3876 5058 0 _1848_.gnd
rlabel metal1 3764 4802 3876 4818 0 _1848_.vdd
rlabel metal2 3853 4933 3867 4947 0 _1848_.A
rlabel metal2 3833 4973 3847 4987 0 _1848_.B
rlabel metal2 3813 4933 3827 4947 0 _1848_.C
rlabel metal2 3793 4953 3807 4967 0 _1848_.Y
rlabel metal1 3864 5042 3976 5058 0 _1849_.gnd
rlabel metal1 3864 4802 3976 4818 0 _1849_.vdd
rlabel metal2 3953 4933 3967 4947 0 _1849_.A
rlabel metal2 3933 4913 3947 4927 0 _1849_.B
rlabel metal2 3913 4933 3927 4947 0 _1849_.C
rlabel metal2 3893 4913 3907 4927 0 _1849_.Y
rlabel metal1 4224 5042 4316 5058 0 _1858_.gnd
rlabel metal1 4224 4802 4316 4818 0 _1858_.vdd
rlabel metal2 4293 4913 4307 4927 0 _1858_.A
rlabel metal2 4253 4913 4267 4927 0 _1858_.B
rlabel metal2 4273 4933 4287 4947 0 _1858_.Y
rlabel metal1 4064 5042 4136 5058 0 _1698_.gnd
rlabel metal1 4064 4802 4136 4818 0 _1698_.vdd
rlabel metal2 4113 4933 4127 4947 0 _1698_.A
rlabel metal2 4093 4953 4107 4967 0 _1698_.Y
rlabel metal1 4124 5042 4236 5058 0 _1921_.gnd
rlabel metal1 4124 4802 4236 4818 0 _1921_.vdd
rlabel metal2 4213 4953 4227 4967 0 _1921_.A
rlabel metal2 4153 4953 4167 4967 0 _1921_.Y
rlabel metal2 4173 4913 4187 4927 0 _1921_.B
rlabel metal1 4404 5042 4516 5058 0 _1866_.gnd
rlabel metal1 4404 4802 4516 4818 0 _1866_.vdd
rlabel metal2 4493 4953 4507 4967 0 _1866_.A
rlabel metal2 4473 4933 4487 4947 0 _1866_.B
rlabel metal2 4433 4933 4447 4947 0 _1866_.C
rlabel metal2 4453 4953 4467 4967 0 _1866_.Y
rlabel metal1 4504 5042 4616 5058 0 _1868_.gnd
rlabel metal1 4504 4802 4616 4818 0 _1868_.vdd
rlabel metal2 4513 4933 4527 4947 0 _1868_.A
rlabel metal2 4533 4913 4547 4927 0 _1868_.B
rlabel metal2 4553 4933 4567 4947 0 _1868_.C
rlabel metal2 4573 4913 4587 4927 0 _1868_.Y
rlabel metal1 4304 5042 4416 5058 0 _1861_.gnd
rlabel metal1 4304 4802 4416 4818 0 _1861_.vdd
rlabel metal2 4313 4953 4327 4967 0 _1861_.A
rlabel metal2 4373 4953 4387 4967 0 _1861_.Y
rlabel metal2 4353 4913 4367 4927 0 _1861_.B
rlabel metal1 4604 5042 4716 5058 0 _1867_.gnd
rlabel metal1 4604 4802 4716 4818 0 _1867_.vdd
rlabel metal2 4613 4953 4627 4967 0 _1867_.A
rlabel metal2 4633 4933 4647 4947 0 _1867_.B
rlabel metal2 4673 4933 4687 4947 0 _1867_.C
rlabel metal2 4653 4953 4667 4967 0 _1867_.Y
rlabel metal1 4704 5042 4796 5058 0 _1862_.gnd
rlabel metal1 4704 4802 4796 4818 0 _1862_.vdd
rlabel metal2 4773 4913 4787 4927 0 _1862_.A
rlabel metal2 4733 4913 4747 4927 0 _1862_.B
rlabel metal2 4753 4933 4767 4947 0 _1862_.Y
rlabel metal1 4784 5042 4896 5058 0 _1860_.gnd
rlabel metal1 4784 4802 4896 4818 0 _1860_.vdd
rlabel metal2 4873 4953 4887 4967 0 _1860_.A
rlabel metal2 4813 4953 4827 4967 0 _1860_.Y
rlabel metal2 4833 4913 4847 4927 0 _1860_.B
rlabel metal1 4964 5042 5056 5058 0 _1863_.gnd
rlabel metal1 4964 4802 5056 4818 0 _1863_.vdd
rlabel metal2 4973 4913 4987 4927 0 _1863_.A
rlabel metal2 5013 4913 5027 4927 0 _1863_.B
rlabel metal2 4993 4933 5007 4947 0 _1863_.Y
rlabel metal1 4884 5042 4976 5058 0 _1803_.gnd
rlabel metal1 4884 4802 4976 4818 0 _1803_.vdd
rlabel metal2 4953 4913 4967 4927 0 _1803_.A
rlabel metal2 4913 4913 4927 4927 0 _1803_.B
rlabel metal2 4933 4933 4947 4947 0 _1803_.Y
rlabel metal1 5044 5042 5156 5058 0 _1805_.gnd
rlabel metal1 5044 4802 5156 4818 0 _1805_.vdd
rlabel metal2 5053 4953 5067 4967 0 _1805_.A
rlabel metal2 5113 4953 5127 4967 0 _1805_.Y
rlabel metal2 5093 4913 5107 4927 0 _1805_.B
rlabel metal1 5144 5042 5236 5058 0 _1806_.gnd
rlabel metal1 5144 4802 5236 4818 0 _1806_.vdd
rlabel metal2 5213 4913 5227 4927 0 _1806_.A
rlabel metal2 5173 4913 5187 4927 0 _1806_.B
rlabel metal2 5193 4933 5207 4947 0 _1806_.Y
rlabel metal1 5324 5042 5436 5058 0 _1771_.gnd
rlabel metal1 5324 4802 5436 4818 0 _1771_.vdd
rlabel metal2 5333 4953 5347 4967 0 _1771_.A
rlabel metal2 5393 4953 5407 4967 0 _1771_.Y
rlabel metal2 5373 4913 5387 4927 0 _1771_.B
rlabel metal1 5224 5042 5336 5058 0 _1762_.gnd
rlabel metal1 5224 4802 5336 4818 0 _1762_.vdd
rlabel metal2 5313 4953 5327 4967 0 _1762_.A
rlabel metal2 5253 4953 5267 4967 0 _1762_.Y
rlabel metal2 5273 4913 5287 4927 0 _1762_.B
rlabel metal1 5544 5042 5636 5058 0 _1768_.gnd
rlabel metal1 5544 4802 5636 4818 0 _1768_.vdd
rlabel metal2 5613 4913 5627 4927 0 _1768_.A
rlabel metal2 5573 4913 5587 4927 0 _1768_.B
rlabel metal2 5593 4933 5607 4947 0 _1768_.Y
rlabel metal1 5424 5042 5556 5058 0 _1772_.gnd
rlabel metal1 5424 4802 5556 4818 0 _1772_.vdd
rlabel metal2 5533 4953 5547 4967 0 _1772_.A
rlabel metal2 5513 4933 5527 4947 0 _1772_.B
rlabel metal2 5453 4953 5467 4967 0 _1772_.C
rlabel metal2 5473 4933 5487 4947 0 _1772_.D
rlabel metal2 5493 4953 5507 4967 0 _1772_.Y
rlabel metal1 5724 5042 5836 5058 0 _1773_.gnd
rlabel metal1 5724 4802 5836 4818 0 _1773_.vdd
rlabel metal2 5813 4933 5827 4947 0 _1773_.A
rlabel metal2 5793 4973 5807 4987 0 _1773_.B
rlabel metal2 5773 4933 5787 4947 0 _1773_.C
rlabel metal2 5753 4953 5767 4967 0 _1773_.Y
rlabel metal1 5824 5042 5936 5058 0 _1843_.gnd
rlabel metal1 5824 4802 5936 4818 0 _1843_.vdd
rlabel metal2 5913 4933 5927 4947 0 _1843_.A
rlabel metal2 5893 4913 5907 4927 0 _1843_.B
rlabel metal2 5873 4933 5887 4947 0 _1843_.C
rlabel metal2 5853 4913 5867 4927 0 _1843_.Y
rlabel metal1 5624 5042 5736 5058 0 _1769_.gnd
rlabel metal1 5624 4802 5736 4818 0 _1769_.vdd
rlabel metal2 5633 4933 5647 4947 0 _1769_.A
rlabel metal2 5653 4913 5667 4927 0 _1769_.B
rlabel metal2 5673 4933 5687 4947 0 _1769_.C
rlabel metal2 5693 4913 5707 4927 0 _1769_.Y
rlabel metal1 5924 5042 6016 5058 0 _1800_.gnd
rlabel metal1 5924 4802 6016 4818 0 _1800_.vdd
rlabel metal2 5993 4913 6007 4927 0 _1800_.A
rlabel metal2 5953 4913 5967 4927 0 _1800_.B
rlabel metal2 5973 4933 5987 4947 0 _1800_.Y
rlabel metal1 6124 5042 6236 5058 0 _1847_.gnd
rlabel metal1 6124 4802 6236 4818 0 _1847_.vdd
rlabel metal2 6213 4933 6227 4947 0 _1847_.A
rlabel metal2 6193 4913 6207 4927 0 _1847_.B
rlabel metal2 6173 4933 6187 4947 0 _1847_.C
rlabel metal2 6153 4913 6167 4927 0 _1847_.Y
rlabel metal1 6004 5042 6136 5058 0 _1913_.gnd
rlabel metal1 6004 4802 6136 4818 0 _1913_.vdd
rlabel metal2 6013 4953 6027 4967 0 _1913_.A
rlabel metal2 6033 4933 6047 4947 0 _1913_.B
rlabel metal2 6093 4953 6107 4967 0 _1913_.C
rlabel metal2 6073 4933 6087 4947 0 _1913_.D
rlabel metal2 6053 4953 6067 4967 0 _1913_.Y
rlabel metal1 6224 5042 6336 5058 0 _1778_.gnd
rlabel metal1 6224 4802 6336 4818 0 _1778_.vdd
rlabel metal2 6233 4953 6247 4967 0 _1778_.A
rlabel metal2 6253 4933 6267 4947 0 _1778_.B
rlabel metal2 6293 4933 6307 4947 0 _1778_.C
rlabel metal2 6273 4953 6287 4967 0 _1778_.Y
rlabel metal1 6324 5042 6436 5058 0 _1846_.gnd
rlabel metal1 6324 4802 6436 4818 0 _1846_.vdd
rlabel metal2 6413 4933 6427 4947 0 _1846_.A
rlabel metal2 6393 4913 6407 4927 0 _1846_.B
rlabel metal2 6373 4933 6387 4947 0 _1846_.C
rlabel metal2 6353 4913 6367 4927 0 _1846_.Y
rlabel nsubstratencontact 6684 4812 6684 4812 0 FILL100050x72150.vdd
rlabel metal1 6664 5042 6696 5058 0 FILL100050x72150.gnd
rlabel metal1 6604 5042 6676 5058 0 _1780_.gnd
rlabel metal1 6604 4802 6676 4818 0 _1780_.vdd
rlabel metal2 6653 4973 6667 4987 0 _1780_.A
rlabel metal2 6633 4933 6647 4947 0 _1780_.Y
rlabel metal1 6524 5042 6616 5058 0 _1840_.gnd
rlabel metal1 6524 4802 6616 4818 0 _1840_.vdd
rlabel metal2 6533 4913 6547 4927 0 _1840_.A
rlabel metal2 6573 4913 6587 4927 0 _1840_.B
rlabel metal2 6553 4933 6567 4947 0 _1840_.Y
rlabel metal1 6424 5042 6536 5058 0 _1842_.gnd
rlabel metal1 6424 4802 6536 4818 0 _1842_.vdd
rlabel metal2 6513 4933 6527 4947 0 _1842_.A
rlabel metal2 6493 4913 6507 4927 0 _1842_.B
rlabel metal2 6473 4933 6487 4947 0 _1842_.C
rlabel metal2 6453 4913 6467 4927 0 _1842_.Y
rlabel nsubstratencontact 6724 4812 6724 4812 0 FILL100650x72150.vdd
rlabel metal1 6704 5042 6736 5058 0 FILL100650x72150.gnd
rlabel nsubstratencontact 6704 4812 6704 4812 0 FILL100350x72150.vdd
rlabel metal1 6684 5042 6716 5058 0 FILL100350x72150.gnd
rlabel metal1 4 5042 96 5058 0 _3034_.gnd
rlabel metal1 4 5282 96 5298 0 _3034_.vdd
rlabel metal2 73 5133 87 5147 0 _3034_.A
rlabel metal2 33 5133 47 5147 0 _3034_.Y
rlabel metal1 84 5042 336 5058 0 _1619_.gnd
rlabel metal1 84 5282 336 5298 0 _1619_.vdd
rlabel metal2 233 5133 247 5147 0 _1619_.D
rlabel metal2 193 5133 207 5147 0 _1619_.CLK
rlabel metal2 113 5133 127 5147 0 _1619_.Q
rlabel metal1 504 5042 596 5058 0 _1545_.gnd
rlabel metal1 504 5282 596 5298 0 _1545_.vdd
rlabel metal2 573 5173 587 5187 0 _1545_.A
rlabel metal2 533 5173 547 5187 0 _1545_.B
rlabel metal2 553 5153 567 5167 0 _1545_.Y
rlabel metal1 324 5042 416 5058 0 _1543_.gnd
rlabel metal1 324 5282 416 5298 0 _1543_.vdd
rlabel metal2 333 5173 347 5187 0 _1543_.A
rlabel metal2 373 5173 387 5187 0 _1543_.B
rlabel metal2 353 5153 367 5167 0 _1543_.Y
rlabel metal1 404 5042 516 5058 0 _1587_.gnd
rlabel metal1 404 5282 516 5298 0 _1587_.vdd
rlabel metal2 493 5153 507 5167 0 _1587_.A
rlabel metal2 473 5113 487 5127 0 _1587_.B
rlabel metal2 453 5153 467 5167 0 _1587_.C
rlabel metal2 433 5133 447 5147 0 _1587_.Y
rlabel metal1 584 5042 836 5058 0 _2388_.gnd
rlabel metal1 584 5282 836 5298 0 _2388_.vdd
rlabel metal2 673 5133 687 5147 0 _2388_.D
rlabel metal2 713 5133 727 5147 0 _2388_.CLK
rlabel metal2 793 5133 807 5147 0 _2388_.Q
rlabel metal1 904 5042 1016 5058 0 _2272_.gnd
rlabel metal1 904 5282 1016 5298 0 _2272_.vdd
rlabel metal2 993 5133 1007 5147 0 _2272_.A
rlabel metal2 973 5153 987 5167 0 _2272_.B
rlabel metal2 933 5153 947 5167 0 _2272_.C
rlabel metal2 953 5133 967 5147 0 _2272_.Y
rlabel metal1 1004 5042 1116 5058 0 _2271_.gnd
rlabel metal1 1004 5282 1116 5298 0 _2271_.vdd
rlabel metal2 1093 5133 1107 5147 0 _2271_.A
rlabel metal2 1073 5153 1087 5167 0 _2271_.B
rlabel metal2 1033 5153 1047 5167 0 _2271_.C
rlabel metal2 1053 5133 1067 5147 0 _2271_.Y
rlabel metal1 824 5042 916 5058 0 _2258_.gnd
rlabel metal1 824 5282 916 5298 0 _2258_.vdd
rlabel metal2 833 5173 847 5187 0 _2258_.A
rlabel metal2 873 5173 887 5187 0 _2258_.B
rlabel metal2 853 5153 867 5167 0 _2258_.Y
rlabel metal1 1204 5042 1456 5058 0 _2378_.gnd
rlabel metal1 1204 5282 1456 5298 0 _2378_.vdd
rlabel metal2 1353 5133 1367 5147 0 _2378_.D
rlabel metal2 1313 5133 1327 5147 0 _2378_.CLK
rlabel metal2 1233 5133 1247 5147 0 _2378_.Q
rlabel metal1 1104 5042 1216 5058 0 _2270_.gnd
rlabel metal1 1104 5282 1216 5298 0 _2270_.vdd
rlabel metal2 1193 5133 1207 5147 0 _2270_.A
rlabel metal2 1133 5133 1147 5147 0 _2270_.Y
rlabel metal2 1153 5173 1167 5187 0 _2270_.B
rlabel metal1 1604 5042 1856 5058 0 _2379_.gnd
rlabel metal1 1604 5282 1856 5298 0 _2379_.vdd
rlabel metal2 1753 5133 1767 5147 0 _2379_.D
rlabel metal2 1713 5133 1727 5147 0 _2379_.CLK
rlabel metal2 1633 5133 1647 5147 0 _2379_.Q
rlabel metal1 1444 5042 1536 5058 0 _2170_.gnd
rlabel metal1 1444 5282 1536 5298 0 _2170_.vdd
rlabel metal2 1513 5173 1527 5187 0 _2170_.A
rlabel metal2 1473 5173 1487 5187 0 _2170_.B
rlabel metal2 1493 5153 1507 5167 0 _2170_.Y
rlabel metal1 1524 5042 1616 5058 0 _2150_.gnd
rlabel metal1 1524 5282 1616 5298 0 _2150_.vdd
rlabel metal2 1533 5173 1547 5187 0 _2150_.A
rlabel metal2 1573 5173 1587 5187 0 _2150_.B
rlabel metal2 1553 5153 1567 5167 0 _2150_.Y
rlabel metal1 1844 5042 1976 5058 0 _2176_.gnd
rlabel metal1 1844 5282 1976 5298 0 _2176_.vdd
rlabel metal2 1953 5133 1967 5147 0 _2176_.A
rlabel metal2 1933 5153 1947 5167 0 _2176_.B
rlabel metal2 1873 5133 1887 5147 0 _2176_.C
rlabel metal2 1893 5153 1907 5167 0 _2176_.D
rlabel metal2 1913 5133 1927 5147 0 _2176_.Y
rlabel metal1 1964 5042 2036 5058 0 _2171_.gnd
rlabel metal1 1964 5282 2036 5298 0 _2171_.vdd
rlabel metal2 1973 5113 1987 5127 0 _2171_.A
rlabel metal2 1993 5153 2007 5167 0 _2171_.Y
rlabel metal1 2124 5042 2216 5058 0 _2161_.gnd
rlabel metal1 2124 5282 2216 5298 0 _2161_.vdd
rlabel metal2 2133 5173 2147 5187 0 _2161_.A
rlabel metal2 2173 5173 2187 5187 0 _2161_.B
rlabel metal2 2153 5153 2167 5167 0 _2161_.Y
rlabel metal1 2024 5042 2136 5058 0 _2175_.gnd
rlabel metal1 2024 5282 2136 5298 0 _2175_.vdd
rlabel metal2 2113 5133 2127 5147 0 _2175_.A
rlabel metal2 2053 5133 2067 5147 0 _2175_.Y
rlabel metal2 2073 5173 2087 5187 0 _2175_.B
rlabel metal1 2304 5042 2396 5058 0 _2160_.gnd
rlabel metal1 2304 5282 2396 5298 0 _2160_.vdd
rlabel metal2 2373 5173 2387 5187 0 _2160_.A
rlabel metal2 2333 5173 2347 5187 0 _2160_.B
rlabel metal2 2353 5153 2367 5167 0 _2160_.Y
rlabel metal1 2384 5042 2496 5058 0 _1985_.gnd
rlabel metal1 2384 5282 2496 5298 0 _1985_.vdd
rlabel metal2 2473 5153 2487 5167 0 _1985_.A
rlabel metal2 2453 5173 2467 5187 0 _1985_.B
rlabel metal2 2433 5153 2447 5167 0 _1985_.C
rlabel metal2 2413 5173 2427 5187 0 _1985_.Y
rlabel metal1 2204 5042 2316 5058 0 _2159_.gnd
rlabel metal1 2204 5282 2316 5298 0 _2159_.vdd
rlabel metal2 2293 5113 2307 5127 0 _2159_.A
rlabel metal2 2273 5133 2287 5147 0 _2159_.B
rlabel metal2 2233 5153 2247 5167 0 _2159_.Y
rlabel metal1 2484 5042 2576 5058 0 _1912_.gnd
rlabel metal1 2484 5282 2576 5298 0 _1912_.vdd
rlabel metal2 2513 5133 2527 5147 0 _1912_.B
rlabel metal2 2553 5133 2567 5147 0 _1912_.A
rlabel metal2 2533 5113 2547 5127 0 _1912_.Y
rlabel metal1 2564 5042 2636 5058 0 _1911_.gnd
rlabel metal1 2564 5282 2636 5298 0 _1911_.vdd
rlabel metal2 2573 5113 2587 5127 0 _1911_.A
rlabel metal2 2593 5153 2607 5167 0 _1911_.Y
rlabel metal1 2624 5042 2736 5058 0 _2133_.gnd
rlabel metal1 2624 5282 2736 5298 0 _2133_.vdd
rlabel metal2 2713 5133 2727 5147 0 _2133_.A
rlabel metal2 2653 5133 2667 5147 0 _2133_.Y
rlabel metal2 2673 5173 2687 5187 0 _2133_.B
rlabel metal1 2724 5042 2816 5058 0 _2134_.gnd
rlabel metal1 2724 5282 2816 5298 0 _2134_.vdd
rlabel metal2 2773 5133 2787 5147 0 _2134_.B
rlabel metal2 2733 5133 2747 5147 0 _2134_.A
rlabel metal2 2753 5113 2767 5127 0 _2134_.Y
rlabel metal1 2804 5042 2896 5058 0 _2132_.gnd
rlabel metal1 2804 5282 2896 5298 0 _2132_.vdd
rlabel metal2 2873 5173 2887 5187 0 _2132_.A
rlabel metal2 2833 5173 2847 5187 0 _2132_.B
rlabel metal2 2853 5153 2867 5167 0 _2132_.Y
rlabel metal1 2884 5042 2976 5058 0 _2131_.gnd
rlabel metal1 2884 5282 2976 5298 0 _2131_.vdd
rlabel metal2 2953 5173 2967 5187 0 _2131_.A
rlabel metal2 2913 5173 2927 5187 0 _2131_.B
rlabel metal2 2933 5153 2947 5167 0 _2131_.Y
rlabel metal1 3164 5042 3256 5058 0 _2108_.gnd
rlabel metal1 3164 5282 3256 5298 0 _2108_.vdd
rlabel metal2 3173 5173 3187 5187 0 _2108_.A
rlabel metal2 3213 5173 3227 5187 0 _2108_.B
rlabel metal2 3193 5153 3207 5167 0 _2108_.Y
rlabel metal1 2964 5042 3076 5058 0 _2130_.gnd
rlabel metal1 2964 5282 3076 5298 0 _2130_.vdd
rlabel metal2 2973 5113 2987 5127 0 _2130_.A
rlabel metal2 2993 5133 3007 5147 0 _2130_.B
rlabel metal2 3033 5153 3047 5167 0 _2130_.Y
rlabel metal1 3064 5042 3176 5058 0 _2105_.gnd
rlabel metal1 3064 5282 3176 5298 0 _2105_.vdd
rlabel metal2 3153 5133 3167 5147 0 _2105_.A
rlabel metal2 3093 5133 3107 5147 0 _2105_.Y
rlabel metal2 3113 5173 3127 5187 0 _2105_.B
rlabel metal1 3344 5042 3416 5058 0 _2103_.gnd
rlabel metal1 3344 5282 3416 5298 0 _2103_.vdd
rlabel metal2 3393 5113 3407 5127 0 _2103_.A
rlabel metal2 3373 5153 3387 5167 0 _2103_.Y
rlabel metal1 3404 5042 3516 5058 0 _2125_.gnd
rlabel metal1 3404 5282 3516 5298 0 _2125_.vdd
rlabel metal2 3493 5153 3507 5167 0 _2125_.A
rlabel metal2 3473 5113 3487 5127 0 _2125_.B
rlabel metal2 3453 5153 3467 5167 0 _2125_.C
rlabel metal2 3433 5133 3447 5147 0 _2125_.Y
rlabel metal1 3244 5042 3356 5058 0 _2104_.gnd
rlabel metal1 3244 5282 3356 5298 0 _2104_.vdd
rlabel metal2 3333 5153 3347 5167 0 _2104_.A
rlabel metal2 3313 5173 3327 5187 0 _2104_.B
rlabel metal2 3293 5153 3307 5167 0 _2104_.C
rlabel metal2 3273 5173 3287 5187 0 _2104_.Y
rlabel metal1 3584 5042 3696 5058 0 _2100_.gnd
rlabel metal1 3584 5282 3696 5298 0 _2100_.vdd
rlabel metal2 3593 5133 3607 5147 0 _2100_.A
rlabel metal2 3613 5153 3627 5167 0 _2100_.B
rlabel metal2 3653 5153 3667 5167 0 _2100_.C
rlabel metal2 3633 5133 3647 5147 0 _2100_.Y
rlabel metal1 3684 5042 3796 5058 0 _2099_.gnd
rlabel metal1 3684 5282 3796 5298 0 _2099_.vdd
rlabel metal2 3773 5133 3787 5147 0 _2099_.A
rlabel metal2 3753 5153 3767 5167 0 _2099_.B
rlabel metal2 3713 5153 3727 5167 0 _2099_.C
rlabel metal2 3733 5133 3747 5147 0 _2099_.Y
rlabel metal1 3504 5042 3596 5058 0 _2101_.gnd
rlabel metal1 3504 5282 3596 5298 0 _2101_.vdd
rlabel metal2 3533 5133 3547 5147 0 _2101_.B
rlabel metal2 3573 5133 3587 5147 0 _2101_.A
rlabel metal2 3553 5113 3567 5127 0 _2101_.Y
rlabel metal1 3784 5042 3876 5058 0 _2102_.gnd
rlabel metal1 3784 5282 3876 5298 0 _2102_.vdd
rlabel metal2 3833 5133 3847 5147 0 _2102_.B
rlabel metal2 3793 5133 3807 5147 0 _2102_.A
rlabel metal2 3813 5113 3827 5127 0 _2102_.Y
rlabel metal1 3944 5042 4036 5058 0 _2096_.gnd
rlabel metal1 3944 5282 4036 5298 0 _2096_.vdd
rlabel metal2 4013 5173 4027 5187 0 _2096_.A
rlabel metal2 3973 5173 3987 5187 0 _2096_.B
rlabel metal2 3993 5153 4007 5167 0 _2096_.Y
rlabel metal1 3864 5042 3956 5058 0 _2049_.gnd
rlabel metal1 3864 5282 3956 5298 0 _2049_.vdd
rlabel metal2 3873 5173 3887 5187 0 _2049_.A
rlabel metal2 3913 5173 3927 5187 0 _2049_.B
rlabel metal2 3893 5153 3907 5167 0 _2049_.Y
rlabel metal1 4024 5042 4136 5058 0 _1934_.gnd
rlabel metal1 4024 5282 4136 5298 0 _1934_.vdd
rlabel metal2 4033 5133 4047 5147 0 _1934_.A
rlabel metal2 4053 5153 4067 5167 0 _1934_.B
rlabel metal2 4093 5153 4107 5167 0 _1934_.C
rlabel metal2 4073 5133 4087 5147 0 _1934_.Y
rlabel metal1 4124 5042 4216 5058 0 _2051_.gnd
rlabel metal1 4124 5282 4216 5298 0 _2051_.vdd
rlabel metal2 4193 5173 4207 5187 0 _2051_.A
rlabel metal2 4153 5173 4167 5187 0 _2051_.B
rlabel metal2 4173 5153 4187 5167 0 _2051_.Y
rlabel metal1 4204 5042 4316 5058 0 _1929_.gnd
rlabel metal1 4204 5282 4316 5298 0 _1929_.vdd
rlabel metal2 4293 5133 4307 5147 0 _1929_.A
rlabel metal2 4233 5133 4247 5147 0 _1929_.Y
rlabel metal2 4253 5173 4267 5187 0 _1929_.B
rlabel metal1 4484 5042 4596 5058 0 _2053_.gnd
rlabel metal1 4484 5282 4596 5298 0 _2053_.vdd
rlabel metal2 4573 5133 4587 5147 0 _2053_.A
rlabel metal2 4553 5153 4567 5167 0 _2053_.B
rlabel metal2 4513 5153 4527 5167 0 _2053_.C
rlabel metal2 4533 5133 4547 5147 0 _2053_.Y
rlabel metal1 4384 5042 4496 5058 0 _2052_.gnd
rlabel metal1 4384 5282 4496 5298 0 _2052_.vdd
rlabel metal2 4473 5133 4487 5147 0 _2052_.A
rlabel metal2 4453 5153 4467 5167 0 _2052_.B
rlabel metal2 4413 5153 4427 5167 0 _2052_.C
rlabel metal2 4433 5133 4447 5147 0 _2052_.Y
rlabel metal1 4304 5042 4396 5058 0 _1931_.gnd
rlabel metal1 4304 5282 4396 5298 0 _1931_.vdd
rlabel metal2 4373 5173 4387 5187 0 _1931_.A
rlabel metal2 4333 5173 4347 5187 0 _1931_.B
rlabel metal2 4353 5153 4367 5167 0 _1931_.Y
rlabel metal1 4744 5042 4816 5058 0 _1859_.gnd
rlabel metal1 4744 5282 4816 5298 0 _1859_.vdd
rlabel metal2 4753 5113 4767 5127 0 _1859_.A
rlabel metal2 4773 5153 4787 5167 0 _1859_.Y
rlabel metal1 4584 5042 4676 5058 0 _2050_.gnd
rlabel metal1 4584 5282 4676 5298 0 _2050_.vdd
rlabel metal2 4593 5173 4607 5187 0 _2050_.A
rlabel metal2 4633 5173 4647 5187 0 _2050_.B
rlabel metal2 4613 5153 4627 5167 0 _2050_.Y
rlabel metal1 4664 5042 4756 5058 0 _2001_.gnd
rlabel metal1 4664 5282 4756 5298 0 _2001_.vdd
rlabel metal2 4673 5173 4687 5187 0 _2001_.A
rlabel metal2 4713 5173 4727 5187 0 _2001_.B
rlabel metal2 4693 5153 4707 5167 0 _2001_.Y
rlabel metal1 4804 5042 4916 5058 0 _1865_.gnd
rlabel metal1 4804 5282 4916 5298 0 _1865_.vdd
rlabel metal2 4893 5153 4907 5167 0 _1865_.A
rlabel metal2 4873 5173 4887 5187 0 _1865_.B
rlabel metal2 4853 5153 4867 5167 0 _1865_.C
rlabel metal2 4833 5173 4847 5187 0 _1865_.Y
rlabel metal1 4904 5042 5016 5058 0 _1864_.gnd
rlabel metal1 4904 5282 5016 5298 0 _1864_.vdd
rlabel metal2 4913 5133 4927 5147 0 _1864_.A
rlabel metal2 4933 5153 4947 5167 0 _1864_.B
rlabel metal2 4973 5153 4987 5167 0 _1864_.C
rlabel metal2 4953 5133 4967 5147 0 _1864_.Y
rlabel metal1 5064 5042 5156 5058 0 _1810_.gnd
rlabel metal1 5064 5282 5156 5298 0 _1810_.vdd
rlabel metal2 5073 5173 5087 5187 0 _1810_.A
rlabel metal2 5113 5173 5127 5187 0 _1810_.B
rlabel metal2 5093 5153 5107 5167 0 _1810_.Y
rlabel metal1 5004 5042 5076 5058 0 _1680_.gnd
rlabel metal1 5004 5282 5076 5298 0 _1680_.vdd
rlabel metal2 5013 5153 5027 5167 0 _1680_.A
rlabel metal2 5033 5133 5047 5147 0 _1680_.Y
rlabel metal1 5304 5042 5416 5058 0 _1807_.gnd
rlabel metal1 5304 5282 5416 5298 0 _1807_.vdd
rlabel metal2 5313 5133 5327 5147 0 _1807_.A
rlabel metal2 5333 5153 5347 5167 0 _1807_.B
rlabel metal2 5373 5153 5387 5167 0 _1807_.C
rlabel metal2 5353 5133 5367 5147 0 _1807_.Y
rlabel metal1 5224 5042 5316 5058 0 _1811_.gnd
rlabel metal1 5224 5282 5316 5298 0 _1811_.vdd
rlabel metal2 5233 5173 5247 5187 0 _1811_.A
rlabel metal2 5273 5173 5287 5187 0 _1811_.B
rlabel metal2 5253 5153 5267 5167 0 _1811_.Y
rlabel metal1 5144 5042 5236 5058 0 _1668_.gnd
rlabel metal1 5144 5282 5236 5298 0 _1668_.vdd
rlabel metal2 5153 5153 5167 5167 0 _1668_.A
rlabel metal2 5193 5153 5207 5167 0 _1668_.Y
rlabel metal1 5604 5042 5676 5058 0 _1804_.gnd
rlabel metal1 5604 5282 5676 5298 0 _1804_.vdd
rlabel metal2 5613 5113 5627 5127 0 _1804_.A
rlabel metal2 5633 5153 5647 5167 0 _1804_.Y
rlabel metal1 5504 5042 5616 5058 0 _1812_.gnd
rlabel metal1 5504 5282 5616 5298 0 _1812_.vdd
rlabel metal2 5513 5153 5527 5167 0 _1812_.A
rlabel metal2 5533 5173 5547 5187 0 _1812_.B
rlabel metal2 5553 5153 5567 5167 0 _1812_.C
rlabel metal2 5573 5173 5587 5187 0 _1812_.Y
rlabel metal1 5404 5042 5516 5058 0 _1809_.gnd
rlabel metal1 5404 5282 5516 5298 0 _1809_.vdd
rlabel metal2 5413 5153 5427 5167 0 _1809_.A
rlabel metal2 5433 5173 5447 5187 0 _1809_.B
rlabel metal2 5453 5153 5467 5167 0 _1809_.C
rlabel metal2 5473 5173 5487 5187 0 _1809_.Y
rlabel metal1 5764 5042 5876 5058 0 _1899_.gnd
rlabel metal1 5764 5282 5876 5298 0 _1899_.vdd
rlabel metal2 5773 5133 5787 5147 0 _1899_.A
rlabel metal2 5793 5153 5807 5167 0 _1899_.B
rlabel metal2 5833 5153 5847 5167 0 _1899_.C
rlabel metal2 5813 5133 5827 5147 0 _1899_.Y
rlabel metal1 5864 5042 5956 5058 0 _1822_.gnd
rlabel metal1 5864 5282 5956 5298 0 _1822_.vdd
rlabel metal2 5933 5173 5947 5187 0 _1822_.A
rlabel metal2 5893 5173 5907 5187 0 _1822_.B
rlabel metal2 5913 5153 5927 5167 0 _1822_.Y
rlabel metal1 5664 5042 5776 5058 0 _1808_.gnd
rlabel metal1 5664 5282 5776 5298 0 _1808_.vdd
rlabel metal2 5673 5153 5687 5167 0 _1808_.A
rlabel metal2 5693 5173 5707 5187 0 _1808_.B
rlabel metal2 5713 5153 5727 5167 0 _1808_.C
rlabel metal2 5733 5173 5747 5187 0 _1808_.Y
rlabel metal1 6044 5042 6136 5058 0 _1776_.gnd
rlabel metal1 6044 5282 6136 5298 0 _1776_.vdd
rlabel metal2 6053 5173 6067 5187 0 _1776_.A
rlabel metal2 6093 5173 6107 5187 0 _1776_.B
rlabel metal2 6073 5153 6087 5167 0 _1776_.Y
rlabel metal1 6124 5042 6236 5058 0 _1855_.gnd
rlabel metal1 6124 5282 6236 5298 0 _1855_.vdd
rlabel metal2 6213 5153 6227 5167 0 _1855_.A
rlabel metal2 6193 5113 6207 5127 0 _1855_.B
rlabel metal2 6173 5153 6187 5167 0 _1855_.C
rlabel metal2 6153 5133 6167 5147 0 _1855_.Y
rlabel metal1 5944 5042 6056 5058 0 _1823_.gnd
rlabel metal1 5944 5282 6056 5298 0 _1823_.vdd
rlabel metal2 5953 5153 5967 5167 0 _1823_.A
rlabel metal2 5973 5173 5987 5187 0 _1823_.B
rlabel metal2 5993 5153 6007 5167 0 _1823_.C
rlabel metal2 6013 5173 6027 5187 0 _1823_.Y
rlabel metal1 6224 5042 6296 5058 0 _1854_.gnd
rlabel metal1 6224 5282 6296 5298 0 _1854_.vdd
rlabel metal2 6273 5113 6287 5127 0 _1854_.A
rlabel metal2 6253 5153 6267 5167 0 _1854_.Y
rlabel metal1 6384 5042 6496 5058 0 _1845_.gnd
rlabel metal1 6384 5282 6496 5298 0 _1845_.vdd
rlabel metal2 6473 5153 6487 5167 0 _1845_.A
rlabel metal2 6453 5173 6467 5187 0 _1845_.B
rlabel metal2 6433 5153 6447 5167 0 _1845_.C
rlabel metal2 6413 5173 6427 5187 0 _1845_.Y
rlabel metal1 6284 5042 6396 5058 0 _1838_.gnd
rlabel metal1 6284 5282 6396 5298 0 _1838_.vdd
rlabel metal2 6373 5153 6387 5167 0 _1838_.A
rlabel metal2 6353 5173 6367 5187 0 _1838_.B
rlabel metal2 6333 5153 6347 5167 0 _1838_.C
rlabel metal2 6313 5173 6327 5187 0 _1838_.Y
rlabel metal1 6484 5042 6556 5058 0 _1839_.gnd
rlabel metal1 6484 5282 6556 5298 0 _1839_.vdd
rlabel metal2 6493 5113 6507 5127 0 _1839_.A
rlabel metal2 6513 5153 6527 5167 0 _1839_.Y
rlabel metal1 6644 5042 6736 5058 0 _1837_.gnd
rlabel metal1 6644 5282 6736 5298 0 _1837_.vdd
rlabel metal2 6653 5173 6667 5187 0 _1837_.A
rlabel metal2 6693 5173 6707 5187 0 _1837_.B
rlabel metal2 6673 5153 6687 5167 0 _1837_.Y
rlabel metal1 6544 5042 6656 5058 0 _1841_.gnd
rlabel metal1 6544 5282 6656 5298 0 _1841_.vdd
rlabel metal2 6633 5153 6647 5167 0 _1841_.A
rlabel metal2 6613 5173 6627 5187 0 _1841_.B
rlabel metal2 6593 5153 6607 5167 0 _1841_.C
rlabel metal2 6573 5173 6587 5187 0 _1841_.Y
rlabel metal1 4 5522 256 5538 0 _1616_.gnd
rlabel metal1 4 5282 256 5298 0 _1616_.vdd
rlabel metal2 153 5433 167 5447 0 _1616_.D
rlabel metal2 113 5433 127 5447 0 _1616_.CLK
rlabel metal2 33 5433 47 5447 0 _1616_.Q
rlabel metal1 244 5522 336 5538 0 _1534_.gnd
rlabel metal1 244 5282 336 5298 0 _1534_.vdd
rlabel metal2 253 5393 267 5407 0 _1534_.A
rlabel metal2 293 5393 307 5407 0 _1534_.B
rlabel metal2 273 5413 287 5427 0 _1534_.Y
rlabel metal1 424 5522 516 5538 0 _1536_.gnd
rlabel metal1 424 5282 516 5298 0 _1536_.vdd
rlabel metal2 493 5393 507 5407 0 _1536_.A
rlabel metal2 453 5393 467 5407 0 _1536_.B
rlabel metal2 473 5413 487 5427 0 _1536_.Y
rlabel metal1 324 5522 436 5538 0 _1584_.gnd
rlabel metal1 324 5282 436 5298 0 _1584_.vdd
rlabel metal2 413 5413 427 5427 0 _1584_.A
rlabel metal2 393 5453 407 5467 0 _1584_.B
rlabel metal2 373 5413 387 5427 0 _1584_.C
rlabel metal2 353 5433 367 5447 0 _1584_.Y
rlabel metal1 504 5522 616 5538 0 _2301_.gnd
rlabel metal1 504 5282 616 5298 0 _2301_.vdd
rlabel metal2 593 5433 607 5447 0 _2301_.A
rlabel metal2 533 5433 547 5447 0 _2301_.Y
rlabel metal2 553 5393 567 5407 0 _2301_.B
rlabel metal1 684 5522 776 5538 0 _2315_.gnd
rlabel metal1 684 5282 776 5298 0 _2315_.vdd
rlabel metal2 733 5433 747 5447 0 _2315_.B
rlabel metal2 693 5433 707 5447 0 _2315_.A
rlabel metal2 713 5453 727 5467 0 _2315_.Y
rlabel metal1 604 5522 696 5538 0 _2302_.gnd
rlabel metal1 604 5282 696 5298 0 _2302_.vdd
rlabel metal2 653 5433 667 5447 0 _2302_.B
rlabel metal2 613 5433 627 5447 0 _2302_.A
rlabel metal2 633 5453 647 5467 0 _2302_.Y
rlabel metal1 764 5522 856 5538 0 _1535_.gnd
rlabel metal1 764 5282 856 5298 0 _1535_.vdd
rlabel metal2 773 5393 787 5407 0 _1535_.A
rlabel metal2 813 5393 827 5407 0 _1535_.B
rlabel metal2 793 5413 807 5427 0 _1535_.Y
rlabel metal1 924 5522 996 5538 0 _2299_.gnd
rlabel metal1 924 5282 996 5298 0 _2299_.vdd
rlabel metal2 933 5453 947 5467 0 _2299_.A
rlabel metal2 953 5413 967 5427 0 _2299_.Y
rlabel metal1 844 5522 936 5538 0 _1544_.gnd
rlabel metal1 844 5282 936 5298 0 _1544_.vdd
rlabel metal2 853 5393 867 5407 0 _1544_.A
rlabel metal2 893 5393 907 5407 0 _1544_.B
rlabel metal2 873 5413 887 5427 0 _1544_.Y
rlabel metal1 984 5522 1096 5538 0 _2306_.gnd
rlabel metal1 984 5282 1096 5298 0 _2306_.vdd
rlabel metal2 993 5413 1007 5427 0 _2306_.A
rlabel metal2 1013 5453 1027 5467 0 _2306_.B
rlabel metal2 1033 5413 1047 5427 0 _2306_.C
rlabel metal2 1053 5433 1067 5447 0 _2306_.Y
rlabel metal1 1204 5522 1456 5538 0 _2391_.gnd
rlabel metal1 1204 5282 1456 5298 0 _2391_.vdd
rlabel metal2 1353 5433 1367 5447 0 _2391_.D
rlabel metal2 1313 5433 1327 5447 0 _2391_.CLK
rlabel metal2 1233 5433 1247 5447 0 _2391_.Q
rlabel metal1 1084 5522 1216 5538 0 _2307_.gnd
rlabel metal1 1084 5282 1216 5298 0 _2307_.vdd
rlabel metal2 1193 5433 1207 5447 0 _2307_.A
rlabel metal2 1173 5413 1187 5427 0 _2307_.B
rlabel metal2 1113 5433 1127 5447 0 _2307_.C
rlabel metal2 1133 5413 1147 5427 0 _2307_.D
rlabel metal2 1153 5433 1167 5447 0 _2307_.Y
rlabel metal1 1444 5522 1556 5538 0 _2169_.gnd
rlabel metal1 1444 5282 1556 5298 0 _2169_.vdd
rlabel metal2 1533 5413 1547 5427 0 _2169_.A
rlabel metal2 1513 5393 1527 5407 0 _2169_.B
rlabel metal2 1493 5413 1507 5427 0 _2169_.C
rlabel metal2 1473 5393 1487 5407 0 _2169_.Y
rlabel metal1 1544 5522 1656 5538 0 _2162_.gnd
rlabel metal1 1544 5282 1656 5298 0 _2162_.vdd
rlabel metal2 1633 5413 1647 5427 0 _2162_.A
rlabel metal2 1613 5393 1627 5407 0 _2162_.B
rlabel metal2 1593 5413 1607 5427 0 _2162_.C
rlabel metal2 1573 5393 1587 5407 0 _2162_.Y
rlabel metal1 1704 5522 1816 5538 0 _2168_.gnd
rlabel metal1 1704 5282 1816 5298 0 _2168_.vdd
rlabel metal2 1793 5433 1807 5447 0 _2168_.A
rlabel metal2 1773 5413 1787 5427 0 _2168_.B
rlabel metal2 1733 5413 1747 5427 0 _2168_.C
rlabel metal2 1753 5433 1767 5447 0 _2168_.Y
rlabel metal1 1644 5522 1716 5538 0 _2167_.gnd
rlabel metal1 1644 5282 1716 5298 0 _2167_.vdd
rlabel metal2 1693 5453 1707 5467 0 _2167_.A
rlabel metal2 1673 5413 1687 5427 0 _2167_.Y
rlabel metal1 1804 5522 1916 5538 0 _2152_.gnd
rlabel metal1 1804 5282 1916 5298 0 _2152_.vdd
rlabel metal2 1893 5433 1907 5447 0 _2152_.A
rlabel metal2 1833 5433 1847 5447 0 _2152_.Y
rlabel metal2 1853 5393 1867 5407 0 _2152_.B
rlabel metal1 1984 5522 2096 5538 0 _2151_.gnd
rlabel metal1 1984 5282 2096 5298 0 _2151_.vdd
rlabel metal2 2073 5433 2087 5447 0 _2151_.A
rlabel metal2 2053 5413 2067 5427 0 _2151_.B
rlabel metal2 2013 5413 2027 5427 0 _2151_.C
rlabel metal2 2033 5433 2047 5447 0 _2151_.Y
rlabel metal1 1904 5522 1996 5538 0 _2139_.gnd
rlabel metal1 1904 5282 1996 5298 0 _2139_.vdd
rlabel metal2 1973 5393 1987 5407 0 _2139_.A
rlabel metal2 1933 5393 1947 5407 0 _2139_.B
rlabel metal2 1953 5413 1967 5427 0 _2139_.Y
rlabel metal1 2084 5522 2176 5538 0 _2138_.gnd
rlabel metal1 2084 5282 2176 5298 0 _2138_.vdd
rlabel metal2 2093 5393 2107 5407 0 _2138_.A
rlabel metal2 2133 5393 2147 5407 0 _2138_.B
rlabel metal2 2113 5413 2127 5427 0 _2138_.Y
rlabel metal1 2224 5522 2336 5538 0 _2135_.gnd
rlabel metal1 2224 5282 2336 5298 0 _2135_.vdd
rlabel metal2 2313 5433 2327 5447 0 _2135_.A
rlabel metal2 2293 5413 2307 5427 0 _2135_.B
rlabel metal2 2253 5413 2267 5427 0 _2135_.C
rlabel metal2 2273 5433 2287 5447 0 _2135_.Y
rlabel metal1 2324 5522 2416 5538 0 _2137_.gnd
rlabel metal1 2324 5282 2416 5298 0 _2137_.vdd
rlabel metal2 2373 5433 2387 5447 0 _2137_.B
rlabel metal2 2333 5433 2347 5447 0 _2137_.A
rlabel metal2 2353 5453 2367 5467 0 _2137_.Y
rlabel metal1 2164 5522 2236 5538 0 _2136_.gnd
rlabel metal1 2164 5282 2236 5298 0 _2136_.vdd
rlabel metal2 2213 5453 2227 5467 0 _2136_.A
rlabel metal2 2193 5413 2207 5427 0 _2136_.Y
rlabel metal1 2404 5522 2476 5538 0 _1984_.gnd
rlabel metal1 2404 5282 2476 5298 0 _1984_.vdd
rlabel metal2 2453 5453 2467 5467 0 _1984_.A
rlabel metal2 2433 5413 2447 5427 0 _1984_.Y
rlabel metal1 2564 5522 2676 5538 0 _1978_.gnd
rlabel metal1 2564 5282 2676 5298 0 _1978_.vdd
rlabel metal2 2573 5433 2587 5447 0 _1978_.A
rlabel metal2 2593 5413 2607 5427 0 _1978_.B
rlabel metal2 2633 5413 2647 5427 0 _1978_.C
rlabel metal2 2613 5433 2627 5447 0 _1978_.Y
rlabel metal1 2664 5522 2756 5538 0 _2110_.gnd
rlabel metal1 2664 5282 2756 5298 0 _2110_.vdd
rlabel metal2 2673 5393 2687 5407 0 _2110_.A
rlabel metal2 2713 5393 2727 5407 0 _2110_.B
rlabel metal2 2693 5413 2707 5427 0 _2110_.Y
rlabel metal1 2464 5522 2576 5538 0 _1979_.gnd
rlabel metal1 2464 5282 2576 5298 0 _1979_.vdd
rlabel metal2 2553 5413 2567 5427 0 _1979_.A
rlabel metal2 2533 5453 2547 5467 0 _1979_.B
rlabel metal2 2513 5413 2527 5427 0 _1979_.C
rlabel metal2 2493 5433 2507 5447 0 _1979_.Y
rlabel metal1 2924 5522 3016 5538 0 _2107_.gnd
rlabel metal1 2924 5282 3016 5298 0 _2107_.vdd
rlabel metal2 2953 5433 2967 5447 0 _2107_.B
rlabel metal2 2993 5433 3007 5447 0 _2107_.A
rlabel metal2 2973 5453 2987 5467 0 _2107_.Y
rlabel metal1 2844 5522 2936 5538 0 _2109_.gnd
rlabel metal1 2844 5282 2936 5298 0 _2109_.vdd
rlabel metal2 2913 5393 2927 5407 0 _2109_.A
rlabel metal2 2873 5393 2887 5407 0 _2109_.B
rlabel metal2 2893 5413 2907 5427 0 _2109_.Y
rlabel metal1 2744 5522 2856 5538 0 _2113_.gnd
rlabel metal1 2744 5282 2856 5298 0 _2113_.vdd
rlabel metal2 2833 5413 2847 5427 0 _2113_.A
rlabel metal2 2813 5393 2827 5407 0 _2113_.B
rlabel metal2 2793 5413 2807 5427 0 _2113_.C
rlabel metal2 2773 5393 2787 5407 0 _2113_.Y
rlabel metal1 3004 5522 3116 5538 0 _2106_.gnd
rlabel metal1 3004 5282 3116 5298 0 _2106_.vdd
rlabel metal2 3013 5433 3027 5447 0 _2106_.A
rlabel metal2 3033 5413 3047 5427 0 _2106_.B
rlabel metal2 3073 5413 3087 5427 0 _2106_.C
rlabel metal2 3053 5433 3067 5447 0 _2106_.Y
rlabel metal1 3184 5522 3296 5538 0 _2061_.gnd
rlabel metal1 3184 5282 3296 5298 0 _2061_.vdd
rlabel metal2 3193 5433 3207 5447 0 _2061_.A
rlabel metal2 3213 5413 3227 5427 0 _2061_.B
rlabel metal2 3253 5413 3267 5427 0 _2061_.C
rlabel metal2 3233 5433 3247 5447 0 _2061_.Y
rlabel metal1 3104 5522 3196 5538 0 _2044_.gnd
rlabel metal1 3104 5282 3196 5298 0 _2044_.vdd
rlabel metal2 3173 5393 3187 5407 0 _2044_.A
rlabel metal2 3133 5393 3147 5407 0 _2044_.B
rlabel metal2 3153 5413 3167 5427 0 _2044_.Y
rlabel metal1 3384 5522 3476 5538 0 _2057_.gnd
rlabel metal1 3384 5282 3476 5298 0 _2057_.vdd
rlabel metal2 3433 5433 3447 5447 0 _2057_.B
rlabel metal2 3393 5433 3407 5447 0 _2057_.A
rlabel metal2 3413 5453 3427 5467 0 _2057_.Y
rlabel metal1 3464 5522 3576 5538 0 _2054_.gnd
rlabel metal1 3464 5282 3576 5298 0 _2054_.vdd
rlabel metal2 3473 5453 3487 5467 0 _2054_.A
rlabel metal2 3493 5433 3507 5447 0 _2054_.B
rlabel metal2 3533 5413 3547 5427 0 _2054_.Y
rlabel metal1 3284 5522 3396 5538 0 _2058_.gnd
rlabel metal1 3284 5282 3396 5298 0 _2058_.vdd
rlabel metal2 3373 5433 3387 5447 0 _2058_.A
rlabel metal2 3313 5433 3327 5447 0 _2058_.Y
rlabel metal2 3333 5393 3347 5407 0 _2058_.B
rlabel metal1 3564 5522 3676 5538 0 _2055_.gnd
rlabel metal1 3564 5282 3676 5298 0 _2055_.vdd
rlabel metal2 3573 5433 3587 5447 0 _2055_.A
rlabel metal2 3593 5413 3607 5427 0 _2055_.B
rlabel metal2 3633 5413 3647 5427 0 _2055_.C
rlabel metal2 3613 5433 3627 5447 0 _2055_.Y
rlabel metal1 3664 5522 3756 5538 0 _1993_.gnd
rlabel metal1 3664 5282 3756 5298 0 _1993_.vdd
rlabel metal2 3693 5433 3707 5447 0 _1993_.B
rlabel metal2 3733 5433 3747 5447 0 _1993_.A
rlabel metal2 3713 5453 3727 5467 0 _1993_.Y
rlabel metal1 3744 5522 3876 5538 0 _1992_.gnd
rlabel metal1 3744 5282 3876 5298 0 _1992_.vdd
rlabel metal2 3753 5433 3767 5447 0 _1992_.A
rlabel metal2 3773 5413 3787 5427 0 _1992_.B
rlabel metal2 3833 5433 3847 5447 0 _1992_.C
rlabel metal2 3793 5433 3807 5447 0 _1992_.Y
rlabel metal2 3813 5413 3827 5427 0 _1992_.D
rlabel metal1 3944 5522 4056 5538 0 _1935_.gnd
rlabel metal1 3944 5282 4056 5298 0 _1935_.vdd
rlabel metal2 3953 5433 3967 5447 0 _1935_.A
rlabel metal2 3973 5413 3987 5427 0 _1935_.B
rlabel metal2 4013 5413 4027 5427 0 _1935_.C
rlabel metal2 3993 5433 4007 5447 0 _1935_.Y
rlabel metal1 3864 5522 3956 5538 0 _2095_.gnd
rlabel metal1 3864 5282 3956 5298 0 _2095_.vdd
rlabel metal2 3893 5433 3907 5447 0 _2095_.B
rlabel metal2 3933 5433 3947 5447 0 _2095_.A
rlabel metal2 3913 5453 3927 5467 0 _2095_.Y
rlabel metal1 4224 5522 4296 5538 0 _1922_.gnd
rlabel metal1 4224 5282 4296 5298 0 _1922_.vdd
rlabel metal2 4233 5453 4247 5467 0 _1922_.A
rlabel metal2 4253 5413 4267 5427 0 _1922_.Y
rlabel metal1 4144 5522 4236 5538 0 _1930_.gnd
rlabel metal1 4144 5282 4236 5298 0 _1930_.vdd
rlabel metal2 4213 5393 4227 5407 0 _1930_.A
rlabel metal2 4173 5393 4187 5407 0 _1930_.B
rlabel metal2 4193 5413 4207 5427 0 _1930_.Y
rlabel metal1 4044 5522 4156 5538 0 _1936_.gnd
rlabel metal1 4044 5282 4156 5298 0 _1936_.vdd
rlabel metal2 4133 5413 4147 5427 0 _1936_.A
rlabel metal2 4113 5393 4127 5407 0 _1936_.B
rlabel metal2 4093 5413 4107 5427 0 _1936_.C
rlabel metal2 4073 5393 4087 5407 0 _1936_.Y
rlabel metal1 4284 5522 4396 5538 0 _1932_.gnd
rlabel metal1 4284 5282 4396 5298 0 _1932_.vdd
rlabel metal2 4373 5433 4387 5447 0 _1932_.A
rlabel metal2 4353 5413 4367 5427 0 _1932_.B
rlabel metal2 4313 5413 4327 5427 0 _1932_.C
rlabel metal2 4333 5433 4347 5447 0 _1932_.Y
rlabel metal1 4384 5522 4476 5538 0 _2000_.gnd
rlabel metal1 4384 5282 4476 5298 0 _2000_.vdd
rlabel metal2 4453 5393 4467 5407 0 _2000_.A
rlabel metal2 4413 5393 4427 5407 0 _2000_.B
rlabel metal2 4433 5413 4447 5427 0 _2000_.Y
rlabel metal1 4464 5522 4556 5538 0 _1941_.gnd
rlabel metal1 4464 5282 4556 5298 0 _1941_.vdd
rlabel metal2 4473 5393 4487 5407 0 _1941_.A
rlabel metal2 4513 5393 4527 5407 0 _1941_.B
rlabel metal2 4493 5413 4507 5427 0 _1941_.Y
rlabel metal1 4544 5522 4656 5538 0 _2002_.gnd
rlabel metal1 4544 5282 4656 5298 0 _2002_.vdd
rlabel metal2 4633 5433 4647 5447 0 _2002_.A
rlabel metal2 4613 5413 4627 5427 0 _2002_.B
rlabel metal2 4573 5413 4587 5427 0 _2002_.C
rlabel metal2 4593 5433 4607 5447 0 _2002_.Y
rlabel metal1 4644 5522 4756 5538 0 _1923_.gnd
rlabel metal1 4644 5282 4756 5298 0 _1923_.vdd
rlabel metal2 4733 5433 4747 5447 0 _1923_.A
rlabel metal2 4713 5413 4727 5427 0 _1923_.B
rlabel metal2 4673 5413 4687 5427 0 _1923_.C
rlabel metal2 4693 5433 4707 5447 0 _1923_.Y
rlabel metal1 4744 5522 4856 5538 0 _1878_.gnd
rlabel metal1 4744 5282 4856 5298 0 _1878_.vdd
rlabel metal2 4833 5433 4847 5447 0 _1878_.A
rlabel metal2 4773 5433 4787 5447 0 _1878_.Y
rlabel metal2 4793 5393 4807 5407 0 _1878_.B
rlabel metal1 4844 5522 4956 5538 0 _1944_.gnd
rlabel metal1 4844 5282 4956 5298 0 _1944_.vdd
rlabel metal2 4933 5433 4947 5447 0 _1944_.A
rlabel metal2 4913 5413 4927 5427 0 _1944_.B
rlabel metal2 4873 5413 4887 5427 0 _1944_.C
rlabel metal2 4893 5433 4907 5447 0 _1944_.Y
rlabel metal1 4944 5522 5036 5538 0 _1938_.gnd
rlabel metal1 4944 5282 5036 5298 0 _1938_.vdd
rlabel metal2 5013 5393 5027 5407 0 _1938_.A
rlabel metal2 4973 5393 4987 5407 0 _1938_.B
rlabel metal2 4993 5413 5007 5427 0 _1938_.Y
rlabel metal1 5024 5522 5136 5538 0 _1939_.gnd
rlabel metal1 5024 5282 5136 5298 0 _1939_.vdd
rlabel metal2 5113 5433 5127 5447 0 _1939_.A
rlabel metal2 5053 5433 5067 5447 0 _1939_.Y
rlabel metal2 5073 5393 5087 5407 0 _1939_.B
rlabel metal1 5204 5522 5316 5538 0 _1875_.gnd
rlabel metal1 5204 5282 5316 5298 0 _1875_.vdd
rlabel metal2 5213 5433 5227 5447 0 _1875_.A
rlabel metal2 5233 5413 5247 5427 0 _1875_.B
rlabel metal2 5273 5413 5287 5427 0 _1875_.C
rlabel metal2 5253 5433 5267 5447 0 _1875_.Y
rlabel metal1 5124 5522 5216 5538 0 _1873_.gnd
rlabel metal1 5124 5282 5216 5298 0 _1873_.vdd
rlabel metal2 5133 5393 5147 5407 0 _1873_.A
rlabel metal2 5173 5393 5187 5407 0 _1873_.B
rlabel metal2 5153 5413 5167 5427 0 _1873_.Y
rlabel metal1 5304 5522 5416 5538 0 _1817_.gnd
rlabel metal1 5304 5282 5416 5298 0 _1817_.vdd
rlabel metal2 5393 5433 5407 5447 0 _1817_.A
rlabel metal2 5333 5433 5347 5447 0 _1817_.Y
rlabel metal2 5353 5393 5367 5407 0 _1817_.B
rlabel metal1 5404 5522 5516 5538 0 _1820_.gnd
rlabel metal1 5404 5282 5516 5298 0 _1820_.vdd
rlabel metal2 5413 5433 5427 5447 0 _1820_.A
rlabel metal2 5433 5413 5447 5427 0 _1820_.B
rlabel metal2 5473 5413 5487 5427 0 _1820_.C
rlabel metal2 5453 5433 5467 5447 0 _1820_.Y
rlabel metal1 5504 5522 5596 5538 0 _1819_.gnd
rlabel metal1 5504 5282 5596 5298 0 _1819_.vdd
rlabel metal2 5513 5393 5527 5407 0 _1819_.A
rlabel metal2 5553 5393 5567 5407 0 _1819_.B
rlabel metal2 5533 5413 5547 5427 0 _1819_.Y
rlabel metal1 5584 5522 5696 5538 0 _1824_.gnd
rlabel metal1 5584 5282 5696 5298 0 _1824_.vdd
rlabel metal2 5593 5413 5607 5427 0 _1824_.A
rlabel metal2 5613 5393 5627 5407 0 _1824_.B
rlabel metal2 5633 5413 5647 5427 0 _1824_.C
rlabel metal2 5653 5393 5667 5407 0 _1824_.Y
rlabel metal1 5784 5522 5916 5538 0 _1870_.gnd
rlabel metal1 5784 5282 5916 5298 0 _1870_.vdd
rlabel metal2 5893 5433 5907 5447 0 _1870_.A
rlabel metal2 5873 5413 5887 5427 0 _1870_.B
rlabel metal2 5813 5433 5827 5447 0 _1870_.C
rlabel metal2 5833 5413 5847 5427 0 _1870_.D
rlabel metal2 5853 5433 5867 5447 0 _1870_.Y
rlabel metal1 5684 5522 5796 5538 0 _1816_.gnd
rlabel metal1 5684 5282 5796 5298 0 _1816_.vdd
rlabel metal2 5773 5433 5787 5447 0 _1816_.A
rlabel metal2 5713 5433 5727 5447 0 _1816_.Y
rlabel metal2 5733 5393 5747 5407 0 _1816_.B
rlabel metal1 5904 5522 5996 5538 0 _1814_.gnd
rlabel metal1 5904 5282 5996 5298 0 _1814_.vdd
rlabel metal2 5913 5393 5927 5407 0 _1814_.A
rlabel metal2 5953 5393 5967 5407 0 _1814_.B
rlabel metal2 5933 5413 5947 5427 0 _1814_.Y
rlabel metal1 6084 5522 6196 5538 0 _1827_.gnd
rlabel metal1 6084 5282 6196 5298 0 _1827_.vdd
rlabel metal2 6093 5413 6107 5427 0 _1827_.A
rlabel metal2 6113 5453 6127 5467 0 _1827_.B
rlabel metal2 6133 5413 6147 5427 0 _1827_.C
rlabel metal2 6153 5433 6167 5447 0 _1827_.Y
rlabel metal1 5984 5522 6096 5538 0 _1825_.gnd
rlabel metal1 5984 5282 6096 5298 0 _1825_.vdd
rlabel metal2 5993 5413 6007 5427 0 _1825_.A
rlabel metal2 6013 5393 6027 5407 0 _1825_.B
rlabel metal2 6033 5413 6047 5427 0 _1825_.C
rlabel metal2 6053 5393 6067 5407 0 _1825_.Y
rlabel metal1 6384 5522 6496 5538 0 _1905_.gnd
rlabel metal1 6384 5282 6496 5298 0 _1905_.vdd
rlabel metal2 6473 5433 6487 5447 0 _1905_.A
rlabel metal2 6453 5413 6467 5427 0 _1905_.B
rlabel metal2 6413 5413 6427 5427 0 _1905_.C
rlabel metal2 6433 5433 6447 5447 0 _1905_.Y
rlabel metal1 6284 5522 6396 5538 0 _1832_.gnd
rlabel metal1 6284 5282 6396 5298 0 _1832_.vdd
rlabel metal2 6293 5433 6307 5447 0 _1832_.A
rlabel metal2 6313 5413 6327 5427 0 _1832_.B
rlabel metal2 6353 5413 6367 5427 0 _1832_.C
rlabel metal2 6333 5433 6347 5447 0 _1832_.Y
rlabel metal1 6184 5522 6296 5538 0 _1829_.gnd
rlabel metal1 6184 5282 6296 5298 0 _1829_.vdd
rlabel metal2 6273 5433 6287 5447 0 _1829_.A
rlabel metal2 6253 5413 6267 5427 0 _1829_.B
rlabel metal2 6213 5413 6227 5427 0 _1829_.C
rlabel metal2 6233 5433 6247 5447 0 _1829_.Y
rlabel metal1 6584 5522 6696 5538 0 _1904_.gnd
rlabel metal1 6584 5282 6696 5298 0 _1904_.vdd
rlabel metal2 6673 5413 6687 5427 0 _1904_.A
rlabel metal2 6653 5453 6667 5467 0 _1904_.B
rlabel metal2 6633 5413 6647 5427 0 _1904_.C
rlabel metal2 6613 5433 6627 5447 0 _1904_.Y
rlabel metal1 6484 5522 6596 5538 0 _1835_.gnd
rlabel metal1 6484 5282 6596 5298 0 _1835_.vdd
rlabel metal2 6573 5413 6587 5427 0 _1835_.A
rlabel metal2 6553 5393 6567 5407 0 _1835_.B
rlabel metal2 6533 5413 6547 5427 0 _1835_.C
rlabel metal2 6513 5393 6527 5407 0 _1835_.Y
rlabel nsubstratencontact 6724 5292 6724 5292 0 FILL100650x79350.vdd
rlabel metal1 6704 5522 6736 5538 0 FILL100650x79350.gnd
rlabel nsubstratencontact 6704 5292 6704 5292 0 FILL100350x79350.vdd
rlabel metal1 6684 5522 6716 5538 0 FILL100350x79350.gnd
rlabel metal1 4 5522 96 5538 0 _3045_.gnd
rlabel metal1 4 5762 96 5778 0 _3045_.vdd
rlabel metal2 73 5613 87 5627 0 _3045_.A
rlabel metal2 33 5613 47 5627 0 _3045_.Y
rlabel metal1 84 5522 176 5538 0 _3033_.gnd
rlabel metal1 84 5762 176 5778 0 _3033_.vdd
rlabel metal2 153 5613 167 5627 0 _3033_.A
rlabel metal2 113 5613 127 5627 0 _3033_.Y
rlabel metal1 164 5522 416 5538 0 _1618_.gnd
rlabel metal1 164 5762 416 5778 0 _1618_.vdd
rlabel metal2 313 5613 327 5627 0 _1618_.D
rlabel metal2 273 5613 287 5627 0 _1618_.CLK
rlabel metal2 193 5613 207 5627 0 _1618_.Q
rlabel metal1 404 5522 496 5538 0 _2303_.gnd
rlabel metal1 404 5762 496 5778 0 _2303_.vdd
rlabel metal2 433 5613 447 5627 0 _2303_.B
rlabel metal2 473 5613 487 5627 0 _2303_.A
rlabel metal2 453 5593 467 5607 0 _2303_.Y
rlabel metal1 484 5522 596 5538 0 _2309_.gnd
rlabel metal1 484 5762 596 5778 0 _2309_.vdd
rlabel metal2 493 5633 507 5647 0 _2309_.A
rlabel metal2 513 5593 527 5607 0 _2309_.B
rlabel metal2 533 5633 547 5647 0 _2309_.C
rlabel metal2 553 5613 567 5627 0 _2309_.Y
rlabel metal1 584 5522 676 5538 0 _2312_.gnd
rlabel metal1 584 5762 676 5778 0 _2312_.vdd
rlabel metal2 593 5653 607 5667 0 _2312_.A
rlabel metal2 633 5653 647 5667 0 _2312_.B
rlabel metal2 613 5633 627 5647 0 _2312_.Y
rlabel metal1 764 5522 856 5538 0 _2311_.gnd
rlabel metal1 764 5762 856 5778 0 _2311_.vdd
rlabel metal2 773 5653 787 5667 0 _2311_.A
rlabel metal2 813 5653 827 5667 0 _2311_.B
rlabel metal2 793 5633 807 5647 0 _2311_.Y
rlabel metal1 664 5522 776 5538 0 _2310_.gnd
rlabel metal1 664 5762 776 5778 0 _2310_.vdd
rlabel metal2 673 5613 687 5627 0 _2310_.A
rlabel metal2 733 5613 747 5627 0 _2310_.Y
rlabel metal2 713 5653 727 5667 0 _2310_.B
rlabel metal1 924 5522 1016 5538 0 _2314_.gnd
rlabel metal1 924 5762 1016 5778 0 _2314_.vdd
rlabel metal2 973 5613 987 5627 0 _2314_.B
rlabel metal2 933 5613 947 5627 0 _2314_.A
rlabel metal2 953 5593 967 5607 0 _2314_.Y
rlabel metal1 1004 5522 1076 5538 0 _2304_.gnd
rlabel metal1 1004 5762 1076 5778 0 _2304_.vdd
rlabel metal2 1013 5593 1027 5607 0 _2304_.A
rlabel metal2 1033 5633 1047 5647 0 _2304_.Y
rlabel metal1 844 5522 936 5538 0 _2313_.gnd
rlabel metal1 844 5762 936 5778 0 _2313_.vdd
rlabel metal2 853 5653 867 5667 0 _2313_.A
rlabel metal2 893 5653 907 5667 0 _2313_.B
rlabel metal2 873 5633 887 5647 0 _2313_.Y
rlabel metal1 1064 5522 1176 5538 0 _2305_.gnd
rlabel metal1 1064 5762 1176 5778 0 _2305_.vdd
rlabel metal2 1073 5593 1087 5607 0 _2305_.A
rlabel metal2 1093 5613 1107 5627 0 _2305_.B
rlabel metal2 1133 5633 1147 5647 0 _2305_.Y
rlabel metal1 1164 5522 1256 5538 0 _2261_.gnd
rlabel metal1 1164 5762 1256 5778 0 _2261_.vdd
rlabel metal2 1213 5613 1227 5627 0 _2261_.B
rlabel metal2 1173 5613 1187 5627 0 _2261_.A
rlabel metal2 1193 5593 1207 5607 0 _2261_.Y
rlabel metal1 1304 5522 1396 5538 0 _2260_.gnd
rlabel metal1 1304 5762 1396 5778 0 _2260_.vdd
rlabel metal2 1353 5613 1367 5627 0 _2260_.B
rlabel metal2 1313 5613 1327 5627 0 _2260_.A
rlabel metal2 1333 5593 1347 5607 0 _2260_.Y
rlabel metal1 1244 5522 1316 5538 0 _2259_.gnd
rlabel metal1 1244 5762 1316 5778 0 _2259_.vdd
rlabel metal2 1253 5593 1267 5607 0 _2259_.A
rlabel metal2 1273 5633 1287 5647 0 _2259_.Y
rlabel metal1 1444 5522 1696 5538 0 _2374_.gnd
rlabel metal1 1444 5762 1696 5778 0 _2374_.vdd
rlabel metal2 1593 5613 1607 5627 0 _2374_.D
rlabel metal2 1553 5613 1567 5627 0 _2374_.CLK
rlabel metal2 1473 5613 1487 5627 0 _2374_.Q
rlabel metal1 1384 5522 1456 5538 0 _1981_.gnd
rlabel metal1 1384 5762 1456 5778 0 _1981_.vdd
rlabel metal2 1393 5593 1407 5607 0 _1981_.A
rlabel metal2 1413 5633 1427 5647 0 _1981_.Y
rlabel metal1 1684 5522 1816 5538 0 _2042_.gnd
rlabel metal1 1684 5762 1816 5778 0 _2042_.vdd
rlabel metal2 1693 5613 1707 5627 0 _2042_.A
rlabel metal2 1713 5633 1727 5647 0 _2042_.B
rlabel metal2 1773 5613 1787 5627 0 _2042_.C
rlabel metal2 1733 5613 1747 5627 0 _2042_.Y
rlabel metal2 1753 5633 1767 5647 0 _2042_.D
rlabel metal1 1804 5522 1916 5538 0 _2164_.gnd
rlabel metal1 1804 5762 1916 5778 0 _2164_.vdd
rlabel metal2 1893 5613 1907 5627 0 _2164_.A
rlabel metal2 1873 5633 1887 5647 0 _2164_.B
rlabel metal2 1833 5633 1847 5647 0 _2164_.C
rlabel metal2 1853 5613 1867 5627 0 _2164_.Y
rlabel metal1 1984 5522 2056 5538 0 _2146_.gnd
rlabel metal1 1984 5762 2056 5778 0 _2146_.vdd
rlabel metal2 1993 5593 2007 5607 0 _2146_.A
rlabel metal2 2013 5633 2027 5647 0 _2146_.Y
rlabel metal1 1904 5522 1996 5538 0 _2163_.gnd
rlabel metal1 1904 5762 1996 5778 0 _2163_.vdd
rlabel metal2 1973 5653 1987 5667 0 _2163_.A
rlabel metal2 1933 5653 1947 5667 0 _2163_.B
rlabel metal2 1953 5633 1967 5647 0 _2163_.Y
rlabel metal1 2044 5522 2156 5538 0 _2166_.gnd
rlabel metal1 2044 5762 2156 5778 0 _2166_.vdd
rlabel metal2 2133 5633 2147 5647 0 _2166_.A
rlabel metal2 2113 5593 2127 5607 0 _2166_.B
rlabel metal2 2093 5633 2107 5647 0 _2166_.C
rlabel metal2 2073 5613 2087 5627 0 _2166_.Y
rlabel metal1 2144 5522 2236 5538 0 _2037_.gnd
rlabel metal1 2144 5762 2236 5778 0 _2037_.vdd
rlabel metal2 2193 5613 2207 5627 0 _2037_.B
rlabel metal2 2153 5613 2167 5627 0 _2037_.A
rlabel metal2 2173 5593 2187 5607 0 _2037_.Y
rlabel metal1 2224 5522 2316 5538 0 _1986_.gnd
rlabel metal1 2224 5762 2316 5778 0 _1986_.vdd
rlabel metal2 2233 5653 2247 5667 0 _1986_.A
rlabel metal2 2273 5653 2287 5667 0 _1986_.B
rlabel metal2 2253 5633 2267 5647 0 _1986_.Y
rlabel metal1 2304 5762 2496 5778 0 _2039_.vdd
rlabel metal2 2453 5613 2467 5627 0 _2039_.A
rlabel metal2 2413 5633 2427 5647 0 _2039_.B
rlabel metal2 2393 5613 2407 5627 0 _2039_.C
rlabel metal2 2353 5633 2367 5647 0 _2039_.Y
rlabel metal1 2304 5522 2496 5538 0 _2039_.gnd
rlabel metal1 2484 5522 2576 5538 0 _2114_.gnd
rlabel metal1 2484 5762 2576 5778 0 _2114_.vdd
rlabel metal2 2553 5653 2567 5667 0 _2114_.A
rlabel metal2 2513 5653 2527 5667 0 _2114_.B
rlabel metal2 2533 5633 2547 5647 0 _2114_.Y
rlabel metal1 2564 5522 2676 5538 0 _2117_.gnd
rlabel metal1 2564 5762 2676 5778 0 _2117_.vdd
rlabel metal2 2653 5633 2667 5647 0 _2117_.A
rlabel metal2 2633 5653 2647 5667 0 _2117_.B
rlabel metal2 2613 5633 2627 5647 0 _2117_.C
rlabel metal2 2593 5653 2607 5667 0 _2117_.Y
rlabel metal1 2664 5522 2776 5538 0 _2111_.gnd
rlabel metal1 2664 5762 2776 5778 0 _2111_.vdd
rlabel metal2 2753 5633 2767 5647 0 _2111_.A
rlabel metal2 2733 5653 2747 5667 0 _2111_.B
rlabel metal2 2713 5633 2727 5647 0 _2111_.C
rlabel metal2 2693 5653 2707 5667 0 _2111_.Y
rlabel metal1 2844 5522 2956 5538 0 _1918_.gnd
rlabel metal1 2844 5762 2956 5778 0 _1918_.vdd
rlabel metal2 2853 5613 2867 5627 0 _1918_.A
rlabel metal2 2873 5633 2887 5647 0 _1918_.B
rlabel metal2 2913 5633 2927 5647 0 _1918_.C
rlabel metal2 2893 5613 2907 5627 0 _1918_.Y
rlabel metal1 2764 5522 2856 5538 0 _2112_.gnd
rlabel metal1 2764 5762 2856 5778 0 _2112_.vdd
rlabel metal2 2773 5653 2787 5667 0 _2112_.A
rlabel metal2 2813 5653 2827 5667 0 _2112_.B
rlabel metal2 2793 5633 2807 5647 0 _2112_.Y
rlabel metal1 3144 5522 3256 5538 0 _2059_.gnd
rlabel metal1 3144 5762 3256 5778 0 _2059_.vdd
rlabel metal2 3233 5613 3247 5627 0 _2059_.A
rlabel metal2 3213 5633 3227 5647 0 _2059_.B
rlabel metal2 3173 5633 3187 5647 0 _2059_.C
rlabel metal2 3193 5613 3207 5627 0 _2059_.Y
rlabel metal1 3044 5522 3156 5538 0 _2068_.gnd
rlabel metal1 3044 5762 3156 5778 0 _2068_.vdd
rlabel metal2 3053 5633 3067 5647 0 _2068_.A
rlabel metal2 3073 5593 3087 5607 0 _2068_.B
rlabel metal2 3093 5633 3107 5647 0 _2068_.C
rlabel metal2 3113 5613 3127 5627 0 _2068_.Y
rlabel metal1 2944 5522 3056 5538 0 _2060_.gnd
rlabel metal1 2944 5762 3056 5778 0 _2060_.vdd
rlabel metal2 3033 5633 3047 5647 0 _2060_.A
rlabel metal2 3013 5653 3027 5667 0 _2060_.B
rlabel metal2 2993 5633 3007 5647 0 _2060_.C
rlabel metal2 2973 5653 2987 5667 0 _2060_.Y
rlabel metal1 3244 5522 3316 5538 0 _2048_.gnd
rlabel metal1 3244 5762 3316 5778 0 _2048_.vdd
rlabel metal2 3293 5593 3307 5607 0 _2048_.A
rlabel metal2 3273 5633 3287 5647 0 _2048_.Y
rlabel metal1 3404 5522 3516 5538 0 _2063_.gnd
rlabel metal1 3404 5762 3516 5778 0 _2063_.vdd
rlabel metal2 3493 5633 3507 5647 0 _2063_.A
rlabel metal2 3473 5653 3487 5667 0 _2063_.B
rlabel metal2 3453 5633 3467 5647 0 _2063_.C
rlabel metal2 3433 5653 3447 5667 0 _2063_.Y
rlabel metal1 3304 5522 3416 5538 0 _2056_.gnd
rlabel metal1 3304 5762 3416 5778 0 _2056_.vdd
rlabel metal2 3313 5633 3327 5647 0 _2056_.A
rlabel metal2 3333 5653 3347 5667 0 _2056_.B
rlabel metal2 3353 5633 3367 5647 0 _2056_.C
rlabel metal2 3373 5653 3387 5667 0 _2056_.Y
rlabel metal1 3664 5522 3776 5538 0 _1995_.gnd
rlabel metal1 3664 5762 3776 5778 0 _1995_.vdd
rlabel metal2 3753 5613 3767 5627 0 _1995_.A
rlabel metal2 3733 5633 3747 5647 0 _1995_.B
rlabel metal2 3693 5633 3707 5647 0 _1995_.C
rlabel metal2 3713 5613 3727 5627 0 _1995_.Y
rlabel metal1 3604 5522 3676 5538 0 _1994_.gnd
rlabel metal1 3604 5762 3676 5778 0 _1994_.vdd
rlabel metal2 3653 5593 3667 5607 0 _1994_.A
rlabel metal2 3633 5633 3647 5647 0 _1994_.Y
rlabel metal1 3504 5522 3616 5538 0 _2062_.gnd
rlabel metal1 3504 5762 3616 5778 0 _2062_.vdd
rlabel metal2 3593 5633 3607 5647 0 _2062_.A
rlabel metal2 3573 5653 3587 5667 0 _2062_.B
rlabel metal2 3553 5633 3567 5647 0 _2062_.C
rlabel metal2 3533 5653 3547 5667 0 _2062_.Y
rlabel metal1 3844 5522 3956 5538 0 _2012_.gnd
rlabel metal1 3844 5762 3956 5778 0 _2012_.vdd
rlabel metal2 3853 5613 3867 5627 0 _2012_.A
rlabel metal2 3873 5633 3887 5647 0 _2012_.B
rlabel metal2 3913 5633 3927 5647 0 _2012_.C
rlabel metal2 3893 5613 3907 5627 0 _2012_.Y
rlabel metal1 3764 5522 3856 5538 0 _1998_.gnd
rlabel metal1 3764 5762 3856 5778 0 _1998_.vdd
rlabel metal2 3793 5613 3807 5627 0 _1998_.B
rlabel metal2 3833 5613 3847 5627 0 _1998_.A
rlabel metal2 3813 5593 3827 5607 0 _1998_.Y
rlabel metal1 3944 5522 4016 5538 0 _2005_.gnd
rlabel metal1 3944 5762 4016 5778 0 _2005_.vdd
rlabel metal2 3993 5593 4007 5607 0 _2005_.A
rlabel metal2 3973 5633 3987 5647 0 _2005_.Y
rlabel metal1 4004 5522 4136 5538 0 _2047_.gnd
rlabel metal1 4004 5762 4136 5778 0 _2047_.vdd
rlabel metal2 4113 5613 4127 5627 0 _2047_.A
rlabel metal2 4093 5633 4107 5647 0 _2047_.B
rlabel metal2 4033 5613 4047 5627 0 _2047_.C
rlabel metal2 4053 5633 4067 5647 0 _2047_.D
rlabel metal2 4073 5613 4087 5627 0 _2047_.Y
rlabel metal1 4124 5522 4236 5538 0 _1988_.gnd
rlabel metal1 4124 5762 4236 5778 0 _1988_.vdd
rlabel metal2 4213 5613 4227 5627 0 _1988_.A
rlabel metal2 4193 5633 4207 5647 0 _1988_.B
rlabel metal2 4153 5633 4167 5647 0 _1988_.C
rlabel metal2 4173 5613 4187 5627 0 _1988_.Y
rlabel metal1 4224 5522 4336 5538 0 _1933_.gnd
rlabel metal1 4224 5762 4336 5778 0 _1933_.vdd
rlabel metal2 4313 5633 4327 5647 0 _1933_.A
rlabel metal2 4293 5653 4307 5667 0 _1933_.B
rlabel metal2 4273 5633 4287 5647 0 _1933_.C
rlabel metal2 4253 5653 4267 5667 0 _1933_.Y
rlabel metal1 4384 5522 4496 5538 0 _2003_.gnd
rlabel metal1 4384 5762 4496 5778 0 _2003_.vdd
rlabel metal2 4473 5613 4487 5627 0 _2003_.A
rlabel metal2 4453 5633 4467 5647 0 _2003_.B
rlabel metal2 4413 5633 4427 5647 0 _2003_.C
rlabel metal2 4433 5613 4447 5627 0 _2003_.Y
rlabel metal1 4324 5522 4396 5538 0 _1928_.gnd
rlabel metal1 4324 5762 4396 5778 0 _1928_.vdd
rlabel metal2 4333 5593 4347 5607 0 _1928_.A
rlabel metal2 4353 5633 4367 5647 0 _1928_.Y
rlabel metal1 4484 5522 4596 5538 0 _1942_.gnd
rlabel metal1 4484 5762 4596 5778 0 _1942_.vdd
rlabel metal2 4573 5613 4587 5627 0 _1942_.A
rlabel metal2 4513 5613 4527 5627 0 _1942_.Y
rlabel metal2 4533 5653 4547 5667 0 _1942_.B
rlabel metal1 4664 5522 4776 5538 0 _1949_.gnd
rlabel metal1 4664 5762 4776 5778 0 _1949_.vdd
rlabel metal2 4753 5613 4767 5627 0 _1949_.A
rlabel metal2 4733 5633 4747 5647 0 _1949_.B
rlabel metal2 4693 5633 4707 5647 0 _1949_.C
rlabel metal2 4713 5613 4727 5627 0 _1949_.Y
rlabel metal1 4764 5522 4876 5538 0 _1943_.gnd
rlabel metal1 4764 5762 4876 5778 0 _1943_.vdd
rlabel metal2 4773 5613 4787 5627 0 _1943_.A
rlabel metal2 4793 5633 4807 5647 0 _1943_.B
rlabel metal2 4833 5633 4847 5647 0 _1943_.C
rlabel metal2 4813 5613 4827 5627 0 _1943_.Y
rlabel metal1 4584 5522 4676 5538 0 _1948_.gnd
rlabel metal1 4584 5762 4676 5778 0 _1948_.vdd
rlabel metal2 4593 5653 4607 5667 0 _1948_.A
rlabel metal2 4633 5653 4647 5667 0 _1948_.B
rlabel metal2 4613 5633 4627 5647 0 _1948_.Y
rlabel metal1 5064 5522 5176 5538 0 _1880_.gnd
rlabel metal1 5064 5762 5176 5778 0 _1880_.vdd
rlabel metal2 5073 5613 5087 5627 0 _1880_.A
rlabel metal2 5093 5633 5107 5647 0 _1880_.B
rlabel metal2 5133 5633 5147 5647 0 _1880_.C
rlabel metal2 5113 5613 5127 5627 0 _1880_.Y
rlabel metal1 4964 5522 5076 5538 0 _1945_.gnd
rlabel metal1 4964 5762 5076 5778 0 _1945_.vdd
rlabel metal2 4973 5633 4987 5647 0 _1945_.A
rlabel metal2 4993 5593 5007 5607 0 _1945_.B
rlabel metal2 5013 5633 5027 5647 0 _1945_.C
rlabel metal2 5033 5613 5047 5627 0 _1945_.Y
rlabel metal1 4864 5522 4976 5538 0 _1954_.gnd
rlabel metal1 4864 5762 4976 5778 0 _1954_.vdd
rlabel metal2 4953 5633 4967 5647 0 _1954_.A
rlabel metal2 4933 5653 4947 5667 0 _1954_.B
rlabel metal2 4913 5633 4927 5647 0 _1954_.C
rlabel metal2 4893 5653 4907 5667 0 _1954_.Y
rlabel metal1 5264 5522 5356 5538 0 _1872_.gnd
rlabel metal1 5264 5762 5356 5778 0 _1872_.vdd
rlabel metal2 5273 5653 5287 5667 0 _1872_.A
rlabel metal2 5313 5653 5327 5667 0 _1872_.B
rlabel metal2 5293 5633 5307 5647 0 _1872_.Y
rlabel metal1 5164 5522 5276 5538 0 _1874_.gnd
rlabel metal1 5164 5762 5276 5778 0 _1874_.vdd
rlabel metal2 5173 5633 5187 5647 0 _1874_.A
rlabel metal2 5193 5653 5207 5667 0 _1874_.B
rlabel metal2 5213 5633 5227 5647 0 _1874_.C
rlabel metal2 5233 5653 5247 5667 0 _1874_.Y
rlabel metal1 5544 5522 5636 5538 0 _1910_.gnd
rlabel metal1 5544 5762 5636 5778 0 _1910_.vdd
rlabel metal2 5553 5653 5567 5667 0 _1910_.A
rlabel metal2 5593 5653 5607 5667 0 _1910_.B
rlabel metal2 5573 5633 5587 5647 0 _1910_.Y
rlabel metal1 5444 5522 5556 5538 0 _1876_.gnd
rlabel metal1 5444 5762 5556 5778 0 _1876_.vdd
rlabel metal2 5453 5633 5467 5647 0 _1876_.A
rlabel metal2 5473 5593 5487 5607 0 _1876_.B
rlabel metal2 5493 5633 5507 5647 0 _1876_.C
rlabel metal2 5513 5613 5527 5627 0 _1876_.Y
rlabel metal1 5344 5522 5456 5538 0 _1885_.gnd
rlabel metal1 5344 5762 5456 5778 0 _1885_.vdd
rlabel metal2 5353 5633 5367 5647 0 _1885_.A
rlabel metal2 5373 5653 5387 5667 0 _1885_.B
rlabel metal2 5393 5633 5407 5647 0 _1885_.C
rlabel metal2 5413 5653 5427 5667 0 _1885_.Y
rlabel metal1 5824 5522 5936 5538 0 _1871_.gnd
rlabel metal1 5824 5762 5936 5778 0 _1871_.vdd
rlabel metal2 5913 5613 5927 5627 0 _1871_.A
rlabel metal2 5893 5633 5907 5647 0 _1871_.B
rlabel metal2 5853 5633 5867 5647 0 _1871_.C
rlabel metal2 5873 5613 5887 5627 0 _1871_.Y
rlabel metal1 5624 5522 5716 5538 0 _1818_.gnd
rlabel metal1 5624 5762 5716 5778 0 _1818_.vdd
rlabel metal2 5693 5653 5707 5667 0 _1818_.A
rlabel metal2 5653 5653 5667 5667 0 _1818_.B
rlabel metal2 5673 5633 5687 5647 0 _1818_.Y
rlabel metal1 5704 5522 5836 5538 0 _1883_.gnd
rlabel metal1 5704 5762 5836 5778 0 _1883_.vdd
rlabel metal2 5713 5613 5727 5627 0 _1883_.A
rlabel metal2 5733 5633 5747 5647 0 _1883_.B
rlabel metal2 5793 5613 5807 5627 0 _1883_.C
rlabel metal2 5773 5633 5787 5647 0 _1883_.D
rlabel metal2 5753 5613 5767 5627 0 _1883_.Y
rlabel metal1 5924 5522 5996 5538 0 _1815_.gnd
rlabel metal1 5924 5762 5996 5778 0 _1815_.vdd
rlabel metal2 5933 5593 5947 5607 0 _1815_.A
rlabel metal2 5953 5633 5967 5647 0 _1815_.Y
rlabel metal1 6104 5522 6216 5538 0 _1821_.gnd
rlabel metal1 6104 5762 6216 5778 0 _1821_.vdd
rlabel metal2 6113 5633 6127 5647 0 _1821_.A
rlabel metal2 6133 5653 6147 5667 0 _1821_.B
rlabel metal2 6153 5633 6167 5647 0 _1821_.C
rlabel metal2 6173 5653 6187 5667 0 _1821_.Y
rlabel metal1 5984 5522 6116 5538 0 _1828_.gnd
rlabel metal1 5984 5762 6116 5778 0 _1828_.vdd
rlabel metal2 5993 5613 6007 5627 0 _1828_.A
rlabel metal2 6013 5633 6027 5647 0 _1828_.B
rlabel metal2 6073 5613 6087 5627 0 _1828_.C
rlabel metal2 6053 5633 6067 5647 0 _1828_.D
rlabel metal2 6033 5613 6047 5627 0 _1828_.Y
rlabel metal1 6204 5522 6276 5538 0 _1777_.gnd
rlabel metal1 6204 5762 6276 5778 0 _1777_.vdd
rlabel metal2 6253 5593 6267 5607 0 _1777_.A
rlabel metal2 6233 5633 6247 5647 0 _1777_.Y
rlabel metal1 6264 5522 6376 5538 0 _1856_.gnd
rlabel metal1 6264 5762 6376 5778 0 _1856_.vdd
rlabel metal2 6273 5633 6287 5647 0 _1856_.A
rlabel metal2 6293 5593 6307 5607 0 _1856_.B
rlabel metal2 6313 5633 6327 5647 0 _1856_.C
rlabel metal2 6333 5613 6347 5627 0 _1856_.Y
rlabel metal1 6364 5522 6476 5538 0 _1826_.gnd
rlabel metal1 6364 5762 6476 5778 0 _1826_.vdd
rlabel metal2 6373 5633 6387 5647 0 _1826_.A
rlabel metal2 6393 5653 6407 5667 0 _1826_.B
rlabel metal2 6413 5633 6427 5647 0 _1826_.C
rlabel metal2 6433 5653 6447 5667 0 _1826_.Y
rlabel nsubstratencontact 6676 5768 6676 5768 0 FILL100050x82950.vdd
rlabel metal1 6664 5522 6696 5538 0 FILL100050x82950.gnd
rlabel metal1 6564 5522 6676 5538 0 _1834_.gnd
rlabel metal1 6564 5762 6676 5778 0 _1834_.vdd
rlabel metal2 6573 5633 6587 5647 0 _1834_.A
rlabel metal2 6593 5653 6607 5667 0 _1834_.B
rlabel metal2 6613 5633 6627 5647 0 _1834_.C
rlabel metal2 6633 5653 6647 5667 0 _1834_.Y
rlabel metal1 6464 5522 6576 5538 0 _1833_.gnd
rlabel metal1 6464 5762 6576 5778 0 _1833_.vdd
rlabel metal2 6473 5633 6487 5647 0 _1833_.A
rlabel metal2 6493 5653 6507 5667 0 _1833_.B
rlabel metal2 6513 5633 6527 5647 0 _1833_.C
rlabel metal2 6533 5653 6547 5667 0 _1833_.Y
rlabel nsubstratencontact 6716 5768 6716 5768 0 FILL100650x82950.vdd
rlabel metal1 6704 5522 6736 5538 0 FILL100650x82950.gnd
rlabel nsubstratencontact 6696 5768 6696 5768 0 FILL100350x82950.vdd
rlabel metal1 6684 5522 6716 5538 0 FILL100350x82950.gnd
rlabel metal1 4 6002 96 6018 0 _3046_.gnd
rlabel metal1 4 5762 96 5778 0 _3046_.vdd
rlabel metal2 73 5913 87 5927 0 _3046_.A
rlabel metal2 33 5913 47 5927 0 _3046_.Y
rlabel metal1 164 6002 256 6018 0 _1540_.gnd
rlabel metal1 164 5762 256 5778 0 _1540_.vdd
rlabel metal2 173 5873 187 5887 0 _1540_.A
rlabel metal2 213 5873 227 5887 0 _1540_.B
rlabel metal2 193 5893 207 5907 0 _1540_.Y
rlabel metal1 84 6002 176 6018 0 _1537_.gnd
rlabel metal1 84 5762 176 5778 0 _1537_.vdd
rlabel metal2 93 5873 107 5887 0 _1537_.A
rlabel metal2 133 5873 147 5887 0 _1537_.B
rlabel metal2 113 5893 127 5907 0 _1537_.Y
rlabel metal1 244 6002 356 6018 0 _1586_.gnd
rlabel metal1 244 5762 356 5778 0 _1586_.vdd
rlabel metal2 333 5893 347 5907 0 _1586_.A
rlabel metal2 313 5933 327 5947 0 _1586_.B
rlabel metal2 293 5893 307 5907 0 _1586_.C
rlabel metal2 273 5913 287 5927 0 _1586_.Y
rlabel metal1 484 6002 576 6018 0 _2295_.gnd
rlabel metal1 484 5762 576 5778 0 _2295_.vdd
rlabel metal2 513 5913 527 5927 0 _2295_.B
rlabel metal2 553 5913 567 5927 0 _2295_.A
rlabel metal2 533 5933 547 5947 0 _2295_.Y
rlabel metal1 424 6002 496 6018 0 _2291_.gnd
rlabel metal1 424 5762 496 5778 0 _2291_.vdd
rlabel metal2 433 5933 447 5947 0 _2291_.A
rlabel metal2 453 5893 467 5907 0 _2291_.Y
rlabel metal1 344 6002 436 6018 0 _1542_.gnd
rlabel metal1 344 5762 436 5778 0 _1542_.vdd
rlabel metal2 413 5873 427 5887 0 _1542_.A
rlabel metal2 373 5873 387 5887 0 _1542_.B
rlabel metal2 393 5893 407 5907 0 _1542_.Y
rlabel metal1 644 6002 756 6018 0 _2300_.gnd
rlabel metal1 644 5762 756 5778 0 _2300_.vdd
rlabel metal2 653 5913 667 5927 0 _2300_.A
rlabel metal2 673 5893 687 5907 0 _2300_.B
rlabel metal2 713 5893 727 5907 0 _2300_.C
rlabel metal2 693 5913 707 5927 0 _2300_.Y
rlabel metal1 564 6002 656 6018 0 _2292_.gnd
rlabel metal1 564 5762 656 5778 0 _2292_.vdd
rlabel metal2 613 5913 627 5927 0 _2292_.B
rlabel metal2 573 5913 587 5927 0 _2292_.A
rlabel metal2 593 5933 607 5947 0 _2292_.Y
rlabel metal1 744 6002 816 6018 0 _2286_.gnd
rlabel metal1 744 5762 816 5778 0 _2286_.vdd
rlabel metal2 793 5933 807 5947 0 _2286_.A
rlabel metal2 773 5893 787 5907 0 _2286_.Y
rlabel metal1 964 6002 1076 6018 0 _2275_.gnd
rlabel metal1 964 5762 1076 5778 0 _2275_.vdd
rlabel metal2 1053 5913 1067 5927 0 _2275_.A
rlabel metal2 1033 5893 1047 5907 0 _2275_.B
rlabel metal2 993 5893 1007 5907 0 _2275_.C
rlabel metal2 1013 5913 1027 5927 0 _2275_.Y
rlabel metal1 804 6002 896 6018 0 _2287_.gnd
rlabel metal1 804 5762 896 5778 0 _2287_.vdd
rlabel metal2 853 5913 867 5927 0 _2287_.B
rlabel metal2 813 5913 827 5927 0 _2287_.A
rlabel metal2 833 5933 847 5947 0 _2287_.Y
rlabel metal1 1064 6002 1156 6018 0 _2262_.gnd
rlabel metal1 1064 5762 1156 5778 0 _2262_.vdd
rlabel metal2 1113 5913 1127 5927 0 _2262_.B
rlabel metal2 1073 5913 1087 5927 0 _2262_.A
rlabel metal2 1093 5933 1107 5947 0 _2262_.Y
rlabel metal1 884 6002 976 6018 0 _2122_.gnd
rlabel metal1 884 5762 976 5778 0 _2122_.vdd
rlabel metal2 953 5873 967 5887 0 _2122_.A
rlabel metal2 913 5873 927 5887 0 _2122_.B
rlabel metal2 933 5893 947 5907 0 _2122_.Y
rlabel metal1 1204 6002 1456 6018 0 _2377_.gnd
rlabel metal1 1204 5762 1456 5778 0 _2377_.vdd
rlabel metal2 1353 5913 1367 5927 0 _2377_.D
rlabel metal2 1313 5913 1327 5927 0 _2377_.CLK
rlabel metal2 1233 5913 1247 5927 0 _2377_.Q
rlabel metal1 1144 6002 1216 6018 0 _2274_.gnd
rlabel metal1 1144 5762 1216 5778 0 _2274_.vdd
rlabel metal2 1193 5933 1207 5947 0 _2274_.A
rlabel metal2 1173 5893 1187 5907 0 _2274_.Y
rlabel metal1 1444 6002 1536 6018 0 _2149_.gnd
rlabel metal1 1444 5762 1536 5778 0 _2149_.vdd
rlabel metal2 1453 5873 1467 5887 0 _2149_.A
rlabel metal2 1493 5873 1507 5887 0 _2149_.B
rlabel metal2 1473 5893 1487 5907 0 _2149_.Y
rlabel metal1 1524 6002 1636 6018 0 _2148_.gnd
rlabel metal1 1524 5762 1636 5778 0 _2148_.vdd
rlabel metal2 1613 5893 1627 5907 0 _2148_.A
rlabel metal2 1593 5873 1607 5887 0 _2148_.B
rlabel metal2 1573 5893 1587 5907 0 _2148_.C
rlabel metal2 1553 5873 1567 5887 0 _2148_.Y
rlabel metal1 1624 6002 1736 6018 0 _2154_.gnd
rlabel metal1 1624 5762 1736 5778 0 _2154_.vdd
rlabel metal2 1713 5913 1727 5927 0 _2154_.A
rlabel metal2 1693 5893 1707 5907 0 _2154_.B
rlabel metal2 1653 5893 1667 5907 0 _2154_.C
rlabel metal2 1673 5913 1687 5927 0 _2154_.Y
rlabel metal1 1724 6002 1816 6018 0 _2153_.gnd
rlabel metal1 1724 5762 1816 5778 0 _2153_.vdd
rlabel metal2 1753 5913 1767 5927 0 _2153_.B
rlabel metal2 1793 5913 1807 5927 0 _2153_.A
rlabel metal2 1773 5933 1787 5947 0 _2153_.Y
rlabel metal1 1804 6002 1916 6018 0 _2140_.gnd
rlabel metal1 1804 5762 1916 5778 0 _2140_.vdd
rlabel metal2 1893 5893 1907 5907 0 _2140_.A
rlabel metal2 1873 5873 1887 5887 0 _2140_.B
rlabel metal2 1853 5893 1867 5907 0 _2140_.C
rlabel metal2 1833 5873 1847 5887 0 _2140_.Y
rlabel metal1 1964 6002 2076 6018 0 _2147_.gnd
rlabel metal1 1964 5762 2076 5778 0 _2147_.vdd
rlabel metal2 2053 5913 2067 5927 0 _2147_.A
rlabel metal2 2033 5893 2047 5907 0 _2147_.B
rlabel metal2 1993 5893 2007 5907 0 _2147_.C
rlabel metal2 2013 5913 2027 5927 0 _2147_.Y
rlabel metal1 1904 6002 1976 6018 0 _2144_.gnd
rlabel metal1 1904 5762 1976 5778 0 _2144_.vdd
rlabel metal2 1913 5933 1927 5947 0 _2144_.A
rlabel metal2 1933 5893 1947 5907 0 _2144_.Y
rlabel metal1 2064 6002 2176 6018 0 _2165_.gnd
rlabel metal1 2064 5762 2176 5778 0 _2165_.vdd
rlabel metal2 2073 5893 2087 5907 0 _2165_.A
rlabel metal2 2093 5873 2107 5887 0 _2165_.B
rlabel metal2 2113 5893 2127 5907 0 _2165_.C
rlabel metal2 2133 5873 2147 5887 0 _2165_.Y
rlabel metal1 2264 6002 2376 6018 0 _2143_.gnd
rlabel metal1 2264 5762 2376 5778 0 _2143_.vdd
rlabel metal2 2273 5913 2287 5927 0 _2143_.A
rlabel metal2 2293 5893 2307 5907 0 _2143_.B
rlabel metal2 2333 5893 2347 5907 0 _2143_.C
rlabel metal2 2313 5913 2327 5927 0 _2143_.Y
rlabel metal1 2364 6002 2456 6018 0 _2118_.gnd
rlabel metal1 2364 5762 2456 5778 0 _2118_.vdd
rlabel metal2 2433 5873 2447 5887 0 _2118_.A
rlabel metal2 2393 5873 2407 5887 0 _2118_.B
rlabel metal2 2413 5893 2427 5907 0 _2118_.Y
rlabel metal1 2164 6002 2276 6018 0 _2145_.gnd
rlabel metal1 2164 5762 2276 5778 0 _2145_.vdd
rlabel metal2 2253 5893 2267 5907 0 _2145_.A
rlabel metal2 2233 5933 2247 5947 0 _2145_.B
rlabel metal2 2213 5893 2227 5907 0 _2145_.C
rlabel metal2 2193 5913 2207 5927 0 _2145_.Y
rlabel metal1 2644 6002 2736 6018 0 _2116_.gnd
rlabel metal1 2644 5762 2736 5778 0 _2116_.vdd
rlabel metal2 2653 5873 2667 5887 0 _2116_.A
rlabel metal2 2693 5873 2707 5887 0 _2116_.B
rlabel metal2 2673 5893 2687 5907 0 _2116_.Y
rlabel metal1 2544 6002 2656 6018 0 _2141_.gnd
rlabel metal1 2544 5762 2656 5778 0 _2141_.vdd
rlabel metal2 2633 5893 2647 5907 0 _2141_.A
rlabel metal2 2613 5933 2627 5947 0 _2141_.B
rlabel metal2 2593 5893 2607 5907 0 _2141_.C
rlabel metal2 2573 5913 2587 5927 0 _2141_.Y
rlabel metal1 2444 6002 2556 6018 0 _2115_.gnd
rlabel metal1 2444 5762 2556 5778 0 _2115_.vdd
rlabel metal2 2533 5893 2547 5907 0 _2115_.A
rlabel metal2 2513 5873 2527 5887 0 _2115_.B
rlabel metal2 2493 5893 2507 5907 0 _2115_.C
rlabel metal2 2473 5873 2487 5887 0 _2115_.Y
rlabel metal1 2924 6002 3036 6018 0 _2078_.gnd
rlabel metal1 2924 5762 3036 5778 0 _2078_.vdd
rlabel metal2 3013 5893 3027 5907 0 _2078_.A
rlabel metal2 2993 5873 3007 5887 0 _2078_.B
rlabel metal2 2973 5893 2987 5907 0 _2078_.C
rlabel metal2 2953 5873 2967 5887 0 _2078_.Y
rlabel metal1 2724 6002 2836 6018 0 _2077_.gnd
rlabel metal1 2724 5762 2836 5778 0 _2077_.vdd
rlabel metal2 2813 5893 2827 5907 0 _2077_.A
rlabel metal2 2793 5873 2807 5887 0 _2077_.B
rlabel metal2 2773 5893 2787 5907 0 _2077_.C
rlabel metal2 2753 5873 2767 5887 0 _2077_.Y
rlabel metal1 2824 6002 2936 6018 0 _2070_.gnd
rlabel metal1 2824 5762 2936 5778 0 _2070_.vdd
rlabel metal2 2913 5893 2927 5907 0 _2070_.A
rlabel metal2 2893 5873 2907 5887 0 _2070_.B
rlabel metal2 2873 5893 2887 5907 0 _2070_.C
rlabel metal2 2853 5873 2867 5887 0 _2070_.Y
rlabel metal1 3124 6002 3236 6018 0 _2073_.gnd
rlabel metal1 3124 5762 3236 5778 0 _2073_.vdd
rlabel metal2 3133 5893 3147 5907 0 _2073_.A
rlabel metal2 3153 5873 3167 5887 0 _2073_.B
rlabel metal2 3173 5893 3187 5907 0 _2073_.C
rlabel metal2 3193 5873 3207 5887 0 _2073_.Y
rlabel metal1 3024 6002 3136 6018 0 _2064_.gnd
rlabel metal1 3024 5762 3136 5778 0 _2064_.vdd
rlabel metal2 3113 5893 3127 5907 0 _2064_.A
rlabel metal2 3093 5873 3107 5887 0 _2064_.B
rlabel metal2 3073 5893 3087 5907 0 _2064_.C
rlabel metal2 3053 5873 3067 5887 0 _2064_.Y
rlabel metal1 3324 6002 3436 6018 0 _2072_.gnd
rlabel metal1 3324 5762 3436 5778 0 _2072_.vdd
rlabel metal2 3333 5913 3347 5927 0 _2072_.A
rlabel metal2 3353 5893 3367 5907 0 _2072_.B
rlabel metal2 3393 5893 3407 5907 0 _2072_.C
rlabel metal2 3373 5913 3387 5927 0 _2072_.Y
rlabel metal1 3224 6002 3336 6018 0 _2069_.gnd
rlabel metal1 3224 5762 3336 5778 0 _2069_.vdd
rlabel metal2 3313 5913 3327 5927 0 _2069_.A
rlabel metal2 3293 5893 3307 5907 0 _2069_.B
rlabel metal2 3253 5893 3267 5907 0 _2069_.C
rlabel metal2 3273 5913 3287 5927 0 _2069_.Y
rlabel metal1 3424 6002 3536 6018 0 _2067_.gnd
rlabel metal1 3424 5762 3536 5778 0 _2067_.vdd
rlabel metal2 3513 5893 3527 5907 0 _2067_.A
rlabel metal2 3493 5933 3507 5947 0 _2067_.B
rlabel metal2 3473 5893 3487 5907 0 _2067_.C
rlabel metal2 3453 5913 3467 5927 0 _2067_.Y
rlabel metal1 3524 6002 3636 6018 0 _2046_.gnd
rlabel metal1 3524 5762 3636 5778 0 _2046_.vdd
rlabel metal2 3613 5913 3627 5927 0 _2046_.A
rlabel metal2 3593 5893 3607 5907 0 _2046_.B
rlabel metal2 3553 5893 3567 5907 0 _2046_.C
rlabel metal2 3573 5913 3587 5927 0 _2046_.Y
rlabel metal1 3724 6002 3836 6018 0 _2014_.gnd
rlabel metal1 3724 5762 3836 5778 0 _2014_.vdd
rlabel metal2 3733 5893 3747 5907 0 _2014_.A
rlabel metal2 3753 5933 3767 5947 0 _2014_.B
rlabel metal2 3773 5893 3787 5907 0 _2014_.C
rlabel metal2 3793 5913 3807 5927 0 _2014_.Y
rlabel metal1 3624 6002 3736 6018 0 _2022_.gnd
rlabel metal1 3624 5762 3736 5778 0 _2022_.vdd
rlabel metal2 3713 5893 3727 5907 0 _2022_.A
rlabel metal2 3693 5873 3707 5887 0 _2022_.B
rlabel metal2 3673 5893 3687 5907 0 _2022_.C
rlabel metal2 3653 5873 3667 5887 0 _2022_.Y
rlabel metal1 3924 6002 4036 6018 0 _2045_.gnd
rlabel metal1 3924 5762 4036 5778 0 _2045_.vdd
rlabel metal2 4013 5893 4027 5907 0 _2045_.A
rlabel metal2 3993 5933 4007 5947 0 _2045_.B
rlabel metal2 3973 5893 3987 5907 0 _2045_.C
rlabel metal2 3953 5913 3967 5927 0 _2045_.Y
rlabel metal1 3824 6002 3936 6018 0 _2016_.gnd
rlabel metal1 3824 5762 3936 5778 0 _2016_.vdd
rlabel metal2 3913 5893 3927 5907 0 _2016_.A
rlabel metal2 3893 5873 3907 5887 0 _2016_.B
rlabel metal2 3873 5893 3887 5907 0 _2016_.C
rlabel metal2 3853 5873 3867 5887 0 _2016_.Y
rlabel metal1 4124 6002 4236 6018 0 _2007_.gnd
rlabel metal1 4124 5762 4236 5778 0 _2007_.vdd
rlabel metal2 4213 5893 4227 5907 0 _2007_.A
rlabel metal2 4193 5933 4207 5947 0 _2007_.B
rlabel metal2 4173 5893 4187 5907 0 _2007_.C
rlabel metal2 4153 5913 4167 5927 0 _2007_.Y
rlabel metal1 4024 6002 4136 6018 0 _2013_.gnd
rlabel metal1 4024 5762 4136 5778 0 _2013_.vdd
rlabel metal2 4113 5893 4127 5907 0 _2013_.A
rlabel metal2 4093 5873 4107 5887 0 _2013_.B
rlabel metal2 4073 5893 4087 5907 0 _2013_.C
rlabel metal2 4053 5873 4067 5887 0 _2013_.Y
rlabel metal1 4224 6002 4336 6018 0 _2011_.gnd
rlabel metal1 4224 5762 4336 5778 0 _2011_.vdd
rlabel metal2 4233 5893 4247 5907 0 _2011_.A
rlabel metal2 4253 5873 4267 5887 0 _2011_.B
rlabel metal2 4273 5893 4287 5907 0 _2011_.C
rlabel metal2 4293 5873 4307 5887 0 _2011_.Y
rlabel metal1 4404 6002 4516 6018 0 _1997_.gnd
rlabel metal1 4404 5762 4516 5778 0 _1997_.vdd
rlabel metal2 4493 5913 4507 5927 0 _1997_.A
rlabel metal2 4473 5893 4487 5907 0 _1997_.B
rlabel metal2 4433 5893 4447 5907 0 _1997_.C
rlabel metal2 4453 5913 4467 5927 0 _1997_.Y
rlabel metal1 4504 6002 4596 6018 0 _1996_.gnd
rlabel metal1 4504 5762 4596 5778 0 _1996_.vdd
rlabel metal2 4533 5913 4547 5927 0 _1996_.B
rlabel metal2 4573 5913 4587 5927 0 _1996_.A
rlabel metal2 4553 5933 4567 5947 0 _1996_.Y
rlabel metal1 4324 6002 4416 6018 0 _2006_.gnd
rlabel metal1 4324 5762 4416 5778 0 _2006_.vdd
rlabel metal2 4333 5873 4347 5887 0 _2006_.A
rlabel metal2 4373 5873 4387 5887 0 _2006_.B
rlabel metal2 4353 5893 4367 5907 0 _2006_.Y
rlabel metal1 4784 6002 4876 6018 0 _1947_.gnd
rlabel metal1 4784 5762 4876 5778 0 _1947_.vdd
rlabel metal2 4793 5873 4807 5887 0 _1947_.A
rlabel metal2 4833 5873 4847 5887 0 _1947_.B
rlabel metal2 4813 5893 4827 5907 0 _1947_.Y
rlabel metal1 4684 6002 4796 6018 0 _2010_.gnd
rlabel metal1 4684 5762 4796 5778 0 _2010_.vdd
rlabel metal2 4773 5893 4787 5907 0 _2010_.A
rlabel metal2 4753 5933 4767 5947 0 _2010_.B
rlabel metal2 4733 5893 4747 5907 0 _2010_.C
rlabel metal2 4713 5913 4727 5927 0 _2010_.Y
rlabel metal1 4584 6002 4696 6018 0 _2009_.gnd
rlabel metal1 4584 5762 4696 5778 0 _2009_.vdd
rlabel metal2 4593 5913 4607 5927 0 _2009_.A
rlabel metal2 4653 5913 4667 5927 0 _2009_.Y
rlabel metal2 4633 5873 4647 5887 0 _2009_.B
rlabel metal1 4864 6002 4936 6018 0 _1946_.gnd
rlabel metal1 4864 5762 4936 5778 0 _1946_.vdd
rlabel metal2 4913 5933 4927 5947 0 _1946_.A
rlabel metal2 4893 5893 4907 5907 0 _1946_.Y
rlabel metal1 5024 6002 5136 6018 0 _1950_.gnd
rlabel metal1 5024 5762 5136 5778 0 _1950_.vdd
rlabel metal2 5033 5893 5047 5907 0 _1950_.A
rlabel metal2 5053 5933 5067 5947 0 _1950_.B
rlabel metal2 5073 5893 5087 5907 0 _1950_.C
rlabel metal2 5093 5913 5107 5927 0 _1950_.Y
rlabel metal1 4924 6002 5036 6018 0 _1953_.gnd
rlabel metal1 4924 5762 5036 5778 0 _1953_.vdd
rlabel metal2 5013 5893 5027 5907 0 _1953_.A
rlabel metal2 4993 5873 5007 5887 0 _1953_.B
rlabel metal2 4973 5893 4987 5907 0 _1953_.C
rlabel metal2 4953 5873 4967 5887 0 _1953_.Y
rlabel metal1 5124 6002 5236 6018 0 _1959_.gnd
rlabel metal1 5124 5762 5236 5778 0 _1959_.vdd
rlabel metal2 5133 5913 5147 5927 0 _1959_.A
rlabel metal2 5153 5893 5167 5907 0 _1959_.B
rlabel metal2 5193 5893 5207 5907 0 _1959_.C
rlabel metal2 5173 5913 5187 5927 0 _1959_.Y
rlabel metal1 5224 6002 5336 6018 0 _1940_.gnd
rlabel metal1 5224 5762 5336 5778 0 _1940_.vdd
rlabel metal2 5233 5913 5247 5927 0 _1940_.A
rlabel metal2 5253 5893 5267 5907 0 _1940_.B
rlabel metal2 5293 5893 5307 5907 0 _1940_.C
rlabel metal2 5273 5913 5287 5927 0 _1940_.Y
rlabel metal1 5324 6002 5456 6018 0 _1952_.gnd
rlabel metal1 5324 5762 5456 5778 0 _1952_.vdd
rlabel metal2 5333 5913 5347 5927 0 _1952_.A
rlabel metal2 5353 5893 5367 5907 0 _1952_.B
rlabel metal2 5413 5913 5427 5927 0 _1952_.C
rlabel metal2 5393 5893 5407 5907 0 _1952_.D
rlabel metal2 5373 5913 5387 5927 0 _1952_.Y
rlabel metal1 5524 6002 5596 6018 0 _1877_.gnd
rlabel metal1 5524 5762 5596 5778 0 _1877_.vdd
rlabel metal2 5533 5933 5547 5947 0 _1877_.A
rlabel metal2 5553 5893 5567 5907 0 _1877_.Y
rlabel metal1 5444 6002 5536 6018 0 _1879_.gnd
rlabel metal1 5444 5762 5536 5778 0 _1879_.vdd
rlabel metal2 5513 5873 5527 5887 0 _1879_.A
rlabel metal2 5473 5873 5487 5887 0 _1879_.B
rlabel metal2 5493 5893 5507 5907 0 _1879_.Y
rlabel metal1 5584 6002 5696 6018 0 _1884_.gnd
rlabel metal1 5584 5762 5696 5778 0 _1884_.vdd
rlabel metal2 5673 5893 5687 5907 0 _1884_.A
rlabel metal2 5653 5873 5667 5887 0 _1884_.B
rlabel metal2 5633 5893 5647 5907 0 _1884_.C
rlabel metal2 5613 5873 5627 5887 0 _1884_.Y
rlabel metal1 5784 6002 5896 6018 0 _1890_.gnd
rlabel metal1 5784 5762 5896 5778 0 _1890_.vdd
rlabel metal2 5873 5913 5887 5927 0 _1890_.A
rlabel metal2 5853 5893 5867 5907 0 _1890_.B
rlabel metal2 5813 5893 5827 5907 0 _1890_.C
rlabel metal2 5833 5913 5847 5927 0 _1890_.Y
rlabel metal1 5684 6002 5796 6018 0 _1881_.gnd
rlabel metal1 5684 5762 5796 5778 0 _1881_.vdd
rlabel metal2 5693 5893 5707 5907 0 _1881_.A
rlabel metal2 5713 5933 5727 5947 0 _1881_.B
rlabel metal2 5733 5893 5747 5907 0 _1881_.C
rlabel metal2 5753 5913 5767 5927 0 _1881_.Y
rlabel metal1 5984 6002 6096 6018 0 _1903_.gnd
rlabel metal1 5984 5762 6096 5778 0 _1903_.vdd
rlabel metal2 6073 5913 6087 5927 0 _1903_.A
rlabel metal2 6053 5893 6067 5907 0 _1903_.B
rlabel metal2 6013 5893 6027 5907 0 _1903_.C
rlabel metal2 6033 5913 6047 5927 0 _1903_.Y
rlabel metal1 5884 6002 5996 6018 0 _1882_.gnd
rlabel metal1 5884 5762 5996 5778 0 _1882_.vdd
rlabel metal2 5893 5913 5907 5927 0 _1882_.A
rlabel metal2 5913 5893 5927 5907 0 _1882_.B
rlabel metal2 5953 5893 5967 5907 0 _1882_.C
rlabel metal2 5933 5913 5947 5927 0 _1882_.Y
rlabel metal1 6084 6002 6216 6018 0 _1898_.gnd
rlabel metal1 6084 5762 6216 5778 0 _1898_.vdd
rlabel metal2 6093 5913 6107 5927 0 _1898_.A
rlabel metal2 6113 5893 6127 5907 0 _1898_.B
rlabel metal2 6173 5913 6187 5927 0 _1898_.C
rlabel metal2 6153 5893 6167 5907 0 _1898_.D
rlabel metal2 6133 5913 6147 5927 0 _1898_.Y
rlabel metal1 6384 6002 6496 6018 0 _1857_.gnd
rlabel metal1 6384 5762 6496 5778 0 _1857_.vdd
rlabel metal2 6393 5913 6407 5927 0 _1857_.A
rlabel metal2 6413 5893 6427 5907 0 _1857_.B
rlabel metal2 6453 5893 6467 5907 0 _1857_.C
rlabel metal2 6433 5913 6447 5927 0 _1857_.Y
rlabel metal1 6204 6002 6296 6018 0 _1831_.gnd
rlabel metal1 6204 5762 6296 5778 0 _1831_.vdd
rlabel metal2 6273 5873 6287 5887 0 _1831_.A
rlabel metal2 6233 5873 6247 5887 0 _1831_.B
rlabel metal2 6253 5893 6267 5907 0 _1831_.Y
rlabel metal1 6284 6002 6396 6018 0 _1813_.gnd
rlabel metal1 6284 5762 6396 5778 0 _1813_.vdd
rlabel metal2 6293 5913 6307 5927 0 _1813_.A
rlabel metal2 6353 5913 6367 5927 0 _1813_.Y
rlabel metal2 6333 5873 6347 5887 0 _1813_.B
rlabel nsubstratencontact 6684 5772 6684 5772 0 FILL100050x86550.vdd
rlabel metal1 6664 6002 6696 6018 0 FILL100050x86550.gnd
rlabel metal1 6584 6002 6676 6018 0 _1836_.gnd
rlabel metal1 6584 5762 6676 5778 0 _1836_.vdd
rlabel metal2 6593 5873 6607 5887 0 _1836_.A
rlabel metal2 6633 5873 6647 5887 0 _1836_.B
rlabel metal2 6613 5893 6627 5907 0 _1836_.Y
rlabel metal1 6484 6002 6596 6018 0 _1830_.gnd
rlabel metal1 6484 5762 6596 5778 0 _1830_.vdd
rlabel metal2 6493 5893 6507 5907 0 _1830_.A
rlabel metal2 6513 5873 6527 5887 0 _1830_.B
rlabel metal2 6533 5893 6547 5907 0 _1830_.C
rlabel metal2 6553 5873 6567 5887 0 _1830_.Y
rlabel nsubstratencontact 6724 5772 6724 5772 0 FILL100650x86550.vdd
rlabel metal1 6704 6002 6736 6018 0 FILL100650x86550.gnd
rlabel nsubstratencontact 6704 5772 6704 5772 0 FILL100350x86550.vdd
rlabel metal1 6684 6002 6716 6018 0 FILL100350x86550.gnd
rlabel metal1 4 6482 256 6498 0 _2390_.gnd
rlabel metal1 4 6242 256 6258 0 _2390_.vdd
rlabel metal2 93 6393 107 6407 0 _2390_.D
rlabel metal2 133 6393 147 6407 0 _2390_.CLK
rlabel metal2 213 6393 227 6407 0 _2390_.Q
rlabel metal1 4 6002 256 6018 0 _1617_.gnd
rlabel metal1 4 6242 256 6258 0 _1617_.vdd
rlabel metal2 153 6093 167 6107 0 _1617_.D
rlabel metal2 113 6093 127 6107 0 _1617_.CLK
rlabel metal2 33 6093 47 6107 0 _1617_.Q
rlabel metal1 244 6482 356 6498 0 _2298_.gnd
rlabel metal1 244 6242 356 6258 0 _2298_.vdd
rlabel metal2 333 6393 347 6407 0 _2298_.A
rlabel metal2 313 6373 327 6387 0 _2298_.B
rlabel metal2 273 6373 287 6387 0 _2298_.C
rlabel metal2 293 6393 307 6407 0 _2298_.Y
rlabel metal1 244 6002 356 6018 0 _1585_.gnd
rlabel metal1 244 6242 356 6258 0 _1585_.vdd
rlabel metal2 333 6113 347 6127 0 _1585_.A
rlabel metal2 313 6073 327 6087 0 _1585_.B
rlabel metal2 293 6113 307 6127 0 _1585_.C
rlabel metal2 273 6093 287 6107 0 _1585_.Y
rlabel metal1 424 6002 516 6018 0 _2293_.gnd
rlabel metal1 424 6242 516 6258 0 _2293_.vdd
rlabel metal2 473 6093 487 6107 0 _2293_.B
rlabel metal2 433 6093 447 6107 0 _2293_.A
rlabel metal2 453 6073 467 6087 0 _2293_.Y
rlabel metal1 504 6002 596 6018 0 _2297_.gnd
rlabel metal1 504 6242 596 6258 0 _2297_.vdd
rlabel metal2 573 6133 587 6147 0 _2297_.A
rlabel metal2 533 6133 547 6147 0 _2297_.B
rlabel metal2 553 6113 567 6127 0 _2297_.Y
rlabel metal1 344 6482 436 6498 0 _2284_.gnd
rlabel metal1 344 6242 436 6258 0 _2284_.vdd
rlabel metal2 353 6353 367 6367 0 _2284_.A
rlabel metal2 393 6353 407 6367 0 _2284_.B
rlabel metal2 373 6373 387 6387 0 _2284_.Y
rlabel metal1 424 6482 516 6498 0 _1541_.gnd
rlabel metal1 424 6242 516 6258 0 _1541_.vdd
rlabel metal2 493 6353 507 6367 0 _1541_.A
rlabel metal2 453 6353 467 6367 0 _1541_.B
rlabel metal2 473 6373 487 6387 0 _1541_.Y
rlabel metal1 344 6002 436 6018 0 _1539_.gnd
rlabel metal1 344 6242 436 6258 0 _1539_.vdd
rlabel metal2 413 6133 427 6147 0 _1539_.A
rlabel metal2 373 6133 387 6147 0 _1539_.B
rlabel metal2 393 6113 407 6127 0 _1539_.Y
rlabel metal1 504 6482 596 6498 0 _1538_.gnd
rlabel metal1 504 6242 596 6258 0 _1538_.vdd
rlabel metal2 513 6353 527 6367 0 _1538_.A
rlabel metal2 553 6353 567 6367 0 _1538_.B
rlabel metal2 533 6373 547 6387 0 _1538_.Y
rlabel metal1 584 6482 836 6498 0 _2389_.gnd
rlabel metal1 584 6242 836 6258 0 _2389_.vdd
rlabel metal2 733 6393 747 6407 0 _2389_.D
rlabel metal2 693 6393 707 6407 0 _2389_.CLK
rlabel metal2 613 6393 627 6407 0 _2389_.Q
rlabel metal1 684 6002 796 6018 0 _2296_.gnd
rlabel metal1 684 6242 796 6258 0 _2296_.vdd
rlabel metal2 773 6093 787 6107 0 _2296_.A
rlabel metal2 753 6113 767 6127 0 _2296_.B
rlabel metal2 713 6113 727 6127 0 _2296_.C
rlabel metal2 733 6093 747 6107 0 _2296_.Y
rlabel metal1 584 6002 696 6018 0 _2294_.gnd
rlabel metal1 584 6242 696 6258 0 _2294_.vdd
rlabel metal2 593 6093 607 6107 0 _2294_.A
rlabel metal2 613 6113 627 6127 0 _2294_.B
rlabel metal2 653 6113 667 6127 0 _2294_.C
rlabel metal2 633 6093 647 6107 0 _2294_.Y
rlabel metal1 784 6002 876 6018 0 _2290_.gnd
rlabel metal1 784 6242 876 6258 0 _2290_.vdd
rlabel metal2 833 6093 847 6107 0 _2290_.B
rlabel metal2 793 6093 807 6107 0 _2290_.A
rlabel metal2 813 6073 827 6087 0 _2290_.Y
rlabel metal1 1064 6482 1316 6498 0 _2376_.gnd
rlabel metal1 1064 6242 1316 6258 0 _2376_.vdd
rlabel metal2 1213 6393 1227 6407 0 _2376_.D
rlabel metal2 1173 6393 1187 6407 0 _2376_.CLK
rlabel metal2 1093 6393 1107 6407 0 _2376_.Q
rlabel metal1 824 6482 896 6498 0 _2273_.gnd
rlabel metal1 824 6242 896 6258 0 _2273_.vdd
rlabel metal2 833 6413 847 6427 0 _2273_.A
rlabel metal2 853 6373 867 6387 0 _2273_.Y
rlabel metal1 1064 6002 1136 6018 0 _2263_.gnd
rlabel metal1 1064 6242 1136 6258 0 _2263_.vdd
rlabel metal2 1113 6073 1127 6087 0 _2263_.A
rlabel metal2 1093 6113 1107 6127 0 _2263_.Y
rlabel metal1 1004 6482 1076 6498 0 _2090_.gnd
rlabel metal1 1004 6242 1076 6258 0 _2090_.vdd
rlabel metal2 1053 6413 1067 6427 0 _2090_.A
rlabel metal2 1033 6373 1047 6387 0 _2090_.Y
rlabel metal1 864 6002 976 6018 0 _2282_.gnd
rlabel metal1 864 6242 976 6258 0 _2282_.vdd
rlabel metal2 953 6113 967 6127 0 _2282_.A
rlabel metal2 933 6073 947 6087 0 _2282_.B
rlabel metal2 913 6113 927 6127 0 _2282_.C
rlabel metal2 893 6093 907 6107 0 _2282_.Y
rlabel metal1 964 6002 1076 6018 0 _2281_.gnd
rlabel metal1 964 6242 1076 6258 0 _2281_.vdd
rlabel metal2 973 6073 987 6087 0 _2281_.A
rlabel metal2 993 6093 1007 6107 0 _2281_.B
rlabel metal2 1033 6113 1047 6127 0 _2281_.Y
rlabel metal1 884 6482 1016 6498 0 _2283_.gnd
rlabel metal1 884 6242 1016 6258 0 _2283_.vdd
rlabel metal2 893 6393 907 6407 0 _2283_.A
rlabel metal2 913 6373 927 6387 0 _2283_.B
rlabel metal2 973 6393 987 6407 0 _2283_.C
rlabel metal2 953 6373 967 6387 0 _2283_.D
rlabel metal2 933 6393 947 6407 0 _2283_.Y
rlabel metal1 1304 6482 1436 6498 0 _2121_.gnd
rlabel metal1 1304 6242 1436 6258 0 _2121_.vdd
rlabel metal2 1313 6393 1327 6407 0 _2121_.A
rlabel metal2 1333 6373 1347 6387 0 _2121_.B
rlabel metal2 1393 6393 1407 6407 0 _2121_.C
rlabel metal2 1353 6393 1367 6407 0 _2121_.Y
rlabel metal2 1373 6373 1387 6387 0 _2121_.D
rlabel metal1 1204 6002 1316 6018 0 _2289_.gnd
rlabel metal1 1204 6242 1316 6258 0 _2289_.vdd
rlabel metal2 1293 6093 1307 6107 0 _2289_.A
rlabel metal2 1273 6113 1287 6127 0 _2289_.B
rlabel metal2 1233 6113 1247 6127 0 _2289_.C
rlabel metal2 1253 6093 1267 6107 0 _2289_.Y
rlabel metal1 1124 6002 1216 6018 0 _2285_.gnd
rlabel metal1 1124 6242 1216 6258 0 _2285_.vdd
rlabel metal2 1173 6093 1187 6107 0 _2285_.B
rlabel metal2 1133 6093 1147 6107 0 _2285_.A
rlabel metal2 1153 6073 1167 6087 0 _2285_.Y
rlabel metal1 1304 6002 1376 6018 0 _2288_.gnd
rlabel metal1 1304 6242 1376 6258 0 _2288_.vdd
rlabel metal2 1353 6073 1367 6087 0 _2288_.A
rlabel metal2 1333 6113 1347 6127 0 _2288_.Y
rlabel metal1 1424 6482 1536 6498 0 _2120_.gnd
rlabel metal1 1424 6242 1536 6258 0 _2120_.vdd
rlabel metal2 1513 6393 1527 6407 0 _2120_.A
rlabel metal2 1493 6373 1507 6387 0 _2120_.B
rlabel metal2 1453 6373 1467 6387 0 _2120_.C
rlabel metal2 1473 6393 1487 6407 0 _2120_.Y
rlabel metal1 1424 6002 1516 6018 0 _2279_.gnd
rlabel metal1 1424 6242 1516 6258 0 _2279_.vdd
rlabel metal2 1473 6093 1487 6107 0 _2279_.B
rlabel metal2 1433 6093 1447 6107 0 _2279_.A
rlabel metal2 1453 6073 1467 6087 0 _2279_.Y
rlabel metal1 1504 6002 1596 6018 0 _2278_.gnd
rlabel metal1 1504 6242 1596 6258 0 _2278_.vdd
rlabel metal2 1553 6093 1567 6107 0 _2278_.B
rlabel metal2 1513 6093 1527 6107 0 _2278_.A
rlabel metal2 1533 6073 1547 6087 0 _2278_.Y
rlabel metal1 1364 6002 1436 6018 0 _2280_.gnd
rlabel metal1 1364 6242 1436 6258 0 _2280_.vdd
rlabel metal2 1413 6073 1427 6087 0 _2280_.A
rlabel metal2 1393 6113 1407 6127 0 _2280_.Y
rlabel metal1 1584 6002 1656 6018 0 _2276_.gnd
rlabel metal1 1584 6242 1656 6258 0 _2276_.vdd
rlabel metal2 1593 6073 1607 6087 0 _2276_.A
rlabel metal2 1613 6113 1627 6127 0 _2276_.Y
rlabel metal1 1524 6482 1636 6498 0 _2119_.gnd
rlabel metal1 1524 6242 1636 6258 0 _2119_.vdd
rlabel metal2 1613 6393 1627 6407 0 _2119_.A
rlabel metal2 1553 6393 1567 6407 0 _2119_.Y
rlabel metal2 1573 6353 1587 6367 0 _2119_.B
rlabel metal1 1684 6482 1936 6498 0 _2375_.gnd
rlabel metal1 1684 6242 1936 6258 0 _2375_.vdd
rlabel metal2 1833 6393 1847 6407 0 _2375_.D
rlabel metal2 1793 6393 1807 6407 0 _2375_.CLK
rlabel metal2 1713 6393 1727 6407 0 _2375_.Q
rlabel metal1 1804 6002 1916 6018 0 _2124_.gnd
rlabel metal1 1804 6242 1916 6258 0 _2124_.vdd
rlabel metal2 1813 6093 1827 6107 0 _2124_.A
rlabel metal2 1833 6113 1847 6127 0 _2124_.B
rlabel metal2 1873 6113 1887 6127 0 _2124_.C
rlabel metal2 1853 6093 1867 6107 0 _2124_.Y
rlabel metal1 1644 6002 1736 6018 0 _2277_.gnd
rlabel metal1 1644 6242 1736 6258 0 _2277_.vdd
rlabel metal2 1693 6093 1707 6107 0 _2277_.B
rlabel metal2 1653 6093 1667 6107 0 _2277_.A
rlabel metal2 1673 6073 1687 6087 0 _2277_.Y
rlabel metal1 1724 6002 1816 6018 0 _2094_.gnd
rlabel metal1 1724 6242 1816 6258 0 _2094_.vdd
rlabel metal2 1773 6093 1787 6107 0 _2094_.B
rlabel metal2 1733 6093 1747 6107 0 _2094_.A
rlabel metal2 1753 6073 1767 6087 0 _2094_.Y
rlabel metal1 1624 6482 1696 6498 0 _2043_.gnd
rlabel metal1 1624 6242 1696 6258 0 _2043_.vdd
rlabel metal2 1673 6413 1687 6427 0 _2043_.A
rlabel metal2 1653 6373 1667 6387 0 _2043_.Y
rlabel metal1 1924 6482 2036 6498 0 _2089_.gnd
rlabel metal1 1924 6242 2036 6258 0 _2089_.vdd
rlabel metal2 1933 6393 1947 6407 0 _2089_.A
rlabel metal2 1953 6373 1967 6387 0 _2089_.B
rlabel metal2 1993 6373 2007 6387 0 _2089_.C
rlabel metal2 1973 6393 1987 6407 0 _2089_.Y
rlabel metal1 2104 6482 2216 6498 0 _2088_.gnd
rlabel metal1 2104 6242 2216 6258 0 _2088_.vdd
rlabel metal2 2193 6393 2207 6407 0 _2088_.A
rlabel metal2 2173 6373 2187 6387 0 _2088_.B
rlabel metal2 2133 6373 2147 6387 0 _2088_.C
rlabel metal2 2153 6393 2167 6407 0 _2088_.Y
rlabel metal1 2124 6002 2236 6018 0 _2040_.gnd
rlabel metal1 2124 6242 2236 6258 0 _2040_.vdd
rlabel metal2 2213 6093 2227 6107 0 _2040_.A
rlabel metal2 2193 6113 2207 6127 0 _2040_.B
rlabel metal2 2153 6113 2167 6127 0 _2040_.C
rlabel metal2 2173 6093 2187 6107 0 _2040_.Y
rlabel metal1 1904 6002 1976 6018 0 _2123_.gnd
rlabel metal1 1904 6242 1976 6258 0 _2123_.vdd
rlabel metal2 1913 6073 1927 6087 0 _2123_.A
rlabel metal2 1933 6113 1947 6127 0 _2123_.Y
rlabel metal1 2064 6002 2136 6018 0 _2036_.gnd
rlabel metal1 2064 6242 2136 6258 0 _2036_.vdd
rlabel metal2 2073 6073 2087 6087 0 _2036_.A
rlabel metal2 2093 6113 2107 6127 0 _2036_.Y
rlabel metal1 2024 6482 2116 6498 0 _2041_.gnd
rlabel metal1 2024 6242 2116 6258 0 _2041_.vdd
rlabel metal2 2033 6353 2047 6367 0 _2041_.A
rlabel metal2 2073 6353 2087 6367 0 _2041_.B
rlabel metal2 2053 6373 2067 6387 0 _2041_.Y
rlabel metal1 1964 6002 2076 6018 0 _2092_.gnd
rlabel metal1 1964 6242 2076 6258 0 _2092_.vdd
rlabel metal2 2053 6113 2067 6127 0 _2092_.A
rlabel metal2 2033 6073 2047 6087 0 _2092_.B
rlabel metal2 2013 6113 2027 6127 0 _2092_.C
rlabel metal2 1993 6093 2007 6107 0 _2092_.Y
rlabel metal1 2284 6002 2396 6018 0 _2093_.gnd
rlabel metal1 2284 6242 2396 6258 0 _2093_.vdd
rlabel metal2 2373 6093 2387 6107 0 _2093_.A
rlabel metal2 2353 6113 2367 6127 0 _2093_.B
rlabel metal2 2313 6113 2327 6127 0 _2093_.C
rlabel metal2 2333 6093 2347 6107 0 _2093_.Y
rlabel metal1 2384 6482 2476 6498 0 _2087_.gnd
rlabel metal1 2384 6242 2476 6258 0 _2087_.vdd
rlabel metal2 2413 6393 2427 6407 0 _2087_.B
rlabel metal2 2453 6393 2467 6407 0 _2087_.A
rlabel metal2 2433 6413 2447 6427 0 _2087_.Y
rlabel metal1 2224 6002 2296 6018 0 _2038_.gnd
rlabel metal1 2224 6242 2296 6258 0 _2038_.vdd
rlabel metal2 2233 6073 2247 6087 0 _2038_.A
rlabel metal2 2253 6113 2267 6127 0 _2038_.Y
rlabel metal1 2304 6482 2396 6498 0 _2082_.gnd
rlabel metal1 2304 6242 2396 6258 0 _2082_.vdd
rlabel metal2 2373 6353 2387 6367 0 _2082_.A
rlabel metal2 2333 6353 2347 6367 0 _2082_.B
rlabel metal2 2353 6373 2367 6387 0 _2082_.Y
rlabel metal1 2204 6482 2316 6498 0 _2081_.gnd
rlabel metal1 2204 6242 2316 6258 0 _2081_.vdd
rlabel metal2 2293 6373 2307 6387 0 _2081_.A
rlabel metal2 2273 6413 2287 6427 0 _2081_.B
rlabel metal2 2253 6373 2267 6387 0 _2081_.C
rlabel metal2 2233 6393 2247 6407 0 _2081_.Y
rlabel metal1 2384 6002 2496 6018 0 _2083_.gnd
rlabel metal1 2384 6242 2496 6258 0 _2083_.vdd
rlabel metal2 2473 6113 2487 6127 0 _2083_.A
rlabel metal2 2453 6133 2467 6147 0 _2083_.B
rlabel metal2 2433 6113 2447 6127 0 _2083_.C
rlabel metal2 2413 6133 2427 6147 0 _2083_.Y
rlabel metal1 2464 6482 2556 6498 0 _2142_.gnd
rlabel metal1 2464 6242 2556 6258 0 _2142_.vdd
rlabel metal2 2513 6393 2527 6407 0 _2142_.B
rlabel metal2 2473 6393 2487 6407 0 _2142_.A
rlabel metal2 2493 6413 2507 6427 0 _2142_.Y
rlabel metal1 2584 6002 2676 6018 0 _2080_.gnd
rlabel metal1 2584 6242 2676 6258 0 _2080_.vdd
rlabel metal2 2613 6093 2627 6107 0 _2080_.B
rlabel metal2 2653 6093 2667 6107 0 _2080_.A
rlabel metal2 2633 6073 2647 6087 0 _2080_.Y
rlabel metal1 2544 6482 2636 6498 0 _2086_.gnd
rlabel metal1 2544 6242 2636 6258 0 _2086_.vdd
rlabel metal2 2553 6353 2567 6367 0 _2086_.A
rlabel metal2 2593 6353 2607 6367 0 _2086_.B
rlabel metal2 2573 6373 2587 6387 0 _2086_.Y
rlabel metal1 2484 6002 2596 6018 0 _2079_.gnd
rlabel metal1 2484 6242 2596 6258 0 _2079_.vdd
rlabel metal2 2573 6113 2587 6127 0 _2079_.A
rlabel metal2 2553 6073 2567 6087 0 _2079_.B
rlabel metal2 2533 6113 2547 6127 0 _2079_.C
rlabel metal2 2513 6093 2527 6107 0 _2079_.Y
rlabel metal1 2624 6482 2736 6498 0 _2091_.gnd
rlabel metal1 2624 6242 2736 6258 0 _2091_.vdd
rlabel metal2 2713 6373 2727 6387 0 _2091_.A
rlabel metal2 2693 6353 2707 6367 0 _2091_.B
rlabel metal2 2673 6373 2687 6387 0 _2091_.C
rlabel metal2 2653 6353 2667 6367 0 _2091_.Y
rlabel metal1 2664 6002 2776 6018 0 _2085_.gnd
rlabel metal1 2664 6242 2776 6258 0 _2085_.vdd
rlabel metal2 2753 6113 2767 6127 0 _2085_.A
rlabel metal2 2733 6133 2747 6147 0 _2085_.B
rlabel metal2 2713 6113 2727 6127 0 _2085_.C
rlabel metal2 2693 6133 2707 6147 0 _2085_.Y
rlabel metal1 2904 6482 3016 6498 0 _2076_.gnd
rlabel metal1 2904 6242 3016 6258 0 _2076_.vdd
rlabel metal2 2993 6393 3007 6407 0 _2076_.A
rlabel metal2 2973 6373 2987 6387 0 _2076_.B
rlabel metal2 2933 6373 2947 6387 0 _2076_.C
rlabel metal2 2953 6393 2967 6407 0 _2076_.Y
rlabel metal1 2884 6002 2956 6018 0 _2071_.gnd
rlabel metal1 2884 6242 2956 6258 0 _2071_.vdd
rlabel metal2 2933 6073 2947 6087 0 _2071_.A
rlabel metal2 2913 6113 2927 6127 0 _2071_.Y
rlabel metal1 2724 6482 2816 6498 0 _2035_.gnd
rlabel metal1 2724 6242 2816 6258 0 _2035_.vdd
rlabel metal2 2733 6353 2747 6367 0 _2035_.A
rlabel metal2 2773 6353 2787 6367 0 _2035_.B
rlabel metal2 2753 6373 2767 6387 0 _2035_.Y
rlabel metal1 2804 6482 2916 6498 0 _2034_.gnd
rlabel metal1 2804 6242 2916 6258 0 _2034_.vdd
rlabel metal2 2893 6373 2907 6387 0 _2034_.A
rlabel metal2 2873 6353 2887 6367 0 _2034_.B
rlabel metal2 2853 6373 2867 6387 0 _2034_.C
rlabel metal2 2833 6353 2847 6367 0 _2034_.Y
rlabel metal1 2764 6002 2896 6018 0 _2075_.gnd
rlabel metal1 2764 6242 2896 6258 0 _2075_.vdd
rlabel metal2 2873 6093 2887 6107 0 _2075_.A
rlabel metal2 2853 6113 2867 6127 0 _2075_.B
rlabel metal2 2793 6093 2807 6107 0 _2075_.C
rlabel metal2 2813 6113 2827 6127 0 _2075_.D
rlabel metal2 2833 6093 2847 6107 0 _2075_.Y
rlabel metal1 3004 6482 3116 6498 0 _2033_.gnd
rlabel metal1 3004 6242 3116 6258 0 _2033_.vdd
rlabel metal2 3093 6393 3107 6407 0 _2033_.A
rlabel metal2 3073 6373 3087 6387 0 _2033_.B
rlabel metal2 3033 6373 3047 6387 0 _2033_.C
rlabel metal2 3053 6393 3067 6407 0 _2033_.Y
rlabel metal1 3104 6482 3176 6498 0 _2031_.gnd
rlabel metal1 3104 6242 3176 6258 0 _2031_.vdd
rlabel metal2 3153 6413 3167 6427 0 _2031_.A
rlabel metal2 3133 6373 3147 6387 0 _2031_.Y
rlabel metal1 3164 6482 3236 6498 0 _1989_.gnd
rlabel metal1 3164 6242 3236 6258 0 _1989_.vdd
rlabel metal2 3213 6413 3227 6427 0 _1989_.A
rlabel metal2 3193 6373 3207 6387 0 _1989_.Y
rlabel metal1 3044 6002 3156 6018 0 _2084_.gnd
rlabel metal1 3044 6242 3156 6258 0 _2084_.vdd
rlabel metal2 3133 6113 3147 6127 0 _2084_.A
rlabel metal2 3113 6073 3127 6087 0 _2084_.B
rlabel metal2 3093 6113 3107 6127 0 _2084_.C
rlabel metal2 3073 6093 3087 6107 0 _2084_.Y
rlabel metal1 2944 6002 3056 6018 0 _2074_.gnd
rlabel metal1 2944 6242 3056 6258 0 _2074_.vdd
rlabel metal2 2953 6113 2967 6127 0 _2074_.A
rlabel metal2 2973 6133 2987 6147 0 _2074_.B
rlabel metal2 2993 6113 3007 6127 0 _2074_.C
rlabel metal2 3013 6133 3027 6147 0 _2074_.Y
rlabel metal1 3144 6002 3256 6018 0 _2030_.gnd
rlabel metal1 3144 6242 3256 6258 0 _2030_.vdd
rlabel metal2 3233 6113 3247 6127 0 _2030_.A
rlabel metal2 3213 6133 3227 6147 0 _2030_.B
rlabel metal2 3193 6113 3207 6127 0 _2030_.C
rlabel metal2 3173 6133 3187 6147 0 _2030_.Y
rlabel metal1 3324 6482 3436 6498 0 _2028_.gnd
rlabel metal1 3324 6242 3436 6258 0 _2028_.vdd
rlabel metal2 3333 6393 3347 6407 0 _2028_.A
rlabel metal2 3353 6373 3367 6387 0 _2028_.B
rlabel metal2 3393 6373 3407 6387 0 _2028_.C
rlabel metal2 3373 6393 3387 6407 0 _2028_.Y
rlabel metal1 3344 6002 3416 6018 0 _2065_.gnd
rlabel metal1 3344 6242 3416 6258 0 _2065_.vdd
rlabel metal2 3393 6073 3407 6087 0 _2065_.A
rlabel metal2 3373 6113 3387 6127 0 _2065_.Y
rlabel metal1 3244 6002 3356 6018 0 _2066_.gnd
rlabel metal1 3244 6242 3356 6258 0 _2066_.vdd
rlabel metal2 3333 6113 3347 6127 0 _2066_.A
rlabel metal2 3313 6073 3327 6087 0 _2066_.B
rlabel metal2 3293 6113 3307 6127 0 _2066_.C
rlabel metal2 3273 6093 3287 6107 0 _2066_.Y
rlabel metal1 3424 6482 3536 6498 0 _2032_.gnd
rlabel metal1 3424 6242 3536 6258 0 _2032_.vdd
rlabel metal2 3513 6373 3527 6387 0 _2032_.A
rlabel metal2 3493 6413 3507 6427 0 _2032_.B
rlabel metal2 3473 6373 3487 6387 0 _2032_.C
rlabel metal2 3453 6393 3467 6407 0 _2032_.Y
rlabel metal1 3224 6482 3336 6498 0 _2027_.gnd
rlabel metal1 3224 6242 3336 6258 0 _2027_.vdd
rlabel metal2 3233 6373 3247 6387 0 _2027_.A
rlabel metal2 3253 6413 3267 6427 0 _2027_.B
rlabel metal2 3273 6373 3287 6387 0 _2027_.C
rlabel metal2 3293 6393 3307 6407 0 _2027_.Y
rlabel metal1 3404 6002 3516 6018 0 _2025_.gnd
rlabel metal1 3404 6242 3516 6258 0 _2025_.vdd
rlabel metal2 3493 6113 3507 6127 0 _2025_.A
rlabel metal2 3473 6133 3487 6147 0 _2025_.B
rlabel metal2 3453 6113 3467 6127 0 _2025_.C
rlabel metal2 3433 6133 3447 6147 0 _2025_.Y
rlabel metal1 3724 6482 3836 6498 0 _2026_.gnd
rlabel metal1 3724 6242 3836 6258 0 _2026_.vdd
rlabel metal2 3813 6393 3827 6407 0 _2026_.A
rlabel metal2 3793 6373 3807 6387 0 _2026_.B
rlabel metal2 3753 6373 3767 6387 0 _2026_.C
rlabel metal2 3773 6393 3787 6407 0 _2026_.Y
rlabel metal1 3604 6002 3676 6018 0 _2015_.gnd
rlabel metal1 3604 6242 3676 6258 0 _2015_.vdd
rlabel metal2 3613 6073 3627 6087 0 _2015_.A
rlabel metal2 3633 6113 3647 6127 0 _2015_.Y
rlabel metal1 3524 6482 3636 6498 0 _2024_.gnd
rlabel metal1 3524 6242 3636 6258 0 _2024_.vdd
rlabel metal2 3613 6373 3627 6387 0 _2024_.A
rlabel metal2 3593 6413 3607 6427 0 _2024_.B
rlabel metal2 3573 6373 3587 6387 0 _2024_.C
rlabel metal2 3553 6393 3567 6407 0 _2024_.Y
rlabel metal1 3664 6002 3776 6018 0 _2018_.gnd
rlabel metal1 3664 6242 3776 6258 0 _2018_.vdd
rlabel metal2 3673 6113 3687 6127 0 _2018_.A
rlabel metal2 3693 6073 3707 6087 0 _2018_.B
rlabel metal2 3713 6113 3727 6127 0 _2018_.C
rlabel metal2 3733 6093 3747 6107 0 _2018_.Y
rlabel metal1 3624 6482 3736 6498 0 _2023_.gnd
rlabel metal1 3624 6242 3736 6258 0 _2023_.vdd
rlabel metal2 3633 6373 3647 6387 0 _2023_.A
rlabel metal2 3653 6353 3667 6367 0 _2023_.B
rlabel metal2 3673 6373 3687 6387 0 _2023_.C
rlabel metal2 3693 6353 3707 6367 0 _2023_.Y
rlabel metal1 3504 6002 3616 6018 0 _2021_.gnd
rlabel metal1 3504 6242 3616 6258 0 _2021_.vdd
rlabel metal2 3513 6113 3527 6127 0 _2021_.A
rlabel metal2 3533 6133 3547 6147 0 _2021_.B
rlabel metal2 3553 6113 3567 6127 0 _2021_.C
rlabel metal2 3573 6133 3587 6147 0 _2021_.Y
rlabel metal1 3824 6482 3936 6498 0 _2019_.gnd
rlabel metal1 3824 6242 3936 6258 0 _2019_.vdd
rlabel metal2 3833 6393 3847 6407 0 _2019_.A
rlabel metal2 3853 6373 3867 6387 0 _2019_.B
rlabel metal2 3893 6373 3907 6387 0 _2019_.C
rlabel metal2 3873 6393 3887 6407 0 _2019_.Y
rlabel metal1 3924 6002 4036 6018 0 _2008_.gnd
rlabel metal1 3924 6242 4036 6258 0 _2008_.vdd
rlabel metal2 4013 6093 4027 6107 0 _2008_.A
rlabel metal2 3993 6113 4007 6127 0 _2008_.B
rlabel metal2 3953 6113 3967 6127 0 _2008_.C
rlabel metal2 3973 6093 3987 6107 0 _2008_.Y
rlabel metal1 3924 6482 3996 6498 0 _2020_.gnd
rlabel metal1 3924 6242 3996 6258 0 _2020_.vdd
rlabel metal2 3933 6413 3947 6427 0 _2020_.A
rlabel metal2 3953 6373 3967 6387 0 _2020_.Y
rlabel metal1 3764 6002 3856 6018 0 _1983_.gnd
rlabel metal1 3764 6242 3856 6258 0 _1983_.vdd
rlabel metal2 3833 6133 3847 6147 0 _1983_.A
rlabel metal2 3793 6133 3807 6147 0 _1983_.B
rlabel metal2 3813 6113 3827 6127 0 _1983_.Y
rlabel metal1 3844 6002 3936 6018 0 _1982_.gnd
rlabel metal1 3844 6242 3936 6258 0 _1982_.vdd
rlabel metal2 3853 6133 3867 6147 0 _1982_.A
rlabel metal2 3893 6133 3907 6147 0 _1982_.B
rlabel metal2 3873 6113 3887 6127 0 _1982_.Y
rlabel metal1 3984 6482 4076 6498 0 _1977_.gnd
rlabel metal1 3984 6242 4076 6258 0 _1977_.vdd
rlabel metal2 3993 6353 4007 6367 0 _1977_.A
rlabel metal2 4033 6353 4047 6367 0 _1977_.B
rlabel metal2 4013 6373 4027 6387 0 _1977_.Y
rlabel metal1 4024 6002 4136 6018 0 _2017_.gnd
rlabel metal1 4024 6242 4136 6258 0 _2017_.vdd
rlabel metal2 4033 6093 4047 6107 0 _2017_.A
rlabel metal2 4053 6113 4067 6127 0 _2017_.B
rlabel metal2 4093 6113 4107 6127 0 _2017_.C
rlabel metal2 4073 6093 4087 6107 0 _2017_.Y
rlabel metal1 4124 6002 4216 6018 0 _2004_.gnd
rlabel metal1 4124 6242 4216 6258 0 _2004_.vdd
rlabel metal2 4153 6093 4167 6107 0 _2004_.B
rlabel metal2 4193 6093 4207 6107 0 _2004_.A
rlabel metal2 4173 6073 4187 6087 0 _2004_.Y
rlabel metal1 4204 6002 4276 6018 0 _1999_.gnd
rlabel metal1 4204 6242 4276 6258 0 _1999_.vdd
rlabel metal2 4213 6073 4227 6087 0 _1999_.A
rlabel metal2 4233 6113 4247 6127 0 _1999_.Y
rlabel metal1 4164 6482 4256 6498 0 _2029_.gnd
rlabel metal1 4164 6242 4256 6258 0 _2029_.vdd
rlabel metal2 4173 6353 4187 6367 0 _2029_.A
rlabel metal2 4213 6353 4227 6367 0 _2029_.B
rlabel metal2 4193 6373 4207 6387 0 _2029_.Y
rlabel metal1 4264 6002 4356 6018 0 _1937_.gnd
rlabel metal1 4264 6242 4356 6258 0 _1937_.vdd
rlabel metal2 4333 6133 4347 6147 0 _1937_.A
rlabel metal2 4293 6133 4307 6147 0 _1937_.B
rlabel metal2 4313 6113 4327 6127 0 _1937_.Y
rlabel metal1 4244 6482 4356 6498 0 _1976_.gnd
rlabel metal1 4244 6242 4356 6258 0 _1976_.vdd
rlabel metal2 4333 6373 4347 6387 0 _1976_.A
rlabel metal2 4313 6353 4327 6367 0 _1976_.B
rlabel metal2 4293 6373 4307 6387 0 _1976_.C
rlabel metal2 4273 6353 4287 6367 0 _1976_.Y
rlabel metal1 4064 6482 4176 6498 0 _1987_.gnd
rlabel metal1 4064 6242 4176 6258 0 _1987_.vdd
rlabel metal2 4153 6393 4167 6407 0 _1987_.A
rlabel metal2 4093 6393 4107 6407 0 _1987_.Y
rlabel metal2 4113 6353 4127 6367 0 _1987_.B
rlabel metal1 4444 6002 4556 6018 0 _1991_.gnd
rlabel metal1 4444 6242 4556 6258 0 _1991_.vdd
rlabel metal2 4533 6093 4547 6107 0 _1991_.A
rlabel metal2 4513 6113 4527 6127 0 _1991_.B
rlabel metal2 4473 6113 4487 6127 0 _1991_.C
rlabel metal2 4493 6093 4507 6107 0 _1991_.Y
rlabel metal1 4444 6482 4556 6498 0 _1975_.gnd
rlabel metal1 4444 6242 4556 6258 0 _1975_.vdd
rlabel metal2 4533 6373 4547 6387 0 _1975_.A
rlabel metal2 4513 6353 4527 6367 0 _1975_.B
rlabel metal2 4493 6373 4507 6387 0 _1975_.C
rlabel metal2 4473 6353 4487 6367 0 _1975_.Y
rlabel metal1 4344 6482 4456 6498 0 _1974_.gnd
rlabel metal1 4344 6242 4456 6258 0 _1974_.vdd
rlabel metal2 4433 6373 4447 6387 0 _1974_.A
rlabel metal2 4413 6353 4427 6367 0 _1974_.B
rlabel metal2 4393 6373 4407 6387 0 _1974_.C
rlabel metal2 4373 6353 4387 6367 0 _1974_.Y
rlabel metal1 4344 6002 4456 6018 0 _1957_.gnd
rlabel metal1 4344 6242 4456 6258 0 _1957_.vdd
rlabel metal2 4353 6093 4367 6107 0 _1957_.A
rlabel metal2 4413 6093 4427 6107 0 _1957_.Y
rlabel metal2 4393 6133 4407 6147 0 _1957_.B
rlabel metal1 4804 6482 4916 6498 0 _1971_.gnd
rlabel metal1 4804 6242 4916 6258 0 _1971_.vdd
rlabel metal2 4813 6393 4827 6407 0 _1971_.A
rlabel metal2 4833 6373 4847 6387 0 _1971_.B
rlabel metal2 4873 6373 4887 6387 0 _1971_.C
rlabel metal2 4853 6393 4867 6407 0 _1971_.Y
rlabel metal1 4544 6482 4616 6498 0 _1924_.gnd
rlabel metal1 4544 6242 4616 6258 0 _1924_.vdd
rlabel metal2 4553 6413 4567 6427 0 _1924_.A
rlabel metal2 4573 6373 4587 6387 0 _1924_.Y
rlabel metal1 4744 6002 4856 6018 0 _1990_.gnd
rlabel metal1 4744 6242 4856 6258 0 _1990_.vdd
rlabel metal2 4833 6113 4847 6127 0 _1990_.A
rlabel metal2 4813 6073 4827 6087 0 _1990_.B
rlabel metal2 4793 6113 4807 6127 0 _1990_.C
rlabel metal2 4773 6093 4787 6107 0 _1990_.Y
rlabel metal1 4704 6482 4816 6498 0 _1970_.gnd
rlabel metal1 4704 6242 4816 6258 0 _1970_.vdd
rlabel metal2 4713 6373 4727 6387 0 _1970_.A
rlabel metal2 4733 6413 4747 6427 0 _1970_.B
rlabel metal2 4753 6373 4767 6387 0 _1970_.C
rlabel metal2 4773 6393 4787 6407 0 _1970_.Y
rlabel metal1 4604 6482 4716 6498 0 _1967_.gnd
rlabel metal1 4604 6242 4716 6258 0 _1967_.vdd
rlabel metal2 4613 6373 4627 6387 0 _1967_.A
rlabel metal2 4633 6413 4647 6427 0 _1967_.B
rlabel metal2 4653 6373 4667 6387 0 _1967_.C
rlabel metal2 4673 6393 4687 6407 0 _1967_.Y
rlabel metal1 4544 6002 4656 6018 0 _1960_.gnd
rlabel metal1 4544 6242 4656 6258 0 _1960_.vdd
rlabel metal2 4633 6113 4647 6127 0 _1960_.A
rlabel metal2 4613 6073 4627 6087 0 _1960_.B
rlabel metal2 4593 6113 4607 6127 0 _1960_.C
rlabel metal2 4573 6093 4587 6107 0 _1960_.Y
rlabel metal1 4644 6002 4756 6018 0 _1964_.gnd
rlabel metal1 4644 6242 4756 6258 0 _1964_.vdd
rlabel metal2 4653 6113 4667 6127 0 _1964_.A
rlabel metal2 4673 6133 4687 6147 0 _1964_.B
rlabel metal2 4693 6113 4707 6127 0 _1964_.C
rlabel metal2 4713 6133 4727 6147 0 _1964_.Y
rlabel metal1 4904 6482 5016 6498 0 _1969_.gnd
rlabel metal1 4904 6242 5016 6258 0 _1969_.vdd
rlabel metal2 4993 6393 5007 6407 0 _1969_.A
rlabel metal2 4973 6373 4987 6387 0 _1969_.B
rlabel metal2 4933 6373 4947 6387 0 _1969_.C
rlabel metal2 4953 6393 4967 6407 0 _1969_.Y
rlabel metal1 5004 6482 5116 6498 0 _1961_.gnd
rlabel metal1 5004 6242 5116 6258 0 _1961_.vdd
rlabel metal2 5013 6393 5027 6407 0 _1961_.A
rlabel metal2 5033 6373 5047 6387 0 _1961_.B
rlabel metal2 5073 6373 5087 6387 0 _1961_.C
rlabel metal2 5053 6393 5067 6407 0 _1961_.Y
rlabel metal1 5044 6002 5156 6018 0 _1951_.gnd
rlabel metal1 5044 6242 5156 6258 0 _1951_.vdd
rlabel metal2 5133 6093 5147 6107 0 _1951_.A
rlabel metal2 5113 6113 5127 6127 0 _1951_.B
rlabel metal2 5073 6113 5087 6127 0 _1951_.C
rlabel metal2 5093 6093 5107 6107 0 _1951_.Y
rlabel metal1 4844 6002 4956 6018 0 _1958_.gnd
rlabel metal1 4844 6242 4956 6258 0 _1958_.vdd
rlabel metal2 4933 6113 4947 6127 0 _1958_.A
rlabel metal2 4913 6133 4927 6147 0 _1958_.B
rlabel metal2 4893 6113 4907 6127 0 _1958_.C
rlabel metal2 4873 6133 4887 6147 0 _1958_.Y
rlabel metal1 4944 6002 5056 6018 0 _1955_.gnd
rlabel metal1 4944 6242 5056 6258 0 _1955_.vdd
rlabel metal2 4953 6113 4967 6127 0 _1955_.A
rlabel metal2 4973 6133 4987 6147 0 _1955_.B
rlabel metal2 4993 6113 5007 6127 0 _1955_.C
rlabel metal2 5013 6133 5027 6147 0 _1955_.Y
rlabel metal1 5324 6002 5436 6018 0 _1926_.gnd
rlabel metal1 5324 6242 5436 6258 0 _1926_.vdd
rlabel metal2 5333 6093 5347 6107 0 _1926_.A
rlabel metal2 5353 6113 5367 6127 0 _1926_.B
rlabel metal2 5393 6113 5407 6127 0 _1926_.C
rlabel metal2 5373 6093 5387 6107 0 _1926_.Y
rlabel metal1 5144 6002 5236 6018 0 _1869_.gnd
rlabel metal1 5144 6242 5236 6258 0 _1869_.vdd
rlabel metal2 5213 6133 5227 6147 0 _1869_.A
rlabel metal2 5173 6133 5187 6147 0 _1869_.B
rlabel metal2 5193 6113 5207 6127 0 _1869_.Y
rlabel metal1 5204 6482 5316 6498 0 _1968_.gnd
rlabel metal1 5204 6242 5316 6258 0 _1968_.vdd
rlabel metal2 5293 6373 5307 6387 0 _1968_.A
rlabel metal2 5273 6353 5287 6367 0 _1968_.B
rlabel metal2 5253 6373 5267 6387 0 _1968_.C
rlabel metal2 5233 6353 5247 6367 0 _1968_.Y
rlabel metal1 5104 6482 5216 6498 0 _1966_.gnd
rlabel metal1 5104 6242 5216 6258 0 _1966_.vdd
rlabel metal2 5193 6373 5207 6387 0 _1966_.A
rlabel metal2 5173 6353 5187 6367 0 _1966_.B
rlabel metal2 5153 6373 5167 6387 0 _1966_.C
rlabel metal2 5133 6353 5147 6367 0 _1966_.Y
rlabel metal1 5304 6482 5416 6498 0 _1965_.gnd
rlabel metal1 5304 6242 5416 6258 0 _1965_.vdd
rlabel metal2 5393 6373 5407 6387 0 _1965_.A
rlabel metal2 5373 6353 5387 6367 0 _1965_.B
rlabel metal2 5353 6373 5367 6387 0 _1965_.C
rlabel metal2 5333 6353 5347 6367 0 _1965_.Y
rlabel metal1 5224 6002 5336 6018 0 _1888_.gnd
rlabel metal1 5224 6242 5336 6258 0 _1888_.vdd
rlabel metal2 5233 6093 5247 6107 0 _1888_.A
rlabel metal2 5293 6093 5307 6107 0 _1888_.Y
rlabel metal2 5273 6133 5287 6147 0 _1888_.B
rlabel metal1 5604 6482 5676 6498 0 _1962_.gnd
rlabel metal1 5604 6242 5676 6258 0 _1962_.vdd
rlabel metal2 5653 6413 5667 6427 0 _1962_.A
rlabel metal2 5633 6373 5647 6387 0 _1962_.Y
rlabel metal1 5504 6482 5616 6498 0 _1963_.gnd
rlabel metal1 5504 6242 5616 6258 0 _1963_.vdd
rlabel metal2 5593 6373 5607 6387 0 _1963_.A
rlabel metal2 5573 6413 5587 6427 0 _1963_.B
rlabel metal2 5553 6373 5567 6387 0 _1963_.C
rlabel metal2 5533 6393 5547 6407 0 _1963_.Y
rlabel metal1 5404 6482 5516 6498 0 _1956_.gnd
rlabel metal1 5404 6242 5516 6258 0 _1956_.vdd
rlabel metal2 5413 6373 5427 6387 0 _1956_.A
rlabel metal2 5433 6413 5447 6427 0 _1956_.B
rlabel metal2 5453 6373 5467 6387 0 _1956_.C
rlabel metal2 5473 6393 5487 6407 0 _1956_.Y
rlabel metal1 5424 6002 5536 6018 0 _1925_.gnd
rlabel metal1 5424 6242 5536 6258 0 _1925_.vdd
rlabel metal2 5513 6113 5527 6127 0 _1925_.A
rlabel metal2 5493 6073 5507 6087 0 _1925_.B
rlabel metal2 5473 6113 5487 6127 0 _1925_.C
rlabel metal2 5453 6093 5467 6107 0 _1925_.Y
rlabel metal1 5524 6002 5636 6018 0 _1889_.gnd
rlabel metal1 5524 6242 5636 6258 0 _1889_.vdd
rlabel metal2 5613 6113 5627 6127 0 _1889_.A
rlabel metal2 5593 6133 5607 6147 0 _1889_.B
rlabel metal2 5573 6113 5587 6127 0 _1889_.C
rlabel metal2 5553 6133 5567 6147 0 _1889_.Y
rlabel metal1 5864 6482 5976 6498 0 _1920_.gnd
rlabel metal1 5864 6242 5976 6258 0 _1920_.vdd
rlabel metal2 5953 6373 5967 6387 0 _1920_.A
rlabel metal2 5933 6413 5947 6427 0 _1920_.B
rlabel metal2 5913 6373 5927 6387 0 _1920_.C
rlabel metal2 5893 6393 5907 6407 0 _1920_.Y
rlabel metal1 5664 6482 5776 6498 0 _1891_.gnd
rlabel metal1 5664 6242 5776 6258 0 _1891_.vdd
rlabel metal2 5673 6373 5687 6387 0 _1891_.A
rlabel metal2 5693 6413 5707 6427 0 _1891_.B
rlabel metal2 5713 6373 5727 6387 0 _1891_.C
rlabel metal2 5733 6393 5747 6407 0 _1891_.Y
rlabel metal1 5724 6002 5836 6018 0 _1887_.gnd
rlabel metal1 5724 6242 5836 6258 0 _1887_.vdd
rlabel metal2 5813 6113 5827 6127 0 _1887_.A
rlabel metal2 5793 6073 5807 6087 0 _1887_.B
rlabel metal2 5773 6113 5787 6127 0 _1887_.C
rlabel metal2 5753 6093 5767 6107 0 _1887_.Y
rlabel metal1 5824 6002 5936 6018 0 _1896_.gnd
rlabel metal1 5824 6242 5936 6258 0 _1896_.vdd
rlabel metal2 5833 6113 5847 6127 0 _1896_.A
rlabel metal2 5853 6133 5867 6147 0 _1896_.B
rlabel metal2 5873 6113 5887 6127 0 _1896_.C
rlabel metal2 5893 6133 5907 6147 0 _1896_.Y
rlabel metal1 5764 6482 5876 6498 0 _1895_.gnd
rlabel metal1 5764 6242 5876 6258 0 _1895_.vdd
rlabel metal2 5773 6373 5787 6387 0 _1895_.A
rlabel metal2 5793 6353 5807 6367 0 _1895_.B
rlabel metal2 5813 6373 5827 6387 0 _1895_.C
rlabel metal2 5833 6353 5847 6367 0 _1895_.Y
rlabel metal1 5624 6002 5736 6018 0 _1886_.gnd
rlabel metal1 5624 6242 5736 6258 0 _1886_.vdd
rlabel metal2 5633 6113 5647 6127 0 _1886_.A
rlabel metal2 5653 6133 5667 6147 0 _1886_.B
rlabel metal2 5673 6113 5687 6127 0 _1886_.C
rlabel metal2 5693 6133 5707 6147 0 _1886_.Y
rlabel metal1 6124 6482 6236 6498 0 _1973_.gnd
rlabel metal1 6124 6242 6236 6258 0 _1973_.vdd
rlabel metal2 6213 6393 6227 6407 0 _1973_.A
rlabel metal2 6193 6373 6207 6387 0 _1973_.B
rlabel metal2 6153 6373 6167 6387 0 _1973_.C
rlabel metal2 6173 6393 6187 6407 0 _1973_.Y
rlabel metal1 5924 6002 6036 6018 0 _1901_.gnd
rlabel metal1 5924 6242 6036 6258 0 _1901_.vdd
rlabel metal2 5933 6093 5947 6107 0 _1901_.A
rlabel metal2 5953 6113 5967 6127 0 _1901_.B
rlabel metal2 5993 6113 6007 6127 0 _1901_.C
rlabel metal2 5973 6093 5987 6107 0 _1901_.Y
rlabel metal1 6024 6002 6136 6018 0 _1892_.gnd
rlabel metal1 6024 6242 6136 6258 0 _1892_.vdd
rlabel metal2 6033 6093 6047 6107 0 _1892_.A
rlabel metal2 6053 6113 6067 6127 0 _1892_.B
rlabel metal2 6093 6113 6107 6127 0 _1892_.C
rlabel metal2 6073 6093 6087 6107 0 _1892_.Y
rlabel metal1 5964 6482 6036 6498 0 _1919_.gnd
rlabel metal1 5964 6242 6036 6258 0 _1919_.vdd
rlabel metal2 6013 6413 6027 6427 0 _1919_.A
rlabel metal2 5993 6373 6007 6387 0 _1919_.Y
rlabel metal1 6024 6482 6136 6498 0 _1902_.gnd
rlabel metal1 6024 6242 6136 6258 0 _1902_.vdd
rlabel metal2 6113 6373 6127 6387 0 _1902_.A
rlabel metal2 6093 6413 6107 6427 0 _1902_.B
rlabel metal2 6073 6373 6087 6387 0 _1902_.C
rlabel metal2 6053 6393 6067 6407 0 _1902_.Y
rlabel metal1 6124 6002 6236 6018 0 _1897_.gnd
rlabel metal1 6124 6242 6236 6258 0 _1897_.vdd
rlabel metal2 6133 6113 6147 6127 0 _1897_.A
rlabel metal2 6153 6133 6167 6147 0 _1897_.B
rlabel metal2 6173 6113 6187 6127 0 _1897_.C
rlabel metal2 6193 6133 6207 6147 0 _1897_.Y
rlabel metal1 6224 6482 6336 6498 0 _1972_.gnd
rlabel metal1 6224 6242 6336 6258 0 _1972_.vdd
rlabel metal2 6313 6373 6327 6387 0 _1972_.A
rlabel metal2 6293 6413 6307 6427 0 _1972_.B
rlabel metal2 6273 6373 6287 6387 0 _1972_.C
rlabel metal2 6253 6393 6267 6407 0 _1972_.Y
rlabel metal1 6324 6002 6436 6018 0 _1909_.gnd
rlabel metal1 6324 6242 6436 6258 0 _1909_.vdd
rlabel metal2 6413 6113 6427 6127 0 _1909_.A
rlabel metal2 6393 6133 6407 6147 0 _1909_.B
rlabel metal2 6373 6113 6387 6127 0 _1909_.C
rlabel metal2 6353 6133 6367 6147 0 _1909_.Y
rlabel metal1 6224 6002 6336 6018 0 _1908_.gnd
rlabel metal1 6224 6242 6336 6258 0 _1908_.vdd
rlabel metal2 6233 6113 6247 6127 0 _1908_.A
rlabel metal2 6253 6133 6267 6147 0 _1908_.B
rlabel metal2 6273 6113 6287 6127 0 _1908_.C
rlabel metal2 6293 6133 6307 6147 0 _1908_.Y
rlabel metal1 6324 6482 6436 6498 0 _1900_.gnd
rlabel metal1 6324 6242 6436 6258 0 _1900_.vdd
rlabel metal2 6333 6373 6347 6387 0 _1900_.A
rlabel metal2 6353 6353 6367 6367 0 _1900_.B
rlabel metal2 6373 6373 6387 6387 0 _1900_.C
rlabel metal2 6393 6353 6407 6367 0 _1900_.Y
rlabel nsubstratencontact 6676 6248 6676 6248 0 FILL100050x90150.vdd
rlabel metal1 6664 6002 6696 6018 0 FILL100050x90150.gnd
rlabel nsubstratencontact 6656 6248 6656 6248 0 FILL99750x90150.vdd
rlabel metal1 6644 6002 6676 6018 0 FILL99750x90150.gnd
rlabel metal1 6584 6002 6656 6018 0 _2581_.gnd
rlabel metal1 6584 6242 6656 6258 0 _2581_.vdd
rlabel metal2 6593 6073 6607 6087 0 _2581_.A
rlabel metal2 6613 6113 6627 6127 0 _2581_.Y
rlabel metal1 6524 6482 6596 6498 0 _1907_.gnd
rlabel metal1 6524 6242 6596 6258 0 _1907_.vdd
rlabel metal2 6533 6413 6547 6427 0 _1907_.A
rlabel metal2 6553 6373 6567 6387 0 _1907_.Y
rlabel metal1 6524 6002 6596 6018 0 _1893_.gnd
rlabel metal1 6524 6242 6596 6258 0 _1893_.vdd
rlabel metal2 6533 6073 6547 6087 0 _1893_.A
rlabel metal2 6553 6113 6567 6127 0 _1893_.Y
rlabel metal1 6424 6002 6536 6018 0 _1894_.gnd
rlabel metal1 6424 6242 6536 6258 0 _1894_.vdd
rlabel metal2 6513 6113 6527 6127 0 _1894_.A
rlabel metal2 6493 6073 6507 6087 0 _1894_.B
rlabel metal2 6473 6113 6487 6127 0 _1894_.C
rlabel metal2 6453 6093 6467 6107 0 _1894_.Y
rlabel metal1 6424 6482 6536 6498 0 _1906_.gnd
rlabel metal1 6424 6242 6536 6258 0 _1906_.vdd
rlabel metal2 6513 6373 6527 6387 0 _1906_.A
rlabel metal2 6493 6353 6507 6367 0 _1906_.B
rlabel metal2 6473 6373 6487 6387 0 _1906_.C
rlabel metal2 6453 6353 6467 6367 0 _1906_.Y
rlabel metal1 6584 6482 6716 6498 0 _2707_.gnd
rlabel metal1 6584 6242 6716 6258 0 _2707_.vdd
rlabel metal2 6593 6393 6607 6407 0 _2707_.A
rlabel metal2 6613 6373 6627 6387 0 _2707_.B
rlabel metal2 6673 6393 6687 6407 0 _2707_.C
rlabel metal2 6653 6373 6667 6387 0 _2707_.D
rlabel metal2 6633 6393 6647 6407 0 _2707_.Y
rlabel nsubstratencontact 6724 6252 6724 6252 0 FILL100650x93750.vdd
rlabel metal1 6704 6482 6736 6498 0 FILL100650x93750.gnd
rlabel nsubstratencontact 6716 6248 6716 6248 0 FILL100650x90150.vdd
rlabel metal1 6704 6002 6736 6018 0 FILL100650x90150.gnd
rlabel nsubstratencontact 6696 6248 6696 6248 0 FILL100350x90150.vdd
rlabel metal1 6684 6002 6716 6018 0 FILL100350x90150.gnd
<< end >>
