magic
tech scmos
magscale 1 2
timestamp 1726480912
<< nwell >>
rect -14 154 132 272
<< ntransistor >>
rect 22 14 26 54
rect 32 14 36 54
rect 52 14 56 54
rect 62 14 66 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 32 54
rect 36 14 38 54
rect 50 14 52 54
rect 56 14 62 54
rect 66 14 68 54
<< pdiffusion >>
rect 18 168 20 246
rect 6 166 20 168
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 168 46 246
rect 58 168 60 246
rect 44 166 60 168
rect 64 234 80 246
rect 64 166 66 234
rect 78 166 80 234
rect 84 166 86 246
<< ndcontact >>
rect 8 14 20 54
rect 38 14 50 54
rect 68 14 80 54
<< pdcontact >>
rect 6 168 18 246
rect 26 180 38 246
rect 46 168 58 246
rect 66 166 78 234
rect 86 166 98 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 20 144 24 166
rect 40 144 44 166
rect 6 138 24 144
rect 32 138 44 144
rect 60 144 64 166
rect 80 144 84 166
rect 60 138 68 144
rect 80 138 88 144
rect 6 102 12 138
rect 32 128 36 138
rect 6 62 12 90
rect 6 58 26 62
rect 22 54 26 58
rect 32 54 36 116
rect 62 128 68 138
rect 62 116 64 128
rect 62 76 68 116
rect 52 72 68 76
rect 84 102 88 138
rect 52 54 56 72
rect 84 62 88 90
rect 62 58 88 62
rect 62 54 66 58
rect 22 10 26 14
rect 32 10 36 14
rect 52 10 56 14
rect 62 10 66 14
<< polycontact >>
rect 24 116 36 128
rect 4 90 16 102
rect 64 116 76 128
rect 84 90 96 102
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 26 246 38 252
rect 18 168 46 174
rect 58 240 86 246
rect 66 160 78 166
rect 44 154 78 160
rect 44 116 50 154
rect 43 54 50 102
rect 8 8 20 14
rect 68 8 80 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 102 17 116
rect 23 102 37 116
rect 43 102 57 116
rect 63 102 77 116
rect 83 102 97 116
<< metal2 >>
rect 6 116 14 134
rect 46 116 54 134
rect 86 116 94 134
rect 26 86 34 102
rect 66 86 74 102
<< m1p >>
rect -6 252 126 268
rect -6 -8 126 8
<< m2p >>
rect 6 118 14 134
rect 46 118 54 134
rect 86 118 94 134
rect 26 86 34 100
rect 66 86 74 100
<< labels >>
rlabel metal2 10 130 10 130 5 A
port 1 n signal input
rlabel metal2 30 88 30 88 7 B
port 2 n signal input
rlabel metal2 90 130 90 130 1 C
port 3 n signal input
rlabel metal2 70 88 70 88 5 D
port 4 n signal input
rlabel metal2 50 130 50 130 5 Y
port 5 n signal output
rlabel metal1 -6 252 106 268 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
