magic
tech scmos
magscale 1 3
timestamp 1725923597
<< checkpaint >>
rect -50 530 1124 870
rect -50 410 2264 530
rect -10 390 2264 410
rect -10 380 2254 390
rect -60 300 2254 380
rect -60 240 2244 300
rect -60 100 2354 240
rect -60 -60 2244 100
use ndiode  ndiode_0
timestamp 1554524574
transform 1 0 500 0 1 470
box 10 10 240 240
use NMOS4  NMOS4_0
timestamp 1554524574
transform 1 0 55 0 1 478
box 5 2 76 134
use p2res  p2res_0
timestamp 1554524574
transform 1 0 42 0 1 422
box 8 8 1032 28
use pdiode  pdiode_0
timestamp 1554524574
transform 1 0 790 0 1 480
box 0 0 270 270
use pipcap  pipcap_0
timestamp 1554524574
transform 1 0 318 0 1 478
box 2 2 142 122
use PMOS4  PMOS4_0
timestamp 1554524574
transform 1 0 180 0 1 480
box 0 0 88 142
use pnp2  pnp2_0
timestamp 1554524574
transform 1 0 -45 0 1 -45
box 45 45 365 365
use pnp5  pnp5_0
timestamp 1554524574
transform 1 0 305 0 1 -45
box 45 45 395 395
use pnp10  pnp10_0
timestamp 1554524574
transform 1 0 685 0 1 -45
box 45 45 445 445
<< end >>
