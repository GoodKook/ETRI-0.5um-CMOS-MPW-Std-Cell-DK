magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -56 -56 164 164
<< genericcontact >>
rect 23 79 29 85
rect 51 79 57 85
rect 79 79 85 85
rect 23 51 29 57
rect 51 51 57 57
rect 79 51 85 57
rect 23 23 29 29
rect 51 23 57 29
rect 79 23 85 29
<< metal1 >>
rect 4 4 104 104
<< end >>
