magic
tech scmos
magscale 1 2
timestamp 1727839497
<< nwell >>
rect 172 252 192 253
rect -12 134 192 252
<< ntransistor >>
rect 40 14 44 34
rect 60 14 64 34
rect 80 14 84 34
<< ptransistor >>
rect 20 166 24 226
rect 40 166 44 226
rect 60 166 64 226
rect 80 166 84 226
rect 124 158 128 218
rect 144 158 148 218
<< ndiffusion >>
rect 38 14 40 34
rect 44 14 46 34
rect 58 14 60 34
rect 64 14 66 34
rect 78 14 80 34
rect 84 14 86 34
<< pdiffusion >>
rect 18 166 20 226
rect 24 166 26 226
rect 38 166 40 226
rect 44 166 46 226
rect 58 166 60 226
rect 64 214 80 226
rect 64 166 66 214
rect 78 166 80 214
rect 84 168 86 226
rect 84 166 98 168
rect 122 158 124 218
rect 128 214 144 218
rect 128 162 130 214
rect 142 162 144 214
rect 128 158 144 162
rect 148 158 150 218
<< ndcontact >>
rect 24 14 38 34
rect 46 14 58 34
rect 66 14 78 34
rect 86 14 98 34
<< pdcontact >>
rect 6 166 18 226
rect 26 166 38 226
rect 46 166 58 226
rect 66 166 78 214
rect 86 168 98 226
rect 110 158 122 218
rect 130 162 142 214
rect 150 158 162 218
<< psubstratepcontact >>
rect -6 -6 186 6
<< nsubstratencontact >>
rect -6 234 186 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 60 226 64 230
rect 80 226 84 230
rect 124 218 128 222
rect 144 218 148 222
rect 20 162 24 166
rect 40 162 44 166
rect 20 158 44 162
rect 40 122 44 158
rect 36 110 44 122
rect 40 34 44 110
rect 60 162 64 166
rect 80 162 84 166
rect 60 158 84 162
rect 60 34 64 158
rect 124 150 128 158
rect 144 150 148 158
rect 98 146 148 150
rect 98 122 104 146
rect 96 110 104 122
rect 98 56 104 110
rect 80 50 104 56
rect 80 34 84 50
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 24 110 36 122
rect 84 110 96 122
rect 64 76 76 88
<< metal1 >>
rect -6 246 186 248
rect -6 232 186 234
rect 26 226 38 232
rect 58 220 86 226
rect 6 160 18 166
rect 46 160 58 166
rect 6 154 58 160
rect 110 220 162 226
rect 110 218 122 220
rect 66 162 78 166
rect 66 158 110 162
rect 150 218 162 220
rect 66 156 122 158
rect 130 146 138 162
rect 115 138 138 146
rect 115 46 123 138
rect 51 40 123 46
rect 51 34 58 40
rect 91 34 98 40
rect 24 8 38 14
rect 66 8 78 14
rect -6 6 186 8
rect -6 -8 186 -6
<< m2contact >>
rect 23 96 37 110
rect 63 88 77 102
rect 83 96 97 110
rect 123 88 137 102
<< metal2 >>
rect 23 82 37 96
rect 63 102 77 116
rect 83 82 97 96
rect 123 102 137 116
<< m2p >>
rect 63 102 77 116
rect 123 102 137 116
rect 23 82 37 96
rect 83 82 97 96
<< labels >>
rlabel metal1 -6 -8 186 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 -6 232 186 248 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal2 23 82 37 96 0 A
port 0 nsew signal input
rlabel metal2 63 102 77 116 0 B
port 1 nsew signal input
rlabel metal2 83 82 97 96 0 C
port 2 nsew signal input
rlabel metal2 123 102 137 116 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
