magic
tech scmos
magscale 1 2
timestamp 1749781447
<< error_s >>
rect 4 5524 5756 5536
rect 4 5284 5756 5296
rect 4 5044 5756 5056
rect 4 4804 5756 4816
rect 4 4564 5756 4576
rect 4 4324 5756 4336
rect 4 4084 5756 4096
rect 4 3844 5756 3856
rect 4 3604 5756 3616
rect 4 3364 5756 3376
rect 4 3124 5756 3136
rect 4 2884 5756 2896
rect 4 2644 5756 2656
rect 4 2404 5756 2416
rect 4 2164 5756 2176
rect 4 1924 5756 1936
rect 4 1684 5756 1696
rect 4 1444 5756 1456
rect 4 1204 5756 1216
rect 4 964 5756 976
rect 4 724 5756 736
rect 4 484 5756 496
rect 4 244 5756 256
rect 4 4 5756 16
<< metal1 >>
rect -62 5298 -2 5538
rect 5730 5522 5822 5538
rect 5257 5383 5263 5453
rect 5257 5377 5283 5383
rect 5277 5363 5283 5377
rect 5277 5357 5293 5363
rect -62 5282 30 5298
rect -62 4818 -2 5282
rect 2767 5217 2783 5223
rect 2777 5143 2783 5217
rect 4687 5217 4713 5223
rect 2767 5137 2783 5143
rect 3017 5197 3033 5203
rect 3017 5123 3023 5197
rect 2987 5117 3023 5123
rect 5762 5058 5822 5522
rect 5730 5042 5822 5058
rect 1887 4977 1903 4983
rect 1897 4923 1903 4977
rect 4347 4957 4393 4963
rect 1897 4917 1913 4923
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 3727 4737 3743 4743
rect 3627 4697 3643 4703
rect 2337 4623 2343 4633
rect 3637 4627 3643 4697
rect 3737 4663 3743 4737
rect 3727 4657 3743 4663
rect 4177 4737 4213 4743
rect 4177 4643 4183 4737
rect 4197 4717 4213 4723
rect 4197 4667 4203 4717
rect 4177 4637 4213 4643
rect 2337 4617 2393 4623
rect 5762 4578 5822 5042
rect 5730 4562 5822 4578
rect 1767 4497 1793 4503
rect 1887 4497 1913 4503
rect 3457 4497 3493 4503
rect 3457 4443 3463 4497
rect 3547 4497 3563 4503
rect 3447 4437 3463 4443
rect 3557 4407 3563 4497
rect 3647 4497 3693 4503
rect 5407 4497 5433 4503
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 1247 4237 1263 4243
rect 1257 4163 1263 4237
rect 2657 4237 2673 4243
rect 1257 4157 1293 4163
rect 2657 4163 2663 4237
rect 2727 4237 2753 4243
rect 3247 4237 3293 4243
rect 3347 4237 3363 4243
rect 2607 4157 2663 4163
rect 3357 4163 3363 4237
rect 3357 4157 3373 4163
rect 5762 4098 5822 4562
rect 5730 4082 5822 4098
rect 587 4017 603 4023
rect 597 3963 603 4017
rect 2767 3997 2793 4003
rect 597 3957 613 3963
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 2257 3717 2273 3723
rect 2257 3703 2263 3717
rect 2247 3697 2263 3703
rect 2347 3677 2413 3683
rect 5762 3618 5822 4082
rect 5730 3602 5822 3618
rect 4047 3537 4063 3543
rect 4057 3527 4063 3537
rect 5037 3537 5053 3543
rect 5037 3467 5043 3537
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 2877 3277 2893 3283
rect 567 3217 593 3223
rect 2877 3203 2883 3277
rect 2877 3197 2893 3203
rect 5762 3138 5822 3602
rect 5730 3122 5822 3138
rect 3157 3077 3173 3083
rect 647 3057 673 3063
rect 2617 3057 2633 3063
rect 2057 3037 2093 3043
rect 2057 2987 2063 3037
rect 2197 2983 2203 3053
rect 2617 3023 2623 3057
rect 2587 3017 2623 3023
rect 3157 3003 3163 3077
rect 3217 3037 3253 3043
rect 3157 2997 3173 3003
rect 2197 2977 2213 2983
rect 3217 2963 3223 3037
rect 3317 2983 3323 3053
rect 3507 3037 3533 3043
rect 4647 3037 4693 3043
rect 3357 3023 3363 3033
rect 3347 3017 3363 3023
rect 3317 2977 3353 2983
rect 3217 2957 3233 2963
rect 5727 2917 5743 2923
rect -62 2882 30 2898
rect 5737 2897 5743 2917
rect -62 2418 -2 2882
rect 647 2797 663 2803
rect 657 2727 663 2797
rect 4117 2743 4123 2813
rect 4797 2797 4813 2803
rect 4117 2737 4133 2743
rect 4797 2723 4803 2797
rect 4797 2717 4813 2723
rect 5762 2658 5822 3122
rect 5730 2642 5822 2658
rect 4587 2557 4613 2563
rect 5287 2557 5313 2563
rect 987 2497 1053 2503
rect 1107 2497 1133 2503
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 847 2317 893 2323
rect 947 2317 973 2323
rect 1207 2297 1283 2303
rect 1277 2243 1283 2297
rect 1277 2237 1293 2243
rect 3017 2243 3023 2293
rect 5247 2257 5273 2263
rect 3007 2237 3023 2243
rect 5762 2178 5822 2642
rect 5730 2162 5822 2178
rect 1047 2077 1083 2083
rect 1077 2047 1083 2077
rect 1107 2077 1133 2083
rect 1577 2043 1583 2133
rect 3487 2097 3553 2103
rect 3957 2097 3973 2103
rect 1577 2037 1593 2043
rect 3957 2023 3963 2097
rect 4527 2097 4543 2103
rect 4537 2027 4543 2097
rect 3947 2017 3963 2023
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 2337 1837 2353 1843
rect 2337 1783 2343 1837
rect 3097 1837 3113 1843
rect 2307 1777 2343 1783
rect 2437 1783 2443 1833
rect 2527 1817 2543 1823
rect 2437 1777 2453 1783
rect 2537 1767 2543 1817
rect 2637 1763 2643 1813
rect 2877 1783 2883 1833
rect 2867 1777 2883 1783
rect 3097 1767 3103 1837
rect 3417 1837 3433 1843
rect 3277 1767 3283 1833
rect 3417 1823 3423 1837
rect 3397 1817 3423 1823
rect 2637 1757 2653 1763
rect 3397 1763 3403 1817
rect 3887 1817 3903 1823
rect 3387 1757 3403 1763
rect 3437 1757 3453 1763
rect 3437 1743 3443 1757
rect 3657 1757 3673 1763
rect 3407 1737 3443 1743
rect 3657 1743 3663 1757
rect 3777 1763 3783 1773
rect 3897 1767 3903 1817
rect 4037 1817 4053 1823
rect 4037 1783 4043 1817
rect 4027 1777 4043 1783
rect 3767 1757 3783 1763
rect 3627 1737 3663 1743
rect 4257 1743 4263 1853
rect 4897 1837 4913 1843
rect 4557 1783 4563 1813
rect 4557 1777 4573 1783
rect 4897 1763 4903 1837
rect 4867 1757 4903 1763
rect 4257 1737 4313 1743
rect 5762 1698 5822 2162
rect 5730 1682 5822 1698
rect 477 1567 483 1613
rect 717 1587 723 1653
rect 3397 1617 3413 1623
rect 937 1523 943 1613
rect 927 1517 943 1523
rect 2957 1483 2963 1613
rect 3397 1563 3403 1617
rect 3907 1617 3943 1623
rect 3487 1597 3503 1603
rect 3387 1557 3403 1563
rect 3497 1563 3503 1597
rect 3497 1557 3553 1563
rect 3937 1563 3943 1617
rect 5067 1617 5093 1623
rect 5187 1597 5253 1603
rect 3937 1557 3953 1563
rect 4147 1557 4193 1563
rect 2947 1477 2963 1483
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 137 1423 143 1443
rect 107 1417 143 1423
rect 3347 1377 3393 1383
rect 417 1357 433 1363
rect 417 1303 423 1357
rect 3137 1337 3193 1343
rect 367 1297 423 1303
rect 947 1297 973 1303
rect 1597 1303 1603 1333
rect 1597 1297 1633 1303
rect 2097 1303 2103 1333
rect 2087 1297 2103 1303
rect 3137 1283 3143 1337
rect 3987 1337 4003 1343
rect 3997 1307 4003 1337
rect 3377 1297 3413 1303
rect 3377 1287 3383 1297
rect 3127 1277 3143 1283
rect 3667 1257 3733 1263
rect 5762 1218 5822 1682
rect 5730 1202 5822 1218
rect 987 1157 1003 1163
rect 437 1117 453 1123
rect 437 1107 443 1117
rect 997 1083 1003 1157
rect 2147 1137 2163 1143
rect 1117 1103 1123 1113
rect 1117 1097 1133 1103
rect 997 1077 1033 1083
rect 2157 1083 2163 1137
rect 2157 1077 2173 1083
rect 2237 1083 2243 1153
rect 2707 1137 2723 1143
rect 2717 1087 2723 1137
rect 2847 1137 2863 1143
rect 2227 1077 2243 1083
rect 2137 1043 2143 1053
rect 2137 1037 2173 1043
rect 2857 1043 2863 1137
rect 2877 1137 2893 1143
rect 2877 1067 2883 1137
rect 4037 1137 4053 1143
rect 4037 1107 4043 1137
rect 4057 1117 4073 1123
rect 4057 1083 4063 1117
rect 4037 1077 4063 1083
rect 4037 1067 4043 1077
rect 2857 1037 2873 1043
rect 3447 1037 3473 1043
rect 4477 1043 4483 1113
rect 4477 1037 4493 1043
rect -62 962 30 978
rect -62 498 -2 962
rect 2217 823 2223 873
rect 2217 817 2233 823
rect 2397 823 2403 893
rect 3747 877 3793 883
rect 2447 857 2463 863
rect 2387 817 2403 823
rect 2457 823 2463 857
rect 2457 817 2473 823
rect 3237 823 3243 873
rect 3207 817 3243 823
rect 4797 807 4803 873
rect 3107 797 3133 803
rect 5762 738 5822 1202
rect 5730 722 5822 738
rect 5057 657 5073 663
rect 1257 637 1273 643
rect 1257 563 1263 637
rect 3457 637 3513 643
rect 3457 603 3463 637
rect 5057 607 5063 657
rect 5247 637 5293 643
rect 3447 597 3463 603
rect 1257 557 1273 563
rect -62 482 30 498
rect -62 18 -2 482
rect 4707 397 4753 403
rect 2267 317 2313 323
rect 5762 258 5822 722
rect 5730 242 5822 258
rect 847 157 873 163
rect -62 2 30 18
rect 5762 2 5822 242
<< m2contact >>
rect 5253 5453 5267 5467
rect 5293 5353 5307 5367
rect 413 5273 427 5287
rect 2753 5213 2767 5227
rect 2753 5133 2767 5147
rect 4673 5213 4687 5227
rect 4713 5213 4727 5227
rect 2973 5113 2987 5127
rect 3033 5193 3047 5207
rect 1873 4973 1887 4987
rect 4333 4953 4347 4967
rect 4393 4953 4407 4967
rect 1913 4913 1927 4927
rect 1813 4813 1827 4827
rect 113 4793 127 4807
rect 1333 4793 1347 4807
rect 4613 4793 4627 4807
rect 5733 4793 5747 4807
rect 3713 4733 3727 4747
rect 3613 4693 3627 4707
rect 2333 4633 2347 4647
rect 3713 4653 3727 4667
rect 4213 4733 4227 4747
rect 4213 4713 4227 4727
rect 4193 4653 4207 4667
rect 4213 4633 4227 4647
rect 2393 4613 2407 4627
rect 3633 4613 3647 4627
rect 1753 4493 1767 4507
rect 1793 4493 1807 4507
rect 1873 4493 1887 4507
rect 1913 4493 1927 4507
rect 3433 4433 3447 4447
rect 3493 4493 3507 4507
rect 3533 4493 3547 4507
rect 3633 4493 3647 4507
rect 3693 4493 3707 4507
rect 5393 4493 5407 4507
rect 5433 4493 5447 4507
rect 3553 4393 3567 4407
rect 5113 4333 5127 4347
rect 513 4313 527 4327
rect 5733 4313 5747 4327
rect 1233 4233 1247 4247
rect 1293 4153 1307 4167
rect 2593 4153 2607 4167
rect 2673 4233 2687 4247
rect 2713 4233 2727 4247
rect 2753 4233 2767 4247
rect 3233 4233 3247 4247
rect 3293 4233 3307 4247
rect 3333 4233 3347 4247
rect 3373 4153 3387 4167
rect 573 4013 587 4027
rect 2753 3993 2767 4007
rect 2793 3993 2807 4007
rect 613 3953 627 3967
rect 93 3833 107 3847
rect 3133 3833 3147 3847
rect 4053 3833 4067 3847
rect 5033 3833 5047 3847
rect 5733 3833 5747 3847
rect 2233 3693 2247 3707
rect 2273 3713 2287 3727
rect 2333 3673 2347 3687
rect 2413 3673 2427 3687
rect 4033 3533 4047 3547
rect 4053 3513 4067 3527
rect 5053 3533 5067 3547
rect 5033 3453 5047 3467
rect 5733 3373 5747 3387
rect 3073 3353 3087 3367
rect 4813 3353 4827 3367
rect 4973 3353 4987 3367
rect 553 3213 567 3227
rect 593 3213 607 3227
rect 2893 3273 2907 3287
rect 2893 3193 2907 3207
rect 633 3053 647 3067
rect 673 3053 687 3067
rect 2193 3053 2207 3067
rect 2093 3033 2107 3047
rect 2053 2973 2067 2987
rect 2573 3013 2587 3027
rect 2633 3053 2647 3067
rect 3173 3073 3187 3087
rect 3313 3053 3327 3067
rect 3173 2993 3187 3007
rect 2213 2973 2227 2987
rect 3253 3033 3267 3047
rect 3353 3033 3367 3047
rect 3493 3033 3507 3047
rect 3533 3033 3547 3047
rect 4633 3033 4647 3047
rect 4693 3033 4707 3047
rect 3333 3013 3347 3027
rect 3353 2973 3367 2987
rect 3233 2953 3247 2967
rect 5713 2913 5727 2927
rect 1473 2893 1487 2907
rect 993 2873 1007 2887
rect 4093 2873 4107 2887
rect 4113 2813 4127 2827
rect 633 2793 647 2807
rect 4133 2733 4147 2747
rect 653 2713 667 2727
rect 4813 2793 4827 2807
rect 4813 2713 4827 2727
rect 4573 2553 4587 2567
rect 4613 2553 4627 2567
rect 5273 2553 5287 2567
rect 5313 2553 5327 2567
rect 973 2493 987 2507
rect 1053 2493 1067 2507
rect 1093 2493 1107 2507
rect 1133 2493 1147 2507
rect 4593 2413 4607 2427
rect 3113 2393 3127 2407
rect 833 2313 847 2327
rect 893 2313 907 2327
rect 933 2313 947 2327
rect 973 2313 987 2327
rect 1193 2293 1207 2307
rect 3013 2293 3027 2307
rect 1293 2233 1307 2247
rect 2993 2233 3007 2247
rect 5233 2253 5247 2267
rect 5273 2253 5287 2267
rect 1573 2133 1587 2147
rect 1033 2073 1047 2087
rect 1093 2073 1107 2087
rect 1133 2073 1147 2087
rect 1073 2033 1087 2047
rect 3473 2093 3487 2107
rect 3553 2093 3567 2107
rect 1593 2033 1607 2047
rect 3933 2013 3947 2027
rect 3973 2093 3987 2107
rect 4513 2093 4527 2107
rect 4533 2013 4547 2027
rect 5093 1913 5107 1927
rect 4253 1853 4267 1867
rect 2293 1773 2307 1787
rect 2353 1833 2367 1847
rect 2433 1833 2447 1847
rect 2873 1833 2887 1847
rect 2513 1813 2527 1827
rect 2453 1773 2467 1787
rect 2633 1813 2647 1827
rect 2533 1753 2547 1767
rect 2853 1773 2867 1787
rect 3113 1833 3127 1847
rect 3273 1833 3287 1847
rect 3433 1833 3447 1847
rect 2653 1753 2667 1767
rect 3093 1753 3107 1767
rect 3273 1753 3287 1767
rect 3373 1753 3387 1767
rect 3873 1813 3887 1827
rect 3773 1773 3787 1787
rect 3393 1733 3407 1747
rect 3453 1753 3467 1767
rect 3613 1733 3627 1747
rect 3673 1753 3687 1767
rect 3753 1753 3767 1767
rect 4013 1773 4027 1787
rect 4053 1813 4067 1827
rect 3893 1753 3907 1767
rect 4553 1813 4567 1827
rect 4573 1773 4587 1787
rect 4853 1753 4867 1767
rect 4913 1833 4927 1847
rect 4313 1733 4327 1747
rect 713 1653 727 1667
rect 473 1613 487 1627
rect 933 1613 947 1627
rect 2953 1613 2967 1627
rect 713 1573 727 1587
rect 473 1553 487 1567
rect 913 1513 927 1527
rect 2933 1473 2947 1487
rect 3373 1553 3387 1567
rect 3413 1613 3427 1627
rect 3893 1613 3907 1627
rect 3473 1593 3487 1607
rect 3553 1553 3567 1567
rect 5053 1613 5067 1627
rect 5093 1613 5107 1627
rect 5173 1593 5187 1607
rect 5253 1593 5267 1607
rect 3953 1553 3967 1567
rect 4133 1553 4147 1567
rect 4193 1553 4207 1567
rect 93 1413 107 1427
rect 2233 1433 2247 1447
rect 5573 1433 5587 1447
rect 3333 1373 3347 1387
rect 3393 1373 3407 1387
rect 353 1293 367 1307
rect 433 1353 447 1367
rect 1593 1333 1607 1347
rect 2093 1333 2107 1347
rect 933 1293 947 1307
rect 973 1293 987 1307
rect 1633 1293 1647 1307
rect 2073 1293 2087 1307
rect 3113 1273 3127 1287
rect 3193 1333 3207 1347
rect 3973 1333 3987 1347
rect 3413 1293 3427 1307
rect 3993 1293 4007 1307
rect 3373 1273 3387 1287
rect 3653 1253 3667 1267
rect 3733 1253 3747 1267
rect 973 1153 987 1167
rect 453 1113 467 1127
rect 433 1093 447 1107
rect 2233 1153 2247 1167
rect 2133 1133 2147 1147
rect 1113 1113 1127 1127
rect 1133 1093 1147 1107
rect 1033 1073 1047 1087
rect 2173 1073 2187 1087
rect 2213 1073 2227 1087
rect 2693 1133 2707 1147
rect 2833 1133 2847 1147
rect 2713 1073 2727 1087
rect 2133 1053 2147 1067
rect 2173 1033 2187 1047
rect 2893 1133 2907 1147
rect 4053 1133 4067 1147
rect 4033 1093 4047 1107
rect 4073 1113 4087 1127
rect 4473 1113 4487 1127
rect 2873 1053 2887 1067
rect 4033 1053 4047 1067
rect 2873 1033 2887 1047
rect 3433 1033 3447 1047
rect 3473 1033 3487 1047
rect 4493 1033 4507 1047
rect 513 953 527 967
rect 2393 893 2407 907
rect 2213 873 2227 887
rect 2233 813 2247 827
rect 2373 813 2387 827
rect 3233 873 3247 887
rect 3733 873 3747 887
rect 3793 873 3807 887
rect 4793 873 4807 887
rect 2433 853 2447 867
rect 2473 813 2487 827
rect 3193 813 3207 827
rect 3093 793 3107 807
rect 3133 793 3147 807
rect 4793 793 4807 807
rect 1273 633 1287 647
rect 3433 593 3447 607
rect 3513 633 3527 647
rect 5073 653 5087 667
rect 5233 633 5247 647
rect 5293 633 5307 647
rect 5053 593 5067 607
rect 1273 553 1287 567
rect 493 473 507 487
rect 1273 473 1287 487
rect 3353 473 3367 487
rect 4613 473 4627 487
rect 5733 473 5747 487
rect 4693 393 4707 407
rect 4753 393 4767 407
rect 2253 313 2267 327
rect 2313 313 2327 327
rect 833 153 847 167
rect 873 153 887 167
rect 673 13 687 27
rect 5733 13 5747 27
<< metal2 >>
rect 76 5436 83 5453
rect 116 5436 143 5443
rect 56 5416 63 5433
rect 96 5387 103 5423
rect 136 5403 143 5436
rect 156 5407 163 5453
rect 196 5416 203 5453
rect 256 5436 263 5453
rect 296 5436 343 5443
rect 116 5396 143 5403
rect 56 5183 63 5373
rect 116 5183 123 5396
rect 176 5367 183 5403
rect 36 5176 63 5183
rect 96 5176 123 5183
rect 36 5127 43 5176
rect 116 5087 123 5176
rect 196 5156 203 5173
rect 156 5087 163 5143
rect 296 5127 303 5163
rect 336 5147 343 5436
rect 396 5416 423 5423
rect 356 5327 363 5403
rect 416 5287 423 5416
rect 796 5423 803 5453
rect 776 5416 803 5423
rect 427 5276 443 5283
rect 436 5167 443 5276
rect 456 5183 463 5313
rect 456 5176 483 5183
rect 356 5127 363 5143
rect 76 4936 103 4943
rect 36 4767 43 4923
rect 96 4803 103 4936
rect 96 4796 113 4803
rect 96 4696 103 4713
rect 116 4667 123 4793
rect 176 4727 183 5113
rect 376 5047 383 5123
rect 196 4976 203 5033
rect 376 4936 383 5013
rect 396 4987 403 5133
rect 396 4787 403 4973
rect 456 4927 463 4943
rect 196 4663 203 4773
rect 476 4767 483 5176
rect 816 5163 823 5413
rect 796 5156 823 5163
rect 616 5067 623 5123
rect 516 4976 523 5053
rect 496 4956 503 4973
rect 616 4923 623 4993
rect 776 4956 783 5113
rect 796 5047 803 5156
rect 836 5087 843 5393
rect 796 5027 803 5033
rect 656 4936 663 4953
rect 696 4923 703 4953
rect 616 4916 643 4923
rect 676 4916 703 4923
rect 236 4696 243 4753
rect 276 4667 283 4683
rect 76 4456 83 4653
rect 136 4647 143 4663
rect 176 4656 203 4663
rect 36 4223 43 4443
rect 36 4216 63 4223
rect 56 4007 63 4216
rect 176 4187 183 4656
rect 556 4496 563 4693
rect 576 4607 583 4683
rect 656 4676 663 4693
rect 736 4676 743 4893
rect 756 4787 763 4943
rect 576 4467 583 4593
rect 636 4476 643 4673
rect 776 4643 783 4913
rect 796 4887 803 4973
rect 836 4907 843 5073
rect 896 4983 903 5153
rect 876 4976 903 4983
rect 816 4696 823 4713
rect 916 4707 923 5453
rect 996 5436 1023 5443
rect 976 5407 983 5423
rect 1016 5387 1023 5436
rect 1036 5407 1043 5423
rect 1216 5403 1223 5473
rect 1416 5456 1483 5463
rect 1256 5416 1263 5453
rect 1196 5396 1223 5403
rect 936 5147 943 5173
rect 976 5156 983 5173
rect 996 5007 1003 5173
rect 1016 5007 1023 5153
rect 1036 5147 1043 5183
rect 1096 5167 1103 5393
rect 1136 5176 1143 5253
rect 1196 5183 1203 5396
rect 1296 5403 1303 5433
rect 1336 5416 1343 5433
rect 1276 5396 1303 5403
rect 1356 5367 1363 5393
rect 1176 5176 1203 5183
rect 1156 5127 1163 5153
rect 1196 5083 1203 5176
rect 1236 5107 1243 5143
rect 1396 5143 1403 5373
rect 1416 5167 1423 5456
rect 1476 5436 1483 5456
rect 1516 5456 1543 5463
rect 1616 5456 1623 5473
rect 1456 5407 1463 5423
rect 1496 5416 1503 5433
rect 1376 5136 1403 5143
rect 1196 5076 1223 5083
rect 996 4983 1003 4993
rect 996 4976 1023 4983
rect 1056 4956 1063 4973
rect 1096 4943 1103 4953
rect 956 4707 963 4713
rect 756 4636 783 4643
rect 756 4527 763 4636
rect 356 4456 373 4463
rect 356 4203 363 4456
rect 456 4427 463 4463
rect 536 4447 543 4463
rect 596 4456 623 4463
rect 596 4447 603 4456
rect 656 4407 663 4463
rect 716 4443 723 4473
rect 756 4456 763 4473
rect 796 4443 803 4673
rect 856 4667 863 4693
rect 876 4643 883 4683
rect 876 4636 893 4643
rect 856 4476 863 4493
rect 716 4436 743 4443
rect 776 4436 803 4443
rect 516 4207 523 4313
rect 356 4196 383 4203
rect 456 4196 483 4203
rect 196 4147 203 4163
rect 56 3963 63 3993
rect 376 3987 383 4196
rect 476 4167 483 4196
rect 716 4196 723 4436
rect 776 4247 783 4436
rect 536 3996 543 4173
rect 796 4167 803 4413
rect 836 4367 843 4463
rect 896 4447 903 4633
rect 916 4487 923 4653
rect 996 4443 1003 4893
rect 1036 4887 1043 4943
rect 1096 4936 1123 4943
rect 1196 4936 1203 5033
rect 1056 4787 1063 4913
rect 1116 4807 1123 4936
rect 1056 4696 1063 4773
rect 1076 4667 1083 4683
rect 1096 4667 1103 4703
rect 1116 4567 1123 4673
rect 1136 4527 1143 4733
rect 1196 4696 1203 4733
rect 1216 4667 1223 5076
rect 1236 4927 1243 5093
rect 1396 4887 1403 5136
rect 1456 5107 1463 5393
rect 1516 5267 1523 5456
rect 1716 5436 1723 5453
rect 1756 5436 1783 5443
rect 1576 5423 1583 5433
rect 1556 5416 1583 5423
rect 1776 5387 1783 5436
rect 1836 5427 1843 5473
rect 1856 5416 1883 5423
rect 2156 5416 2183 5423
rect 1816 5387 1823 5403
rect 1496 4936 1503 5173
rect 1576 4967 1583 5253
rect 1256 4727 1263 4773
rect 1256 4663 1263 4713
rect 1336 4687 1343 4793
rect 1396 4707 1403 4753
rect 1236 4647 1243 4663
rect 1256 4656 1283 4663
rect 1256 4603 1263 4656
rect 1396 4663 1403 4693
rect 1436 4663 1443 4753
rect 1376 4656 1403 4663
rect 1416 4656 1443 4663
rect 1236 4596 1263 4603
rect 1056 4476 1063 4513
rect 976 4436 1003 4443
rect 896 4427 903 4433
rect 976 4423 983 4436
rect 956 4416 983 4423
rect 956 4407 963 4416
rect 556 4147 563 4163
rect 596 4016 623 4023
rect 576 3996 583 4013
rect 596 3987 603 4016
rect 76 3976 103 3983
rect 36 3956 63 3963
rect 96 3847 103 3976
rect 636 3963 643 3983
rect 627 3956 643 3963
rect 176 3736 203 3743
rect 16 3716 43 3723
rect 16 3687 23 3716
rect 56 3627 63 3683
rect 116 3627 123 3723
rect 196 3707 203 3736
rect 216 3687 223 3723
rect 216 3667 223 3673
rect 76 3496 83 3513
rect 56 3427 63 3483
rect 96 3447 103 3483
rect 56 3236 63 3253
rect 96 3203 103 3413
rect 116 3367 123 3493
rect 176 3476 183 3533
rect 196 3496 203 3513
rect 236 3487 243 3733
rect 296 3716 323 3723
rect 256 3507 263 3713
rect 296 3707 303 3716
rect 296 3496 303 3533
rect 276 3467 283 3483
rect 156 3227 163 3433
rect 176 3236 183 3353
rect 316 3347 323 3473
rect 336 3447 343 3683
rect 376 3567 383 3703
rect 516 3687 523 3703
rect 556 3683 563 3773
rect 576 3736 603 3743
rect 636 3736 643 3773
rect 576 3687 583 3736
rect 536 3676 563 3683
rect 616 3547 623 3723
rect 656 3607 663 4153
rect 676 3787 683 4133
rect 836 4127 843 4333
rect 856 4183 863 4193
rect 856 4176 873 4183
rect 936 4183 943 4213
rect 956 4207 963 4393
rect 1076 4227 1083 4353
rect 1116 4243 1123 4473
rect 1136 4447 1143 4493
rect 1216 4476 1223 4493
rect 1096 4236 1123 4243
rect 996 4196 1003 4213
rect 916 4176 943 4183
rect 856 4127 863 4153
rect 736 3996 743 4113
rect 756 4027 763 4093
rect 896 4087 903 4163
rect 1016 4087 1023 4113
rect 716 3767 723 3993
rect 676 3647 683 3703
rect 456 3496 483 3503
rect 376 3483 383 3493
rect 376 3476 403 3483
rect 476 3467 483 3496
rect 536 3467 543 3483
rect 76 3047 83 3203
rect 96 3196 123 3203
rect 76 3016 83 3033
rect 56 2987 63 3003
rect 56 2756 63 2933
rect 96 2747 103 2993
rect 116 2947 123 3196
rect 176 3056 183 3173
rect 256 3047 263 3243
rect 376 3236 383 3253
rect 316 3207 323 3223
rect 336 3187 343 3233
rect 356 3187 363 3223
rect 416 3207 423 3243
rect 436 3227 443 3333
rect 476 3247 483 3453
rect 536 3367 543 3453
rect 556 3287 563 3493
rect 576 3487 583 3513
rect 596 3496 603 3513
rect 696 3496 703 3653
rect 736 3527 743 3733
rect 756 3647 763 4013
rect 796 4003 803 4053
rect 816 4016 823 4033
rect 776 3996 803 4003
rect 836 3996 843 4073
rect 896 4047 903 4073
rect 776 3747 783 3996
rect 856 3947 863 4033
rect 916 4027 923 4053
rect 936 4016 943 4033
rect 916 3996 923 4013
rect 976 4007 983 4053
rect 1016 3996 1023 4073
rect 1036 4067 1043 4203
rect 1056 4167 1063 4213
rect 676 3463 683 3493
rect 656 3456 683 3463
rect 656 3267 663 3456
rect 756 3447 763 3483
rect 776 3327 783 3493
rect 796 3307 803 3753
rect 856 3627 863 3933
rect 916 3727 923 3953
rect 956 3867 963 3983
rect 876 3687 883 3703
rect 976 3687 983 3993
rect 856 3503 863 3613
rect 916 3536 963 3543
rect 836 3496 863 3503
rect 916 3483 923 3536
rect 896 3476 923 3483
rect 1016 3367 1023 3713
rect 1036 3427 1043 3973
rect 1056 3716 1063 3733
rect 1076 3667 1083 4193
rect 1096 4027 1103 4236
rect 1156 4216 1163 4233
rect 1136 4183 1143 4203
rect 1116 4176 1143 4183
rect 1096 3647 1103 4013
rect 1076 3507 1083 3553
rect 1116 3407 1123 4176
rect 1136 3747 1143 4033
rect 1176 3976 1183 4413
rect 1196 4367 1203 4473
rect 1236 4263 1243 4596
rect 1276 4456 1283 4573
rect 1296 4507 1303 4643
rect 1416 4483 1423 4656
rect 1456 4523 1463 4653
rect 1476 4647 1483 4793
rect 1336 4476 1363 4483
rect 1356 4447 1363 4476
rect 1396 4476 1423 4483
rect 1436 4516 1463 4523
rect 1396 4347 1403 4476
rect 1436 4456 1443 4516
rect 1456 4436 1463 4493
rect 1476 4456 1483 4633
rect 1516 4607 1523 4673
rect 1596 4667 1603 5013
rect 1636 4976 1643 5013
rect 1656 4956 1663 4993
rect 1756 4983 1763 5273
rect 1816 5187 1823 5373
rect 1776 5147 1783 5163
rect 1776 5047 1783 5133
rect 1756 4976 1783 4983
rect 1756 4907 1763 4943
rect 1576 4496 1583 4593
rect 1596 4567 1603 4613
rect 1616 4607 1623 4643
rect 1756 4627 1763 4713
rect 1556 4476 1563 4493
rect 1596 4476 1603 4553
rect 1656 4496 1663 4513
rect 1616 4463 1623 4493
rect 1716 4476 1723 4533
rect 1756 4463 1763 4493
rect 1616 4456 1643 4463
rect 1236 4256 1263 4263
rect 1236 4216 1243 4233
rect 1216 4147 1223 4203
rect 1156 3947 1163 3963
rect 1256 3747 1263 4256
rect 1276 4187 1283 4233
rect 1356 4196 1383 4203
rect 1336 4163 1343 4183
rect 1307 4156 1343 4163
rect 1196 3703 1203 3733
rect 1276 3707 1283 4073
rect 1356 4027 1363 4173
rect 1376 4147 1383 4196
rect 1396 4107 1403 4193
rect 1416 4047 1423 4253
rect 1576 4227 1583 4453
rect 1696 4427 1703 4463
rect 1736 4456 1763 4463
rect 1656 4216 1663 4393
rect 1476 4127 1483 4203
rect 1316 3996 1343 4003
rect 1376 3996 1403 4003
rect 1416 3996 1423 4013
rect 1456 3996 1463 4033
rect 1316 3987 1323 3996
rect 1316 3767 1323 3973
rect 1396 3887 1403 3996
rect 1476 3967 1483 4013
rect 1496 3947 1503 4153
rect 1516 3967 1523 4203
rect 1556 4196 1563 4213
rect 1576 4147 1583 4153
rect 1636 4127 1643 4203
rect 1536 3976 1543 4013
rect 1556 3996 1563 4113
rect 1596 4067 1603 4073
rect 1596 3996 1603 4053
rect 1616 4007 1623 4073
rect 1676 4003 1683 4333
rect 1656 3996 1683 4003
rect 1696 3996 1703 4373
rect 1776 4267 1783 4976
rect 1796 4727 1803 4933
rect 1816 4927 1823 5053
rect 1836 4967 1843 5413
rect 1856 5156 1863 5253
rect 1876 5167 1883 5416
rect 2176 5407 2183 5416
rect 1976 5163 1983 5393
rect 1896 5156 1923 5163
rect 1976 5156 2003 5163
rect 1876 5067 1883 5153
rect 1896 5103 1903 5156
rect 1976 5147 1983 5156
rect 1896 5096 1923 5103
rect 1856 4976 1863 5033
rect 1876 4956 1883 4973
rect 1816 4827 1823 4913
rect 1816 4527 1823 4673
rect 1807 4496 1843 4503
rect 1836 4476 1843 4496
rect 1876 4476 1883 4493
rect 1816 4387 1823 4463
rect 1856 4427 1863 4463
rect 1896 4367 1903 5053
rect 1916 4947 1923 5096
rect 1936 4936 1943 4973
rect 1956 4916 1963 5013
rect 1976 4936 1983 5033
rect 1916 4747 1923 4913
rect 1936 4663 1943 4873
rect 1976 4676 1983 4893
rect 1996 4727 2003 4923
rect 2016 4907 2023 5073
rect 2036 4956 2043 5053
rect 2156 5007 2163 5013
rect 2076 4956 2103 4963
rect 2156 4956 2163 4993
rect 2196 4983 2203 5433
rect 2276 5267 2283 5453
rect 2336 5436 2363 5443
rect 2336 5387 2343 5436
rect 2276 5123 2283 5253
rect 2276 5116 2303 5123
rect 2176 4976 2203 4983
rect 2096 4787 2103 4956
rect 2176 4767 2183 4976
rect 2216 4967 2223 4993
rect 2296 4987 2303 5116
rect 2316 5007 2323 5213
rect 2336 5176 2343 5373
rect 2416 5176 2423 5513
rect 2536 5443 2543 5533
rect 2516 5436 2543 5443
rect 2536 5383 2543 5436
rect 2736 5423 2743 5583
rect 2776 5527 2783 5583
rect 2816 5547 2823 5583
rect 2616 5407 2623 5423
rect 2736 5416 2763 5423
rect 2516 5376 2543 5383
rect 2516 5143 2523 5376
rect 2756 5287 2763 5416
rect 2756 5207 2763 5213
rect 2396 5127 2403 5143
rect 2236 4976 2283 4983
rect 2096 4696 2103 4713
rect 2016 4676 2043 4683
rect 2036 4667 2043 4676
rect 2076 4667 2083 4683
rect 1936 4656 1963 4663
rect 1756 4216 1763 4233
rect 1796 4216 1803 4293
rect 1776 4167 1783 4203
rect 1816 4127 1823 4353
rect 1916 4307 1923 4493
rect 1736 4027 1743 4033
rect 1736 4007 1743 4013
rect 1776 4007 1783 4113
rect 1836 4047 1843 4273
rect 1936 4227 1943 4593
rect 1996 4507 2003 4643
rect 2036 4476 2043 4513
rect 1996 4267 2003 4463
rect 2056 4427 2063 4453
rect 2096 4267 2103 4513
rect 2116 4247 2123 4733
rect 2196 4703 2203 4943
rect 2236 4707 2243 4976
rect 2316 4976 2323 4993
rect 2296 4956 2303 4973
rect 2196 4696 2223 4703
rect 2136 4647 2143 4693
rect 2216 4683 2223 4696
rect 2216 4676 2243 4683
rect 2256 4676 2263 4713
rect 2156 4507 2163 4673
rect 2336 4667 2343 4933
rect 2176 4587 2183 4663
rect 2156 4387 2163 4453
rect 2176 4287 2183 4443
rect 2216 4436 2223 4553
rect 2236 4456 2243 4613
rect 2316 4587 2323 4663
rect 2336 4627 2343 4633
rect 2316 4496 2323 4513
rect 2356 4476 2363 4613
rect 2376 4547 2383 5093
rect 2436 4916 2443 5113
rect 2456 5087 2463 5143
rect 2516 5136 2543 5143
rect 2556 5136 2583 5143
rect 2456 4936 2463 4993
rect 2476 4727 2483 4923
rect 2496 4696 2503 4973
rect 2536 4803 2543 5033
rect 2556 4927 2563 5136
rect 2596 4983 2603 5173
rect 2736 5147 2743 5183
rect 2776 5167 2783 5413
rect 2836 5407 2843 5423
rect 2956 5403 2963 5473
rect 3016 5456 3023 5473
rect 2936 5396 2963 5403
rect 2976 5387 2983 5453
rect 3056 5436 3083 5443
rect 2996 5407 3003 5423
rect 3016 5207 3023 5413
rect 3036 5367 3043 5423
rect 3076 5407 3083 5436
rect 3096 5383 3103 5583
rect 3136 5527 3143 5583
rect 3236 5447 3243 5453
rect 3076 5376 3103 5383
rect 3116 5436 3143 5443
rect 3076 5347 3083 5376
rect 2836 5176 2843 5193
rect 2916 5176 2943 5183
rect 2976 5176 3003 5183
rect 2756 5147 2763 5163
rect 2656 4987 2663 5013
rect 2576 4976 2603 4983
rect 2576 4956 2583 4976
rect 2656 4956 2663 4973
rect 2596 4923 2603 4943
rect 2576 4916 2603 4923
rect 2536 4796 2563 4803
rect 2536 4707 2543 4773
rect 2396 4647 2403 4663
rect 2416 4623 2423 4643
rect 2407 4616 2423 4623
rect 2416 4496 2423 4553
rect 2396 4476 2403 4493
rect 2296 4447 2303 4453
rect 1616 3987 1623 3993
rect 1336 3736 1343 3773
rect 1356 3736 1363 3873
rect 1396 3736 1403 3753
rect 1416 3727 1423 3773
rect 1516 3747 1523 3953
rect 1136 3627 1143 3703
rect 1176 3696 1203 3703
rect 1156 3547 1163 3683
rect 1156 3516 1183 3523
rect 1176 3367 1183 3516
rect 1196 3387 1203 3503
rect 536 3236 563 3243
rect 556 3227 563 3236
rect 596 3227 603 3243
rect 616 3227 623 3263
rect 796 3243 803 3273
rect 776 3236 803 3243
rect 496 3207 503 3223
rect 476 3183 483 3193
rect 476 3176 503 3183
rect 136 3036 163 3043
rect 196 3036 223 3043
rect 136 2987 143 3036
rect 216 3007 223 3036
rect 396 3036 403 3053
rect 436 3047 443 3153
rect 496 3056 503 3176
rect 636 3147 643 3233
rect 676 3207 683 3233
rect 816 3227 823 3313
rect 836 3256 843 3293
rect 596 3067 603 3133
rect 676 3067 683 3193
rect 716 3147 723 3223
rect 796 3056 823 3063
rect 516 3036 543 3043
rect 376 3016 383 3033
rect 536 3027 543 3036
rect 596 3036 603 3053
rect 636 3036 643 3053
rect 156 2767 163 2973
rect 216 2763 223 2833
rect 336 2827 343 2993
rect 256 2776 283 2783
rect 196 2756 223 2763
rect 76 2627 83 2723
rect 136 2607 143 2733
rect 76 2536 83 2573
rect 56 2503 63 2523
rect 96 2507 103 2523
rect 56 2496 83 2503
rect 16 2047 23 2373
rect 36 2276 63 2283
rect 36 2083 43 2276
rect 76 2207 83 2496
rect 116 2283 123 2593
rect 156 2287 163 2543
rect 176 2307 183 2713
rect 236 2707 243 2753
rect 256 2727 263 2776
rect 336 2767 343 2813
rect 416 2807 423 3013
rect 396 2767 403 2773
rect 356 2747 363 2763
rect 416 2727 423 2743
rect 416 2687 423 2713
rect 256 2536 263 2613
rect 436 2567 443 2913
rect 456 2723 463 2793
rect 496 2756 503 2773
rect 456 2716 483 2723
rect 296 2523 303 2553
rect 356 2536 363 2553
rect 396 2523 403 2553
rect 476 2527 483 2716
rect 516 2647 523 2743
rect 536 2576 543 2763
rect 556 2747 563 2773
rect 556 2556 563 2573
rect 276 2516 303 2523
rect 336 2367 343 2523
rect 376 2516 403 2523
rect 416 2467 423 2523
rect 216 2296 223 2313
rect 116 2276 143 2283
rect 36 2076 63 2083
rect 96 2076 103 2113
rect 136 2083 143 2276
rect 156 2247 163 2273
rect 196 2267 203 2283
rect 236 2267 243 2293
rect 196 2227 203 2253
rect 256 2247 263 2313
rect 136 2076 163 2083
rect 196 2076 203 2093
rect 16 1487 23 1913
rect 36 1816 43 1893
rect 56 1767 63 2033
rect 76 1947 83 2063
rect 156 2063 163 2076
rect 156 2056 183 2063
rect 56 1603 63 1753
rect 76 1623 83 1803
rect 96 1647 103 1893
rect 176 1807 183 2056
rect 216 2047 223 2093
rect 236 1967 243 2233
rect 256 2007 263 2193
rect 276 2107 283 2253
rect 316 2247 323 2263
rect 296 2187 303 2243
rect 296 2087 303 2133
rect 316 1987 323 2043
rect 336 1927 343 2353
rect 396 2276 403 2293
rect 436 2267 443 2493
rect 456 2487 463 2523
rect 376 2227 383 2243
rect 416 2167 423 2263
rect 436 2147 443 2253
rect 456 2187 463 2293
rect 476 2127 483 2513
rect 576 2507 583 3033
rect 596 2776 603 2933
rect 636 2807 643 2993
rect 656 2947 663 3013
rect 676 2847 683 3053
rect 736 3016 743 3053
rect 636 2776 643 2793
rect 616 2747 623 2763
rect 656 2743 663 2813
rect 676 2807 683 2833
rect 696 2756 703 2793
rect 656 2736 683 2743
rect 656 2627 663 2713
rect 736 2667 743 2763
rect 756 2647 763 3003
rect 796 2927 803 3056
rect 836 2787 843 3013
rect 856 3007 863 3293
rect 896 3183 903 3253
rect 1156 3243 1163 3353
rect 1216 3327 1223 3653
rect 1236 3527 1243 3683
rect 1256 3647 1263 3703
rect 1316 3687 1323 3723
rect 1516 3667 1523 3703
rect 1276 3516 1283 3533
rect 1236 3487 1243 3513
rect 1156 3236 1183 3243
rect 876 3176 903 3183
rect 596 2576 643 2583
rect 596 2567 603 2576
rect 656 2556 663 2573
rect 496 2263 503 2273
rect 496 2256 523 2263
rect 556 2243 563 2263
rect 556 2236 603 2243
rect 416 2076 443 2083
rect 456 2076 463 2113
rect 496 2076 503 2093
rect 516 2087 523 2233
rect 596 2143 603 2213
rect 616 2207 623 2263
rect 596 2136 623 2143
rect 176 1707 183 1773
rect 76 1616 103 1623
rect 36 1596 63 1603
rect 16 863 23 1333
rect 36 1083 43 1596
rect 56 1347 63 1553
rect 96 1427 103 1616
rect 116 1563 123 1653
rect 176 1596 183 1673
rect 196 1667 203 1763
rect 196 1576 203 1633
rect 116 1556 143 1563
rect 76 1316 83 1333
rect 56 1127 63 1303
rect 116 1127 123 1533
rect 116 1083 123 1113
rect 36 1076 63 1083
rect 16 856 43 863
rect 16 383 23 856
rect 56 667 63 1076
rect 96 1076 123 1083
rect 96 647 103 1076
rect 136 1067 143 1556
rect 156 1387 163 1573
rect 216 1407 223 1653
rect 236 1387 243 1693
rect 336 1663 343 1713
rect 316 1656 343 1663
rect 256 1607 263 1613
rect 296 1596 303 1653
rect 276 1387 283 1583
rect 316 1576 323 1656
rect 176 1327 183 1373
rect 236 1336 243 1373
rect 296 1347 303 1553
rect 336 1467 343 1633
rect 356 1583 363 1793
rect 376 1607 383 1803
rect 396 1596 403 2033
rect 416 1847 423 1993
rect 416 1707 423 1833
rect 436 1747 443 2076
rect 476 1967 483 2063
rect 456 1807 463 1953
rect 356 1576 383 1583
rect 356 1443 363 1553
rect 336 1436 363 1443
rect 316 1336 323 1373
rect 336 1367 343 1436
rect 216 1303 223 1333
rect 196 1296 223 1303
rect 176 1227 183 1283
rect 196 1136 203 1253
rect 156 1103 163 1133
rect 216 1107 223 1153
rect 256 1143 263 1323
rect 296 1147 303 1333
rect 336 1316 363 1323
rect 356 1307 363 1316
rect 236 1136 263 1143
rect 156 1096 183 1103
rect 196 887 203 1093
rect 236 967 243 1136
rect 316 1116 323 1173
rect 276 1007 283 1093
rect 296 1027 303 1103
rect 336 947 343 1133
rect 356 987 363 1293
rect 376 883 383 1293
rect 396 1247 403 1553
rect 416 1507 423 1583
rect 436 1487 443 1553
rect 456 1547 463 1693
rect 476 1627 483 1933
rect 496 1603 503 1973
rect 536 1887 543 2113
rect 596 2096 603 2113
rect 556 2076 583 2083
rect 616 2076 623 2136
rect 556 1927 563 2076
rect 636 1847 643 2493
rect 656 2187 663 2243
rect 696 2187 703 2633
rect 756 2576 763 2613
rect 736 2556 743 2573
rect 716 2127 723 2553
rect 796 2547 803 2773
rect 816 2747 823 2763
rect 856 2756 863 2813
rect 876 2787 883 3176
rect 896 3056 903 3153
rect 976 3043 983 3233
rect 1176 3207 1183 3236
rect 996 3187 1003 3203
rect 1136 3056 1143 3073
rect 976 3036 1003 3043
rect 996 3023 1003 3036
rect 916 2967 923 3023
rect 996 3016 1023 3023
rect 916 2827 923 2953
rect 996 2887 1003 3016
rect 1276 2987 1283 3353
rect 1296 3227 1303 3533
rect 1336 3516 1343 3573
rect 1436 3496 1443 3533
rect 1476 3483 1483 3553
rect 1536 3536 1543 3913
rect 1596 3743 1603 3813
rect 1576 3736 1603 3743
rect 1636 3736 1643 3893
rect 1576 3687 1583 3736
rect 1656 3707 1663 3996
rect 1796 3996 1823 4003
rect 1856 3996 1863 4213
rect 1916 4196 1923 4213
rect 1876 4147 1883 4193
rect 1956 4183 1963 4213
rect 1976 4187 1983 4233
rect 1996 4196 2003 4213
rect 1936 4176 1963 4183
rect 2036 4083 2043 4233
rect 2116 4223 2123 4233
rect 2096 4216 2123 4223
rect 2156 4216 2183 4223
rect 2136 4187 2143 4203
rect 2036 4076 2063 4083
rect 1896 3996 1923 4003
rect 1716 3867 1723 3983
rect 1576 3647 1583 3673
rect 1596 3567 1603 3633
rect 1676 3587 1683 3793
rect 1716 3716 1723 3833
rect 1776 3827 1783 3993
rect 1796 3867 1803 3996
rect 1916 3907 1923 3996
rect 1936 3987 1943 4073
rect 1996 3996 2023 4003
rect 1976 3767 1983 3973
rect 2016 3907 2023 3996
rect 2036 3967 2043 4053
rect 2056 4007 2063 4076
rect 2076 3976 2083 4153
rect 2176 4127 2183 4216
rect 2216 4183 2223 4233
rect 2256 4207 2263 4373
rect 2296 4247 2303 4433
rect 2336 4407 2343 4463
rect 2456 4443 2463 4573
rect 2476 4467 2483 4693
rect 2436 4436 2463 4443
rect 2216 4176 2243 4183
rect 2236 4067 2243 4176
rect 2276 4107 2283 4183
rect 2296 4167 2303 4203
rect 2316 4067 2323 4353
rect 2376 4216 2403 4223
rect 2396 4207 2403 4216
rect 2356 4147 2363 4203
rect 2056 3827 2063 3963
rect 1776 3727 1783 3753
rect 2076 3747 2083 3853
rect 2096 3747 2103 3953
rect 2036 3736 2063 3743
rect 1816 3716 1843 3723
rect 1696 3687 1703 3713
rect 1696 3627 1703 3673
rect 1516 3516 1523 3533
rect 1556 3516 1583 3523
rect 1456 3476 1483 3483
rect 1576 3483 1583 3516
rect 1576 3476 1603 3483
rect 1636 3476 1643 3533
rect 1716 3523 1723 3593
rect 1776 3563 1783 3613
rect 1756 3556 1783 3563
rect 1696 3516 1723 3523
rect 1756 3516 1763 3556
rect 1816 3547 1823 3653
rect 1836 3547 1843 3716
rect 1916 3703 1923 3713
rect 1896 3696 1923 3703
rect 1876 3587 1883 3683
rect 1656 3496 1663 3513
rect 1296 3023 1303 3193
rect 1316 3167 1323 3243
rect 1336 3027 1343 3263
rect 1376 3256 1403 3263
rect 1356 3227 1363 3243
rect 1396 3227 1403 3256
rect 1416 3167 1423 3333
rect 1296 3016 1323 3023
rect 896 2747 903 2813
rect 836 2727 843 2743
rect 876 2687 883 2743
rect 916 2723 923 2793
rect 976 2727 983 2743
rect 916 2716 963 2723
rect 796 2487 803 2533
rect 816 2487 823 2673
rect 876 2556 903 2563
rect 776 2287 783 2303
rect 816 2296 823 2413
rect 756 2247 763 2283
rect 536 1796 563 1803
rect 476 1596 503 1603
rect 476 1587 483 1596
rect 516 1587 523 1693
rect 536 1576 543 1773
rect 556 1767 563 1796
rect 576 1727 583 1793
rect 476 1527 483 1553
rect 416 1147 423 1453
rect 436 1367 443 1453
rect 476 1367 483 1393
rect 436 1336 443 1353
rect 476 1336 483 1353
rect 496 1347 503 1393
rect 456 1287 463 1323
rect 516 1307 523 1513
rect 536 1343 543 1373
rect 556 1367 563 1563
rect 576 1427 583 1593
rect 596 1487 603 1833
rect 616 1623 623 1653
rect 636 1647 643 1783
rect 656 1707 663 2093
rect 776 2076 783 2133
rect 836 2107 843 2313
rect 856 2287 863 2333
rect 896 2327 903 2556
rect 956 2536 963 2653
rect 936 2487 943 2523
rect 976 2507 983 2523
rect 876 2267 883 2313
rect 936 2296 943 2313
rect 916 2267 923 2283
rect 816 2076 843 2083
rect 716 2056 733 2063
rect 756 2047 763 2063
rect 676 1767 683 1873
rect 696 1727 703 2033
rect 756 1887 763 2033
rect 756 1807 763 1833
rect 796 1827 803 2053
rect 836 2007 843 2076
rect 916 2056 923 2073
rect 956 2067 963 2453
rect 976 2327 983 2493
rect 996 2327 1003 2753
rect 1096 2747 1103 2763
rect 1116 2747 1123 2783
rect 1016 2487 1023 2713
rect 1036 2707 1043 2743
rect 1036 2507 1043 2693
rect 1096 2576 1103 2613
rect 1056 2507 1063 2553
rect 1076 2503 1083 2543
rect 1096 2507 1103 2533
rect 1067 2496 1083 2503
rect 1096 2467 1103 2493
rect 1116 2327 1123 2613
rect 1156 2536 1163 2733
rect 1176 2667 1183 2893
rect 1216 2787 1223 2913
rect 1136 2507 1143 2523
rect 1176 2487 1183 2523
rect 976 2147 983 2313
rect 816 1807 823 1873
rect 856 1787 863 2053
rect 876 1847 883 2033
rect 896 2007 903 2043
rect 936 2027 943 2043
rect 976 2027 983 2133
rect 1016 2087 1023 2283
rect 1036 2087 1043 2233
rect 1056 2127 1063 2313
rect 1076 2307 1083 2313
rect 1116 2296 1143 2303
rect 1136 2263 1143 2296
rect 1116 2256 1143 2263
rect 1016 2056 1023 2073
rect 1076 2067 1083 2253
rect 1096 2227 1103 2253
rect 1116 2247 1123 2256
rect 1096 2107 1103 2213
rect 1156 2127 1163 2473
rect 1196 2307 1203 2773
rect 1216 2756 1223 2773
rect 1236 2627 1243 2913
rect 1296 2803 1303 3016
rect 1276 2796 1303 2803
rect 1276 2763 1283 2796
rect 1276 2756 1303 2763
rect 1256 2536 1263 2673
rect 1316 2627 1323 2973
rect 1436 2907 1443 3223
rect 1496 3207 1503 3473
rect 1696 3467 1703 3516
rect 1596 3267 1603 3393
rect 1536 3167 1543 3253
rect 1556 3207 1563 3243
rect 1596 3236 1603 3253
rect 1576 3187 1583 3223
rect 1616 3187 1623 3223
rect 1456 2867 1463 3093
rect 1476 2927 1483 3133
rect 1496 3016 1503 3053
rect 1516 3036 1523 3073
rect 1556 3036 1563 3113
rect 1336 2667 1343 2773
rect 1476 2767 1483 2893
rect 1536 2887 1543 3023
rect 1576 2887 1583 3153
rect 1636 3087 1643 3353
rect 1676 3236 1683 3353
rect 1656 3107 1663 3213
rect 1696 3207 1703 3223
rect 1596 3007 1603 3073
rect 1656 3063 1663 3093
rect 1716 3067 1723 3233
rect 1736 3187 1743 3253
rect 1756 3227 1763 3313
rect 1756 3147 1763 3193
rect 1776 3107 1783 3533
rect 1816 3516 1833 3523
rect 1876 3516 1883 3553
rect 1976 3527 1983 3723
rect 2016 3687 2023 3723
rect 2056 3707 2063 3736
rect 2116 3727 2123 4033
rect 2136 4016 2143 4033
rect 2216 3996 2243 4003
rect 2276 3996 2283 4013
rect 2296 4007 2303 4053
rect 2316 4047 2323 4053
rect 2216 3867 2223 3996
rect 2296 3976 2303 3993
rect 2256 3847 2263 3973
rect 2316 3963 2323 4013
rect 2356 3976 2363 3993
rect 2316 3956 2343 3963
rect 2156 3736 2183 3743
rect 2156 3703 2163 3736
rect 2216 3727 2223 3743
rect 2136 3696 2163 3703
rect 2196 3687 2203 3723
rect 2236 3707 2243 3723
rect 1896 3516 1943 3523
rect 1836 3463 1843 3513
rect 1896 3483 1903 3516
rect 1856 3476 1903 3483
rect 1936 3476 1943 3516
rect 1956 3496 1963 3513
rect 1996 3483 2003 3593
rect 1976 3476 2003 3483
rect 1836 3456 1863 3463
rect 1836 3167 1843 3213
rect 1836 3123 1843 3153
rect 1816 3116 1843 3123
rect 1656 3056 1683 3063
rect 1636 3036 1643 3053
rect 1676 3036 1683 3056
rect 1756 3056 1763 3073
rect 1716 3036 1743 3043
rect 1776 3036 1783 3053
rect 1616 3027 1623 3033
rect 1656 3007 1663 3023
rect 1656 2927 1663 2993
rect 1636 2776 1643 2793
rect 1656 2747 1663 2853
rect 1296 2587 1303 2593
rect 1236 2507 1243 2523
rect 1176 2227 1183 2263
rect 1196 2203 1203 2233
rect 1176 2196 1203 2203
rect 996 2027 1003 2043
rect 1076 1987 1083 2033
rect 1096 2027 1103 2073
rect 716 1776 743 1783
rect 616 1616 643 1623
rect 676 1596 683 1693
rect 616 1467 623 1583
rect 636 1447 643 1573
rect 536 1336 563 1343
rect 596 1336 603 1353
rect 436 1123 443 1213
rect 456 1127 463 1133
rect 416 1116 443 1123
rect 416 1096 423 1116
rect 436 1087 443 1093
rect 396 1047 403 1083
rect 356 876 383 883
rect 176 796 203 803
rect 136 627 143 633
rect 176 616 183 796
rect 136 603 143 613
rect 76 567 83 603
rect 116 596 143 603
rect 216 603 223 633
rect 276 616 283 633
rect 196 596 223 603
rect 296 547 303 603
rect 316 507 323 733
rect 336 607 343 853
rect 356 843 363 876
rect 356 836 383 843
rect 356 727 363 773
rect 376 747 383 836
rect 396 787 403 973
rect 416 807 423 1053
rect 456 883 463 1053
rect 436 876 463 883
rect 356 603 363 713
rect 436 667 443 876
rect 456 836 463 853
rect 476 827 483 1233
rect 496 1147 503 1273
rect 536 1267 543 1336
rect 556 1183 563 1293
rect 576 1207 583 1323
rect 616 1267 623 1303
rect 636 1267 643 1413
rect 656 1387 663 1583
rect 696 1567 703 1673
rect 716 1667 723 1776
rect 756 1727 763 1763
rect 716 1607 723 1633
rect 736 1596 743 1633
rect 756 1616 763 1653
rect 776 1596 783 1753
rect 796 1707 803 1783
rect 836 1727 843 1783
rect 876 1727 883 1833
rect 936 1816 943 1953
rect 896 1707 903 1813
rect 976 1807 983 1823
rect 956 1783 963 1793
rect 996 1787 1003 1803
rect 936 1776 963 1783
rect 936 1767 943 1776
rect 896 1687 903 1693
rect 656 1336 663 1353
rect 696 1327 703 1513
rect 616 1247 623 1253
rect 636 1227 643 1253
rect 676 1227 683 1303
rect 716 1287 723 1573
rect 796 1547 803 1633
rect 756 1267 763 1343
rect 776 1307 783 1323
rect 556 1176 583 1183
rect 496 1027 503 1073
rect 516 983 523 1053
rect 536 1047 543 1073
rect 556 1047 563 1093
rect 516 976 543 983
rect 496 867 503 933
rect 516 847 523 953
rect 396 647 403 653
rect 396 616 403 633
rect 436 616 443 653
rect 456 647 463 733
rect 496 636 503 793
rect 536 707 543 976
rect 576 887 583 1176
rect 596 1087 603 1133
rect 616 1083 623 1153
rect 656 1107 663 1133
rect 716 1096 723 1153
rect 736 1107 743 1253
rect 756 1096 763 1213
rect 616 1076 643 1083
rect 596 1027 603 1073
rect 556 856 563 873
rect 596 856 603 953
rect 576 807 583 843
rect 356 596 383 603
rect 416 596 423 613
rect 476 567 483 623
rect 516 616 523 633
rect 536 627 543 673
rect 556 636 563 793
rect 576 656 583 673
rect 596 636 623 643
rect 16 376 43 383
rect 16 123 23 376
rect 16 116 43 123
rect 36 67 43 116
rect 356 107 363 533
rect 396 363 403 493
rect 476 407 483 553
rect 376 356 403 363
rect 456 356 463 373
rect 496 367 503 473
rect 576 367 583 393
rect 376 136 383 356
rect 516 156 523 353
rect 536 347 543 363
rect 556 327 563 343
rect 596 327 603 343
rect 616 247 623 636
rect 456 127 463 143
rect 496 107 503 143
rect 576 127 583 213
rect 636 207 643 693
rect 656 447 663 993
rect 696 847 703 1053
rect 716 907 723 1053
rect 696 663 703 803
rect 736 787 743 973
rect 756 947 763 1053
rect 776 987 783 1083
rect 796 967 803 1253
rect 816 1227 823 1673
rect 836 1596 863 1603
rect 896 1596 903 1633
rect 916 1603 923 1713
rect 936 1627 943 1633
rect 916 1596 943 1603
rect 836 1587 843 1596
rect 876 1567 883 1583
rect 836 1507 843 1553
rect 836 1203 843 1493
rect 916 1367 923 1513
rect 936 1507 943 1596
rect 856 1336 863 1353
rect 936 1307 943 1333
rect 956 1287 963 1753
rect 1016 1747 1023 1803
rect 1036 1796 1063 1803
rect 1036 1747 1043 1796
rect 1096 1787 1103 1953
rect 1116 1867 1123 2113
rect 1176 2103 1183 2196
rect 1216 2167 1223 2243
rect 1256 2183 1263 2473
rect 1296 2303 1303 2573
rect 1316 2427 1323 2593
rect 1356 2556 1363 2593
rect 1356 2427 1363 2513
rect 1276 2296 1303 2303
rect 1276 2263 1283 2296
rect 1316 2276 1323 2373
rect 1276 2256 1303 2263
rect 1276 2207 1283 2233
rect 1236 2176 1263 2183
rect 1156 2096 1183 2103
rect 1156 2076 1163 2096
rect 1236 2103 1243 2176
rect 1216 2096 1243 2103
rect 1196 2076 1203 2093
rect 1136 2056 1143 2073
rect 996 1616 1003 1633
rect 976 1596 983 1613
rect 1016 1596 1023 1673
rect 996 1487 1003 1573
rect 1036 1343 1043 1633
rect 1056 1547 1063 1773
rect 1116 1687 1123 1833
rect 1136 1727 1143 1913
rect 1076 1603 1083 1653
rect 1096 1627 1103 1653
rect 1076 1596 1103 1603
rect 1136 1596 1143 1633
rect 1036 1336 1063 1343
rect 976 1307 983 1323
rect 1056 1303 1063 1336
rect 1076 1327 1083 1553
rect 1156 1523 1163 1993
rect 1176 1967 1183 2053
rect 1216 1947 1223 2096
rect 1256 2027 1263 2063
rect 1276 2007 1283 2193
rect 1296 2147 1303 2233
rect 1356 2207 1363 2283
rect 1296 1927 1303 2113
rect 1376 2107 1383 2653
rect 1436 2523 1443 2653
rect 1436 2516 1463 2523
rect 1396 2247 1403 2333
rect 1456 2227 1463 2263
rect 1476 2247 1483 2393
rect 1496 2267 1503 2523
rect 1516 2407 1523 2593
rect 1556 2576 1563 2593
rect 1596 2556 1603 2593
rect 1516 2227 1523 2263
rect 1556 2247 1563 2263
rect 1576 2147 1583 2283
rect 1596 2247 1603 2513
rect 1636 2467 1643 2673
rect 1676 2643 1683 2893
rect 1696 2827 1703 3033
rect 1716 2967 1723 3036
rect 1716 2756 1723 2913
rect 1736 2687 1743 2743
rect 1756 2727 1763 2753
rect 1656 2636 1683 2643
rect 1656 2536 1663 2636
rect 1676 2556 1683 2613
rect 1696 2527 1703 2543
rect 1616 2276 1643 2283
rect 1616 2207 1623 2276
rect 1696 2247 1703 2263
rect 1656 2187 1663 2243
rect 1716 2187 1723 2273
rect 1736 2143 1743 2453
rect 1756 2247 1763 2693
rect 1776 2687 1783 2753
rect 1776 2563 1783 2633
rect 1796 2587 1803 3053
rect 1816 3036 1823 3116
rect 1816 2707 1823 2953
rect 1836 2807 1843 3093
rect 1856 3087 1863 3456
rect 1876 3207 1883 3476
rect 2016 3467 2023 3493
rect 1876 3036 1883 3073
rect 1856 2787 1863 2993
rect 1876 2756 1883 2873
rect 1896 2847 1903 3453
rect 2036 3447 2043 3573
rect 2056 3523 2063 3673
rect 2116 3587 2123 3683
rect 2196 3587 2203 3613
rect 2176 3527 2183 3573
rect 2056 3516 2083 3523
rect 2116 3516 2143 3523
rect 1936 3247 1943 3273
rect 1916 3167 1923 3223
rect 1956 3207 1963 3223
rect 1916 3047 1923 3153
rect 1976 3147 1983 3433
rect 2076 3363 2083 3516
rect 2136 3487 2143 3516
rect 2156 3503 2163 3513
rect 2156 3496 2183 3503
rect 2216 3496 2223 3553
rect 2096 3476 2123 3483
rect 2116 3467 2123 3476
rect 2156 3467 2163 3496
rect 2256 3483 2263 3813
rect 2276 3727 2283 3833
rect 2356 3707 2363 3733
rect 2376 3707 2383 3953
rect 2336 3687 2343 3703
rect 2376 3647 2383 3693
rect 2396 3627 2403 4173
rect 2416 4147 2423 4313
rect 2436 4187 2443 4436
rect 2496 4347 2503 4493
rect 2516 4287 2523 4683
rect 2556 4667 2563 4796
rect 2576 4696 2583 4916
rect 2636 4887 2643 4943
rect 2676 4923 2683 5013
rect 2716 4936 2723 5033
rect 2676 4916 2703 4923
rect 2736 4916 2743 5033
rect 2776 4983 2783 5153
rect 2816 5047 2823 5143
rect 2916 5143 2923 5176
rect 2916 5136 2943 5143
rect 2756 4976 2783 4983
rect 2796 4976 2803 5013
rect 2756 4936 2763 4976
rect 2836 4956 2863 4963
rect 2816 4927 2823 4943
rect 2556 4507 2563 4633
rect 2576 4487 2583 4633
rect 2596 4627 2603 4683
rect 2616 4527 2623 4673
rect 2656 4663 2663 4913
rect 2856 4707 2863 4956
rect 2896 4947 2903 5073
rect 2936 5007 2943 5136
rect 2956 5123 2963 5163
rect 2996 5127 3003 5176
rect 3036 5176 3043 5193
rect 3076 5176 3083 5213
rect 2956 5116 2973 5123
rect 3016 5023 3023 5173
rect 3056 5147 3063 5163
rect 3096 5147 3103 5353
rect 3016 5016 3043 5023
rect 2936 4943 2943 4993
rect 2976 4976 3003 4983
rect 2916 4936 2943 4943
rect 2687 4676 2703 4683
rect 2796 4683 2803 4693
rect 2796 4676 2823 4683
rect 2636 4656 2663 4663
rect 2596 4487 2603 4513
rect 2536 4327 2543 4443
rect 2576 4436 2583 4473
rect 2616 4367 2623 4513
rect 2467 4216 2483 4223
rect 2516 4216 2523 4233
rect 2456 4167 2463 4213
rect 2496 4187 2503 4203
rect 2536 4187 2543 4293
rect 2556 4167 2563 4183
rect 2576 4156 2593 4163
rect 2416 3687 2423 4053
rect 2436 4047 2443 4153
rect 2436 3787 2443 4033
rect 2456 3996 2463 4093
rect 2516 3987 2523 4153
rect 2536 4016 2543 4133
rect 2576 3963 2583 4053
rect 2556 3956 2583 3963
rect 2436 3727 2443 3773
rect 2476 3747 2483 3793
rect 2556 3736 2563 3956
rect 2236 3476 2263 3483
rect 2076 3356 2103 3363
rect 2036 3263 2043 3333
rect 2016 3256 2043 3263
rect 1956 3123 1963 3133
rect 1956 3116 1983 3123
rect 1936 3016 1943 3053
rect 1976 3027 1983 3116
rect 1996 3067 2003 3223
rect 2016 3007 2023 3256
rect 2056 3187 2063 3223
rect 1996 2987 2003 3003
rect 2036 2947 2043 3133
rect 2056 3007 2063 3053
rect 2076 3016 2083 3153
rect 2096 3047 2103 3356
rect 2116 3227 2123 3453
rect 2176 3247 2183 3263
rect 2156 3227 2163 3243
rect 2116 3147 2123 3193
rect 2116 3016 2123 3073
rect 2136 3047 2143 3173
rect 2156 3047 2163 3213
rect 2096 2996 2103 3013
rect 2056 2947 2063 2973
rect 1936 2767 1943 2913
rect 1836 2667 1843 2693
rect 1776 2556 1803 2563
rect 1876 2556 1883 2613
rect 1716 2136 1743 2143
rect 1496 2107 1503 2133
rect 1516 2116 1643 2123
rect 1416 2076 1443 2083
rect 1176 1847 1183 1913
rect 1196 1816 1203 1873
rect 1176 1747 1183 1783
rect 1216 1687 1223 1813
rect 1256 1647 1263 1853
rect 1316 1847 1323 2073
rect 1356 2027 1363 2063
rect 1276 1816 1303 1823
rect 1336 1816 1343 1873
rect 1276 1767 1283 1816
rect 1316 1787 1323 1793
rect 1176 1616 1183 1633
rect 1216 1567 1223 1613
rect 1236 1596 1263 1603
rect 1296 1596 1303 1613
rect 1236 1587 1243 1596
rect 1156 1516 1183 1523
rect 976 1287 983 1293
rect 816 1196 843 1203
rect 816 1007 823 1196
rect 856 1107 863 1273
rect 996 1267 1003 1303
rect 1036 1296 1063 1303
rect 1096 1287 1103 1323
rect 836 1027 843 1073
rect 876 1063 883 1083
rect 856 1056 883 1063
rect 856 1047 863 1056
rect 896 1047 903 1253
rect 916 1107 923 1213
rect 976 1147 983 1153
rect 956 1096 963 1133
rect 796 836 803 873
rect 676 656 703 663
rect 676 636 683 656
rect 756 627 763 813
rect 656 407 663 413
rect 656 376 663 393
rect 696 376 703 393
rect 676 347 683 363
rect 716 287 723 593
rect 736 376 743 433
rect 776 387 783 813
rect 816 807 823 823
rect 836 687 843 843
rect 856 807 863 1033
rect 876 663 883 953
rect 916 836 923 873
rect 936 807 943 823
rect 956 787 963 843
rect 976 707 983 1053
rect 996 787 1003 1233
rect 1076 1116 1083 1153
rect 1016 1087 1023 1103
rect 1056 1087 1063 1103
rect 1096 1087 1103 1193
rect 1116 1127 1123 1253
rect 1156 1116 1163 1213
rect 1176 1147 1183 1516
rect 1196 1323 1203 1353
rect 1236 1347 1243 1573
rect 1276 1367 1283 1583
rect 1316 1576 1323 1593
rect 1336 1527 1343 1633
rect 1196 1316 1223 1323
rect 1256 1316 1263 1353
rect 1196 1187 1203 1293
rect 1236 1127 1243 1303
rect 1296 1267 1303 1493
rect 1336 1316 1343 1353
rect 1356 1247 1363 1973
rect 1376 1783 1383 1993
rect 1396 1987 1403 2063
rect 1436 1967 1443 2076
rect 1436 1827 1443 1953
rect 1456 1807 1463 2093
rect 1476 2076 1483 2093
rect 1516 2076 1523 2116
rect 1636 2096 1643 2116
rect 1556 2076 1583 2083
rect 1496 2027 1503 2063
rect 1536 1887 1543 2053
rect 1576 1967 1583 2076
rect 1596 2063 1603 2093
rect 1676 2076 1703 2083
rect 1596 2056 1623 2063
rect 1596 1943 1603 2033
rect 1576 1936 1603 1943
rect 1556 1887 1563 1913
rect 1476 1807 1483 1833
rect 1556 1787 1563 1803
rect 1376 1776 1403 1783
rect 1487 1776 1503 1783
rect 1476 1763 1483 1773
rect 1536 1767 1543 1783
rect 1576 1767 1583 1936
rect 1596 1816 1623 1823
rect 1656 1816 1663 1933
rect 1596 1807 1603 1816
rect 1436 1667 1443 1763
rect 1456 1756 1483 1763
rect 1276 1136 1283 1153
rect 1376 1147 1383 1513
rect 1396 1303 1403 1613
rect 1436 1596 1443 1613
rect 1416 1347 1423 1533
rect 1456 1387 1463 1756
rect 1476 1487 1483 1713
rect 1596 1667 1603 1793
rect 1516 1576 1523 1593
rect 1496 1527 1503 1553
rect 1436 1316 1443 1333
rect 1516 1307 1523 1353
rect 1396 1296 1423 1303
rect 1316 1116 1343 1123
rect 1036 1063 1043 1073
rect 1036 1056 1063 1063
rect 856 656 883 663
rect 876 647 883 656
rect 896 636 903 693
rect 936 636 983 643
rect 836 447 843 623
rect 756 307 763 363
rect 796 343 803 433
rect 876 343 883 373
rect 796 336 823 343
rect 856 336 883 343
rect 716 156 723 173
rect 776 156 783 193
rect 836 187 843 323
rect 856 227 863 336
rect 896 307 903 553
rect 916 327 923 613
rect 976 407 983 636
rect 996 387 1003 693
rect 1016 687 1023 993
rect 1036 847 1043 953
rect 1056 856 1063 1056
rect 1116 887 1123 1093
rect 1076 807 1083 843
rect 1096 767 1103 853
rect 1136 827 1143 1093
rect 1176 1067 1183 1103
rect 1216 1096 1243 1103
rect 1236 1087 1243 1096
rect 1196 1027 1203 1073
rect 1256 1047 1263 1103
rect 1176 847 1183 873
rect 1216 836 1243 843
rect 1156 787 1163 823
rect 1236 807 1243 836
rect 1256 827 1263 1013
rect 1016 347 1023 673
rect 1036 636 1043 653
rect 1076 636 1083 693
rect 1096 647 1103 673
rect 1096 616 1103 633
rect 1116 627 1123 773
rect 1196 767 1203 803
rect 1276 787 1283 1053
rect 1296 947 1303 1073
rect 1336 947 1343 1116
rect 1396 1116 1403 1213
rect 1416 1096 1423 1193
rect 1376 987 1383 1093
rect 1436 1007 1443 1273
rect 1456 987 1463 1303
rect 1496 1296 1513 1303
rect 1496 1136 1503 1233
rect 1516 1116 1523 1173
rect 1536 1063 1543 1393
rect 1556 1367 1563 1633
rect 1636 1603 1643 1803
rect 1676 1647 1683 2033
rect 1696 1927 1703 2076
rect 1716 2007 1723 2136
rect 1776 2127 1783 2313
rect 1816 2287 1823 2543
rect 1856 2347 1863 2543
rect 1896 2327 1903 2653
rect 1956 2536 1963 2933
rect 1976 2667 1983 2813
rect 1996 2707 2003 2833
rect 2036 2807 2043 2873
rect 2076 2843 2083 2973
rect 2076 2836 2103 2843
rect 2036 2647 2043 2753
rect 2056 2727 2063 2783
rect 2096 2763 2103 2836
rect 2076 2756 2103 2763
rect 2016 2567 2023 2613
rect 2116 2607 2123 2933
rect 2156 2887 2163 3033
rect 2176 3007 2183 3073
rect 2196 3067 2203 3243
rect 2216 3043 2223 3413
rect 2296 3367 2303 3613
rect 2316 3483 2323 3513
rect 2356 3496 2363 3553
rect 2396 3536 2403 3553
rect 2416 3516 2423 3593
rect 2316 3476 2343 3483
rect 2396 3223 2403 3253
rect 2316 3207 2323 3223
rect 2356 3216 2403 3223
rect 2236 3187 2243 3203
rect 2196 3036 2223 3043
rect 2136 2747 2143 2763
rect 2176 2756 2183 2853
rect 2196 2787 2203 3036
rect 2236 3016 2243 3153
rect 2216 2807 2223 2973
rect 2276 2927 2283 3193
rect 2416 3147 2423 3233
rect 2316 3016 2323 3033
rect 2336 2996 2343 3033
rect 2356 3016 2363 3053
rect 2376 3007 2383 3113
rect 2416 3067 2423 3133
rect 2436 3087 2443 3573
rect 2456 3567 2463 3673
rect 2456 3447 2463 3503
rect 2476 3463 2483 3513
rect 2496 3487 2503 3693
rect 2476 3456 2503 3463
rect 2216 2776 2243 2783
rect 2276 2776 2283 2853
rect 2216 2743 2223 2776
rect 2296 2747 2303 2913
rect 2316 2827 2323 2933
rect 2396 2887 2403 3053
rect 2416 3036 2423 3053
rect 2476 3016 2483 3033
rect 2436 2987 2443 3013
rect 2336 2747 2343 2783
rect 2156 2727 2163 2743
rect 2196 2736 2223 2743
rect 2196 2707 2203 2736
rect 2356 2743 2363 2763
rect 2356 2736 2383 2743
rect 2276 2727 2283 2733
rect 1996 2487 2003 2543
rect 2136 2543 2143 2693
rect 2176 2567 2183 2613
rect 2196 2547 2203 2693
rect 2256 2576 2263 2593
rect 2216 2556 2243 2563
rect 2276 2556 2283 2713
rect 2356 2556 2363 2653
rect 2376 2576 2383 2736
rect 2396 2567 2403 2793
rect 2136 2536 2163 2543
rect 2156 2527 2163 2536
rect 2176 2447 2183 2453
rect 1916 2296 1943 2303
rect 1996 2296 2023 2303
rect 1936 2287 1943 2296
rect 2016 2287 2023 2296
rect 2056 2287 2063 2293
rect 2096 2276 2103 2293
rect 1936 2263 1943 2273
rect 2056 2263 2063 2273
rect 1736 2076 1743 2113
rect 1796 2107 1803 2263
rect 1836 2247 1843 2263
rect 1916 2256 1943 2263
rect 1816 2076 1823 2113
rect 1696 1847 1703 1893
rect 1696 1747 1703 1833
rect 1716 1823 1723 1993
rect 1756 1967 1763 2063
rect 1716 1816 1743 1823
rect 1756 1647 1763 1803
rect 1796 1727 1803 2063
rect 1836 1847 1843 2093
rect 1856 2047 1863 2213
rect 1916 2096 1923 2256
rect 1976 2207 1983 2263
rect 2036 2256 2063 2263
rect 2076 2243 2083 2263
rect 2076 2236 2103 2243
rect 1876 2076 1903 2083
rect 1936 2076 1943 2133
rect 1956 2076 1983 2083
rect 2016 2076 2023 2133
rect 1856 1887 1863 1893
rect 1856 1816 1863 1873
rect 1876 1787 1883 2076
rect 1956 2043 1963 2076
rect 1956 2036 1983 2043
rect 1896 1807 1903 2033
rect 1956 1816 1963 1853
rect 1636 1596 1663 1603
rect 1576 1327 1583 1593
rect 1616 1576 1623 1593
rect 1596 1547 1603 1563
rect 1636 1547 1643 1563
rect 1656 1367 1663 1596
rect 1676 1363 1683 1593
rect 1696 1567 1703 1633
rect 1716 1576 1723 1613
rect 1756 1567 1763 1583
rect 1796 1407 1803 1653
rect 1816 1616 1823 1773
rect 1836 1627 1843 1773
rect 1676 1356 1703 1363
rect 1596 1347 1603 1353
rect 1596 1283 1603 1313
rect 1616 1307 1623 1323
rect 1636 1307 1643 1343
rect 1696 1307 1703 1356
rect 1576 1276 1603 1283
rect 1556 1136 1563 1173
rect 1576 1087 1583 1103
rect 1596 1063 1603 1133
rect 1536 1056 1563 1063
rect 1296 856 1303 933
rect 1316 807 1323 843
rect 1336 823 1343 853
rect 1336 816 1363 823
rect 1236 667 1243 713
rect 1236 627 1243 653
rect 1336 647 1343 753
rect 1356 727 1363 816
rect 1287 636 1303 643
rect 1256 616 1283 623
rect 1196 603 1203 613
rect 1176 596 1203 603
rect 1036 376 1043 593
rect 1176 367 1183 596
rect 1256 447 1263 616
rect 1276 567 1283 573
rect 1056 347 1063 363
rect 936 307 943 343
rect 1096 327 1103 363
rect 1136 356 1163 363
rect 1156 347 1163 356
rect 1196 347 1203 433
rect 1216 327 1223 343
rect 856 207 863 213
rect 936 187 943 293
rect 956 267 963 323
rect 816 156 833 163
rect 916 156 923 173
rect 616 136 623 153
rect 696 136 703 153
rect 587 116 603 123
rect 636 107 643 113
rect 676 27 683 133
rect 736 87 743 143
rect 796 107 803 143
rect 856 127 863 153
rect 876 87 883 153
rect 976 143 983 313
rect 1116 267 1123 323
rect 1156 267 1163 313
rect 1116 247 1123 253
rect 1116 147 1123 213
rect 1156 176 1163 253
rect 1236 187 1243 323
rect 976 136 1003 143
rect 996 107 1003 136
rect 1276 136 1283 473
rect 1356 367 1363 713
rect 1376 627 1383 893
rect 1396 856 1423 863
rect 1396 807 1403 856
rect 1436 827 1443 833
rect 1496 827 1503 863
rect 1536 856 1543 993
rect 1456 636 1463 813
rect 1516 707 1523 843
rect 1556 687 1563 1056
rect 1576 1056 1603 1063
rect 1576 747 1583 1056
rect 1616 887 1623 1113
rect 1636 1083 1643 1153
rect 1676 1096 1683 1153
rect 1636 1076 1663 1083
rect 1656 867 1663 1013
rect 1716 887 1723 1373
rect 1736 1303 1743 1333
rect 1736 1296 1763 1303
rect 1776 1207 1783 1283
rect 1816 1187 1823 1573
rect 1836 1547 1843 1583
rect 1776 1136 1783 1173
rect 1736 907 1743 1133
rect 1836 1123 1843 1473
rect 1856 1467 1863 1613
rect 1876 1587 1883 1733
rect 1916 1603 1923 1773
rect 1936 1627 1943 1773
rect 1916 1596 1943 1603
rect 1896 1563 1903 1593
rect 1936 1576 1943 1596
rect 1976 1563 1983 2036
rect 2036 2027 2043 2113
rect 1996 1796 2003 1853
rect 2016 1807 2023 1873
rect 2036 1796 2043 1973
rect 2056 1823 2063 2113
rect 2076 2067 2083 2093
rect 2096 2076 2103 2236
rect 2116 2187 2123 2263
rect 2136 2167 2143 2283
rect 2156 2187 2163 2293
rect 2176 2127 2183 2433
rect 2216 2387 2223 2556
rect 2416 2547 2423 2893
rect 2436 2787 2443 2853
rect 2496 2847 2503 3456
rect 2516 3107 2523 3713
rect 2536 3707 2543 3723
rect 2576 3567 2583 3733
rect 2596 3587 2603 4013
rect 2616 3747 2623 4273
rect 2636 3747 2643 4656
rect 2676 4643 2683 4673
rect 2656 4636 2683 4643
rect 2656 4476 2663 4636
rect 2716 4607 2723 4643
rect 2776 4627 2783 4673
rect 2836 4627 2843 4663
rect 2876 4607 2883 4663
rect 2696 4496 2703 4513
rect 2676 4247 2683 4463
rect 2656 4216 2673 4223
rect 2656 4027 2663 4216
rect 2716 4216 2723 4233
rect 2696 4187 2703 4203
rect 2736 4183 2743 4533
rect 2756 4467 2763 4553
rect 2756 4187 2763 4233
rect 2776 4196 2783 4573
rect 2876 4527 2883 4593
rect 2896 4587 2903 4733
rect 2996 4727 3003 4976
rect 3016 4767 3023 4993
rect 3036 4967 3043 5016
rect 3056 4956 3063 5113
rect 3116 5087 3123 5436
rect 3156 5407 3163 5423
rect 3196 5387 3203 5423
rect 3236 5403 3243 5433
rect 3236 5396 3263 5403
rect 3296 5387 3303 5403
rect 3296 5367 3303 5373
rect 3136 5103 3143 5143
rect 3136 5096 3163 5103
rect 3096 4956 3103 4993
rect 3116 4987 3123 5053
rect 3036 4936 3043 4953
rect 3016 4747 3023 4753
rect 2916 4696 2923 4713
rect 2916 4487 2923 4653
rect 2936 4567 2943 4673
rect 2976 4667 2983 4713
rect 3016 4696 3023 4733
rect 3076 4707 3083 4943
rect 3136 4907 3143 4943
rect 2796 4447 2803 4463
rect 2716 4176 2743 4183
rect 2716 4047 2723 4176
rect 2816 4163 2823 4253
rect 2796 4156 2823 4163
rect 2676 4016 2703 4023
rect 2696 3947 2703 4016
rect 2736 3987 2743 4073
rect 2756 3956 2763 3993
rect 2776 3987 2783 4113
rect 2836 4027 2843 4233
rect 2856 4216 2863 4473
rect 2936 4443 2943 4513
rect 2956 4476 2963 4653
rect 2976 4527 2983 4653
rect 2916 4436 2943 4443
rect 2976 4247 2983 4473
rect 2896 4216 2923 4223
rect 2856 3996 2863 4173
rect 2876 4167 2883 4203
rect 2916 4187 2923 4216
rect 2796 3907 2803 3993
rect 2836 3967 2843 3983
rect 2876 3976 2883 4013
rect 2836 3947 2843 3953
rect 2896 3887 2903 3993
rect 2936 3827 2943 4233
rect 2996 4227 3003 4613
rect 3016 4456 3023 4513
rect 3076 4476 3083 4553
rect 3096 4267 3103 4713
rect 3136 4676 3143 4693
rect 3116 4627 3123 4643
rect 3156 4607 3163 5096
rect 3176 5007 3183 5143
rect 3176 4587 3183 4933
rect 3196 4923 3203 5013
rect 3196 4916 3223 4923
rect 3196 4667 3203 4733
rect 3216 4696 3223 4713
rect 3236 4667 3243 4683
rect 3116 4476 3123 4533
rect 3156 4476 3163 4513
rect 3196 4476 3203 4533
rect 3216 4507 3223 4513
rect 3276 4507 3283 5333
rect 3316 5327 3323 5513
rect 3356 5436 3363 5473
rect 3396 5207 3403 5473
rect 3416 5436 3423 5453
rect 3436 5436 3463 5443
rect 3496 5436 3503 5473
rect 5256 5467 5263 5473
rect 3856 5456 3883 5463
rect 3536 5436 3563 5443
rect 3436 5227 3443 5436
rect 3396 5156 3403 5173
rect 3336 5107 3343 5143
rect 3436 5143 3443 5213
rect 3416 5136 3443 5143
rect 3456 5107 3463 5393
rect 3476 5187 3483 5413
rect 3516 5387 3523 5423
rect 3556 5367 3563 5436
rect 3596 5416 3603 5453
rect 3656 5436 3683 5443
rect 3636 5407 3643 5423
rect 3536 5147 3543 5163
rect 3516 5027 3523 5143
rect 3556 5127 3563 5353
rect 3616 5156 3623 5373
rect 3676 5367 3683 5436
rect 3736 5436 3743 5453
rect 3716 5367 3723 5423
rect 3756 5416 3783 5423
rect 3776 5387 3783 5416
rect 3876 5403 3883 5456
rect 3956 5456 3983 5463
rect 3956 5403 3963 5456
rect 3876 5396 3903 5403
rect 3936 5396 3963 5403
rect 3716 5243 3723 5353
rect 3696 5236 3723 5243
rect 3696 5167 3703 5236
rect 3816 5156 3823 5173
rect 3576 5067 3583 5153
rect 3596 5127 3603 5143
rect 3676 5107 3683 5113
rect 3296 4956 3323 4963
rect 3296 4927 3303 4956
rect 3396 4947 3403 4993
rect 3436 4976 3443 4993
rect 3456 4956 3483 4963
rect 3376 4907 3383 4943
rect 3296 4627 3303 4693
rect 3136 4327 3143 4463
rect 3176 4447 3183 4463
rect 3016 4196 3043 4203
rect 2956 3987 2963 4093
rect 2996 4087 3003 4163
rect 3036 4107 3043 4196
rect 3076 4167 3083 4183
rect 3036 3987 3043 4073
rect 3076 3967 3083 4073
rect 3096 4023 3103 4213
rect 3116 4196 3123 4233
rect 3096 4016 3123 4023
rect 3136 4016 3143 4153
rect 3156 4023 3163 4353
rect 3176 4196 3183 4213
rect 3196 4187 3203 4313
rect 3216 4023 3223 4493
rect 3236 4476 3263 4483
rect 3296 4476 3303 4553
rect 3316 4507 3323 4753
rect 3336 4647 3343 4893
rect 3356 4696 3363 4833
rect 3336 4476 3343 4633
rect 3376 4627 3383 4683
rect 3396 4667 3403 4703
rect 3236 4447 3243 4476
rect 3316 4447 3323 4463
rect 3236 4167 3243 4233
rect 3156 4016 3183 4023
rect 2996 3867 3003 3953
rect 3016 3887 3023 3963
rect 3096 3947 3103 3993
rect 2616 3716 2643 3723
rect 2536 3507 2543 3553
rect 2556 3516 2563 3533
rect 2596 3256 2603 3493
rect 2616 3487 2623 3503
rect 2616 3467 2623 3473
rect 2616 3287 2623 3413
rect 2636 3347 2643 3716
rect 2676 3687 2683 3793
rect 2696 3647 2703 3723
rect 2696 3516 2703 3533
rect 2776 3516 2783 3553
rect 2676 3407 2683 3503
rect 2716 3496 2723 3513
rect 2756 3467 2763 3473
rect 2536 3187 2543 3243
rect 2536 3167 2543 3173
rect 2556 3056 2563 3233
rect 2576 3227 2583 3243
rect 2616 3207 2623 3273
rect 2636 3247 2643 3333
rect 2656 3227 2663 3293
rect 2716 3287 2723 3353
rect 2716 3236 2723 3273
rect 2516 2827 2523 3053
rect 2576 3047 2583 3153
rect 2536 2987 2543 3023
rect 2536 2867 2543 2973
rect 2576 2967 2583 3013
rect 2596 2907 2603 3073
rect 2616 3067 2623 3113
rect 2636 3067 2643 3093
rect 2656 3056 2663 3113
rect 2456 2707 2463 2763
rect 2476 2556 2483 2653
rect 2496 2607 2503 2763
rect 2536 2723 2543 2833
rect 2616 2807 2623 3053
rect 2676 3036 2683 3133
rect 2696 2803 2703 3073
rect 2716 3036 2723 3133
rect 2736 3027 2743 3153
rect 2756 3147 2763 3453
rect 2776 3223 2783 3353
rect 2796 3287 2803 3503
rect 2836 3236 2843 3393
rect 2856 3327 2863 3553
rect 2876 3367 2883 3683
rect 2896 3427 2903 3493
rect 2936 3403 2943 3613
rect 2956 3503 2963 3633
rect 2976 3527 2983 3813
rect 3016 3736 3043 3743
rect 3016 3667 3023 3736
rect 2956 3496 2983 3503
rect 2956 3427 2963 3496
rect 3016 3467 3023 3653
rect 3056 3627 3063 3933
rect 3096 3716 3103 3893
rect 3116 3607 3123 4016
rect 3136 3947 3143 3973
rect 3136 3727 3143 3833
rect 3156 3687 3163 3873
rect 3176 3767 3183 4016
rect 3196 4016 3223 4023
rect 3236 4016 3243 4033
rect 3196 3763 3203 4016
rect 3256 4007 3263 4433
rect 3276 4227 3283 4273
rect 3336 4247 3343 4433
rect 3356 4287 3363 4553
rect 3376 4367 3383 4573
rect 3396 4503 3403 4593
rect 3416 4587 3423 4673
rect 3436 4527 3443 4933
rect 3476 4927 3483 4956
rect 3396 4496 3443 4503
rect 3376 4243 3383 4333
rect 3396 4247 3403 4496
rect 3416 4447 3423 4463
rect 3436 4447 3443 4453
rect 3456 4247 3463 4653
rect 3356 4236 3383 4243
rect 3296 4216 3303 4233
rect 3276 4007 3283 4213
rect 3316 4187 3323 4203
rect 3216 3967 3223 3983
rect 3296 3976 3303 4073
rect 3316 4047 3323 4173
rect 3356 3983 3363 4236
rect 3416 4216 3423 4233
rect 3476 4227 3483 4913
rect 3556 4883 3563 4943
rect 3556 4876 3583 4883
rect 3496 4627 3503 4663
rect 3496 4507 3503 4533
rect 3516 4523 3523 4643
rect 3556 4607 3563 4853
rect 3576 4687 3583 4876
rect 3596 4676 3603 4913
rect 3636 4907 3643 4923
rect 3676 4847 3683 5093
rect 3696 4747 3703 5153
rect 3716 5127 3723 5143
rect 3736 4963 3743 5113
rect 3756 5007 3763 5133
rect 3776 4983 3783 5013
rect 3716 4956 3743 4963
rect 3756 4976 3783 4983
rect 3716 4747 3723 4956
rect 3756 4936 3763 4976
rect 3836 4963 3843 5193
rect 3856 5147 3863 5393
rect 3856 4987 3863 5133
rect 3876 5107 3883 5396
rect 3916 5023 3923 5163
rect 3956 5067 3963 5396
rect 3996 5387 4003 5423
rect 3996 5367 4003 5373
rect 4016 5207 4023 5433
rect 4256 5423 4263 5433
rect 4256 5416 4283 5423
rect 4276 5407 4283 5416
rect 4216 5363 4223 5373
rect 4216 5356 4243 5363
rect 4116 5176 4143 5183
rect 3896 5016 3923 5023
rect 3816 4956 3843 4963
rect 3796 4923 3803 4933
rect 3776 4916 3803 4923
rect 3616 4707 3623 4713
rect 3636 4667 3643 4713
rect 3696 4667 3703 4703
rect 3636 4643 3643 4653
rect 3616 4636 3643 4643
rect 3576 4583 3583 4633
rect 3716 4627 3723 4653
rect 3556 4576 3583 4583
rect 3516 4516 3543 4523
rect 3536 4507 3543 4516
rect 3507 4496 3523 4503
rect 3556 4463 3563 4576
rect 3576 4487 3583 4513
rect 3596 4476 3603 4553
rect 3636 4507 3643 4613
rect 3716 4496 3723 4513
rect 3636 4476 3643 4493
rect 3556 4456 3583 4463
rect 3516 4427 3523 4453
rect 3556 4447 3563 4456
rect 3376 3987 3383 4153
rect 3396 4047 3403 4153
rect 3336 3976 3363 3983
rect 3276 3956 3283 3973
rect 3196 3756 3223 3763
rect 3216 3747 3223 3756
rect 3156 3647 3163 3673
rect 2936 3396 2963 3403
rect 2856 3267 2863 3313
rect 2776 3216 2823 3223
rect 2696 2796 2713 2803
rect 2656 2776 2683 2783
rect 2716 2776 2723 2793
rect 2576 2756 2583 2773
rect 2536 2716 2563 2723
rect 2456 2323 2463 2553
rect 2556 2547 2563 2716
rect 2576 2583 2583 2713
rect 2596 2647 2603 2743
rect 2616 2707 2623 2763
rect 2656 2607 2663 2776
rect 2696 2707 2703 2763
rect 2736 2627 2743 2993
rect 2776 2927 2783 2953
rect 2756 2756 2763 2793
rect 2776 2683 2783 2713
rect 2756 2676 2783 2683
rect 2576 2576 2603 2583
rect 2616 2576 2623 2593
rect 2456 2316 2483 2323
rect 2236 2276 2263 2283
rect 2056 1816 2083 1823
rect 2076 1807 2083 1816
rect 2076 1787 2083 1793
rect 2056 1767 2063 1783
rect 2016 1747 2023 1763
rect 2016 1576 2023 1593
rect 1896 1556 1923 1563
rect 1956 1556 1983 1563
rect 1856 1316 1863 1333
rect 1876 1327 1883 1553
rect 1896 1147 1903 1333
rect 1916 1307 1923 1433
rect 1956 1367 1963 1556
rect 1976 1336 1983 1373
rect 1816 1116 1843 1123
rect 1816 967 1823 1116
rect 1856 1107 1863 1113
rect 1596 856 1623 863
rect 1596 827 1603 856
rect 1676 856 1703 863
rect 1736 856 1743 893
rect 1836 887 1843 1083
rect 1916 1083 1923 1273
rect 1996 1187 2003 1513
rect 2016 1336 2023 1373
rect 2036 1367 2043 1563
rect 2056 1547 2063 1733
rect 2076 1627 2083 1773
rect 2096 1603 2103 2013
rect 2156 2007 2163 2063
rect 2176 2027 2183 2093
rect 2216 2087 2223 2253
rect 2256 2227 2263 2276
rect 2136 1796 2143 1993
rect 2156 1827 2163 1993
rect 2176 1887 2183 2013
rect 2076 1596 2103 1603
rect 2076 1567 2083 1596
rect 2096 1347 2103 1533
rect 2116 1527 2123 1713
rect 2036 1307 2043 1323
rect 2076 1316 2103 1323
rect 1896 1076 1923 1083
rect 1936 1116 1963 1123
rect 1996 1116 2003 1133
rect 1676 823 1683 856
rect 1676 816 1703 823
rect 1376 387 1383 613
rect 1396 567 1403 623
rect 1436 567 1443 623
rect 1576 616 1583 693
rect 1696 623 1703 816
rect 1696 616 1723 623
rect 1756 616 1763 813
rect 1776 787 1783 873
rect 1856 867 1863 1053
rect 1896 887 1903 1076
rect 1936 1027 1943 1116
rect 2036 967 2043 1213
rect 2056 907 2063 1313
rect 2076 1147 2083 1293
rect 2096 1287 2103 1316
rect 2116 1127 2123 1453
rect 2136 1427 2143 1533
rect 2156 1407 2163 1783
rect 2176 1707 2183 1803
rect 2196 1667 2203 2073
rect 2236 2056 2243 2133
rect 2216 1667 2223 2043
rect 2256 1796 2263 1893
rect 2276 1847 2283 2313
rect 2356 2276 2363 2293
rect 2376 2263 2383 2293
rect 2456 2267 2463 2283
rect 2376 2256 2403 2263
rect 2316 2207 2323 2233
rect 2316 2007 2323 2043
rect 2356 2027 2363 2043
rect 2376 1887 2383 2256
rect 2436 2207 2443 2263
rect 2396 1907 2403 2133
rect 2416 2056 2423 2093
rect 2436 2076 2443 2173
rect 2456 2107 2463 2193
rect 2476 2187 2483 2316
rect 2496 2247 2503 2433
rect 2516 2227 2523 2533
rect 2536 2447 2543 2543
rect 2556 2296 2563 2433
rect 2576 2407 2583 2576
rect 2596 2556 2603 2576
rect 2536 2207 2543 2263
rect 2476 2076 2483 2093
rect 2456 2047 2463 2063
rect 2456 2027 2463 2033
rect 2496 2027 2503 2093
rect 2316 1787 2323 1833
rect 2276 1776 2293 1783
rect 2336 1743 2343 1833
rect 2356 1816 2363 1833
rect 2336 1736 2353 1743
rect 2316 1687 2323 1713
rect 2236 1447 2243 1573
rect 2156 1336 2183 1343
rect 2176 1327 2183 1336
rect 2136 1147 2143 1273
rect 2176 1143 2183 1313
rect 2156 1136 2183 1143
rect 2076 1067 2083 1113
rect 2136 1067 2143 1083
rect 1796 856 1823 863
rect 1676 607 1683 613
rect 1416 376 1443 383
rect 1436 367 1443 376
rect 1296 207 1303 343
rect 1436 327 1443 353
rect 1456 347 1463 373
rect 1476 367 1483 593
rect 1556 587 1563 603
rect 1716 547 1723 616
rect 1736 587 1743 603
rect 1516 356 1523 433
rect 1556 343 1563 393
rect 1536 336 1563 343
rect 1456 327 1463 333
rect 1396 176 1403 213
rect 1576 136 1583 493
rect 1616 367 1623 383
rect 1596 327 1603 363
rect 1636 347 1643 363
rect 1656 207 1663 333
rect 1676 307 1683 533
rect 1776 447 1783 603
rect 1796 567 1803 856
rect 1876 856 1903 863
rect 1936 856 1943 893
rect 1816 616 1823 733
rect 1876 707 1883 856
rect 1916 827 1923 843
rect 1836 596 1843 673
rect 1676 143 1683 293
rect 1696 147 1703 413
rect 1716 327 1723 433
rect 1776 387 1783 393
rect 1796 376 1803 553
rect 1876 487 1883 603
rect 1896 587 1903 653
rect 1836 376 1863 383
rect 1896 376 1903 513
rect 1916 407 1923 773
rect 1936 636 1943 753
rect 1956 667 1963 873
rect 2076 803 2083 853
rect 2096 827 2103 1053
rect 2136 836 2143 1033
rect 2156 807 2163 1136
rect 2216 1107 2223 1433
rect 2256 1423 2263 1573
rect 2396 1523 2403 1753
rect 2416 1543 2423 2013
rect 2436 1847 2443 1993
rect 2436 1767 2443 1813
rect 2456 1807 2463 1933
rect 2516 1827 2523 2173
rect 2536 2143 2543 2173
rect 2556 2167 2563 2193
rect 2536 2136 2563 2143
rect 2556 2056 2563 2136
rect 2576 2107 2583 2373
rect 2596 2167 2603 2253
rect 2616 2087 2623 2473
rect 2636 2147 2643 2513
rect 2656 2327 2663 2573
rect 2696 2487 2703 2543
rect 2696 2307 2703 2473
rect 2716 2263 2723 2433
rect 2736 2307 2743 2613
rect 2756 2487 2763 2676
rect 2776 2536 2783 2613
rect 2796 2567 2803 3193
rect 2856 3167 2863 3223
rect 2876 3207 2883 3333
rect 2896 3256 2903 3273
rect 2936 3256 2943 3293
rect 2896 3143 2903 3193
rect 2916 3167 2923 3243
rect 2956 3207 2963 3396
rect 3087 3356 3093 3363
rect 2996 3236 3003 3273
rect 3056 3243 3063 3253
rect 3036 3236 3063 3243
rect 2976 3167 2983 3213
rect 2896 3136 2923 3143
rect 2816 2767 2823 3023
rect 2836 2947 2843 3053
rect 2856 3007 2863 3133
rect 2916 2987 2923 3136
rect 2836 2847 2843 2933
rect 2936 2787 2943 3033
rect 2956 3016 2963 3073
rect 3016 3036 3023 3093
rect 3036 3067 3043 3236
rect 3076 3087 3083 3273
rect 3136 3247 3143 3393
rect 3156 3367 3163 3493
rect 3176 3287 3183 3593
rect 3196 3587 3203 3723
rect 3236 3707 3243 3933
rect 3276 3807 3283 3813
rect 3316 3807 3323 3963
rect 3336 3827 3343 3976
rect 3396 3976 3403 4033
rect 3256 3607 3263 3753
rect 3276 3703 3283 3793
rect 3316 3727 3323 3753
rect 3356 3716 3363 3733
rect 3396 3703 3403 3733
rect 3276 3696 3303 3703
rect 3336 3627 3343 3703
rect 3376 3696 3403 3703
rect 3196 3256 3203 3333
rect 3096 3227 3103 3243
rect 3216 3243 3223 3353
rect 3216 3236 3243 3243
rect 3116 3167 3123 3223
rect 3156 3207 3163 3223
rect 3096 3027 3103 3093
rect 2896 2776 2923 2783
rect 2836 2727 2843 2763
rect 2916 2747 2923 2776
rect 2956 2623 2963 2953
rect 2996 2887 3003 3023
rect 3056 2987 3063 3023
rect 3116 2807 3123 3073
rect 3136 2967 3143 3193
rect 3156 2987 3163 3173
rect 3176 3087 3183 3233
rect 3196 3127 3203 3193
rect 2976 2647 2983 2753
rect 3016 2747 3023 2763
rect 2956 2616 2983 2623
rect 2956 2576 2963 2593
rect 2976 2447 2983 2616
rect 3076 2567 3083 2793
rect 3116 2756 3123 2773
rect 3136 2607 3143 2743
rect 3156 2727 3163 2763
rect 3176 2747 3183 2993
rect 3216 2827 3223 3133
rect 3236 3087 3243 3213
rect 3256 3147 3263 3533
rect 3296 3507 3303 3613
rect 3316 3467 3323 3483
rect 3316 3347 3323 3453
rect 3236 3016 3243 3053
rect 3256 2996 3263 3033
rect 3276 3016 3283 3093
rect 3316 3067 3323 3073
rect 3336 3047 3343 3573
rect 3356 3516 3363 3533
rect 3396 3516 3403 3553
rect 3416 3547 3423 3963
rect 3436 3747 3443 4213
rect 3476 4107 3483 4183
rect 3476 4087 3483 4093
rect 3476 3976 3483 4033
rect 3456 3767 3463 3963
rect 3516 3827 3523 4173
rect 3536 3967 3543 4433
rect 3556 4407 3563 4413
rect 3656 4247 3663 4493
rect 3696 4476 3703 4493
rect 3736 4487 3743 4733
rect 3816 4703 3823 4956
rect 3836 4727 3843 4913
rect 3876 4847 3883 4923
rect 3896 4887 3903 5016
rect 3916 4987 3923 4993
rect 3956 4976 3983 4983
rect 4016 4976 4023 5113
rect 4036 4987 4043 5163
rect 4056 5147 4063 5173
rect 4116 5127 4123 5176
rect 4156 5127 4163 5163
rect 3916 4943 3923 4973
rect 3976 4967 3983 4976
rect 3987 4956 4003 4963
rect 4056 4956 4063 4973
rect 3976 4943 3983 4953
rect 3916 4936 3943 4943
rect 3956 4936 3983 4943
rect 3796 4696 3843 4703
rect 3776 4627 3783 4683
rect 3816 4647 3823 4673
rect 3836 4643 3843 4696
rect 3876 4647 3883 4663
rect 3836 4636 3863 4643
rect 3556 4187 3563 4213
rect 3596 4087 3603 4153
rect 3556 3996 3563 4073
rect 3576 4016 3583 4033
rect 3616 4003 3623 4233
rect 3716 4183 3723 4453
rect 3756 4227 3763 4513
rect 3796 4476 3803 4493
rect 3836 4476 3843 4513
rect 3656 4147 3663 4183
rect 3696 4167 3703 4183
rect 3716 4176 3743 4183
rect 3656 4016 3663 4033
rect 3596 3996 3623 4003
rect 3456 3716 3463 3733
rect 3496 3687 3503 3713
rect 3436 3516 3443 3593
rect 3516 3523 3523 3793
rect 3576 3627 3583 3683
rect 3616 3607 3623 3773
rect 3676 3747 3683 3983
rect 3656 3587 3663 3683
rect 3496 3516 3523 3523
rect 3376 3483 3383 3503
rect 3356 3476 3383 3483
rect 3356 3247 3363 3476
rect 3476 3387 3483 3493
rect 3496 3343 3503 3516
rect 3536 3476 3543 3553
rect 3696 3547 3703 4033
rect 3716 4027 3723 4176
rect 3736 4007 3743 4153
rect 3756 4027 3763 4073
rect 3776 4016 3783 4093
rect 3796 4047 3803 4433
rect 3876 4247 3883 4553
rect 3896 4547 3903 4713
rect 3916 4676 3923 4693
rect 3936 4627 3943 4713
rect 3956 4667 3963 4936
rect 4076 4927 4083 4943
rect 4116 4936 4123 4953
rect 4136 4927 4143 4973
rect 4076 4907 4083 4913
rect 3976 4696 3983 4713
rect 4036 4647 4043 4693
rect 4056 4687 4063 4713
rect 3896 4223 3903 4493
rect 3956 4476 3963 4493
rect 3976 4467 3983 4633
rect 3996 4476 4003 4573
rect 4076 4527 4083 4893
rect 4116 4676 4123 4693
rect 4096 4587 4103 4663
rect 4136 4647 4143 4663
rect 4036 4476 4043 4493
rect 3976 4327 3983 4453
rect 4056 4243 4063 4493
rect 4096 4247 4103 4573
rect 4116 4456 4123 4533
rect 4156 4507 4163 4673
rect 4176 4567 4183 5113
rect 4196 4687 4203 5333
rect 4236 5156 4243 5356
rect 4276 5047 4283 5393
rect 4316 5387 4323 5413
rect 4356 5403 4363 5433
rect 4356 5396 4383 5403
rect 4296 5107 4303 5213
rect 4376 5187 4383 5396
rect 4416 5367 4423 5403
rect 4436 5367 4443 5413
rect 4456 5347 4463 5413
rect 4476 5387 4483 5403
rect 4516 5396 4523 5433
rect 4536 5416 4563 5423
rect 4616 5416 4623 5453
rect 5247 5436 5263 5443
rect 4336 5107 4343 5143
rect 4376 5067 4383 5143
rect 4396 5127 4403 5153
rect 4416 5143 4423 5173
rect 4516 5163 4523 5193
rect 4556 5167 4563 5416
rect 4656 5403 4663 5413
rect 4596 5367 4603 5403
rect 4636 5396 4663 5403
rect 4676 5227 4683 5403
rect 4756 5403 4763 5433
rect 5176 5416 5183 5433
rect 4756 5396 4783 5403
rect 4816 5347 4823 5403
rect 4656 5176 4683 5183
rect 4496 5156 4523 5163
rect 4416 5136 4443 5143
rect 4276 4923 4283 5013
rect 4296 4976 4303 5013
rect 4336 4943 4343 4953
rect 4316 4936 4343 4943
rect 4256 4916 4283 4923
rect 4356 4907 4363 5033
rect 4416 4987 4423 5136
rect 4476 5127 4483 5143
rect 4516 5107 4523 5133
rect 4536 5027 4543 5143
rect 4556 5107 4563 5123
rect 4576 5107 4583 5143
rect 4396 4936 4403 4953
rect 4436 4936 4443 4953
rect 4316 4847 4323 4893
rect 4227 4736 4233 4743
rect 4216 4696 4223 4713
rect 4256 4696 4263 4733
rect 4316 4707 4323 4833
rect 4376 4703 4383 4833
rect 4496 4743 4503 4973
rect 4536 4936 4543 4973
rect 4636 4967 4643 5163
rect 4676 5127 4683 5176
rect 4576 4956 4603 4963
rect 4576 4947 4583 4956
rect 4656 4956 4683 4963
rect 4576 4923 4583 4933
rect 4556 4916 4583 4923
rect 4496 4736 4523 4743
rect 4356 4696 4383 4703
rect 4196 4647 4203 4653
rect 4336 4647 4343 4683
rect 4376 4667 4383 4696
rect 4396 4696 4423 4703
rect 4176 4476 4203 4483
rect 4036 4236 4063 4243
rect 3816 4216 3843 4223
rect 3876 4216 3903 4223
rect 3816 4147 3823 4216
rect 3856 4127 3863 4203
rect 3896 4167 3903 4216
rect 3756 3996 3763 4013
rect 3816 3996 3823 4013
rect 3736 3727 3743 3743
rect 3716 3567 3723 3723
rect 3836 3687 3843 3713
rect 3556 3496 3563 3513
rect 3496 3336 3523 3343
rect 3356 3167 3363 3203
rect 3356 3047 3363 3133
rect 3236 2847 3243 2953
rect 3216 2647 3223 2793
rect 3256 2756 3263 2793
rect 3276 2727 3283 2743
rect 3216 2576 3223 2593
rect 3056 2543 3063 2553
rect 3056 2536 3083 2543
rect 2636 2056 2643 2113
rect 2656 2076 2663 2233
rect 2676 2207 2683 2243
rect 2696 2207 2703 2263
rect 2716 2256 2743 2263
rect 2716 2187 2723 2256
rect 2696 2076 2723 2083
rect 2536 2027 2543 2043
rect 2576 1867 2583 2013
rect 2496 1816 2513 1823
rect 2496 1796 2503 1816
rect 2456 1743 2463 1773
rect 2476 1763 2483 1773
rect 2476 1756 2503 1763
rect 2436 1736 2463 1743
rect 2436 1607 2443 1736
rect 2456 1547 2463 1693
rect 2416 1536 2443 1543
rect 2396 1516 2423 1523
rect 2236 1416 2263 1423
rect 2236 1167 2243 1416
rect 2276 1307 2283 1343
rect 2316 1336 2323 1353
rect 2276 1147 2283 1293
rect 2296 1287 2303 1323
rect 2176 1067 2183 1073
rect 2196 1067 2203 1103
rect 2236 1087 2243 1133
rect 2316 1116 2323 1253
rect 2336 1127 2343 1493
rect 2356 1316 2363 1373
rect 2396 1316 2403 1433
rect 2416 1427 2423 1516
rect 2436 1347 2443 1536
rect 2476 1523 2483 1733
rect 2456 1516 2483 1523
rect 2076 796 2123 803
rect 1976 636 1983 753
rect 1776 323 1783 373
rect 1856 347 1863 376
rect 1916 347 1923 363
rect 1756 316 1783 323
rect 1716 156 1723 313
rect 1756 156 1763 213
rect 1656 136 1683 143
rect 1836 123 1843 273
rect 1916 267 1923 313
rect 1936 267 1943 383
rect 1976 363 1983 393
rect 1996 367 2003 573
rect 2016 383 2023 693
rect 2036 467 2043 673
rect 2096 636 2103 796
rect 2076 603 2083 623
rect 2116 616 2123 653
rect 2056 596 2083 603
rect 2016 376 2043 383
rect 1956 356 1983 363
rect 1976 347 1983 356
rect 1996 267 2003 323
rect 1916 147 1923 253
rect 1936 207 1943 253
rect 1996 227 2003 253
rect 1956 156 1963 173
rect 1996 167 2003 193
rect 1236 67 1243 123
rect 1836 116 1863 123
rect 1896 87 1903 123
rect 2016 107 2023 173
rect 2036 156 2043 376
rect 2056 367 2063 596
rect 2076 387 2083 533
rect 2136 407 2143 713
rect 2176 687 2183 1033
rect 2196 827 2203 893
rect 2216 887 2223 1073
rect 2256 1047 2263 1103
rect 2296 1067 2303 1103
rect 2336 1027 2343 1093
rect 2316 887 2323 913
rect 2216 803 2223 853
rect 2276 836 2283 853
rect 2336 836 2343 873
rect 2356 867 2363 1273
rect 2376 1267 2383 1283
rect 2436 1267 2443 1313
rect 2456 1287 2463 1516
rect 2496 1507 2503 1756
rect 2516 1707 2523 1793
rect 2536 1783 2543 1853
rect 2596 1807 2603 1973
rect 2616 1803 2623 1873
rect 2636 1827 2643 2013
rect 2676 2007 2683 2063
rect 2716 1947 2723 2076
rect 2616 1796 2643 1803
rect 2676 1796 2683 1813
rect 2636 1783 2643 1796
rect 2536 1776 2563 1783
rect 2636 1776 2653 1783
rect 2696 1776 2723 1783
rect 2547 1756 2563 1763
rect 2536 1583 2543 1733
rect 2556 1647 2563 1756
rect 2587 1756 2603 1763
rect 2516 1576 2543 1583
rect 2516 1483 2523 1553
rect 2496 1476 2523 1483
rect 2476 1287 2483 1353
rect 2496 1307 2503 1476
rect 2536 1367 2543 1493
rect 2556 1447 2563 1593
rect 2576 1387 2583 1573
rect 2596 1563 2603 1756
rect 2636 1727 2643 1753
rect 2616 1596 2623 1713
rect 2656 1627 2663 1753
rect 2696 1596 2703 1753
rect 2716 1707 2723 1776
rect 2736 1747 2743 2213
rect 2756 2107 2763 2133
rect 2796 2127 2803 2293
rect 2816 2227 2823 2273
rect 2836 2207 2843 2263
rect 2856 2167 2863 2243
rect 2876 2167 2883 2253
rect 2896 2187 2903 2373
rect 2916 2267 2923 2393
rect 2796 2076 2803 2093
rect 2856 2067 2863 2113
rect 2896 2103 2903 2173
rect 2936 2127 2943 2433
rect 2976 2367 2983 2393
rect 3016 2307 3023 2313
rect 3056 2287 3063 2493
rect 3096 2447 3103 2513
rect 3116 2407 3123 2523
rect 2956 2247 2963 2263
rect 2996 2247 3003 2263
rect 2876 2096 2903 2103
rect 2876 2076 2883 2096
rect 2916 2076 2923 2093
rect 2956 2087 2963 2233
rect 2976 2167 2983 2243
rect 2776 1967 2783 2033
rect 2816 2027 2823 2063
rect 2896 2047 2903 2063
rect 2756 1747 2763 1953
rect 2776 1827 2783 1893
rect 2796 1847 2803 1993
rect 2816 1987 2823 2013
rect 2796 1823 2803 1833
rect 2836 1827 2843 1853
rect 2856 1847 2863 2033
rect 2936 1987 2943 2063
rect 2976 2043 2983 2113
rect 2956 2036 2983 2043
rect 2956 1963 2963 2036
rect 2936 1956 2963 1963
rect 2936 1847 2943 1956
rect 2976 1847 2983 1993
rect 2996 1907 3003 2093
rect 3016 1887 3023 2273
rect 3036 2107 3043 2253
rect 3056 2207 3063 2243
rect 3076 2187 3083 2263
rect 3047 2096 3063 2103
rect 2887 1836 2923 1843
rect 2796 1816 2823 1823
rect 2816 1796 2823 1816
rect 2916 1816 2923 1836
rect 2736 1667 2743 1733
rect 2776 1687 2783 1793
rect 2856 1787 2863 1803
rect 2836 1727 2843 1783
rect 2876 1727 2883 1813
rect 2596 1556 2623 1563
rect 2616 1547 2623 1556
rect 2596 1447 2603 1533
rect 2376 1047 2383 1173
rect 2476 1123 2483 1253
rect 2516 1247 2523 1303
rect 2556 1287 2563 1303
rect 2616 1247 2623 1373
rect 2476 1116 2503 1123
rect 2536 1116 2543 1133
rect 2576 1116 2603 1123
rect 2456 1096 2463 1113
rect 2476 1083 2483 1116
rect 2476 1076 2503 1083
rect 2396 887 2403 893
rect 2196 796 2223 803
rect 2196 656 2203 796
rect 2216 787 2223 796
rect 2236 783 2243 813
rect 2256 807 2263 823
rect 2236 776 2263 783
rect 2167 636 2183 643
rect 2216 636 2223 673
rect 2236 636 2243 713
rect 2256 647 2263 776
rect 2296 747 2303 823
rect 2296 636 2303 733
rect 2156 547 2163 633
rect 2076 343 2083 373
rect 2176 347 2183 533
rect 2076 336 2103 343
rect 2196 343 2203 393
rect 2196 336 2223 343
rect 2056 267 2063 333
rect 2236 316 2253 323
rect 2096 136 2103 173
rect 2116 87 2123 153
rect 2136 107 2143 153
rect 2156 147 2163 233
rect 2196 156 2203 173
rect 2236 156 2243 293
rect 2176 136 2183 153
rect 2256 47 2263 253
rect 2276 187 2283 593
rect 2296 287 2303 593
rect 2316 387 2323 813
rect 2376 707 2383 813
rect 2396 707 2403 853
rect 2416 767 2423 1053
rect 2436 867 2443 1013
rect 2436 787 2443 833
rect 2336 607 2343 623
rect 2376 467 2383 613
rect 2376 347 2383 393
rect 2316 327 2323 343
rect 2356 327 2363 343
rect 2336 267 2343 323
rect 2276 123 2283 133
rect 2356 123 2363 173
rect 2396 156 2403 553
rect 2416 387 2423 653
rect 2436 467 2443 693
rect 2456 507 2463 1053
rect 2496 867 2503 1076
rect 2516 967 2523 1103
rect 2556 1027 2563 1103
rect 2596 1087 2603 1116
rect 2536 927 2543 953
rect 2556 887 2563 1013
rect 2616 887 2623 1093
rect 2636 1067 2643 1513
rect 2656 1327 2663 1553
rect 2676 1547 2683 1583
rect 2716 1563 2723 1633
rect 2756 1576 2763 1673
rect 2716 1556 2743 1563
rect 2716 1467 2723 1556
rect 2656 1287 2663 1313
rect 2676 1263 2683 1303
rect 2676 1256 2703 1263
rect 2696 1227 2703 1256
rect 2716 1247 2723 1303
rect 2736 1267 2743 1513
rect 2756 1347 2763 1533
rect 2776 1527 2783 1563
rect 2796 1467 2803 1613
rect 2816 1387 2823 1613
rect 2836 1576 2843 1593
rect 2856 1556 2863 1653
rect 2896 1647 2903 1813
rect 2876 1576 2883 1613
rect 2896 1547 2903 1563
rect 2836 1367 2843 1433
rect 2856 1387 2863 1513
rect 2876 1447 2883 1493
rect 2756 1316 2763 1333
rect 2776 1307 2783 1353
rect 2796 1247 2803 1303
rect 2816 1227 2823 1283
rect 2836 1267 2843 1303
rect 2836 1223 2843 1253
rect 2856 1247 2863 1283
rect 2836 1216 2863 1223
rect 2676 1096 2683 1173
rect 2696 1147 2703 1213
rect 2716 1107 2723 1133
rect 2656 1027 2663 1083
rect 2696 1063 2703 1073
rect 2676 1056 2703 1063
rect 2636 863 2643 913
rect 2616 856 2643 863
rect 2476 827 2483 843
rect 2556 827 2563 843
rect 2476 607 2483 813
rect 2496 807 2503 813
rect 2516 616 2523 793
rect 2536 747 2543 823
rect 2596 807 2603 843
rect 2556 627 2563 653
rect 2576 636 2603 643
rect 2636 636 2643 833
rect 2656 823 2663 873
rect 2676 867 2683 1056
rect 2716 1027 2723 1073
rect 2736 1067 2743 1153
rect 2756 1087 2763 1113
rect 2776 1096 2783 1173
rect 2796 1116 2803 1173
rect 2836 1147 2843 1153
rect 2756 927 2763 1073
rect 2816 947 2823 1103
rect 2856 1083 2863 1216
rect 2836 1076 2863 1083
rect 2876 1083 2883 1303
rect 2896 1187 2903 1513
rect 2916 1327 2923 1713
rect 2936 1687 2943 1793
rect 2956 1763 2963 1823
rect 2976 1787 2983 1803
rect 2956 1756 2983 1763
rect 2976 1707 2983 1756
rect 2996 1687 3003 1873
rect 3036 1863 3043 2053
rect 3056 1947 3063 2053
rect 3076 1867 3083 2093
rect 3036 1856 3063 1863
rect 3056 1843 3063 1856
rect 3056 1836 3083 1843
rect 3036 1816 3043 1833
rect 3076 1816 3083 1836
rect 3016 1787 3023 1813
rect 3056 1787 3063 1803
rect 3096 1787 3103 2173
rect 3116 2107 3123 2213
rect 3136 2107 3143 2553
rect 3176 2527 3183 2573
rect 3236 2556 3243 2693
rect 3296 2687 3303 2763
rect 3176 2276 3183 2473
rect 3156 2167 3163 2263
rect 3176 2147 3183 2193
rect 3116 1903 3123 2033
rect 3136 1927 3143 2063
rect 3176 2056 3203 2063
rect 3196 2027 3203 2056
rect 3216 2003 3223 2513
rect 3256 2487 3263 2673
rect 3276 2556 3283 2633
rect 3296 2523 3303 2593
rect 3316 2567 3323 3033
rect 3356 3016 3383 3023
rect 3336 2987 3343 3013
rect 3356 3007 3363 3016
rect 3396 2996 3403 3013
rect 3356 2967 3363 2973
rect 3336 2767 3343 2813
rect 3376 2723 3383 2973
rect 3416 2723 3423 2953
rect 3456 2783 3463 3053
rect 3476 3007 3483 3113
rect 3496 3047 3503 3293
rect 3516 3067 3523 3336
rect 3576 3303 3583 3483
rect 3556 3296 3583 3303
rect 3536 3227 3543 3243
rect 3556 3047 3563 3296
rect 3576 3247 3583 3273
rect 3596 3227 3603 3413
rect 3616 3287 3623 3533
rect 3636 3516 3663 3523
rect 3636 3487 3643 3516
rect 3736 3516 3743 3593
rect 3756 3507 3763 3533
rect 3776 3507 3783 3673
rect 3676 3467 3683 3503
rect 3616 3236 3623 3253
rect 3496 2807 3503 3033
rect 3516 3016 3523 3033
rect 3536 3023 3543 3033
rect 3536 3016 3563 3023
rect 3516 2787 3523 2973
rect 3336 2707 3343 2723
rect 3356 2716 3383 2723
rect 3396 2716 3423 2723
rect 3436 2776 3463 2783
rect 3296 2516 3323 2523
rect 3256 2276 3263 2353
rect 3296 2276 3303 2293
rect 3236 2247 3243 2263
rect 3256 2056 3263 2233
rect 3276 2007 3283 2043
rect 3196 1996 3223 2003
rect 3156 1927 3163 1973
rect 3116 1896 3143 1903
rect 3136 1847 3143 1896
rect 3116 1816 3123 1833
rect 3107 1756 3113 1763
rect 2967 1616 3003 1623
rect 2936 1507 2943 1613
rect 3036 1596 3043 1653
rect 2956 1503 2963 1593
rect 3056 1587 3063 1753
rect 3076 1596 3083 1713
rect 3136 1627 3143 1713
rect 3116 1596 3123 1613
rect 3156 1596 3163 1773
rect 2976 1527 2983 1583
rect 2956 1496 2983 1503
rect 2936 1447 2943 1473
rect 2956 1316 2963 1453
rect 2976 1447 2983 1496
rect 2976 1307 2983 1333
rect 2936 1247 2943 1283
rect 2936 1167 2943 1233
rect 2896 1116 2903 1133
rect 2976 1116 2983 1273
rect 2916 1087 2923 1103
rect 2956 1087 2963 1103
rect 2876 1076 2903 1083
rect 2836 947 2843 1076
rect 2867 1056 2873 1063
rect 2696 823 2703 843
rect 2656 816 2703 823
rect 2676 727 2683 816
rect 2676 636 2683 693
rect 2496 547 2503 603
rect 2536 527 2543 603
rect 2576 547 2583 636
rect 2696 627 2703 773
rect 2716 767 2723 863
rect 2736 787 2743 843
rect 2716 636 2723 733
rect 2756 667 2763 873
rect 2836 807 2843 823
rect 2596 507 2603 533
rect 2616 527 2623 623
rect 2776 616 2783 773
rect 2796 747 2803 793
rect 2816 747 2823 803
rect 2796 527 2803 673
rect 2416 267 2423 353
rect 2416 247 2423 253
rect 2436 167 2443 433
rect 2536 327 2543 373
rect 2636 347 2643 493
rect 2756 367 2763 453
rect 2816 387 2823 653
rect 2836 387 2843 633
rect 2856 627 2863 853
rect 2876 807 2883 1033
rect 2896 767 2903 1076
rect 2876 596 2883 753
rect 2916 747 2923 1013
rect 2936 967 2943 1033
rect 2956 847 2963 1013
rect 2996 943 3003 1553
rect 3016 1507 3023 1583
rect 3016 1287 3023 1433
rect 3056 1327 3063 1473
rect 3136 1467 3143 1583
rect 3156 1316 3163 1413
rect 3176 1327 3183 1933
rect 3196 1607 3203 1996
rect 3236 1847 3243 1893
rect 3276 1847 3283 1873
rect 3296 1827 3303 2153
rect 3316 2147 3323 2263
rect 3336 2083 3343 2313
rect 3356 2247 3363 2716
rect 3376 2276 3383 2353
rect 3396 2287 3403 2716
rect 3416 2556 3423 2693
rect 3316 2076 3343 2083
rect 3316 1947 3323 2076
rect 3356 2056 3363 2093
rect 3396 2087 3403 2243
rect 3336 1887 3343 2043
rect 3256 1816 3283 1823
rect 3196 1347 3203 1573
rect 3216 1527 3223 1773
rect 3236 1767 3243 1803
rect 3276 1783 3283 1816
rect 3316 1796 3323 1833
rect 3356 1796 3363 1813
rect 3256 1776 3283 1783
rect 3256 1727 3263 1776
rect 3296 1763 3303 1783
rect 3336 1767 3343 1783
rect 3396 1767 3403 2013
rect 3416 2003 3423 2153
rect 3436 2127 3443 2776
rect 3556 2756 3563 2973
rect 3576 2767 3583 3003
rect 3596 2756 3603 2773
rect 3456 2743 3463 2753
rect 3536 2743 3543 2753
rect 3456 2736 3483 2743
rect 3516 2736 3543 2743
rect 3536 2727 3543 2736
rect 3496 2687 3503 2723
rect 3576 2667 3583 2723
rect 3456 2556 3463 2593
rect 3616 2567 3623 2743
rect 3476 2367 3483 2553
rect 3496 2287 3503 2553
rect 3636 2543 3643 3453
rect 3696 3287 3703 3473
rect 3756 3283 3763 3493
rect 3756 3276 3783 3283
rect 3716 3256 3743 3263
rect 3696 3223 3703 3243
rect 3696 3216 3723 3223
rect 3676 2907 3683 3023
rect 3716 2767 3723 3216
rect 3736 3067 3743 3256
rect 3776 3236 3783 3276
rect 3756 3023 3763 3053
rect 3736 3016 3763 3023
rect 3676 2756 3703 2763
rect 3696 2723 3703 2756
rect 3736 2756 3743 2773
rect 3696 2716 3723 2723
rect 3636 2536 3663 2543
rect 3516 2387 3523 2513
rect 3456 2256 3483 2263
rect 3456 2147 3463 2256
rect 3476 2236 3503 2243
rect 3476 2107 3483 2236
rect 3516 2223 3523 2263
rect 3556 2247 3563 2413
rect 3596 2263 3603 2353
rect 3616 2307 3623 2533
rect 3496 2216 3523 2223
rect 3496 2207 3503 2216
rect 3496 2087 3503 2193
rect 3416 1996 3443 2003
rect 3416 1787 3423 1973
rect 3436 1847 3443 1996
rect 3476 1967 3483 2053
rect 3296 1756 3323 1763
rect 3256 1576 3263 1613
rect 3236 1427 3243 1563
rect 3276 1556 3283 1753
rect 3296 1627 3303 1693
rect 3296 1576 3303 1593
rect 3016 1147 3023 1253
rect 3036 1147 3043 1293
rect 3056 1116 3063 1153
rect 3076 1096 3083 1303
rect 2996 936 3023 943
rect 2976 827 2983 933
rect 2936 727 2943 813
rect 2996 723 3003 913
rect 3016 827 3023 936
rect 3056 867 3063 933
rect 2976 716 3003 723
rect 2896 627 2903 713
rect 2936 647 2943 713
rect 2936 587 2943 613
rect 2956 607 2963 693
rect 2876 376 2883 453
rect 2896 407 2903 493
rect 2936 367 2943 433
rect 2956 407 2963 513
rect 2976 467 2983 716
rect 3036 667 3043 843
rect 3076 836 3083 953
rect 3096 927 3103 1273
rect 3116 1096 3123 1273
rect 3136 1247 3143 1313
rect 3236 1307 3243 1333
rect 3216 1287 3223 1303
rect 3156 1163 3163 1233
rect 3176 1187 3183 1283
rect 3156 1156 3183 1163
rect 3136 1107 3143 1153
rect 3156 1096 3163 1133
rect 3176 1127 3183 1156
rect 3176 967 3183 1083
rect 3196 967 3203 1153
rect 3216 1027 3223 1253
rect 3256 1247 3263 1513
rect 3296 1316 3303 1433
rect 3316 1347 3323 1756
rect 3376 1727 3383 1753
rect 3336 1387 3343 1713
rect 3396 1687 3403 1733
rect 3416 1647 3423 1773
rect 3436 1707 3443 1813
rect 3476 1796 3483 1953
rect 3536 1827 3543 2233
rect 3576 2167 3583 2263
rect 3596 2256 3623 2263
rect 3636 2127 3643 2473
rect 3656 2367 3663 2536
rect 3556 2076 3563 2093
rect 3576 2067 3583 2093
rect 3616 2076 3623 2113
rect 3656 2103 3663 2263
rect 3636 2096 3663 2103
rect 3467 1756 3473 1763
rect 3496 1743 3503 1783
rect 3496 1736 3523 1743
rect 3436 1623 3443 1673
rect 3427 1616 3443 1623
rect 3476 1607 3483 1713
rect 3356 1567 3363 1583
rect 3356 1527 3363 1553
rect 3376 1447 3383 1553
rect 3396 1467 3403 1593
rect 3436 1576 3443 1593
rect 3416 1547 3423 1563
rect 3196 887 3203 933
rect 3056 707 3063 823
rect 3036 636 3043 653
rect 3056 616 3063 633
rect 3096 627 3103 793
rect 3116 767 3123 833
rect 3216 827 3223 913
rect 3236 887 3243 1213
rect 3276 1127 3283 1273
rect 3316 1247 3323 1303
rect 3336 1287 3343 1323
rect 3356 1167 3363 1373
rect 3376 1307 3383 1413
rect 3407 1376 3413 1383
rect 3456 1336 3463 1373
rect 3476 1367 3483 1573
rect 3496 1447 3503 1713
rect 3516 1707 3523 1736
rect 3536 1687 3543 1753
rect 3556 1687 3563 1933
rect 3576 1707 3583 1993
rect 3616 1807 3623 1833
rect 3596 1756 3623 1763
rect 3596 1647 3603 1756
rect 3616 1707 3623 1733
rect 3616 1687 3623 1693
rect 3616 1623 3623 1633
rect 3576 1616 3623 1623
rect 3576 1596 3583 1616
rect 3516 1567 3523 1583
rect 3536 1547 3543 1573
rect 3376 1187 3383 1273
rect 3396 1227 3403 1313
rect 3416 1307 3423 1333
rect 3436 1307 3443 1323
rect 3376 1167 3383 1173
rect 3316 1116 3323 1133
rect 3276 1076 3303 1083
rect 3256 1047 3263 1073
rect 3276 1007 3283 1076
rect 3136 807 3143 823
rect 3176 807 3183 823
rect 3116 636 3123 753
rect 3156 636 3163 793
rect 3176 616 3183 633
rect 2716 347 2723 363
rect 2647 336 2663 343
rect 2476 187 2483 213
rect 2516 176 2523 193
rect 2476 143 2483 173
rect 2556 156 2563 213
rect 2576 143 2583 293
rect 2616 267 2623 323
rect 2476 136 2503 143
rect 2276 116 2303 123
rect 2336 116 2363 123
rect 2536 107 2543 143
rect 2576 136 2603 143
rect 2636 107 2643 213
rect 2656 147 2663 253
rect 2696 243 2703 343
rect 2736 267 2743 353
rect 2696 236 2743 243
rect 2676 156 2683 193
rect 2716 156 2723 213
rect 2736 167 2743 236
rect 2756 67 2763 353
rect 2776 243 2783 333
rect 2796 267 2803 333
rect 2816 243 2823 343
rect 2776 236 2823 243
rect 2796 123 2803 193
rect 2876 123 2883 193
rect 2936 176 2943 193
rect 2916 156 2923 173
rect 2956 156 2963 393
rect 3016 383 3023 593
rect 3076 487 3083 613
rect 2996 376 3023 383
rect 2976 267 2983 373
rect 2996 347 3003 376
rect 3056 367 3063 383
rect 3096 367 3103 553
rect 3136 507 3143 613
rect 3196 587 3203 813
rect 3216 627 3223 753
rect 3236 747 3243 853
rect 3256 767 3263 843
rect 3296 836 3303 1033
rect 3336 927 3343 1113
rect 3356 1007 3363 1133
rect 3416 1116 3423 1273
rect 3436 1127 3443 1273
rect 3476 1267 3483 1333
rect 3396 1047 3403 1103
rect 3436 1047 3443 1053
rect 3356 863 3363 953
rect 3396 867 3403 913
rect 3336 856 3363 863
rect 3236 667 3243 713
rect 3276 687 3283 823
rect 3336 787 3343 856
rect 3416 847 3423 933
rect 3236 636 3243 653
rect 3316 607 3323 753
rect 3216 467 3223 593
rect 2996 147 3003 313
rect 3036 187 3043 363
rect 3096 156 3103 233
rect 3116 167 3123 413
rect 3136 387 3143 453
rect 3136 247 3143 353
rect 2796 116 2823 123
rect 2856 116 2883 123
rect 3076 87 3083 143
rect 3156 136 3163 363
rect 3196 356 3203 413
rect 3216 327 3223 343
rect 3236 307 3243 593
rect 3276 356 3283 393
rect 3236 176 3243 193
rect 3116 123 3123 133
rect 3196 123 3203 153
rect 3116 116 3143 123
rect 3176 116 3203 123
rect 3216 87 3223 153
rect 3276 67 3283 293
rect 3296 247 3303 333
rect 3336 307 3343 613
rect 3356 607 3363 733
rect 3376 636 3383 813
rect 3396 667 3403 753
rect 3416 656 3423 733
rect 3436 667 3443 993
rect 3456 967 3463 1233
rect 3476 1047 3483 1173
rect 3496 1127 3503 1373
rect 3516 1227 3523 1533
rect 3536 1347 3543 1433
rect 3556 1247 3563 1553
rect 3616 1547 3623 1593
rect 3576 1367 3583 1513
rect 3576 1316 3583 1353
rect 3596 1347 3603 1433
rect 3596 1247 3603 1303
rect 3516 1096 3523 1173
rect 3496 927 3503 1073
rect 3496 856 3523 863
rect 3367 476 3373 483
rect 3396 447 3403 613
rect 3436 607 3443 623
rect 3456 427 3463 813
rect 3516 747 3523 856
rect 3356 327 3363 353
rect 3296 127 3303 173
rect 3316 156 3323 253
rect 3376 167 3383 373
rect 3416 367 3423 373
rect 3456 356 3463 413
rect 3396 307 3403 343
rect 3436 176 3443 193
rect 3456 156 3463 253
rect 3376 136 3383 153
rect 3476 27 3483 653
rect 3536 643 3543 1073
rect 3556 807 3563 1213
rect 3576 1087 3583 1113
rect 3596 1027 3603 1213
rect 3616 1187 3623 1473
rect 3636 1347 3643 2096
rect 3656 1927 3663 2063
rect 3676 1867 3683 2633
rect 3696 2487 3703 2593
rect 3716 2527 3723 2693
rect 3756 2627 3763 2893
rect 3756 2543 3763 2613
rect 3736 2536 3763 2543
rect 3776 2487 3783 3173
rect 3796 2667 3803 3613
rect 3816 3067 3823 3393
rect 3856 3283 3863 3813
rect 3916 3707 3923 4233
rect 3956 4167 3963 4183
rect 3936 4147 3943 4163
rect 3976 4143 3983 4193
rect 4036 4187 4043 4236
rect 3956 4136 3983 4143
rect 3956 3987 3963 4136
rect 4036 4047 4043 4173
rect 4056 4027 4063 4203
rect 4076 4107 4083 4223
rect 4116 4216 4123 4413
rect 4156 4267 4163 4463
rect 4196 4443 4203 4476
rect 4176 4436 4203 4443
rect 4096 4167 4103 4203
rect 4016 3947 4023 3993
rect 4036 3963 4043 4013
rect 4036 3956 4063 3963
rect 3936 3716 3963 3723
rect 3876 3467 3883 3633
rect 3896 3607 3903 3683
rect 3936 3567 3943 3716
rect 4036 3707 4043 3956
rect 4116 3927 4123 4173
rect 4156 4107 4163 4253
rect 4136 3967 4143 4093
rect 4176 4067 4183 4436
rect 4216 4427 4223 4633
rect 4256 4476 4263 4493
rect 4236 4456 4243 4473
rect 4316 4463 4323 4533
rect 4316 4456 4343 4463
rect 4356 4447 4363 4473
rect 4396 4467 4403 4696
rect 4496 4687 4503 4713
rect 4516 4707 4523 4736
rect 4576 4696 4583 4713
rect 4436 4667 4443 4683
rect 4476 4676 4493 4683
rect 4236 4167 4243 4223
rect 4256 4187 4263 4203
rect 4236 4127 4243 4153
rect 4256 4147 4263 4173
rect 4016 3607 4023 3703
rect 3936 3496 3943 3553
rect 4016 3536 4033 3543
rect 4056 3543 4063 3833
rect 4116 3767 4123 3913
rect 4136 3716 4143 3773
rect 4096 3647 4103 3673
rect 4056 3536 4083 3543
rect 3916 3407 3923 3483
rect 3956 3467 3963 3483
rect 3976 3407 3983 3533
rect 3856 3276 3883 3283
rect 3836 3236 3863 3243
rect 3836 3227 3843 3236
rect 3836 3023 3843 3213
rect 3876 3127 3883 3276
rect 4056 3203 4063 3513
rect 4076 3487 4083 3536
rect 4096 3516 4103 3633
rect 4116 3587 4123 3713
rect 4116 3536 4123 3573
rect 4136 3516 4143 3533
rect 4136 3243 4143 3473
rect 4156 3447 4163 4013
rect 4196 3976 4203 3993
rect 4216 3947 4223 3963
rect 4236 3847 4243 4093
rect 4276 4027 4283 4433
rect 4436 4223 4443 4613
rect 4556 4567 4563 4683
rect 4596 4647 4603 4893
rect 4627 4796 4633 4803
rect 4676 4707 4683 4956
rect 4696 4947 4703 5313
rect 4716 5067 4723 5213
rect 4736 5167 4743 5173
rect 4756 5107 4763 5123
rect 4716 4976 4743 4983
rect 4716 4907 4723 4976
rect 4776 4943 4783 4973
rect 4756 4936 4783 4943
rect 4676 4676 4683 4693
rect 4656 4627 4663 4663
rect 4416 4216 4463 4223
rect 4296 4127 4303 4213
rect 4396 4167 4403 4193
rect 4296 4007 4303 4073
rect 4296 3976 4303 3993
rect 4276 3956 4283 3973
rect 4316 3947 4323 3963
rect 4336 3887 4343 4053
rect 4356 3987 4363 3993
rect 4176 3627 4183 3693
rect 4216 3667 4223 3723
rect 4276 3716 4283 3833
rect 4336 3723 4343 3853
rect 4316 3716 4343 3723
rect 4236 3647 4243 3693
rect 4336 3647 4343 3716
rect 4356 3667 4363 3973
rect 4376 3727 4383 3873
rect 4396 3787 4403 3953
rect 4416 3743 4423 4216
rect 4456 4196 4463 4216
rect 4516 4207 4523 4373
rect 4616 4287 4623 4553
rect 4716 4456 4723 4793
rect 4496 4187 4503 4203
rect 4616 4196 4623 4253
rect 4436 4127 4443 4183
rect 4476 4167 4483 4183
rect 4456 3947 4463 4153
rect 4476 3996 4503 4003
rect 4536 3996 4543 4093
rect 4636 4067 4643 4183
rect 4636 4047 4643 4053
rect 4476 3907 4483 3996
rect 4516 3947 4523 3983
rect 4416 3736 4433 3743
rect 4396 3707 4403 3723
rect 4436 3716 4443 3733
rect 4176 3536 4183 3553
rect 4276 3516 4283 3573
rect 4316 3516 4323 3633
rect 4336 3507 4343 3593
rect 4376 3516 4383 3633
rect 4396 3536 4403 3613
rect 4416 3547 4423 3703
rect 4416 3516 4443 3523
rect 4436 3487 4443 3516
rect 4136 3236 4163 3243
rect 4036 3196 4063 3203
rect 3996 3056 4003 3073
rect 4116 3027 4123 3153
rect 3816 3016 3843 3023
rect 3836 2907 3843 3016
rect 3916 2756 3923 2893
rect 4087 2876 4093 2883
rect 3816 2687 3823 2743
rect 3856 2647 3863 2743
rect 3916 2576 3943 2583
rect 3696 2167 3703 2453
rect 3716 2247 3723 2453
rect 3936 2447 3943 2576
rect 4036 2536 4043 2873
rect 4116 2827 4123 2973
rect 4136 2803 4143 3213
rect 4156 2887 4163 3003
rect 4116 2796 4143 2803
rect 4056 2756 4063 2773
rect 3736 2327 3743 2373
rect 3736 2267 3743 2313
rect 3796 2296 3803 2313
rect 3696 1827 3703 2153
rect 3716 1827 3723 2173
rect 3776 2147 3783 2283
rect 3816 2167 3823 2313
rect 3836 2263 3843 2293
rect 3856 2283 3863 2353
rect 3856 2276 3883 2283
rect 3836 2256 3863 2263
rect 3736 2007 3743 2113
rect 3776 2107 3783 2133
rect 3756 2047 3763 2063
rect 3656 1727 3663 1813
rect 3736 1796 3743 1893
rect 3776 1787 3783 2053
rect 3836 1907 3843 2213
rect 3856 1887 3863 2256
rect 3876 1947 3883 2233
rect 3916 2056 3923 2213
rect 3936 2187 3943 2253
rect 3956 2247 3963 2273
rect 3976 2227 3983 2433
rect 4016 2287 4023 2333
rect 3936 2027 3943 2043
rect 3796 1796 3803 1833
rect 3836 1796 3843 1873
rect 3876 1827 3883 1853
rect 3676 1767 3683 1783
rect 3656 1607 3663 1693
rect 3676 1576 3683 1733
rect 3696 1683 3703 1753
rect 3716 1747 3723 1783
rect 3736 1727 3743 1753
rect 3696 1676 3723 1683
rect 3656 1407 3663 1563
rect 3716 1547 3723 1676
rect 3736 1567 3743 1673
rect 3756 1647 3763 1753
rect 3776 1667 3783 1753
rect 3816 1747 3823 1763
rect 3776 1576 3783 1633
rect 3796 1627 3803 1653
rect 3816 1603 3823 1693
rect 3836 1667 3843 1713
rect 3876 1663 3883 1793
rect 3896 1787 3903 2013
rect 3956 1827 3963 2173
rect 3976 2107 3983 2133
rect 3976 1867 3983 2073
rect 3996 2027 4003 2153
rect 4036 2083 4043 2353
rect 4056 2307 4063 2653
rect 4076 2587 4083 2793
rect 4096 2187 4103 2773
rect 4116 2763 4123 2796
rect 4176 2787 4183 3333
rect 4236 3167 4243 3253
rect 4256 3023 4263 3053
rect 4236 3016 4263 3023
rect 4116 2756 4143 2763
rect 4147 2736 4163 2743
rect 4116 2187 4123 2733
rect 4136 2576 4143 2653
rect 4196 2647 4203 2743
rect 4216 2687 4223 3013
rect 4236 2787 4243 2793
rect 4236 2756 4243 2773
rect 4176 2543 4183 2573
rect 4156 2536 4183 2543
rect 4196 2407 4203 2593
rect 4236 2556 4243 2713
rect 4256 2627 4263 2913
rect 4276 2607 4283 3433
rect 4356 3243 4363 3473
rect 4336 3236 4363 3243
rect 4336 3203 4343 3236
rect 4456 3223 4463 3613
rect 4496 3527 4503 3933
rect 4536 3703 4543 3773
rect 4536 3696 4563 3703
rect 4596 3687 4603 3913
rect 4576 3667 4583 3683
rect 4556 3503 4563 3633
rect 4556 3496 4583 3503
rect 4556 3483 4563 3496
rect 4536 3476 4563 3483
rect 4596 3367 4603 3513
rect 4616 3287 4623 4033
rect 4656 3987 4663 4273
rect 4676 4207 4683 4233
rect 4696 4103 4703 4293
rect 4676 4096 4703 4103
rect 4636 3927 4643 3983
rect 4676 3727 4683 4096
rect 4696 3927 4703 4073
rect 4716 3976 4723 4053
rect 4636 3716 4663 3723
rect 4636 3503 4643 3716
rect 4636 3496 4653 3503
rect 4636 3247 4643 3496
rect 4676 3347 4683 3713
rect 4736 3627 4743 4933
rect 4776 4203 4783 4453
rect 4796 4307 4803 5273
rect 4876 5207 4883 5413
rect 4916 5387 4923 5403
rect 4887 5196 4903 5203
rect 4836 5147 4843 5183
rect 4896 5167 4903 5196
rect 4956 5176 4983 5183
rect 4836 4943 4843 5093
rect 4896 4956 4903 4993
rect 4836 4936 4863 4943
rect 4936 4707 4943 5163
rect 4976 5143 4983 5176
rect 4996 5163 5003 5393
rect 5116 5347 5123 5403
rect 5156 5387 5163 5403
rect 5196 5396 5203 5433
rect 4996 5156 5023 5163
rect 5056 5156 5063 5213
rect 4976 5136 5003 5143
rect 4956 4947 4963 4993
rect 4996 4987 5003 5136
rect 5016 4987 5023 5156
rect 4976 4956 4983 4973
rect 5036 4936 5043 5113
rect 5076 5067 5083 5143
rect 5096 5123 5103 5333
rect 5136 5127 5143 5143
rect 5156 5127 5163 5373
rect 5176 5156 5183 5173
rect 5096 5116 5123 5123
rect 5196 5067 5203 5213
rect 5236 5203 5243 5403
rect 5256 5387 5263 5436
rect 5276 5427 5283 5453
rect 5316 5436 5323 5473
rect 5296 5416 5303 5433
rect 5276 5207 5283 5413
rect 5336 5403 5343 5423
rect 5376 5403 5383 5433
rect 5456 5423 5463 5433
rect 5436 5416 5463 5423
rect 5336 5396 5383 5403
rect 5236 5196 5263 5203
rect 5256 5176 5263 5196
rect 5296 5176 5303 5353
rect 5356 5176 5363 5193
rect 5076 5047 5083 5053
rect 5096 4976 5103 4993
rect 5056 4956 5083 4963
rect 5116 4956 5123 4973
rect 5056 4847 5063 4956
rect 4996 4696 5003 4713
rect 5016 4707 5023 4773
rect 4836 4676 4843 4693
rect 4876 4647 4883 4663
rect 4836 4456 4843 4633
rect 4916 4503 4923 4693
rect 4976 4667 4983 4683
rect 5016 4627 5023 4673
rect 5096 4647 5103 4683
rect 5116 4627 5123 4833
rect 5136 4787 5143 4973
rect 4916 4496 4943 4503
rect 4816 4387 4823 4443
rect 4856 4407 4863 4443
rect 4916 4307 4923 4463
rect 4936 4207 4943 4496
rect 5016 4427 5023 4613
rect 4756 4196 4783 4203
rect 4756 4067 4763 4196
rect 4776 4187 4783 4196
rect 4796 4087 4803 4193
rect 5036 4147 5043 4513
rect 4896 4016 4903 4093
rect 4756 3947 4763 4013
rect 4916 3787 4923 4073
rect 4876 3736 4883 3773
rect 4996 3767 5003 4053
rect 5076 4003 5083 4613
rect 5096 4447 5103 4573
rect 5116 4467 5123 4593
rect 5136 4527 5143 4713
rect 5156 4687 5163 5053
rect 5196 4943 5203 5033
rect 5176 4936 5203 4943
rect 5136 4456 5143 4493
rect 5156 4476 5163 4633
rect 5176 4507 5183 4936
rect 5196 4667 5203 4913
rect 5176 4447 5183 4463
rect 5096 4227 5103 4433
rect 5116 4207 5123 4333
rect 5136 4087 5143 4373
rect 5156 4247 5163 4313
rect 5176 4267 5183 4433
rect 5156 4196 5163 4233
rect 5076 3996 5103 4003
rect 5016 3976 5043 3983
rect 5036 3847 5043 3976
rect 5076 3963 5083 3973
rect 5056 3956 5083 3963
rect 4916 3736 4923 3753
rect 4896 3707 4903 3723
rect 4436 3216 4463 3223
rect 4316 3196 4343 3203
rect 4316 3036 4323 3053
rect 4356 3036 4363 3073
rect 4296 2667 4303 3033
rect 4376 3016 4383 3033
rect 4316 2607 4323 2763
rect 4336 2727 4343 3013
rect 4416 2987 4423 3193
rect 4436 3007 4443 3216
rect 4456 3036 4463 3113
rect 4496 3036 4503 3113
rect 4556 3036 4583 3043
rect 4516 3016 4523 3033
rect 4536 2863 4543 3033
rect 4556 2867 4563 3036
rect 4636 3016 4643 3033
rect 4516 2856 4543 2863
rect 4516 2723 4523 2856
rect 4596 2727 4603 2993
rect 4656 2776 4663 3133
rect 4496 2716 4523 2723
rect 4296 2447 4303 2543
rect 4316 2463 4323 2553
rect 4356 2536 4363 2553
rect 4336 2487 4343 2523
rect 4376 2516 4383 2573
rect 4396 2536 4403 2553
rect 4416 2487 4423 2653
rect 4436 2567 4443 2653
rect 4476 2583 4483 2633
rect 4476 2576 4503 2583
rect 4436 2543 4443 2553
rect 4496 2547 4503 2576
rect 4516 2563 4523 2673
rect 4516 2556 4543 2563
rect 4556 2556 4563 2613
rect 4616 2583 4623 2763
rect 4596 2576 4623 2583
rect 4436 2536 4463 2543
rect 4496 2487 4503 2533
rect 4536 2527 4543 2556
rect 4316 2456 4343 2463
rect 4076 2096 4083 2113
rect 4036 2076 4063 2083
rect 4016 2047 4023 2063
rect 4036 2047 4043 2076
rect 4116 2056 4123 2133
rect 4136 2087 4143 2253
rect 4176 2143 4183 2293
rect 4316 2207 4323 2243
rect 4336 2187 4343 2456
rect 4176 2136 4203 2143
rect 4016 1927 4023 1973
rect 3996 1827 4003 1913
rect 3956 1767 3963 1783
rect 3856 1656 3883 1663
rect 3896 1663 3903 1753
rect 3936 1747 3943 1763
rect 3896 1656 3923 1663
rect 3856 1627 3863 1656
rect 3876 1616 3883 1633
rect 3896 1627 3903 1633
rect 3816 1596 3863 1603
rect 3816 1576 3843 1583
rect 3676 1383 3683 1533
rect 3656 1376 3683 1383
rect 3636 1227 3643 1273
rect 3656 1267 3663 1376
rect 3676 1147 3683 1333
rect 3616 836 3623 913
rect 3636 867 3643 1053
rect 3656 1027 3663 1103
rect 3696 1067 3703 1373
rect 3716 1327 3723 1413
rect 3776 1387 3783 1533
rect 3816 1487 3823 1533
rect 3836 1507 3843 1576
rect 3876 1527 3883 1573
rect 3816 1467 3823 1473
rect 3836 1467 3843 1493
rect 3716 1007 3723 1273
rect 3736 927 3743 1253
rect 3756 1143 3763 1293
rect 3796 1283 3803 1313
rect 3776 1276 3803 1283
rect 3776 1167 3783 1276
rect 3816 1247 3823 1413
rect 3756 1136 3783 1143
rect 3756 1047 3763 1103
rect 3776 1067 3783 1136
rect 3796 1116 3803 1213
rect 3816 1187 3823 1213
rect 3856 1143 3863 1493
rect 3876 1347 3883 1353
rect 3876 1316 3883 1333
rect 3916 1287 3923 1656
rect 3936 1487 3943 1633
rect 3976 1623 3983 1633
rect 3996 1623 4003 1753
rect 4016 1743 4023 1773
rect 4036 1763 4043 2033
rect 4056 1827 4063 1933
rect 4076 1796 4083 1813
rect 4096 1763 4103 1833
rect 4116 1816 4123 1853
rect 4156 1816 4163 2093
rect 4176 2047 4183 2113
rect 4196 2067 4203 2136
rect 4216 2076 4223 2173
rect 4256 2096 4263 2153
rect 4356 2076 4363 2193
rect 4276 2027 4283 2063
rect 4336 2007 4343 2063
rect 4036 1756 4063 1763
rect 4076 1756 4103 1763
rect 4016 1736 4043 1743
rect 3976 1616 4003 1623
rect 3956 1567 3963 1583
rect 3976 1576 4003 1583
rect 3976 1467 3983 1576
rect 3976 1347 3983 1453
rect 3996 1327 4003 1513
rect 4016 1447 4023 1553
rect 4036 1507 4043 1736
rect 4056 1576 4063 1613
rect 4076 1587 4083 1756
rect 4136 1747 4143 1803
rect 4116 1647 4123 1733
rect 4176 1643 4183 1993
rect 4256 1867 4263 1973
rect 4396 1963 4403 2173
rect 4416 1987 4423 2433
rect 4496 2107 4503 2453
rect 4516 2147 4523 2333
rect 4536 2307 4543 2513
rect 4576 2467 4583 2553
rect 4596 2547 4603 2576
rect 4636 2556 4643 2693
rect 4676 2663 4683 3053
rect 4716 3043 4723 3353
rect 4776 3256 4803 3263
rect 4796 3227 4803 3256
rect 4816 3247 4823 3353
rect 4876 3247 4883 3393
rect 4796 3147 4803 3213
rect 4836 3067 4843 3233
rect 4916 3223 4923 3373
rect 4936 3267 4943 3753
rect 4976 3716 4983 3733
rect 5016 3707 5023 3723
rect 4996 3647 5003 3703
rect 4956 3496 4983 3503
rect 4976 3367 4983 3496
rect 4996 3343 5003 3483
rect 5016 3387 5023 3673
rect 5036 3667 5043 3813
rect 5056 3687 5063 3933
rect 5096 3787 5103 3996
rect 5116 3947 5123 4053
rect 5116 3883 5123 3933
rect 5116 3876 5143 3883
rect 5096 3763 5103 3773
rect 5076 3756 5103 3763
rect 5076 3723 5083 3756
rect 5076 3716 5103 3723
rect 5136 3716 5143 3876
rect 5156 3743 5163 4093
rect 5176 4067 5183 4253
rect 5196 4107 5203 4193
rect 5196 3747 5203 4033
rect 5156 3736 5183 3743
rect 5036 3487 5043 3653
rect 5056 3516 5063 3533
rect 5176 3523 5183 3736
rect 5216 3643 5223 4953
rect 5236 4727 5243 5033
rect 5276 4987 5283 5163
rect 5376 5047 5383 5163
rect 5416 5147 5423 5413
rect 5476 5387 5483 5453
rect 5596 5416 5603 5453
rect 5576 5227 5583 5403
rect 5536 5143 5543 5213
rect 5616 5143 5623 5393
rect 5516 5127 5523 5143
rect 5536 5136 5563 5143
rect 5596 5136 5623 5143
rect 5676 5007 5683 5143
rect 5436 4976 5463 4983
rect 5256 4936 5283 4943
rect 5276 4903 5283 4936
rect 5456 4927 5463 4976
rect 5256 4896 5283 4903
rect 5256 4683 5263 4896
rect 5236 4676 5263 4683
rect 5236 4607 5243 4676
rect 5236 4496 5243 4513
rect 5276 4507 5283 4713
rect 5416 4607 5423 4643
rect 5436 4523 5443 4713
rect 5416 4516 5443 4523
rect 5256 4387 5263 4453
rect 5276 4407 5283 4493
rect 5336 4476 5363 4483
rect 5356 4467 5363 4476
rect 5396 4463 5403 4493
rect 5376 4456 5403 4463
rect 5236 4187 5243 4203
rect 5256 4127 5263 4353
rect 5236 4016 5243 4073
rect 5256 3996 5263 4093
rect 5276 4007 5283 4213
rect 5416 4207 5423 4516
rect 5436 4476 5443 4493
rect 5476 4476 5483 4593
rect 5456 4427 5463 4463
rect 5496 4456 5503 4493
rect 5416 4127 5423 4163
rect 5236 3727 5243 3773
rect 5276 3767 5283 3993
rect 5256 3723 5263 3753
rect 5256 3716 5283 3723
rect 5216 3636 5243 3643
rect 5156 3516 5183 3523
rect 5076 3487 5083 3503
rect 5116 3496 5143 3503
rect 5036 3423 5043 3453
rect 5036 3416 5063 3423
rect 4976 3336 5003 3343
rect 4976 3307 4983 3336
rect 4976 3227 4983 3293
rect 4856 3207 4863 3223
rect 4896 3216 4923 3223
rect 4856 3187 4863 3193
rect 4716 3036 4743 3043
rect 4696 3003 4703 3033
rect 4736 3027 4743 3036
rect 4776 3016 4803 3023
rect 4696 2996 4723 3003
rect 4796 2987 4803 3016
rect 4836 3007 4843 3023
rect 4696 2767 4703 2793
rect 4736 2747 4743 2763
rect 4676 2656 4703 2663
rect 4676 2556 4683 2633
rect 4616 2536 4623 2553
rect 4596 2427 4603 2533
rect 4656 2523 4663 2543
rect 4656 2516 4683 2523
rect 4676 2487 4683 2516
rect 4556 2307 4563 2413
rect 4556 2127 4563 2293
rect 4596 2287 4603 2413
rect 4676 2203 4683 2473
rect 4696 2307 4703 2656
rect 4736 2447 4743 2713
rect 4776 2647 4783 2773
rect 4796 2667 4803 2953
rect 4856 2823 4863 3013
rect 4896 2987 4903 3013
rect 4916 2927 4923 3216
rect 5056 3223 5063 3416
rect 5136 3407 5143 3496
rect 5136 3283 5143 3353
rect 5156 3303 5163 3516
rect 5196 3496 5203 3533
rect 5176 3367 5183 3483
rect 5156 3296 5183 3303
rect 5136 3276 5163 3283
rect 4996 3207 5003 3223
rect 5036 3216 5063 3223
rect 4936 3003 4943 3053
rect 5016 3047 5023 3203
rect 5016 3003 5023 3033
rect 5036 3007 5043 3216
rect 5096 3207 5103 3243
rect 5116 3147 5123 3263
rect 5156 3256 5163 3276
rect 5076 3016 5083 3053
rect 5116 3027 5123 3133
rect 5156 3056 5163 3133
rect 5136 3007 5143 3023
rect 4936 2996 4963 3003
rect 4996 2996 5023 3003
rect 4856 2816 4883 2823
rect 4816 2776 4823 2793
rect 4856 2776 4863 2793
rect 4836 2747 4843 2763
rect 4816 2727 4823 2733
rect 4876 2627 4883 2816
rect 4896 2747 4903 2833
rect 4916 2783 4923 2853
rect 4956 2847 4963 2996
rect 5056 2967 5063 3003
rect 4916 2776 4943 2783
rect 4976 2776 5003 2783
rect 4916 2747 4923 2776
rect 4996 2727 5003 2776
rect 5036 2756 5043 2773
rect 5096 2763 5103 2973
rect 5076 2756 5103 2763
rect 5156 2756 5163 2773
rect 5176 2767 5183 3296
rect 5216 3236 5223 3273
rect 5196 2756 5223 2763
rect 4776 2367 4783 2613
rect 4856 2327 4863 2513
rect 5016 2507 5023 2733
rect 5056 2607 5063 2743
rect 5036 2576 5083 2583
rect 5036 2567 5043 2576
rect 5076 2567 5083 2576
rect 5056 2536 5063 2553
rect 4656 2196 4683 2203
rect 4476 2076 4483 2093
rect 4516 2076 4523 2093
rect 4396 1956 4423 1963
rect 4276 1843 4283 1873
rect 4256 1836 4283 1843
rect 4236 1816 4243 1833
rect 4216 1783 4223 1803
rect 4256 1783 4263 1836
rect 4216 1776 4263 1783
rect 4196 1727 4203 1753
rect 4276 1747 4283 1813
rect 4296 1787 4303 1853
rect 4316 1767 4323 1833
rect 4356 1796 4363 1853
rect 4396 1796 4403 1833
rect 4416 1787 4423 1956
rect 4456 1847 4463 2073
rect 4536 2043 4543 2093
rect 4576 2056 4583 2073
rect 4536 2036 4563 2043
rect 4436 1783 4443 1833
rect 4436 1776 4463 1783
rect 4176 1636 4203 1643
rect 4196 1627 4203 1636
rect 4236 1627 4243 1693
rect 4096 1587 4103 1593
rect 4136 1567 4143 1613
rect 4216 1596 4243 1603
rect 4116 1507 4123 1563
rect 3936 1316 3963 1323
rect 3836 1136 3863 1143
rect 3756 947 3763 1013
rect 3676 847 3683 863
rect 3716 856 3723 873
rect 3736 847 3743 873
rect 3656 823 3663 843
rect 3696 827 3703 843
rect 3756 827 3763 933
rect 3596 807 3603 823
rect 3636 816 3683 823
rect 3527 636 3543 643
rect 3536 616 3543 636
rect 3496 47 3503 573
rect 3516 187 3523 553
rect 3556 527 3563 603
rect 3536 267 3543 433
rect 3576 287 3583 653
rect 3656 647 3663 693
rect 3596 567 3603 613
rect 3656 587 3663 603
rect 3596 387 3603 533
rect 3596 356 3603 373
rect 3516 123 3523 153
rect 3556 136 3563 173
rect 3576 167 3583 273
rect 3516 116 3543 123
rect 3576 107 3583 113
rect 3596 87 3603 193
rect 3616 136 3623 333
rect 3636 307 3643 473
rect 3656 367 3663 533
rect 3676 347 3683 816
rect 3696 647 3703 673
rect 3656 147 3663 153
rect 3696 127 3703 393
rect 3676 107 3683 123
rect 3556 -24 3563 73
rect 3596 -24 3603 33
rect 3716 27 3723 673
rect 3776 663 3783 953
rect 3796 887 3803 1053
rect 3836 983 3843 1136
rect 3896 1127 3903 1283
rect 3936 1247 3943 1316
rect 3976 1207 3983 1283
rect 3936 1143 3943 1173
rect 3996 1167 4003 1293
rect 3916 1136 3943 1143
rect 3856 1116 3883 1123
rect 3876 1087 3883 1116
rect 3816 976 3843 983
rect 3816 847 3823 976
rect 3836 856 3843 953
rect 3876 907 3883 1073
rect 3796 707 3803 823
rect 3856 667 3863 823
rect 3876 747 3883 873
rect 3776 656 3803 663
rect 3756 636 3783 643
rect 3736 527 3743 593
rect 3756 527 3763 573
rect 3776 567 3783 636
rect 3796 487 3803 656
rect 3876 647 3883 733
rect 3896 687 3903 993
rect 3916 827 3923 1136
rect 3936 1116 3983 1123
rect 3996 1116 4003 1133
rect 3956 1067 3963 1083
rect 3956 1047 3963 1053
rect 3976 947 3983 1116
rect 4016 947 4023 1253
rect 4036 1167 4043 1393
rect 4056 1267 4063 1323
rect 4096 1316 4103 1393
rect 4116 1347 4123 1473
rect 4156 1387 4163 1573
rect 4176 1567 4183 1573
rect 4196 1567 4203 1583
rect 4207 1556 4223 1563
rect 4176 1367 4183 1553
rect 4056 1147 4063 1153
rect 4036 1123 4043 1133
rect 4076 1127 4083 1303
rect 4136 1227 4143 1293
rect 4156 1267 4163 1343
rect 4196 1336 4203 1493
rect 4216 1463 4223 1556
rect 4236 1527 4243 1596
rect 4236 1487 4243 1513
rect 4216 1456 4243 1463
rect 4236 1387 4243 1456
rect 4256 1427 4263 1593
rect 4216 1327 4223 1373
rect 4236 1347 4243 1373
rect 4276 1347 4283 1593
rect 4296 1576 4303 1633
rect 4316 1596 4323 1733
rect 4356 1623 4363 1733
rect 4376 1647 4383 1763
rect 4356 1616 4383 1623
rect 4376 1587 4383 1616
rect 4316 1367 4323 1553
rect 4236 1247 4243 1313
rect 4036 1116 4063 1123
rect 4056 1103 4063 1116
rect 4096 1116 4103 1173
rect 4136 1116 4143 1153
rect 4196 1116 4203 1133
rect 4056 1096 4083 1103
rect 4036 1087 4043 1093
rect 3956 847 3963 863
rect 3996 856 4003 873
rect 4036 863 4043 1053
rect 4056 1027 4063 1096
rect 4176 1087 4183 1103
rect 4216 1096 4223 1153
rect 4256 1147 4263 1303
rect 4076 967 4083 1013
rect 4036 856 4063 863
rect 4096 856 4103 873
rect 3936 767 3943 843
rect 3976 807 3983 843
rect 4036 827 4043 856
rect 3956 767 3963 793
rect 3856 596 3863 633
rect 3876 616 3883 633
rect 3896 587 3903 603
rect 3916 507 3923 753
rect 3936 607 3943 653
rect 3956 636 3963 673
rect 3996 667 4003 813
rect 3976 587 3983 623
rect 4016 587 4023 623
rect 3756 207 3763 473
rect 4016 407 4023 573
rect 4036 447 4043 733
rect 4076 707 4083 843
rect 4116 747 4123 933
rect 4196 927 4203 1073
rect 4176 856 4183 873
rect 4196 867 4203 913
rect 4176 627 4183 793
rect 4216 667 4223 833
rect 4236 807 4243 1133
rect 4276 1096 4283 1113
rect 4147 616 4163 623
rect 4196 616 4203 633
rect 4056 587 4063 603
rect 4216 587 4223 603
rect 4236 567 4243 633
rect 4256 463 4263 933
rect 4276 856 4283 1053
rect 4296 967 4303 1083
rect 4316 947 4323 1273
rect 4336 887 4343 1583
rect 4396 1563 4403 1613
rect 4416 1583 4423 1753
rect 4476 1667 4483 1773
rect 4496 1767 4503 2033
rect 4516 1747 4523 1783
rect 4536 1723 4543 2013
rect 4596 1967 4603 2043
rect 4556 1827 4563 1953
rect 4616 1887 4623 2133
rect 4656 2087 4663 2196
rect 4656 2047 4663 2073
rect 4676 2056 4683 2093
rect 4696 2076 4703 2243
rect 4736 2076 4743 2093
rect 4716 2047 4723 2063
rect 4636 1816 4643 2013
rect 4756 2007 4763 2053
rect 4556 1796 4583 1803
rect 4556 1747 4563 1796
rect 4516 1716 4543 1723
rect 4516 1596 4523 1716
rect 4416 1576 4443 1583
rect 4396 1556 4423 1563
rect 4356 1327 4363 1553
rect 4356 1047 4363 1293
rect 4376 1127 4383 1553
rect 4416 1507 4423 1556
rect 4396 1287 4403 1353
rect 4416 1347 4423 1493
rect 4456 1407 4463 1573
rect 4496 1527 4503 1583
rect 4556 1507 4563 1733
rect 4576 1587 4583 1773
rect 4596 1747 4603 1793
rect 4616 1667 4623 1803
rect 4656 1747 4663 1893
rect 4676 1807 4683 1913
rect 4696 1796 4703 1813
rect 4616 1647 4623 1653
rect 4636 1616 4643 1733
rect 4676 1687 4683 1763
rect 4596 1596 4623 1603
rect 4436 1327 4443 1393
rect 4396 1136 4403 1253
rect 4416 1116 4423 1153
rect 4436 1007 4443 1233
rect 4296 687 4303 833
rect 4316 807 4323 863
rect 4336 827 4343 843
rect 4316 507 4323 623
rect 4356 607 4363 993
rect 4376 767 4383 843
rect 4396 827 4403 863
rect 4436 856 4443 933
rect 4416 803 4423 843
rect 4407 796 4423 803
rect 4376 467 4383 733
rect 4236 456 4263 463
rect 4076 376 4083 393
rect 4136 367 4143 433
rect 3736 123 3743 173
rect 3776 136 3783 153
rect 3856 136 3863 173
rect 3736 116 3763 123
rect 3896 123 3903 153
rect 3936 127 3943 143
rect 4016 136 4023 353
rect 4036 307 4043 363
rect 4216 327 4223 363
rect 4236 223 4243 456
rect 4396 447 4403 793
rect 4456 747 4463 1273
rect 4476 1127 4483 1493
rect 4496 1387 4503 1393
rect 4496 1316 4503 1373
rect 4516 1227 4523 1333
rect 4576 1247 4583 1573
rect 4596 1527 4603 1596
rect 4596 1287 4603 1493
rect 4616 1247 4623 1303
rect 4656 1267 4663 1303
rect 4476 1096 4493 1103
rect 4476 847 4483 1096
rect 4516 1076 4523 1193
rect 4676 1187 4683 1653
rect 4696 1507 4703 1673
rect 4716 1627 4723 1833
rect 4736 1727 4743 1933
rect 4756 1647 4763 1993
rect 4776 1867 4783 2113
rect 4796 2076 4803 2133
rect 4816 1847 4823 2173
rect 4856 1987 4863 2313
rect 4876 2247 4883 2283
rect 4836 1816 4843 1953
rect 4776 1787 4783 1803
rect 4796 1687 4803 1793
rect 4816 1783 4823 1803
rect 4856 1783 4863 1813
rect 4816 1776 4863 1783
rect 4716 1567 4723 1613
rect 4756 1576 4763 1593
rect 4736 1547 4743 1563
rect 4716 1507 4723 1533
rect 4716 1316 4723 1473
rect 4736 1307 4743 1533
rect 4756 1287 4763 1333
rect 4796 1327 4803 1633
rect 4836 1616 4843 1776
rect 4856 1687 4863 1753
rect 4876 1647 4883 2233
rect 4896 2187 4903 2433
rect 4916 2147 4923 2353
rect 4896 1907 4903 2093
rect 4896 1707 4903 1853
rect 4916 1847 4923 2113
rect 4936 2103 4943 2393
rect 5016 2247 5023 2433
rect 5036 2147 5043 2533
rect 5096 2483 5103 2733
rect 5076 2476 5103 2483
rect 5076 2287 5083 2476
rect 5116 2287 5123 2753
rect 5196 2723 5203 2756
rect 5236 2747 5243 3636
rect 5256 3487 5263 3513
rect 5256 2747 5263 3433
rect 5276 3407 5283 3503
rect 5296 3447 5303 3953
rect 5316 3827 5323 4073
rect 5336 3927 5343 4093
rect 5356 3996 5363 4033
rect 5396 3996 5403 4053
rect 5416 3967 5423 4093
rect 5436 3987 5443 4413
rect 5516 4367 5523 4833
rect 5536 4727 5543 4993
rect 5616 4956 5643 4963
rect 5676 4956 5683 4973
rect 5696 4967 5703 5153
rect 5576 4916 5603 4923
rect 5576 4703 5583 4916
rect 5616 4907 5623 4956
rect 5656 4847 5663 4943
rect 5696 4936 5703 4953
rect 5556 4696 5583 4703
rect 5536 4667 5543 4683
rect 5556 4587 5563 4696
rect 5547 4476 5563 4483
rect 5596 4476 5603 4493
rect 5516 4203 5523 4313
rect 5536 4283 5543 4473
rect 5576 4447 5583 4463
rect 5616 4456 5623 4673
rect 5536 4276 5563 4283
rect 5516 4196 5543 4203
rect 5496 3996 5503 4113
rect 5516 3976 5523 3993
rect 5536 3823 5543 4053
rect 5556 4047 5563 4276
rect 5576 3996 5583 4033
rect 5596 4027 5603 4233
rect 5616 4047 5623 4413
rect 5636 4183 5643 4633
rect 5696 4427 5703 4893
rect 5716 4243 5723 4973
rect 5736 4807 5743 4933
rect 5736 4667 5743 4793
rect 5736 4307 5743 4313
rect 5716 4236 5743 4243
rect 5696 4216 5723 4223
rect 5636 4176 5663 4183
rect 5596 3947 5603 3983
rect 5636 3976 5643 4013
rect 5656 3943 5663 4176
rect 5676 4067 5683 4203
rect 5716 4183 5723 4216
rect 5696 4176 5723 4183
rect 5636 3936 5663 3943
rect 5536 3816 5563 3823
rect 5456 3647 5463 3683
rect 5316 3243 5323 3493
rect 5556 3347 5563 3816
rect 5616 3736 5623 3753
rect 5296 3236 5323 3243
rect 5296 3023 5303 3236
rect 5476 3127 5483 3203
rect 5496 3103 5503 3333
rect 5616 3287 5623 3393
rect 5636 3383 5643 3936
rect 5656 3547 5663 3853
rect 5656 3407 5663 3453
rect 5636 3376 5663 3383
rect 5636 3263 5643 3293
rect 5616 3256 5643 3263
rect 5476 3096 5503 3103
rect 5276 3016 5303 3023
rect 5296 2803 5303 3016
rect 5276 2796 5303 2803
rect 5276 2763 5283 2796
rect 5476 2763 5483 3096
rect 5596 3023 5603 3243
rect 5616 3043 5623 3256
rect 5616 3036 5643 3043
rect 5576 3016 5603 3023
rect 5276 2756 5303 2763
rect 5476 2756 5503 2763
rect 5187 2716 5203 2723
rect 5276 2587 5283 2756
rect 5196 2556 5223 2563
rect 5136 2527 5143 2543
rect 5196 2487 5203 2556
rect 5276 2536 5283 2553
rect 5296 2527 5303 2733
rect 5476 2707 5483 2723
rect 5316 2523 5323 2553
rect 5356 2536 5363 2553
rect 5396 2547 5403 2613
rect 5316 2516 5343 2523
rect 5136 2387 5143 2473
rect 5056 2127 5063 2253
rect 5096 2247 5103 2263
rect 5076 2227 5083 2243
rect 4936 2096 4983 2103
rect 4936 2007 4943 2063
rect 4936 1847 4943 1873
rect 4956 1823 4963 1873
rect 4976 1847 4983 2096
rect 4996 1827 5003 2073
rect 5036 2056 5043 2113
rect 5076 2067 5083 2133
rect 5096 1967 5103 2233
rect 5116 2167 5123 2273
rect 5136 2207 5143 2373
rect 5156 2227 5163 2263
rect 5196 2187 5203 2263
rect 5216 2247 5223 2293
rect 5236 2267 5243 2353
rect 5116 2107 5123 2153
rect 5136 2096 5143 2173
rect 5116 2076 5123 2093
rect 4956 1816 4983 1823
rect 4836 1487 4843 1573
rect 4536 1096 4543 1133
rect 4556 1067 4563 1083
rect 4496 1047 4503 1053
rect 4496 807 4503 973
rect 4576 963 4583 1133
rect 4656 1096 4663 1133
rect 4596 987 4603 1073
rect 4576 956 4603 963
rect 4536 836 4543 853
rect 4596 827 4603 956
rect 4656 856 4663 933
rect 4676 867 4683 1053
rect 4476 636 4483 653
rect 4416 616 4423 633
rect 4456 607 4463 623
rect 4496 587 4503 673
rect 4536 547 4543 653
rect 4576 636 4583 753
rect 4616 636 4623 693
rect 4636 656 4643 813
rect 4676 767 4683 853
rect 4656 636 4683 643
rect 4556 587 4563 603
rect 4596 587 4603 633
rect 4396 247 4403 323
rect 4216 216 4243 223
rect 3836 107 3843 123
rect 3876 116 3903 123
rect 4216 47 4223 216
rect 4416 187 4423 393
rect 4556 376 4563 393
rect 4436 176 4443 213
rect 4316 136 4323 153
rect 4376 123 4383 173
rect 4476 156 4483 173
rect 4496 147 4503 353
rect 4516 167 4523 363
rect 4556 176 4563 233
rect 4536 156 4543 173
rect 4576 156 4583 173
rect 4616 167 4623 473
rect 4636 156 4643 493
rect 4656 376 4663 573
rect 4676 467 4683 636
rect 4696 423 4703 1213
rect 4776 1147 4783 1293
rect 4816 1207 4823 1303
rect 4836 1287 4843 1323
rect 4716 1096 4743 1103
rect 4716 947 4723 1096
rect 4816 1083 4823 1173
rect 4796 1076 4823 1083
rect 4836 927 4843 1253
rect 4807 876 4813 883
rect 4856 883 4863 1313
rect 4876 1287 4883 1633
rect 4896 1527 4903 1673
rect 4916 1547 4923 1733
rect 4936 1727 4943 1803
rect 4956 1667 4963 1773
rect 4976 1687 4983 1816
rect 4936 1596 4943 1613
rect 4976 1596 4983 1673
rect 4996 1427 5003 1813
rect 5036 1796 5043 1833
rect 5056 1807 5063 1853
rect 5076 1823 5083 1893
rect 5096 1847 5103 1913
rect 5076 1816 5103 1823
rect 5016 1747 5023 1783
rect 5056 1727 5063 1763
rect 5016 1596 5023 1653
rect 5036 1616 5043 1653
rect 5096 1627 5103 1816
rect 5116 1807 5123 2033
rect 5176 1887 5183 2113
rect 5216 2107 5223 2233
rect 5256 2187 5263 2513
rect 5336 2296 5343 2313
rect 5276 2267 5283 2283
rect 5316 2263 5323 2283
rect 5356 2263 5363 2333
rect 5416 2307 5423 2513
rect 5456 2307 5463 2543
rect 5476 2527 5483 2593
rect 5476 2347 5483 2513
rect 5496 2323 5503 2756
rect 5576 2743 5583 2973
rect 5596 2927 5603 3016
rect 5636 3003 5643 3036
rect 5616 2996 5643 3003
rect 5616 2763 5623 2996
rect 5636 2776 5643 2913
rect 5596 2756 5623 2763
rect 5576 2736 5603 2743
rect 5516 2487 5523 2523
rect 5576 2507 5583 2713
rect 5516 2367 5523 2473
rect 5596 2467 5603 2736
rect 5616 2527 5623 2733
rect 5656 2727 5663 3376
rect 5636 2443 5643 2573
rect 5616 2436 5643 2443
rect 5476 2316 5503 2323
rect 5376 2283 5383 2293
rect 5376 2276 5403 2283
rect 5316 2256 5363 2263
rect 5207 2076 5223 2083
rect 5196 2027 5203 2073
rect 5116 1707 5123 1773
rect 5136 1747 5143 1803
rect 5176 1796 5183 1853
rect 5156 1767 5163 1783
rect 5196 1627 5203 1783
rect 5056 1596 5063 1613
rect 5076 1547 5083 1593
rect 5096 1587 5103 1613
rect 5196 1607 5203 1613
rect 5156 1596 5173 1603
rect 4896 1307 4903 1353
rect 4936 1307 4943 1323
rect 4956 1307 4963 1343
rect 4876 1147 4883 1153
rect 4876 1116 4883 1133
rect 4916 1116 4923 1133
rect 4896 1047 4903 1103
rect 4936 1096 4943 1113
rect 4856 876 4883 883
rect 4756 856 4783 863
rect 4736 827 4743 843
rect 4776 807 4783 856
rect 4796 856 4823 863
rect 4796 827 4803 856
rect 4716 627 4723 793
rect 4776 787 4783 793
rect 4796 787 4803 793
rect 4836 707 4843 843
rect 4736 636 4743 693
rect 4796 636 4803 673
rect 4776 467 4783 623
rect 4696 416 4723 423
rect 4696 376 4703 393
rect 4716 387 4723 416
rect 4736 367 4743 453
rect 4767 396 4783 403
rect 4776 376 4783 396
rect 4796 307 4803 363
rect 4416 127 4423 133
rect 4356 116 4383 123
rect 4696 107 4703 213
rect 4716 127 4723 273
rect 4756 136 4763 153
rect 4796 123 4803 133
rect 4736 107 4743 123
rect 4776 116 4803 123
rect 4816 107 4823 373
rect 4836 287 4843 363
rect 4856 347 4863 753
rect 4876 627 4883 876
rect 4876 527 4883 613
rect 4876 327 4883 353
rect 4896 307 4903 873
rect 4916 856 4923 913
rect 4956 887 4963 1133
rect 4976 1107 4983 1273
rect 4936 787 4943 843
rect 4936 616 4943 633
rect 4916 583 4923 593
rect 4916 576 4943 583
rect 4916 356 4923 413
rect 4856 136 4863 153
rect 4936 147 4943 576
rect 4956 547 4963 603
rect 4976 367 4983 1093
rect 4996 1087 5003 1393
rect 5136 1343 5143 1573
rect 5116 1336 5143 1343
rect 5016 1227 5023 1313
rect 5036 1287 5043 1323
rect 5036 1136 5043 1213
rect 5016 1116 5023 1133
rect 5056 1116 5063 1153
rect 5076 967 5083 1233
rect 5096 1087 5103 1153
rect 5116 1147 5123 1336
rect 5136 1136 5143 1293
rect 5156 1207 5163 1283
rect 5176 1227 5183 1303
rect 5156 1116 5163 1153
rect 5196 1143 5203 1333
rect 5216 1167 5223 1913
rect 5256 1727 5263 1973
rect 5236 1307 5243 1673
rect 5276 1596 5283 1773
rect 5296 1627 5303 2233
rect 5416 2227 5423 2263
rect 5456 2207 5463 2263
rect 5316 1907 5323 2073
rect 5376 2036 5383 2113
rect 5416 2087 5423 2193
rect 5476 2163 5483 2316
rect 5516 2307 5523 2353
rect 5496 2247 5503 2293
rect 5536 2287 5543 2313
rect 5456 2156 5483 2163
rect 5396 2056 5423 2063
rect 5416 2007 5423 2056
rect 5376 1763 5383 1893
rect 5396 1807 5403 1993
rect 5456 1927 5463 2156
rect 5476 2107 5483 2133
rect 5496 2103 5503 2213
rect 5516 2123 5523 2233
rect 5536 2207 5543 2243
rect 5556 2187 5563 2263
rect 5576 2227 5583 2293
rect 5616 2287 5623 2436
rect 5596 2207 5603 2263
rect 5616 2227 5623 2243
rect 5516 2116 5543 2123
rect 5496 2096 5523 2103
rect 5476 2076 5483 2093
rect 5476 1947 5483 2033
rect 5496 1987 5503 2053
rect 5516 2007 5523 2096
rect 5536 1907 5543 2116
rect 5556 2087 5563 2133
rect 5576 2056 5583 2113
rect 5596 2007 5603 2043
rect 5376 1756 5403 1763
rect 5356 1627 5363 1713
rect 5376 1616 5383 1713
rect 5396 1683 5403 1733
rect 5396 1676 5423 1683
rect 5256 1587 5263 1593
rect 5256 1367 5263 1533
rect 5256 1316 5263 1353
rect 5196 1136 5223 1143
rect 4996 607 5003 953
rect 5016 767 5023 893
rect 5036 667 5043 913
rect 5176 847 5183 1133
rect 5196 1087 5203 1103
rect 5216 1027 5223 1136
rect 5236 1127 5243 1293
rect 5296 1227 5303 1303
rect 5316 1267 5323 1273
rect 5336 1247 5343 1613
rect 5396 1607 5403 1653
rect 5376 1316 5383 1513
rect 5396 1287 5403 1553
rect 5416 1347 5423 1676
rect 5436 1567 5443 1693
rect 5416 1247 5423 1303
rect 5456 1207 5463 1693
rect 5496 1603 5503 1673
rect 5476 1596 5503 1603
rect 5476 1467 5483 1596
rect 5236 867 5243 1113
rect 5056 643 5063 793
rect 5076 787 5083 803
rect 5096 767 5103 823
rect 5156 767 5163 823
rect 5076 667 5083 673
rect 5056 636 5083 643
rect 5116 636 5123 673
rect 5056 623 5063 636
rect 5016 616 5063 623
rect 5136 616 5143 673
rect 4896 123 4903 133
rect 4876 116 4903 123
rect 4976 123 4983 293
rect 5016 136 5023 533
rect 5056 403 5063 593
rect 5056 396 5083 403
rect 5076 327 5083 396
rect 5116 363 5123 593
rect 5156 487 5163 653
rect 5176 636 5183 753
rect 5196 667 5203 823
rect 5236 807 5243 853
rect 5256 847 5263 1153
rect 5456 1136 5463 1173
rect 5476 1087 5483 1413
rect 5496 1336 5503 1553
rect 5516 1507 5523 1583
rect 5536 1567 5543 1833
rect 5556 1707 5563 1973
rect 5576 1847 5583 1893
rect 5596 1807 5603 1953
rect 5576 1647 5583 1803
rect 5576 1596 5583 1613
rect 5596 1507 5603 1793
rect 5616 1587 5623 2193
rect 5636 1727 5643 2233
rect 5656 2107 5663 2493
rect 5676 2447 5683 4033
rect 5696 3527 5703 4176
rect 5696 3307 5703 3483
rect 5696 2747 5703 3273
rect 5716 2987 5723 4153
rect 5736 3867 5743 4236
rect 5736 3727 5743 3833
rect 5736 3387 5743 3493
rect 5716 2927 5723 2933
rect 5716 2576 5723 2593
rect 5676 2096 5683 2253
rect 5696 2207 5703 2513
rect 5716 2487 5723 2533
rect 5696 2076 5703 2153
rect 5676 1687 5683 2013
rect 5696 1947 5703 2033
rect 5696 1627 5703 1933
rect 5536 1207 5543 1343
rect 5556 1107 5563 1323
rect 5576 1096 5583 1433
rect 5616 1316 5623 1473
rect 5696 1367 5703 1573
rect 5656 1316 5663 1333
rect 5636 1267 5643 1303
rect 5296 856 5323 863
rect 5256 767 5263 833
rect 5296 647 5303 856
rect 5236 616 5243 633
rect 5096 356 5123 363
rect 5056 136 5063 293
rect 4956 116 4983 123
rect 4916 107 4923 113
rect 5096 67 5103 356
rect 5116 107 5123 153
rect 5156 136 5163 433
rect 5196 356 5203 473
rect 5256 187 5263 633
rect 5316 627 5323 813
rect 5356 767 5363 863
rect 5376 827 5383 843
rect 5636 836 5643 1113
rect 5696 1107 5703 1333
rect 5716 1127 5723 2453
rect 5736 1567 5743 3353
rect 5736 1327 5743 1353
rect 5736 1307 5743 1313
rect 5736 1136 5743 1293
rect 5756 1227 5763 4673
rect 5336 636 5343 673
rect 5376 636 5383 673
rect 5396 607 5403 823
rect 5436 807 5443 823
rect 5416 783 5423 803
rect 5456 783 5463 813
rect 5596 803 5603 833
rect 5476 787 5483 803
rect 5596 796 5623 803
rect 5416 776 5463 783
rect 5416 636 5423 693
rect 5436 656 5443 673
rect 5456 636 5463 653
rect 5516 636 5523 653
rect 5536 603 5543 693
rect 5636 636 5643 693
rect 5656 656 5663 1093
rect 5676 867 5683 1103
rect 5676 636 5683 833
rect 5536 596 5563 603
rect 5616 387 5623 393
rect 5696 387 5703 1073
rect 5176 107 5183 123
rect 5236 67 5243 143
rect 5316 136 5323 353
rect 5696 127 5703 373
rect 5736 367 5743 473
rect 5736 27 5743 133
rect 3636 -24 3643 13
rect 3836 -24 3843 13
<< m3contact >>
rect 2533 5533 2547 5547
rect 2413 5513 2427 5527
rect 1213 5473 1227 5487
rect 1613 5473 1627 5487
rect 1833 5473 1847 5487
rect 73 5453 87 5467
rect 153 5453 167 5467
rect 193 5453 207 5467
rect 253 5453 267 5467
rect 273 5453 287 5467
rect 513 5453 527 5467
rect 793 5453 807 5467
rect 873 5453 887 5467
rect 913 5453 927 5467
rect 53 5433 67 5447
rect 53 5373 67 5387
rect 93 5373 107 5387
rect 153 5393 167 5407
rect 213 5393 227 5407
rect 173 5353 187 5367
rect 73 5153 87 5167
rect 33 5113 47 5127
rect 193 5173 207 5187
rect 273 5173 287 5187
rect 313 5173 327 5187
rect 133 5113 147 5127
rect 353 5313 367 5327
rect 693 5413 707 5427
rect 813 5413 827 5427
rect 853 5413 867 5427
rect 453 5313 467 5327
rect 433 5153 447 5167
rect 333 5133 347 5147
rect 393 5133 407 5147
rect 173 5113 187 5127
rect 293 5113 307 5127
rect 353 5113 367 5127
rect 113 5073 127 5087
rect 153 5073 167 5087
rect 33 4753 47 4767
rect 93 4713 107 4727
rect 53 4693 67 4707
rect 73 4673 87 4687
rect 193 5033 207 5047
rect 373 5033 387 5047
rect 373 5013 387 5027
rect 393 4973 407 4987
rect 453 4913 467 4927
rect 193 4773 207 4787
rect 393 4773 407 4787
rect 173 4713 187 4727
rect 73 4653 87 4667
rect 113 4653 127 4667
rect 493 5153 507 5167
rect 833 5393 847 5407
rect 773 5113 787 5127
rect 513 5053 527 5067
rect 613 5053 627 5067
rect 493 4973 507 4987
rect 613 4993 627 5007
rect 533 4953 547 4967
rect 653 4953 667 4967
rect 693 4953 707 4967
rect 733 4953 747 4967
rect 873 5153 887 5167
rect 893 5153 907 5167
rect 833 5073 847 5087
rect 793 5033 807 5047
rect 793 5013 807 5027
rect 793 4973 807 4987
rect 713 4933 727 4947
rect 733 4893 747 4907
rect 233 4753 247 4767
rect 473 4753 487 4767
rect 553 4693 567 4707
rect 653 4693 667 4707
rect 133 4633 147 4647
rect 153 4633 167 4647
rect 73 4193 87 4207
rect 273 4653 287 4667
rect 393 4633 407 4647
rect 193 4493 207 4507
rect 633 4673 647 4687
rect 773 4913 787 4927
rect 753 4773 767 4787
rect 573 4593 587 4607
rect 853 4933 867 4947
rect 833 4893 847 4907
rect 793 4873 807 4887
rect 813 4713 827 4727
rect 933 5433 947 5447
rect 973 5393 987 5407
rect 1173 5413 1187 5427
rect 1033 5393 1047 5407
rect 1093 5393 1107 5407
rect 1153 5393 1167 5407
rect 1253 5453 1267 5467
rect 1293 5433 1307 5447
rect 1333 5433 1347 5447
rect 1013 5373 1027 5387
rect 933 5173 947 5187
rect 973 5173 987 5187
rect 993 5173 1007 5187
rect 933 5133 947 5147
rect 953 5113 967 5127
rect 1013 5153 1027 5167
rect 1073 5173 1087 5187
rect 1133 5253 1147 5267
rect 1233 5393 1247 5407
rect 1313 5393 1327 5407
rect 1353 5393 1367 5407
rect 1393 5373 1407 5387
rect 1353 5353 1367 5367
rect 1053 5153 1067 5167
rect 1093 5153 1107 5167
rect 1153 5153 1167 5167
rect 1033 5133 1047 5147
rect 1153 5113 1167 5127
rect 1253 5153 1267 5167
rect 1293 5153 1307 5167
rect 1273 5133 1287 5147
rect 1333 5133 1347 5147
rect 1433 5433 1447 5447
rect 1493 5433 1507 5447
rect 1453 5393 1467 5407
rect 1433 5173 1447 5187
rect 1413 5153 1427 5167
rect 1353 5113 1367 5127
rect 1233 5093 1247 5107
rect 1193 5033 1207 5047
rect 993 4993 1007 5007
rect 1013 4993 1027 5007
rect 973 4973 987 4987
rect 1053 4973 1067 4987
rect 1093 4953 1107 4967
rect 953 4933 967 4947
rect 993 4933 1007 4947
rect 993 4893 1007 4907
rect 953 4713 967 4727
rect 853 4693 867 4707
rect 913 4693 927 4707
rect 953 4693 967 4707
rect 793 4673 807 4687
rect 833 4673 847 4687
rect 753 4513 767 4527
rect 673 4473 687 4487
rect 713 4473 727 4487
rect 753 4473 767 4487
rect 373 4453 387 4467
rect 573 4453 587 4467
rect 533 4433 547 4447
rect 593 4433 607 4447
rect 453 4413 467 4427
rect 853 4653 867 4667
rect 913 4653 927 4667
rect 973 4653 987 4667
rect 893 4633 907 4647
rect 853 4493 867 4507
rect 813 4473 827 4487
rect 653 4393 667 4407
rect 173 4173 187 4187
rect 193 4133 207 4147
rect 193 4013 207 4027
rect 53 3993 67 4007
rect 513 4193 527 4207
rect 633 4193 647 4207
rect 793 4413 807 4427
rect 773 4233 787 4247
rect 773 4193 787 4207
rect 533 4173 547 4187
rect 573 4173 587 4187
rect 473 4153 487 4167
rect 873 4453 887 4467
rect 913 4473 927 4487
rect 953 4453 967 4467
rect 893 4433 907 4447
rect 933 4433 947 4447
rect 1053 4913 1067 4927
rect 1033 4873 1047 4887
rect 1113 4793 1127 4807
rect 1053 4773 1067 4787
rect 1133 4733 1147 4747
rect 1193 4733 1207 4747
rect 1113 4673 1127 4687
rect 1073 4653 1087 4667
rect 1093 4653 1107 4667
rect 1113 4553 1127 4567
rect 1373 4973 1387 4987
rect 1233 4913 1247 4927
rect 1713 5453 1727 5467
rect 1733 5453 1747 5467
rect 1573 5433 1587 5447
rect 1633 5413 1647 5427
rect 1973 5453 1987 5467
rect 2273 5453 2287 5467
rect 2193 5433 2207 5447
rect 1833 5413 1847 5427
rect 1773 5373 1787 5387
rect 1813 5373 1827 5387
rect 1753 5273 1767 5287
rect 1513 5253 1527 5267
rect 1573 5253 1587 5267
rect 1493 5173 1507 5187
rect 1473 5153 1487 5167
rect 1453 5093 1467 5107
rect 1593 5113 1607 5127
rect 1593 5013 1607 5027
rect 1633 5013 1647 5027
rect 1573 4953 1587 4967
rect 1533 4913 1547 4927
rect 1393 4873 1407 4887
rect 1473 4793 1487 4807
rect 1253 4773 1267 4787
rect 1253 4713 1267 4727
rect 1173 4653 1187 4667
rect 1213 4653 1227 4667
rect 1393 4753 1407 4767
rect 1433 4753 1447 4767
rect 1393 4693 1407 4707
rect 1333 4673 1347 4687
rect 1233 4633 1247 4647
rect 1313 4653 1327 4667
rect 1453 4693 1467 4707
rect 1053 4513 1067 4527
rect 1133 4513 1147 4527
rect 1073 4493 1087 4507
rect 1133 4493 1147 4507
rect 1213 4493 1227 4507
rect 1093 4473 1107 4487
rect 1113 4473 1127 4487
rect 893 4413 907 4427
rect 953 4393 967 4407
rect 833 4353 847 4367
rect 833 4333 847 4347
rect 653 4153 667 4167
rect 733 4153 747 4167
rect 753 4153 767 4167
rect 793 4153 807 4167
rect 553 4133 567 4147
rect 553 4013 567 4027
rect 373 3973 387 3987
rect 453 3973 467 3987
rect 593 3973 607 3987
rect 553 3773 567 3787
rect 633 3773 647 3787
rect 133 3733 147 3747
rect 13 3673 27 3687
rect 153 3713 167 3727
rect 233 3733 247 3747
rect 273 3733 287 3747
rect 193 3693 207 3707
rect 213 3673 227 3687
rect 213 3653 227 3667
rect 53 3613 67 3627
rect 113 3613 127 3627
rect 173 3533 187 3547
rect 73 3513 87 3527
rect 113 3493 127 3507
rect 153 3493 167 3507
rect 93 3433 107 3447
rect 53 3413 67 3427
rect 93 3413 107 3427
rect 53 3253 67 3267
rect 133 3473 147 3487
rect 193 3513 207 3527
rect 253 3713 267 3727
rect 353 3713 367 3727
rect 473 3713 487 3727
rect 293 3693 307 3707
rect 293 3533 307 3547
rect 253 3493 267 3507
rect 233 3473 247 3487
rect 313 3473 327 3487
rect 273 3453 287 3467
rect 153 3433 167 3447
rect 113 3353 127 3367
rect 173 3353 187 3367
rect 513 3673 527 3687
rect 573 3673 587 3687
rect 373 3553 387 3567
rect 673 4133 687 4147
rect 933 4213 947 4227
rect 853 4193 867 4207
rect 873 4173 887 4187
rect 1073 4353 1087 4367
rect 1153 4473 1167 4487
rect 1193 4473 1207 4487
rect 1133 4433 1147 4447
rect 1173 4433 1187 4447
rect 1173 4413 1187 4427
rect 993 4213 1007 4227
rect 1053 4213 1067 4227
rect 1073 4213 1087 4227
rect 953 4193 967 4207
rect 973 4173 987 4187
rect 1013 4173 1027 4187
rect 853 4153 867 4167
rect 733 4113 747 4127
rect 833 4113 847 4127
rect 853 4113 867 4127
rect 693 3993 707 4007
rect 713 3993 727 4007
rect 753 4093 767 4107
rect 1013 4113 1027 4127
rect 833 4073 847 4087
rect 893 4073 907 4087
rect 1013 4073 1027 4087
rect 793 4053 807 4067
rect 753 4013 767 4027
rect 673 3773 687 3787
rect 713 3753 727 3767
rect 733 3733 747 3747
rect 713 3693 727 3707
rect 693 3673 707 3687
rect 693 3653 707 3667
rect 673 3633 687 3647
rect 653 3593 667 3607
rect 613 3533 627 3547
rect 573 3513 587 3527
rect 593 3513 607 3527
rect 373 3493 387 3507
rect 413 3493 427 3507
rect 433 3473 447 3487
rect 513 3493 527 3507
rect 553 3493 567 3507
rect 493 3473 507 3487
rect 473 3453 487 3467
rect 533 3453 547 3467
rect 333 3433 347 3447
rect 313 3333 327 3347
rect 433 3333 447 3347
rect 373 3253 387 3267
rect 133 3213 147 3227
rect 153 3213 167 3227
rect 73 3033 87 3047
rect 93 2993 107 3007
rect 53 2973 67 2987
rect 53 2933 67 2947
rect 173 3173 187 3187
rect 293 3233 307 3247
rect 333 3233 347 3247
rect 273 3213 287 3227
rect 313 3193 327 3207
rect 393 3213 407 3227
rect 533 3353 547 3367
rect 633 3493 647 3507
rect 673 3493 687 3507
rect 813 4033 827 4047
rect 913 4053 927 4067
rect 973 4053 987 4067
rect 853 4033 867 4047
rect 893 4033 907 4047
rect 933 4033 947 4047
rect 893 4013 907 4027
rect 913 4013 927 4027
rect 873 3993 887 4007
rect 973 3993 987 4007
rect 1073 4193 1087 4207
rect 1053 4153 1067 4167
rect 1033 4053 1047 4067
rect 1033 4013 1047 4027
rect 1053 3993 1067 4007
rect 913 3953 927 3967
rect 853 3933 867 3947
rect 793 3753 807 3767
rect 773 3733 787 3747
rect 753 3633 767 3647
rect 733 3513 747 3527
rect 733 3493 747 3507
rect 773 3493 787 3507
rect 573 3473 587 3487
rect 613 3473 627 3487
rect 653 3473 667 3487
rect 713 3473 727 3487
rect 553 3273 567 3287
rect 753 3433 767 3447
rect 773 3313 787 3327
rect 833 3733 847 3747
rect 813 3693 827 3707
rect 953 3853 967 3867
rect 913 3713 927 3727
rect 1033 3973 1047 3987
rect 1013 3713 1027 3727
rect 873 3673 887 3687
rect 973 3673 987 3687
rect 853 3613 867 3627
rect 873 3493 887 3507
rect 853 3473 867 3487
rect 993 3513 1007 3527
rect 933 3493 947 3507
rect 973 3493 987 3507
rect 1053 3733 1067 3747
rect 1153 4233 1167 4247
rect 1113 4213 1127 4227
rect 1093 4013 1107 4027
rect 1073 3653 1087 3667
rect 1093 3633 1107 3647
rect 1073 3553 1087 3567
rect 1093 3513 1107 3527
rect 1073 3493 1087 3507
rect 1033 3413 1047 3427
rect 1133 4033 1147 4047
rect 1193 4353 1207 4367
rect 1273 4573 1287 4587
rect 1293 4493 1307 4507
rect 1293 4473 1307 4487
rect 1453 4653 1467 4667
rect 1493 4673 1507 4687
rect 1513 4673 1527 4687
rect 1473 4633 1487 4647
rect 1313 4453 1327 4467
rect 1353 4433 1367 4447
rect 1453 4493 1467 4507
rect 1413 4433 1427 4447
rect 1653 4993 1667 5007
rect 1613 4953 1627 4967
rect 1813 5173 1827 5187
rect 1773 5133 1787 5147
rect 1813 5053 1827 5067
rect 1773 5033 1787 5047
rect 1753 4893 1767 4907
rect 1753 4713 1767 4727
rect 1593 4653 1607 4667
rect 1593 4613 1607 4627
rect 1513 4593 1527 4607
rect 1573 4593 1587 4607
rect 1553 4493 1567 4507
rect 1753 4613 1767 4627
rect 1613 4593 1627 4607
rect 1593 4553 1607 4567
rect 1713 4533 1727 4547
rect 1653 4513 1667 4527
rect 1613 4493 1627 4507
rect 1573 4453 1587 4467
rect 1673 4473 1687 4487
rect 1393 4333 1407 4347
rect 1193 4213 1207 4227
rect 1213 4133 1227 4147
rect 1213 4013 1227 4027
rect 1233 3973 1247 3987
rect 1193 3953 1207 3967
rect 1153 3933 1167 3947
rect 1413 4253 1427 4267
rect 1273 4233 1287 4247
rect 1313 4193 1327 4207
rect 1273 4173 1287 4187
rect 1293 4173 1307 4187
rect 1353 4173 1367 4187
rect 1273 4073 1287 4087
rect 1133 3733 1147 3747
rect 1193 3733 1207 3747
rect 1253 3733 1267 3747
rect 1393 4193 1407 4207
rect 1373 4133 1387 4147
rect 1393 4093 1407 4107
rect 1693 4413 1707 4427
rect 1653 4393 1667 4407
rect 1453 4213 1467 4227
rect 1493 4213 1507 4227
rect 1553 4213 1567 4227
rect 1573 4213 1587 4227
rect 1613 4213 1627 4227
rect 1693 4373 1707 4387
rect 1673 4333 1687 4347
rect 1493 4153 1507 4167
rect 1473 4113 1487 4127
rect 1413 4033 1427 4047
rect 1453 4033 1467 4047
rect 1353 4013 1367 4027
rect 1413 4013 1427 4027
rect 1433 4013 1447 4027
rect 1473 4013 1487 4027
rect 1313 3973 1327 3987
rect 1473 3953 1487 3967
rect 1593 4193 1607 4207
rect 1573 4153 1587 4167
rect 1573 4133 1587 4147
rect 1553 4113 1567 4127
rect 1633 4113 1647 4127
rect 1533 4013 1547 4027
rect 1593 4073 1607 4087
rect 1613 4073 1627 4087
rect 1593 4053 1607 4067
rect 1613 3993 1627 4007
rect 1793 4933 1807 4947
rect 1853 5253 1867 5267
rect 1973 5393 1987 5407
rect 2173 5393 2187 5407
rect 1873 5153 1887 5167
rect 1973 5133 1987 5147
rect 2173 5113 2187 5127
rect 1873 5053 1887 5067
rect 1893 5053 1907 5067
rect 1853 5033 1867 5047
rect 1833 4953 1847 4967
rect 1813 4913 1827 4927
rect 1793 4713 1807 4727
rect 1793 4673 1807 4687
rect 1813 4673 1827 4687
rect 1873 4673 1887 4687
rect 1813 4513 1827 4527
rect 1793 4473 1807 4487
rect 1853 4413 1867 4427
rect 1813 4373 1827 4387
rect 2013 5073 2027 5087
rect 1973 5033 1987 5047
rect 1953 5013 1967 5027
rect 1933 4973 1947 4987
rect 1913 4933 1927 4947
rect 1973 4893 1987 4907
rect 1933 4873 1947 4887
rect 1913 4733 1927 4747
rect 2033 5053 2047 5067
rect 2153 5013 2167 5027
rect 2153 4993 2167 5007
rect 2053 4973 2067 4987
rect 2133 4973 2147 4987
rect 2233 5413 2247 5427
rect 2313 5433 2327 5447
rect 2333 5373 2347 5387
rect 2273 5253 2287 5267
rect 2313 5213 2327 5227
rect 2293 5153 2307 5167
rect 2213 4993 2227 5007
rect 2013 4893 2027 4907
rect 2093 4773 2107 4787
rect 2473 5433 2487 5447
rect 2813 5533 2827 5547
rect 2773 5513 2787 5527
rect 2953 5473 2967 5487
rect 3013 5473 3027 5487
rect 2813 5453 2827 5467
rect 2613 5393 2627 5407
rect 2773 5413 2787 5427
rect 2753 5273 2767 5287
rect 2753 5193 2767 5207
rect 2593 5173 2607 5187
rect 2693 5173 2707 5187
rect 2393 5113 2407 5127
rect 2433 5113 2447 5127
rect 2373 5093 2387 5107
rect 2313 4993 2327 5007
rect 2213 4953 2227 4967
rect 2173 4753 2187 4767
rect 2113 4733 2127 4747
rect 1993 4713 2007 4727
rect 2093 4713 2107 4727
rect 2053 4693 2067 4707
rect 2033 4653 2047 4667
rect 2073 4653 2087 4667
rect 1933 4593 1947 4607
rect 1813 4353 1827 4367
rect 1893 4353 1907 4367
rect 1793 4293 1807 4307
rect 1773 4253 1787 4267
rect 1753 4233 1767 4247
rect 1773 4153 1787 4167
rect 1913 4293 1927 4307
rect 1833 4273 1847 4287
rect 1773 4113 1787 4127
rect 1813 4113 1827 4127
rect 1733 4033 1747 4047
rect 1733 4013 1747 4027
rect 2033 4513 2047 4527
rect 2093 4513 2107 4527
rect 1993 4493 2007 4507
rect 1973 4473 1987 4487
rect 2013 4473 2027 4487
rect 2053 4493 2067 4507
rect 2073 4473 2087 4487
rect 1953 4453 1967 4467
rect 2053 4453 2067 4467
rect 2053 4413 2067 4427
rect 1993 4253 2007 4267
rect 2093 4253 2107 4267
rect 2133 4693 2147 4707
rect 2293 4973 2307 4987
rect 2253 4953 2267 4967
rect 2333 4933 2347 4947
rect 2253 4713 2267 4727
rect 2153 4673 2167 4687
rect 2193 4673 2207 4687
rect 2233 4693 2247 4707
rect 2293 4673 2307 4687
rect 2133 4633 2147 4647
rect 2213 4633 2227 4647
rect 2273 4633 2287 4647
rect 2233 4613 2247 4627
rect 2173 4573 2187 4587
rect 2213 4553 2227 4567
rect 2153 4493 2167 4507
rect 2153 4453 2167 4467
rect 2193 4453 2207 4467
rect 2153 4373 2167 4387
rect 2333 4653 2347 4667
rect 2333 4613 2347 4627
rect 2353 4613 2367 4627
rect 2313 4573 2327 4587
rect 2313 4513 2327 4527
rect 2413 4933 2427 4947
rect 2453 5073 2467 5087
rect 2533 5033 2547 5047
rect 2453 4993 2467 5007
rect 2493 4973 2507 4987
rect 2473 4713 2487 4727
rect 2473 4693 2487 4707
rect 2713 5153 2727 5167
rect 2913 5413 2927 5427
rect 2833 5393 2847 5407
rect 2893 5393 2907 5407
rect 2973 5453 2987 5467
rect 3013 5413 3027 5427
rect 2993 5393 3007 5407
rect 2973 5373 2987 5387
rect 3073 5393 3087 5407
rect 3133 5513 3147 5527
rect 3313 5513 3327 5527
rect 3173 5453 3187 5467
rect 3233 5453 3247 5467
rect 3033 5353 3047 5367
rect 3093 5353 3107 5367
rect 3073 5333 3087 5347
rect 3073 5213 3087 5227
rect 2833 5193 2847 5207
rect 3013 5193 3027 5207
rect 2773 5153 2787 5167
rect 2733 5133 2747 5147
rect 2713 5033 2727 5047
rect 2733 5033 2747 5047
rect 2653 5013 2667 5027
rect 2673 5013 2687 5027
rect 2653 4973 2667 4987
rect 2613 4953 2627 4967
rect 2553 4913 2567 4927
rect 2533 4773 2547 4787
rect 2533 4693 2547 4707
rect 2433 4653 2447 4667
rect 2393 4633 2407 4647
rect 2453 4573 2467 4587
rect 2413 4553 2427 4567
rect 2373 4533 2387 4547
rect 2393 4493 2407 4507
rect 2433 4473 2447 4487
rect 2293 4453 2307 4467
rect 2293 4433 2307 4447
rect 2253 4373 2267 4387
rect 2173 4273 2187 4287
rect 1973 4233 1987 4247
rect 2033 4233 2047 4247
rect 2113 4233 2127 4247
rect 2213 4233 2227 4247
rect 1853 4213 1867 4227
rect 1913 4213 1927 4227
rect 1933 4213 1947 4227
rect 1953 4213 1967 4227
rect 1833 4033 1847 4047
rect 1573 3973 1587 3987
rect 1613 3973 1627 3987
rect 1513 3953 1527 3967
rect 1493 3933 1507 3947
rect 1353 3873 1367 3887
rect 1393 3873 1407 3887
rect 1333 3773 1347 3787
rect 1313 3753 1327 3767
rect 1293 3733 1307 3747
rect 1413 3773 1427 3787
rect 1393 3753 1407 3767
rect 1533 3913 1547 3927
rect 1513 3733 1527 3747
rect 1213 3693 1227 3707
rect 1133 3613 1147 3627
rect 1213 3653 1227 3667
rect 1153 3533 1167 3547
rect 1133 3493 1147 3507
rect 1113 3393 1127 3407
rect 1193 3373 1207 3387
rect 1013 3353 1027 3367
rect 1153 3353 1167 3367
rect 1173 3353 1187 3367
rect 813 3313 827 3327
rect 793 3293 807 3307
rect 793 3273 807 3287
rect 473 3233 487 3247
rect 653 3253 667 3267
rect 633 3233 647 3247
rect 673 3233 687 3247
rect 733 3233 747 3247
rect 433 3213 447 3227
rect 613 3213 627 3227
rect 413 3193 427 3207
rect 473 3193 487 3207
rect 493 3193 507 3207
rect 333 3173 347 3187
rect 353 3173 367 3187
rect 433 3153 447 3167
rect 393 3053 407 3067
rect 233 3033 247 3047
rect 253 3033 267 3047
rect 293 3033 307 3047
rect 373 3033 387 3047
rect 833 3293 847 3307
rect 853 3293 867 3307
rect 673 3193 687 3207
rect 593 3133 607 3147
rect 633 3133 647 3147
rect 753 3213 767 3227
rect 813 3213 827 3227
rect 713 3133 727 3147
rect 593 3053 607 3067
rect 613 3053 627 3067
rect 733 3053 747 3067
rect 433 3033 447 3047
rect 473 3033 487 3047
rect 573 3033 587 3047
rect 413 3013 427 3027
rect 533 3013 547 3027
rect 213 2993 227 3007
rect 273 2993 287 3007
rect 333 2993 347 3007
rect 133 2973 147 2987
rect 153 2973 167 2987
rect 113 2933 127 2947
rect 213 2833 227 2847
rect 153 2753 167 2767
rect 333 2813 347 2827
rect 233 2753 247 2767
rect 93 2733 107 2747
rect 133 2733 147 2747
rect 173 2733 187 2747
rect 73 2613 87 2627
rect 173 2713 187 2727
rect 113 2593 127 2607
rect 133 2593 147 2607
rect 73 2573 87 2587
rect 13 2373 27 2387
rect 93 2493 107 2507
rect 133 2573 147 2587
rect 313 2773 327 2787
rect 433 2913 447 2927
rect 413 2793 427 2807
rect 393 2773 407 2787
rect 293 2753 307 2767
rect 333 2753 347 2767
rect 393 2753 407 2767
rect 353 2733 367 2747
rect 373 2733 387 2747
rect 253 2713 267 2727
rect 413 2713 427 2727
rect 233 2693 247 2707
rect 413 2673 427 2687
rect 253 2613 267 2627
rect 453 2793 467 2807
rect 493 2773 507 2787
rect 553 2773 567 2787
rect 473 2733 487 2747
rect 293 2553 307 2567
rect 353 2553 367 2567
rect 393 2553 407 2567
rect 433 2553 447 2567
rect 233 2513 247 2527
rect 433 2533 447 2547
rect 513 2633 527 2647
rect 553 2733 567 2747
rect 553 2573 567 2587
rect 513 2553 527 2567
rect 433 2493 447 2507
rect 413 2453 427 2467
rect 333 2353 347 2367
rect 213 2313 227 2327
rect 253 2313 267 2327
rect 173 2293 187 2307
rect 233 2293 247 2307
rect 93 2253 107 2267
rect 113 2233 127 2247
rect 73 2193 87 2207
rect 93 2113 107 2127
rect 153 2273 167 2287
rect 193 2253 207 2267
rect 233 2253 247 2267
rect 153 2233 167 2247
rect 273 2253 287 2267
rect 233 2233 247 2247
rect 253 2233 267 2247
rect 193 2213 207 2227
rect 193 2093 207 2107
rect 213 2093 227 2107
rect 13 2033 27 2047
rect 53 2033 67 2047
rect 13 1913 27 1927
rect 33 1893 47 1907
rect 113 2053 127 2067
rect 73 1933 87 1947
rect 93 1893 107 1907
rect 53 1753 67 1767
rect 213 2033 227 2047
rect 253 2193 267 2207
rect 313 2233 327 2247
rect 293 2173 307 2187
rect 293 2133 307 2147
rect 273 2093 287 2107
rect 293 2073 307 2087
rect 293 2053 307 2067
rect 273 2033 287 2047
rect 253 1993 267 2007
rect 313 1973 327 1987
rect 233 1953 247 1967
rect 393 2293 407 2307
rect 353 2273 367 2287
rect 473 2513 487 2527
rect 453 2473 467 2487
rect 453 2293 467 2307
rect 373 2213 387 2227
rect 433 2253 447 2267
rect 413 2153 427 2167
rect 453 2173 467 2187
rect 433 2133 447 2147
rect 653 3013 667 3027
rect 633 2993 647 3007
rect 593 2933 607 2947
rect 653 2933 667 2947
rect 693 3013 707 3027
rect 713 2993 727 3007
rect 673 2833 687 2847
rect 653 2813 667 2827
rect 613 2733 627 2747
rect 673 2793 687 2807
rect 693 2793 707 2807
rect 713 2733 727 2747
rect 733 2653 747 2667
rect 833 3013 847 3027
rect 793 2913 807 2927
rect 893 3253 907 3267
rect 873 3233 887 3247
rect 973 3233 987 3247
rect 1273 3693 1287 3707
rect 1373 3713 1387 3727
rect 1413 3713 1427 3727
rect 1473 3693 1487 3707
rect 1313 3673 1327 3687
rect 1513 3653 1527 3667
rect 1253 3633 1267 3647
rect 1333 3573 1347 3587
rect 1273 3533 1287 3547
rect 1293 3533 1307 3547
rect 1233 3513 1247 3527
rect 1233 3473 1247 3487
rect 1273 3353 1287 3367
rect 1213 3313 1227 3327
rect 853 2993 867 3007
rect 853 2813 867 2827
rect 793 2773 807 2787
rect 833 2773 847 2787
rect 693 2633 707 2647
rect 753 2633 767 2647
rect 653 2613 667 2627
rect 653 2573 667 2587
rect 593 2553 607 2567
rect 613 2553 627 2567
rect 573 2493 587 2507
rect 633 2493 647 2507
rect 493 2273 507 2287
rect 513 2233 527 2247
rect 533 2233 547 2247
rect 573 2253 587 2267
rect 453 2113 467 2127
rect 473 2113 487 2127
rect 373 2093 387 2107
rect 493 2093 507 2107
rect 593 2213 607 2227
rect 613 2193 627 2207
rect 533 2113 547 2127
rect 593 2113 607 2127
rect 353 2053 367 2067
rect 393 2053 407 2067
rect 393 2033 407 2047
rect 333 1913 347 1927
rect 173 1793 187 1807
rect 353 1793 367 1807
rect 173 1773 187 1787
rect 173 1693 187 1707
rect 173 1673 187 1687
rect 113 1653 127 1667
rect 93 1633 107 1647
rect 13 1473 27 1487
rect 13 1333 27 1347
rect 73 1573 87 1587
rect 53 1553 67 1567
rect 133 1593 147 1607
rect 333 1713 347 1727
rect 233 1693 247 1707
rect 193 1653 207 1667
rect 213 1653 227 1667
rect 193 1633 207 1647
rect 153 1573 167 1587
rect 113 1533 127 1547
rect 53 1333 67 1347
rect 73 1333 87 1347
rect 53 1113 67 1127
rect 113 1113 127 1127
rect 73 1093 87 1107
rect 73 833 87 847
rect 53 653 67 667
rect 213 1393 227 1407
rect 293 1653 307 1667
rect 253 1613 267 1627
rect 253 1593 267 1607
rect 333 1633 347 1647
rect 293 1553 307 1567
rect 153 1373 167 1387
rect 173 1373 187 1387
rect 233 1373 247 1387
rect 273 1373 287 1387
rect 213 1333 227 1347
rect 373 1593 387 1607
rect 413 1993 427 2007
rect 413 1833 427 1847
rect 513 2073 527 2087
rect 513 2053 527 2067
rect 493 1973 507 1987
rect 453 1953 467 1967
rect 473 1953 487 1967
rect 473 1933 487 1947
rect 453 1793 467 1807
rect 433 1733 447 1747
rect 413 1693 427 1707
rect 453 1693 467 1707
rect 433 1593 447 1607
rect 353 1553 367 1567
rect 393 1553 407 1567
rect 333 1453 347 1467
rect 313 1373 327 1387
rect 273 1333 287 1347
rect 293 1333 307 1347
rect 333 1353 347 1367
rect 353 1333 367 1347
rect 173 1313 187 1327
rect 153 1293 167 1307
rect 193 1253 207 1267
rect 173 1213 187 1227
rect 153 1133 167 1147
rect 213 1153 227 1167
rect 373 1313 387 1327
rect 373 1293 387 1307
rect 313 1173 327 1187
rect 193 1093 207 1107
rect 213 1093 227 1107
rect 133 1053 147 1067
rect 273 1133 287 1147
rect 293 1133 307 1147
rect 333 1133 347 1147
rect 253 1093 267 1107
rect 273 1093 287 1107
rect 293 1013 307 1027
rect 273 993 287 1007
rect 233 953 247 967
rect 353 973 367 987
rect 333 933 347 947
rect 193 873 207 887
rect 433 1553 447 1567
rect 413 1493 427 1507
rect 553 1913 567 1927
rect 533 1873 547 1887
rect 673 2273 687 2287
rect 753 2613 767 2627
rect 733 2573 747 2587
rect 713 2553 727 2567
rect 773 2553 787 2567
rect 653 2173 667 2187
rect 693 2173 707 2187
rect 893 3153 907 3167
rect 1253 3233 1267 3247
rect 1173 3193 1187 3207
rect 993 3173 1007 3187
rect 1133 3073 1147 3087
rect 973 2993 987 3007
rect 913 2953 927 2967
rect 1473 3553 1487 3567
rect 1433 3533 1447 3547
rect 1313 3473 1327 3487
rect 1413 3473 1427 3487
rect 1513 3533 1527 3547
rect 1633 3893 1647 3907
rect 1593 3813 1607 3827
rect 1613 3713 1627 3727
rect 1733 3993 1747 4007
rect 1773 3993 1787 4007
rect 1873 4193 1887 4207
rect 1893 4173 1907 4187
rect 1993 4213 2007 4227
rect 1973 4173 1987 4187
rect 2013 4153 2027 4167
rect 1873 4133 1887 4147
rect 1933 4073 1947 4087
rect 2053 4213 2067 4227
rect 2073 4193 2087 4207
rect 2133 4173 2147 4187
rect 2073 4153 2087 4167
rect 1673 3973 1687 3987
rect 1713 3853 1727 3867
rect 1713 3833 1727 3847
rect 1673 3793 1687 3807
rect 1653 3693 1667 3707
rect 1573 3673 1587 3687
rect 1573 3633 1587 3647
rect 1593 3633 1607 3647
rect 1693 3713 1707 3727
rect 1833 3973 1847 3987
rect 1873 3973 1887 3987
rect 2033 4053 2047 4067
rect 1973 4013 1987 4027
rect 1953 3993 1967 4007
rect 1933 3973 1947 3987
rect 1973 3973 1987 3987
rect 1913 3893 1927 3907
rect 1793 3853 1807 3867
rect 1773 3813 1787 3827
rect 2053 3993 2067 4007
rect 2493 4493 2507 4507
rect 2473 4453 2487 4467
rect 2333 4393 2347 4407
rect 2313 4353 2327 4367
rect 2293 4233 2307 4247
rect 2253 4193 2267 4207
rect 2173 4113 2187 4127
rect 2293 4153 2307 4167
rect 2273 4093 2287 4107
rect 2413 4313 2427 4327
rect 2333 4213 2347 4227
rect 2393 4193 2407 4207
rect 2393 4173 2407 4187
rect 2353 4133 2367 4147
rect 2233 4053 2247 4067
rect 2293 4053 2307 4067
rect 2313 4053 2327 4067
rect 2113 4033 2127 4047
rect 2133 4033 2147 4047
rect 2033 3953 2047 3967
rect 2013 3893 2027 3907
rect 2093 3953 2107 3967
rect 2073 3853 2087 3867
rect 2053 3813 2067 3827
rect 1773 3753 1787 3767
rect 1973 3753 1987 3767
rect 1993 3733 2007 3747
rect 1773 3713 1787 3727
rect 1753 3693 1767 3707
rect 1793 3693 1807 3707
rect 1693 3673 1707 3687
rect 1733 3673 1747 3687
rect 1813 3653 1827 3667
rect 1693 3613 1707 3627
rect 1773 3613 1787 3627
rect 1713 3593 1727 3607
rect 1673 3573 1687 3587
rect 1593 3553 1607 3567
rect 1633 3533 1647 3547
rect 1493 3473 1507 3487
rect 1613 3493 1627 3507
rect 1653 3513 1667 3527
rect 1733 3533 1747 3547
rect 1913 3713 1927 3727
rect 1853 3693 1867 3707
rect 1873 3573 1887 3587
rect 1873 3553 1887 3567
rect 1773 3533 1787 3547
rect 1813 3533 1827 3547
rect 1833 3533 1847 3547
rect 1413 3333 1427 3347
rect 1293 3213 1307 3227
rect 1293 3193 1307 3207
rect 1313 3153 1327 3167
rect 1353 3213 1367 3227
rect 1393 3213 1407 3227
rect 1413 3153 1427 3167
rect 1273 2973 1287 2987
rect 1213 2913 1227 2927
rect 1233 2913 1247 2927
rect 1173 2893 1187 2907
rect 893 2813 907 2827
rect 913 2813 927 2827
rect 873 2773 887 2787
rect 913 2793 927 2807
rect 813 2733 827 2747
rect 833 2713 847 2727
rect 893 2733 907 2747
rect 993 2753 1007 2767
rect 1013 2753 1027 2767
rect 933 2733 947 2747
rect 973 2713 987 2727
rect 813 2673 827 2687
rect 873 2673 887 2687
rect 793 2533 807 2547
rect 953 2653 967 2667
rect 853 2573 867 2587
rect 833 2553 847 2567
rect 793 2473 807 2487
rect 813 2473 827 2487
rect 813 2413 827 2427
rect 853 2333 867 2347
rect 773 2273 787 2287
rect 793 2273 807 2287
rect 753 2233 767 2247
rect 773 2133 787 2147
rect 713 2113 727 2127
rect 653 2093 667 2107
rect 733 2093 747 2107
rect 593 1833 607 1847
rect 633 1833 647 1847
rect 513 1813 527 1827
rect 553 1813 567 1827
rect 533 1773 547 1787
rect 513 1693 527 1707
rect 473 1573 487 1587
rect 493 1573 507 1587
rect 513 1573 527 1587
rect 573 1793 587 1807
rect 553 1753 567 1767
rect 573 1713 587 1727
rect 573 1593 587 1607
rect 513 1553 527 1567
rect 453 1533 467 1547
rect 473 1513 487 1527
rect 513 1513 527 1527
rect 433 1473 447 1487
rect 413 1453 427 1467
rect 433 1453 447 1467
rect 393 1233 407 1247
rect 473 1393 487 1407
rect 493 1393 507 1407
rect 473 1353 487 1367
rect 493 1333 507 1347
rect 533 1373 547 1387
rect 613 1793 627 1807
rect 613 1653 627 1667
rect 693 2073 707 2087
rect 933 2473 947 2487
rect 953 2453 967 2467
rect 873 2313 887 2327
rect 853 2273 867 2287
rect 893 2293 907 2307
rect 873 2253 887 2267
rect 913 2253 927 2267
rect 793 2093 807 2107
rect 833 2093 847 2107
rect 733 2053 747 2067
rect 793 2053 807 2067
rect 693 2033 707 2047
rect 753 2033 767 2047
rect 673 1873 687 1887
rect 673 1753 687 1767
rect 753 1873 767 1887
rect 753 1833 767 1847
rect 913 2073 927 2087
rect 853 2053 867 2067
rect 1153 2773 1167 2787
rect 1133 2753 1147 2767
rect 1013 2713 1027 2727
rect 1093 2733 1107 2747
rect 1113 2733 1127 2747
rect 1153 2733 1167 2747
rect 1033 2693 1047 2707
rect 1093 2613 1107 2627
rect 1113 2613 1127 2627
rect 1053 2553 1067 2567
rect 1033 2493 1047 2507
rect 1093 2533 1107 2547
rect 1013 2473 1027 2487
rect 1093 2453 1107 2467
rect 1193 2773 1207 2787
rect 1213 2773 1227 2787
rect 1173 2653 1187 2667
rect 1153 2473 1167 2487
rect 1173 2473 1187 2487
rect 993 2313 1007 2327
rect 1053 2313 1067 2327
rect 1073 2313 1087 2327
rect 1113 2313 1127 2327
rect 993 2293 1007 2307
rect 1033 2293 1047 2307
rect 973 2133 987 2147
rect 953 2053 967 2067
rect 833 1993 847 2007
rect 813 1873 827 1887
rect 793 1813 807 1827
rect 753 1793 767 1807
rect 813 1793 827 1807
rect 873 2033 887 2047
rect 1033 2233 1047 2247
rect 1073 2293 1087 2307
rect 1093 2273 1107 2287
rect 1073 2253 1087 2267
rect 1093 2253 1107 2267
rect 1053 2113 1067 2127
rect 1013 2073 1027 2087
rect 1113 2233 1127 2247
rect 1093 2213 1107 2227
rect 1333 3013 1347 3027
rect 1393 3013 1407 3027
rect 1313 2973 1327 2987
rect 1253 2673 1267 2687
rect 1233 2613 1247 2627
rect 1473 3213 1487 3227
rect 1693 3453 1707 3467
rect 1593 3393 1607 3407
rect 1633 3353 1647 3367
rect 1673 3353 1687 3367
rect 1533 3253 1547 3267
rect 1593 3253 1607 3267
rect 1453 3193 1467 3207
rect 1493 3193 1507 3207
rect 1553 3193 1567 3207
rect 1573 3173 1587 3187
rect 1613 3173 1627 3187
rect 1533 3153 1547 3167
rect 1573 3153 1587 3167
rect 1473 3133 1487 3147
rect 1453 3093 1467 3107
rect 1433 2893 1447 2907
rect 1553 3113 1567 3127
rect 1513 3073 1527 3087
rect 1493 3053 1507 3067
rect 1473 2913 1487 2927
rect 1453 2853 1467 2867
rect 1333 2773 1347 2787
rect 1753 3313 1767 3327
rect 1733 3253 1747 3267
rect 1713 3233 1727 3247
rect 1653 3213 1667 3227
rect 1693 3193 1707 3207
rect 1653 3093 1667 3107
rect 1593 3073 1607 3087
rect 1633 3073 1647 3087
rect 1633 3053 1647 3067
rect 1753 3213 1767 3227
rect 1753 3193 1767 3207
rect 1733 3173 1747 3187
rect 1753 3133 1767 3147
rect 1833 3513 1847 3527
rect 2073 3733 2087 3747
rect 2093 3733 2107 3747
rect 2273 4013 2287 4027
rect 2313 4033 2327 4047
rect 2313 4013 2327 4027
rect 2153 3973 2167 3987
rect 2293 3993 2307 4007
rect 2253 3973 2267 3987
rect 2213 3853 2227 3867
rect 2353 3993 2367 4007
rect 2373 3953 2387 3967
rect 2253 3833 2267 3847
rect 2273 3833 2287 3847
rect 2253 3813 2267 3827
rect 2113 3713 2127 3727
rect 2053 3693 2067 3707
rect 2093 3693 2107 3707
rect 2213 3713 2227 3727
rect 2013 3673 2027 3687
rect 2053 3673 2067 3687
rect 1993 3593 2007 3607
rect 1913 3493 1927 3507
rect 1953 3513 1967 3527
rect 1973 3513 1987 3527
rect 2033 3573 2047 3587
rect 2013 3493 2027 3507
rect 1793 3213 1807 3227
rect 1833 3213 1847 3227
rect 1813 3193 1827 3207
rect 1833 3153 1847 3167
rect 1773 3093 1787 3107
rect 1753 3073 1767 3087
rect 1613 3033 1627 3047
rect 1713 3053 1727 3067
rect 1773 3053 1787 3067
rect 1793 3053 1807 3067
rect 1693 3033 1707 3047
rect 1613 3013 1627 3027
rect 1593 2993 1607 3007
rect 1653 2993 1667 3007
rect 1653 2913 1667 2927
rect 1673 2893 1687 2907
rect 1533 2873 1547 2887
rect 1573 2873 1587 2887
rect 1653 2853 1667 2867
rect 1633 2793 1647 2807
rect 1473 2753 1487 2767
rect 1593 2753 1607 2767
rect 1653 2733 1667 2747
rect 1473 2713 1487 2727
rect 1633 2673 1647 2687
rect 1333 2653 1347 2667
rect 1373 2653 1387 2667
rect 1433 2653 1447 2667
rect 1313 2613 1327 2627
rect 1293 2593 1307 2607
rect 1313 2593 1327 2607
rect 1353 2593 1367 2607
rect 1293 2573 1307 2587
rect 1273 2513 1287 2527
rect 1233 2493 1247 2507
rect 1253 2473 1267 2487
rect 1193 2273 1207 2287
rect 1233 2273 1247 2287
rect 1193 2233 1207 2247
rect 1173 2213 1187 2227
rect 1113 2113 1127 2127
rect 1153 2113 1167 2127
rect 1093 2093 1107 2107
rect 1053 2053 1067 2067
rect 1073 2053 1087 2067
rect 1033 2033 1047 2047
rect 933 2013 947 2027
rect 973 2013 987 2027
rect 993 2013 1007 2027
rect 893 1993 907 2007
rect 1093 2013 1107 2027
rect 1073 1973 1087 1987
rect 933 1953 947 1967
rect 1093 1953 1107 1967
rect 873 1833 887 1847
rect 693 1713 707 1727
rect 653 1693 667 1707
rect 673 1693 687 1707
rect 633 1633 647 1647
rect 693 1673 707 1687
rect 593 1473 607 1487
rect 633 1573 647 1587
rect 613 1453 627 1467
rect 633 1433 647 1447
rect 573 1413 587 1427
rect 633 1413 647 1427
rect 553 1353 567 1367
rect 593 1353 607 1367
rect 513 1293 527 1307
rect 453 1273 467 1287
rect 493 1273 507 1287
rect 473 1233 487 1247
rect 433 1213 447 1227
rect 413 1133 427 1147
rect 453 1133 467 1147
rect 453 1093 467 1107
rect 433 1073 447 1087
rect 413 1053 427 1067
rect 453 1053 467 1067
rect 393 1033 407 1047
rect 393 973 407 987
rect 333 853 347 867
rect 93 633 107 647
rect 133 633 147 647
rect 93 613 107 627
rect 133 613 147 627
rect 313 733 327 747
rect 213 633 227 647
rect 273 633 287 647
rect 153 593 167 607
rect 253 593 267 607
rect 73 553 87 567
rect 293 533 307 547
rect 353 773 367 787
rect 413 793 427 807
rect 393 773 407 787
rect 373 733 387 747
rect 353 713 367 727
rect 333 593 347 607
rect 453 853 467 867
rect 553 1293 567 1307
rect 533 1253 547 1267
rect 773 1773 787 1787
rect 773 1753 787 1767
rect 753 1713 767 1727
rect 753 1653 767 1667
rect 713 1633 727 1647
rect 733 1633 747 1647
rect 713 1593 727 1607
rect 813 1753 827 1767
rect 853 1773 867 1787
rect 893 1813 907 1827
rect 833 1713 847 1727
rect 873 1713 887 1727
rect 1033 1813 1047 1827
rect 1073 1813 1087 1827
rect 953 1793 967 1807
rect 973 1793 987 1807
rect 993 1773 1007 1787
rect 933 1753 947 1767
rect 953 1753 967 1767
rect 913 1713 927 1727
rect 793 1693 807 1707
rect 893 1693 907 1707
rect 813 1673 827 1687
rect 893 1673 907 1687
rect 793 1633 807 1647
rect 693 1553 707 1567
rect 693 1513 707 1527
rect 653 1373 667 1387
rect 653 1353 667 1367
rect 693 1313 707 1327
rect 613 1253 627 1267
rect 633 1253 647 1267
rect 613 1233 627 1247
rect 793 1533 807 1547
rect 733 1313 747 1327
rect 713 1273 727 1287
rect 793 1333 807 1347
rect 773 1293 787 1307
rect 733 1253 747 1267
rect 753 1253 767 1267
rect 793 1253 807 1267
rect 633 1213 647 1227
rect 673 1213 687 1227
rect 573 1193 587 1207
rect 493 1133 507 1147
rect 533 1133 547 1147
rect 493 1113 507 1127
rect 513 1093 527 1107
rect 553 1093 567 1107
rect 493 1073 507 1087
rect 533 1073 547 1087
rect 513 1053 527 1067
rect 493 1013 507 1027
rect 533 1033 547 1047
rect 553 1033 567 1047
rect 493 933 507 947
rect 493 853 507 867
rect 513 833 527 847
rect 473 813 487 827
rect 493 793 507 807
rect 453 733 467 747
rect 393 653 407 667
rect 433 653 447 667
rect 393 633 407 647
rect 413 613 427 627
rect 453 633 467 647
rect 613 1153 627 1167
rect 713 1153 727 1167
rect 593 1133 607 1147
rect 593 1073 607 1087
rect 653 1133 667 1147
rect 653 1093 667 1107
rect 693 1093 707 1107
rect 753 1213 767 1227
rect 733 1093 747 1107
rect 673 1073 687 1087
rect 733 1073 747 1087
rect 693 1053 707 1067
rect 713 1053 727 1067
rect 753 1053 767 1067
rect 593 1013 607 1027
rect 653 993 667 1007
rect 593 953 607 967
rect 553 873 567 887
rect 573 873 587 887
rect 633 833 647 847
rect 553 793 567 807
rect 573 793 587 807
rect 613 793 627 807
rect 533 693 547 707
rect 533 673 547 687
rect 513 633 527 647
rect 633 693 647 707
rect 573 673 587 687
rect 533 613 547 627
rect 473 553 487 567
rect 353 533 367 547
rect 313 493 327 507
rect 73 353 87 367
rect 193 313 207 327
rect 193 173 207 187
rect 73 133 87 147
rect 393 493 407 507
rect 473 393 487 407
rect 453 373 467 387
rect 573 393 587 407
rect 493 353 507 367
rect 513 353 527 367
rect 573 353 587 367
rect 533 333 547 347
rect 553 313 567 327
rect 593 313 607 327
rect 613 233 627 247
rect 573 213 587 227
rect 453 113 467 127
rect 733 973 747 987
rect 713 893 727 907
rect 693 833 707 847
rect 673 813 687 827
rect 713 813 727 827
rect 773 973 787 987
rect 893 1633 907 1647
rect 933 1633 947 1647
rect 833 1573 847 1587
rect 913 1573 927 1587
rect 833 1553 847 1567
rect 873 1553 887 1567
rect 833 1493 847 1507
rect 813 1213 827 1227
rect 933 1493 947 1507
rect 853 1353 867 1367
rect 913 1353 927 1367
rect 893 1333 907 1347
rect 933 1333 947 1347
rect 873 1313 887 1327
rect 1353 2513 1367 2527
rect 1313 2413 1327 2427
rect 1353 2413 1367 2427
rect 1313 2373 1327 2387
rect 1333 2253 1347 2267
rect 1273 2233 1287 2247
rect 1273 2193 1287 2207
rect 1213 2153 1227 2167
rect 1193 2093 1207 2107
rect 1173 2053 1187 2067
rect 1153 1993 1167 2007
rect 1133 1913 1147 1927
rect 1113 1853 1127 1867
rect 1113 1833 1127 1847
rect 1053 1773 1067 1787
rect 1093 1773 1107 1787
rect 1013 1733 1027 1747
rect 1033 1733 1047 1747
rect 1013 1673 1027 1687
rect 993 1633 1007 1647
rect 973 1613 987 1627
rect 1033 1633 1047 1647
rect 993 1573 1007 1587
rect 993 1473 1007 1487
rect 1133 1713 1147 1727
rect 1113 1673 1127 1687
rect 1073 1653 1087 1667
rect 1093 1653 1107 1667
rect 1133 1633 1147 1647
rect 1093 1613 1107 1627
rect 1113 1613 1127 1627
rect 1073 1553 1087 1567
rect 1053 1533 1067 1547
rect 1013 1313 1027 1327
rect 1173 1953 1187 1967
rect 1253 2013 1267 2027
rect 1353 2193 1367 2207
rect 1293 2133 1307 2147
rect 1293 2113 1307 2127
rect 1273 1993 1287 2007
rect 1213 1933 1227 1947
rect 1413 2553 1427 2567
rect 1393 2513 1407 2527
rect 1513 2593 1527 2607
rect 1553 2593 1567 2607
rect 1593 2593 1607 2607
rect 1473 2533 1487 2547
rect 1473 2393 1487 2407
rect 1393 2333 1407 2347
rect 1413 2253 1427 2267
rect 1393 2233 1407 2247
rect 1433 2233 1447 2247
rect 1533 2533 1547 2547
rect 1573 2533 1587 2547
rect 1593 2513 1607 2527
rect 1513 2393 1527 2407
rect 1533 2273 1547 2287
rect 1493 2253 1507 2267
rect 1473 2233 1487 2247
rect 1553 2233 1567 2247
rect 1453 2213 1467 2227
rect 1513 2213 1527 2227
rect 1713 2953 1727 2967
rect 1713 2913 1727 2927
rect 1693 2813 1707 2827
rect 1753 2753 1767 2767
rect 1773 2753 1787 2767
rect 1693 2733 1707 2747
rect 1753 2713 1767 2727
rect 1753 2693 1767 2707
rect 1733 2673 1747 2687
rect 1673 2613 1687 2627
rect 1713 2553 1727 2567
rect 1693 2513 1707 2527
rect 1633 2453 1647 2467
rect 1733 2453 1747 2467
rect 1593 2233 1607 2247
rect 1673 2273 1687 2287
rect 1713 2273 1727 2287
rect 1613 2193 1627 2207
rect 1693 2233 1707 2247
rect 1653 2173 1667 2187
rect 1713 2173 1727 2187
rect 1493 2133 1507 2147
rect 1773 2673 1787 2687
rect 1773 2633 1787 2647
rect 1833 3093 1847 3107
rect 1813 2953 1827 2967
rect 1893 3453 1907 3467
rect 2013 3453 2027 3467
rect 1873 3193 1887 3207
rect 1853 3073 1867 3087
rect 1873 3073 1887 3087
rect 1853 2993 1867 3007
rect 1833 2793 1847 2807
rect 1873 2873 1887 2887
rect 1853 2773 1867 2787
rect 1833 2753 1847 2767
rect 2193 3673 2207 3687
rect 2193 3613 2207 3627
rect 2113 3573 2127 3587
rect 2173 3573 2187 3587
rect 2193 3573 2207 3587
rect 2213 3553 2227 3567
rect 1973 3433 1987 3447
rect 2033 3433 2047 3447
rect 1933 3273 1947 3287
rect 1933 3233 1947 3247
rect 1933 3193 1947 3207
rect 1953 3193 1967 3207
rect 1913 3153 1927 3167
rect 2153 3513 2167 3527
rect 2173 3513 2187 3527
rect 2133 3473 2147 3487
rect 2193 3473 2207 3487
rect 2353 3733 2367 3747
rect 2293 3693 2307 3707
rect 2353 3693 2367 3707
rect 2373 3693 2387 3707
rect 2313 3673 2327 3687
rect 2373 3633 2387 3647
rect 2493 4333 2507 4347
rect 2653 4913 2667 4927
rect 2873 5133 2887 5147
rect 2893 5073 2907 5087
rect 2813 5033 2827 5047
rect 2793 5013 2807 5027
rect 2773 4933 2787 4947
rect 2813 4913 2827 4927
rect 2633 4873 2647 4887
rect 2613 4693 2627 4707
rect 2553 4653 2567 4667
rect 2553 4633 2567 4647
rect 2573 4633 2587 4647
rect 2553 4493 2567 4507
rect 2613 4673 2627 4687
rect 2633 4673 2647 4687
rect 2593 4613 2607 4627
rect 3013 5173 3027 5187
rect 2993 5113 3007 5127
rect 3053 5133 3067 5147
rect 3093 5133 3107 5147
rect 3053 5113 3067 5127
rect 2933 4993 2947 5007
rect 3013 4993 3027 5007
rect 2893 4933 2907 4947
rect 2953 4953 2967 4967
rect 2893 4733 2907 4747
rect 2793 4693 2807 4707
rect 2853 4693 2867 4707
rect 2673 4673 2687 4687
rect 2733 4673 2747 4687
rect 2773 4673 2787 4687
rect 2853 4673 2867 4687
rect 2593 4513 2607 4527
rect 2613 4513 2627 4527
rect 2573 4473 2587 4487
rect 2593 4473 2607 4487
rect 2553 4453 2567 4467
rect 2593 4453 2607 4467
rect 2613 4353 2627 4367
rect 2533 4313 2547 4327
rect 2533 4293 2547 4307
rect 2513 4273 2527 4287
rect 2513 4233 2527 4247
rect 2453 4213 2467 4227
rect 2433 4173 2447 4187
rect 2613 4273 2627 4287
rect 2493 4173 2507 4187
rect 2533 4173 2547 4187
rect 2593 4173 2607 4187
rect 2433 4153 2447 4167
rect 2453 4153 2467 4167
rect 2513 4153 2527 4167
rect 2553 4153 2567 4167
rect 2413 4133 2427 4147
rect 2413 4053 2427 4067
rect 2453 4093 2467 4107
rect 2433 4033 2447 4047
rect 2473 4013 2487 4027
rect 2493 3993 2507 4007
rect 2533 4133 2547 4147
rect 2573 4053 2587 4067
rect 2513 3973 2527 3987
rect 2553 3973 2567 3987
rect 2593 4013 2607 4027
rect 2473 3793 2487 3807
rect 2433 3773 2447 3787
rect 2473 3733 2487 3747
rect 2513 3733 2527 3747
rect 2573 3733 2587 3747
rect 2433 3713 2447 3727
rect 2493 3713 2507 3727
rect 2513 3713 2527 3727
rect 2493 3693 2507 3707
rect 2453 3673 2467 3687
rect 2293 3613 2307 3627
rect 2393 3613 2407 3627
rect 2113 3453 2127 3467
rect 2153 3453 2167 3467
rect 2033 3333 2047 3347
rect 1953 3133 1967 3147
rect 1973 3133 1987 3147
rect 1933 3053 1947 3067
rect 1913 3033 1927 3047
rect 1993 3053 2007 3067
rect 1973 3013 1987 3027
rect 2053 3173 2067 3187
rect 2073 3153 2087 3167
rect 2033 3133 2047 3147
rect 1953 2993 1967 3007
rect 2013 2993 2027 3007
rect 1993 2973 2007 2987
rect 2053 3053 2067 3067
rect 2213 3413 2227 3427
rect 2133 3253 2147 3267
rect 2173 3233 2187 3247
rect 2113 3213 2127 3227
rect 2153 3213 2167 3227
rect 2113 3193 2127 3207
rect 2133 3173 2147 3187
rect 2113 3133 2127 3147
rect 2113 3073 2127 3087
rect 2093 3013 2107 3027
rect 2173 3073 2187 3087
rect 2133 3033 2147 3047
rect 2153 3033 2167 3047
rect 2053 2993 2067 3007
rect 2133 2993 2147 3007
rect 2073 2973 2087 2987
rect 1953 2933 1967 2947
rect 2033 2933 2047 2947
rect 2053 2933 2067 2947
rect 1933 2913 1947 2927
rect 1893 2833 1907 2847
rect 1933 2753 1947 2767
rect 1853 2733 1867 2747
rect 1893 2733 1907 2747
rect 1913 2713 1927 2727
rect 1813 2693 1827 2707
rect 1833 2693 1847 2707
rect 1833 2653 1847 2667
rect 1893 2653 1907 2667
rect 1873 2613 1887 2627
rect 1793 2573 1807 2587
rect 1833 2553 1847 2567
rect 1773 2313 1787 2327
rect 1753 2233 1767 2247
rect 1373 2093 1387 2107
rect 1453 2093 1467 2107
rect 1473 2093 1487 2107
rect 1493 2093 1507 2107
rect 1313 2073 1327 2087
rect 1333 2073 1347 2087
rect 1373 2073 1387 2087
rect 1173 1913 1187 1927
rect 1293 1913 1307 1927
rect 1193 1873 1207 1887
rect 1173 1833 1187 1847
rect 1253 1853 1267 1867
rect 1213 1813 1227 1827
rect 1173 1733 1187 1747
rect 1233 1773 1247 1787
rect 1213 1673 1227 1687
rect 1353 2013 1367 2027
rect 1373 1993 1387 2007
rect 1353 1973 1367 1987
rect 1333 1873 1347 1887
rect 1313 1833 1327 1847
rect 1313 1793 1327 1807
rect 1313 1773 1327 1787
rect 1273 1753 1287 1767
rect 1173 1633 1187 1647
rect 1253 1633 1267 1647
rect 1333 1633 1347 1647
rect 1213 1613 1227 1627
rect 1293 1613 1307 1627
rect 1193 1573 1207 1587
rect 1313 1593 1327 1607
rect 1233 1573 1247 1587
rect 1213 1553 1227 1567
rect 1113 1333 1127 1347
rect 1153 1333 1167 1347
rect 1073 1313 1087 1327
rect 853 1273 867 1287
rect 953 1273 967 1287
rect 973 1273 987 1287
rect 1133 1313 1147 1327
rect 1093 1273 1107 1287
rect 893 1253 907 1267
rect 993 1253 1007 1267
rect 1113 1253 1127 1267
rect 853 1093 867 1107
rect 833 1073 847 1087
rect 993 1233 1007 1247
rect 913 1213 927 1227
rect 953 1133 967 1147
rect 973 1133 987 1147
rect 913 1093 927 1107
rect 933 1073 947 1087
rect 973 1073 987 1087
rect 973 1053 987 1067
rect 853 1033 867 1047
rect 893 1033 907 1047
rect 833 1013 847 1027
rect 813 993 827 1007
rect 793 953 807 967
rect 753 933 767 947
rect 793 873 807 887
rect 753 813 767 827
rect 773 813 787 827
rect 733 773 747 787
rect 713 633 727 647
rect 693 613 707 627
rect 733 613 747 627
rect 753 613 767 627
rect 713 593 727 607
rect 653 433 667 447
rect 653 413 667 427
rect 653 393 667 407
rect 693 393 707 407
rect 673 333 687 347
rect 733 433 747 447
rect 813 793 827 807
rect 873 953 887 967
rect 853 793 867 807
rect 833 673 847 687
rect 913 873 927 887
rect 893 813 907 827
rect 933 793 947 807
rect 953 773 967 787
rect 1093 1193 1107 1207
rect 1073 1153 1087 1167
rect 1033 1133 1047 1147
rect 1153 1213 1167 1227
rect 1193 1353 1207 1367
rect 1333 1513 1347 1527
rect 1293 1493 1307 1507
rect 1253 1353 1267 1367
rect 1273 1353 1287 1367
rect 1233 1333 1247 1347
rect 1193 1293 1207 1307
rect 1193 1173 1207 1187
rect 1173 1133 1187 1147
rect 1273 1293 1287 1307
rect 1333 1353 1347 1367
rect 1313 1273 1327 1287
rect 1293 1253 1307 1267
rect 1393 1973 1407 1987
rect 1433 1953 1447 1967
rect 1433 1813 1447 1827
rect 1593 2093 1607 2107
rect 1533 2053 1547 2067
rect 1493 2013 1507 2027
rect 1653 2053 1667 2067
rect 1673 2033 1687 2047
rect 1573 1953 1587 1967
rect 1553 1913 1567 1927
rect 1533 1873 1547 1887
rect 1553 1873 1567 1887
rect 1473 1833 1487 1847
rect 1413 1793 1427 1807
rect 1453 1793 1467 1807
rect 1473 1793 1487 1807
rect 1513 1793 1527 1807
rect 1473 1773 1487 1787
rect 1553 1773 1567 1787
rect 1653 1933 1667 1947
rect 1593 1793 1607 1807
rect 1433 1653 1447 1667
rect 1393 1613 1407 1627
rect 1433 1613 1447 1627
rect 1373 1593 1387 1607
rect 1373 1513 1387 1527
rect 1353 1233 1367 1247
rect 1273 1153 1287 1167
rect 1413 1553 1427 1567
rect 1413 1533 1427 1547
rect 1533 1753 1547 1767
rect 1573 1753 1587 1767
rect 1473 1713 1487 1727
rect 1593 1653 1607 1667
rect 1553 1633 1567 1647
rect 1513 1593 1527 1607
rect 1493 1553 1507 1567
rect 1533 1553 1547 1567
rect 1493 1513 1507 1527
rect 1473 1473 1487 1487
rect 1533 1393 1547 1407
rect 1453 1373 1467 1387
rect 1513 1353 1527 1367
rect 1413 1333 1427 1347
rect 1433 1333 1447 1347
rect 1473 1313 1487 1327
rect 1433 1273 1447 1287
rect 1393 1213 1407 1227
rect 1373 1133 1387 1147
rect 1193 1113 1207 1127
rect 1233 1113 1247 1127
rect 1113 1093 1127 1107
rect 1013 1073 1027 1087
rect 1053 1073 1067 1087
rect 1093 1073 1107 1087
rect 1013 993 1027 1007
rect 993 773 1007 787
rect 893 693 907 707
rect 973 693 987 707
rect 993 693 1007 707
rect 873 633 887 647
rect 913 613 927 627
rect 953 613 967 627
rect 893 553 907 567
rect 793 433 807 447
rect 833 433 847 447
rect 773 373 787 387
rect 873 373 887 387
rect 753 293 767 307
rect 713 273 727 287
rect 633 193 647 207
rect 773 193 787 207
rect 713 173 727 187
rect 613 153 627 167
rect 693 153 707 167
rect 753 153 767 167
rect 973 393 987 407
rect 1033 953 1047 967
rect 1113 873 1127 887
rect 1093 853 1107 867
rect 1033 833 1047 847
rect 1073 793 1087 807
rect 1113 833 1127 847
rect 1193 1073 1207 1087
rect 1233 1073 1247 1087
rect 1173 1053 1187 1067
rect 1293 1093 1307 1107
rect 1293 1073 1307 1087
rect 1273 1053 1287 1067
rect 1253 1033 1267 1047
rect 1193 1013 1207 1027
rect 1253 1013 1267 1027
rect 1173 873 1187 887
rect 1173 833 1187 847
rect 1133 813 1147 827
rect 1253 813 1267 827
rect 1113 773 1127 787
rect 1153 773 1167 787
rect 1093 753 1107 767
rect 1073 693 1087 707
rect 1013 673 1027 687
rect 993 373 1007 387
rect 1033 653 1047 667
rect 1093 673 1107 687
rect 1093 633 1107 647
rect 1053 613 1067 627
rect 1233 793 1247 807
rect 1353 1113 1367 1127
rect 1413 1193 1427 1207
rect 1373 1093 1387 1107
rect 1433 993 1447 1007
rect 1513 1293 1527 1307
rect 1493 1233 1507 1247
rect 1513 1173 1527 1187
rect 1473 1113 1487 1127
rect 1573 1593 1587 1607
rect 1613 1593 1627 1607
rect 1853 2333 1867 2347
rect 2033 2873 2047 2887
rect 1993 2833 2007 2847
rect 1973 2813 1987 2827
rect 2113 2933 2127 2947
rect 2033 2793 2047 2807
rect 2013 2773 2027 2787
rect 2033 2753 2047 2767
rect 1993 2693 2007 2707
rect 1973 2653 1987 2667
rect 2053 2713 2067 2727
rect 2033 2633 2047 2647
rect 2013 2613 2027 2627
rect 2413 3593 2427 3607
rect 2353 3553 2367 3567
rect 2393 3553 2407 3567
rect 2313 3513 2327 3527
rect 2433 3573 2447 3587
rect 2373 3473 2387 3487
rect 2293 3353 2307 3367
rect 2393 3253 2407 3267
rect 2253 3233 2267 3247
rect 2333 3233 2347 3247
rect 2373 3233 2387 3247
rect 2413 3233 2427 3247
rect 2273 3193 2287 3207
rect 2313 3193 2327 3207
rect 2233 3173 2247 3187
rect 2233 3153 2247 3167
rect 2173 2993 2187 3007
rect 2153 2873 2167 2887
rect 2173 2853 2187 2867
rect 2213 2993 2227 3007
rect 2253 2993 2267 3007
rect 2413 3133 2427 3147
rect 2373 3113 2387 3127
rect 2353 3053 2367 3067
rect 2313 3033 2327 3047
rect 2333 3033 2347 3047
rect 2293 2993 2307 3007
rect 2453 3553 2467 3567
rect 2473 3513 2487 3527
rect 2493 3473 2507 3487
rect 2453 3433 2467 3447
rect 2473 3233 2487 3247
rect 2453 3193 2467 3207
rect 2433 3073 2447 3087
rect 2393 3053 2407 3067
rect 2413 3053 2427 3067
rect 2373 2993 2387 3007
rect 2313 2933 2327 2947
rect 2273 2913 2287 2927
rect 2293 2913 2307 2927
rect 2273 2853 2287 2867
rect 2213 2793 2227 2807
rect 2193 2773 2207 2787
rect 2133 2733 2147 2747
rect 2253 2753 2267 2767
rect 2453 3033 2467 3047
rect 2473 3033 2487 3047
rect 2433 3013 2447 3027
rect 2433 2973 2447 2987
rect 2413 2893 2427 2907
rect 2393 2873 2407 2887
rect 2313 2813 2327 2827
rect 2393 2793 2407 2807
rect 2313 2753 2327 2767
rect 2373 2773 2387 2787
rect 2153 2713 2167 2727
rect 2273 2733 2287 2747
rect 2293 2733 2307 2747
rect 2333 2733 2347 2747
rect 2273 2713 2287 2727
rect 2133 2693 2147 2707
rect 2193 2693 2207 2707
rect 2113 2593 2127 2607
rect 2073 2573 2087 2587
rect 1973 2553 1987 2567
rect 2013 2553 2027 2567
rect 2093 2533 2107 2547
rect 2173 2613 2187 2627
rect 2173 2553 2187 2567
rect 2253 2593 2267 2607
rect 2353 2653 2367 2667
rect 2193 2533 2207 2547
rect 2153 2513 2167 2527
rect 1993 2473 2007 2487
rect 2173 2453 2187 2467
rect 2173 2433 2187 2447
rect 1893 2313 1907 2327
rect 1873 2293 1887 2307
rect 2053 2293 2067 2307
rect 2093 2293 2107 2307
rect 2153 2293 2167 2307
rect 1813 2273 1827 2287
rect 1893 2273 1907 2287
rect 1933 2273 1947 2287
rect 2013 2273 2027 2287
rect 2053 2273 2067 2287
rect 1733 2113 1747 2127
rect 1773 2113 1787 2127
rect 1833 2233 1847 2247
rect 1853 2213 1867 2227
rect 1813 2113 1827 2127
rect 1793 2093 1807 2107
rect 1773 2073 1787 2087
rect 1833 2093 1847 2107
rect 1713 1993 1727 2007
rect 1693 1913 1707 1927
rect 1693 1893 1707 1907
rect 1693 1833 1707 1847
rect 1753 1953 1767 1967
rect 1773 1813 1787 1827
rect 1693 1733 1707 1747
rect 1973 2193 1987 2207
rect 1933 2133 1947 2147
rect 2013 2133 2027 2147
rect 1993 2093 2007 2107
rect 2033 2113 2047 2127
rect 2053 2113 2067 2127
rect 1853 2033 1867 2047
rect 1853 1893 1867 1907
rect 1853 1873 1867 1887
rect 1833 1833 1847 1847
rect 1813 1813 1827 1827
rect 1833 1793 1847 1807
rect 1893 2033 1907 2047
rect 1953 1853 1967 1867
rect 1913 1813 1927 1827
rect 1893 1793 1907 1807
rect 1933 1793 1947 1807
rect 1813 1773 1827 1787
rect 1833 1773 1847 1787
rect 1873 1773 1887 1787
rect 1913 1773 1927 1787
rect 1933 1773 1947 1787
rect 1793 1713 1807 1727
rect 1793 1653 1807 1667
rect 1673 1633 1687 1647
rect 1693 1633 1707 1647
rect 1753 1633 1767 1647
rect 1553 1353 1567 1367
rect 1593 1533 1607 1547
rect 1633 1533 1647 1547
rect 1673 1593 1687 1607
rect 1593 1353 1607 1367
rect 1653 1353 1667 1367
rect 1713 1613 1727 1627
rect 1733 1593 1747 1607
rect 1773 1593 1787 1607
rect 1693 1553 1707 1567
rect 1753 1553 1767 1567
rect 1873 1733 1887 1747
rect 1833 1613 1847 1627
rect 1853 1613 1867 1627
rect 1813 1573 1827 1587
rect 1793 1393 1807 1407
rect 1713 1373 1727 1387
rect 1553 1313 1567 1327
rect 1573 1313 1587 1327
rect 1593 1313 1607 1327
rect 1673 1333 1687 1347
rect 1653 1313 1667 1327
rect 1613 1293 1627 1307
rect 1693 1293 1707 1307
rect 1553 1173 1567 1187
rect 1633 1153 1647 1167
rect 1673 1153 1687 1167
rect 1593 1133 1607 1147
rect 1573 1073 1587 1087
rect 1613 1113 1627 1127
rect 1533 993 1547 1007
rect 1373 973 1387 987
rect 1453 973 1467 987
rect 1293 933 1307 947
rect 1333 933 1347 947
rect 1373 893 1387 907
rect 1333 853 1347 867
rect 1353 833 1367 847
rect 1313 793 1327 807
rect 1273 773 1287 787
rect 1193 753 1207 767
rect 1333 753 1347 767
rect 1233 713 1247 727
rect 1233 653 1247 667
rect 1173 633 1187 647
rect 1353 713 1367 727
rect 1333 633 1347 647
rect 1113 613 1127 627
rect 1193 613 1207 627
rect 1233 613 1247 627
rect 1033 593 1047 607
rect 1073 373 1087 387
rect 1313 613 1327 627
rect 1273 573 1287 587
rect 1193 433 1207 447
rect 1253 433 1267 447
rect 913 313 927 327
rect 973 333 987 347
rect 1013 333 1027 347
rect 1053 333 1067 347
rect 1173 353 1187 367
rect 1153 333 1167 347
rect 1193 333 1207 347
rect 1253 333 1267 347
rect 893 293 907 307
rect 933 293 947 307
rect 853 213 867 227
rect 853 193 867 207
rect 973 313 987 327
rect 1093 313 1107 327
rect 953 253 967 267
rect 833 173 847 187
rect 913 173 927 187
rect 933 173 947 187
rect 853 153 867 167
rect 953 153 967 167
rect 673 133 687 147
rect 573 113 587 127
rect 633 113 647 127
rect 353 93 367 107
rect 493 93 507 107
rect 633 93 647 107
rect 33 53 47 67
rect 833 133 847 147
rect 853 113 867 127
rect 793 93 807 107
rect 933 133 947 147
rect 1153 313 1167 327
rect 1213 313 1227 327
rect 1113 253 1127 267
rect 1153 253 1167 267
rect 1113 233 1127 247
rect 1113 213 1127 227
rect 1093 173 1107 187
rect 1233 173 1247 187
rect 1073 133 1087 147
rect 1113 133 1127 147
rect 1173 133 1187 147
rect 1453 853 1467 867
rect 1433 833 1447 847
rect 1473 833 1487 847
rect 1433 813 1447 827
rect 1453 813 1467 827
rect 1493 813 1507 827
rect 1393 793 1407 807
rect 1413 653 1427 667
rect 1513 693 1527 707
rect 1693 1073 1707 1087
rect 1653 1013 1667 1027
rect 1613 873 1627 887
rect 1733 1333 1747 1347
rect 1793 1293 1807 1307
rect 1773 1193 1787 1207
rect 1833 1533 1847 1547
rect 1833 1473 1847 1487
rect 1773 1173 1787 1187
rect 1813 1173 1827 1187
rect 1733 1133 1747 1147
rect 1753 1113 1767 1127
rect 1793 1113 1807 1127
rect 1893 1593 1907 1607
rect 1933 1613 1947 1627
rect 1873 1573 1887 1587
rect 1873 1553 1887 1567
rect 2033 2013 2047 2027
rect 2033 1973 2047 1987
rect 2013 1873 2027 1887
rect 1993 1853 2007 1867
rect 2013 1793 2027 1807
rect 2073 2093 2087 2107
rect 2113 2173 2127 2187
rect 2153 2173 2167 2187
rect 2133 2153 2147 2167
rect 2393 2553 2407 2567
rect 2433 2853 2447 2867
rect 2533 3693 2547 3707
rect 2753 4653 2767 4667
rect 2773 4613 2787 4627
rect 2833 4613 2847 4627
rect 2713 4593 2727 4607
rect 2873 4593 2887 4607
rect 2773 4573 2787 4587
rect 2753 4553 2767 4567
rect 2733 4533 2747 4547
rect 2693 4513 2707 4527
rect 2713 4453 2727 4467
rect 2673 4213 2687 4227
rect 2693 4173 2707 4187
rect 2753 4453 2767 4467
rect 3033 4953 3047 4967
rect 3233 5433 3247 5447
rect 3153 5393 3167 5407
rect 3273 5413 3287 5427
rect 3193 5373 3207 5387
rect 3293 5373 3307 5387
rect 3293 5353 3307 5367
rect 3273 5333 3287 5347
rect 3233 5153 3247 5167
rect 3153 5113 3167 5127
rect 3113 5073 3127 5087
rect 3113 5053 3127 5067
rect 3093 4993 3107 5007
rect 3113 4973 3127 4987
rect 3013 4753 3027 4767
rect 3013 4733 3027 4747
rect 2913 4713 2927 4727
rect 2973 4713 2987 4727
rect 2993 4713 3007 4727
rect 2953 4693 2967 4707
rect 2933 4673 2947 4687
rect 2913 4653 2927 4667
rect 2893 4573 2907 4587
rect 2873 4513 2887 4527
rect 2813 4493 2827 4507
rect 3133 4893 3147 4907
rect 3093 4713 3107 4727
rect 3053 4693 3067 4707
rect 3073 4693 3087 4707
rect 3033 4673 3047 4687
rect 2953 4653 2967 4667
rect 2973 4653 2987 4667
rect 2933 4553 2947 4567
rect 2933 4513 2947 4527
rect 2853 4473 2867 4487
rect 2893 4473 2907 4487
rect 2913 4473 2927 4487
rect 2793 4433 2807 4447
rect 2813 4253 2827 4267
rect 2753 4173 2767 4187
rect 2833 4233 2847 4247
rect 2773 4113 2787 4127
rect 2733 4073 2747 4087
rect 2713 4033 2727 4047
rect 2653 4013 2667 4027
rect 2653 3973 2667 3987
rect 2733 3973 2747 3987
rect 2713 3953 2727 3967
rect 2993 4613 3007 4627
rect 2973 4513 2987 4527
rect 2973 4473 2987 4487
rect 2933 4233 2947 4247
rect 2973 4233 2987 4247
rect 2853 4173 2867 4187
rect 2833 4013 2847 4027
rect 2813 3993 2827 4007
rect 2913 4173 2927 4187
rect 2873 4153 2887 4167
rect 2873 4013 2887 4027
rect 2773 3973 2787 3987
rect 2693 3933 2707 3947
rect 2893 3993 2907 4007
rect 2833 3953 2847 3967
rect 2833 3933 2847 3947
rect 2793 3893 2807 3907
rect 2893 3873 2907 3887
rect 3073 4553 3087 4567
rect 3013 4513 3027 4527
rect 3033 4473 3047 4487
rect 3053 4453 3067 4467
rect 3133 4693 3147 4707
rect 3113 4613 3127 4627
rect 3213 5113 3227 5127
rect 3193 5013 3207 5027
rect 3173 4993 3187 5007
rect 3173 4933 3187 4947
rect 3153 4593 3167 4607
rect 3233 4933 3247 4947
rect 3253 4913 3267 4927
rect 3193 4733 3207 4747
rect 3213 4713 3227 4727
rect 3253 4693 3267 4707
rect 3193 4653 3207 4667
rect 3233 4653 3247 4667
rect 3173 4573 3187 4587
rect 3113 4533 3127 4547
rect 3193 4533 3207 4547
rect 3153 4513 3167 4527
rect 3213 4513 3227 4527
rect 3353 5473 3367 5487
rect 3393 5473 3407 5487
rect 3493 5473 3507 5487
rect 5253 5473 5267 5487
rect 5313 5473 5327 5487
rect 3373 5393 3387 5407
rect 3313 5313 3327 5327
rect 3413 5453 3427 5467
rect 3593 5453 3607 5467
rect 3733 5453 3747 5467
rect 3473 5413 3487 5427
rect 3453 5393 3467 5407
rect 3433 5213 3447 5227
rect 3393 5193 3407 5207
rect 3393 5173 3407 5187
rect 3353 5153 3367 5167
rect 3373 5133 3387 5147
rect 3513 5373 3527 5387
rect 3613 5433 3627 5447
rect 3633 5393 3647 5407
rect 3613 5373 3627 5387
rect 3553 5353 3567 5367
rect 3473 5173 3487 5187
rect 3493 5153 3507 5167
rect 3473 5133 3487 5147
rect 3333 5093 3347 5107
rect 3453 5093 3467 5107
rect 3533 5133 3547 5147
rect 3573 5153 3587 5167
rect 3693 5433 3707 5447
rect 3833 5413 3847 5427
rect 3853 5393 3867 5407
rect 3913 5413 3927 5427
rect 4613 5453 4627 5467
rect 5033 5453 5047 5467
rect 5273 5453 5287 5467
rect 4013 5433 4027 5447
rect 4093 5433 4107 5447
rect 4133 5433 4147 5447
rect 4253 5433 4267 5447
rect 4293 5433 4307 5447
rect 4353 5433 4367 5447
rect 4513 5433 4527 5447
rect 3773 5373 3787 5387
rect 3673 5353 3687 5367
rect 3713 5353 3727 5367
rect 3833 5193 3847 5207
rect 3813 5173 3827 5187
rect 3653 5153 3667 5167
rect 3693 5153 3707 5167
rect 3553 5113 3567 5127
rect 3633 5133 3647 5147
rect 3673 5133 3687 5147
rect 3593 5113 3607 5127
rect 3673 5113 3687 5127
rect 3673 5093 3687 5107
rect 3573 5053 3587 5067
rect 3513 5013 3527 5027
rect 3393 4993 3407 5007
rect 3433 4993 3447 5007
rect 3353 4973 3367 4987
rect 3573 4973 3587 4987
rect 3413 4953 3427 4967
rect 3333 4933 3347 4947
rect 3293 4913 3307 4927
rect 3393 4933 3407 4947
rect 3433 4933 3447 4947
rect 3333 4893 3347 4907
rect 3373 4893 3387 4907
rect 3313 4753 3327 4767
rect 3293 4693 3307 4707
rect 3293 4613 3307 4627
rect 3293 4553 3307 4567
rect 3213 4493 3227 4507
rect 3273 4493 3287 4507
rect 3173 4433 3187 4447
rect 3153 4353 3167 4367
rect 3133 4313 3147 4327
rect 3093 4253 3107 4267
rect 3113 4233 3127 4247
rect 2993 4213 3007 4227
rect 3093 4213 3107 4227
rect 2973 4193 2987 4207
rect 2953 4173 2967 4187
rect 2953 4093 2967 4107
rect 3073 4153 3087 4167
rect 3033 4093 3047 4107
rect 2993 4073 3007 4087
rect 3033 4073 3047 4087
rect 3073 4073 3087 4087
rect 2993 4013 3007 4027
rect 2953 3973 2967 3987
rect 2973 3973 2987 3987
rect 3033 3973 3047 3987
rect 3133 4173 3147 4187
rect 3133 4153 3147 4167
rect 3193 4313 3207 4327
rect 3173 4213 3187 4227
rect 3193 4173 3207 4187
rect 3353 4833 3367 4847
rect 3333 4633 3347 4647
rect 3313 4493 3327 4507
rect 3413 4673 3427 4687
rect 3393 4653 3407 4667
rect 3373 4613 3387 4627
rect 3393 4593 3407 4607
rect 3373 4573 3387 4587
rect 3353 4553 3367 4567
rect 3273 4453 3287 4467
rect 3233 4433 3247 4447
rect 3253 4433 3267 4447
rect 3313 4433 3327 4447
rect 3333 4433 3347 4447
rect 3233 4153 3247 4167
rect 3233 4033 3247 4047
rect 3093 3993 3107 4007
rect 2993 3953 3007 3967
rect 3053 3953 3067 3967
rect 3073 3953 3087 3967
rect 3053 3933 3067 3947
rect 3093 3933 3107 3947
rect 3013 3873 3027 3887
rect 2993 3853 3007 3867
rect 2933 3813 2947 3827
rect 2973 3813 2987 3827
rect 2673 3793 2687 3807
rect 2613 3733 2627 3747
rect 2633 3733 2647 3747
rect 2593 3573 2607 3587
rect 2533 3553 2547 3567
rect 2573 3553 2587 3567
rect 2553 3533 2567 3547
rect 2593 3533 2607 3547
rect 2533 3493 2547 3507
rect 2573 3493 2587 3507
rect 2593 3493 2607 3507
rect 2553 3253 2567 3267
rect 2613 3473 2627 3487
rect 2613 3453 2627 3467
rect 2613 3413 2627 3427
rect 2673 3673 2687 3687
rect 2693 3633 2707 3647
rect 2773 3553 2787 3567
rect 2853 3553 2867 3567
rect 2693 3533 2707 3547
rect 2653 3513 2667 3527
rect 2713 3513 2727 3527
rect 2813 3513 2827 3527
rect 2753 3473 2767 3487
rect 2753 3453 2767 3467
rect 2673 3393 2687 3407
rect 2713 3353 2727 3367
rect 2633 3333 2647 3347
rect 2613 3273 2627 3287
rect 2553 3233 2567 3247
rect 2533 3173 2547 3187
rect 2533 3153 2547 3167
rect 2513 3093 2527 3107
rect 2513 3053 2527 3067
rect 2573 3213 2587 3227
rect 2653 3293 2667 3307
rect 2633 3233 2647 3247
rect 2713 3273 2727 3287
rect 2673 3233 2687 3247
rect 2653 3213 2667 3227
rect 2693 3213 2707 3227
rect 2733 3213 2747 3227
rect 2613 3193 2627 3207
rect 2573 3153 2587 3167
rect 2733 3153 2747 3167
rect 2493 2833 2507 2847
rect 2673 3133 2687 3147
rect 2713 3133 2727 3147
rect 2613 3113 2627 3127
rect 2653 3113 2667 3127
rect 2593 3073 2607 3087
rect 2573 3033 2587 3047
rect 2533 2973 2547 2987
rect 2573 2953 2587 2967
rect 2633 3093 2647 3107
rect 2613 3053 2627 3067
rect 2593 2893 2607 2907
rect 2533 2853 2547 2867
rect 2533 2833 2547 2847
rect 2513 2813 2527 2827
rect 2433 2773 2447 2787
rect 2473 2773 2487 2787
rect 2513 2773 2527 2787
rect 2453 2693 2467 2707
rect 2473 2653 2487 2667
rect 2453 2553 2467 2567
rect 2633 3033 2647 3047
rect 2693 3073 2707 3087
rect 2613 2793 2627 2807
rect 2773 3353 2787 3367
rect 2833 3493 2847 3507
rect 2833 3393 2847 3407
rect 2793 3273 2807 3287
rect 2793 3233 2807 3247
rect 2953 3633 2967 3647
rect 2933 3613 2947 3627
rect 2893 3493 2907 3507
rect 2893 3413 2907 3427
rect 2993 3713 3007 3727
rect 3013 3653 3027 3667
rect 2973 3513 2987 3527
rect 3093 3893 3107 3907
rect 3073 3673 3087 3687
rect 3053 3613 3067 3627
rect 3133 3973 3147 3987
rect 3153 3973 3167 3987
rect 3133 3933 3147 3947
rect 3153 3873 3167 3887
rect 3133 3713 3147 3727
rect 3173 3753 3187 3767
rect 3273 4273 3287 4287
rect 3413 4573 3427 4587
rect 3473 4913 3487 4927
rect 3453 4653 3467 4667
rect 3433 4513 3447 4527
rect 3373 4353 3387 4367
rect 3373 4333 3387 4347
rect 3353 4273 3367 4287
rect 3433 4453 3447 4467
rect 3413 4433 3427 4447
rect 3273 4213 3287 4227
rect 3333 4213 3347 4227
rect 3313 4173 3327 4187
rect 3293 4073 3307 4087
rect 3253 3993 3267 4007
rect 3273 3993 3287 4007
rect 3253 3973 3267 3987
rect 3273 3973 3287 3987
rect 3313 4033 3327 4047
rect 3393 4233 3407 4247
rect 3413 4233 3427 4247
rect 3453 4233 3467 4247
rect 3373 4213 3387 4227
rect 3613 4933 3627 4947
rect 3593 4913 3607 4927
rect 3553 4853 3567 4867
rect 3533 4653 3547 4667
rect 3493 4613 3507 4627
rect 3493 4533 3507 4547
rect 3573 4673 3587 4687
rect 3633 4893 3647 4907
rect 3673 4833 3687 4847
rect 3753 5133 3767 5147
rect 3713 5113 3727 5127
rect 3733 5113 3747 5127
rect 3793 5113 3807 5127
rect 3773 5013 3787 5027
rect 3753 4993 3767 5007
rect 3853 5133 3867 5147
rect 3893 5173 3907 5187
rect 3933 5173 3947 5187
rect 3873 5093 3887 5107
rect 3993 5373 4007 5387
rect 3993 5353 4007 5367
rect 4073 5413 4087 5427
rect 4113 5413 4127 5427
rect 4213 5413 4227 5427
rect 4313 5413 4327 5427
rect 4193 5393 4207 5407
rect 4233 5393 4247 5407
rect 4273 5393 4287 5407
rect 4213 5373 4227 5387
rect 4193 5333 4207 5347
rect 4013 5193 4027 5207
rect 4053 5173 4067 5187
rect 3993 5153 4007 5167
rect 3973 5133 3987 5147
rect 4013 5133 4027 5147
rect 4013 5113 4027 5127
rect 3953 5053 3967 5067
rect 3853 4973 3867 4987
rect 3793 4933 3807 4947
rect 3733 4913 3747 4927
rect 3693 4733 3707 4747
rect 3733 4733 3747 4747
rect 3613 4713 3627 4727
rect 3633 4713 3647 4727
rect 3653 4693 3667 4707
rect 3673 4673 3687 4687
rect 3713 4673 3727 4687
rect 3633 4653 3647 4667
rect 3693 4653 3707 4667
rect 3573 4633 3587 4647
rect 3553 4593 3567 4607
rect 3713 4613 3727 4627
rect 3493 4473 3507 4487
rect 3533 4473 3547 4487
rect 3513 4453 3527 4467
rect 3593 4553 3607 4567
rect 3573 4513 3587 4527
rect 3573 4473 3587 4487
rect 3713 4513 3727 4527
rect 3653 4493 3667 4507
rect 3613 4453 3627 4467
rect 3533 4433 3547 4447
rect 3553 4433 3567 4447
rect 3513 4413 3527 4427
rect 3433 4213 3447 4227
rect 3473 4213 3487 4227
rect 3393 4193 3407 4207
rect 3393 4153 3407 4167
rect 3393 4033 3407 4047
rect 3213 3953 3227 3967
rect 3233 3933 3247 3947
rect 3173 3733 3187 3747
rect 3213 3733 3227 3747
rect 3153 3673 3167 3687
rect 3153 3633 3167 3647
rect 3113 3593 3127 3607
rect 3173 3593 3187 3607
rect 3153 3533 3167 3547
rect 3153 3493 3167 3507
rect 3013 3453 3027 3467
rect 2953 3413 2967 3427
rect 2873 3353 2887 3367
rect 2873 3333 2887 3347
rect 2853 3313 2867 3327
rect 2853 3253 2867 3267
rect 2793 3193 2807 3207
rect 2753 3133 2767 3147
rect 2773 3033 2787 3047
rect 2733 3013 2747 3027
rect 2753 3013 2767 3027
rect 2733 2993 2747 3007
rect 2713 2793 2727 2807
rect 2573 2773 2587 2787
rect 2553 2733 2567 2747
rect 2493 2593 2507 2607
rect 2513 2573 2527 2587
rect 2413 2533 2427 2547
rect 2213 2373 2227 2387
rect 2273 2313 2287 2327
rect 2573 2713 2587 2727
rect 2613 2693 2627 2707
rect 2593 2633 2607 2647
rect 2693 2693 2707 2707
rect 2773 2953 2787 2967
rect 2773 2913 2787 2927
rect 2753 2793 2767 2807
rect 2773 2713 2787 2727
rect 2733 2613 2747 2627
rect 2613 2593 2627 2607
rect 2653 2593 2667 2607
rect 2493 2533 2507 2547
rect 2513 2533 2527 2547
rect 2493 2433 2507 2447
rect 2213 2253 2227 2267
rect 2173 2113 2187 2127
rect 2133 2093 2147 2107
rect 2173 2093 2187 2107
rect 2073 2053 2087 2067
rect 2113 2053 2127 2067
rect 2093 2013 2107 2027
rect 2073 1793 2087 1807
rect 2073 1773 2087 1787
rect 2053 1753 2067 1767
rect 2013 1733 2027 1747
rect 2053 1733 2067 1747
rect 2013 1593 2027 1607
rect 1853 1453 1867 1467
rect 1853 1333 1867 1347
rect 1913 1433 1927 1447
rect 1893 1333 1907 1347
rect 1873 1313 1887 1327
rect 1873 1273 1887 1287
rect 1993 1553 2007 1567
rect 1993 1513 2007 1527
rect 1973 1373 1987 1387
rect 1953 1353 1967 1367
rect 1933 1333 1947 1347
rect 1953 1313 1967 1327
rect 1913 1293 1927 1307
rect 1913 1273 1927 1287
rect 1893 1133 1907 1147
rect 1853 1113 1867 1127
rect 1853 1093 1867 1107
rect 1813 953 1827 967
rect 1733 893 1747 907
rect 1713 873 1727 887
rect 1653 853 1667 867
rect 1873 1073 1887 1087
rect 2013 1373 2027 1387
rect 2073 1613 2087 1627
rect 2253 2213 2267 2227
rect 2233 2133 2247 2147
rect 2193 2073 2207 2087
rect 2213 2073 2227 2087
rect 2173 2013 2187 2027
rect 2133 1993 2147 2007
rect 2153 1993 2167 2007
rect 2173 1873 2187 1887
rect 2153 1813 2167 1827
rect 2113 1773 2127 1787
rect 2113 1713 2127 1727
rect 2073 1553 2087 1567
rect 2093 1553 2107 1567
rect 2053 1533 2067 1547
rect 2093 1533 2107 1547
rect 2033 1353 2047 1367
rect 2133 1573 2147 1587
rect 2133 1533 2147 1547
rect 2113 1513 2127 1527
rect 2113 1453 2127 1467
rect 2053 1333 2067 1347
rect 2053 1313 2067 1327
rect 2033 1293 2047 1307
rect 2033 1213 2047 1227
rect 1993 1173 2007 1187
rect 1993 1133 2007 1147
rect 1853 1053 1867 1067
rect 1773 873 1787 887
rect 1833 873 1847 887
rect 1633 833 1647 847
rect 1593 813 1607 827
rect 1713 833 1727 847
rect 1573 733 1587 747
rect 1573 693 1587 707
rect 1553 673 1567 687
rect 1373 613 1387 627
rect 1653 613 1667 627
rect 1673 613 1687 627
rect 1753 813 1767 827
rect 1973 1093 1987 1107
rect 2013 1093 2027 1107
rect 1933 1013 1947 1027
rect 2033 953 2047 967
rect 2093 1273 2107 1287
rect 2073 1133 2087 1147
rect 2133 1413 2147 1427
rect 2173 1693 2187 1707
rect 2253 2033 2267 2047
rect 2253 1893 2267 1907
rect 2353 2293 2367 2307
rect 2373 2293 2387 2307
rect 2313 2273 2327 2287
rect 2293 2253 2307 2267
rect 2413 2273 2427 2287
rect 2313 2233 2327 2247
rect 2333 2233 2347 2247
rect 2313 2193 2327 2207
rect 2333 2053 2347 2067
rect 2353 2013 2367 2027
rect 2313 1993 2327 2007
rect 2453 2253 2467 2267
rect 2433 2193 2447 2207
rect 2453 2193 2467 2207
rect 2433 2173 2447 2187
rect 2393 2133 2407 2147
rect 2413 2093 2427 2107
rect 2493 2233 2507 2247
rect 2553 2533 2567 2547
rect 2533 2433 2547 2447
rect 2553 2433 2567 2447
rect 2653 2573 2667 2587
rect 2633 2553 2647 2567
rect 2633 2513 2647 2527
rect 2613 2473 2627 2487
rect 2573 2393 2587 2407
rect 2573 2373 2587 2387
rect 2513 2213 2527 2227
rect 2533 2193 2547 2207
rect 2553 2193 2567 2207
rect 2473 2173 2487 2187
rect 2513 2173 2527 2187
rect 2533 2173 2547 2187
rect 2453 2093 2467 2107
rect 2473 2093 2487 2107
rect 2493 2093 2507 2107
rect 2453 2033 2467 2047
rect 2413 2013 2427 2027
rect 2453 2013 2467 2027
rect 2493 2013 2507 2027
rect 2393 1893 2407 1907
rect 2373 1873 2387 1887
rect 2273 1833 2287 1847
rect 2313 1833 2327 1847
rect 2333 1833 2347 1847
rect 2293 1793 2307 1807
rect 2233 1773 2247 1787
rect 2313 1773 2327 1787
rect 2393 1813 2407 1827
rect 2373 1793 2387 1807
rect 2393 1753 2407 1767
rect 2353 1733 2367 1747
rect 2313 1713 2327 1727
rect 2313 1673 2327 1687
rect 2193 1653 2207 1667
rect 2213 1653 2227 1667
rect 2253 1613 2267 1627
rect 2233 1573 2247 1587
rect 2253 1573 2267 1587
rect 2213 1433 2227 1447
rect 2153 1393 2167 1407
rect 2173 1313 2187 1327
rect 2133 1293 2147 1307
rect 2133 1273 2147 1287
rect 2193 1293 2207 1307
rect 2073 1113 2087 1127
rect 2113 1113 2127 1127
rect 2113 1093 2127 1107
rect 2093 1073 2107 1087
rect 2073 1053 2087 1067
rect 2093 1053 2107 1067
rect 1933 893 1947 907
rect 2053 893 2067 907
rect 1893 873 1907 887
rect 1773 773 1787 787
rect 1473 593 1487 607
rect 1393 553 1407 567
rect 1433 553 1447 567
rect 1373 373 1387 387
rect 1453 373 1467 387
rect 1353 353 1367 367
rect 1393 353 1407 367
rect 1433 353 1447 367
rect 1333 333 1347 347
rect 1593 593 1607 607
rect 1633 593 1647 607
rect 1673 593 1687 607
rect 1553 573 1567 587
rect 1733 573 1747 587
rect 1673 533 1687 547
rect 1713 533 1727 547
rect 1573 493 1587 507
rect 1513 433 1527 447
rect 1473 353 1487 367
rect 1553 393 1567 407
rect 1453 333 1467 347
rect 1313 313 1327 327
rect 1433 313 1447 327
rect 1453 313 1467 327
rect 1493 313 1507 327
rect 1393 213 1407 227
rect 1293 193 1307 207
rect 1653 373 1667 387
rect 1613 353 1627 367
rect 1633 333 1647 347
rect 1653 333 1667 347
rect 1593 313 1607 327
rect 1853 853 1867 867
rect 1953 873 1967 887
rect 1833 833 1847 847
rect 1813 733 1827 747
rect 1913 813 1927 827
rect 1913 773 1927 787
rect 1873 693 1887 707
rect 1833 673 1847 687
rect 1893 653 1907 667
rect 1853 613 1867 627
rect 1793 553 1807 567
rect 1713 433 1727 447
rect 1773 433 1787 447
rect 1693 413 1707 427
rect 1673 293 1687 307
rect 1653 193 1667 207
rect 1773 393 1787 407
rect 1773 373 1787 387
rect 1893 573 1907 587
rect 1893 513 1907 527
rect 1873 473 1887 487
rect 1933 753 1947 767
rect 2033 853 2047 867
rect 2073 853 2087 867
rect 1993 813 2007 827
rect 2053 813 2067 827
rect 2133 1033 2147 1047
rect 2093 813 2107 827
rect 2433 1993 2447 2007
rect 2453 1933 2467 1947
rect 2433 1813 2447 1827
rect 2553 2153 2567 2167
rect 2593 2253 2607 2267
rect 2593 2153 2607 2167
rect 2573 2093 2587 2107
rect 2693 2473 2707 2487
rect 2653 2313 2667 2327
rect 2713 2433 2727 2447
rect 2693 2293 2707 2307
rect 2653 2253 2667 2267
rect 2773 2613 2787 2627
rect 2933 3293 2947 3307
rect 2873 3193 2887 3207
rect 2853 3153 2867 3167
rect 2853 3133 2867 3147
rect 3133 3393 3147 3407
rect 3093 3353 3107 3367
rect 2993 3273 3007 3287
rect 3073 3273 3087 3287
rect 3053 3253 3067 3267
rect 2973 3213 2987 3227
rect 3013 3213 3027 3227
rect 2953 3193 2967 3207
rect 2913 3153 2927 3167
rect 2973 3153 2987 3167
rect 2833 3053 2847 3067
rect 2873 3053 2887 3067
rect 2893 3013 2907 3027
rect 2853 2993 2867 3007
rect 3013 3093 3027 3107
rect 2953 3073 2967 3087
rect 2933 3033 2947 3047
rect 2913 2973 2927 2987
rect 2833 2933 2847 2947
rect 2833 2833 2847 2847
rect 2973 3033 2987 3047
rect 3153 3353 3167 3367
rect 3273 3813 3287 3827
rect 3373 3973 3387 3987
rect 3373 3953 3387 3967
rect 3333 3813 3347 3827
rect 3273 3793 3287 3807
rect 3313 3793 3327 3807
rect 3253 3753 3267 3767
rect 3233 3693 3247 3707
rect 3313 3753 3327 3767
rect 3353 3733 3367 3747
rect 3393 3733 3407 3747
rect 3313 3713 3327 3727
rect 3293 3613 3307 3627
rect 3333 3613 3347 3627
rect 3253 3593 3267 3607
rect 3193 3573 3207 3587
rect 3253 3533 3267 3547
rect 3213 3353 3227 3367
rect 3193 3333 3207 3347
rect 3173 3273 3187 3287
rect 3133 3233 3147 3247
rect 3173 3233 3187 3247
rect 3093 3213 3107 3227
rect 3133 3193 3147 3207
rect 3153 3193 3167 3207
rect 3113 3153 3127 3167
rect 3093 3093 3107 3107
rect 3073 3073 3087 3087
rect 3033 3053 3047 3067
rect 3033 3033 3047 3047
rect 3073 3033 3087 3047
rect 3113 3073 3127 3087
rect 2953 2953 2967 2967
rect 2853 2773 2867 2787
rect 2813 2753 2827 2767
rect 2873 2753 2887 2767
rect 2933 2773 2947 2787
rect 2913 2733 2927 2747
rect 2833 2713 2847 2727
rect 3093 3013 3107 3027
rect 3053 2973 3067 2987
rect 2993 2873 3007 2887
rect 3153 3173 3167 3187
rect 3233 3213 3247 3227
rect 3193 3193 3207 3207
rect 3213 3133 3227 3147
rect 3193 3113 3207 3127
rect 3173 3053 3187 3067
rect 3193 3013 3207 3027
rect 3153 2973 3167 2987
rect 3133 2953 3147 2967
rect 3073 2793 3087 2807
rect 3113 2793 3127 2807
rect 2993 2773 3007 2787
rect 3033 2773 3047 2787
rect 2973 2753 2987 2767
rect 3013 2733 3027 2747
rect 2973 2633 2987 2647
rect 2953 2593 2967 2607
rect 2793 2553 2807 2567
rect 2753 2473 2767 2487
rect 3113 2773 3127 2787
rect 3093 2733 3107 2747
rect 3333 3573 3347 3587
rect 3273 3493 3287 3507
rect 3293 3493 3307 3507
rect 3313 3453 3327 3467
rect 3313 3333 3327 3347
rect 3253 3133 3267 3147
rect 3273 3093 3287 3107
rect 3233 3073 3247 3087
rect 3233 3053 3247 3067
rect 3313 3073 3327 3087
rect 3393 3553 3407 3567
rect 3353 3533 3367 3547
rect 3513 4173 3527 4187
rect 3493 4153 3507 4167
rect 3473 4093 3487 4107
rect 3473 4073 3487 4087
rect 3473 4033 3487 4047
rect 3493 3953 3507 3967
rect 3553 4413 3567 4427
rect 3753 4693 3767 4707
rect 3853 4933 3867 4947
rect 3833 4913 3847 4927
rect 3913 4993 3927 5007
rect 3913 4973 3927 4987
rect 4053 5133 4067 5147
rect 4173 5173 4187 5187
rect 4113 5113 4127 5127
rect 4153 5113 4167 5127
rect 4173 5113 4187 5127
rect 4033 4973 4047 4987
rect 4053 4973 4067 4987
rect 4133 4973 4147 4987
rect 3973 4953 3987 4967
rect 4033 4953 4047 4967
rect 4093 4953 4107 4967
rect 4113 4953 4127 4967
rect 3893 4873 3907 4887
rect 3873 4833 3887 4847
rect 3833 4713 3847 4727
rect 3893 4713 3907 4727
rect 3933 4713 3947 4727
rect 3813 4673 3827 4687
rect 3813 4633 3827 4647
rect 3873 4633 3887 4647
rect 3773 4613 3787 4627
rect 3873 4553 3887 4567
rect 3753 4513 3767 4527
rect 3833 4513 3847 4527
rect 3733 4473 3747 4487
rect 3713 4453 3727 4467
rect 3613 4233 3627 4247
rect 3653 4233 3667 4247
rect 3553 4213 3567 4227
rect 3573 4193 3587 4207
rect 3553 4173 3567 4187
rect 3593 4153 3607 4167
rect 3553 4073 3567 4087
rect 3593 4073 3607 4087
rect 3573 4033 3587 4047
rect 3633 4193 3647 4207
rect 3673 4193 3687 4207
rect 3793 4493 3807 4507
rect 3813 4493 3827 4507
rect 3793 4433 3807 4447
rect 3753 4213 3767 4227
rect 3693 4153 3707 4167
rect 3653 4133 3667 4147
rect 3653 4033 3667 4047
rect 3693 4033 3707 4047
rect 3533 3953 3547 3967
rect 3513 3813 3527 3827
rect 3513 3793 3527 3807
rect 3453 3753 3467 3767
rect 3433 3733 3447 3747
rect 3453 3733 3467 3747
rect 3493 3713 3507 3727
rect 3433 3693 3447 3707
rect 3473 3693 3487 3707
rect 3493 3673 3507 3687
rect 3433 3593 3447 3607
rect 3413 3533 3427 3547
rect 3613 3773 3627 3787
rect 3553 3693 3567 3707
rect 3593 3693 3607 3707
rect 3573 3613 3587 3627
rect 3673 3733 3687 3747
rect 3633 3713 3647 3727
rect 3613 3593 3627 3607
rect 3653 3573 3667 3587
rect 3533 3553 3547 3567
rect 3413 3493 3427 3507
rect 3473 3493 3487 3507
rect 3473 3373 3487 3387
rect 3513 3493 3527 3507
rect 3773 4173 3787 4187
rect 3733 4153 3747 4167
rect 3753 4153 3767 4167
rect 3713 4013 3727 4027
rect 3773 4093 3787 4107
rect 3753 4073 3767 4087
rect 3753 4013 3767 4027
rect 3913 4693 3927 4707
rect 4073 4913 4087 4927
rect 4133 4913 4147 4927
rect 4073 4893 4087 4907
rect 3973 4713 3987 4727
rect 4053 4713 4067 4727
rect 4013 4693 4027 4707
rect 4033 4693 4047 4707
rect 3993 4673 4007 4687
rect 3953 4653 3967 4667
rect 4053 4673 4067 4687
rect 3973 4633 3987 4647
rect 4033 4633 4047 4647
rect 3933 4613 3947 4627
rect 3893 4533 3907 4547
rect 3893 4493 3907 4507
rect 3933 4493 3947 4507
rect 3953 4493 3967 4507
rect 3873 4233 3887 4247
rect 3913 4473 3927 4487
rect 3993 4573 4007 4587
rect 4113 4693 4127 4707
rect 4153 4673 4167 4687
rect 4133 4633 4147 4647
rect 4093 4573 4107 4587
rect 4073 4513 4087 4527
rect 4013 4493 4027 4507
rect 4033 4493 4047 4507
rect 4053 4493 4067 4507
rect 3973 4453 3987 4467
rect 3973 4313 3987 4327
rect 3913 4233 3927 4247
rect 4113 4533 4127 4547
rect 4213 5113 4227 5127
rect 4393 5413 4407 5427
rect 4433 5413 4447 5427
rect 4453 5413 4467 5427
rect 4493 5413 4507 5427
rect 4313 5373 4327 5387
rect 4293 5213 4307 5227
rect 4413 5353 4427 5367
rect 4433 5353 4447 5367
rect 4753 5433 4767 5447
rect 4893 5433 4907 5447
rect 4953 5433 4967 5447
rect 5173 5433 5187 5447
rect 5193 5433 5207 5447
rect 5233 5433 5247 5447
rect 4473 5373 4487 5387
rect 4453 5333 4467 5347
rect 4513 5193 4527 5207
rect 4373 5173 4387 5187
rect 4413 5173 4427 5187
rect 4393 5153 4407 5167
rect 4353 5113 4367 5127
rect 4293 5093 4307 5107
rect 4333 5093 4347 5107
rect 4453 5153 4467 5167
rect 4653 5413 4667 5427
rect 4693 5413 4707 5427
rect 4593 5353 4607 5367
rect 4713 5393 4727 5407
rect 4793 5413 4807 5427
rect 4873 5413 4887 5427
rect 5013 5413 5027 5427
rect 5133 5413 5147 5427
rect 4813 5333 4827 5347
rect 4693 5313 4707 5327
rect 4613 5173 4627 5187
rect 4553 5153 4567 5167
rect 4393 5113 4407 5127
rect 4373 5053 4387 5067
rect 4273 5033 4287 5047
rect 4353 5033 4367 5047
rect 4273 5013 4287 5027
rect 4293 5013 4307 5027
rect 4233 4933 4247 4947
rect 4213 4913 4227 4927
rect 4513 5133 4527 5147
rect 4473 5113 4487 5127
rect 4513 5093 4527 5107
rect 4553 5093 4567 5107
rect 4573 5093 4587 5107
rect 4533 5013 4547 5027
rect 4413 4973 4427 4987
rect 4493 4973 4507 4987
rect 4533 4973 4547 4987
rect 4433 4953 4447 4967
rect 4413 4913 4427 4927
rect 4453 4913 4467 4927
rect 4313 4893 4327 4907
rect 4353 4893 4367 4907
rect 4313 4833 4327 4847
rect 4373 4833 4387 4847
rect 4233 4733 4247 4747
rect 4253 4733 4267 4747
rect 4313 4693 4327 4707
rect 4673 5113 4687 5127
rect 4633 4953 4647 4967
rect 4573 4933 4587 4947
rect 4513 4913 4527 4927
rect 4633 4913 4647 4927
rect 4593 4893 4607 4907
rect 4493 4713 4507 4727
rect 4193 4673 4207 4687
rect 4233 4673 4247 4687
rect 4373 4653 4387 4667
rect 4193 4633 4207 4647
rect 4333 4633 4347 4647
rect 4173 4553 4187 4567
rect 4153 4493 4167 4507
rect 4133 4473 4147 4487
rect 4113 4413 4127 4427
rect 3813 4133 3827 4147
rect 3893 4153 3907 4167
rect 3853 4113 3867 4127
rect 3793 4033 3807 4047
rect 3813 4013 3827 4027
rect 3733 3993 3747 4007
rect 3793 3993 3807 4007
rect 3853 3993 3867 4007
rect 3833 3973 3847 3987
rect 3873 3973 3887 3987
rect 3853 3813 3867 3827
rect 3773 3733 3787 3747
rect 3733 3713 3747 3727
rect 3753 3713 3767 3727
rect 3833 3713 3847 3727
rect 3773 3673 3787 3687
rect 3833 3673 3847 3687
rect 3733 3593 3747 3607
rect 3713 3553 3727 3567
rect 3613 3533 3627 3547
rect 3693 3533 3707 3547
rect 3553 3513 3567 3527
rect 3493 3293 3507 3307
rect 3353 3233 3367 3247
rect 3353 3153 3367 3167
rect 3353 3133 3367 3147
rect 3473 3113 3487 3127
rect 3453 3053 3467 3067
rect 3313 3033 3327 3047
rect 3333 3033 3347 3047
rect 3293 2993 3307 3007
rect 3233 2833 3247 2847
rect 3213 2813 3227 2827
rect 3213 2793 3227 2807
rect 3253 2793 3267 2807
rect 3173 2733 3187 2747
rect 3153 2713 3167 2727
rect 3233 2733 3247 2747
rect 3273 2713 3287 2727
rect 3233 2693 3247 2707
rect 3213 2633 3227 2647
rect 3133 2593 3147 2607
rect 3213 2593 3227 2607
rect 3173 2573 3187 2587
rect 3053 2553 3067 2567
rect 3073 2553 3087 2567
rect 3133 2553 3147 2567
rect 3093 2513 3107 2527
rect 3053 2493 3067 2507
rect 2933 2433 2947 2447
rect 2973 2433 2987 2447
rect 2913 2393 2927 2407
rect 2893 2373 2907 2387
rect 2733 2293 2747 2307
rect 2793 2293 2807 2307
rect 2653 2233 2667 2247
rect 2633 2133 2647 2147
rect 2633 2113 2647 2127
rect 2613 2073 2627 2087
rect 2673 2193 2687 2207
rect 2693 2193 2707 2207
rect 2773 2253 2787 2267
rect 2753 2233 2767 2247
rect 2733 2213 2747 2227
rect 2713 2173 2727 2187
rect 2573 2033 2587 2047
rect 2533 2013 2547 2027
rect 2573 2013 2587 2027
rect 2633 2013 2647 2027
rect 2593 1973 2607 1987
rect 2533 1853 2547 1867
rect 2573 1853 2587 1867
rect 2453 1793 2467 1807
rect 2513 1793 2527 1807
rect 2473 1773 2487 1787
rect 2433 1753 2447 1767
rect 2473 1733 2487 1747
rect 2453 1693 2467 1707
rect 2433 1593 2447 1607
rect 2433 1573 2447 1587
rect 2333 1493 2347 1507
rect 2313 1353 2327 1367
rect 2253 1313 2267 1327
rect 2273 1293 2287 1307
rect 2293 1273 2307 1287
rect 2313 1253 2327 1267
rect 2233 1133 2247 1147
rect 2273 1133 2287 1147
rect 2213 1093 2227 1107
rect 2393 1433 2407 1447
rect 2353 1373 2367 1387
rect 2413 1413 2427 1427
rect 2453 1533 2467 1547
rect 2433 1333 2447 1347
rect 2433 1313 2447 1327
rect 2413 1293 2427 1307
rect 2353 1273 2367 1287
rect 2333 1113 2347 1127
rect 2233 1073 2247 1087
rect 2173 1053 2187 1067
rect 2193 1053 2207 1067
rect 1973 753 1987 767
rect 1953 653 1967 667
rect 2013 693 2027 707
rect 1953 613 1967 627
rect 1993 613 2007 627
rect 1993 573 2007 587
rect 1913 393 1927 407
rect 1973 393 1987 407
rect 1733 353 1747 367
rect 1713 313 1727 327
rect 1813 353 1827 367
rect 1853 333 1867 347
rect 1913 333 1927 347
rect 1913 313 1927 327
rect 1833 273 1847 287
rect 1753 213 1767 227
rect 1693 133 1707 147
rect 1733 133 1747 147
rect 1773 133 1787 147
rect 2033 673 2047 687
rect 2053 633 2067 647
rect 2153 793 2167 807
rect 2133 713 2147 727
rect 2113 653 2127 667
rect 2033 453 2047 467
rect 1993 353 2007 367
rect 2013 353 2027 367
rect 1973 333 1987 347
rect 1913 253 1927 267
rect 1933 253 1947 267
rect 1993 253 2007 267
rect 1993 213 2007 227
rect 1933 193 1947 207
rect 1993 193 2007 207
rect 1953 173 1967 187
rect 1973 173 1987 187
rect 2013 173 2027 187
rect 1993 153 2007 167
rect 1873 133 1887 147
rect 1913 133 1927 147
rect 993 93 1007 107
rect 733 73 747 87
rect 873 73 887 87
rect 2073 533 2087 547
rect 2193 893 2207 907
rect 2333 1093 2347 1107
rect 2293 1053 2307 1067
rect 2253 1033 2267 1047
rect 2333 1013 2347 1027
rect 2313 913 2327 927
rect 2313 873 2327 887
rect 2333 873 2347 887
rect 2213 853 2227 867
rect 2273 853 2287 867
rect 2193 813 2207 827
rect 2233 833 2247 847
rect 2613 1873 2627 1887
rect 2573 1793 2587 1807
rect 2593 1793 2607 1807
rect 2673 1993 2687 2007
rect 2713 1933 2727 1947
rect 2673 1813 2687 1827
rect 2713 1793 2727 1807
rect 2653 1773 2667 1787
rect 2533 1733 2547 1747
rect 2513 1693 2527 1707
rect 2573 1753 2587 1767
rect 2553 1633 2567 1647
rect 2553 1593 2567 1607
rect 2513 1553 2527 1567
rect 2493 1493 2507 1507
rect 2533 1493 2547 1507
rect 2473 1353 2487 1367
rect 2573 1573 2587 1587
rect 2553 1433 2567 1447
rect 2633 1753 2647 1767
rect 2693 1753 2707 1767
rect 2613 1713 2627 1727
rect 2633 1713 2647 1727
rect 2653 1613 2667 1627
rect 2653 1593 2667 1607
rect 2753 2133 2767 2147
rect 2813 2273 2827 2287
rect 2813 2213 2827 2227
rect 2873 2253 2887 2267
rect 2833 2193 2847 2207
rect 2913 2253 2927 2267
rect 2893 2173 2907 2187
rect 2853 2153 2867 2167
rect 2873 2153 2887 2167
rect 2793 2113 2807 2127
rect 2853 2113 2867 2127
rect 2753 2093 2767 2107
rect 2793 2093 2807 2107
rect 2753 2073 2767 2087
rect 2833 2073 2847 2087
rect 2973 2393 2987 2407
rect 2973 2353 2987 2367
rect 3013 2313 3027 2327
rect 3093 2433 3107 2447
rect 3013 2273 3027 2287
rect 3053 2273 3067 2287
rect 2953 2233 2967 2247
rect 2933 2113 2947 2127
rect 2913 2093 2927 2107
rect 2973 2153 2987 2167
rect 2973 2113 2987 2127
rect 2953 2073 2967 2087
rect 2773 2053 2787 2067
rect 2773 2033 2787 2047
rect 2853 2053 2867 2067
rect 2853 2033 2867 2047
rect 2893 2033 2907 2047
rect 2813 2013 2827 2027
rect 2793 1993 2807 2007
rect 2753 1953 2767 1967
rect 2773 1953 2787 1967
rect 2773 1893 2787 1907
rect 2813 1973 2827 1987
rect 2833 1853 2847 1867
rect 2793 1833 2807 1847
rect 2773 1813 2787 1827
rect 2993 2093 3007 2107
rect 2933 1973 2947 1987
rect 2973 1993 2987 2007
rect 2993 1893 3007 1907
rect 3033 2253 3047 2267
rect 3053 2193 3067 2207
rect 3113 2213 3127 2227
rect 3073 2173 3087 2187
rect 3093 2173 3107 2187
rect 3033 2093 3047 2107
rect 3073 2093 3087 2107
rect 3033 2053 3047 2067
rect 3053 2053 3067 2067
rect 2993 1873 3007 1887
rect 3013 1873 3027 1887
rect 2853 1833 2867 1847
rect 2773 1793 2787 1807
rect 2833 1813 2847 1827
rect 2873 1813 2887 1827
rect 2893 1813 2907 1827
rect 2933 1833 2947 1847
rect 2973 1833 2987 1847
rect 2733 1733 2747 1747
rect 2753 1733 2767 1747
rect 2713 1693 2727 1707
rect 2793 1773 2807 1787
rect 2833 1713 2847 1727
rect 2873 1713 2887 1727
rect 2753 1673 2767 1687
rect 2773 1673 2787 1687
rect 2733 1653 2747 1667
rect 2713 1633 2727 1647
rect 2633 1573 2647 1587
rect 2653 1553 2667 1567
rect 2593 1533 2607 1547
rect 2613 1533 2627 1547
rect 2633 1513 2647 1527
rect 2593 1433 2607 1447
rect 2573 1373 2587 1387
rect 2613 1373 2627 1387
rect 2533 1353 2547 1367
rect 2533 1313 2547 1327
rect 2573 1313 2587 1327
rect 2493 1293 2507 1307
rect 2453 1273 2467 1287
rect 2473 1273 2487 1287
rect 2373 1253 2387 1267
rect 2433 1253 2447 1267
rect 2473 1253 2487 1267
rect 2373 1173 2387 1187
rect 2453 1113 2467 1127
rect 2593 1293 2607 1307
rect 2553 1273 2567 1287
rect 2513 1233 2527 1247
rect 2613 1233 2627 1247
rect 2533 1133 2547 1147
rect 2413 1093 2427 1107
rect 2393 1073 2407 1087
rect 2433 1073 2447 1087
rect 2413 1053 2427 1067
rect 2453 1053 2467 1067
rect 2373 1033 2387 1047
rect 2393 873 2407 887
rect 2353 853 2367 867
rect 2393 853 2407 867
rect 2373 833 2387 847
rect 2173 673 2187 687
rect 2213 773 2227 787
rect 2253 793 2267 807
rect 2233 713 2247 727
rect 2213 673 2227 687
rect 2153 633 2167 647
rect 2313 813 2327 827
rect 2353 813 2367 827
rect 2293 733 2307 747
rect 2253 633 2267 647
rect 2273 593 2287 607
rect 2293 593 2307 607
rect 2153 533 2167 547
rect 2173 533 2187 547
rect 2133 393 2147 407
rect 2073 373 2087 387
rect 2053 353 2067 367
rect 2053 333 2067 347
rect 2113 353 2127 367
rect 2153 353 2167 367
rect 2193 393 2207 407
rect 2133 333 2147 347
rect 2173 333 2187 347
rect 2253 333 2267 347
rect 2233 293 2247 307
rect 2053 253 2067 267
rect 2153 233 2167 247
rect 2093 173 2107 187
rect 2073 153 2087 167
rect 2053 133 2067 147
rect 2113 153 2127 167
rect 2133 153 2147 167
rect 2013 93 2027 107
rect 2193 173 2207 187
rect 2173 153 2187 167
rect 2253 253 2267 267
rect 2153 133 2167 147
rect 2213 133 2227 147
rect 2133 93 2147 107
rect 1893 73 1907 87
rect 2113 73 2127 87
rect 1233 53 1247 67
rect 2433 1013 2447 1027
rect 2433 833 2447 847
rect 2433 773 2447 787
rect 2413 753 2427 767
rect 2373 693 2387 707
rect 2393 693 2407 707
rect 2433 693 2447 707
rect 2353 653 2367 667
rect 2413 653 2427 667
rect 2393 633 2407 647
rect 2373 613 2387 627
rect 2333 593 2347 607
rect 2393 553 2407 567
rect 2373 453 2387 467
rect 2373 393 2387 407
rect 2313 373 2327 387
rect 2373 333 2387 347
rect 2293 273 2307 287
rect 2353 313 2367 327
rect 2333 253 2347 267
rect 2273 173 2287 187
rect 2353 173 2367 187
rect 2273 133 2287 147
rect 2313 133 2327 147
rect 2613 1093 2627 1107
rect 2593 1073 2607 1087
rect 2553 1013 2567 1027
rect 2513 953 2527 967
rect 2533 953 2547 967
rect 2533 913 2547 927
rect 2853 1653 2867 1667
rect 2793 1613 2807 1627
rect 2813 1613 2827 1627
rect 2673 1533 2687 1547
rect 2753 1533 2767 1547
rect 2733 1513 2747 1527
rect 2713 1453 2727 1467
rect 2653 1313 2667 1327
rect 2653 1273 2667 1287
rect 2693 1273 2707 1287
rect 2773 1513 2787 1527
rect 2793 1453 2807 1467
rect 2833 1593 2847 1607
rect 2933 1793 2947 1807
rect 2913 1713 2927 1727
rect 2893 1633 2907 1647
rect 2873 1613 2887 1627
rect 2893 1533 2907 1547
rect 2853 1513 2867 1527
rect 2893 1513 2907 1527
rect 2833 1433 2847 1447
rect 2813 1373 2827 1387
rect 2873 1493 2887 1507
rect 2873 1433 2887 1447
rect 2853 1373 2867 1387
rect 2773 1353 2787 1367
rect 2833 1353 2847 1367
rect 2753 1333 2767 1347
rect 2773 1293 2787 1307
rect 2733 1253 2747 1267
rect 2713 1233 2727 1247
rect 2793 1233 2807 1247
rect 2833 1253 2847 1267
rect 2693 1213 2707 1227
rect 2813 1213 2827 1227
rect 2853 1233 2867 1247
rect 2673 1173 2687 1187
rect 2773 1173 2787 1187
rect 2793 1173 2807 1187
rect 2733 1153 2747 1167
rect 2713 1133 2727 1147
rect 2713 1093 2727 1107
rect 2633 1053 2647 1067
rect 2693 1073 2707 1087
rect 2653 1013 2667 1027
rect 2633 913 2647 927
rect 2553 873 2567 887
rect 2613 873 2627 887
rect 2493 853 2507 867
rect 2573 853 2587 867
rect 2653 873 2667 887
rect 2513 833 2527 847
rect 2493 813 2507 827
rect 2493 793 2507 807
rect 2513 793 2527 807
rect 2553 813 2567 827
rect 2633 833 2647 847
rect 2593 793 2607 807
rect 2533 733 2547 747
rect 2553 653 2567 667
rect 2753 1113 2767 1127
rect 2833 1153 2847 1167
rect 2833 1113 2847 1127
rect 2753 1073 2767 1087
rect 2733 1053 2747 1067
rect 2713 1013 2727 1027
rect 2973 1773 2987 1787
rect 2973 1693 2987 1707
rect 3053 1933 3067 1947
rect 3033 1833 3047 1847
rect 3073 1853 3087 1867
rect 3013 1813 3027 1827
rect 3193 2553 3207 2567
rect 3253 2673 3267 2687
rect 3293 2673 3307 2687
rect 3173 2513 3187 2527
rect 3213 2513 3227 2527
rect 3173 2473 3187 2487
rect 3173 2193 3187 2207
rect 3153 2153 3167 2167
rect 3173 2133 3187 2147
rect 3113 2093 3127 2107
rect 3133 2093 3147 2107
rect 3113 2073 3127 2087
rect 3153 2073 3167 2087
rect 3113 2033 3127 2047
rect 3193 2013 3207 2027
rect 3273 2633 3287 2647
rect 3293 2593 3307 2607
rect 3393 3013 3407 3027
rect 3413 3013 3427 3027
rect 3353 2993 3367 3007
rect 3433 2993 3447 3007
rect 3333 2973 3347 2987
rect 3373 2973 3387 2987
rect 3353 2953 3367 2967
rect 3333 2813 3347 2827
rect 3333 2753 3347 2767
rect 3353 2733 3367 2747
rect 3413 2953 3427 2967
rect 3393 2753 3407 2767
rect 3593 3413 3607 3427
rect 3533 3213 3547 3227
rect 3513 3053 3527 3067
rect 3573 3273 3587 3287
rect 3573 3233 3587 3247
rect 3693 3513 3707 3527
rect 3753 3533 3767 3547
rect 3793 3613 3807 3627
rect 3633 3473 3647 3487
rect 3713 3493 3727 3507
rect 3753 3493 3767 3507
rect 3773 3493 3787 3507
rect 3693 3473 3707 3487
rect 3633 3453 3647 3467
rect 3673 3453 3687 3467
rect 3613 3273 3627 3287
rect 3613 3253 3627 3267
rect 3593 3213 3607 3227
rect 3513 3033 3527 3047
rect 3553 3033 3567 3047
rect 3473 2993 3487 3007
rect 3533 2993 3547 3007
rect 3513 2973 3527 2987
rect 3553 2973 3567 2987
rect 3493 2793 3507 2807
rect 3333 2693 3347 2707
rect 3313 2553 3327 2567
rect 3333 2553 3347 2567
rect 3253 2473 3267 2487
rect 3253 2353 3267 2367
rect 3333 2313 3347 2327
rect 3293 2293 3307 2307
rect 3273 2253 3287 2267
rect 3233 2233 3247 2247
rect 3253 2233 3267 2247
rect 3293 2153 3307 2167
rect 3233 2033 3247 2047
rect 3153 1973 3167 1987
rect 3173 1933 3187 1947
rect 3133 1913 3147 1927
rect 3153 1913 3167 1927
rect 3133 1833 3147 1847
rect 3153 1813 3167 1827
rect 3133 1793 3147 1807
rect 3013 1773 3027 1787
rect 3053 1773 3067 1787
rect 3093 1773 3107 1787
rect 3153 1773 3167 1787
rect 3053 1753 3067 1767
rect 3113 1753 3127 1767
rect 2933 1673 2947 1687
rect 2993 1673 3007 1687
rect 3033 1653 3047 1667
rect 2933 1613 2947 1627
rect 2953 1593 2967 1607
rect 2933 1493 2947 1507
rect 3073 1713 3087 1727
rect 3133 1713 3147 1727
rect 3113 1613 3127 1627
rect 3133 1613 3147 1627
rect 2993 1553 3007 1567
rect 2973 1513 2987 1527
rect 2953 1453 2967 1467
rect 2933 1433 2947 1447
rect 2913 1313 2927 1327
rect 2973 1433 2987 1447
rect 2973 1333 2987 1347
rect 2973 1293 2987 1307
rect 2973 1273 2987 1287
rect 2933 1233 2947 1247
rect 2893 1173 2907 1187
rect 2933 1153 2947 1167
rect 2933 1113 2947 1127
rect 2853 1053 2867 1067
rect 2813 933 2827 947
rect 2833 933 2847 947
rect 2753 913 2767 927
rect 2753 873 2767 887
rect 2673 853 2687 867
rect 2693 773 2707 787
rect 2673 713 2687 727
rect 2673 693 2687 707
rect 2553 613 2567 627
rect 2473 593 2487 607
rect 2493 533 2507 547
rect 2733 773 2747 787
rect 2713 753 2727 767
rect 2713 733 2727 747
rect 2853 853 2867 867
rect 2793 813 2807 827
rect 2793 793 2807 807
rect 2773 773 2787 787
rect 2753 653 2767 667
rect 2753 633 2767 647
rect 2573 533 2587 547
rect 2593 533 2607 547
rect 2533 513 2547 527
rect 2653 613 2667 627
rect 2693 613 2707 627
rect 2733 613 2747 627
rect 2833 793 2847 807
rect 2793 733 2807 747
rect 2813 733 2827 747
rect 2793 673 2807 687
rect 2813 653 2827 667
rect 2613 513 2627 527
rect 2793 513 2807 527
rect 2453 493 2467 507
rect 2593 493 2607 507
rect 2633 493 2647 507
rect 2433 453 2447 467
rect 2433 433 2447 447
rect 2413 373 2427 387
rect 2413 353 2427 367
rect 2413 253 2427 267
rect 2413 233 2427 247
rect 2413 173 2427 187
rect 2533 373 2547 387
rect 2473 353 2487 367
rect 2513 353 2527 367
rect 2453 333 2467 347
rect 2553 353 2567 367
rect 2753 453 2767 467
rect 2833 633 2847 647
rect 2873 793 2887 807
rect 2913 1073 2927 1087
rect 2953 1073 2967 1087
rect 2933 1033 2947 1047
rect 2913 1013 2927 1027
rect 2873 753 2887 767
rect 2893 753 2907 767
rect 2853 613 2867 627
rect 2953 1013 2967 1027
rect 2933 953 2947 967
rect 2973 933 2987 947
rect 3053 1573 3067 1587
rect 3093 1573 3107 1587
rect 3013 1493 3027 1507
rect 3053 1473 3067 1487
rect 3013 1433 3027 1447
rect 3133 1453 3147 1467
rect 3153 1413 3167 1427
rect 3053 1313 3067 1327
rect 3093 1313 3107 1327
rect 3133 1313 3147 1327
rect 3273 1993 3287 2007
rect 3233 1893 3247 1907
rect 3273 1873 3287 1887
rect 3233 1833 3247 1847
rect 3313 2133 3327 2147
rect 3373 2353 3387 2367
rect 3413 2693 3427 2707
rect 3393 2273 3407 2287
rect 3353 2233 3367 2247
rect 3353 2093 3367 2107
rect 3413 2153 3427 2167
rect 3393 2073 3407 2087
rect 3393 2053 3407 2067
rect 3313 1933 3327 1947
rect 3373 2033 3387 2047
rect 3393 2013 3407 2027
rect 3333 1873 3347 1887
rect 3313 1833 3327 1847
rect 3213 1813 3227 1827
rect 3213 1773 3227 1787
rect 3193 1593 3207 1607
rect 3193 1573 3207 1587
rect 3293 1813 3307 1827
rect 3353 1813 3367 1827
rect 3233 1753 3247 1767
rect 3373 1773 3387 1787
rect 3513 2773 3527 2787
rect 3453 2753 3467 2767
rect 3533 2753 3547 2767
rect 3593 2773 3607 2787
rect 3573 2753 3587 2767
rect 3533 2713 3547 2727
rect 3493 2673 3507 2687
rect 3573 2653 3587 2667
rect 3453 2593 3467 2607
rect 3473 2553 3487 2567
rect 3493 2553 3507 2567
rect 3613 2553 3627 2567
rect 3473 2353 3487 2367
rect 3533 2533 3547 2547
rect 3573 2533 3587 2547
rect 3613 2533 3627 2547
rect 3693 3273 3707 3287
rect 3673 3253 3687 3267
rect 3653 3233 3667 3247
rect 3693 3053 3707 3067
rect 3673 2893 3687 2907
rect 3773 3173 3787 3187
rect 3733 3053 3747 3067
rect 3753 3053 3767 3067
rect 3753 2893 3767 2907
rect 3733 2773 3747 2787
rect 3653 2713 3667 2727
rect 3713 2753 3727 2767
rect 3713 2693 3727 2707
rect 3673 2633 3687 2647
rect 3513 2513 3527 2527
rect 3553 2513 3567 2527
rect 3593 2513 3607 2527
rect 3553 2413 3567 2427
rect 3513 2373 3527 2387
rect 3493 2273 3507 2287
rect 3453 2133 3467 2147
rect 3433 2113 3447 2127
rect 3533 2253 3547 2267
rect 3593 2353 3607 2367
rect 3633 2473 3647 2487
rect 3613 2293 3627 2307
rect 3533 2233 3547 2247
rect 3553 2233 3567 2247
rect 3493 2193 3507 2207
rect 3433 2093 3447 2107
rect 3493 2073 3507 2087
rect 3453 2053 3467 2067
rect 3473 2053 3487 2067
rect 3413 1973 3427 1987
rect 3473 1953 3487 1967
rect 3433 1813 3447 1827
rect 3413 1773 3427 1787
rect 3253 1713 3267 1727
rect 3253 1613 3267 1627
rect 3213 1513 3227 1527
rect 3293 1693 3307 1707
rect 3293 1613 3307 1627
rect 3293 1593 3307 1607
rect 3253 1513 3267 1527
rect 3233 1413 3247 1427
rect 3233 1333 3247 1347
rect 3173 1313 3187 1327
rect 3193 1313 3207 1327
rect 3033 1293 3047 1307
rect 3013 1273 3027 1287
rect 3013 1253 3027 1267
rect 3053 1153 3067 1167
rect 3013 1133 3027 1147
rect 3033 1133 3047 1147
rect 3013 1113 3027 1127
rect 3033 1093 3047 1107
rect 3113 1293 3127 1307
rect 3093 1273 3107 1287
rect 3073 953 3087 967
rect 2953 833 2967 847
rect 2993 913 3007 927
rect 2933 813 2947 827
rect 2973 813 2987 827
rect 2913 733 2927 747
rect 2893 713 2907 727
rect 2933 713 2947 727
rect 3053 933 3067 947
rect 3053 853 3067 867
rect 3013 813 3027 827
rect 2953 693 2967 707
rect 2933 633 2947 647
rect 2893 613 2907 627
rect 2933 613 2947 627
rect 2913 593 2927 607
rect 2953 593 2967 607
rect 2933 573 2947 587
rect 2953 513 2967 527
rect 2893 493 2907 507
rect 2873 453 2887 467
rect 2813 373 2827 387
rect 2833 373 2847 387
rect 2933 433 2947 447
rect 2893 393 2907 407
rect 2913 373 2927 387
rect 3233 1293 3247 1307
rect 3133 1233 3147 1247
rect 3153 1233 3167 1247
rect 3133 1153 3147 1167
rect 3213 1273 3227 1287
rect 3213 1253 3227 1267
rect 3173 1173 3187 1187
rect 3153 1133 3167 1147
rect 3133 1093 3147 1107
rect 3193 1153 3207 1167
rect 3173 1113 3187 1127
rect 3133 1073 3147 1087
rect 3293 1433 3307 1447
rect 3333 1753 3347 1767
rect 3393 1753 3407 1767
rect 3333 1713 3347 1727
rect 3373 1713 3387 1727
rect 3393 1673 3407 1687
rect 3573 2153 3587 2167
rect 3653 2353 3667 2367
rect 3613 2113 3627 2127
rect 3633 2113 3647 2127
rect 3573 2093 3587 2107
rect 3573 2053 3587 2067
rect 3593 2053 3607 2067
rect 3573 1993 3587 2007
rect 3553 1933 3567 1947
rect 3533 1813 3547 1827
rect 3513 1793 3527 1807
rect 3453 1773 3467 1787
rect 3473 1753 3487 1767
rect 3533 1773 3547 1787
rect 3533 1753 3547 1767
rect 3473 1713 3487 1727
rect 3493 1713 3507 1727
rect 3433 1693 3447 1707
rect 3433 1673 3447 1687
rect 3413 1633 3427 1647
rect 3373 1613 3387 1627
rect 3393 1593 3407 1607
rect 3433 1593 3447 1607
rect 3353 1553 3367 1567
rect 3353 1513 3367 1527
rect 3473 1573 3487 1587
rect 3453 1553 3467 1567
rect 3413 1533 3427 1547
rect 3393 1453 3407 1467
rect 3373 1433 3387 1447
rect 3373 1413 3387 1427
rect 3353 1373 3367 1387
rect 3313 1333 3327 1347
rect 3273 1293 3287 1307
rect 3273 1273 3287 1287
rect 3253 1233 3267 1247
rect 3233 1213 3247 1227
rect 3213 1013 3227 1027
rect 3173 953 3187 967
rect 3193 953 3207 967
rect 3193 933 3207 947
rect 3093 913 3107 927
rect 3213 913 3227 927
rect 3193 873 3207 887
rect 3113 833 3127 847
rect 3153 833 3167 847
rect 3193 833 3207 847
rect 3093 813 3107 827
rect 3053 693 3067 707
rect 3033 653 3047 667
rect 2993 633 3007 647
rect 3053 633 3067 647
rect 3013 613 3027 627
rect 3333 1273 3347 1287
rect 3313 1233 3327 1247
rect 3413 1373 3427 1387
rect 3453 1373 3467 1387
rect 3413 1333 3427 1347
rect 3513 1693 3527 1707
rect 3613 1833 3627 1847
rect 3593 1793 3607 1807
rect 3613 1793 3627 1807
rect 3573 1693 3587 1707
rect 3533 1673 3547 1687
rect 3553 1673 3567 1687
rect 3613 1693 3627 1707
rect 3613 1673 3627 1687
rect 3593 1633 3607 1647
rect 3613 1633 3627 1647
rect 3533 1613 3547 1627
rect 3613 1593 3627 1607
rect 3533 1573 3547 1587
rect 3553 1573 3567 1587
rect 3513 1553 3527 1567
rect 3513 1533 3527 1547
rect 3533 1533 3547 1547
rect 3493 1433 3507 1447
rect 3493 1373 3507 1387
rect 3473 1353 3487 1367
rect 3473 1333 3487 1347
rect 3393 1313 3407 1327
rect 3373 1293 3387 1307
rect 3433 1293 3447 1307
rect 3413 1273 3427 1287
rect 3433 1273 3447 1287
rect 3393 1213 3407 1227
rect 3373 1173 3387 1187
rect 3353 1153 3367 1167
rect 3373 1153 3387 1167
rect 3313 1133 3327 1147
rect 3353 1133 3367 1147
rect 3253 1113 3267 1127
rect 3273 1113 3287 1127
rect 3333 1113 3347 1127
rect 3253 1073 3267 1087
rect 3253 1033 3267 1047
rect 3293 1033 3307 1047
rect 3273 993 3287 1007
rect 3233 853 3247 867
rect 3213 813 3227 827
rect 3153 793 3167 807
rect 3173 793 3187 807
rect 3113 753 3127 767
rect 3173 633 3187 647
rect 3073 613 3087 627
rect 3093 613 3107 627
rect 3133 613 3147 627
rect 3013 593 3027 607
rect 2973 453 2987 467
rect 2953 393 2967 407
rect 2673 353 2687 367
rect 2733 353 2747 367
rect 2753 353 2767 367
rect 2793 353 2807 367
rect 2833 353 2847 367
rect 2893 353 2907 367
rect 2933 353 2947 367
rect 2593 333 2607 347
rect 2633 333 2647 347
rect 2493 313 2507 327
rect 2533 313 2547 327
rect 2573 293 2587 307
rect 2473 213 2487 227
rect 2553 213 2567 227
rect 2513 193 2527 207
rect 2473 173 2487 187
rect 2433 153 2447 167
rect 2613 253 2627 267
rect 2653 253 2667 267
rect 2633 213 2647 227
rect 2613 153 2627 167
rect 2713 333 2727 347
rect 2733 253 2747 267
rect 2713 213 2727 227
rect 2673 193 2687 207
rect 2733 153 2747 167
rect 2653 133 2667 147
rect 2693 133 2707 147
rect 2733 133 2747 147
rect 2533 93 2547 107
rect 2633 93 2647 107
rect 2773 333 2787 347
rect 2793 333 2807 347
rect 2793 253 2807 267
rect 2853 333 2867 347
rect 2793 193 2807 207
rect 2873 193 2887 207
rect 2933 193 2947 207
rect 2833 133 2847 147
rect 2913 173 2927 187
rect 2973 373 2987 387
rect 3093 553 3107 567
rect 3073 473 3087 487
rect 3213 753 3227 767
rect 3373 1113 3387 1127
rect 3473 1253 3487 1267
rect 3453 1233 3467 1247
rect 3433 1113 3447 1127
rect 3433 1093 3447 1107
rect 3433 1053 3447 1067
rect 3393 1033 3407 1047
rect 3353 993 3367 1007
rect 3433 993 3447 1007
rect 3353 953 3367 967
rect 3333 913 3347 927
rect 3413 933 3427 947
rect 3393 913 3407 927
rect 3253 753 3267 767
rect 3233 733 3247 747
rect 3233 713 3247 727
rect 3313 813 3327 827
rect 3393 853 3407 867
rect 3373 833 3387 847
rect 3413 833 3427 847
rect 3373 813 3387 827
rect 3333 773 3347 787
rect 3313 753 3327 767
rect 3273 673 3287 687
rect 3233 653 3247 667
rect 3273 633 3287 647
rect 3213 613 3227 627
rect 3253 613 3267 627
rect 3293 613 3307 627
rect 3353 733 3367 747
rect 3333 613 3347 627
rect 3213 593 3227 607
rect 3233 593 3247 607
rect 3313 593 3327 607
rect 3193 573 3207 587
rect 3133 493 3147 507
rect 3133 453 3147 467
rect 3213 453 3227 467
rect 3113 413 3127 427
rect 2993 333 3007 347
rect 2993 313 3007 327
rect 2973 253 2987 267
rect 3053 353 3067 367
rect 3073 353 3087 367
rect 3093 353 3107 367
rect 3093 233 3107 247
rect 3033 173 3047 187
rect 3013 153 3027 167
rect 3053 153 3067 167
rect 3193 413 3207 427
rect 3133 373 3147 387
rect 3133 353 3147 367
rect 3133 233 3147 247
rect 3113 153 3127 167
rect 2993 133 3007 147
rect 3033 133 3047 147
rect 3113 133 3127 147
rect 3173 333 3187 347
rect 3213 313 3227 327
rect 3273 393 3287 407
rect 3293 333 3307 347
rect 3233 293 3247 307
rect 3273 293 3287 307
rect 3233 193 3247 207
rect 3193 153 3207 167
rect 3213 153 3227 167
rect 3253 133 3267 147
rect 3073 73 3087 87
rect 3213 73 3227 87
rect 3393 753 3407 767
rect 3413 733 3427 747
rect 3393 653 3407 667
rect 3473 1173 3487 1187
rect 3533 1433 3547 1447
rect 3533 1333 3547 1347
rect 3533 1293 3547 1307
rect 3613 1533 3627 1547
rect 3573 1513 3587 1527
rect 3613 1473 3627 1487
rect 3593 1433 3607 1447
rect 3573 1353 3587 1367
rect 3593 1333 3607 1347
rect 3553 1233 3567 1247
rect 3593 1233 3607 1247
rect 3513 1213 3527 1227
rect 3553 1213 3567 1227
rect 3593 1213 3607 1227
rect 3513 1173 3527 1187
rect 3493 1113 3507 1127
rect 3493 1073 3507 1087
rect 3533 1073 3547 1087
rect 3453 953 3467 967
rect 3493 913 3507 927
rect 3453 853 3467 867
rect 3473 833 3487 847
rect 3453 813 3467 827
rect 3433 653 3447 667
rect 3393 613 3407 627
rect 3353 593 3367 607
rect 3373 473 3387 487
rect 3393 433 3407 447
rect 3513 733 3527 747
rect 3473 653 3487 667
rect 3453 413 3467 427
rect 3373 373 3387 387
rect 3413 373 3427 387
rect 3353 353 3367 367
rect 3353 313 3367 327
rect 3333 293 3347 307
rect 3313 253 3327 267
rect 3293 233 3307 247
rect 3293 173 3307 187
rect 3413 353 3427 367
rect 3393 293 3407 307
rect 3453 253 3467 267
rect 3433 193 3447 207
rect 3353 153 3367 167
rect 3373 153 3387 167
rect 3413 153 3427 167
rect 3333 133 3347 147
rect 3293 113 3307 127
rect 2753 53 2767 67
rect 3273 53 3287 67
rect 2253 33 2267 47
rect 3573 1113 3587 1127
rect 3573 1073 3587 1087
rect 3653 1913 3667 1927
rect 3693 2593 3707 2607
rect 3753 2613 3767 2627
rect 3713 2513 3727 2527
rect 3813 3533 3827 3547
rect 3833 3493 3847 3507
rect 3813 3393 3827 3407
rect 3873 3713 3887 3727
rect 3973 4193 3987 4207
rect 3993 4193 4007 4207
rect 3953 4153 3967 4167
rect 3933 4133 3947 4147
rect 4093 4233 4107 4247
rect 4033 4173 4047 4187
rect 4033 4033 4047 4047
rect 4153 4253 4167 4267
rect 4113 4173 4127 4187
rect 4093 4153 4107 4167
rect 4073 4093 4087 4107
rect 3993 4013 4007 4027
rect 4033 4013 4047 4027
rect 4053 4013 4067 4027
rect 4013 3993 4027 4007
rect 3953 3973 3967 3987
rect 3973 3973 3987 3987
rect 4073 3973 4087 3987
rect 4013 3933 4027 3947
rect 3913 3693 3927 3707
rect 3873 3633 3887 3647
rect 3893 3593 3907 3607
rect 3993 3713 4007 3727
rect 4093 3953 4107 3967
rect 4133 4093 4147 4107
rect 4153 4093 4167 4107
rect 4313 4533 4327 4547
rect 4253 4493 4267 4507
rect 4233 4473 4247 4487
rect 4293 4473 4307 4487
rect 4273 4453 4287 4467
rect 4353 4473 4367 4487
rect 4453 4693 4467 4707
rect 4573 4713 4587 4727
rect 4513 4693 4527 4707
rect 4533 4693 4547 4707
rect 4493 4673 4507 4687
rect 4433 4653 4447 4667
rect 4433 4613 4447 4627
rect 4393 4453 4407 4467
rect 4413 4453 4427 4467
rect 4273 4433 4287 4447
rect 4353 4433 4367 4447
rect 4213 4413 4227 4427
rect 4193 4213 4207 4227
rect 4213 4193 4227 4207
rect 4253 4173 4267 4187
rect 4233 4153 4247 4167
rect 4253 4133 4267 4147
rect 4233 4113 4247 4127
rect 4233 4093 4247 4107
rect 4173 4053 4187 4067
rect 4153 4013 4167 4027
rect 4133 3953 4147 3967
rect 4113 3913 4127 3927
rect 3973 3693 3987 3707
rect 4033 3693 4047 3707
rect 4013 3593 4027 3607
rect 3933 3553 3947 3567
rect 3973 3533 3987 3547
rect 4133 3773 4147 3787
rect 4113 3753 4127 3767
rect 4113 3713 4127 3727
rect 4093 3693 4107 3707
rect 4073 3673 4087 3687
rect 4093 3673 4107 3687
rect 4093 3633 4107 3647
rect 3873 3453 3887 3467
rect 3953 3453 3967 3467
rect 3993 3513 4007 3527
rect 4033 3513 4047 3527
rect 3913 3393 3927 3407
rect 3973 3393 3987 3407
rect 3833 3213 3847 3227
rect 3813 3053 3827 3067
rect 4113 3573 4127 3587
rect 4133 3533 4147 3547
rect 4073 3473 4087 3487
rect 4133 3473 4147 3487
rect 4193 3993 4207 4007
rect 4173 3953 4187 3967
rect 4213 3933 4227 3947
rect 4293 4213 4307 4227
rect 4633 4793 4647 4807
rect 4793 5273 4807 5287
rect 4733 5173 4747 5187
rect 4733 5153 4747 5167
rect 4753 5093 4767 5107
rect 4713 5053 4727 5067
rect 4693 4933 4707 4947
rect 4773 4973 4787 4987
rect 4733 4933 4747 4947
rect 4713 4893 4727 4907
rect 4713 4793 4727 4807
rect 4673 4693 4687 4707
rect 4633 4673 4647 4687
rect 4593 4633 4607 4647
rect 4693 4653 4707 4667
rect 4653 4613 4667 4627
rect 4553 4553 4567 4567
rect 4613 4553 4627 4567
rect 4593 4493 4607 4507
rect 4513 4373 4527 4387
rect 4313 4193 4327 4207
rect 4353 4193 4367 4207
rect 4393 4193 4407 4207
rect 4373 4173 4387 4187
rect 4333 4153 4347 4167
rect 4393 4153 4407 4167
rect 4293 4113 4307 4127
rect 4293 4073 4307 4087
rect 4273 4013 4287 4027
rect 4333 4053 4347 4067
rect 4293 3993 4307 4007
rect 4253 3973 4267 3987
rect 4273 3973 4287 3987
rect 4313 3933 4327 3947
rect 4373 4013 4387 4027
rect 4353 3993 4367 4007
rect 4393 3993 4407 4007
rect 4353 3973 4367 3987
rect 4333 3873 4347 3887
rect 4333 3853 4347 3867
rect 4233 3833 4247 3847
rect 4273 3833 4287 3847
rect 4193 3733 4207 3747
rect 4233 3733 4247 3747
rect 4173 3693 4187 3707
rect 4233 3693 4247 3707
rect 4253 3693 4267 3707
rect 4293 3693 4307 3707
rect 4213 3653 4227 3667
rect 4393 3953 4407 3967
rect 4373 3873 4387 3887
rect 4393 3773 4407 3787
rect 4693 4293 4707 4307
rect 4613 4273 4627 4287
rect 4653 4273 4667 4287
rect 4613 4253 4627 4267
rect 4513 4193 4527 4207
rect 4573 4193 4587 4207
rect 4493 4173 4507 4187
rect 4593 4173 4607 4187
rect 4453 4153 4467 4167
rect 4473 4153 4487 4167
rect 4433 4113 4447 4127
rect 4433 3973 4447 3987
rect 4533 4093 4547 4107
rect 4633 4053 4647 4067
rect 4613 4033 4627 4047
rect 4633 4033 4647 4047
rect 4453 3933 4467 3947
rect 4573 3993 4587 4007
rect 4553 3973 4567 3987
rect 4493 3933 4507 3947
rect 4513 3933 4527 3947
rect 4473 3893 4487 3907
rect 4433 3733 4447 3747
rect 4373 3713 4387 3727
rect 4393 3693 4407 3707
rect 4353 3653 4367 3667
rect 4233 3633 4247 3647
rect 4313 3633 4327 3647
rect 4333 3633 4347 3647
rect 4373 3633 4387 3647
rect 4173 3613 4187 3627
rect 4273 3573 4287 3587
rect 4173 3553 4187 3567
rect 4333 3593 4347 3607
rect 4393 3613 4407 3627
rect 4453 3693 4467 3707
rect 4453 3613 4467 3627
rect 4413 3533 4427 3547
rect 4193 3493 4207 3507
rect 4293 3493 4307 3507
rect 4333 3493 4347 3507
rect 4353 3473 4367 3487
rect 4433 3473 4447 3487
rect 4153 3433 4167 3447
rect 4273 3433 4287 3447
rect 4173 3333 4187 3347
rect 4133 3213 4147 3227
rect 4113 3153 4127 3167
rect 3873 3113 3887 3127
rect 3993 3073 4007 3087
rect 4113 3013 4127 3027
rect 4113 2973 4127 2987
rect 3833 2893 3847 2907
rect 3913 2893 3927 2907
rect 4033 2873 4047 2887
rect 4073 2873 4087 2887
rect 3813 2673 3827 2687
rect 3793 2653 3807 2667
rect 3853 2633 3867 2647
rect 3693 2473 3707 2487
rect 3773 2473 3787 2487
rect 3693 2453 3707 2467
rect 3713 2453 3727 2467
rect 4073 2793 4087 2807
rect 4153 2873 4167 2887
rect 4053 2773 4067 2787
rect 4053 2653 4067 2667
rect 3933 2433 3947 2447
rect 3973 2433 3987 2447
rect 3733 2373 3747 2387
rect 3853 2353 3867 2367
rect 3733 2313 3747 2327
rect 3793 2313 3807 2327
rect 3813 2313 3827 2327
rect 3753 2293 3767 2307
rect 3733 2253 3747 2267
rect 3713 2233 3727 2247
rect 3713 2173 3727 2187
rect 3693 2153 3707 2167
rect 3673 1853 3687 1867
rect 3833 2293 3847 2307
rect 3913 2273 3927 2287
rect 3953 2273 3967 2287
rect 3833 2213 3847 2227
rect 3813 2153 3827 2167
rect 3773 2133 3787 2147
rect 3733 2113 3747 2127
rect 3773 2093 3787 2107
rect 3813 2093 3827 2107
rect 3793 2073 3807 2087
rect 3773 2053 3787 2067
rect 3753 2033 3767 2047
rect 3733 1993 3747 2007
rect 3733 1893 3747 1907
rect 3653 1813 3667 1827
rect 3693 1813 3707 1827
rect 3713 1813 3727 1827
rect 3693 1793 3707 1807
rect 3833 1893 3847 1907
rect 3893 2253 3907 2267
rect 3933 2253 3947 2267
rect 3873 2233 3887 2247
rect 3913 2213 3927 2227
rect 3953 2233 3967 2247
rect 4033 2353 4047 2367
rect 4013 2333 4027 2347
rect 4013 2273 4027 2287
rect 3993 2253 4007 2267
rect 3973 2213 3987 2227
rect 3933 2173 3947 2187
rect 3953 2173 3967 2187
rect 3893 2033 3907 2047
rect 3893 2013 3907 2027
rect 3873 1933 3887 1947
rect 3833 1873 3847 1887
rect 3853 1873 3867 1887
rect 3793 1833 3807 1847
rect 3873 1853 3887 1867
rect 3873 1793 3887 1807
rect 3693 1753 3707 1767
rect 3673 1733 3687 1747
rect 3653 1713 3667 1727
rect 3653 1693 3667 1707
rect 3653 1593 3667 1607
rect 3753 1773 3767 1787
rect 3853 1773 3867 1787
rect 3733 1753 3747 1767
rect 3773 1753 3787 1767
rect 3713 1733 3727 1747
rect 3733 1713 3747 1727
rect 3693 1553 3707 1567
rect 3733 1673 3747 1687
rect 3813 1733 3827 1747
rect 3833 1713 3847 1727
rect 3813 1693 3827 1707
rect 3773 1653 3787 1667
rect 3793 1653 3807 1667
rect 3753 1633 3767 1647
rect 3773 1633 3787 1647
rect 3793 1613 3807 1627
rect 3833 1653 3847 1667
rect 3993 2153 4007 2167
rect 3973 2133 3987 2147
rect 3973 2073 3987 2087
rect 4093 2773 4107 2787
rect 4073 2573 4087 2587
rect 4073 2513 4087 2527
rect 4053 2293 4067 2307
rect 4053 2273 4067 2287
rect 4193 3253 4207 3267
rect 4233 3253 4247 3267
rect 4233 3153 4247 3167
rect 4213 3053 4227 3067
rect 4253 3053 4267 3067
rect 4213 3013 4227 3027
rect 4173 2773 4187 2787
rect 4173 2753 4187 2767
rect 4113 2733 4127 2747
rect 4133 2653 4147 2667
rect 4253 2913 4267 2927
rect 4233 2793 4247 2807
rect 4233 2773 4247 2787
rect 4233 2713 4247 2727
rect 4213 2673 4227 2687
rect 4193 2633 4207 2647
rect 4193 2593 4207 2607
rect 4173 2573 4187 2587
rect 4253 2613 4267 2627
rect 4293 3233 4307 3247
rect 4433 3233 4447 3247
rect 4593 3913 4607 3927
rect 4533 3773 4547 3787
rect 4513 3713 4527 3727
rect 4593 3673 4607 3687
rect 4573 3653 4587 3667
rect 4553 3633 4567 3647
rect 4493 3513 4507 3527
rect 4513 3493 4527 3507
rect 4593 3513 4607 3527
rect 4493 3473 4507 3487
rect 4593 3353 4607 3367
rect 4673 4233 4687 4247
rect 4673 4193 4687 4207
rect 4653 3973 4667 3987
rect 4633 3913 4647 3927
rect 4693 4073 4707 4087
rect 4713 4053 4727 4067
rect 4693 3913 4707 3927
rect 4673 3713 4687 3727
rect 4613 3273 4627 3287
rect 4653 3493 4667 3507
rect 4773 4673 4787 4687
rect 4773 4453 4787 4467
rect 4753 4433 4767 4447
rect 4993 5393 5007 5407
rect 4913 5373 4927 5387
rect 4873 5193 4887 5207
rect 4813 5153 4827 5167
rect 4873 5173 4887 5187
rect 4913 5173 4927 5187
rect 4853 5153 4867 5167
rect 4893 5153 4907 5167
rect 4833 5133 4847 5147
rect 4833 5093 4847 5107
rect 4893 4993 4907 5007
rect 4913 4973 4927 4987
rect 5213 5413 5227 5427
rect 5153 5373 5167 5387
rect 5093 5333 5107 5347
rect 5113 5333 5127 5347
rect 5053 5213 5067 5227
rect 4953 4993 4967 5007
rect 5033 5133 5047 5147
rect 5033 5113 5047 5127
rect 4973 4973 4987 4987
rect 4993 4973 5007 4987
rect 5013 4973 5027 4987
rect 5013 4953 5027 4967
rect 4953 4933 4967 4947
rect 4993 4933 5007 4947
rect 5193 5213 5207 5227
rect 5173 5173 5187 5187
rect 5133 5113 5147 5127
rect 5153 5113 5167 5127
rect 5293 5433 5307 5447
rect 5413 5453 5427 5467
rect 5473 5453 5487 5467
rect 5533 5453 5547 5467
rect 5593 5453 5607 5467
rect 5353 5433 5367 5447
rect 5373 5433 5387 5447
rect 5453 5433 5467 5447
rect 5273 5413 5287 5427
rect 5253 5373 5267 5387
rect 5413 5413 5427 5427
rect 5273 5193 5287 5207
rect 5353 5193 5367 5207
rect 5393 5173 5407 5187
rect 5073 5053 5087 5067
rect 5153 5053 5167 5067
rect 5193 5053 5207 5067
rect 5073 5033 5087 5047
rect 5093 4993 5107 5007
rect 5113 4973 5127 4987
rect 5133 4973 5147 4987
rect 5053 4833 5067 4847
rect 5113 4833 5127 4847
rect 5013 4773 5027 4787
rect 4993 4713 5007 4727
rect 4833 4693 4847 4707
rect 4913 4693 4927 4707
rect 4933 4693 4947 4707
rect 4953 4693 4967 4707
rect 5013 4693 5027 4707
rect 4813 4653 4827 4667
rect 4833 4633 4847 4647
rect 4873 4633 4887 4647
rect 5013 4673 5027 4687
rect 5053 4673 5067 4687
rect 4973 4653 4987 4667
rect 5033 4653 5047 4667
rect 5073 4653 5087 4667
rect 5093 4633 5107 4647
rect 5133 4773 5147 4787
rect 5133 4713 5147 4727
rect 5013 4613 5027 4627
rect 5073 4613 5087 4627
rect 5113 4613 5127 4627
rect 4853 4393 4867 4407
rect 4813 4373 4827 4387
rect 4793 4293 4807 4307
rect 4913 4293 4927 4307
rect 5033 4513 5047 4527
rect 5013 4413 5027 4427
rect 4793 4193 4807 4207
rect 4933 4193 4947 4207
rect 4773 4173 4787 4187
rect 4933 4153 4947 4167
rect 5053 4453 5067 4467
rect 5053 4193 5067 4207
rect 5033 4133 5047 4147
rect 4893 4093 4907 4107
rect 4793 4073 4807 4087
rect 4753 4053 4767 4067
rect 4753 4013 4767 4027
rect 4913 4073 4927 4087
rect 4753 3933 4767 3947
rect 4993 4053 5007 4067
rect 4873 3773 4887 3787
rect 4913 3773 4927 3787
rect 5113 4593 5127 4607
rect 5093 4573 5107 4587
rect 5193 5033 5207 5047
rect 5233 5033 5247 5047
rect 5213 4953 5227 4967
rect 5153 4673 5167 4687
rect 5153 4633 5167 4647
rect 5133 4513 5147 4527
rect 5133 4493 5147 4507
rect 5113 4453 5127 4467
rect 5193 4913 5207 4927
rect 5193 4653 5207 4667
rect 5173 4493 5187 4507
rect 5193 4473 5207 4487
rect 5093 4433 5107 4447
rect 5173 4433 5187 4447
rect 5133 4373 5147 4387
rect 5093 4213 5107 4227
rect 5113 4193 5127 4207
rect 5153 4313 5167 4327
rect 5173 4253 5187 4267
rect 5153 4233 5167 4247
rect 5153 4093 5167 4107
rect 5133 4073 5147 4087
rect 5113 4053 5127 4067
rect 5073 3973 5087 3987
rect 5053 3933 5067 3947
rect 5033 3813 5047 3827
rect 4913 3753 4927 3767
rect 4933 3753 4947 3767
rect 4993 3753 5007 3767
rect 4793 3713 4807 3727
rect 4893 3693 4907 3707
rect 4733 3613 4747 3627
rect 4833 3533 4847 3547
rect 4873 3393 4887 3407
rect 4713 3353 4727 3367
rect 4673 3333 4687 3347
rect 4633 3233 4647 3247
rect 4413 3193 4427 3207
rect 4353 3073 4367 3087
rect 4313 3053 4327 3067
rect 4293 3033 4307 3047
rect 4373 3033 4387 3047
rect 4333 3013 4347 3027
rect 4293 2653 4307 2667
rect 4613 3193 4627 3207
rect 4653 3133 4667 3147
rect 4453 3113 4467 3127
rect 4493 3113 4507 3127
rect 4513 3033 4527 3047
rect 4533 3033 4547 3047
rect 4473 3013 4487 3027
rect 4433 2993 4447 3007
rect 4413 2973 4427 2987
rect 4613 3033 4627 3047
rect 4593 3013 4607 3027
rect 4593 2993 4607 3007
rect 4333 2713 4347 2727
rect 4553 2853 4567 2867
rect 4673 3053 4687 3067
rect 4593 2713 4607 2727
rect 4513 2673 4527 2687
rect 4413 2653 4427 2667
rect 4433 2653 4447 2667
rect 4273 2593 4287 2607
rect 4313 2593 4327 2607
rect 4273 2573 4287 2587
rect 4373 2573 4387 2587
rect 4313 2553 4327 2567
rect 4353 2553 4367 2567
rect 4253 2533 4267 2547
rect 4393 2553 4407 2567
rect 4473 2633 4487 2647
rect 4433 2553 4447 2567
rect 4553 2613 4567 2627
rect 4633 2693 4647 2707
rect 4493 2533 4507 2547
rect 4533 2513 4547 2527
rect 4333 2473 4347 2487
rect 4413 2473 4427 2487
rect 4493 2473 4507 2487
rect 4293 2433 4307 2447
rect 4193 2393 4207 2407
rect 4173 2293 4187 2307
rect 4133 2273 4147 2287
rect 4133 2253 4147 2267
rect 4093 2173 4107 2187
rect 4113 2173 4127 2187
rect 4113 2133 4127 2147
rect 4073 2113 4087 2127
rect 4313 2193 4327 2207
rect 4493 2453 4507 2467
rect 4413 2433 4427 2447
rect 4353 2193 4367 2207
rect 4213 2173 4227 2187
rect 4333 2173 4347 2187
rect 4173 2113 4187 2127
rect 4153 2093 4167 2107
rect 4133 2073 4147 2087
rect 4013 2033 4027 2047
rect 4033 2033 4047 2047
rect 4093 2033 4107 2047
rect 4133 2033 4147 2047
rect 3993 2013 4007 2027
rect 4013 1973 4027 1987
rect 3993 1913 4007 1927
rect 4013 1913 4027 1927
rect 3973 1853 3987 1867
rect 3953 1813 3967 1827
rect 3993 1813 4007 1827
rect 3913 1793 3927 1807
rect 3973 1793 3987 1807
rect 4013 1793 4027 1807
rect 3893 1773 3907 1787
rect 3993 1773 4007 1787
rect 3953 1753 3967 1767
rect 3993 1753 4007 1767
rect 3933 1733 3947 1747
rect 3873 1633 3887 1647
rect 3893 1633 3907 1647
rect 3853 1613 3867 1627
rect 3893 1593 3907 1607
rect 3733 1553 3747 1567
rect 3753 1553 3767 1567
rect 3793 1553 3807 1567
rect 3673 1533 3687 1547
rect 3713 1533 3727 1547
rect 3773 1533 3787 1547
rect 3813 1533 3827 1547
rect 3653 1393 3667 1407
rect 3713 1413 3727 1427
rect 3633 1333 3647 1347
rect 3633 1313 3647 1327
rect 3633 1273 3647 1287
rect 3693 1373 3707 1387
rect 3673 1333 3687 1347
rect 3633 1213 3647 1227
rect 3613 1173 3627 1187
rect 3673 1133 3687 1147
rect 3633 1113 3647 1127
rect 3673 1113 3687 1127
rect 3613 1093 3627 1107
rect 3633 1053 3647 1067
rect 3593 1013 3607 1027
rect 3613 913 3627 927
rect 3573 833 3587 847
rect 3873 1573 3887 1587
rect 3873 1513 3887 1527
rect 3833 1493 3847 1507
rect 3853 1493 3867 1507
rect 3813 1473 3827 1487
rect 3813 1453 3827 1467
rect 3833 1453 3847 1467
rect 3813 1413 3827 1427
rect 3773 1373 3787 1387
rect 3733 1333 3747 1347
rect 3773 1333 3787 1347
rect 3713 1313 3727 1327
rect 3753 1313 3767 1327
rect 3793 1313 3807 1327
rect 3753 1293 3767 1307
rect 3713 1273 3727 1287
rect 3693 1053 3707 1067
rect 3653 1013 3667 1027
rect 3713 993 3727 1007
rect 3813 1233 3827 1247
rect 3793 1213 3807 1227
rect 3813 1213 3827 1227
rect 3773 1153 3787 1167
rect 3813 1173 3827 1187
rect 3873 1353 3887 1367
rect 3873 1333 3887 1347
rect 3933 1633 3947 1647
rect 3973 1633 3987 1647
rect 4053 1933 4067 1947
rect 4113 1853 4127 1867
rect 4093 1833 4107 1847
rect 4073 1813 4087 1827
rect 4253 2153 4267 2167
rect 4313 2073 4327 2087
rect 4393 2173 4407 2187
rect 4193 2053 4207 2067
rect 4233 2053 4247 2067
rect 4173 2033 4187 2047
rect 4273 2013 4287 2027
rect 4373 2053 4387 2067
rect 4173 1993 4187 2007
rect 4333 1993 4347 2007
rect 4013 1593 4027 1607
rect 3933 1473 3947 1487
rect 4013 1553 4027 1567
rect 3993 1513 4007 1527
rect 3973 1453 3987 1467
rect 4053 1613 4067 1627
rect 4113 1733 4127 1747
rect 4133 1733 4147 1747
rect 4113 1633 4127 1647
rect 4253 1973 4267 1987
rect 4473 2293 4487 2307
rect 4433 2273 4447 2287
rect 4513 2333 4527 2347
rect 4733 3233 4747 3247
rect 4913 3373 4927 3387
rect 4813 3233 4827 3247
rect 4833 3233 4847 3247
rect 4873 3233 4887 3247
rect 4793 3213 4807 3227
rect 4793 3133 4807 3147
rect 4973 3733 4987 3747
rect 4953 3693 4967 3707
rect 5013 3693 5027 3707
rect 5013 3673 5027 3687
rect 4993 3633 5007 3647
rect 5133 3993 5147 4007
rect 5113 3933 5127 3947
rect 5093 3773 5107 3787
rect 5193 4193 5207 4207
rect 5193 4093 5207 4107
rect 5173 4053 5187 4067
rect 5193 4033 5207 4047
rect 5173 3993 5187 4007
rect 5113 3693 5127 3707
rect 5153 3693 5167 3707
rect 5053 3673 5067 3687
rect 5033 3653 5047 3667
rect 5093 3513 5107 3527
rect 5193 3733 5207 3747
rect 5193 3713 5207 3727
rect 5513 5413 5527 5427
rect 5473 5373 5487 5387
rect 5613 5393 5627 5407
rect 5533 5213 5547 5227
rect 5573 5213 5587 5227
rect 5413 5133 5427 5147
rect 5473 5133 5487 5147
rect 5653 5153 5667 5167
rect 5693 5153 5707 5167
rect 5493 5113 5507 5127
rect 5513 5113 5527 5127
rect 5573 5113 5587 5127
rect 5373 5033 5387 5047
rect 5533 4993 5547 5007
rect 5673 4993 5687 5007
rect 5273 4973 5287 4987
rect 5453 4913 5467 4927
rect 5233 4713 5247 4727
rect 5513 4833 5527 4847
rect 5273 4713 5287 4727
rect 5433 4713 5447 4727
rect 5233 4593 5247 4607
rect 5233 4513 5247 4527
rect 5413 4593 5427 4607
rect 5473 4593 5487 4607
rect 5273 4493 5287 4507
rect 5313 4493 5327 4507
rect 5253 4453 5267 4467
rect 5353 4453 5367 4467
rect 5273 4393 5287 4407
rect 5253 4373 5267 4387
rect 5253 4353 5267 4367
rect 5233 4173 5247 4187
rect 5273 4213 5287 4227
rect 5253 4113 5267 4127
rect 5253 4093 5267 4107
rect 5233 4073 5247 4087
rect 5493 4493 5507 4507
rect 5433 4413 5447 4427
rect 5453 4413 5467 4427
rect 5413 4193 5427 4207
rect 5413 4113 5427 4127
rect 5333 4093 5347 4107
rect 5413 4093 5427 4107
rect 5313 4073 5327 4087
rect 5273 3993 5287 4007
rect 5233 3773 5247 3787
rect 5293 3973 5307 3987
rect 5293 3953 5307 3967
rect 5253 3753 5267 3767
rect 5273 3753 5287 3767
rect 5233 3713 5247 3727
rect 5193 3533 5207 3547
rect 5033 3473 5047 3487
rect 5073 3473 5087 3487
rect 5013 3373 5027 3387
rect 4973 3293 4987 3307
rect 4933 3253 4947 3267
rect 4853 3193 4867 3207
rect 4853 3173 4867 3187
rect 4833 3053 4847 3067
rect 4893 3053 4907 3067
rect 4873 3033 4887 3047
rect 4733 3013 4747 3027
rect 4753 2993 4767 3007
rect 4853 3013 4867 3027
rect 4893 3013 4907 3027
rect 4833 2993 4847 3007
rect 4793 2973 4807 2987
rect 4793 2953 4807 2967
rect 4693 2793 4707 2807
rect 4713 2773 4727 2787
rect 4753 2773 4767 2787
rect 4773 2773 4787 2787
rect 4693 2753 4707 2767
rect 4733 2733 4747 2747
rect 4733 2713 4747 2727
rect 4673 2633 4687 2647
rect 4593 2533 4607 2547
rect 4573 2453 4587 2467
rect 4673 2473 4687 2487
rect 4553 2413 4567 2427
rect 4533 2293 4547 2307
rect 4553 2293 4567 2307
rect 4513 2133 4527 2147
rect 4573 2273 4587 2287
rect 4593 2273 4607 2287
rect 4713 2513 4727 2527
rect 4893 2973 4907 2987
rect 4933 3213 4947 3227
rect 4973 3213 4987 3227
rect 5133 3393 5147 3407
rect 5133 3353 5147 3367
rect 5213 3473 5227 3487
rect 5173 3353 5187 3367
rect 4993 3193 5007 3207
rect 4933 3053 4947 3067
rect 5013 3033 5027 3047
rect 4973 3013 4987 3027
rect 5093 3193 5107 3207
rect 5133 3233 5147 3247
rect 5113 3133 5127 3147
rect 5153 3133 5167 3147
rect 5073 3053 5087 3067
rect 5113 3013 5127 3027
rect 4913 2913 4927 2927
rect 4913 2853 4927 2867
rect 4893 2833 4907 2847
rect 4853 2793 4867 2807
rect 4813 2733 4827 2747
rect 4833 2733 4847 2747
rect 4793 2653 4807 2667
rect 4773 2633 4787 2647
rect 5033 2993 5047 3007
rect 5093 2993 5107 3007
rect 5133 2993 5147 3007
rect 5093 2973 5107 2987
rect 5053 2953 5067 2967
rect 4953 2833 4967 2847
rect 4953 2753 4967 2767
rect 4893 2733 4907 2747
rect 4913 2733 4927 2747
rect 5033 2773 5047 2787
rect 5153 2773 5167 2787
rect 5113 2753 5127 2767
rect 5213 3273 5227 3287
rect 5193 3013 5207 3027
rect 5173 2753 5187 2767
rect 5013 2733 5027 2747
rect 4993 2713 5007 2727
rect 4773 2613 4787 2627
rect 4873 2613 4887 2627
rect 4753 2533 4767 2547
rect 4733 2433 4747 2447
rect 4873 2573 4887 2587
rect 4853 2513 4867 2527
rect 4773 2353 4787 2367
rect 5093 2733 5107 2747
rect 5053 2593 5067 2607
rect 5033 2553 5047 2567
rect 5053 2553 5067 2567
rect 5073 2553 5087 2567
rect 5033 2533 5047 2547
rect 5013 2493 5027 2507
rect 4893 2433 4907 2447
rect 5013 2433 5027 2447
rect 4853 2313 4867 2327
rect 4693 2293 4707 2307
rect 4613 2133 4627 2147
rect 4553 2113 4567 2127
rect 4473 2093 4487 2107
rect 4493 2093 4507 2107
rect 4533 2093 4547 2107
rect 4453 2073 4467 2087
rect 4413 1973 4427 1987
rect 4273 1873 4287 1887
rect 4233 1833 4247 1847
rect 4293 1853 4307 1867
rect 4353 1853 4367 1867
rect 4193 1813 4207 1827
rect 4273 1813 4287 1827
rect 4193 1753 4207 1767
rect 4313 1833 4327 1847
rect 4293 1773 4307 1787
rect 4393 1833 4407 1847
rect 4493 2033 4507 2047
rect 4573 2073 4587 2087
rect 4433 1833 4447 1847
rect 4453 1833 4467 1847
rect 4333 1773 4347 1787
rect 4413 1773 4427 1787
rect 4473 1813 4487 1827
rect 4473 1773 4487 1787
rect 4313 1753 4327 1767
rect 4273 1733 4287 1747
rect 4353 1733 4367 1747
rect 4193 1713 4207 1727
rect 4233 1693 4247 1707
rect 4293 1633 4307 1647
rect 4133 1613 4147 1627
rect 4173 1613 4187 1627
rect 4193 1613 4207 1627
rect 4233 1613 4247 1627
rect 4093 1593 4107 1607
rect 4073 1573 4087 1587
rect 4093 1573 4107 1587
rect 4153 1573 4167 1587
rect 4173 1573 4187 1587
rect 4073 1553 4087 1567
rect 4033 1493 4047 1507
rect 4113 1493 4127 1507
rect 4113 1473 4127 1487
rect 4013 1433 4027 1447
rect 4033 1393 4047 1407
rect 4093 1393 4107 1407
rect 3813 1093 3827 1107
rect 3773 1053 3787 1067
rect 3793 1053 3807 1067
rect 3753 1033 3767 1047
rect 3753 1013 3767 1027
rect 3773 953 3787 967
rect 3753 933 3767 947
rect 3733 913 3747 927
rect 3713 873 3727 887
rect 3633 853 3647 867
rect 3673 833 3687 847
rect 3733 833 3747 847
rect 3553 793 3567 807
rect 3593 793 3607 807
rect 3653 693 3667 707
rect 3573 653 3587 667
rect 3493 613 3507 627
rect 3513 593 3527 607
rect 3493 573 3507 587
rect 3513 553 3527 567
rect 3553 513 3567 527
rect 3533 433 3547 447
rect 3653 633 3667 647
rect 3593 613 3607 627
rect 3633 613 3647 627
rect 3613 593 3627 607
rect 3653 573 3667 587
rect 3593 553 3607 567
rect 3593 533 3607 547
rect 3653 533 3667 547
rect 3633 473 3647 487
rect 3593 373 3607 387
rect 3613 333 3627 347
rect 3573 273 3587 287
rect 3533 253 3547 267
rect 3513 173 3527 187
rect 3553 173 3567 187
rect 3513 153 3527 167
rect 3593 193 3607 207
rect 3573 153 3587 167
rect 3573 113 3587 127
rect 3573 93 3587 107
rect 3653 353 3667 367
rect 3693 813 3707 827
rect 3753 813 3767 827
rect 3693 673 3707 687
rect 3713 673 3727 687
rect 3693 633 3707 647
rect 3693 393 3707 407
rect 3673 333 3687 347
rect 3633 293 3647 307
rect 3653 153 3667 167
rect 3653 133 3667 147
rect 3633 113 3647 127
rect 3693 113 3707 127
rect 3673 93 3687 107
rect 3553 73 3567 87
rect 3593 73 3607 87
rect 3493 33 3507 47
rect 3473 13 3487 27
rect 3593 33 3607 47
rect 3913 1273 3927 1287
rect 3993 1313 4007 1327
rect 3933 1233 3947 1247
rect 3973 1193 3987 1207
rect 3933 1173 3947 1187
rect 4013 1253 4027 1267
rect 3993 1153 4007 1167
rect 3893 1113 3907 1127
rect 3873 1073 3887 1087
rect 3833 953 3847 967
rect 3893 993 3907 1007
rect 3873 893 3887 907
rect 3873 873 3887 887
rect 3813 833 3827 847
rect 3793 693 3807 707
rect 3873 733 3887 747
rect 3733 593 3747 607
rect 3753 573 3767 587
rect 3773 553 3787 567
rect 3733 513 3747 527
rect 3753 513 3767 527
rect 3853 653 3867 667
rect 3993 1133 4007 1147
rect 3953 1053 3967 1067
rect 3953 1033 3967 1047
rect 4173 1553 4187 1567
rect 4153 1373 4167 1387
rect 4193 1493 4207 1507
rect 4173 1353 4187 1367
rect 4113 1333 4127 1347
rect 4133 1313 4147 1327
rect 4053 1253 4067 1267
rect 4033 1153 4047 1167
rect 4053 1153 4067 1167
rect 4033 1133 4047 1147
rect 4113 1293 4127 1307
rect 4133 1293 4147 1307
rect 4253 1593 4267 1607
rect 4273 1593 4287 1607
rect 4233 1513 4247 1527
rect 4233 1473 4247 1487
rect 4253 1413 4267 1427
rect 4213 1373 4227 1387
rect 4233 1373 4247 1387
rect 4413 1753 4427 1767
rect 4373 1633 4387 1647
rect 4353 1593 4367 1607
rect 4393 1613 4407 1627
rect 4313 1553 4327 1567
rect 4313 1353 4327 1367
rect 4233 1333 4247 1347
rect 4273 1333 4287 1347
rect 4173 1313 4187 1327
rect 4213 1313 4227 1327
rect 4233 1313 4247 1327
rect 4273 1313 4287 1327
rect 4313 1313 4327 1327
rect 4153 1253 4167 1267
rect 4233 1233 4247 1247
rect 4133 1213 4147 1227
rect 4093 1173 4107 1187
rect 4133 1153 4147 1167
rect 4213 1153 4227 1167
rect 4193 1133 4207 1147
rect 4153 1113 4167 1127
rect 4033 1073 4047 1087
rect 3973 933 3987 947
rect 4013 933 4027 947
rect 3993 873 4007 887
rect 4113 1093 4127 1107
rect 4293 1293 4307 1307
rect 4313 1273 4327 1287
rect 4233 1133 4247 1147
rect 4253 1133 4267 1147
rect 4173 1073 4187 1087
rect 4193 1073 4207 1087
rect 4053 1013 4067 1027
rect 4073 1013 4087 1027
rect 4073 953 4087 967
rect 4113 933 4127 947
rect 4093 873 4107 887
rect 3913 813 3927 827
rect 3953 833 3967 847
rect 3993 813 4007 827
rect 4033 813 4047 827
rect 3953 793 3967 807
rect 3973 793 3987 807
rect 3913 753 3927 767
rect 3933 753 3947 767
rect 3953 753 3967 767
rect 3893 673 3907 687
rect 3853 633 3867 647
rect 3873 633 3887 647
rect 3833 613 3847 627
rect 3893 573 3907 587
rect 3953 673 3967 687
rect 3933 653 3947 667
rect 4033 733 4047 747
rect 3993 653 4007 667
rect 3933 593 3947 607
rect 3973 573 3987 587
rect 4013 573 4027 587
rect 3913 493 3927 507
rect 3753 473 3767 487
rect 3793 473 3807 487
rect 3733 353 3747 367
rect 4193 913 4207 927
rect 4173 873 4187 887
rect 4193 853 4207 867
rect 4213 833 4227 847
rect 4133 813 4147 827
rect 4193 813 4207 827
rect 4173 793 4187 807
rect 4113 733 4127 747
rect 4073 693 4087 707
rect 4273 1113 4287 1127
rect 4253 1073 4267 1087
rect 4273 1053 4287 1067
rect 4253 933 4267 947
rect 4233 793 4247 807
rect 4213 653 4227 667
rect 4193 633 4207 647
rect 4233 633 4247 647
rect 4073 613 4087 627
rect 4133 613 4147 627
rect 4173 613 4187 627
rect 4093 593 4107 607
rect 4173 593 4187 607
rect 4053 573 4067 587
rect 4213 573 4227 587
rect 4233 553 4247 567
rect 4293 953 4307 967
rect 4313 933 4327 947
rect 4373 1573 4387 1587
rect 4353 1553 4367 1567
rect 4373 1553 4387 1567
rect 4493 1753 4507 1767
rect 4513 1733 4527 1747
rect 4553 1953 4567 1967
rect 4593 1953 4607 1967
rect 4673 2093 4687 2107
rect 4653 2073 4667 2087
rect 4813 2173 4827 2187
rect 4793 2133 4807 2147
rect 4773 2113 4787 2127
rect 4733 2093 4747 2107
rect 4753 2053 4767 2067
rect 4653 2033 4667 2047
rect 4713 2033 4727 2047
rect 4633 2013 4647 2027
rect 4613 1873 4627 1887
rect 4593 1813 4607 1827
rect 4753 1993 4767 2007
rect 4733 1933 4747 1947
rect 4673 1913 4687 1927
rect 4653 1893 4667 1907
rect 4593 1793 4607 1807
rect 4553 1733 4567 1747
rect 4473 1653 4487 1667
rect 4453 1613 4467 1627
rect 4473 1593 4487 1607
rect 4453 1573 4467 1587
rect 4353 1313 4367 1327
rect 4353 1293 4367 1307
rect 4413 1493 4427 1507
rect 4393 1353 4407 1367
rect 4533 1573 4547 1587
rect 4493 1513 4507 1527
rect 4593 1733 4607 1747
rect 4713 1833 4727 1847
rect 4693 1813 4707 1827
rect 4673 1793 4687 1807
rect 4633 1733 4647 1747
rect 4653 1733 4667 1747
rect 4613 1653 4627 1667
rect 4613 1633 4627 1647
rect 4673 1673 4687 1687
rect 4693 1673 4707 1687
rect 4673 1653 4687 1667
rect 4573 1573 4587 1587
rect 4473 1493 4487 1507
rect 4553 1493 4567 1507
rect 4433 1393 4447 1407
rect 4453 1393 4467 1407
rect 4413 1333 4427 1347
rect 4433 1313 4447 1327
rect 4413 1293 4427 1307
rect 4453 1293 4467 1307
rect 4393 1273 4407 1287
rect 4433 1273 4447 1287
rect 4453 1273 4467 1287
rect 4393 1253 4407 1267
rect 4433 1233 4447 1247
rect 4413 1153 4427 1167
rect 4373 1113 4387 1127
rect 4353 1033 4367 1047
rect 4353 993 4367 1007
rect 4433 993 4447 1007
rect 4333 873 4347 887
rect 4293 833 4307 847
rect 4333 813 4347 827
rect 4313 793 4327 807
rect 4293 673 4307 687
rect 4293 653 4307 667
rect 4333 633 4347 647
rect 4273 613 4287 627
rect 4433 933 4447 947
rect 4393 813 4407 827
rect 4393 793 4407 807
rect 4373 753 4387 767
rect 4373 733 4387 747
rect 4353 593 4367 607
rect 4313 493 4327 507
rect 4033 433 4047 447
rect 4133 433 4147 447
rect 4013 393 4027 407
rect 4073 393 4087 407
rect 4013 353 4027 367
rect 3913 313 3927 327
rect 3753 193 3767 207
rect 3733 173 3747 187
rect 3853 173 3867 187
rect 3773 153 3787 167
rect 3893 153 3907 167
rect 3793 113 3807 127
rect 4133 353 4147 367
rect 4213 313 4227 327
rect 4033 293 4047 307
rect 4373 453 4387 467
rect 4493 1393 4507 1407
rect 4493 1373 4507 1387
rect 4513 1333 4527 1347
rect 4533 1313 4547 1327
rect 4653 1593 4667 1607
rect 4593 1513 4607 1527
rect 4593 1493 4607 1507
rect 4593 1273 4607 1287
rect 4633 1273 4647 1287
rect 4653 1253 4667 1267
rect 4573 1233 4587 1247
rect 4613 1233 4627 1247
rect 4513 1213 4527 1227
rect 4513 1193 4527 1207
rect 4493 1093 4507 1107
rect 4733 1713 4747 1727
rect 4773 1853 4787 1867
rect 4833 2073 4847 2087
rect 4873 2233 4887 2247
rect 4853 1973 4867 1987
rect 4833 1953 4847 1967
rect 4813 1833 4827 1847
rect 4793 1813 4807 1827
rect 4853 1813 4867 1827
rect 4793 1793 4807 1807
rect 4773 1773 4787 1787
rect 4793 1673 4807 1687
rect 4753 1633 4767 1647
rect 4793 1633 4807 1647
rect 4713 1613 4727 1627
rect 4753 1593 4767 1607
rect 4713 1553 4727 1567
rect 4773 1553 4787 1567
rect 4713 1533 4727 1547
rect 4733 1533 4747 1547
rect 4693 1493 4707 1507
rect 4713 1493 4727 1507
rect 4713 1473 4727 1487
rect 4753 1333 4767 1347
rect 4733 1293 4747 1307
rect 4853 1673 4867 1687
rect 4933 2393 4947 2407
rect 4913 2353 4927 2367
rect 4893 2173 4907 2187
rect 4913 2133 4927 2147
rect 4913 2113 4927 2127
rect 4893 2093 4907 2107
rect 4893 1893 4907 1907
rect 4893 1853 4907 1867
rect 4953 2273 4967 2287
rect 5013 2233 5027 2247
rect 5173 2713 5187 2727
rect 5253 3513 5267 3527
rect 5253 3473 5267 3487
rect 5253 3433 5267 3447
rect 5393 4053 5407 4067
rect 5353 4033 5367 4047
rect 5373 4013 5387 4027
rect 5673 4973 5687 4987
rect 5713 4973 5727 4987
rect 5553 4933 5567 4947
rect 5533 4713 5547 4727
rect 5693 4953 5707 4967
rect 5613 4893 5627 4907
rect 5693 4893 5707 4907
rect 5653 4833 5667 4847
rect 5533 4653 5547 4667
rect 5613 4673 5627 4687
rect 5653 4673 5667 4687
rect 5553 4573 5567 4587
rect 5593 4493 5607 4507
rect 5533 4473 5547 4487
rect 5513 4353 5527 4367
rect 5513 4313 5527 4327
rect 5633 4633 5647 4647
rect 5673 4633 5687 4647
rect 5573 4433 5587 4447
rect 5613 4413 5627 4427
rect 5493 4113 5507 4127
rect 5453 3993 5467 4007
rect 5533 4053 5547 4067
rect 5513 3993 5527 4007
rect 5433 3973 5447 3987
rect 5473 3973 5487 3987
rect 5413 3953 5427 3967
rect 5333 3913 5347 3927
rect 5313 3813 5327 3827
rect 5593 4233 5607 4247
rect 5573 4213 5587 4227
rect 5553 4033 5567 4047
rect 5573 4033 5587 4047
rect 5693 4413 5707 4427
rect 5733 4933 5747 4947
rect 5753 4673 5767 4687
rect 5733 4653 5747 4667
rect 5733 4293 5747 4307
rect 5653 4213 5667 4227
rect 5613 4033 5627 4047
rect 5593 4013 5607 4027
rect 5633 4013 5647 4027
rect 5613 3993 5627 4007
rect 5593 3933 5607 3947
rect 5673 4053 5687 4067
rect 5673 4033 5687 4047
rect 5453 3633 5467 3647
rect 5533 3533 5547 3547
rect 5313 3493 5327 3507
rect 5353 3493 5367 3507
rect 5293 3433 5307 3447
rect 5273 3393 5287 3407
rect 5613 3753 5627 3767
rect 5573 3713 5587 3727
rect 5613 3393 5627 3407
rect 5493 3333 5507 3347
rect 5553 3333 5567 3347
rect 5473 3113 5487 3127
rect 5653 3853 5667 3867
rect 5653 3533 5667 3547
rect 5653 3493 5667 3507
rect 5653 3453 5667 3467
rect 5653 3393 5667 3407
rect 5633 3293 5647 3307
rect 5613 3273 5627 3287
rect 5453 3053 5467 3067
rect 5573 2973 5587 2987
rect 5233 2733 5247 2747
rect 5253 2733 5267 2747
rect 5293 2733 5307 2747
rect 5273 2573 5287 2587
rect 5133 2513 5147 2527
rect 5253 2553 5267 2567
rect 5233 2533 5247 2547
rect 5473 2693 5487 2707
rect 5393 2613 5407 2627
rect 5353 2553 5367 2567
rect 5253 2513 5267 2527
rect 5293 2513 5307 2527
rect 5473 2593 5487 2607
rect 5433 2573 5447 2587
rect 5393 2533 5407 2547
rect 5373 2513 5387 2527
rect 5413 2513 5427 2527
rect 5133 2473 5147 2487
rect 5193 2473 5207 2487
rect 5133 2373 5147 2387
rect 5073 2273 5087 2287
rect 5113 2273 5127 2287
rect 5053 2253 5067 2267
rect 5033 2133 5047 2147
rect 5093 2233 5107 2247
rect 5073 2213 5087 2227
rect 5073 2133 5087 2147
rect 5033 2113 5047 2127
rect 5053 2113 5067 2127
rect 4933 1993 4947 2007
rect 4933 1873 4947 1887
rect 4953 1873 4967 1887
rect 4933 1833 4947 1847
rect 4913 1813 4927 1827
rect 4993 2073 5007 2087
rect 4973 1833 4987 1847
rect 5073 2053 5087 2067
rect 5013 2033 5027 2047
rect 5053 2033 5067 2047
rect 5233 2353 5247 2367
rect 5213 2293 5227 2307
rect 5173 2233 5187 2247
rect 5153 2213 5167 2227
rect 5133 2193 5147 2207
rect 5213 2233 5227 2247
rect 5133 2173 5147 2187
rect 5193 2173 5207 2187
rect 5113 2153 5127 2167
rect 5113 2093 5127 2107
rect 5173 2113 5187 2127
rect 5153 2073 5167 2087
rect 5113 2033 5127 2047
rect 5093 1953 5107 1967
rect 5073 1893 5087 1907
rect 5053 1853 5067 1867
rect 5033 1833 5047 1847
rect 4913 1733 4927 1747
rect 4893 1693 4907 1707
rect 4893 1673 4907 1687
rect 4873 1633 4887 1647
rect 4813 1593 4827 1607
rect 4853 1593 4867 1607
rect 4833 1573 4847 1587
rect 4833 1473 4847 1487
rect 4793 1313 4807 1327
rect 4773 1293 4787 1307
rect 4693 1273 4707 1287
rect 4753 1273 4767 1287
rect 4693 1213 4707 1227
rect 4673 1173 4687 1187
rect 4533 1133 4547 1147
rect 4573 1133 4587 1147
rect 4653 1133 4667 1147
rect 4493 1053 4507 1067
rect 4553 1053 4567 1067
rect 4493 973 4507 987
rect 4473 833 4487 847
rect 4613 1093 4627 1107
rect 4593 1073 4607 1087
rect 4633 1073 4647 1087
rect 4673 1073 4687 1087
rect 4673 1053 4687 1067
rect 4593 973 4607 987
rect 4533 853 4547 867
rect 4573 833 4587 847
rect 4653 933 4667 947
rect 4613 853 4627 867
rect 4673 853 4687 867
rect 4633 833 4647 847
rect 4513 813 4527 827
rect 4593 813 4607 827
rect 4633 813 4647 827
rect 4493 793 4507 807
rect 4553 793 4567 807
rect 4573 753 4587 767
rect 4453 733 4467 747
rect 4493 673 4507 687
rect 4473 653 4487 667
rect 4413 633 4427 647
rect 4433 633 4447 647
rect 4453 593 4467 607
rect 4533 653 4547 667
rect 4513 633 4527 647
rect 4493 573 4507 587
rect 4613 693 4627 707
rect 4593 633 4607 647
rect 4673 753 4687 767
rect 4553 573 4567 587
rect 4593 573 4607 587
rect 4653 573 4667 587
rect 4533 533 4547 547
rect 4633 493 4647 507
rect 4393 433 4407 447
rect 4413 393 4427 407
rect 4553 393 4567 407
rect 4393 233 4407 247
rect 4193 173 4207 187
rect 3933 113 3947 127
rect 3833 93 3847 107
rect 4493 353 4507 367
rect 4433 213 4447 227
rect 4373 173 4387 187
rect 4413 173 4427 187
rect 4473 173 4487 187
rect 4313 153 4327 167
rect 4553 233 4567 247
rect 4533 173 4547 187
rect 4573 173 4587 187
rect 4513 153 4527 167
rect 4613 153 4627 167
rect 4673 453 4687 467
rect 4853 1313 4867 1327
rect 4833 1273 4847 1287
rect 4833 1253 4847 1267
rect 4813 1193 4827 1207
rect 4813 1173 4827 1187
rect 4773 1133 4787 1147
rect 4773 1093 4787 1107
rect 4753 1073 4767 1087
rect 4713 933 4727 947
rect 4833 913 4847 927
rect 4813 873 4827 887
rect 4953 1773 4967 1787
rect 4933 1713 4947 1727
rect 4993 1813 5007 1827
rect 4973 1673 4987 1687
rect 4953 1653 4967 1667
rect 4933 1613 4947 1627
rect 4953 1613 4967 1627
rect 4913 1533 4927 1547
rect 4893 1513 4907 1527
rect 5093 1833 5107 1847
rect 5053 1793 5067 1807
rect 5073 1793 5087 1807
rect 5013 1733 5027 1747
rect 5053 1713 5067 1727
rect 5013 1653 5027 1667
rect 5033 1653 5047 1667
rect 5353 2333 5367 2347
rect 5333 2313 5347 2327
rect 5293 2293 5307 2307
rect 5473 2513 5487 2527
rect 5473 2333 5487 2347
rect 5593 2913 5607 2927
rect 5633 2913 5647 2927
rect 5573 2713 5587 2727
rect 5533 2533 5547 2547
rect 5553 2513 5567 2527
rect 5573 2493 5587 2507
rect 5513 2473 5527 2487
rect 5613 2733 5627 2747
rect 5653 2713 5667 2727
rect 5633 2573 5647 2587
rect 5613 2513 5627 2527
rect 5593 2453 5607 2467
rect 5653 2533 5667 2547
rect 5653 2493 5667 2507
rect 5513 2353 5527 2367
rect 5373 2293 5387 2307
rect 5413 2293 5427 2307
rect 5453 2293 5467 2307
rect 5433 2273 5447 2287
rect 5293 2233 5307 2247
rect 5253 2173 5267 2187
rect 5213 2093 5227 2107
rect 5193 2073 5207 2087
rect 5253 2073 5267 2087
rect 5233 2053 5247 2067
rect 5273 2053 5287 2067
rect 5193 2013 5207 2027
rect 5253 1973 5267 1987
rect 5213 1913 5227 1927
rect 5173 1873 5187 1887
rect 5173 1853 5187 1867
rect 5113 1793 5127 1807
rect 5113 1773 5127 1787
rect 5153 1753 5167 1767
rect 5133 1733 5147 1747
rect 5113 1693 5127 1707
rect 5193 1613 5207 1627
rect 5073 1593 5087 1607
rect 5113 1593 5127 1607
rect 5193 1593 5207 1607
rect 5093 1573 5107 1587
rect 5133 1573 5147 1587
rect 5173 1573 5187 1587
rect 5073 1533 5087 1547
rect 4993 1413 5007 1427
rect 4993 1393 5007 1407
rect 4893 1353 4907 1367
rect 4913 1333 4927 1347
rect 4973 1313 4987 1327
rect 4893 1293 4907 1307
rect 4933 1293 4947 1307
rect 4953 1293 4967 1307
rect 4873 1273 4887 1287
rect 4973 1273 4987 1287
rect 4873 1153 4887 1167
rect 4873 1133 4887 1147
rect 4913 1133 4927 1147
rect 4953 1133 4967 1147
rect 4933 1113 4947 1127
rect 4893 1033 4907 1047
rect 4913 913 4927 927
rect 4713 853 4727 867
rect 4733 813 4747 827
rect 4853 853 4867 867
rect 4793 813 4807 827
rect 4713 793 4727 807
rect 4773 793 4787 807
rect 4773 773 4787 787
rect 4793 773 4807 787
rect 4853 753 4867 767
rect 4733 693 4747 707
rect 4833 693 4847 707
rect 4793 673 4807 687
rect 4713 613 4727 627
rect 4833 613 4847 627
rect 4733 453 4747 467
rect 4773 453 4787 467
rect 4713 373 4727 387
rect 4813 373 4827 387
rect 4673 353 4687 367
rect 4733 353 4747 367
rect 4793 293 4807 307
rect 4713 273 4727 287
rect 4693 213 4707 227
rect 4653 173 4667 187
rect 4673 153 4687 167
rect 4413 133 4427 147
rect 4453 133 4467 147
rect 4493 133 4507 147
rect 4413 113 4427 127
rect 4753 153 4767 167
rect 4793 133 4807 147
rect 4713 113 4727 127
rect 4893 873 4907 887
rect 4873 613 4887 627
rect 4873 513 4887 527
rect 4873 353 4887 367
rect 4853 333 4867 347
rect 4873 313 4887 327
rect 4973 1093 4987 1107
rect 4953 873 4967 887
rect 4953 853 4967 867
rect 4933 773 4947 787
rect 4933 633 4947 647
rect 4913 593 4927 607
rect 4913 413 4927 427
rect 4893 293 4907 307
rect 4833 273 4847 287
rect 4853 153 4867 167
rect 4953 533 4967 547
rect 5013 1313 5027 1327
rect 5073 1313 5087 1327
rect 5053 1293 5067 1307
rect 5093 1293 5107 1307
rect 5033 1273 5047 1287
rect 5073 1233 5087 1247
rect 5013 1213 5027 1227
rect 5033 1213 5047 1227
rect 5013 1133 5027 1147
rect 5053 1153 5067 1167
rect 4993 1073 5007 1087
rect 5093 1153 5107 1167
rect 5193 1333 5207 1347
rect 5133 1293 5147 1307
rect 5113 1133 5127 1147
rect 5173 1213 5187 1227
rect 5153 1193 5167 1207
rect 5153 1153 5167 1167
rect 5113 1113 5127 1127
rect 5173 1133 5187 1147
rect 5233 1813 5247 1827
rect 5273 1793 5287 1807
rect 5273 1773 5287 1787
rect 5253 1713 5267 1727
rect 5233 1673 5247 1687
rect 5413 2213 5427 2227
rect 5413 2193 5427 2207
rect 5453 2193 5467 2207
rect 5373 2113 5387 2127
rect 5313 2073 5327 2087
rect 5353 2053 5367 2067
rect 5333 2033 5347 2047
rect 5533 2313 5547 2327
rect 5493 2293 5507 2307
rect 5513 2293 5527 2307
rect 5573 2293 5587 2307
rect 5533 2273 5547 2287
rect 5513 2253 5527 2267
rect 5493 2233 5507 2247
rect 5513 2233 5527 2247
rect 5493 2213 5507 2227
rect 5413 2073 5427 2087
rect 5433 2053 5447 2067
rect 5393 1993 5407 2007
rect 5413 1993 5427 2007
rect 5313 1893 5327 1907
rect 5373 1893 5387 1907
rect 5473 2133 5487 2147
rect 5473 2093 5487 2107
rect 5533 2193 5547 2207
rect 5613 2273 5627 2287
rect 5573 2213 5587 2227
rect 5633 2253 5647 2267
rect 5633 2233 5647 2247
rect 5613 2213 5627 2227
rect 5593 2193 5607 2207
rect 5613 2193 5627 2207
rect 5553 2173 5567 2187
rect 5553 2133 5567 2147
rect 5493 2053 5507 2067
rect 5473 2033 5487 2047
rect 5513 1993 5527 2007
rect 5493 1973 5507 1987
rect 5473 1933 5487 1947
rect 5453 1913 5467 1927
rect 5573 2113 5587 2127
rect 5553 2073 5567 2087
rect 5553 2033 5567 2047
rect 5593 1993 5607 2007
rect 5553 1973 5567 1987
rect 5533 1893 5547 1907
rect 5533 1833 5547 1847
rect 5393 1793 5407 1807
rect 5393 1733 5407 1747
rect 5353 1713 5367 1727
rect 5373 1713 5387 1727
rect 5293 1613 5307 1627
rect 5333 1613 5347 1627
rect 5353 1613 5367 1627
rect 5433 1693 5447 1707
rect 5453 1693 5467 1707
rect 5393 1653 5407 1667
rect 5313 1593 5327 1607
rect 5253 1573 5267 1587
rect 5293 1573 5307 1587
rect 5253 1533 5267 1547
rect 5253 1353 5267 1367
rect 5233 1293 5247 1307
rect 5213 1153 5227 1167
rect 5093 1073 5107 1087
rect 4993 953 5007 967
rect 5073 953 5087 967
rect 5033 913 5047 927
rect 5013 893 5027 907
rect 5013 753 5027 767
rect 5193 1073 5207 1087
rect 5313 1273 5327 1287
rect 5313 1253 5327 1267
rect 5353 1593 5367 1607
rect 5393 1593 5407 1607
rect 5393 1553 5407 1567
rect 5373 1513 5387 1527
rect 5433 1553 5447 1567
rect 5413 1333 5427 1347
rect 5393 1273 5407 1287
rect 5433 1273 5447 1287
rect 5333 1233 5347 1247
rect 5413 1233 5427 1247
rect 5293 1213 5307 1227
rect 5493 1673 5507 1687
rect 5493 1553 5507 1567
rect 5473 1453 5487 1467
rect 5473 1413 5487 1427
rect 5453 1193 5467 1207
rect 5453 1173 5467 1187
rect 5253 1153 5267 1167
rect 5233 1113 5247 1127
rect 5213 1013 5227 1027
rect 5233 853 5247 867
rect 5173 833 5187 847
rect 5213 833 5227 847
rect 5053 813 5067 827
rect 5053 793 5067 807
rect 5033 653 5047 667
rect 5073 773 5087 787
rect 5093 753 5107 767
rect 5153 753 5167 767
rect 5173 753 5187 767
rect 5073 673 5087 687
rect 5113 673 5127 687
rect 5133 673 5147 687
rect 5093 613 5107 627
rect 5153 653 5167 667
rect 4993 593 5007 607
rect 5113 593 5127 607
rect 5013 533 5027 547
rect 4973 353 4987 367
rect 4973 293 4987 307
rect 4893 133 4907 147
rect 4933 133 4947 147
rect 4833 113 4847 127
rect 4913 113 4927 127
rect 5053 353 5067 367
rect 5273 1093 5287 1107
rect 5593 1953 5607 1967
rect 5573 1893 5587 1907
rect 5573 1833 5587 1847
rect 5553 1693 5567 1707
rect 5593 1793 5607 1807
rect 5573 1633 5587 1647
rect 5573 1613 5587 1627
rect 5553 1573 5567 1587
rect 5533 1553 5547 1567
rect 5713 4153 5727 4167
rect 5693 3513 5707 3527
rect 5693 3293 5707 3307
rect 5693 3273 5707 3287
rect 5733 3853 5747 3867
rect 5733 3713 5747 3727
rect 5733 3493 5747 3507
rect 5733 3353 5747 3367
rect 5713 2973 5727 2987
rect 5713 2933 5727 2947
rect 5693 2733 5707 2747
rect 5713 2593 5727 2607
rect 5693 2553 5707 2567
rect 5713 2533 5727 2547
rect 5693 2513 5707 2527
rect 5673 2433 5687 2447
rect 5673 2253 5687 2267
rect 5653 2093 5667 2107
rect 5713 2473 5727 2487
rect 5713 2453 5727 2467
rect 5693 2193 5707 2207
rect 5693 2153 5707 2167
rect 5653 2073 5667 2087
rect 5693 2033 5707 2047
rect 5673 2013 5687 2027
rect 5653 1793 5667 1807
rect 5633 1713 5647 1727
rect 5693 1933 5707 1947
rect 5673 1673 5687 1687
rect 5693 1613 5707 1627
rect 5613 1573 5627 1587
rect 5653 1573 5667 1587
rect 5693 1573 5707 1587
rect 5633 1553 5647 1567
rect 5673 1553 5687 1567
rect 5513 1493 5527 1507
rect 5593 1493 5607 1507
rect 5613 1473 5627 1487
rect 5513 1313 5527 1327
rect 5533 1193 5547 1207
rect 5553 1093 5567 1107
rect 5693 1353 5707 1367
rect 5653 1333 5667 1347
rect 5693 1333 5707 1347
rect 5593 1293 5607 1307
rect 5673 1293 5687 1307
rect 5633 1253 5647 1267
rect 5633 1113 5647 1127
rect 5473 1073 5487 1087
rect 5613 1073 5627 1087
rect 5253 833 5267 847
rect 5233 793 5247 807
rect 5253 753 5267 767
rect 5193 653 5207 667
rect 5333 833 5347 847
rect 5313 813 5327 827
rect 5213 633 5227 647
rect 5253 633 5267 647
rect 5193 613 5207 627
rect 5153 473 5167 487
rect 5193 473 5207 487
rect 5153 433 5167 447
rect 5073 313 5087 327
rect 5053 293 5067 307
rect 5033 113 5047 127
rect 5073 113 5087 127
rect 4693 93 4707 107
rect 4733 93 4747 107
rect 4813 93 4827 107
rect 4913 93 4927 107
rect 5133 333 5147 347
rect 5113 153 5127 167
rect 5533 833 5547 847
rect 5593 833 5607 847
rect 5733 1553 5747 1567
rect 5733 1353 5747 1367
rect 5733 1313 5747 1327
rect 5733 1293 5747 1307
rect 5753 1213 5767 1227
rect 5713 1113 5727 1127
rect 5653 1093 5667 1107
rect 5373 813 5387 827
rect 5353 753 5367 767
rect 5333 673 5347 687
rect 5373 673 5387 687
rect 5313 613 5327 627
rect 5353 613 5367 627
rect 5453 813 5467 827
rect 5493 813 5507 827
rect 5433 793 5447 807
rect 5473 773 5487 787
rect 5413 693 5427 707
rect 5533 693 5547 707
rect 5633 693 5647 707
rect 5433 673 5447 687
rect 5453 653 5467 667
rect 5513 653 5527 667
rect 5393 593 5407 607
rect 5573 633 5587 647
rect 5693 1093 5707 1107
rect 5693 1073 5707 1087
rect 5673 853 5687 867
rect 5673 833 5687 847
rect 5613 393 5627 407
rect 5613 373 5627 387
rect 5693 373 5707 387
rect 5273 353 5287 367
rect 5313 353 5327 367
rect 5573 353 5587 367
rect 5253 173 5267 187
rect 5133 113 5147 127
rect 5113 93 5127 107
rect 5173 93 5187 107
rect 5453 313 5467 327
rect 5493 173 5507 187
rect 5613 133 5627 147
rect 5733 353 5747 367
rect 5733 133 5747 147
rect 5653 113 5667 127
rect 5693 113 5707 127
rect 5093 53 5107 67
rect 5233 53 5247 67
rect 4213 33 4227 47
rect 3633 13 3647 27
rect 3713 13 3727 27
rect 3833 13 3847 27
<< metal3 >>
rect 2547 5536 2813 5544
rect 2427 5516 2773 5524
rect 3147 5516 3313 5524
rect 1227 5476 1613 5484
rect 1627 5476 1833 5484
rect 2967 5476 3013 5484
rect 3027 5476 3353 5484
rect 3407 5476 3493 5484
rect 5267 5476 5313 5484
rect 87 5456 153 5464
rect 207 5456 253 5464
rect 287 5456 513 5464
rect 807 5456 873 5464
rect 887 5456 913 5464
rect 1267 5456 1713 5464
rect 1747 5456 1973 5464
rect 2287 5456 2813 5464
rect 2827 5456 2973 5464
rect 3187 5456 3233 5464
rect 3427 5456 3593 5464
rect 3607 5456 3733 5464
rect 4627 5456 5033 5464
rect 5047 5456 5264 5464
rect 67 5436 933 5444
rect 1307 5436 1333 5444
rect 1507 5436 1573 5444
rect 2207 5436 2313 5444
rect 2327 5436 2473 5444
rect 3247 5436 3613 5444
rect 4027 5436 4093 5444
rect 4147 5436 4253 5444
rect 4307 5436 4353 5444
rect 4527 5436 4753 5444
rect 4767 5436 4893 5444
rect 4967 5436 5173 5444
rect 5207 5436 5233 5444
rect 5256 5444 5264 5456
rect 5287 5456 5413 5464
rect 5487 5456 5533 5464
rect 5547 5456 5593 5464
rect 5256 5436 5293 5444
rect 5387 5436 5453 5444
rect 707 5416 813 5424
rect 936 5424 944 5433
rect 867 5416 944 5424
rect 1436 5424 1444 5433
rect 1187 5416 1244 5424
rect 1236 5407 1244 5416
rect 1316 5416 1633 5424
rect 1316 5407 1324 5416
rect 1847 5416 2233 5424
rect 2787 5416 2913 5424
rect 3027 5416 3273 5424
rect 3696 5424 3704 5433
rect 3487 5416 3833 5424
rect 3856 5416 3913 5424
rect 3856 5407 3864 5416
rect 4127 5416 4213 5424
rect 4227 5416 4313 5424
rect 4407 5416 4433 5424
rect 4467 5416 4493 5424
rect 4667 5416 4693 5424
rect 4807 5416 4873 5424
rect 4956 5424 4964 5433
rect 4956 5416 5013 5424
rect 5147 5416 5213 5424
rect 5227 5416 5273 5424
rect 5356 5424 5364 5433
rect 5356 5416 5413 5424
rect 5427 5416 5513 5424
rect 167 5396 213 5404
rect 847 5396 973 5404
rect 1047 5396 1093 5404
rect 1107 5396 1153 5404
rect 1367 5396 1453 5404
rect 1987 5396 2173 5404
rect 2187 5396 2613 5404
rect 2847 5396 2893 5404
rect 2907 5396 2993 5404
rect 3087 5396 3153 5404
rect 3387 5396 3453 5404
rect 3647 5396 3853 5404
rect 4076 5404 4084 5413
rect 4076 5396 4193 5404
rect 4287 5396 4713 5404
rect 4727 5396 4993 5404
rect 5007 5396 5613 5404
rect 67 5376 93 5384
rect 107 5376 1013 5384
rect 1407 5376 1773 5384
rect 1827 5376 2333 5384
rect 2987 5376 3193 5384
rect 3207 5376 3293 5384
rect 3527 5376 3613 5384
rect 3627 5376 3773 5384
rect 3787 5376 3993 5384
rect 4236 5384 4244 5393
rect 4227 5376 4244 5384
rect 4327 5376 4473 5384
rect 4927 5376 5153 5384
rect 5267 5376 5473 5384
rect 187 5356 1353 5364
rect 3047 5356 3093 5364
rect 3307 5356 3553 5364
rect 3687 5356 3713 5364
rect 4007 5356 4413 5364
rect 4447 5356 4593 5364
rect 3087 5336 3273 5344
rect 4207 5336 4453 5344
rect 4467 5336 4813 5344
rect 4827 5336 5093 5344
rect 5107 5336 5113 5344
rect 367 5316 453 5324
rect 3327 5316 4693 5324
rect 1767 5276 2753 5284
rect 2767 5276 4793 5284
rect 1147 5256 1513 5264
rect 1527 5256 1573 5264
rect 1587 5256 1853 5264
rect 1867 5256 2273 5264
rect 2327 5216 3073 5224
rect 3087 5216 3433 5224
rect 4307 5216 5053 5224
rect 5067 5216 5193 5224
rect 5207 5216 5533 5224
rect 5547 5216 5573 5224
rect 2767 5196 2833 5204
rect 2847 5196 3013 5204
rect 3407 5196 3524 5204
rect 207 5176 273 5184
rect 947 5176 973 5184
rect 1007 5176 1073 5184
rect 1447 5176 1493 5184
rect 1507 5176 1813 5184
rect 2607 5176 2693 5184
rect 3027 5176 3393 5184
rect 3407 5176 3473 5184
rect 316 5164 324 5173
rect 87 5156 324 5164
rect 447 5156 493 5164
rect 887 5156 893 5164
rect 907 5156 1013 5164
rect 1067 5156 1093 5164
rect 1167 5156 1253 5164
rect 1307 5156 1413 5164
rect 1487 5156 1873 5164
rect 1887 5156 2293 5164
rect 2727 5156 2773 5164
rect 3247 5156 3353 5164
rect 3456 5156 3493 5164
rect 347 5136 393 5144
rect 947 5136 1033 5144
rect 1287 5136 1333 5144
rect 1787 5136 1973 5144
rect 2747 5136 2873 5144
rect 2887 5136 3053 5144
rect 3067 5136 3093 5144
rect 3456 5144 3464 5156
rect 3387 5136 3464 5144
rect 3516 5144 3524 5196
rect 3847 5196 4013 5204
rect 4527 5196 4873 5204
rect 5287 5196 5353 5204
rect 3827 5176 3893 5184
rect 3947 5176 4053 5184
rect 4387 5176 4413 5184
rect 4627 5176 4733 5184
rect 4887 5176 4913 5184
rect 5187 5176 5393 5184
rect 3587 5156 3653 5164
rect 3707 5156 3993 5164
rect 4176 5164 4184 5173
rect 4176 5156 4393 5164
rect 4407 5156 4453 5164
rect 4747 5156 4813 5164
rect 4867 5156 4893 5164
rect 5667 5156 5693 5164
rect 3487 5136 3524 5144
rect 3547 5136 3633 5144
rect 3687 5136 3753 5144
rect 3867 5136 3973 5144
rect 4027 5136 4053 5144
rect 4556 5144 4564 5153
rect 4527 5136 4564 5144
rect 4847 5136 5033 5144
rect 5427 5136 5473 5144
rect 47 5116 133 5124
rect 147 5116 173 5124
rect 307 5116 353 5124
rect 787 5116 953 5124
rect 967 5116 1153 5124
rect 1367 5116 1593 5124
rect 2187 5116 2393 5124
rect 2447 5116 2993 5124
rect 3007 5116 3053 5124
rect 3167 5116 3213 5124
rect 3567 5116 3593 5124
rect 3687 5116 3713 5124
rect 3747 5116 3793 5124
rect 4027 5116 4113 5124
rect 4167 5116 4173 5124
rect 4187 5116 4213 5124
rect 4367 5116 4393 5124
rect 4487 5116 4673 5124
rect 4687 5116 5033 5124
rect 5147 5116 5153 5124
rect 5167 5116 5493 5124
rect 5527 5116 5573 5124
rect 1247 5096 1453 5104
rect 2387 5096 3333 5104
rect 3467 5096 3673 5104
rect 3887 5096 4293 5104
rect 4307 5096 4333 5104
rect 4527 5096 4553 5104
rect 4587 5096 4753 5104
rect 4767 5096 4833 5104
rect 127 5076 153 5084
rect 167 5076 833 5084
rect 2027 5076 2453 5084
rect 2907 5076 3113 5084
rect 527 5056 613 5064
rect 1827 5056 1873 5064
rect 1907 5056 2033 5064
rect 3127 5056 3573 5064
rect 3967 5056 4373 5064
rect 4387 5056 4713 5064
rect 4727 5056 5073 5064
rect 5167 5056 5193 5064
rect 207 5036 373 5044
rect 807 5036 1193 5044
rect 1207 5036 1773 5044
rect 1867 5036 1973 5044
rect 2547 5036 2713 5044
rect 2747 5036 2813 5044
rect 4287 5036 4353 5044
rect 5087 5036 5193 5044
rect 5247 5036 5373 5044
rect 387 5016 793 5024
rect 1607 5016 1633 5024
rect 1647 5016 1953 5024
rect 2167 5016 2653 5024
rect 2687 5016 2793 5024
rect 3207 5016 3513 5024
rect 3787 5016 4273 5024
rect 4287 5016 4293 5024
rect 4307 5016 4533 5024
rect 627 4996 993 5004
rect 1027 4996 1653 5004
rect 1667 4996 2153 5004
rect 2227 4996 2313 5004
rect 2467 4996 2933 5004
rect 3027 4996 3093 5004
rect 3107 4996 3173 5004
rect 3407 4996 3433 5004
rect 3767 4996 3913 5004
rect 4907 4996 4953 5004
rect 4967 4996 5093 5004
rect 5547 4996 5673 5004
rect 407 4976 493 4984
rect 507 4976 793 4984
rect 987 4976 1004 4984
rect 547 4956 653 4964
rect 707 4956 733 4964
rect 996 4964 1004 4976
rect 1067 4976 1373 4984
rect 1947 4976 2053 4984
rect 2147 4976 2293 4984
rect 2307 4976 2493 4984
rect 2667 4976 3113 4984
rect 3367 4976 3444 4984
rect 996 4956 1093 4964
rect 1587 4956 1613 4964
rect 1847 4956 2213 4964
rect 2227 4956 2253 4964
rect 2627 4956 2724 4964
rect 727 4936 853 4944
rect 967 4936 993 4944
rect 1807 4936 1913 4944
rect 2347 4936 2413 4944
rect 467 4916 773 4924
rect 1067 4916 1233 4924
rect 1547 4916 1813 4924
rect 2567 4916 2653 4924
rect 2716 4924 2724 4956
rect 2967 4956 3033 4964
rect 3436 4964 3444 4976
rect 3587 4976 3853 4984
rect 3927 4976 4033 4984
rect 4047 4976 4053 4984
rect 4147 4976 4413 4984
rect 4507 4976 4533 4984
rect 4787 4976 4913 4984
rect 4927 4976 4973 4984
rect 5027 4976 5113 4984
rect 5147 4976 5273 4984
rect 5687 4976 5713 4984
rect 3436 4956 3973 4964
rect 3996 4956 4033 4964
rect 2787 4936 2893 4944
rect 3187 4936 3233 4944
rect 3347 4936 3393 4944
rect 3416 4944 3424 4953
rect 3416 4936 3433 4944
rect 3627 4936 3744 4944
rect 3736 4927 3744 4936
rect 3807 4936 3853 4944
rect 2716 4916 2813 4924
rect 3267 4916 3293 4924
rect 3487 4916 3593 4924
rect 3996 4924 4004 4956
rect 4127 4956 4433 4964
rect 4447 4956 4633 4964
rect 4996 4964 5004 4973
rect 4996 4956 5013 4964
rect 5227 4956 5693 4964
rect 4096 4944 4104 4953
rect 4096 4936 4224 4944
rect 4216 4927 4224 4936
rect 4247 4936 4573 4944
rect 4707 4936 4733 4944
rect 4967 4936 4993 4944
rect 5567 4936 5733 4944
rect 3847 4916 4004 4924
rect 4087 4916 4133 4924
rect 4467 4916 4513 4924
rect 4527 4916 4633 4924
rect 5207 4916 5453 4924
rect 747 4896 833 4904
rect 1007 4896 1753 4904
rect 1767 4896 1973 4904
rect 1987 4896 2013 4904
rect 3147 4896 3333 4904
rect 3347 4896 3373 4904
rect 3647 4896 4073 4904
rect 4327 4896 4353 4904
rect 4416 4904 4424 4913
rect 4416 4896 4593 4904
rect 4607 4896 4713 4904
rect 5627 4896 5693 4904
rect 807 4876 1033 4884
rect 1047 4876 1393 4884
rect 1407 4876 1933 4884
rect 2647 4876 3893 4884
rect 3556 4867 3564 4876
rect 3367 4836 3673 4844
rect 3887 4836 4313 4844
rect 4387 4836 5053 4844
rect 5067 4836 5113 4844
rect 5527 4836 5653 4844
rect 1127 4796 1473 4804
rect 4647 4796 4713 4804
rect 207 4776 393 4784
rect 767 4776 1053 4784
rect 1267 4776 2093 4784
rect 2107 4776 2533 4784
rect 5027 4776 5133 4784
rect 47 4756 233 4764
rect 247 4756 473 4764
rect 487 4756 1393 4764
rect 1447 4756 2173 4764
rect 3027 4756 3313 4764
rect 1147 4736 1193 4744
rect 1207 4736 1913 4744
rect 1927 4736 2113 4744
rect 2907 4736 3013 4744
rect 3207 4736 3693 4744
rect 3707 4736 3733 4744
rect 4216 4736 4233 4744
rect 4247 4736 4253 4744
rect 107 4716 173 4724
rect 187 4716 813 4724
rect 967 4716 1253 4724
rect 1767 4716 1793 4724
rect 2007 4716 2093 4724
rect 2107 4716 2253 4724
rect 2487 4716 2624 4724
rect 2616 4707 2624 4716
rect 2927 4716 2973 4724
rect 2987 4716 2993 4724
rect 3107 4716 3213 4724
rect 3227 4716 3424 4724
rect 67 4696 104 4704
rect 56 4676 73 4684
rect 56 4644 64 4676
rect 96 4684 104 4696
rect 567 4696 653 4704
rect 667 4696 853 4704
rect 927 4696 953 4704
rect 1407 4696 1453 4704
rect 2067 4696 2133 4704
rect 2247 4696 2473 4704
rect 2547 4696 2604 4704
rect 96 4676 633 4684
rect 807 4676 833 4684
rect 847 4676 1113 4684
rect 1347 4676 1493 4684
rect 1527 4676 1793 4684
rect 1827 4676 1873 4684
rect 1887 4676 2153 4684
rect 2167 4676 2193 4684
rect 2207 4676 2293 4684
rect 2596 4684 2604 4696
rect 2627 4696 2793 4704
rect 2836 4696 2853 4704
rect 2596 4676 2613 4684
rect 2647 4676 2673 4684
rect 2747 4676 2773 4684
rect 87 4656 113 4664
rect 127 4656 273 4664
rect 867 4656 913 4664
rect 987 4656 1073 4664
rect 1107 4656 1173 4664
rect 1227 4656 1313 4664
rect 1467 4656 1593 4664
rect 2047 4656 2073 4664
rect 2347 4656 2433 4664
rect 2567 4656 2753 4664
rect 2836 4664 2844 4696
rect 3067 4696 3073 4704
rect 3087 4696 3133 4704
rect 3267 4696 3293 4704
rect 2867 4676 2933 4684
rect 2956 4684 2964 4693
rect 3416 4687 3424 4716
rect 3647 4716 3833 4724
rect 3616 4704 3624 4713
rect 3616 4696 3653 4704
rect 2956 4676 3033 4684
rect 2956 4667 2964 4676
rect 3436 4676 3573 4684
rect 2836 4656 2913 4664
rect 2987 4656 3193 4664
rect 3207 4656 3233 4664
rect 3436 4664 3444 4676
rect 3587 4676 3673 4684
rect 3736 4684 3744 4716
rect 3847 4716 3893 4724
rect 3947 4716 3973 4724
rect 4067 4716 4493 4724
rect 4507 4716 4573 4724
rect 5007 4716 5133 4724
rect 5247 4716 5273 4724
rect 5447 4716 5533 4724
rect 3927 4696 4013 4704
rect 4047 4696 4113 4704
rect 4156 4696 4313 4704
rect 3727 4676 3744 4684
rect 3756 4684 3764 4693
rect 4156 4687 4164 4696
rect 4467 4696 4513 4704
rect 4547 4696 4673 4704
rect 4847 4696 4913 4704
rect 4927 4696 4933 4704
rect 4967 4696 5013 4704
rect 3756 4676 3813 4684
rect 4007 4676 4053 4684
rect 4207 4676 4233 4684
rect 4507 4676 4633 4684
rect 4696 4676 4773 4684
rect 4696 4667 4704 4676
rect 4956 4684 4964 4693
rect 4816 4676 4964 4684
rect 4816 4667 4824 4676
rect 5027 4676 5053 4684
rect 5167 4676 5613 4684
rect 5667 4676 5753 4684
rect 3407 4656 3453 4664
rect 3547 4656 3633 4664
rect 3707 4656 3953 4664
rect 3967 4656 4373 4664
rect 4447 4656 4693 4664
rect 4987 4656 5033 4664
rect 5087 4656 5193 4664
rect 5547 4656 5733 4664
rect 56 4636 133 4644
rect 167 4636 393 4644
rect 907 4636 1233 4644
rect 1487 4636 2133 4644
rect 2147 4636 2213 4644
rect 2227 4636 2273 4644
rect 2287 4636 2393 4644
rect 2407 4636 2553 4644
rect 2587 4636 3333 4644
rect 3587 4636 3813 4644
rect 3827 4636 3873 4644
rect 3987 4636 4033 4644
rect 4147 4636 4193 4644
rect 4347 4636 4593 4644
rect 4847 4636 4873 4644
rect 5107 4636 5153 4644
rect 5647 4636 5673 4644
rect 1607 4616 1753 4624
rect 2247 4616 2333 4624
rect 2367 4616 2593 4624
rect 2787 4616 2833 4624
rect 3007 4616 3113 4624
rect 3127 4616 3293 4624
rect 3307 4616 3373 4624
rect 3507 4616 3713 4624
rect 3787 4616 3933 4624
rect 4447 4616 4653 4624
rect 4667 4616 5013 4624
rect 5087 4616 5113 4624
rect 587 4596 1513 4604
rect 1587 4596 1613 4604
rect 1947 4596 2713 4604
rect 2887 4596 3153 4604
rect 3407 4596 3553 4604
rect 5127 4596 5233 4604
rect 5427 4596 5473 4604
rect 1287 4576 2173 4584
rect 2327 4576 2453 4584
rect 2787 4576 2893 4584
rect 3187 4576 3373 4584
rect 3427 4576 3993 4584
rect 4007 4576 4093 4584
rect 5107 4576 5553 4584
rect 1127 4556 1593 4564
rect 2227 4556 2413 4564
rect 2767 4556 2933 4564
rect 3087 4556 3293 4564
rect 3367 4556 3593 4564
rect 3887 4556 4173 4564
rect 4567 4556 4613 4564
rect 1727 4536 2373 4544
rect 2747 4536 3113 4544
rect 3207 4536 3493 4544
rect 3907 4536 4113 4544
rect 4127 4536 4313 4544
rect 767 4516 1053 4524
rect 1067 4516 1133 4524
rect 1667 4516 1813 4524
rect 2047 4516 2093 4524
rect 2327 4516 2593 4524
rect 2627 4516 2693 4524
rect 2707 4516 2873 4524
rect 2947 4516 2973 4524
rect 3027 4516 3153 4524
rect 3227 4516 3433 4524
rect 3587 4516 3713 4524
rect 3767 4516 3833 4524
rect 3847 4516 4073 4524
rect 5047 4516 5133 4524
rect 5147 4516 5233 4524
rect 207 4496 853 4504
rect 1087 4496 1133 4504
rect 1227 4496 1293 4504
rect 1467 4496 1553 4504
rect 1567 4496 1613 4504
rect 1627 4496 1993 4504
rect 2167 4496 2393 4504
rect 2407 4496 2493 4504
rect 2567 4496 2813 4504
rect 2827 4496 3213 4504
rect 3327 4496 3653 4504
rect 3667 4496 3793 4504
rect 3827 4496 3884 4504
rect 687 4476 713 4484
rect 767 4476 813 4484
rect 927 4476 1093 4484
rect 1107 4476 1113 4484
rect 1167 4476 1184 4484
rect 387 4456 573 4464
rect 887 4456 953 4464
rect 1176 4464 1184 4476
rect 1207 4476 1293 4484
rect 1687 4476 1793 4484
rect 1807 4476 1973 4484
rect 1176 4456 1313 4464
rect 1587 4456 1953 4464
rect 547 4436 593 4444
rect 907 4436 933 4444
rect 1147 4436 1173 4444
rect 1367 4436 1413 4444
rect 2016 4444 2024 4473
rect 2056 4467 2064 4493
rect 2087 4476 2284 4484
rect 2167 4456 2193 4464
rect 2276 4464 2284 4476
rect 2447 4476 2573 4484
rect 2607 4476 2853 4484
rect 2867 4476 2893 4484
rect 2927 4476 2964 4484
rect 2276 4456 2293 4464
rect 2487 4456 2553 4464
rect 2727 4456 2753 4464
rect 2956 4464 2964 4476
rect 2987 4476 3033 4484
rect 3276 4484 3284 4493
rect 3256 4476 3284 4484
rect 2956 4456 3053 4464
rect 2016 4436 2293 4444
rect 2596 4444 2604 4453
rect 3256 4447 3264 4476
rect 3547 4476 3573 4484
rect 3616 4476 3733 4484
rect 3287 4456 3433 4464
rect 3496 4464 3504 4473
rect 3496 4456 3513 4464
rect 3536 4447 3544 4473
rect 3616 4467 3624 4476
rect 3876 4484 3884 4496
rect 3907 4496 3933 4504
rect 3967 4496 4013 4504
rect 4047 4496 4053 4504
rect 4067 4496 4153 4504
rect 4267 4496 4593 4504
rect 5147 4496 5173 4504
rect 5287 4496 5313 4504
rect 5507 4496 5593 4504
rect 3876 4476 3913 4484
rect 4147 4476 4233 4484
rect 4307 4476 4353 4484
rect 5207 4476 5533 4484
rect 3727 4456 3973 4464
rect 4287 4456 4393 4464
rect 4427 4456 4773 4464
rect 4787 4456 5053 4464
rect 5067 4456 5113 4464
rect 5267 4456 5353 4464
rect 2596 4436 2793 4444
rect 2807 4436 3173 4444
rect 3187 4436 3233 4444
rect 3327 4436 3333 4444
rect 3347 4436 3413 4444
rect 3567 4436 3793 4444
rect 4287 4436 4353 4444
rect 4767 4436 5093 4444
rect 5187 4436 5573 4444
rect 467 4416 793 4424
rect 807 4416 893 4424
rect 1187 4416 1693 4424
rect 1867 4416 2053 4424
rect 3527 4416 3553 4424
rect 4127 4416 4213 4424
rect 5027 4416 5433 4424
rect 5447 4416 5453 4424
rect 5627 4416 5693 4424
rect 667 4396 953 4404
rect 1667 4396 2333 4404
rect 4867 4396 5273 4404
rect 1707 4376 1813 4384
rect 2167 4376 2253 4384
rect 4527 4376 4813 4384
rect 5147 4376 5253 4384
rect 847 4356 1073 4364
rect 1087 4356 1193 4364
rect 1827 4356 1893 4364
rect 2327 4356 2613 4364
rect 3167 4356 3373 4364
rect 5267 4356 5513 4364
rect 847 4336 1393 4344
rect 1407 4336 1673 4344
rect 2507 4336 3373 4344
rect 2427 4316 2533 4324
rect 3147 4316 3193 4324
rect 3987 4316 5153 4324
rect 5527 4316 5744 4324
rect 5736 4307 5744 4316
rect 1807 4296 1913 4304
rect 1927 4296 2533 4304
rect 4707 4296 4793 4304
rect 4807 4296 4913 4304
rect 1847 4276 2173 4284
rect 2527 4276 2613 4284
rect 3287 4276 3353 4284
rect 4627 4276 4653 4284
rect 1427 4256 1773 4264
rect 2007 4256 2093 4264
rect 2107 4256 2813 4264
rect 2827 4256 3093 4264
rect 4167 4256 4613 4264
rect 4627 4256 5173 4264
rect 787 4236 1153 4244
rect 1287 4236 1624 4244
rect 1616 4227 1624 4236
rect 1767 4236 1973 4244
rect 2047 4236 2113 4244
rect 2227 4236 2293 4244
rect 2527 4236 2833 4244
rect 2947 4236 2973 4244
rect 3127 4236 3393 4244
rect 3427 4236 3453 4244
rect 3627 4236 3653 4244
rect 3887 4236 3913 4244
rect 4107 4236 4673 4244
rect 5167 4236 5593 4244
rect 947 4216 993 4224
rect 1007 4216 1053 4224
rect 1087 4216 1113 4224
rect 1207 4216 1453 4224
rect 1507 4216 1553 4224
rect 1567 4216 1573 4224
rect 1867 4216 1913 4224
rect 1967 4216 1993 4224
rect 2007 4216 2053 4224
rect 2347 4216 2453 4224
rect 2687 4216 2993 4224
rect 3107 4216 3173 4224
rect 3287 4216 3333 4224
rect 3387 4216 3433 4224
rect 3447 4216 3473 4224
rect 3567 4216 3753 4224
rect 4207 4216 4293 4224
rect 5107 4216 5273 4224
rect 5287 4216 5573 4224
rect 87 4196 513 4204
rect 576 4196 633 4204
rect 576 4187 584 4196
rect 787 4196 853 4204
rect 967 4196 1073 4204
rect 1327 4196 1393 4204
rect 1607 4196 1873 4204
rect 187 4176 533 4184
rect 887 4176 973 4184
rect 1027 4176 1273 4184
rect 1307 4176 1353 4184
rect 1936 4184 1944 4213
rect 2087 4196 2253 4204
rect 2407 4196 2564 4204
rect 1907 4176 1944 4184
rect 1987 4176 2133 4184
rect 2407 4176 2433 4184
rect 2507 4176 2533 4184
rect 2556 4184 2564 4196
rect 2987 4196 3393 4204
rect 3587 4196 3633 4204
rect 3687 4196 3973 4204
rect 4007 4196 4213 4204
rect 4227 4196 4313 4204
rect 4367 4196 4393 4204
rect 4476 4196 4513 4204
rect 2556 4176 2593 4184
rect 2607 4176 2693 4184
rect 2767 4176 2853 4184
rect 2927 4176 2953 4184
rect 3147 4176 3193 4184
rect 3207 4176 3313 4184
rect 3527 4176 3553 4184
rect 3787 4176 4033 4184
rect 4127 4176 4253 4184
rect 4476 4184 4484 4196
rect 4587 4196 4673 4204
rect 4807 4196 4933 4204
rect 5067 4196 5113 4204
rect 5207 4196 5413 4204
rect 4387 4176 4484 4184
rect 4507 4176 4593 4184
rect 4787 4176 5233 4184
rect 487 4156 653 4164
rect 747 4156 753 4164
rect 767 4156 793 4164
rect 807 4156 853 4164
rect 1067 4156 1493 4164
rect 1587 4156 1773 4164
rect 2027 4156 2073 4164
rect 2307 4156 2433 4164
rect 2467 4156 2513 4164
rect 2527 4156 2553 4164
rect 2887 4156 3073 4164
rect 3087 4156 3133 4164
rect 3247 4156 3393 4164
rect 3507 4156 3593 4164
rect 3707 4156 3733 4164
rect 3747 4156 3753 4164
rect 3907 4156 3953 4164
rect 3967 4156 4093 4164
rect 4247 4156 4333 4164
rect 4407 4156 4453 4164
rect 4487 4156 4933 4164
rect 5656 4164 5664 4213
rect 5656 4156 5713 4164
rect 207 4136 553 4144
rect 687 4136 1213 4144
rect 1387 4136 1573 4144
rect 1887 4136 2353 4144
rect 2427 4136 2533 4144
rect 3667 4136 3813 4144
rect 3827 4136 3933 4144
rect 4267 4136 5033 4144
rect 747 4116 833 4124
rect 867 4116 1013 4124
rect 1487 4116 1553 4124
rect 1567 4116 1633 4124
rect 1787 4116 1813 4124
rect 2187 4116 2773 4124
rect 3867 4116 4233 4124
rect 4307 4116 4433 4124
rect 5267 4116 5364 4124
rect 767 4096 1393 4104
rect 2287 4096 2453 4104
rect 2967 4096 3033 4104
rect 3047 4096 3473 4104
rect 3787 4096 4073 4104
rect 4087 4096 4133 4104
rect 4167 4096 4233 4104
rect 4547 4096 4893 4104
rect 5167 4096 5193 4104
rect 5267 4096 5333 4104
rect 5356 4104 5364 4116
rect 5427 4116 5493 4124
rect 5356 4096 5413 4104
rect 847 4076 893 4084
rect 1027 4076 1273 4084
rect 1287 4076 1593 4084
rect 1627 4076 1933 4084
rect 1947 4076 2733 4084
rect 3007 4076 3033 4084
rect 3087 4076 3293 4084
rect 3487 4076 3553 4084
rect 3607 4076 3753 4084
rect 4307 4076 4693 4084
rect 4807 4076 4913 4084
rect 5147 4076 5233 4084
rect 5247 4076 5313 4084
rect 807 4056 913 4064
rect 987 4056 1033 4064
rect 1607 4056 2033 4064
rect 2247 4056 2293 4064
rect 2327 4056 2413 4064
rect 2587 4056 4173 4064
rect 4187 4056 4333 4064
rect 4347 4056 4633 4064
rect 4727 4056 4753 4064
rect 4767 4056 4993 4064
rect 5127 4056 5173 4064
rect 5187 4056 5393 4064
rect 5547 4056 5673 4064
rect 827 4036 853 4044
rect 907 4036 933 4044
rect 1147 4036 1413 4044
rect 1467 4036 1733 4044
rect 1847 4036 2113 4044
rect 2147 4036 2313 4044
rect 2447 4036 2713 4044
rect 3247 4036 3313 4044
rect 3407 4036 3473 4044
rect 3587 4036 3653 4044
rect 3707 4036 3793 4044
rect 4047 4036 4613 4044
rect 4647 4036 5193 4044
rect 5207 4036 5353 4044
rect 5367 4036 5553 4044
rect 5567 4036 5573 4044
rect 5627 4036 5673 4044
rect 207 4016 553 4024
rect 767 4016 893 4024
rect 927 4016 1033 4024
rect 1107 4016 1213 4024
rect 1367 4016 1413 4024
rect 1447 4016 1473 4024
rect 1487 4016 1533 4024
rect 1747 4016 1973 4024
rect 2287 4016 2313 4024
rect 2487 4016 2593 4024
rect 2847 4016 2873 4024
rect 2887 4016 2993 4024
rect 3007 4016 3713 4024
rect 3767 4016 3813 4024
rect 4007 4016 4033 4024
rect 4047 4016 4053 4024
rect 4167 4016 4273 4024
rect 4287 4016 4373 4024
rect 4767 4016 5373 4024
rect 5607 4016 5633 4024
rect 67 3996 693 4004
rect 707 3996 713 4004
rect 887 3996 973 4004
rect 1067 3996 1613 4004
rect 1747 3996 1764 4004
rect 467 3976 593 3984
rect 607 3976 1033 3984
rect 1247 3976 1313 3984
rect 1587 3976 1613 3984
rect 1756 3984 1764 3996
rect 1787 3996 1953 4004
rect 1976 3996 2053 4004
rect 1976 3987 1984 3996
rect 2236 3996 2293 4004
rect 1756 3976 1833 3984
rect 1887 3976 1933 3984
rect 2236 3984 2244 3996
rect 2367 3996 2493 4004
rect 2656 4004 2664 4013
rect 2656 3996 2764 4004
rect 2167 3976 2244 3984
rect 2267 3976 2513 3984
rect 2536 3976 2553 3984
rect 376 3964 384 3973
rect 376 3956 913 3964
rect 1207 3956 1473 3964
rect 1676 3964 1684 3973
rect 1527 3956 1684 3964
rect 2047 3956 2093 3964
rect 2536 3964 2544 3976
rect 2667 3976 2733 3984
rect 2387 3956 2544 3964
rect 2756 3964 2764 3996
rect 2827 3996 2893 4004
rect 3107 3996 3253 4004
rect 3287 3996 3404 4004
rect 2787 3976 2953 3984
rect 2967 3976 2973 3984
rect 3047 3976 3133 3984
rect 3167 3976 3253 3984
rect 3287 3976 3373 3984
rect 2727 3956 2764 3964
rect 2847 3956 2993 3964
rect 3007 3956 3053 3964
rect 3087 3956 3213 3964
rect 3396 3964 3404 3996
rect 3747 3996 3793 4004
rect 3807 3996 3844 4004
rect 3836 3987 3844 3996
rect 3867 3996 4013 4004
rect 4207 3996 4293 4004
rect 4367 3996 4393 4004
rect 4536 3996 4573 4004
rect 3887 3976 3953 3984
rect 3967 3976 3973 3984
rect 4087 3976 4184 3984
rect 4176 3967 4184 3976
rect 4287 3976 4353 3984
rect 4536 3984 4544 3996
rect 5056 3996 5133 4004
rect 4447 3976 4544 3984
rect 4567 3976 4653 3984
rect 3387 3956 3404 3964
rect 3507 3956 3533 3964
rect 4107 3956 4133 3964
rect 4256 3964 4264 3973
rect 4256 3956 4393 3964
rect 5056 3947 5064 3996
rect 5156 3996 5173 4004
rect 5156 3984 5164 3996
rect 5187 3996 5273 4004
rect 5416 3996 5453 4004
rect 5087 3976 5164 3984
rect 5416 3984 5424 3996
rect 5527 3996 5613 4004
rect 5307 3976 5424 3984
rect 5447 3976 5473 3984
rect 5307 3956 5413 3964
rect 867 3936 1153 3944
rect 1507 3936 2693 3944
rect 2707 3936 2833 3944
rect 3067 3936 3093 3944
rect 3147 3936 3233 3944
rect 4027 3936 4213 3944
rect 4327 3936 4453 3944
rect 4507 3936 4513 3944
rect 4527 3936 4753 3944
rect 5127 3936 5593 3944
rect 1547 3916 4113 3924
rect 4607 3916 4633 3924
rect 4707 3916 5333 3924
rect 1647 3896 1913 3904
rect 1927 3896 2013 3904
rect 2027 3896 2793 3904
rect 2807 3896 3093 3904
rect 3107 3896 4473 3904
rect 1367 3876 1393 3884
rect 1407 3876 2893 3884
rect 2907 3876 3013 3884
rect 3027 3876 3153 3884
rect 4347 3876 4373 3884
rect 967 3856 1713 3864
rect 1727 3856 1793 3864
rect 2087 3856 2213 3864
rect 3007 3856 4333 3864
rect 5667 3856 5733 3864
rect 1727 3836 2253 3844
rect 2267 3836 2273 3844
rect 2436 3836 4233 3844
rect 1607 3816 1773 3824
rect 1787 3816 2053 3824
rect 2436 3824 2444 3836
rect 4247 3836 4273 3844
rect 2267 3816 2444 3824
rect 2947 3816 2973 3824
rect 3287 3816 3333 3824
rect 3527 3816 3853 3824
rect 5047 3816 5313 3824
rect 1687 3796 2473 3804
rect 2687 3796 3273 3804
rect 3327 3796 3513 3804
rect 567 3776 633 3784
rect 647 3776 673 3784
rect 1347 3776 1413 3784
rect 2447 3776 3613 3784
rect 4147 3776 4393 3784
rect 4407 3776 4533 3784
rect 4887 3776 4913 3784
rect 5107 3776 5233 3784
rect 727 3756 793 3764
rect 1327 3756 1393 3764
rect 1407 3756 1684 3764
rect 147 3736 233 3744
rect 287 3736 733 3744
rect 787 3736 833 3744
rect 1067 3736 1133 3744
rect 1207 3736 1253 3744
rect 1307 3736 1513 3744
rect 167 3716 253 3724
rect 367 3716 473 3724
rect 927 3716 1013 3724
rect 1387 3716 1413 3724
rect 1436 3724 1444 3736
rect 1676 3744 1684 3756
rect 1787 3756 1973 3764
rect 2456 3756 3164 3764
rect 1676 3736 1993 3744
rect 2007 3736 2073 3744
rect 2107 3736 2353 3744
rect 2456 3744 2464 3756
rect 2367 3736 2464 3744
rect 2487 3736 2513 3744
rect 2587 3736 2613 3744
rect 3156 3744 3164 3756
rect 3187 3756 3253 3764
rect 3327 3756 3453 3764
rect 4127 3756 4913 3764
rect 4927 3756 4933 3764
rect 5007 3756 5253 3764
rect 5287 3756 5613 3764
rect 3156 3736 3173 3744
rect 3227 3736 3353 3744
rect 3407 3736 3433 3744
rect 3467 3736 3673 3744
rect 3787 3736 4193 3744
rect 4447 3736 4973 3744
rect 5156 3736 5193 3744
rect 1436 3716 1613 3724
rect 1707 3716 1773 3724
rect 1927 3716 2113 3724
rect 2227 3716 2433 3724
rect 2447 3716 2493 3724
rect 2636 3724 2644 3733
rect 2527 3716 2644 3724
rect 3007 3716 3133 3724
rect 3327 3716 3493 3724
rect 3647 3716 3733 3724
rect 3767 3716 3833 3724
rect 3847 3716 3873 3724
rect 4007 3716 4113 3724
rect 4236 3707 4244 3733
rect 4256 3716 4373 3724
rect 4256 3707 4264 3716
rect 4456 3716 4513 3724
rect 4456 3707 4464 3716
rect 4687 3716 4793 3724
rect 5156 3707 5164 3736
rect 5207 3716 5233 3724
rect 5587 3716 5733 3724
rect 207 3696 293 3704
rect 727 3696 813 3704
rect 1227 3696 1273 3704
rect 1487 3696 1653 3704
rect 1676 3696 1753 3704
rect 27 3676 213 3684
rect 527 3676 573 3684
rect 587 3676 693 3684
rect 887 3676 973 3684
rect 987 3676 1313 3684
rect 1676 3684 1684 3696
rect 1807 3696 1853 3704
rect 2067 3696 2093 3704
rect 2307 3696 2353 3704
rect 2387 3696 2493 3704
rect 2507 3696 2533 3704
rect 3247 3696 3433 3704
rect 3487 3696 3553 3704
rect 3607 3696 3913 3704
rect 3987 3696 4033 3704
rect 4107 3696 4173 3704
rect 4307 3696 4393 3704
rect 4907 3696 4953 3704
rect 5027 3696 5113 3704
rect 1587 3676 1684 3684
rect 1707 3676 1733 3684
rect 2027 3676 2053 3684
rect 2207 3676 2313 3684
rect 2467 3676 2673 3684
rect 3087 3676 3153 3684
rect 3507 3676 3773 3684
rect 3847 3676 4073 3684
rect 4107 3676 4593 3684
rect 5027 3676 5053 3684
rect 227 3656 693 3664
rect 1087 3656 1213 3664
rect 1527 3656 1813 3664
rect 1827 3656 3013 3664
rect 4227 3656 4353 3664
rect 4587 3656 5033 3664
rect 687 3636 753 3644
rect 1107 3636 1253 3644
rect 1267 3636 1573 3644
rect 1607 3636 2373 3644
rect 2707 3636 2953 3644
rect 3167 3636 3873 3644
rect 3887 3636 4093 3644
rect 4247 3636 4313 3644
rect 4347 3636 4373 3644
rect 4387 3636 4553 3644
rect 5007 3636 5453 3644
rect 67 3616 113 3624
rect 127 3616 853 3624
rect 1147 3616 1693 3624
rect 1787 3616 2193 3624
rect 2307 3616 2393 3624
rect 2947 3616 3053 3624
rect 3307 3616 3333 3624
rect 3587 3616 3793 3624
rect 4187 3616 4393 3624
rect 4467 3616 4733 3624
rect 667 3596 1713 3604
rect 2007 3596 2413 3604
rect 3127 3596 3173 3604
rect 3267 3596 3433 3604
rect 3627 3596 3733 3604
rect 3907 3596 4013 3604
rect 4027 3596 4333 3604
rect 1347 3576 1673 3584
rect 1887 3576 2033 3584
rect 2127 3576 2173 3584
rect 2207 3576 2424 3584
rect 387 3556 1073 3564
rect 1487 3556 1593 3564
rect 1887 3556 2213 3564
rect 2367 3556 2393 3564
rect 2416 3564 2424 3576
rect 2447 3576 2593 3584
rect 3207 3576 3333 3584
rect 3667 3576 4113 3584
rect 4127 3576 4273 3584
rect 2416 3556 2453 3564
rect 2547 3556 2573 3564
rect 2787 3556 2853 3564
rect 3407 3556 3533 3564
rect 3727 3556 3933 3564
rect 3947 3556 4173 3564
rect 187 3536 293 3544
rect 627 3536 984 3544
rect 87 3516 193 3524
rect 207 3516 573 3524
rect 587 3516 593 3524
rect 747 3516 944 3524
rect 936 3507 944 3516
rect 976 3507 984 3536
rect 1167 3536 1273 3544
rect 1287 3536 1293 3544
rect 1447 3536 1513 3544
rect 1647 3536 1733 3544
rect 1787 3536 1813 3544
rect 1847 3536 2553 3544
rect 2707 3536 3153 3544
rect 3267 3536 3353 3544
rect 3427 3536 3613 3544
rect 3707 3536 3753 3544
rect 3767 3536 3813 3544
rect 3987 3536 4133 3544
rect 4427 3536 4833 3544
rect 5207 3536 5533 3544
rect 5616 3536 5653 3544
rect 1007 3516 1093 3524
rect 1247 3516 1653 3524
rect 1847 3516 1953 3524
rect 1987 3516 2153 3524
rect 2187 3516 2313 3524
rect 2596 3524 2604 3533
rect 2487 3516 2604 3524
rect 2727 3516 2813 3524
rect 2987 3516 3553 3524
rect 4047 3516 4493 3524
rect 4507 3516 4593 3524
rect 5107 3516 5253 3524
rect 127 3496 153 3504
rect 267 3496 373 3504
rect 427 3496 513 3504
rect 527 3496 553 3504
rect 647 3496 673 3504
rect 747 3496 773 3504
rect 787 3496 873 3504
rect 1087 3496 1133 3504
rect 1927 3496 2013 3504
rect 2547 3496 2573 3504
rect 2656 3504 2664 3513
rect 2607 3496 2664 3504
rect 2847 3496 2893 3504
rect 3167 3496 3273 3504
rect 3307 3496 3413 3504
rect 3487 3496 3513 3504
rect 147 3476 233 3484
rect 327 3476 433 3484
rect 507 3476 573 3484
rect 667 3476 713 3484
rect 727 3476 853 3484
rect 1247 3476 1313 3484
rect 1427 3476 1493 3484
rect 1616 3484 1624 3493
rect 3696 3487 3704 3513
rect 3727 3496 3753 3504
rect 3787 3496 3833 3504
rect 3996 3504 4004 3513
rect 3847 3496 4004 3504
rect 4207 3496 4293 3504
rect 4347 3496 4513 3504
rect 4667 3496 5313 3504
rect 5327 3496 5353 3504
rect 1616 3476 2133 3484
rect 2147 3476 2193 3484
rect 2387 3476 2493 3484
rect 2627 3476 2753 3484
rect 2996 3476 3633 3484
rect 287 3456 473 3464
rect 616 3464 624 3473
rect 547 3456 624 3464
rect 1707 3456 1893 3464
rect 2027 3456 2113 3464
rect 2167 3456 2613 3464
rect 2996 3464 3004 3476
rect 4087 3476 4133 3484
rect 4367 3476 4433 3484
rect 4447 3476 4493 3484
rect 5047 3476 5073 3484
rect 5227 3476 5253 3484
rect 2767 3456 3004 3464
rect 3027 3456 3313 3464
rect 3647 3456 3673 3464
rect 3887 3456 3953 3464
rect 107 3436 153 3444
rect 347 3436 753 3444
rect 1987 3436 2033 3444
rect 2467 3436 4153 3444
rect 4167 3436 4273 3444
rect 5267 3436 5293 3444
rect 5616 3444 5624 3536
rect 5636 3516 5693 3524
rect 5636 3464 5644 3516
rect 5667 3496 5733 3504
rect 5636 3456 5653 3464
rect 5616 3436 5744 3444
rect 67 3416 93 3424
rect 1047 3416 2213 3424
rect 2627 3416 2893 3424
rect 2967 3416 3593 3424
rect 1127 3396 1593 3404
rect 1607 3396 2673 3404
rect 2687 3396 2833 3404
rect 2847 3396 3133 3404
rect 3827 3396 3913 3404
rect 3927 3396 3973 3404
rect 4887 3396 5133 3404
rect 5147 3396 5273 3404
rect 5627 3396 5653 3404
rect 1207 3376 3473 3384
rect 4927 3376 5013 3384
rect 5736 3367 5744 3436
rect 127 3356 173 3364
rect 187 3356 533 3364
rect 1027 3356 1153 3364
rect 1187 3356 1273 3364
rect 1647 3356 1673 3364
rect 1687 3356 2293 3364
rect 2307 3356 2713 3364
rect 2787 3356 2873 3364
rect 3107 3356 3153 3364
rect 3167 3356 3213 3364
rect 4607 3356 4713 3364
rect 5147 3356 5173 3364
rect 327 3336 433 3344
rect 1427 3336 2033 3344
rect 2047 3336 2633 3344
rect 2887 3336 3193 3344
rect 3207 3336 3313 3344
rect 4187 3336 4673 3344
rect 5507 3336 5553 3344
rect 787 3316 813 3324
rect 1227 3316 1753 3324
rect 1767 3316 2853 3324
rect 807 3296 833 3304
rect 847 3296 853 3304
rect 2667 3296 2933 3304
rect 3056 3296 3493 3304
rect 567 3276 793 3284
rect 1947 3276 2613 3284
rect 2727 3276 2793 3284
rect 2807 3276 2993 3284
rect 3056 3284 3064 3296
rect 4987 3296 5633 3304
rect 5647 3296 5693 3304
rect 3007 3276 3064 3284
rect 3087 3276 3173 3284
rect 3587 3276 3613 3284
rect 3676 3276 3693 3284
rect 3676 3267 3684 3276
rect 4627 3276 5213 3284
rect 5627 3276 5693 3284
rect 67 3256 373 3264
rect 667 3256 893 3264
rect 1547 3256 1593 3264
rect 1747 3256 2133 3264
rect 2407 3256 2553 3264
rect 3067 3256 3613 3264
rect 4207 3256 4233 3264
rect 4947 3256 5144 3264
rect 307 3236 333 3244
rect 487 3236 633 3244
rect 687 3236 733 3244
rect 887 3236 973 3244
rect 1267 3236 1713 3244
rect 1836 3236 1933 3244
rect 1836 3227 1844 3236
rect 2187 3236 2253 3244
rect 2267 3236 2333 3244
rect 2387 3236 2413 3244
rect 2427 3236 2473 3244
rect 2567 3236 2633 3244
rect 2647 3236 2673 3244
rect 2716 3236 2793 3244
rect 147 3216 153 3224
rect 167 3216 273 3224
rect 407 3216 433 3224
rect 447 3216 613 3224
rect 767 3216 813 3224
rect 1307 3216 1353 3224
rect 1407 3216 1473 3224
rect 1667 3216 1753 3224
rect 1776 3216 1793 3224
rect 327 3196 413 3204
rect 427 3196 473 3204
rect 507 3196 673 3204
rect 1187 3196 1293 3204
rect 1467 3196 1493 3204
rect 1567 3196 1693 3204
rect 1776 3204 1784 3216
rect 1936 3216 2113 3224
rect 1936 3207 1944 3216
rect 2167 3216 2573 3224
rect 2587 3216 2653 3224
rect 2716 3224 2724 3236
rect 2707 3216 2724 3224
rect 2856 3224 2864 3253
rect 5136 3247 5144 3256
rect 3147 3236 3173 3244
rect 3587 3236 3653 3244
rect 4136 3236 4293 3244
rect 2747 3216 2973 3224
rect 3027 3216 3093 3224
rect 3356 3224 3364 3233
rect 4136 3227 4144 3236
rect 4447 3236 4633 3244
rect 4747 3236 4813 3244
rect 4847 3236 4873 3244
rect 3247 3216 3364 3224
rect 3547 3216 3593 3224
rect 3607 3216 3833 3224
rect 4807 3216 4933 3224
rect 4947 3216 4973 3224
rect 1767 3196 1784 3204
rect 1827 3196 1873 3204
rect 1967 3196 2113 3204
rect 2287 3196 2313 3204
rect 2467 3196 2613 3204
rect 2807 3196 2873 3204
rect 2967 3196 3133 3204
rect 3167 3196 3193 3204
rect 4427 3196 4613 3204
rect 4867 3196 4993 3204
rect 5007 3196 5093 3204
rect 187 3176 333 3184
rect 347 3176 353 3184
rect 1007 3176 1573 3184
rect 1627 3176 1733 3184
rect 2067 3176 2133 3184
rect 2147 3176 2233 3184
rect 2547 3176 3153 3184
rect 3787 3176 4853 3184
rect 447 3156 893 3164
rect 907 3156 1313 3164
rect 1327 3156 1413 3164
rect 1547 3156 1573 3164
rect 1596 3156 1833 3164
rect 607 3136 633 3144
rect 647 3136 713 3144
rect 1596 3144 1604 3156
rect 1927 3156 2073 3164
rect 2247 3156 2533 3164
rect 2587 3156 2733 3164
rect 2867 3156 2913 3164
rect 2987 3156 3104 3164
rect 1487 3136 1604 3144
rect 1767 3136 1953 3144
rect 1987 3136 2033 3144
rect 2127 3136 2404 3144
rect 1567 3116 2373 3124
rect 2396 3124 2404 3136
rect 2427 3136 2673 3144
rect 2687 3136 2713 3144
rect 2767 3136 2853 3144
rect 3096 3144 3104 3156
rect 3127 3156 3353 3164
rect 4127 3156 4233 3164
rect 3096 3136 3213 3144
rect 3267 3136 3353 3144
rect 4667 3136 4793 3144
rect 5127 3136 5153 3144
rect 2396 3116 2613 3124
rect 2667 3116 3184 3124
rect 1467 3096 1653 3104
rect 1787 3096 1833 3104
rect 2527 3096 2633 3104
rect 3027 3096 3093 3104
rect 3176 3104 3184 3116
rect 3207 3116 3473 3124
rect 3887 3116 4453 3124
rect 4507 3116 5473 3124
rect 3176 3096 3273 3104
rect 1147 3076 1513 3084
rect 1607 3076 1633 3084
rect 1767 3076 1853 3084
rect 1887 3076 2113 3084
rect 2127 3076 2173 3084
rect 2447 3076 2593 3084
rect 2707 3076 2953 3084
rect 3087 3076 3113 3084
rect 3247 3076 3313 3084
rect 4007 3076 4353 3084
rect 407 3056 593 3064
rect 627 3056 733 3064
rect 1507 3056 1633 3064
rect 1727 3056 1773 3064
rect 1787 3056 1793 3064
rect 1807 3056 1933 3064
rect 1947 3056 1993 3064
rect 2067 3056 2353 3064
rect 2367 3056 2393 3064
rect 2427 3056 2513 3064
rect 2627 3056 2804 3064
rect 87 3036 233 3044
rect 247 3036 253 3044
rect 307 3036 373 3044
rect 447 3036 473 3044
rect 487 3036 573 3044
rect 1627 3036 1693 3044
rect 1707 3036 1913 3044
rect 2167 3036 2313 3044
rect 2347 3036 2453 3044
rect 2487 3036 2573 3044
rect 2647 3036 2773 3044
rect 2796 3044 2804 3056
rect 2847 3056 2873 3064
rect 2896 3056 3033 3064
rect 2896 3044 2904 3056
rect 3047 3056 3173 3064
rect 3187 3056 3233 3064
rect 3467 3056 3513 3064
rect 3707 3056 3733 3064
rect 3767 3056 3813 3064
rect 3827 3056 4213 3064
rect 4267 3056 4313 3064
rect 4687 3056 4833 3064
rect 4907 3056 4933 3064
rect 5087 3056 5453 3064
rect 2796 3036 2904 3044
rect 2947 3036 2973 3044
rect 3087 3036 3304 3044
rect 427 3016 533 3024
rect 667 3016 693 3024
rect 847 3016 1333 3024
rect 1407 3016 1613 3024
rect 1936 3016 1973 3024
rect 107 2996 213 3004
rect 287 2996 333 3004
rect 647 2996 713 3004
rect 867 2996 973 3004
rect 1607 2996 1653 3004
rect 1936 3004 1944 3016
rect 2136 3024 2144 3033
rect 2107 3016 2244 3024
rect 1867 2996 1944 3004
rect 1967 2996 2013 3004
rect 2067 2996 2133 3004
rect 2187 2996 2213 3004
rect 2236 3004 2244 3016
rect 2636 3024 2644 3033
rect 2447 3016 2644 3024
rect 2747 3016 2753 3024
rect 2767 3016 2893 3024
rect 3036 3024 3044 3033
rect 2907 3016 3044 3024
rect 3107 3016 3193 3024
rect 3296 3024 3304 3036
rect 3327 3036 3333 3044
rect 3347 3036 3513 3044
rect 4307 3036 4373 3044
rect 4387 3036 4513 3044
rect 4547 3036 4613 3044
rect 4887 3036 5013 3044
rect 3296 3016 3393 3024
rect 3427 3016 3544 3024
rect 3536 3007 3544 3016
rect 2236 2996 2253 3004
rect 2307 2996 2373 3004
rect 2747 2996 2853 3004
rect 3307 2996 3353 3004
rect 3447 2996 3473 3004
rect 67 2976 133 2984
rect 147 2976 153 2984
rect 1287 2976 1313 2984
rect 2007 2976 2073 2984
rect 2087 2976 2433 2984
rect 2547 2976 2913 2984
rect 3067 2976 3153 2984
rect 3347 2976 3373 2984
rect 3536 2984 3544 2993
rect 3556 2987 3564 3033
rect 4127 3016 4213 3024
rect 4347 3016 4473 3024
rect 4607 3016 4733 3024
rect 4747 3016 4853 3024
rect 4907 3016 4973 3024
rect 5127 3016 5193 3024
rect 4447 2996 4593 3004
rect 4767 2996 4833 3004
rect 5047 2996 5093 3004
rect 5107 2996 5133 3004
rect 3527 2976 3544 2984
rect 4127 2976 4413 2984
rect 4807 2976 4893 2984
rect 4907 2976 5093 2984
rect 5587 2976 5713 2984
rect 927 2956 1713 2964
rect 1827 2956 2573 2964
rect 2587 2956 2773 2964
rect 2967 2956 3133 2964
rect 3367 2956 3413 2964
rect 4807 2956 5053 2964
rect 67 2936 113 2944
rect 127 2936 593 2944
rect 607 2936 653 2944
rect 1967 2936 2033 2944
rect 2067 2936 2113 2944
rect 2327 2936 2833 2944
rect 447 2916 793 2924
rect 807 2916 1213 2924
rect 1247 2916 1473 2924
rect 1667 2916 1713 2924
rect 1947 2916 2273 2924
rect 2287 2916 2293 2924
rect 2316 2916 2624 2924
rect 1187 2896 1433 2904
rect 2316 2904 2324 2916
rect 1687 2896 2324 2904
rect 2427 2896 2593 2904
rect 2616 2904 2624 2916
rect 2787 2916 4253 2924
rect 4267 2916 4913 2924
rect 5607 2916 5633 2924
rect 5716 2924 5724 2933
rect 5647 2916 5724 2924
rect 2616 2896 3673 2904
rect 3767 2896 3833 2904
rect 3847 2896 3913 2904
rect 1547 2876 1573 2884
rect 1587 2876 1873 2884
rect 2047 2876 2153 2884
rect 2407 2876 2993 2884
rect 4047 2876 4073 2884
rect 4087 2876 4153 2884
rect 1467 2856 1653 2864
rect 2187 2856 2273 2864
rect 2287 2856 2433 2864
rect 2447 2856 2533 2864
rect 4567 2856 4913 2864
rect 227 2836 673 2844
rect 1907 2836 1993 2844
rect 2507 2836 2533 2844
rect 2847 2836 3233 2844
rect 4907 2836 4953 2844
rect 347 2816 653 2824
rect 867 2816 893 2824
rect 907 2816 913 2824
rect 1707 2816 1973 2824
rect 1987 2816 2313 2824
rect 2336 2816 2513 2824
rect 427 2796 453 2804
rect 687 2796 693 2804
rect 707 2796 913 2804
rect 1647 2796 1833 2804
rect 2176 2796 2213 2804
rect 327 2776 393 2784
rect 507 2776 553 2784
rect 807 2776 833 2784
rect 887 2776 1044 2784
rect 167 2756 233 2764
rect 307 2756 333 2764
rect 407 2756 993 2764
rect 1007 2756 1013 2764
rect 1036 2764 1044 2776
rect 1167 2776 1193 2784
rect 1227 2776 1333 2784
rect 1347 2776 1853 2784
rect 1036 2756 1133 2764
rect 1487 2756 1593 2764
rect 1676 2764 1684 2776
rect 1896 2776 2013 2784
rect 1676 2756 1753 2764
rect 1787 2756 1833 2764
rect 1896 2747 1904 2776
rect 2036 2767 2044 2793
rect 1947 2756 2024 2764
rect 107 2736 133 2744
rect 187 2736 353 2744
rect 387 2736 473 2744
rect 567 2736 613 2744
rect 727 2736 813 2744
rect 907 2736 933 2744
rect 956 2736 1093 2744
rect 187 2716 253 2724
rect 267 2716 413 2724
rect 956 2724 964 2736
rect 1127 2736 1153 2744
rect 1667 2736 1693 2744
rect 1736 2736 1853 2744
rect 847 2716 964 2724
rect 987 2716 1013 2724
rect 1736 2724 1744 2736
rect 2016 2744 2024 2756
rect 2176 2764 2184 2796
rect 2336 2804 2344 2816
rect 3227 2816 3333 2824
rect 2316 2796 2344 2804
rect 2207 2776 2284 2784
rect 2176 2756 2253 2764
rect 2276 2747 2284 2776
rect 2316 2767 2324 2796
rect 2407 2796 2613 2804
rect 2627 2796 2704 2804
rect 2387 2776 2424 2784
rect 2416 2764 2424 2776
rect 2447 2776 2473 2784
rect 2527 2776 2573 2784
rect 2696 2784 2704 2796
rect 2727 2796 2753 2804
rect 3087 2796 3113 2804
rect 3227 2796 3253 2804
rect 3267 2796 3493 2804
rect 4087 2796 4233 2804
rect 4707 2796 4853 2804
rect 2696 2776 2853 2784
rect 2947 2776 2993 2784
rect 3047 2776 3113 2784
rect 3316 2776 3513 2784
rect 2416 2756 2444 2764
rect 2016 2736 2133 2744
rect 2307 2736 2333 2744
rect 2436 2744 2444 2756
rect 2827 2756 2873 2764
rect 3316 2764 3324 2776
rect 3607 2776 3733 2784
rect 4067 2776 4093 2784
rect 4107 2776 4173 2784
rect 4247 2776 4713 2784
rect 4767 2776 4773 2784
rect 4787 2776 5033 2784
rect 5047 2776 5153 2784
rect 2987 2756 3324 2764
rect 3347 2756 3364 2764
rect 3356 2747 3364 2756
rect 3407 2756 3453 2764
rect 3547 2756 3573 2764
rect 4707 2756 4953 2764
rect 5127 2756 5173 2764
rect 2436 2736 2553 2744
rect 2927 2736 3013 2744
rect 3107 2736 3173 2744
rect 3247 2736 3353 2744
rect 1487 2716 1744 2724
rect 1767 2716 1913 2724
rect 2067 2716 2153 2724
rect 2287 2716 2573 2724
rect 2787 2716 2833 2724
rect 3167 2716 3273 2724
rect 3547 2716 3653 2724
rect 3716 2707 3724 2753
rect 4176 2744 4184 2753
rect 4127 2736 4184 2744
rect 4747 2736 4813 2744
rect 4847 2736 4893 2744
rect 4927 2736 5013 2744
rect 5107 2736 5233 2744
rect 5267 2736 5293 2744
rect 5627 2736 5693 2744
rect 4247 2716 4333 2724
rect 4607 2716 4733 2724
rect 5007 2716 5173 2724
rect 5587 2716 5653 2724
rect 247 2696 1033 2704
rect 1767 2696 1813 2704
rect 1847 2696 1993 2704
rect 2007 2696 2133 2704
rect 2207 2696 2453 2704
rect 2627 2696 2693 2704
rect 2707 2696 3233 2704
rect 3247 2696 3333 2704
rect 3347 2696 3413 2704
rect 4647 2696 5473 2704
rect 427 2676 813 2684
rect 827 2676 873 2684
rect 896 2676 1253 2684
rect 896 2664 904 2676
rect 1267 2676 1633 2684
rect 1747 2676 1773 2684
rect 3267 2676 3293 2684
rect 3507 2676 3813 2684
rect 4227 2676 4513 2684
rect 747 2656 904 2664
rect 967 2656 1173 2664
rect 1347 2656 1373 2664
rect 1447 2656 1833 2664
rect 1907 2656 1973 2664
rect 1987 2656 2353 2664
rect 2487 2656 3573 2664
rect 3807 2656 4053 2664
rect 4067 2656 4133 2664
rect 4307 2656 4413 2664
rect 4447 2656 4793 2664
rect 527 2636 693 2644
rect 767 2636 1773 2644
rect 2047 2636 2593 2644
rect 2607 2636 2973 2644
rect 3227 2636 3273 2644
rect 3687 2636 3853 2644
rect 4207 2636 4473 2644
rect 4687 2636 4773 2644
rect 87 2616 253 2624
rect 667 2616 753 2624
rect 1107 2616 1113 2624
rect 1127 2616 1233 2624
rect 1327 2616 1673 2624
rect 1887 2616 2013 2624
rect 2187 2616 2733 2624
rect 2787 2616 3753 2624
rect 4267 2616 4553 2624
rect 4567 2616 4773 2624
rect 4887 2616 5393 2624
rect 127 2596 133 2604
rect 147 2596 1293 2604
rect 1327 2596 1353 2604
rect 1527 2596 1553 2604
rect 1607 2596 2104 2604
rect 87 2576 133 2584
rect 567 2576 644 2584
rect 307 2556 353 2564
rect 407 2556 433 2564
rect 527 2556 593 2564
rect 636 2564 644 2576
rect 667 2576 733 2584
rect 747 2576 853 2584
rect 1307 2576 1793 2584
rect 1807 2576 2073 2584
rect 2096 2584 2104 2596
rect 2127 2596 2253 2604
rect 2507 2596 2613 2604
rect 2627 2596 2653 2604
rect 2967 2596 3133 2604
rect 3227 2596 3293 2604
rect 3467 2596 3693 2604
rect 4207 2596 4273 2604
rect 4327 2596 4904 2604
rect 2096 2576 2513 2584
rect 2667 2576 3173 2584
rect 3187 2576 4073 2584
rect 4187 2576 4273 2584
rect 4287 2576 4373 2584
rect 4896 2584 4904 2596
rect 5067 2596 5473 2604
rect 5487 2596 5713 2604
rect 4896 2576 5273 2584
rect 636 2556 713 2564
rect 727 2556 773 2564
rect 847 2556 1053 2564
rect 1427 2556 1544 2564
rect 236 2536 433 2544
rect 236 2527 244 2536
rect 616 2544 624 2553
rect 1536 2547 1544 2556
rect 1727 2556 1833 2564
rect 1856 2556 1973 2564
rect 447 2536 624 2544
rect 807 2536 1093 2544
rect 1396 2536 1473 2544
rect 1396 2527 1404 2536
rect 1856 2544 1864 2556
rect 2027 2556 2173 2564
rect 2407 2556 2453 2564
rect 2807 2556 3053 2564
rect 3087 2556 3133 2564
rect 3207 2556 3313 2564
rect 3347 2556 3473 2564
rect 3507 2556 3613 2564
rect 4327 2556 4353 2564
rect 4407 2556 4433 2564
rect 4876 2564 4884 2573
rect 5056 2567 5064 2576
rect 5447 2576 5633 2584
rect 4876 2556 5033 2564
rect 5087 2556 5253 2564
rect 5367 2556 5564 2564
rect 1587 2536 1864 2544
rect 2107 2536 2193 2544
rect 2427 2536 2493 2544
rect 2527 2536 2553 2544
rect 2636 2544 2644 2553
rect 2616 2536 3533 2544
rect 487 2516 1273 2524
rect 1287 2516 1353 2524
rect 1607 2516 1693 2524
rect 2616 2524 2624 2536
rect 3587 2536 3613 2544
rect 4267 2536 4493 2544
rect 4607 2536 4753 2544
rect 5047 2536 5233 2544
rect 5247 2536 5393 2544
rect 5416 2536 5533 2544
rect 5416 2527 5424 2536
rect 5556 2544 5564 2556
rect 5556 2536 5653 2544
rect 5696 2544 5704 2553
rect 5696 2536 5713 2544
rect 2167 2516 2624 2524
rect 2647 2516 3093 2524
rect 3187 2516 3213 2524
rect 3527 2516 3553 2524
rect 3607 2516 3713 2524
rect 4087 2516 4533 2524
rect 4547 2516 4713 2524
rect 4867 2516 5133 2524
rect 5147 2516 5253 2524
rect 5267 2516 5293 2524
rect 5387 2516 5413 2524
rect 5487 2516 5553 2524
rect 5627 2516 5693 2524
rect 107 2496 433 2504
rect 447 2496 573 2504
rect 647 2496 1033 2504
rect 1047 2496 1233 2504
rect 1247 2496 3053 2504
rect 3067 2496 5013 2504
rect 5587 2496 5653 2504
rect 467 2476 793 2484
rect 827 2476 933 2484
rect 1027 2476 1153 2484
rect 1187 2476 1253 2484
rect 2007 2476 2613 2484
rect 2707 2476 2753 2484
rect 2767 2476 3173 2484
rect 3187 2476 3253 2484
rect 3647 2476 3693 2484
rect 4347 2476 4413 2484
rect 4507 2476 4673 2484
rect 5147 2476 5193 2484
rect 5527 2476 5713 2484
rect 427 2456 904 2464
rect 896 2444 904 2456
rect 967 2456 1093 2464
rect 1647 2456 1733 2464
rect 2187 2456 3693 2464
rect 3776 2464 3784 2473
rect 3727 2456 3784 2464
rect 4507 2456 4573 2464
rect 5607 2456 5713 2464
rect 896 2436 2173 2444
rect 2507 2436 2533 2444
rect 2567 2436 2713 2444
rect 2947 2436 2973 2444
rect 3107 2436 3584 2444
rect 827 2416 1313 2424
rect 1367 2416 3553 2424
rect 3576 2424 3584 2436
rect 3947 2436 3973 2444
rect 4307 2436 4413 2444
rect 4747 2436 4893 2444
rect 5027 2436 5673 2444
rect 3576 2416 4553 2424
rect 1487 2396 1513 2404
rect 2587 2396 2913 2404
rect 2987 2396 3764 2404
rect 27 2376 1313 2384
rect 2227 2376 2573 2384
rect 2587 2376 2893 2384
rect 3527 2376 3733 2384
rect 3756 2384 3764 2396
rect 4207 2396 4933 2404
rect 3756 2376 5133 2384
rect 347 2356 2973 2364
rect 3267 2356 3373 2364
rect 3487 2356 3593 2364
rect 3616 2356 3653 2364
rect 867 2336 1393 2344
rect 3616 2344 3624 2356
rect 3667 2356 3853 2364
rect 3867 2356 4033 2364
rect 4787 2356 4913 2364
rect 5247 2356 5513 2364
rect 1867 2336 3624 2344
rect 3636 2336 4013 2344
rect 227 2316 253 2324
rect 887 2316 984 2324
rect 187 2296 233 2304
rect 407 2296 453 2304
rect 976 2304 984 2316
rect 1007 2316 1053 2324
rect 1087 2316 1113 2324
rect 1787 2316 1893 2324
rect 2287 2316 2653 2324
rect 3027 2316 3333 2324
rect 3636 2324 3644 2336
rect 4027 2336 4513 2344
rect 5367 2336 5473 2344
rect 3347 2316 3644 2324
rect 3747 2316 3793 2324
rect 3827 2316 4853 2324
rect 5347 2316 5533 2324
rect 976 2296 993 2304
rect 1087 2296 1124 2304
rect 167 2276 353 2284
rect 367 2276 493 2284
rect 687 2276 773 2284
rect 807 2276 853 2284
rect 896 2284 904 2293
rect 1036 2284 1044 2293
rect 896 2276 1004 2284
rect 1036 2276 1093 2284
rect 107 2256 193 2264
rect 247 2256 273 2264
rect 447 2256 573 2264
rect 887 2256 913 2264
rect 996 2264 1004 2276
rect 996 2256 1073 2264
rect 1116 2264 1124 2296
rect 1887 2296 2053 2304
rect 2107 2296 2153 2304
rect 2367 2296 2373 2304
rect 2387 2296 2693 2304
rect 2747 2296 2793 2304
rect 2807 2296 3293 2304
rect 3627 2296 3753 2304
rect 3767 2296 3833 2304
rect 4067 2296 4173 2304
rect 4487 2296 4533 2304
rect 4567 2296 4693 2304
rect 5227 2296 5293 2304
rect 5387 2296 5413 2304
rect 5467 2296 5493 2304
rect 5527 2296 5573 2304
rect 1316 2276 1533 2284
rect 1107 2256 1124 2264
rect 1196 2247 1204 2273
rect 1236 2264 1244 2273
rect 1236 2256 1264 2264
rect 127 2236 153 2244
rect 247 2236 253 2244
rect 267 2236 313 2244
rect 527 2236 533 2244
rect 547 2236 753 2244
rect 1047 2236 1113 2244
rect 1256 2244 1264 2256
rect 1256 2236 1273 2244
rect 207 2216 373 2224
rect 607 2216 1093 2224
rect 1316 2224 1324 2276
rect 1687 2276 1713 2284
rect 1827 2276 1893 2284
rect 1947 2276 2013 2284
rect 2067 2276 2244 2284
rect 1347 2256 1413 2264
rect 1507 2256 2213 2264
rect 2236 2264 2244 2276
rect 2427 2276 2813 2284
rect 3027 2276 3053 2284
rect 3507 2276 3544 2284
rect 2236 2256 2293 2264
rect 2316 2247 2324 2273
rect 2416 2264 2424 2273
rect 2336 2256 2424 2264
rect 2336 2247 2344 2256
rect 2467 2256 2593 2264
rect 2667 2256 2684 2264
rect 1407 2236 1433 2244
rect 1487 2236 1553 2244
rect 1607 2236 1693 2244
rect 1767 2236 1833 2244
rect 2507 2236 2653 2244
rect 2676 2244 2684 2256
rect 2787 2256 2873 2264
rect 2927 2256 3033 2264
rect 3396 2264 3404 2273
rect 3536 2267 3544 2276
rect 3927 2276 3953 2284
rect 4027 2276 4053 2284
rect 4147 2276 4164 2284
rect 3287 2256 3404 2264
rect 3747 2256 3893 2264
rect 3947 2256 3993 2264
rect 4007 2256 4133 2264
rect 2676 2236 2753 2244
rect 2967 2236 3233 2244
rect 3267 2236 3353 2244
rect 3547 2236 3553 2244
rect 3567 2236 3713 2244
rect 3887 2236 3953 2244
rect 4156 2244 4164 2276
rect 4447 2276 4573 2284
rect 4587 2276 4593 2284
rect 4967 2276 5073 2284
rect 5056 2267 5064 2276
rect 5127 2276 5433 2284
rect 5067 2256 5513 2264
rect 4156 2236 4873 2244
rect 5027 2236 5093 2244
rect 5187 2236 5213 2244
rect 5307 2236 5493 2244
rect 5536 2244 5544 2273
rect 5527 2236 5544 2244
rect 5616 2244 5624 2273
rect 5647 2256 5673 2264
rect 5616 2236 5633 2244
rect 1187 2216 1324 2224
rect 1467 2216 1513 2224
rect 1527 2216 1853 2224
rect 2267 2216 2513 2224
rect 2527 2216 2733 2224
rect 2827 2216 3113 2224
rect 3127 2216 3833 2224
rect 3927 2216 3973 2224
rect 5087 2216 5153 2224
rect 5427 2216 5493 2224
rect 5587 2216 5613 2224
rect 87 2196 253 2204
rect 267 2196 613 2204
rect 1287 2196 1353 2204
rect 1627 2196 1973 2204
rect 2327 2196 2433 2204
rect 2467 2196 2533 2204
rect 2567 2196 2673 2204
rect 2707 2196 2833 2204
rect 2847 2196 3053 2204
rect 3187 2196 3493 2204
rect 4327 2196 4353 2204
rect 5147 2196 5413 2204
rect 5427 2196 5453 2204
rect 5547 2196 5593 2204
rect 5627 2196 5693 2204
rect 307 2176 453 2184
rect 467 2176 653 2184
rect 707 2176 1653 2184
rect 1727 2176 2113 2184
rect 2167 2176 2433 2184
rect 2487 2176 2513 2184
rect 2547 2176 2713 2184
rect 2907 2176 3024 2184
rect 427 2156 1213 2164
rect 2147 2156 2553 2164
rect 2607 2156 2853 2164
rect 2887 2156 2973 2164
rect 3016 2164 3024 2176
rect 3087 2176 3093 2184
rect 3107 2176 3713 2184
rect 3727 2176 3933 2184
rect 3967 2176 4093 2184
rect 4127 2176 4213 2184
rect 4347 2176 4393 2184
rect 4827 2176 4893 2184
rect 5147 2176 5193 2184
rect 5267 2176 5553 2184
rect 3016 2156 3153 2164
rect 3167 2156 3293 2164
rect 3427 2156 3573 2164
rect 3707 2156 3813 2164
rect 4007 2156 4253 2164
rect 5127 2156 5693 2164
rect 307 2136 433 2144
rect 787 2136 973 2144
rect 1307 2136 1493 2144
rect 1947 2136 2013 2144
rect 2027 2136 2233 2144
rect 2407 2136 2633 2144
rect 2767 2136 3173 2144
rect 3327 2136 3453 2144
rect 3467 2136 3773 2144
rect 3987 2136 4113 2144
rect 4527 2136 4613 2144
rect 4807 2136 4913 2144
rect 5047 2136 5073 2144
rect 5487 2136 5553 2144
rect 107 2116 453 2124
rect 487 2116 533 2124
rect 607 2116 713 2124
rect 1067 2116 1113 2124
rect 1167 2116 1293 2124
rect 1356 2116 1733 2124
rect 207 2096 213 2104
rect 227 2096 273 2104
rect 507 2096 653 2104
rect 756 2096 793 2104
rect 116 2076 293 2084
rect 116 2067 124 2076
rect 307 2056 353 2064
rect 27 2036 53 2044
rect 227 2036 273 2044
rect 376 2044 384 2093
rect 396 2076 513 2084
rect 396 2067 404 2076
rect 536 2076 693 2084
rect 536 2064 544 2076
rect 736 2084 744 2093
rect 716 2076 744 2084
rect 527 2056 544 2064
rect 376 2036 393 2044
rect 716 2044 724 2076
rect 756 2064 764 2096
rect 816 2096 833 2104
rect 816 2084 824 2096
rect 1107 2096 1193 2104
rect 1356 2104 1364 2116
rect 1787 2116 1813 2124
rect 1827 2116 2033 2124
rect 2067 2116 2173 2124
rect 2647 2116 2784 2124
rect 1207 2096 1364 2104
rect 796 2076 824 2084
rect 836 2076 913 2084
rect 796 2067 804 2076
rect 747 2056 764 2064
rect 836 2064 844 2076
rect 1027 2076 1313 2084
rect 816 2056 844 2064
rect 707 2036 724 2044
rect 816 2044 824 2056
rect 867 2056 953 2064
rect 967 2056 1053 2064
rect 1087 2056 1173 2064
rect 767 2036 824 2044
rect 887 2036 1033 2044
rect 1336 2044 1344 2073
rect 1356 2064 1364 2096
rect 1387 2096 1453 2104
rect 1467 2096 1473 2104
rect 1507 2096 1593 2104
rect 1807 2096 1833 2104
rect 2007 2096 2073 2104
rect 2147 2096 2173 2104
rect 2427 2096 2453 2104
rect 2487 2096 2493 2104
rect 2507 2096 2573 2104
rect 2596 2096 2753 2104
rect 1387 2076 1644 2084
rect 1356 2056 1533 2064
rect 1047 2036 1344 2044
rect 1636 2044 1644 2076
rect 1656 2076 1773 2084
rect 1656 2067 1664 2076
rect 2207 2076 2213 2084
rect 2596 2084 2604 2096
rect 2776 2104 2784 2116
rect 2807 2116 2853 2124
rect 2947 2116 2973 2124
rect 3447 2116 3613 2124
rect 3647 2116 3733 2124
rect 4087 2116 4173 2124
rect 4567 2116 4773 2124
rect 4927 2116 5033 2124
rect 5067 2116 5173 2124
rect 5387 2116 5573 2124
rect 2776 2096 2793 2104
rect 2927 2096 2984 2104
rect 2227 2076 2604 2084
rect 2627 2076 2753 2084
rect 2847 2076 2953 2084
rect 2976 2084 2984 2096
rect 3007 2096 3033 2104
rect 3087 2096 3113 2104
rect 3147 2096 3353 2104
rect 3447 2096 3573 2104
rect 3787 2096 3813 2104
rect 3827 2096 4153 2104
rect 4167 2096 4473 2104
rect 4507 2096 4533 2104
rect 4547 2096 4673 2104
rect 4747 2096 4893 2104
rect 4907 2096 5113 2104
rect 5227 2096 5473 2104
rect 5536 2096 5653 2104
rect 2976 2076 3064 2084
rect 2087 2056 2113 2064
rect 2256 2056 2333 2064
rect 2256 2047 2264 2056
rect 1636 2036 1673 2044
rect 1867 2036 1893 2044
rect 2467 2036 2573 2044
rect 2756 2044 2764 2073
rect 2787 2056 2853 2064
rect 2956 2064 2964 2073
rect 3056 2067 3064 2076
rect 3167 2076 3204 2084
rect 2956 2056 3033 2064
rect 3116 2047 3124 2073
rect 2756 2036 2773 2044
rect 2867 2036 2893 2044
rect 3196 2044 3204 2076
rect 3407 2076 3484 2084
rect 3476 2067 3484 2076
rect 3507 2076 3793 2084
rect 3807 2076 3973 2084
rect 4147 2076 4313 2084
rect 4327 2076 4453 2084
rect 4587 2076 4653 2084
rect 4847 2076 4993 2084
rect 5167 2076 5193 2084
rect 5267 2076 5313 2084
rect 5427 2076 5464 2084
rect 3407 2056 3453 2064
rect 3587 2056 3593 2064
rect 3607 2056 3773 2064
rect 4207 2056 4233 2064
rect 4387 2056 4744 2064
rect 3196 2036 3233 2044
rect 3387 2036 3753 2044
rect 3907 2036 4013 2044
rect 4047 2036 4093 2044
rect 4147 2036 4173 2044
rect 4187 2036 4493 2044
rect 4667 2036 4713 2044
rect 4736 2044 4744 2056
rect 4767 2056 5073 2064
rect 5087 2056 5233 2064
rect 5367 2056 5433 2064
rect 4736 2036 5013 2044
rect 5067 2036 5113 2044
rect 5276 2044 5284 2053
rect 5276 2036 5333 2044
rect 5456 2044 5464 2076
rect 5536 2064 5544 2096
rect 5507 2056 5544 2064
rect 5556 2047 5564 2073
rect 5456 2036 5473 2044
rect 5656 2044 5664 2073
rect 5656 2036 5693 2044
rect 947 2016 973 2024
rect 1007 2016 1093 2024
rect 1267 2016 1353 2024
rect 1367 2016 1493 2024
rect 2047 2016 2093 2024
rect 2187 2016 2353 2024
rect 2427 2016 2453 2024
rect 2507 2016 2533 2024
rect 2547 2016 2573 2024
rect 2647 2016 2813 2024
rect 3207 2016 3393 2024
rect 3907 2016 3993 2024
rect 4287 2016 4633 2024
rect 5207 2016 5673 2024
rect 267 1996 413 2004
rect 847 1996 893 2004
rect 907 1996 1153 2004
rect 1287 1996 1373 2004
rect 1727 1996 2133 2004
rect 2167 1996 2313 2004
rect 2447 1996 2673 2004
rect 2807 1996 2973 2004
rect 3287 1996 3573 2004
rect 3747 1996 4173 2004
rect 4347 1996 4753 2004
rect 4947 1996 5393 2004
rect 5407 1996 5413 2004
rect 5527 1996 5593 2004
rect 327 1976 493 1984
rect 1087 1976 1353 1984
rect 1367 1976 1393 1984
rect 2047 1976 2593 1984
rect 2827 1976 2933 1984
rect 2947 1976 3153 1984
rect 3427 1976 4013 1984
rect 4267 1976 4413 1984
rect 4867 1976 5253 1984
rect 5507 1976 5553 1984
rect 247 1956 453 1964
rect 487 1956 933 1964
rect 1107 1956 1173 1964
rect 1447 1956 1573 1964
rect 1587 1956 1753 1964
rect 1767 1956 2753 1964
rect 2787 1956 3344 1964
rect 87 1936 473 1944
rect 1227 1936 1653 1944
rect 1667 1936 2453 1944
rect 2727 1936 3053 1944
rect 3187 1936 3313 1944
rect 3336 1944 3344 1956
rect 3487 1956 4553 1964
rect 4607 1956 4833 1964
rect 5107 1956 5593 1964
rect 3336 1936 3553 1944
rect 3887 1936 4053 1944
rect 4747 1936 5473 1944
rect 5487 1936 5693 1944
rect 27 1916 333 1924
rect 567 1916 1133 1924
rect 1187 1916 1293 1924
rect 1307 1916 1553 1924
rect 1707 1916 3133 1924
rect 3167 1916 3304 1924
rect 47 1896 93 1904
rect 107 1896 1693 1904
rect 1867 1896 2253 1904
rect 2267 1896 2393 1904
rect 2787 1896 2993 1904
rect 3007 1896 3233 1904
rect 3296 1904 3304 1916
rect 3667 1916 3993 1924
rect 4027 1916 4673 1924
rect 5227 1916 5453 1924
rect 3296 1896 3733 1904
rect 3847 1896 4653 1904
rect 4907 1896 5073 1904
rect 5327 1896 5373 1904
rect 5547 1896 5573 1904
rect 547 1876 673 1884
rect 767 1876 813 1884
rect 827 1876 1193 1884
rect 1347 1876 1533 1884
rect 1567 1876 1853 1884
rect 2027 1876 2173 1884
rect 2387 1876 2613 1884
rect 2627 1876 2993 1884
rect 3027 1876 3273 1884
rect 3347 1876 3833 1884
rect 3867 1876 4273 1884
rect 4627 1876 4933 1884
rect 4967 1876 5173 1884
rect 1127 1856 1253 1864
rect 1267 1856 1864 1864
rect 427 1836 564 1844
rect 556 1827 564 1836
rect 607 1836 633 1844
rect 767 1836 873 1844
rect 1127 1836 1173 1844
rect 1327 1836 1473 1844
rect 1707 1836 1833 1844
rect 1856 1844 1864 1856
rect 1967 1856 1993 1864
rect 2007 1856 2533 1864
rect 2587 1856 2833 1864
rect 2876 1856 3073 1864
rect 1856 1836 2273 1844
rect 527 1816 544 1824
rect 187 1796 353 1804
rect 456 1784 464 1793
rect 536 1787 544 1816
rect 807 1816 893 1824
rect 956 1816 1033 1824
rect 956 1807 964 1816
rect 1087 1816 1213 1824
rect 1447 1816 1744 1824
rect 587 1796 613 1804
rect 627 1796 753 1804
rect 827 1796 904 1804
rect 187 1776 464 1784
rect 787 1776 853 1784
rect 896 1784 904 1796
rect 987 1796 1313 1804
rect 1487 1796 1504 1804
rect 896 1776 993 1784
rect 1067 1776 1093 1784
rect 1247 1776 1313 1784
rect 67 1756 553 1764
rect 687 1756 773 1764
rect 827 1756 933 1764
rect 967 1756 1273 1764
rect 1416 1764 1424 1793
rect 1456 1784 1464 1793
rect 1456 1776 1473 1784
rect 1496 1784 1504 1796
rect 1527 1796 1593 1804
rect 1736 1804 1744 1816
rect 1856 1824 1864 1836
rect 2287 1836 2313 1844
rect 2347 1836 2793 1844
rect 2816 1836 2853 1844
rect 1827 1816 1864 1824
rect 1876 1816 1913 1824
rect 1776 1804 1784 1813
rect 1736 1796 1764 1804
rect 1776 1796 1833 1804
rect 1496 1776 1553 1784
rect 1756 1784 1764 1796
rect 1876 1804 1884 1816
rect 2167 1816 2324 1824
rect 1856 1796 1884 1804
rect 1756 1776 1813 1784
rect 1856 1784 1864 1796
rect 1907 1796 1933 1804
rect 1956 1796 2013 1804
rect 1847 1776 1864 1784
rect 1887 1776 1913 1784
rect 1956 1784 1964 1796
rect 2087 1796 2293 1804
rect 2316 1804 2324 1816
rect 2407 1816 2433 1824
rect 2496 1816 2673 1824
rect 2316 1796 2344 1804
rect 1947 1776 1964 1784
rect 2087 1776 2113 1784
rect 2247 1776 2313 1784
rect 2336 1784 2344 1796
rect 2387 1796 2453 1804
rect 2336 1776 2473 1784
rect 1416 1756 1533 1764
rect 1587 1756 2053 1764
rect 2407 1756 2433 1764
rect 2496 1764 2504 1816
rect 2787 1816 2804 1824
rect 2527 1796 2573 1804
rect 2727 1796 2773 1804
rect 2496 1756 2573 1764
rect 2596 1764 2604 1793
rect 2796 1787 2804 1816
rect 2667 1776 2704 1784
rect 2696 1767 2704 1776
rect 2596 1756 2633 1764
rect 2816 1764 2824 1836
rect 2876 1827 2884 1856
rect 3687 1856 3873 1864
rect 3987 1856 4113 1864
rect 4307 1856 4353 1864
rect 4787 1856 4893 1864
rect 5067 1856 5173 1864
rect 2987 1836 3033 1844
rect 3147 1836 3184 1844
rect 2847 1816 2864 1824
rect 2856 1804 2864 1816
rect 2936 1824 2944 1833
rect 2907 1816 2944 1824
rect 3027 1816 3153 1824
rect 2856 1796 2924 1804
rect 2916 1784 2924 1796
rect 2947 1796 3133 1804
rect 2916 1776 2973 1784
rect 3027 1776 3053 1784
rect 3107 1776 3153 1784
rect 3176 1784 3184 1836
rect 3327 1836 3613 1844
rect 3807 1836 4093 1844
rect 4247 1836 4313 1844
rect 4407 1836 4433 1844
rect 4467 1836 4713 1844
rect 4947 1836 4964 1844
rect 3236 1824 3244 1833
rect 3227 1816 3284 1824
rect 3276 1804 3284 1816
rect 3307 1816 3353 1824
rect 3447 1816 3533 1824
rect 3667 1816 3693 1824
rect 3727 1816 3744 1824
rect 3276 1796 3464 1804
rect 3456 1787 3464 1796
rect 3536 1796 3593 1804
rect 3176 1776 3213 1784
rect 3387 1776 3413 1784
rect 2816 1756 3053 1764
rect 3127 1756 3233 1764
rect 3347 1756 3393 1764
rect 3456 1756 3473 1764
rect 3516 1764 3524 1793
rect 3536 1787 3544 1796
rect 3736 1804 3744 1816
rect 3876 1816 3953 1824
rect 3876 1807 3884 1816
rect 4007 1816 4024 1824
rect 4016 1807 4024 1816
rect 4087 1816 4193 1824
rect 4207 1816 4264 1824
rect 3736 1796 3764 1804
rect 3487 1756 3524 1764
rect 3616 1764 3624 1793
rect 3696 1784 3704 1793
rect 3756 1787 3764 1796
rect 3927 1796 3973 1804
rect 4256 1804 4264 1816
rect 4287 1816 4473 1824
rect 4487 1816 4593 1824
rect 4707 1816 4793 1824
rect 4256 1796 4584 1804
rect 3696 1776 3724 1784
rect 3547 1756 3693 1764
rect 3716 1764 3724 1776
rect 3867 1776 3893 1784
rect 3907 1776 3984 1784
rect 3716 1756 3733 1764
rect 3787 1756 3953 1764
rect 447 1736 1013 1744
rect 1047 1736 1173 1744
rect 1707 1736 1873 1744
rect 2027 1736 2053 1744
rect 2367 1736 2473 1744
rect 2547 1736 2733 1744
rect 2767 1736 3673 1744
rect 3727 1736 3813 1744
rect 3827 1736 3933 1744
rect 3976 1744 3984 1776
rect 4007 1776 4293 1784
rect 4347 1776 4413 1784
rect 4576 1784 4584 1796
rect 4607 1796 4673 1804
rect 4816 1804 4824 1833
rect 4867 1816 4913 1824
rect 4807 1796 4824 1804
rect 4956 1787 4964 1836
rect 4987 1836 5033 1844
rect 5107 1836 5284 1844
rect 5007 1816 5233 1824
rect 5276 1807 5284 1836
rect 5547 1836 5573 1844
rect 5067 1796 5073 1804
rect 5127 1796 5144 1804
rect 4487 1776 4773 1784
rect 5076 1784 5084 1793
rect 5076 1776 5113 1784
rect 5136 1784 5144 1796
rect 5607 1796 5653 1804
rect 5136 1776 5273 1784
rect 4007 1756 4193 1764
rect 4327 1756 4413 1764
rect 4507 1756 5153 1764
rect 5396 1747 5404 1793
rect 3976 1736 4113 1744
rect 4147 1736 4273 1744
rect 4287 1736 4353 1744
rect 4527 1736 4553 1744
rect 4607 1736 4633 1744
rect 4667 1736 4913 1744
rect 5027 1736 5133 1744
rect 347 1716 573 1724
rect 707 1716 753 1724
rect 767 1716 833 1724
rect 887 1716 913 1724
rect 1147 1716 1473 1724
rect 1807 1716 2113 1724
rect 2327 1716 2613 1724
rect 2647 1716 2833 1724
rect 2887 1716 2913 1724
rect 2927 1716 3073 1724
rect 3147 1716 3253 1724
rect 3276 1716 3333 1724
rect 187 1696 233 1704
rect 427 1696 453 1704
rect 527 1696 653 1704
rect 687 1696 793 1704
rect 907 1696 2173 1704
rect 2187 1696 2453 1704
rect 2527 1696 2713 1704
rect 3276 1704 3284 1716
rect 3387 1716 3473 1724
rect 3507 1716 3653 1724
rect 3747 1716 3833 1724
rect 4207 1716 4733 1724
rect 4947 1716 5053 1724
rect 5267 1716 5353 1724
rect 5387 1716 5633 1724
rect 2987 1696 3284 1704
rect 3307 1696 3433 1704
rect 3527 1696 3573 1704
rect 3627 1696 3653 1704
rect 3827 1696 4233 1704
rect 4247 1696 4893 1704
rect 5127 1696 5433 1704
rect 5467 1696 5553 1704
rect 187 1676 693 1684
rect 827 1676 893 1684
rect 1027 1676 1113 1684
rect 1227 1676 2313 1684
rect 2336 1676 2753 1684
rect 127 1656 193 1664
rect 227 1656 293 1664
rect 307 1656 613 1664
rect 767 1656 1073 1664
rect 1107 1656 1433 1664
rect 1447 1656 1593 1664
rect 1807 1656 2193 1664
rect 2336 1664 2344 1676
rect 2787 1676 2933 1684
rect 3007 1676 3393 1684
rect 3447 1676 3533 1684
rect 3567 1676 3613 1684
rect 3747 1676 4673 1684
rect 4707 1676 4793 1684
rect 4867 1676 4893 1684
rect 4987 1676 5233 1684
rect 5507 1676 5673 1684
rect 2227 1656 2344 1664
rect 2747 1656 2853 1664
rect 3047 1656 3773 1664
rect 3807 1656 3833 1664
rect 3847 1656 4473 1664
rect 4627 1656 4673 1664
rect 4967 1656 5013 1664
rect 5047 1656 5393 1664
rect 56 1636 93 1644
rect 56 1567 64 1636
rect 207 1636 333 1644
rect 347 1636 633 1644
rect 647 1636 713 1644
rect 747 1636 793 1644
rect 907 1636 933 1644
rect 1007 1636 1033 1644
rect 1047 1636 1133 1644
rect 1147 1636 1173 1644
rect 1267 1636 1333 1644
rect 1567 1636 1673 1644
rect 1707 1636 1753 1644
rect 2567 1636 2713 1644
rect 2907 1636 3164 1644
rect 267 1616 973 1624
rect 1127 1616 1213 1624
rect 1307 1616 1393 1624
rect 1447 1616 1713 1624
rect 1867 1616 1933 1624
rect 2087 1616 2124 1624
rect 147 1596 253 1604
rect 447 1596 573 1604
rect 587 1596 704 1604
rect 87 1576 153 1584
rect 256 1584 264 1593
rect 256 1576 304 1584
rect 296 1567 304 1576
rect 376 1564 384 1593
rect 416 1576 473 1584
rect 367 1556 384 1564
rect 416 1564 424 1576
rect 527 1576 633 1584
rect 696 1584 704 1596
rect 1096 1604 1104 1613
rect 727 1596 1104 1604
rect 1327 1596 1373 1604
rect 1387 1596 1513 1604
rect 1587 1596 1613 1604
rect 1687 1596 1733 1604
rect 696 1576 833 1584
rect 927 1576 993 1584
rect 1207 1576 1233 1584
rect 1776 1584 1784 1593
rect 1516 1576 1784 1584
rect 407 1556 424 1564
rect 496 1564 504 1573
rect 447 1556 504 1564
rect 527 1556 693 1564
rect 847 1556 873 1564
rect 1087 1556 1213 1564
rect 1227 1556 1413 1564
rect 1516 1564 1524 1576
rect 1836 1584 1844 1613
rect 1907 1596 2013 1604
rect 1827 1576 1844 1584
rect 1887 1576 2104 1584
rect 2096 1567 2104 1576
rect 1507 1556 1524 1564
rect 1547 1556 1693 1564
rect 1707 1556 1753 1564
rect 1887 1556 1993 1564
rect 2007 1556 2073 1564
rect 2116 1564 2124 1616
rect 2667 1616 2793 1624
rect 2827 1616 2873 1624
rect 2947 1616 3113 1624
rect 2256 1587 2264 1613
rect 2447 1596 2464 1604
rect 2147 1576 2233 1584
rect 2116 1556 2144 1564
rect 2136 1547 2144 1556
rect 127 1536 453 1544
rect 467 1536 793 1544
rect 1067 1536 1413 1544
rect 1427 1536 1593 1544
rect 1647 1536 1833 1544
rect 2067 1536 2093 1544
rect 487 1516 513 1524
rect 707 1516 1333 1524
rect 1387 1516 1493 1524
rect 2007 1516 2113 1524
rect 2436 1524 2444 1573
rect 2456 1564 2464 1596
rect 2567 1596 2653 1604
rect 2847 1596 2953 1604
rect 3136 1604 3144 1613
rect 2967 1596 3144 1604
rect 2587 1576 2633 1584
rect 2816 1576 3053 1584
rect 2456 1556 2513 1564
rect 2816 1564 2824 1576
rect 3067 1576 3093 1584
rect 3156 1584 3164 1636
rect 3427 1636 3593 1644
rect 3627 1636 3753 1644
rect 3787 1636 3873 1644
rect 3887 1636 3893 1644
rect 3947 1636 3973 1644
rect 4127 1636 4293 1644
rect 4387 1636 4613 1644
rect 4767 1636 4793 1644
rect 4887 1636 5573 1644
rect 3267 1616 3293 1624
rect 3387 1616 3424 1624
rect 3207 1596 3284 1604
rect 3156 1576 3193 1584
rect 3276 1584 3284 1596
rect 3307 1596 3393 1604
rect 3416 1604 3424 1616
rect 3556 1616 3793 1624
rect 3416 1596 3433 1604
rect 3536 1587 3544 1613
rect 3556 1587 3564 1616
rect 3816 1616 3853 1624
rect 3627 1596 3653 1604
rect 3816 1604 3824 1616
rect 4067 1616 4133 1624
rect 4207 1616 4224 1624
rect 3776 1596 3824 1604
rect 3876 1596 3893 1604
rect 3276 1576 3473 1584
rect 2667 1556 2824 1564
rect 3007 1556 3353 1564
rect 3376 1556 3453 1564
rect 2467 1536 2593 1544
rect 2627 1536 2664 1544
rect 2436 1516 2633 1524
rect 2656 1524 2664 1536
rect 2687 1536 2753 1544
rect 3376 1544 3384 1556
rect 3467 1556 3513 1564
rect 3707 1556 3733 1564
rect 3747 1556 3753 1564
rect 3776 1547 3784 1596
rect 3876 1587 3884 1596
rect 4027 1596 4093 1604
rect 4176 1587 4184 1613
rect 4056 1576 4073 1584
rect 4056 1564 4064 1576
rect 4107 1576 4153 1584
rect 4216 1584 4224 1616
rect 4407 1616 4453 1624
rect 4727 1616 4933 1624
rect 4967 1616 5193 1624
rect 5307 1616 5333 1624
rect 5367 1616 5424 1624
rect 4236 1604 4244 1613
rect 4236 1596 4253 1604
rect 4287 1596 4353 1604
rect 4487 1596 4653 1604
rect 4767 1596 4813 1604
rect 5087 1596 5113 1604
rect 5207 1596 5313 1604
rect 5327 1596 5353 1604
rect 5376 1596 5393 1604
rect 4216 1576 4324 1584
rect 4316 1567 4324 1576
rect 4356 1576 4373 1584
rect 4356 1567 4364 1576
rect 4476 1584 4484 1593
rect 4467 1576 4484 1584
rect 4547 1576 4573 1584
rect 4856 1584 4864 1593
rect 4847 1576 4864 1584
rect 5107 1576 5133 1584
rect 5267 1576 5284 1584
rect 4027 1556 4064 1564
rect 4087 1556 4173 1564
rect 4387 1556 4713 1564
rect 4727 1556 4773 1564
rect 2907 1536 3384 1544
rect 3427 1536 3513 1544
rect 3527 1536 3533 1544
rect 3556 1536 3613 1544
rect 2656 1516 2733 1524
rect 2787 1516 2853 1524
rect 2907 1516 2973 1524
rect 3227 1516 3253 1524
rect 3556 1524 3564 1536
rect 3687 1536 3713 1544
rect 3796 1544 3804 1553
rect 3796 1536 3813 1544
rect 4216 1536 4713 1544
rect 3367 1516 3564 1524
rect 3587 1516 3873 1524
rect 4216 1524 4224 1536
rect 4747 1536 4913 1544
rect 4927 1536 5073 1544
rect 5176 1544 5184 1573
rect 5276 1564 5284 1576
rect 5376 1584 5384 1596
rect 5307 1576 5384 1584
rect 5416 1584 5424 1616
rect 5587 1616 5693 1624
rect 5416 1576 5553 1584
rect 5627 1576 5653 1584
rect 5667 1576 5693 1584
rect 5276 1556 5393 1564
rect 5447 1556 5493 1564
rect 5547 1556 5633 1564
rect 5687 1556 5733 1564
rect 5176 1536 5253 1544
rect 4007 1516 4224 1524
rect 4247 1516 4493 1524
rect 4507 1516 4593 1524
rect 4907 1516 5373 1524
rect 427 1496 833 1504
rect 947 1496 1293 1504
rect 2347 1496 2493 1504
rect 2547 1496 2873 1504
rect 2947 1496 3013 1504
rect 3036 1496 3833 1504
rect 27 1476 433 1484
rect 607 1476 993 1484
rect 1487 1476 1833 1484
rect 3036 1484 3044 1496
rect 3867 1496 4033 1504
rect 4047 1496 4113 1504
rect 4207 1496 4413 1504
rect 4487 1496 4553 1504
rect 4607 1496 4693 1504
rect 4727 1496 5513 1504
rect 5527 1496 5593 1504
rect 1847 1476 3044 1484
rect 3067 1476 3613 1484
rect 3827 1476 3933 1484
rect 4127 1476 4233 1484
rect 4727 1476 4833 1484
rect 4847 1476 5613 1484
rect 347 1456 413 1464
rect 447 1456 613 1464
rect 1867 1456 2104 1464
rect 647 1436 1913 1444
rect 2096 1444 2104 1456
rect 2127 1456 2713 1464
rect 2807 1456 2953 1464
rect 2967 1456 3133 1464
rect 3407 1456 3813 1464
rect 3847 1456 3973 1464
rect 3987 1456 5473 1464
rect 2096 1436 2213 1444
rect 2407 1436 2553 1444
rect 2607 1436 2833 1444
rect 2887 1436 2933 1444
rect 2987 1436 3013 1444
rect 3307 1436 3373 1444
rect 3507 1436 3533 1444
rect 3607 1436 4013 1444
rect 587 1416 633 1424
rect 1376 1416 2133 1424
rect 227 1396 473 1404
rect 1376 1404 1384 1416
rect 2427 1416 3153 1424
rect 3167 1416 3233 1424
rect 3247 1416 3373 1424
rect 3387 1416 3713 1424
rect 3827 1416 4253 1424
rect 5007 1416 5473 1424
rect 507 1396 1384 1404
rect 1547 1396 1793 1404
rect 2167 1396 3653 1404
rect 3667 1396 4033 1404
rect 4107 1396 4433 1404
rect 4447 1396 4453 1404
rect 4507 1396 4993 1404
rect 167 1376 173 1384
rect 187 1376 233 1384
rect 247 1376 273 1384
rect 327 1376 533 1384
rect 667 1376 1453 1384
rect 1727 1376 1973 1384
rect 2027 1376 2353 1384
rect 2456 1376 2573 1384
rect 356 1356 473 1364
rect 27 1336 53 1344
rect 87 1336 213 1344
rect 227 1336 273 1344
rect 287 1336 293 1344
rect 176 1304 184 1313
rect 167 1296 184 1304
rect 336 1304 344 1353
rect 356 1347 364 1356
rect 567 1356 593 1364
rect 607 1356 653 1364
rect 867 1356 913 1364
rect 927 1356 1193 1364
rect 1116 1347 1124 1356
rect 1267 1356 1273 1364
rect 1287 1356 1333 1364
rect 1527 1356 1553 1364
rect 1607 1356 1653 1364
rect 2456 1364 2464 1376
rect 2627 1376 2813 1384
rect 2867 1376 3353 1384
rect 3427 1376 3444 1384
rect 2327 1356 2464 1364
rect 2487 1356 2533 1364
rect 2556 1356 2773 1364
rect 376 1336 493 1344
rect 376 1327 384 1336
rect 807 1336 893 1344
rect 907 1336 933 1344
rect 1167 1336 1204 1344
rect 707 1316 733 1324
rect 887 1316 1013 1324
rect 1087 1316 1133 1324
rect 1196 1307 1204 1336
rect 1247 1336 1284 1344
rect 1276 1307 1284 1336
rect 1447 1336 1673 1344
rect 1687 1336 1733 1344
rect 1867 1336 1893 1344
rect 1907 1336 1933 1344
rect 336 1296 373 1304
rect 527 1296 553 1304
rect 567 1296 773 1304
rect 467 1276 493 1284
rect 507 1276 713 1284
rect 867 1276 953 1284
rect 987 1276 1093 1284
rect 1107 1276 1313 1284
rect 1416 1284 1424 1333
rect 1956 1327 1964 1353
rect 1487 1316 1553 1324
rect 1587 1316 1593 1324
rect 1607 1316 1653 1324
rect 2036 1324 2044 1353
rect 2067 1336 2104 1344
rect 2036 1316 2053 1324
rect 1527 1296 1613 1304
rect 1707 1296 1793 1304
rect 1876 1287 1884 1313
rect 1927 1296 2033 1304
rect 2096 1304 2104 1336
rect 2556 1344 2564 1356
rect 2847 1356 3424 1364
rect 3416 1347 3424 1356
rect 2447 1336 2564 1344
rect 2767 1336 2973 1344
rect 3247 1336 3313 1344
rect 3436 1344 3444 1376
rect 3467 1376 3493 1384
rect 3707 1376 3773 1384
rect 4167 1376 4213 1384
rect 4247 1376 4493 1384
rect 3487 1356 3573 1364
rect 3887 1356 4173 1364
rect 3436 1336 3473 1344
rect 3647 1336 3673 1344
rect 3696 1336 3733 1344
rect 2187 1316 2253 1324
rect 2447 1316 2533 1324
rect 2587 1316 2653 1324
rect 2676 1316 2913 1324
rect 2096 1296 2133 1304
rect 2207 1296 2273 1304
rect 2427 1296 2493 1304
rect 2676 1304 2684 1316
rect 2956 1316 3053 1324
rect 2607 1296 2684 1304
rect 2956 1304 2964 1316
rect 3107 1316 3133 1324
rect 3156 1316 3173 1324
rect 2787 1296 2964 1304
rect 1416 1276 1433 1284
rect 1887 1276 1913 1284
rect 2107 1276 2133 1284
rect 2147 1276 2293 1284
rect 2367 1276 2453 1284
rect 2487 1276 2553 1284
rect 2667 1276 2693 1284
rect 2956 1284 2964 1296
rect 2987 1296 3033 1304
rect 3156 1304 3164 1316
rect 3207 1316 3393 1324
rect 3536 1307 3544 1333
rect 3127 1296 3164 1304
rect 3196 1296 3233 1304
rect 2956 1276 2973 1284
rect 3027 1276 3093 1284
rect 207 1256 533 1264
rect 547 1256 613 1264
rect 647 1256 733 1264
rect 767 1256 793 1264
rect 907 1256 993 1264
rect 1127 1256 1293 1264
rect 2327 1256 2373 1264
rect 2447 1256 2473 1264
rect 2747 1256 2833 1264
rect 3196 1264 3204 1296
rect 3247 1296 3273 1304
rect 3387 1296 3433 1304
rect 3227 1276 3273 1284
rect 3347 1276 3413 1284
rect 3596 1284 3604 1333
rect 3636 1287 3644 1313
rect 3696 1304 3704 1336
rect 3787 1336 3873 1344
rect 3727 1316 3753 1324
rect 3807 1316 3993 1324
rect 4116 1307 4124 1333
rect 4136 1327 4144 1356
rect 4327 1356 4393 1364
rect 4907 1356 5253 1364
rect 5707 1356 5733 1364
rect 4156 1336 4233 1344
rect 3696 1296 3753 1304
rect 4156 1304 4164 1336
rect 4287 1336 4304 1344
rect 4187 1316 4213 1324
rect 4247 1316 4273 1324
rect 4296 1307 4304 1336
rect 4427 1336 4513 1344
rect 4767 1336 4913 1344
rect 5207 1336 5413 1344
rect 5667 1336 5693 1344
rect 4327 1316 4353 1324
rect 4456 1316 4533 1324
rect 4147 1296 4164 1304
rect 4367 1296 4413 1304
rect 4436 1287 4444 1313
rect 4456 1307 4464 1316
rect 4807 1316 4853 1324
rect 4867 1316 4973 1324
rect 5027 1316 5073 1324
rect 5527 1316 5733 1324
rect 4467 1296 4733 1304
rect 4747 1296 4773 1304
rect 4907 1296 4933 1304
rect 4967 1296 5053 1304
rect 5107 1296 5133 1304
rect 5247 1296 5593 1304
rect 5687 1296 5733 1304
rect 3447 1276 3604 1284
rect 3727 1276 3913 1284
rect 4327 1276 4393 1284
rect 4467 1276 4593 1284
rect 4647 1276 4693 1284
rect 4767 1276 4833 1284
rect 4887 1276 4973 1284
rect 5047 1276 5313 1284
rect 5407 1276 5433 1284
rect 3027 1256 3204 1264
rect 3227 1256 3473 1264
rect 3487 1256 4013 1264
rect 4027 1256 4053 1264
rect 4167 1256 4393 1264
rect 4667 1256 4833 1264
rect 5327 1256 5633 1264
rect 407 1236 473 1244
rect 627 1236 984 1244
rect 187 1216 433 1224
rect 447 1216 633 1224
rect 687 1216 753 1224
rect 827 1216 913 1224
rect 976 1224 984 1236
rect 1007 1236 1353 1244
rect 1507 1236 2513 1244
rect 2627 1236 2713 1244
rect 2727 1236 2793 1244
rect 2807 1236 2853 1244
rect 2947 1236 3133 1244
rect 3147 1236 3153 1244
rect 3267 1236 3313 1244
rect 3467 1236 3553 1244
rect 3607 1236 3813 1244
rect 3947 1236 4233 1244
rect 4447 1236 4573 1244
rect 4627 1236 5073 1244
rect 5347 1236 5413 1244
rect 976 1216 1153 1224
rect 1407 1216 2033 1224
rect 2707 1216 2813 1224
rect 3247 1216 3393 1224
rect 3527 1216 3553 1224
rect 3607 1216 3633 1224
rect 3647 1216 3793 1224
rect 3827 1216 4133 1224
rect 4527 1216 4693 1224
rect 5027 1216 5033 1224
rect 5047 1216 5173 1224
rect 5307 1216 5753 1224
rect 587 1196 1093 1204
rect 1176 1196 1413 1204
rect 1176 1184 1184 1196
rect 1787 1196 3973 1204
rect 3987 1196 4513 1204
rect 4827 1196 5144 1204
rect 327 1176 1184 1184
rect 1207 1176 1513 1184
rect 1527 1176 1553 1184
rect 1787 1176 1813 1184
rect 2007 1176 2373 1184
rect 2687 1176 2773 1184
rect 2807 1176 2893 1184
rect 3187 1176 3373 1184
rect 3487 1176 3513 1184
rect 3627 1176 3813 1184
rect 3947 1176 4093 1184
rect 4687 1176 4813 1184
rect 5136 1184 5144 1196
rect 5167 1196 5453 1204
rect 5467 1196 5533 1204
rect 5136 1176 5453 1184
rect 227 1156 613 1164
rect 627 1156 713 1164
rect 1087 1156 1273 1164
rect 1287 1156 1633 1164
rect 1687 1156 2733 1164
rect 2847 1156 2933 1164
rect 3067 1156 3133 1164
rect 3207 1156 3353 1164
rect 3387 1156 3773 1164
rect 3936 1156 3993 1164
rect 167 1136 273 1144
rect 307 1136 333 1144
rect 427 1136 453 1144
rect 476 1136 493 1144
rect 67 1116 113 1124
rect 87 1096 193 1104
rect 227 1096 253 1104
rect 287 1096 453 1104
rect 447 1076 464 1084
rect 456 1067 464 1076
rect 147 1056 413 1064
rect 476 1064 484 1136
rect 547 1136 593 1144
rect 667 1136 953 1144
rect 987 1136 1033 1144
rect 1387 1136 1593 1144
rect 1747 1136 1893 1144
rect 2007 1136 2073 1144
rect 2247 1136 2273 1144
rect 2547 1136 2713 1144
rect 2736 1136 3013 1144
rect 516 1116 704 1124
rect 496 1087 504 1113
rect 516 1107 524 1116
rect 696 1107 704 1116
rect 567 1096 653 1104
rect 716 1096 733 1104
rect 547 1076 593 1084
rect 607 1076 673 1084
rect 696 1067 704 1093
rect 716 1067 724 1096
rect 816 1096 853 1104
rect 476 1056 513 1064
rect 736 1064 744 1073
rect 736 1056 753 1064
rect 816 1064 824 1096
rect 927 1096 1113 1104
rect 1176 1104 1184 1133
rect 1207 1116 1224 1124
rect 1216 1104 1224 1116
rect 1247 1116 1353 1124
rect 1627 1116 1753 1124
rect 1807 1116 1853 1124
rect 2087 1116 2113 1124
rect 2136 1116 2333 1124
rect 1176 1096 1204 1104
rect 1216 1096 1293 1104
rect 1196 1087 1204 1096
rect 1476 1104 1484 1113
rect 1387 1096 1484 1104
rect 1867 1096 1973 1104
rect 1996 1096 2013 1104
rect 847 1076 933 1084
rect 987 1076 1013 1084
rect 1067 1076 1093 1084
rect 1247 1076 1293 1084
rect 1587 1076 1693 1084
rect 1996 1084 2004 1096
rect 2027 1096 2113 1104
rect 1887 1076 2004 1084
rect 2136 1084 2144 1116
rect 2347 1116 2453 1124
rect 2736 1124 2744 1136
rect 3047 1136 3124 1144
rect 2467 1116 2744 1124
rect 2767 1116 2833 1124
rect 2947 1116 3013 1124
rect 2227 1096 2333 1104
rect 2427 1096 2613 1104
rect 2727 1096 3033 1104
rect 2107 1076 2144 1084
rect 2247 1076 2393 1084
rect 2607 1076 2693 1084
rect 2767 1076 2913 1084
rect 3116 1084 3124 1136
rect 3167 1136 3313 1144
rect 3367 1136 3673 1144
rect 3936 1144 3944 1156
rect 4047 1156 4053 1164
rect 4067 1156 4133 1164
rect 4227 1156 4413 1164
rect 4427 1156 4873 1164
rect 4887 1156 5053 1164
rect 5107 1156 5153 1164
rect 5227 1156 5253 1164
rect 3796 1136 3944 1144
rect 3187 1116 3253 1124
rect 3287 1116 3333 1124
rect 3347 1116 3373 1124
rect 3416 1116 3433 1124
rect 3416 1104 3424 1116
rect 3587 1116 3633 1124
rect 3796 1124 3804 1136
rect 4007 1136 4033 1144
rect 4207 1136 4233 1144
rect 4267 1136 4304 1144
rect 3687 1116 3824 1124
rect 3147 1096 3424 1104
rect 2967 1076 3133 1084
rect 3436 1084 3444 1093
rect 3496 1087 3504 1113
rect 3816 1107 3824 1116
rect 3907 1116 4153 1124
rect 4116 1107 4124 1116
rect 4167 1116 4273 1124
rect 3267 1076 3444 1084
rect 3547 1076 3573 1084
rect 3616 1084 3624 1093
rect 3616 1076 3873 1084
rect 4047 1076 4173 1084
rect 4207 1076 4253 1084
rect 816 1056 973 1064
rect 1187 1056 1273 1064
rect 1867 1056 2073 1064
rect 2107 1056 2173 1064
rect 2207 1056 2293 1064
rect 2436 1064 2444 1073
rect 2427 1056 2444 1064
rect 2467 1056 2633 1064
rect 2747 1056 2853 1064
rect 2876 1056 3433 1064
rect 407 1036 533 1044
rect 567 1036 853 1044
rect 907 1036 1253 1044
rect 2147 1036 2253 1044
rect 2876 1044 2884 1056
rect 3647 1056 3693 1064
rect 3787 1056 3793 1064
rect 3807 1056 3953 1064
rect 4296 1064 4304 1136
rect 4547 1136 4573 1144
rect 4587 1136 4653 1144
rect 4787 1136 4873 1144
rect 4927 1136 4953 1144
rect 5027 1136 5113 1144
rect 5127 1136 5173 1144
rect 4387 1116 4933 1124
rect 5127 1116 5233 1124
rect 5647 1116 5713 1124
rect 4507 1096 4613 1104
rect 4736 1096 4773 1104
rect 4607 1076 4633 1084
rect 4736 1084 4744 1096
rect 4987 1096 5273 1104
rect 5567 1096 5653 1104
rect 5667 1096 5693 1104
rect 4687 1076 4744 1084
rect 5007 1076 5093 1084
rect 5107 1076 5193 1084
rect 5487 1076 5613 1084
rect 5627 1076 5693 1084
rect 4287 1056 4304 1064
rect 4507 1056 4553 1064
rect 4756 1064 4764 1073
rect 4687 1056 4764 1064
rect 2387 1036 2884 1044
rect 2947 1036 3253 1044
rect 3307 1036 3393 1044
rect 3407 1036 3753 1044
rect 3967 1036 4353 1044
rect 4367 1036 4893 1044
rect 307 1016 493 1024
rect 607 1016 833 1024
rect 1207 1016 1253 1024
rect 1667 1016 1933 1024
rect 2347 1016 2433 1024
rect 2567 1016 2653 1024
rect 2727 1016 2913 1024
rect 2967 1016 3213 1024
rect 3607 1016 3653 1024
rect 3767 1016 4053 1024
rect 4087 1016 5213 1024
rect 287 996 444 1004
rect 367 976 393 984
rect 436 984 444 996
rect 667 996 813 1004
rect 1027 996 1433 1004
rect 1547 996 3273 1004
rect 3367 996 3433 1004
rect 3727 996 3893 1004
rect 4367 996 4433 1004
rect 436 976 733 984
rect 787 976 1373 984
rect 1467 976 4493 984
rect 4507 976 4593 984
rect 247 956 593 964
rect 607 956 793 964
rect 807 956 873 964
rect 1047 956 1813 964
rect 2047 956 2513 964
rect 2547 956 2933 964
rect 3087 956 3173 964
rect 3207 956 3353 964
rect 3467 956 3773 964
rect 3847 956 4073 964
rect 4307 956 4993 964
rect 5007 956 5073 964
rect 347 936 493 944
rect 767 936 1293 944
rect 1347 936 2813 944
rect 2847 936 2973 944
rect 3067 936 3193 944
rect 3427 936 3753 944
rect 3776 936 3973 944
rect 2327 916 2533 924
rect 2647 916 2753 924
rect 3007 916 3093 924
rect 3227 916 3333 924
rect 3407 916 3493 924
rect 3627 916 3733 924
rect 3776 924 3784 936
rect 4027 936 4113 944
rect 4267 936 4313 944
rect 4447 936 4653 944
rect 4667 936 4713 944
rect 3747 916 3784 924
rect 4207 916 4833 924
rect 4847 916 4913 924
rect 4927 916 5033 924
rect 727 896 1373 904
rect 1747 896 1933 904
rect 2067 896 2193 904
rect 2207 896 3873 904
rect 3887 896 5013 904
rect 207 876 553 884
rect 567 876 573 884
rect 587 876 793 884
rect 807 876 913 884
rect 1127 876 1173 884
rect 1727 876 1773 884
rect 1907 876 1953 884
rect 1967 876 2313 884
rect 2347 876 2393 884
rect 2436 876 2553 884
rect 347 856 453 864
rect 467 856 493 864
rect 1107 856 1333 864
rect 1347 856 1453 864
rect 87 836 513 844
rect 647 836 684 844
rect 676 827 684 836
rect 707 836 1033 844
rect 1047 836 1113 844
rect 1187 836 1353 844
rect 1447 836 1473 844
rect 1616 844 1624 873
rect 1616 836 1633 844
rect 1656 844 1664 853
rect 1836 847 1844 873
rect 1867 856 2024 864
rect 1656 836 1713 844
rect 2016 844 2024 856
rect 2047 856 2073 864
rect 2227 856 2273 864
rect 2367 856 2393 864
rect 2436 864 2444 876
rect 2627 876 2653 884
rect 2767 876 3184 884
rect 2416 856 2444 864
rect 2016 836 2233 844
rect 2336 836 2373 844
rect 487 816 673 824
rect 727 816 753 824
rect 787 816 893 824
rect 907 816 1133 824
rect 1267 816 1433 824
rect 1467 816 1493 824
rect 1607 816 1753 824
rect 1927 816 1993 824
rect 2067 816 2093 824
rect 2207 816 2313 824
rect 427 796 493 804
rect 567 796 573 804
rect 587 796 613 804
rect 827 796 853 804
rect 947 796 1073 804
rect 1087 796 1233 804
rect 1247 796 1313 804
rect 1327 796 1393 804
rect 2167 796 2253 804
rect 2336 804 2344 836
rect 2416 824 2424 856
rect 2507 856 2544 864
rect 2447 836 2513 844
rect 2536 844 2544 856
rect 2587 856 2673 864
rect 2867 856 3053 864
rect 3176 864 3184 876
rect 3207 876 3704 884
rect 3176 856 3204 864
rect 3196 847 3204 856
rect 3247 856 3393 864
rect 3616 856 3633 864
rect 2536 836 2633 844
rect 2796 836 2953 844
rect 2796 827 2804 836
rect 3127 836 3153 844
rect 3387 836 3413 844
rect 3456 844 3464 853
rect 3436 836 3464 844
rect 2367 816 2424 824
rect 2507 816 2553 824
rect 2947 816 2973 824
rect 3027 816 3093 824
rect 3227 816 3313 824
rect 3436 824 3444 836
rect 3487 836 3573 844
rect 3616 844 3624 856
rect 3696 864 3704 876
rect 3727 876 3873 884
rect 4007 876 4093 884
rect 4107 876 4173 884
rect 4827 876 4864 884
rect 3696 856 4193 864
rect 4336 864 4344 873
rect 4856 867 4864 876
rect 4907 876 4953 884
rect 4336 856 4504 864
rect 3596 836 3624 844
rect 3387 816 3444 824
rect 3596 824 3604 836
rect 3687 836 3733 844
rect 3827 836 3953 844
rect 3967 836 4213 844
rect 4307 836 4473 844
rect 3467 816 3604 824
rect 3707 816 3753 824
rect 3927 816 3993 824
rect 4047 816 4133 824
rect 4207 816 4333 824
rect 4347 816 4393 824
rect 4496 824 4504 856
rect 4547 856 4604 864
rect 4596 844 4604 856
rect 4627 856 4673 864
rect 4967 856 5233 864
rect 5336 856 5673 864
rect 4596 836 4633 844
rect 4716 844 4724 853
rect 5336 847 5344 856
rect 4716 836 5173 844
rect 4496 816 4513 824
rect 2336 796 2493 804
rect 2527 796 2593 804
rect 2807 796 2833 804
rect 2887 796 3153 804
rect 3187 796 3553 804
rect 3607 796 3953 804
rect 3987 796 4173 804
rect 4187 796 4233 804
rect 4327 796 4393 804
rect 4507 796 4553 804
rect 4576 804 4584 833
rect 5056 827 5064 836
rect 5227 836 5253 844
rect 5547 836 5593 844
rect 5607 836 5673 844
rect 4607 816 4633 824
rect 4747 816 4793 824
rect 5327 816 5373 824
rect 5467 816 5493 824
rect 4576 796 4713 804
rect 4787 796 5053 804
rect 5247 796 5433 804
rect 367 776 393 784
rect 747 776 953 784
rect 967 776 993 784
rect 1007 776 1113 784
rect 1167 776 1273 784
rect 1787 776 1913 784
rect 2227 776 2433 784
rect 2447 776 2693 784
rect 2747 776 2773 784
rect 2787 776 3333 784
rect 3347 776 4773 784
rect 4807 776 4933 784
rect 5087 776 5473 784
rect 1107 756 1193 764
rect 1347 756 1933 764
rect 1987 756 2413 764
rect 2427 756 2713 764
rect 2727 756 2873 764
rect 2887 756 2893 764
rect 2907 756 3113 764
rect 3127 756 3213 764
rect 3267 756 3313 764
rect 3407 756 3913 764
rect 3927 756 3933 764
rect 3967 756 4373 764
rect 4587 756 4673 764
rect 4867 756 5013 764
rect 5027 756 5093 764
rect 5107 756 5153 764
rect 5167 756 5173 764
rect 5267 756 5353 764
rect 327 736 373 744
rect 467 736 1573 744
rect 1587 736 1813 744
rect 2307 736 2533 744
rect 2547 736 2713 744
rect 2727 736 2793 744
rect 2827 736 2913 744
rect 3247 736 3353 744
rect 3367 736 3413 744
rect 3527 736 3873 744
rect 4047 736 4113 744
rect 4387 736 4453 744
rect 367 716 1233 724
rect 1367 716 2133 724
rect 2147 716 2233 724
rect 2687 716 2893 724
rect 2947 716 3233 724
rect 547 696 633 704
rect 907 696 973 704
rect 1007 696 1073 704
rect 1527 696 1573 704
rect 1587 696 1873 704
rect 1887 696 2013 704
rect 2027 696 2373 704
rect 2407 696 2433 704
rect 2687 696 2953 704
rect 3067 696 3653 704
rect 3667 696 3793 704
rect 4087 696 4613 704
rect 4627 696 4733 704
rect 4847 696 5413 704
rect 5427 696 5533 704
rect 5547 696 5633 704
rect 547 676 573 684
rect 847 676 1013 684
rect 1027 676 1093 684
rect 1567 676 1833 684
rect 1847 676 2033 684
rect 2187 676 2213 684
rect 2227 676 2793 684
rect 3287 676 3693 684
rect 3727 676 3893 684
rect 3967 676 4293 684
rect 4507 676 4793 684
rect 5087 676 5113 684
rect 5147 676 5333 684
rect 5387 676 5433 684
rect 67 656 393 664
rect 447 656 1033 664
rect 1247 656 1413 664
rect 1427 656 1824 664
rect 107 636 133 644
rect 227 636 273 644
rect 407 636 453 644
rect 527 636 713 644
rect 887 636 1064 644
rect 1056 627 1064 636
rect 1107 636 1173 644
rect 1196 636 1333 644
rect 1196 627 1204 636
rect 1816 644 1824 656
rect 1907 656 1953 664
rect 1967 656 2113 664
rect 2367 656 2413 664
rect 2567 656 2753 664
rect 2827 656 3033 664
rect 3247 656 3393 664
rect 3447 656 3473 664
rect 3587 656 3853 664
rect 3947 656 3993 664
rect 4227 656 4293 664
rect 4487 656 4533 664
rect 5047 656 5153 664
rect 5207 656 5453 664
rect 5467 656 5513 664
rect 1816 636 1964 644
rect 1956 627 1964 636
rect 2067 636 2153 644
rect 2267 636 2393 644
rect 2656 636 2753 644
rect 2656 627 2664 636
rect 2847 636 2933 644
rect 3067 636 3164 644
rect 107 616 124 624
rect 116 604 124 616
rect 147 616 413 624
rect 547 616 693 624
rect 767 616 913 624
rect 1127 616 1193 624
rect 1247 616 1313 624
rect 1387 616 1653 624
rect 1687 616 1853 624
rect 2387 616 2553 624
rect 2707 616 2733 624
rect 2907 616 2933 624
rect 116 596 153 604
rect 267 596 333 604
rect 736 604 744 613
rect 727 596 744 604
rect 956 604 964 613
rect 956 596 1033 604
rect 1487 596 1584 604
rect 1287 576 1553 584
rect 1576 584 1584 596
rect 1607 596 1633 604
rect 1996 604 2004 613
rect 1996 596 2273 604
rect 2307 596 2333 604
rect 2856 604 2864 613
rect 2487 596 2864 604
rect 2927 596 2953 604
rect 2996 604 3004 633
rect 3027 616 3073 624
rect 3107 616 3133 624
rect 3156 624 3164 636
rect 3187 636 3273 644
rect 3707 636 3853 644
rect 3887 636 4164 644
rect 3156 616 3204 624
rect 2996 596 3013 604
rect 3196 604 3204 616
rect 3227 616 3253 624
rect 3307 616 3333 624
rect 3407 616 3493 624
rect 3607 616 3633 624
rect 3196 596 3213 604
rect 3247 596 3313 604
rect 3367 596 3513 604
rect 3656 604 3664 633
rect 4087 616 4133 624
rect 3627 596 3664 604
rect 3836 604 3844 613
rect 3747 596 3844 604
rect 3947 596 4093 604
rect 4156 604 4164 636
rect 4207 636 4233 644
rect 4347 636 4413 644
rect 4447 636 4513 644
rect 4607 636 4933 644
rect 5227 636 5253 644
rect 5356 636 5573 644
rect 5356 627 5364 636
rect 4187 616 4273 624
rect 4727 616 4833 624
rect 4887 616 5093 624
rect 5107 616 5193 624
rect 5207 616 5313 624
rect 4156 596 4173 604
rect 4367 596 4453 604
rect 4467 596 4913 604
rect 5007 596 5113 604
rect 5127 596 5393 604
rect 1676 584 1684 593
rect 1576 576 1684 584
rect 1747 576 1893 584
rect 2007 576 2933 584
rect 3207 576 3493 584
rect 3667 576 3753 584
rect 3907 576 3973 584
rect 4027 576 4053 584
rect 4227 576 4493 584
rect 4567 576 4593 584
rect 4607 576 4653 584
rect 87 556 473 564
rect 907 556 1393 564
rect 1447 556 1793 564
rect 1807 556 2393 564
rect 2407 556 3093 564
rect 3527 556 3593 564
rect 3787 556 4233 564
rect 307 536 353 544
rect 1687 536 1713 544
rect 2087 536 2153 544
rect 2187 536 2493 544
rect 2507 536 2573 544
rect 2607 536 3593 544
rect 3667 536 4533 544
rect 4547 536 4953 544
rect 4967 536 5013 544
rect 1907 516 2533 524
rect 2547 516 2613 524
rect 2807 516 2953 524
rect 3567 516 3733 524
rect 3767 516 4873 524
rect 327 496 393 504
rect 407 496 1573 504
rect 1587 496 2453 504
rect 2467 496 2593 504
rect 2647 496 2893 504
rect 2907 496 3133 504
rect 3927 496 4313 504
rect 4327 496 4633 504
rect 1887 476 3073 484
rect 3387 476 3633 484
rect 3767 476 3793 484
rect 5167 476 5193 484
rect 2047 456 2373 464
rect 2447 456 2753 464
rect 2887 456 2973 464
rect 2987 456 3133 464
rect 3227 456 4373 464
rect 4687 456 4733 464
rect 4747 456 4773 464
rect 667 436 733 444
rect 747 436 793 444
rect 807 436 833 444
rect 1207 436 1253 444
rect 1267 436 1513 444
rect 1527 436 1713 444
rect 1727 436 1773 444
rect 1787 436 2433 444
rect 2447 436 2933 444
rect 2947 436 3393 444
rect 3547 436 4033 444
rect 4047 436 4133 444
rect 4407 436 5153 444
rect 667 416 1693 424
rect 1707 416 3113 424
rect 3127 416 3193 424
rect 3467 416 4913 424
rect 487 396 573 404
rect 587 396 653 404
rect 707 396 973 404
rect 1567 396 1773 404
rect 1927 396 1973 404
rect 2147 396 2193 404
rect 2387 396 2884 404
rect 467 376 664 384
rect 87 356 493 364
rect 527 356 573 364
rect 656 364 664 376
rect 787 376 873 384
rect 1007 376 1073 384
rect 1387 376 1453 384
rect 1787 376 2073 384
rect 2156 376 2313 384
rect 656 356 1173 364
rect 1187 356 1284 364
rect 547 336 673 344
rect 696 336 973 344
rect 207 316 553 324
rect 696 324 704 336
rect 987 336 1013 344
rect 1067 336 1153 344
rect 1167 336 1184 344
rect 607 316 704 324
rect 927 316 973 324
rect 987 316 1093 324
rect 1107 316 1153 324
rect 1176 324 1184 336
rect 1207 336 1253 344
rect 1276 344 1284 356
rect 1367 356 1393 364
rect 1447 356 1473 364
rect 1487 356 1613 364
rect 1656 347 1664 373
rect 2156 367 2164 376
rect 2396 376 2413 384
rect 1747 356 1804 364
rect 1276 336 1333 344
rect 1467 336 1633 344
rect 1796 344 1804 356
rect 1827 356 1993 364
rect 2027 356 2053 364
rect 2067 356 2113 364
rect 1796 336 1853 344
rect 1867 336 1913 344
rect 1987 336 2053 344
rect 2147 336 2173 344
rect 2267 336 2373 344
rect 2396 344 2404 376
rect 2547 376 2813 384
rect 2847 376 2864 384
rect 2427 356 2473 364
rect 2527 356 2553 364
rect 2687 356 2733 364
rect 2767 356 2793 364
rect 2396 336 2453 344
rect 2607 336 2633 344
rect 2727 336 2773 344
rect 2836 344 2844 353
rect 2856 347 2864 376
rect 2807 336 2844 344
rect 2876 344 2884 396
rect 2967 396 3273 404
rect 3287 396 3693 404
rect 3707 396 4013 404
rect 4087 396 4413 404
rect 4427 396 4553 404
rect 4567 396 5613 404
rect 2896 367 2904 393
rect 2927 376 2973 384
rect 3147 376 3373 384
rect 3387 376 3413 384
rect 3607 376 3744 384
rect 3736 367 3744 376
rect 4727 376 4813 384
rect 5627 376 5693 384
rect 2947 356 3053 364
rect 3087 356 3093 364
rect 3107 356 3133 364
rect 3276 356 3353 364
rect 2876 336 2993 344
rect 3276 344 3284 356
rect 3427 356 3653 364
rect 3747 356 4013 364
rect 4147 356 4493 364
rect 4687 356 4733 364
rect 4887 356 4973 364
rect 4987 356 5053 364
rect 5067 356 5273 364
rect 5287 356 5313 364
rect 5587 356 5733 364
rect 3187 336 3284 344
rect 3307 336 3613 344
rect 3627 336 3673 344
rect 4867 336 5133 344
rect 1176 316 1213 324
rect 1327 316 1433 324
rect 1467 316 1493 324
rect 1607 316 1713 324
rect 1927 316 2353 324
rect 2367 316 2493 324
rect 2507 316 2533 324
rect 2547 316 2993 324
rect 3227 316 3284 324
rect 3276 307 3284 316
rect 3367 316 3913 324
rect 4227 316 4873 324
rect 5087 316 5453 324
rect 767 296 893 304
rect 907 296 933 304
rect 1687 296 2233 304
rect 2247 296 2573 304
rect 2587 296 3233 304
rect 3287 296 3333 304
rect 3347 296 3393 304
rect 3407 296 3624 304
rect 727 276 1833 284
rect 1847 276 2293 284
rect 2307 276 3573 284
rect 3616 284 3624 296
rect 3647 296 4033 304
rect 4807 296 4893 304
rect 4907 296 4973 304
rect 4987 296 5053 304
rect 3616 276 4713 284
rect 4727 276 4833 284
rect 967 256 1113 264
rect 1167 256 1913 264
rect 1947 256 1993 264
rect 2067 256 2253 264
rect 2347 256 2413 264
rect 2627 256 2653 264
rect 2667 256 2733 264
rect 2747 256 2793 264
rect 2987 256 3313 264
rect 3327 256 3453 264
rect 3467 256 3533 264
rect 627 236 884 244
rect 587 216 853 224
rect 876 224 884 236
rect 1127 236 2153 244
rect 2427 236 3093 244
rect 3147 236 3293 244
rect 4407 236 4553 244
rect 876 216 1113 224
rect 1407 216 1753 224
rect 2007 216 2473 224
rect 2567 216 2633 224
rect 2727 216 4433 224
rect 4447 216 4693 224
rect 647 196 773 204
rect 867 196 1293 204
rect 1667 196 1933 204
rect 2007 196 2513 204
rect 2527 196 2673 204
rect 2687 196 2793 204
rect 2887 196 2933 204
rect 2947 196 3233 204
rect 3256 196 3433 204
rect 207 176 713 184
rect 847 176 913 184
rect 947 176 1093 184
rect 1247 176 1953 184
rect 1987 176 2013 184
rect 2107 176 2193 184
rect 2287 176 2353 184
rect 2367 176 2413 184
rect 2487 176 2913 184
rect 3256 184 3264 196
rect 3607 196 3753 204
rect 3047 176 3264 184
rect 3307 176 3513 184
rect 3567 176 3733 184
rect 3867 176 4193 184
rect 4387 176 4413 184
rect 4487 176 4533 184
rect 4587 176 4653 184
rect 5267 176 5493 184
rect 627 156 693 164
rect 767 156 853 164
rect 876 156 953 164
rect 87 136 673 144
rect 876 144 884 156
rect 1676 156 1993 164
rect 847 136 884 144
rect 947 136 1073 144
rect 1127 136 1173 144
rect 1676 144 1684 156
rect 2087 156 2113 164
rect 2147 156 2173 164
rect 2447 156 2613 164
rect 2747 156 3013 164
rect 3067 156 3104 164
rect 1187 136 1684 144
rect 1707 136 1733 144
rect 1787 136 1873 144
rect 1927 136 2053 144
rect 2167 136 2213 144
rect 2227 136 2273 144
rect 2327 136 2653 144
rect 2667 136 2693 144
rect 2747 136 2833 144
rect 3007 136 3033 144
rect 3096 144 3104 156
rect 3127 156 3193 164
rect 3227 156 3353 164
rect 3387 156 3413 164
rect 3527 156 3573 164
rect 3587 156 3653 164
rect 3787 156 3893 164
rect 4327 156 4513 164
rect 4527 156 4613 164
rect 4687 156 4753 164
rect 4867 156 5113 164
rect 3096 136 3113 144
rect 3267 136 3333 144
rect 3667 136 4413 144
rect 4467 136 4493 144
rect 4696 136 4793 144
rect 467 116 573 124
rect 647 116 853 124
rect 867 116 3293 124
rect 3587 116 3633 124
rect 3707 116 3793 124
rect 3807 116 3933 124
rect 4696 124 4704 136
rect 4907 136 4933 144
rect 5627 136 5733 144
rect 4427 116 4704 124
rect 4727 116 4833 124
rect 4927 116 5033 124
rect 5087 116 5133 124
rect 5667 116 5693 124
rect 367 96 493 104
rect 507 96 633 104
rect 807 96 993 104
rect 2027 96 2133 104
rect 2147 96 2533 104
rect 2647 96 3573 104
rect 3687 96 3833 104
rect 4707 96 4733 104
rect 4827 96 4913 104
rect 5127 96 5173 104
rect 747 76 873 84
rect 1907 76 2113 84
rect 3087 76 3213 84
rect 3567 76 3593 84
rect 47 56 1233 64
rect 2767 56 3273 64
rect 3576 56 5093 64
rect 2267 36 3493 44
rect 3576 44 3584 56
rect 5107 56 5233 64
rect 3507 36 3584 44
rect 3607 36 4213 44
rect 3487 16 3633 24
rect 3727 16 3833 24
use NOR2X1  _944_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305106
transform 1 0 2030 0 -1 5050
box -12 -8 92 252
use NOR2X1  _945_
timestamp 1728305106
transform 1 0 1610 0 -1 5050
box -12 -8 92 252
use NOR2X1  _946_
timestamp 1728305106
transform -1 0 1890 0 -1 5050
box -12 -8 92 252
use NAND3X1  _947_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305047
transform 1 0 1930 0 -1 5050
box -12 -8 112 252
use AOI21X1  _948_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304211
transform 1 0 2250 0 1 4570
box -12 -8 112 252
use NAND2X1  _949_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304996
transform 1 0 3170 0 1 3610
box -12 -8 92 252
use INVX1  _950_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1749781103
transform -1 0 2790 0 1 2650
box -12 -8 72 252
use NOR2X1  _951_
timestamp 1728305106
transform 1 0 2590 0 -1 2650
box -12 -8 92 252
use NAND2X1  _952_
timestamp 1728304996
transform -1 0 2730 0 1 2650
box -12 -8 92 252
use NOR2X1  _953_
timestamp 1728305106
transform 1 0 3190 0 -1 2650
box -12 -8 92 252
use AND2X2  _954_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304163
transform 1 0 3270 0 -1 2650
box -12 -8 112 252
use INVX1  _955_
timestamp 1749781103
transform 1 0 2450 0 1 3130
box -12 -8 72 252
use INVX1  _956_
timestamp 1749781103
transform 1 0 1910 0 1 2650
box -12 -8 72 252
use NOR2X1  _957_
timestamp 1728305106
transform -1 0 2410 0 -1 2650
box -12 -8 92 252
use NAND3X1  _958_
timestamp 1728305047
transform 1 0 2310 0 1 2650
box -12 -8 112 252
use INVX1  _959_
timestamp 1749781103
transform 1 0 2070 0 -1 2650
box -12 -8 72 252
use INVX1  _960_
timestamp 1749781103
transform -1 0 2570 0 -1 3130
box -12 -8 72 252
use NAND3X1  _961_
timestamp 1728305047
transform 1 0 2450 0 1 2650
box -12 -8 112 252
use OAI21X1  _962_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305162
transform 1 0 2550 0 1 2650
box -12 -8 112 252
use NAND3X1  _963_
timestamp 1728305047
transform 1 0 3510 0 -1 3130
box -12 -8 112 252
use INVX1  _964_
timestamp 1749781103
transform 1 0 3650 0 1 2650
box -12 -8 72 252
use INVX4  _965_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304878
transform -1 0 1810 0 -1 5050
box -12 -8 92 252
use OR2X2  _966_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305284
transform 1 0 3330 0 1 2650
box -12 -8 112 252
use NOR2X1  _967_
timestamp 1728305106
transform 1 0 3470 0 1 2650
box -12 -8 92 252
use AND2X2  _968_
timestamp 1728304163
transform -1 0 2470 0 1 5050
box -12 -8 112 252
use INVX8  _969_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304916
transform -1 0 2550 0 -1 5530
box -12 -8 133 252
use INVX1  _970_
timestamp 1749781103
transform -1 0 1670 0 -1 4570
box -12 -8 72 252
use NAND3X1  _971_
timestamp 1728305047
transform -1 0 1490 0 -1 4570
box -12 -8 112 252
use NOR2X1  _972_
timestamp 1728305106
transform 1 0 1270 0 1 4570
box -12 -8 92 252
use NOR2X1  _973_
timestamp 1728305106
transform -1 0 1110 0 -1 4570
box -12 -8 92 252
use AND2X2  _974_
timestamp 1728304163
transform -1 0 1230 0 -1 4570
box -12 -8 112 252
use OR2X2  _975_
timestamp 1728305284
transform 1 0 2130 0 -1 5050
box -12 -8 112 252
use AOI21X1  _976_
timestamp 1728304211
transform -1 0 2250 0 1 4570
box -12 -8 112 252
use OAI21X1  _977_
timestamp 1728305162
transform -1 0 1350 0 -1 4570
box -12 -8 112 252
use NAND2X1  _978_
timestamp 1728304996
transform -1 0 1170 0 1 4090
box -12 -8 92 252
use NAND2X1  _979_
timestamp 1728304996
transform 1 0 2890 0 1 3130
box -12 -8 92 252
use OAI21X1  _980_
timestamp 1728305162
transform -1 0 2750 0 1 3130
box -12 -8 112 252
use OAI21X1  _981_
timestamp 1728305162
transform -1 0 2870 0 1 3130
box -12 -8 112 252
use NAND2X1  _982_
timestamp 1728304996
transform 1 0 2230 0 1 2650
box -12 -8 92 252
use AND2X2  _983_
timestamp 1728304163
transform 1 0 1990 0 1 3130
box -12 -8 112 252
use INVX1  _984_
timestamp 1749781103
transform 1 0 2230 0 1 3130
box -12 -8 72 252
use NAND3X1  _985_
timestamp 1728305047
transform -1 0 2210 0 1 3130
box -12 -8 112 252
use OAI21X1  _986_
timestamp 1728305162
transform 1 0 1650 0 1 3130
box -12 -8 112 252
use OAI21X1  _987_
timestamp 1728305162
transform -1 0 1630 0 1 3130
box -12 -8 112 252
use OAI21X1  _988_
timestamp 1728305162
transform 1 0 1690 0 1 2650
box -12 -8 112 252
use NAND3X1  _989_
timestamp 1728305047
transform 1 0 1930 0 -1 3130
box -12 -8 112 252
use OAI21X1  _990_
timestamp 1728305162
transform -1 0 2210 0 1 2650
box -12 -8 112 252
use NAND3X1  _991_
timestamp 1728305047
transform -1 0 2090 0 1 2650
box -12 -8 112 252
use OAI21X1  _992_
timestamp 1728305162
transform -1 0 1910 0 1 2650
box -12 -8 112 252
use OAI21X1  _993_
timestamp 1728305162
transform 1 0 2770 0 -1 3610
box -12 -8 112 252
use AND2X2  _994_
timestamp 1728304163
transform 1 0 1810 0 -1 3130
box -12 -8 112 252
use NAND2X1  _995_
timestamp 1728304996
transform -1 0 2270 0 -1 3130
box -12 -8 92 252
use OAI21X1  _996_
timestamp 1728305162
transform 1 0 2310 0 1 3130
box -12 -8 112 252
use NAND3X1  _997_
timestamp 1728305047
transform 1 0 2530 0 1 3130
box -12 -8 112 252
use OAI21X1  _998_
timestamp 1728305162
transform 1 0 2650 0 -1 3610
box -12 -8 112 252
use OAI21X1  _999_
timestamp 1728305162
transform -1 0 1690 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1000_
timestamp 1728305047
transform 1 0 2070 0 -1 3130
box -12 -8 112 252
use INVX1  _1001_
timestamp 1749781103
transform 1 0 2870 0 -1 3130
box -12 -8 72 252
use OAI21X1  _1002_
timestamp 1728305162
transform 1 0 2410 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1003_
timestamp 1728305047
transform -1 0 2370 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1004_
timestamp 1728305162
transform -1 0 1570 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1005_
timestamp 1728305162
transform 1 0 2970 0 1 3130
box -12 -8 112 252
use NOR2X1  _1006_
timestamp 1728305106
transform -1 0 2690 0 -1 3130
box -12 -8 92 252
use NAND3X1  _1007_
timestamp 1728305047
transform 1 0 3230 0 -1 3130
box -12 -8 112 252
use INVX1  _1008_
timestamp 1749781103
transform 1 0 3170 0 -1 3130
box -12 -8 72 252
use OAI21X1  _1009_
timestamp 1728305162
transform 1 0 3030 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1010_
timestamp 1728305047
transform 1 0 3370 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1011_
timestamp 1728305162
transform -1 0 3170 0 1 3130
box -12 -8 112 252
use OAI21X1  _1012_
timestamp 1728305162
transform 1 0 3230 0 1 2650
box -12 -8 112 252
use NOR3X1  _1013_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728303224
transform 1 0 2690 0 -1 3130
box -12 -8 192 252
use NAND3X1  _1014_
timestamp 1728305047
transform 1 0 2830 0 1 2650
box -12 -8 112 252
use OAI21X1  _1015_
timestamp 1728305162
transform -1 0 3030 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1016_
timestamp 1728305047
transform 1 0 2970 0 1 2650
box -12 -8 112 252
use OAI21X1  _1017_
timestamp 1728305162
transform 1 0 3090 0 1 2650
box -12 -8 112 252
use INVX1  _1018_
timestamp 1749781103
transform 1 0 610 0 -1 4090
box -12 -8 72 252
use NAND2X1  _1019_
timestamp 1728304996
transform 1 0 2050 0 1 4570
box -12 -8 92 252
use AOI21X1  _1020_
timestamp 1728304211
transform -1 0 2030 0 1 4570
box -12 -8 112 252
use NOR2X1  _1021_
timestamp 1728305106
transform -1 0 590 0 -1 4090
box -12 -8 92 252
use INVX1  _1022_
timestamp 1749781103
transform -1 0 670 0 1 4090
box -12 -8 72 252
use NOR2X1  _1023_
timestamp 1728305106
transform -1 0 590 0 1 4090
box -12 -8 92 252
use NAND2X1  _1024_
timestamp 1728304996
transform 1 0 930 0 -1 4570
box -12 -8 92 252
use INVX1  _1025_
timestamp 1749781103
transform -1 0 750 0 1 4090
box -12 -8 72 252
use NAND2X1  _1026_
timestamp 1728304996
transform -1 0 790 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1027_
timestamp 1728305162
transform 1 0 810 0 -1 4570
box -12 -8 112 252
use INVX1  _1028_
timestamp 1749781103
transform -1 0 570 0 -1 4570
box -12 -8 72 252
use OAI21X1  _1029_
timestamp 1728305162
transform -1 0 690 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1030_
timestamp 1728305047
transform -1 0 890 0 1 4570
box -12 -8 112 252
use NAND2X1  _1031_
timestamp 1728304996
transform -1 0 110 0 1 4570
box -12 -8 92 252
use NOR2X1  _1032_
timestamp 1728305106
transform 1 0 130 0 1 4570
box -12 -8 92 252
use INVX1  _1033_
timestamp 1749781103
transform -1 0 770 0 1 4570
box -12 -8 72 252
use NAND2X1  _1034_
timestamp 1728304996
transform -1 0 110 0 1 5050
box -12 -8 92 252
use OR2X2  _1035_
timestamp 1728305284
transform 1 0 130 0 1 5050
box -12 -8 112 252
use NAND2X1  _1036_
timestamp 1728304996
transform -1 0 330 0 1 5050
box -12 -8 92 252
use NOR2X1  _1037_
timestamp 1728305106
transform 1 0 350 0 1 5050
box -12 -8 92 252
use INVX1  _1038_
timestamp 1749781103
transform -1 0 890 0 -1 5530
box -12 -8 72 252
use OAI21X1  _1039_
timestamp 1728305162
transform -1 0 130 0 -1 5530
box -12 -8 112 252
use AND2X2  _1040_
timestamp 1728304163
transform -1 0 1250 0 1 4570
box -12 -8 112 252
use AND2X2  _1041_
timestamp 1728304163
transform 1 0 910 0 1 4570
box -12 -8 112 252
use NAND3X1  _1042_
timestamp 1728305047
transform -1 0 1130 0 1 4570
box -12 -8 112 252
use NAND2X1  _1043_
timestamp 1728304996
transform -1 0 230 0 -1 5530
box -12 -8 92 252
use NOR2X1  _1044_
timestamp 1728305106
transform 1 0 250 0 -1 5530
box -12 -8 92 252
use INVX1  _1045_
timestamp 1749781103
transform 1 0 1610 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1046_
timestamp 1728304996
transform 1 0 1310 0 -1 5530
box -12 -8 92 252
use NOR3X1  _1047_
timestamp 1728303224
transform 1 0 910 0 -1 5530
box -12 -8 192 252
use NAND2X1  _1048_
timestamp 1728304996
transform -1 0 1210 0 -1 5530
box -12 -8 92 252
use NAND2X1  _1049_
timestamp 1728304996
transform -1 0 1290 0 -1 5530
box -12 -8 92 252
use NOR2X1  _1050_
timestamp 1728305106
transform 1 0 1710 0 -1 5530
box -12 -8 92 252
use INVX1  _1051_
timestamp 1749781103
transform 1 0 1530 0 -1 5530
box -12 -8 72 252
use OAI21X1  _1052_
timestamp 1728305162
transform 1 0 1430 0 -1 5530
box -12 -8 112 252
use NAND2X1  _1053_
timestamp 1728304996
transform -1 0 1190 0 1 5050
box -12 -8 92 252
use OAI21X1  _1054_
timestamp 1728305162
transform 1 0 1230 0 1 5050
box -12 -8 112 252
use NOR2X1  _1055_
timestamp 1728305106
transform 1 0 1330 0 1 5050
box -12 -8 92 252
use INVX1  _1056_
timestamp 1749781103
transform 1 0 950 0 1 5050
box -12 -8 72 252
use NAND3X1  _1057_
timestamp 1728305047
transform 1 0 1010 0 1 5050
box -12 -8 112 252
use INVX1  _1058_
timestamp 1749781103
transform -1 0 890 0 -1 5050
box -12 -8 72 252
use OAI21X1  _1059_
timestamp 1728305162
transform -1 0 790 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1060_
timestamp 1728304996
transform -1 0 690 0 -1 5050
box -12 -8 92 252
use NOR2X1  _1061_
timestamp 1728305106
transform 1 0 490 0 -1 5050
box -12 -8 92 252
use INVX1  _1062_
timestamp 1749781103
transform -1 0 990 0 -1 5050
box -12 -8 72 252
use AOI21X1  _1063_
timestamp 1728304211
transform 1 0 990 0 -1 5050
box -12 -8 112 252
use NOR2X1  _1064_
timestamp 1728305106
transform -1 0 1610 0 -1 4570
box -12 -8 92 252
use DFFSR  _1065_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728387359
transform -1 0 3070 0 1 3610
box -12 -8 492 252
use DFFSR  _1066_
timestamp 1728387359
transform 1 0 810 0 1 3130
box -12 -8 492 252
use DFFSR  _1067_
timestamp 1728387359
transform -1 0 1670 0 1 2650
box -12 -8 492 252
use DFFSR  _1068_
timestamp 1728387359
transform -1 0 3350 0 -1 3610
box -12 -8 492 252
use DFFSR  _1069_
timestamp 1728387359
transform 1 0 950 0 -1 3130
box -12 -8 492 252
use DFFSR  _1070_
timestamp 1728387359
transform 1 0 3170 0 1 3130
box -12 -8 492 252
use DFFSR  _1071_
timestamp 1728387359
transform -1 0 3150 0 -1 2650
box -12 -8 492 252
use DFFSR  _1072_
timestamp 1728387359
transform 1 0 10 0 -1 4090
box -12 -8 492 252
use DFFSR  _1073_
timestamp 1728387359
transform 1 0 10 0 1 4090
box -12 -8 492 252
use DFFSR  _1074_
timestamp 1728387359
transform 1 0 10 0 -1 4570
box -12 -8 492 252
use DFFSR  _1075_
timestamp 1728387359
transform 1 0 210 0 1 4570
box -12 -8 492 252
use DFFSR  _1076_
timestamp 1728387359
transform 1 0 10 0 -1 5050
box -12 -8 492 252
use DFFSR  _1077_
timestamp 1728387359
transform 1 0 330 0 -1 5530
box -12 -8 492 252
use DFFSR  _1078_
timestamp 1728387359
transform 1 0 1790 0 -1 5530
box -12 -8 492 252
use DFFSR  _1079_
timestamp 1728387359
transform 1 0 1410 0 1 5050
box -12 -8 492 252
use DFFSR  _1080_
timestamp 1728387359
transform 1 0 430 0 1 5050
box -12 -8 492 252
use DFFSR  _1081_
timestamp 1728387359
transform -1 0 1570 0 -1 5050
box -12 -8 492 252
use DFFSR  _1082_
timestamp 1728387359
transform 1 0 1430 0 1 4570
box -12 -8 492 252
use DFFSR  _1083_
timestamp 1728387359
transform -1 0 2370 0 1 5050
box -12 -8 492 252
use INVX1  _1084_
timestamp 1749781103
transform 1 0 3710 0 1 2650
box -12 -8 72 252
use INVX1  _1085_
timestamp 1749781103
transform -1 0 2830 0 -1 4570
box -12 -8 72 252
use INVX1  _1086_
timestamp 1749781103
transform 1 0 3110 0 -1 5050
box -12 -8 72 252
use INVX1  _1087_
timestamp 1749781103
transform -1 0 3010 0 -1 4090
box -12 -8 72 252
use INVX1  _1088_
timestamp 1749781103
transform 1 0 3070 0 1 3610
box -12 -8 72 252
use INVX1  _1089_
timestamp 1749781103
transform -1 0 2690 0 -1 4090
box -12 -8 72 252
use NAND3X1  _1090_
timestamp 1728305047
transform -1 0 2790 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1091_
timestamp 1728304996
transform 1 0 3210 0 1 4570
box -12 -8 92 252
use NAND2X1  _1092_
timestamp 1728304996
transform -1 0 3950 0 -1 5530
box -12 -8 92 252
use INVX1  _1093_
timestamp 1749781103
transform -1 0 3590 0 -1 5050
box -12 -8 72 252
use NAND3X1  _1094_
timestamp 1728305047
transform -1 0 3730 0 1 4570
box -12 -8 112 252
use NOR2X1  _1095_
timestamp 1728305106
transform 1 0 3690 0 -1 4570
box -12 -8 92 252
use INVX1  _1096_
timestamp 1749781103
transform -1 0 3970 0 -1 5050
box -12 -8 72 252
use NAND3X1  _1097_
timestamp 1728305047
transform -1 0 3430 0 1 4570
box -12 -8 112 252
use NOR2X1  _1098_
timestamp 1728305106
transform -1 0 3770 0 1 5050
box -12 -8 92 252
use NOR2X1  _1099_
timestamp 1728305106
transform -1 0 3550 0 1 4570
box -12 -8 92 252
use NOR2X1  _1100_
timestamp 1728305106
transform -1 0 3550 0 -1 4570
box -12 -8 92 252
use INVX1  _1101_
timestamp 1749781103
transform 1 0 3790 0 1 5050
box -12 -8 72 252
use OAI21X1  _1102_
timestamp 1728305162
transform 1 0 3970 0 1 5050
box -12 -8 112 252
use NAND2X1  _1103_
timestamp 1728304996
transform -1 0 3950 0 1 5050
box -12 -8 92 252
use INVX1  _1104_
timestamp 1749781103
transform -1 0 3450 0 -1 4570
box -12 -8 72 252
use OAI22X1  _1105_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305200
transform 1 0 3250 0 -1 4570
box -12 -8 132 252
use INVX1  _1106_
timestamp 1749781103
transform 1 0 3970 0 -1 5530
box -12 -8 72 252
use INVX1  _1107_
timestamp 1749781103
transform -1 0 3870 0 -1 5530
box -12 -8 72 252
use OAI21X1  _1108_
timestamp 1728305162
transform 1 0 3690 0 -1 5530
box -12 -8 112 252
use OAI21X1  _1109_
timestamp 1728305162
transform -1 0 3670 0 -1 5530
box -12 -8 112 252
use INVX1  _1110_
timestamp 1749781103
transform 1 0 2810 0 -1 5530
box -12 -8 72 252
use AND2X2  _1111_
timestamp 1728304163
transform -1 0 3430 0 -1 5530
box -12 -8 112 252
use OR2X2  _1112_
timestamp 1728305284
transform -1 0 2990 0 -1 5050
box -12 -8 112 252
use INVX1  _1113_
timestamp 1749781103
transform -1 0 2810 0 1 4090
box -12 -8 72 252
use INVX1  _1114_
timestamp 1749781103
transform 1 0 3110 0 1 4570
box -12 -8 72 252
use OAI21X1  _1115_
timestamp 1728305162
transform -1 0 3110 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1116_
timestamp 1728304996
transform -1 0 2990 0 1 5050
box -12 -8 92 252
use NAND2X1  _1117_
timestamp 1728304996
transform -1 0 3090 0 1 5050
box -12 -8 92 252
use AOI21X1  _1118_
timestamp 1728304211
transform 1 0 2990 0 -1 5530
box -12 -8 112 252
use AOI21X1  _1119_
timestamp 1728304211
transform -1 0 3210 0 -1 5530
box -12 -8 112 252
use NAND2X1  _1120_
timestamp 1728304996
transform 1 0 2890 0 -1 5530
box -12 -8 92 252
use NAND2X1  _1121_
timestamp 1728304996
transform -1 0 3310 0 -1 5530
box -12 -8 92 252
use AND2X2  _1122_
timestamp 1728304163
transform -1 0 2890 0 1 5050
box -12 -8 112 252
use NAND2X1  _1123_
timestamp 1728304996
transform 1 0 3010 0 1 4570
box -12 -8 92 252
use NAND2X1  _1124_
timestamp 1728304996
transform 1 0 2910 0 1 4570
box -12 -8 92 252
use INVX1  _1125_
timestamp 1749781103
transform -1 0 1750 0 1 3610
box -12 -8 72 252
use OAI21X1  _1126_
timestamp 1728305162
transform 1 0 2810 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1127_
timestamp 1728304996
transform -1 0 2730 0 1 4090
box -12 -8 92 252
use NOR2X1  _1128_
timestamp 1728305106
transform 1 0 2550 0 1 4090
box -12 -8 92 252
use AOI21X1  _1129_
timestamp 1728304211
transform -1 0 2730 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1130_
timestamp 1728304996
transform 1 0 2050 0 -1 4090
box -12 -8 92 252
use INVX1  _1131_
timestamp 1749781103
transform -1 0 2030 0 1 4090
box -12 -8 72 252
use NOR2X1  _1132_
timestamp 1728305106
transform 1 0 1950 0 -1 4090
box -12 -8 92 252
use INVX1  _1133_
timestamp 1749781103
transform 1 0 750 0 1 4090
box -12 -8 72 252
use NOR2X1  _1134_
timestamp 1728305106
transform -1 0 930 0 1 4090
box -12 -8 92 252
use INVX1  _1135_
timestamp 1749781103
transform 1 0 930 0 -1 4090
box -12 -8 72 252
use AOI22X1  _1136_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304278
transform -1 0 1910 0 -1 4090
box -14 -8 132 252
use NAND2X1  _1137_
timestamp 1728304996
transform 1 0 2330 0 1 4090
box -12 -8 92 252
use OAI21X1  _1138_
timestamp 1728305162
transform -1 0 1950 0 1 4090
box -12 -8 112 252
use INVX1  _1139_
timestamp 1749781103
transform 1 0 2310 0 -1 5050
box -12 -8 72 252
use NAND3X1  _1140_
timestamp 1728305047
transform 1 0 2410 0 -1 5050
box -12 -8 112 252
use OAI21X1  _1141_
timestamp 1728305162
transform -1 0 2890 0 1 4570
box -12 -8 112 252
use AOI21X1  _1142_
timestamp 1728304211
transform 1 0 2690 0 1 4570
box -12 -8 112 252
use NAND3X1  _1143_
timestamp 1728305047
transform -1 0 2770 0 -1 5050
box -12 -8 112 252
use NAND3X1  _1144_
timestamp 1728305047
transform -1 0 2770 0 1 5050
box -12 -8 112 252
use INVX1  _1145_
timestamp 1749781103
transform 1 0 2130 0 -1 4090
box -12 -8 72 252
use AND2X2  _1146_
timestamp 1728304163
transform -1 0 2970 0 -1 4570
box -12 -8 112 252
use INVX1  _1147_
timestamp 1749781103
transform 1 0 1210 0 -1 4090
box -12 -8 72 252
use NOR2X1  _1148_
timestamp 1728305106
transform -1 0 1390 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1149_
timestamp 1728305106
transform -1 0 1470 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1150_
timestamp 1728305162
transform -1 0 1610 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1151_
timestamp 1728304996
transform 1 0 1350 0 1 3610
box -12 -8 92 252
use NAND2X1  _1152_
timestamp 1728304996
transform 1 0 1590 0 1 3610
box -12 -8 92 252
use NAND2X1  _1153_
timestamp 1728304996
transform -1 0 1350 0 1 3610
box -12 -8 92 252
use OAI21X1  _1154_
timestamp 1728305162
transform 1 0 970 0 1 4090
box -12 -8 112 252
use NAND3X1  _1155_
timestamp 1728305047
transform 1 0 1590 0 1 4090
box -12 -8 112 252
use AOI21X1  _1156_
timestamp 1728304211
transform 1 0 2290 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1157_
timestamp 1728305047
transform -1 0 2650 0 1 4570
box -12 -8 112 252
use OAI22X1  _1158_
timestamp 1728305200
transform -1 0 2670 0 -1 5050
box -12 -8 132 252
use AOI21X1  _1159_
timestamp 1728304211
transform 1 0 2770 0 -1 5050
box -12 -8 112 252
use INVX1  _1160_
timestamp 1749781103
transform -1 0 2470 0 1 3610
box -12 -8 72 252
use OAI21X1  _1161_
timestamp 1728305162
transform -1 0 3650 0 -1 4570
box -12 -8 112 252
use INVX1  _1162_
timestamp 1749781103
transform 1 0 3810 0 -1 3610
box -12 -8 72 252
use NAND2X1  _1163_
timestamp 1728304996
transform 1 0 3450 0 -1 4090
box -12 -8 92 252
use NAND2X1  _1164_
timestamp 1728304996
transform -1 0 3350 0 1 4090
box -12 -8 92 252
use AOI22X1  _1165_
timestamp 1728304278
transform 1 0 3110 0 -1 4570
box -14 -8 132 252
use OAI21X1  _1166_
timestamp 1728305162
transform -1 0 3090 0 -1 4570
box -12 -8 112 252
use NOR2X1  _1167_
timestamp 1728305106
transform 1 0 1010 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1168_
timestamp 1728305106
transform -1 0 850 0 -1 4090
box -12 -8 92 252
use INVX2  _1169_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1749781103
transform 1 0 5550 0 -1 1690
box -12 -8 72 252
use NAND2X1  _1170_
timestamp 1728304996
transform -1 0 390 0 -1 2650
box -12 -8 92 252
use INVX1  _1171_
timestamp 1749781103
transform 1 0 810 0 -1 3130
box -12 -8 72 252
use NAND2X1  _1172_
timestamp 1728304996
transform 1 0 410 0 -1 2650
box -12 -8 92 252
use NAND2X1  _1173_
timestamp 1728304996
transform -1 0 290 0 -1 2650
box -12 -8 92 252
use INVX1  _1174_
timestamp 1749781103
transform -1 0 90 0 1 2650
box -12 -8 72 252
use INVX2  _1175_
timestamp 1749781103
transform 1 0 1010 0 1 2650
box -12 -8 72 252
use NAND2X1  _1176_
timestamp 1728304996
transform -1 0 110 0 -1 3130
box -12 -8 92 252
use INVX2  _1177_
timestamp 1749781103
transform -1 0 4890 0 1 3130
box -12 -8 72 252
use NOR2X1  _1178_
timestamp 1728305106
transform 1 0 470 0 -1 3130
box -12 -8 92 252
use NOR2X1  _1179_
timestamp 1728305106
transform -1 0 210 0 -1 3130
box -12 -8 92 252
use OAI21X1  _1180_
timestamp 1728305162
transform -1 0 330 0 1 3130
box -12 -8 112 252
use OR2X2  _1181_
timestamp 1728305284
transform 1 0 110 0 1 3130
box -12 -8 112 252
use NAND2X1  _1182_
timestamp 1728304996
transform -1 0 110 0 -1 3610
box -12 -8 92 252
use INVX2  _1183_
timestamp 1749781103
transform 1 0 170 0 -1 2170
box -12 -8 72 252
use NAND2X1  _1184_
timestamp 1728304996
transform -1 0 330 0 1 2650
box -12 -8 92 252
use AND2X2  _1185_
timestamp 1728304163
transform 1 0 230 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1186_
timestamp 1728305162
transform -1 0 450 0 -1 3130
box -12 -8 112 252
use INVX1  _1187_
timestamp 1749781103
transform 1 0 890 0 -1 3130
box -12 -8 72 252
use NOR2X1  _1188_
timestamp 1728305106
transform -1 0 990 0 1 2650
box -12 -8 92 252
use OR2X2  _1189_
timestamp 1728305284
transform 1 0 470 0 1 3130
box -12 -8 112 252
use INVX1  _1190_
timestamp 1749781103
transform -1 0 90 0 1 3130
box -12 -8 72 252
use OAI21X1  _1191_
timestamp 1728305162
transform 1 0 350 0 1 3130
box -12 -8 112 252
use NAND3X1  _1192_
timestamp 1728305047
transform 1 0 590 0 1 3130
box -12 -8 112 252
use NAND3X1  _1193_
timestamp 1728305047
transform 1 0 590 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1194_
timestamp 1728304996
transform 1 0 490 0 -1 3610
box -12 -8 92 252
use OAI21X1  _1195_
timestamp 1728305162
transform 1 0 710 0 1 3130
box -12 -8 112 252
use NAND3X1  _1196_
timestamp 1728305047
transform 1 0 830 0 -1 3610
box -12 -8 112 252
use INVX1  _1197_
timestamp 1749781103
transform -1 0 70 0 1 3610
box -12 -8 72 252
use NAND2X1  _1198_
timestamp 1728304996
transform -1 0 330 0 -1 3610
box -12 -8 92 252
use NAND3X1  _1199_
timestamp 1728305047
transform -1 0 210 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1200_
timestamp 1728305047
transform -1 0 470 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1201_
timestamp 1728305047
transform 1 0 210 0 1 3610
box -12 -8 112 252
use NAND2X1  _1202_
timestamp 1728304996
transform -1 0 2530 0 1 4090
box -12 -8 92 252
use NAND2X1  _1203_
timestamp 1728304996
transform 1 0 2110 0 1 4090
box -12 -8 92 252
use NAND2X1  _1204_
timestamp 1728304996
transform -1 0 1810 0 1 4090
box -12 -8 92 252
use INVX1  _1205_
timestamp 1749781103
transform -1 0 1590 0 1 4090
box -12 -8 72 252
use NAND3X1  _1206_
timestamp 1728305047
transform -1 0 1530 0 1 4090
box -12 -8 112 252
use NOR2X1  _1207_
timestamp 1728305106
transform -1 0 930 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1208_
timestamp 1728305162
transform 1 0 1290 0 1 4090
box -12 -8 112 252
use NAND2X1  _1209_
timestamp 1728304996
transform -1 0 1250 0 1 4090
box -12 -8 92 252
use AND2X2  _1210_
timestamp 1728304163
transform -1 0 890 0 1 3610
box -12 -8 112 252
use NOR2X1  _1211_
timestamp 1728305106
transform 1 0 670 0 1 3610
box -12 -8 92 252
use NAND2X1  _1212_
timestamp 1728304996
transform 1 0 590 0 1 3610
box -12 -8 92 252
use AOI21X1  _1213_
timestamp 1728304211
transform 1 0 930 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1214_
timestamp 1728305047
transform 1 0 110 0 1 3610
box -12 -8 112 252
use NAND3X1  _1215_
timestamp 1728305047
transform 1 0 690 0 -1 3610
box -12 -8 112 252
use OR2X2  _1216_
timestamp 1728305284
transform -1 0 550 0 1 3610
box -12 -8 112 252
use AOI21X1  _1217_
timestamp 1728304211
transform 1 0 310 0 1 3610
box -12 -8 112 252
use INVX1  _1218_
timestamp 1749781103
transform -1 0 1110 0 -1 2650
box -12 -8 72 252
use NOR2X1  _1219_
timestamp 1728305106
transform -1 0 890 0 -1 2650
box -12 -8 92 252
use INVX2  _1220_
timestamp 1749781103
transform -1 0 5530 0 -1 1690
box -12 -8 72 252
use NOR2X1  _1221_
timestamp 1728305106
transform -1 0 630 0 -1 2170
box -12 -8 92 252
use NOR2X1  _1222_
timestamp 1728305106
transform 1 0 730 0 -1 2650
box -12 -8 92 252
use NAND2X1  _1223_
timestamp 1728304996
transform -1 0 650 0 1 2650
box -12 -8 92 252
use OAI21X1  _1224_
timestamp 1728305162
transform 1 0 130 0 1 2650
box -12 -8 112 252
use OAI21X1  _1225_
timestamp 1728305162
transform -1 0 430 0 1 2650
box -12 -8 112 252
use NOR2X1  _1226_
timestamp 1728305106
transform 1 0 610 0 -1 2650
box -12 -8 92 252
use NOR2X1  _1227_
timestamp 1728305106
transform -1 0 570 0 -1 2650
box -12 -8 92 252
use OAI21X1  _1228_
timestamp 1728305162
transform 1 0 470 0 1 2650
box -12 -8 112 252
use INVX4  _1229_
timestamp 1728304878
transform 1 0 4490 0 1 1210
box -12 -8 92 252
use INVX2  _1230_
timestamp 1749781103
transform -1 0 4030 0 1 2170
box -12 -8 72 252
use NOR2X1  _1231_
timestamp 1728305106
transform 1 0 3030 0 1 2170
box -12 -8 92 252
use INVX1  _1232_
timestamp 1749781103
transform -1 0 3070 0 -1 2170
box -12 -8 72 252
use NOR2X1  _1233_
timestamp 1728305106
transform -1 0 3010 0 1 2170
box -12 -8 92 252
use NOR2X1  _1234_
timestamp 1728305106
transform 1 0 2830 0 1 2170
box -12 -8 92 252
use OAI21X1  _1235_
timestamp 1728305162
transform 1 0 2390 0 1 2170
box -12 -8 112 252
use AOI21X1  _1236_
timestamp 1728304211
transform -1 0 2370 0 1 2170
box -12 -8 112 252
use INVX2  _1237_
timestamp 1749781103
transform -1 0 2510 0 1 1690
box -12 -8 72 252
use NAND2X1  _1238_
timestamp 1728304996
transform -1 0 2370 0 -1 2170
box -12 -8 92 252
use INVX1  _1239_
timestamp 1749781103
transform -1 0 5050 0 -1 730
box -12 -8 72 252
use NAND2X1  _1240_
timestamp 1728304996
transform 1 0 2730 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1241_
timestamp 1728304996
transform -1 0 2270 0 -1 2170
box -12 -8 92 252
use INVX1  _1242_
timestamp 1749781103
transform -1 0 1890 0 1 1210
box -12 -8 72 252
use NAND2X1  _1243_
timestamp 1728304996
transform -1 0 1990 0 1 1210
box -12 -8 92 252
use INVX2  _1244_
timestamp 1749781103
transform 1 0 5110 0 1 250
box -12 -8 72 252
use NAND2X1  _1245_
timestamp 1728304996
transform 1 0 1990 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1246_
timestamp 1728304996
transform -1 0 1970 0 -1 1690
box -12 -8 92 252
use NOR2X1  _1247_
timestamp 1728305106
transform -1 0 1950 0 -1 2170
box -12 -8 92 252
use AND2X2  _1248_
timestamp 1728304163
transform -1 0 2050 0 1 2170
box -12 -8 112 252
use INVX2  _1249_
timestamp 1749781103
transform -1 0 3190 0 1 2170
box -12 -8 72 252
use NAND2X1  _1250_
timestamp 1728304996
transform -1 0 2590 0 -1 2170
box -12 -8 92 252
use AND2X2  _1251_
timestamp 1728304163
transform -1 0 2610 0 1 2170
box -12 -8 112 252
use OAI21X1  _1252_
timestamp 1728305162
transform -1 0 2490 0 -1 2170
box -12 -8 112 252
use NOR2X1  _1253_
timestamp 1728305106
transform 1 0 1970 0 -1 2170
box -12 -8 92 252
use AOI21X1  _1254_
timestamp 1728304211
transform -1 0 2170 0 -1 2170
box -12 -8 112 252
use NOR2X1  _1255_
timestamp 1728305106
transform 1 0 2730 0 1 2170
box -12 -8 92 252
use NOR2X1  _1256_
timestamp 1728305106
transform -1 0 2710 0 1 2170
box -12 -8 92 252
use OAI21X1  _1257_
timestamp 1728305162
transform 1 0 2070 0 1 2170
box -12 -8 112 252
use AOI21X1  _1258_
timestamp 1728304211
transform 1 0 1630 0 1 2170
box -12 -8 112 252
use INVX2  _1259_
timestamp 1749781103
transform 1 0 2150 0 -1 2650
box -12 -8 72 252
use NOR2X1  _1260_
timestamp 1728305106
transform -1 0 650 0 -1 3130
box -12 -8 92 252
use NAND3X1  _1261_
timestamp 1728305047
transform 1 0 690 0 -1 3130
box -12 -8 112 252
use NAND2X1  _1262_
timestamp 1728304996
transform -1 0 1930 0 1 2170
box -12 -8 92 252
use OAI22X1  _1263_
timestamp 1728305200
transform -1 0 1890 0 -1 2650
box -12 -8 132 252
use NOR2X1  _1264_
timestamp 1728305106
transform -1 0 3910 0 -1 1690
box -12 -8 92 252
use AOI21X1  _1265_
timestamp 1728304211
transform 1 0 3950 0 -1 1690
box -12 -8 112 252
use NAND2X1  _1266_
timestamp 1728304996
transform 1 0 4250 0 -1 1210
box -12 -8 92 252
use INVX1  _1267_
timestamp 1749781103
transform -1 0 3910 0 1 1210
box -12 -8 72 252
use NAND3X1  _1268_
timestamp 1728305047
transform 1 0 4050 0 -1 1690
box -12 -8 112 252
use OAI21X1  _1269_
timestamp 1728305162
transform -1 0 3950 0 1 2170
box -12 -8 112 252
use INVX1  _1270_
timestamp 1749781103
transform 1 0 4050 0 1 1690
box -12 -8 72 252
use NOR2X1  _1271_
timestamp 1728305106
transform 1 0 4370 0 -1 1210
box -12 -8 92 252
use NAND3X1  _1272_
timestamp 1728305047
transform 1 0 4130 0 1 1210
box -12 -8 112 252
use INVX1  _1273_
timestamp 1749781103
transform -1 0 4470 0 -1 1690
box -12 -8 72 252
use NAND2X1  _1274_
timestamp 1728304996
transform 1 0 4190 0 1 1690
box -12 -8 92 252
use NAND3X1  _1275_
timestamp 1728305047
transform 1 0 3530 0 -1 2650
box -12 -8 112 252
use NAND3X1  _1276_
timestamp 1728305047
transform 1 0 3350 0 -1 4090
box -12 -8 112 252
use AOI22X1  _1277_
timestamp 1728304278
transform 1 0 3650 0 -1 3610
box -14 -8 132 252
use NAND3X1  _1278_
timestamp 1728305047
transform 1 0 3650 0 1 3130
box -12 -8 112 252
use INVX1  _1279_
timestamp 1749781103
transform -1 0 3710 0 -1 3130
box -12 -8 72 252
use OAI21X1  _1280_
timestamp 1728305162
transform -1 0 1730 0 -1 2650
box -12 -8 112 252
use NOR3X1  _1281_
timestamp 1728303224
transform 1 0 1070 0 -1 3610
box -12 -8 192 252
use OAI22X1  _1282_
timestamp 1728305200
transform -1 0 3550 0 -1 5530
box -12 -8 132 252
use NOR2X1  _1283_
timestamp 1728305106
transform 1 0 3130 0 1 5050
box -12 -8 92 252
use INVX1  _1284_
timestamp 1749781103
transform 1 0 3210 0 1 5050
box -12 -8 72 252
use OAI21X1  _1285_
timestamp 1728305162
transform -1 0 2030 0 -1 4570
box -12 -8 112 252
use NOR2X1  _1286_
timestamp 1728305106
transform 1 0 2030 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1287_
timestamp 1728305162
transform -1 0 1750 0 -1 4090
box -12 -8 112 252
use OAI22X1  _1288_
timestamp 1728305200
transform -1 0 1890 0 -1 4570
box -12 -8 132 252
use NAND2X1  _1289_
timestamp 1728304996
transform -1 0 1210 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1290_
timestamp 1728305162
transform 1 0 1670 0 -1 4570
box -12 -8 112 252
use AOI22X1  _1291_
timestamp 1728304278
transform -1 0 3430 0 1 5050
box -14 -8 132 252
use AOI22X1  _1292_
timestamp 1728304278
transform -1 0 3690 0 1 5050
box -14 -8 132 252
use OAI21X1  _1293_
timestamp 1728305162
transform 1 0 3470 0 1 5050
box -12 -8 112 252
use INVX1  _1294_
timestamp 1749781103
transform -1 0 3630 0 1 4570
box -12 -8 72 252
use NOR2X1  _1295_
timestamp 1728305106
transform 1 0 3410 0 -1 5050
box -12 -8 92 252
use AOI21X1  _1296_
timestamp 1728304211
transform -1 0 3390 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1297_
timestamp 1728304996
transform -1 0 3270 0 -1 5050
box -12 -8 92 252
use AOI22X1  _1298_
timestamp 1728304278
transform -1 0 3390 0 1 3610
box -14 -8 132 252
use NAND2X1  _1299_
timestamp 1728304996
transform 1 0 1230 0 -1 2650
box -12 -8 92 252
use OAI21X1  _1300_
timestamp 1728305162
transform 1 0 670 0 1 2650
box -12 -8 112 252
use OAI21X1  _1301_
timestamp 1728305162
transform -1 0 890 0 1 2650
box -12 -8 112 252
use NAND3X1  _1302_
timestamp 1728305047
transform -1 0 3310 0 -1 1690
box -12 -8 112 252
use OAI21X1  _1303_
timestamp 1728305162
transform 1 0 2230 0 1 1690
box -12 -8 112 252
use NAND2X1  _1304_
timestamp 1728304996
transform 1 0 2350 0 1 1690
box -12 -8 92 252
use NAND2X1  _1305_
timestamp 1728304996
transform 1 0 1130 0 -1 2650
box -12 -8 92 252
use NAND3X1  _1306_
timestamp 1728305047
transform 1 0 1090 0 1 2650
box -12 -8 112 252
use INVX1  _1307_
timestamp 1749781103
transform 1 0 1230 0 -1 2170
box -12 -8 72 252
use OAI21X1  _1308_
timestamp 1728305162
transform 1 0 2110 0 1 1690
box -12 -8 112 252
use NAND3X1  _1309_
timestamp 1728305047
transform -1 0 3830 0 -1 1690
box -12 -8 112 252
use NAND2X1  _1310_
timestamp 1728304996
transform -1 0 3710 0 -1 1690
box -12 -8 92 252
use AOI22X1  _1311_
timestamp 1728304278
transform 1 0 1470 0 -1 2170
box -14 -8 132 252
use NAND3X1  _1312_
timestamp 1728305047
transform 1 0 3390 0 1 1210
box -12 -8 112 252
use NOR3X1  _1313_
timestamp 1728303224
transform 1 0 3510 0 1 1210
box -12 -8 192 252
use OAI21X1  _1314_
timestamp 1728305162
transform -1 0 3690 0 -1 1210
box -12 -8 112 252
use NAND2X1  _1315_
timestamp 1728304996
transform 1 0 3490 0 -1 1210
box -12 -8 92 252
use OAI22X1  _1316_
timestamp 1728305200
transform 1 0 1730 0 -1 2170
box -12 -8 132 252
use AOI21X1  _1317_
timestamp 1728304211
transform 1 0 1610 0 -1 2170
box -12 -8 112 252
use NAND3X1  _1318_
timestamp 1728305047
transform -1 0 3810 0 1 1210
box -12 -8 112 252
use NAND2X1  _1319_
timestamp 1728304996
transform 1 0 3350 0 1 730
box -12 -8 92 252
use AND2X2  _1320_
timestamp 1728304163
transform -1 0 4010 0 -1 1210
box -12 -8 112 252
use NOR3X1  _1321_
timestamp 1728303224
transform -1 0 3890 0 -1 1210
box -12 -8 192 252
use AOI21X1  _1322_
timestamp 1728304211
transform 1 0 3150 0 1 1210
box -12 -8 112 252
use OAI21X1  _1323_
timestamp 1728305162
transform 1 0 3370 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1324_
timestamp 1728305162
transform 1 0 3270 0 1 1210
box -12 -8 112 252
use NOR2X1  _1325_
timestamp 1728305106
transform -1 0 4470 0 1 1210
box -12 -8 92 252
use AOI21X1  _1326_
timestamp 1728304211
transform 1 0 4150 0 -1 1690
box -12 -8 112 252
use NOR2X1  _1327_
timestamp 1728305106
transform 1 0 4610 0 -1 1690
box -12 -8 92 252
use AOI22X1  _1328_
timestamp 1728304278
transform 1 0 3290 0 1 1690
box -14 -8 132 252
use OAI21X1  _1329_
timestamp 1728305162
transform 1 0 3110 0 -1 2170
box -12 -8 112 252
use INVX1  _1330_
timestamp 1749781103
transform -1 0 3630 0 1 1690
box -12 -8 72 252
use OAI21X1  _1331_
timestamp 1728305162
transform 1 0 4870 0 -1 1210
box -12 -8 112 252
use NAND2X1  _1332_
timestamp 1728304996
transform 1 0 4910 0 -1 250
box -12 -8 92 252
use AOI22X1  _1333_
timestamp 1728304278
transform 1 0 3450 0 1 1690
box -14 -8 132 252
use NAND2X1  _1334_
timestamp 1728304996
transform -1 0 3290 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1335_
timestamp 1728304996
transform -1 0 3810 0 1 2170
box -12 -8 92 252
use INVX1  _1336_
timestamp 1749781103
transform -1 0 3410 0 1 2170
box -12 -8 72 252
use AOI22X1  _1337_
timestamp 1728304278
transform 1 0 3230 0 1 2170
box -14 -8 132 252
use AOI22X1  _1338_
timestamp 1728304278
transform 1 0 3350 0 -1 3610
box -14 -8 132 252
use NAND3X1  _1339_
timestamp 1728305047
transform 1 0 3510 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1340_
timestamp 1728304996
transform -1 0 2110 0 1 4090
box -12 -8 92 252
use OAI21X1  _1341_
timestamp 1728305162
transform 1 0 2230 0 1 4090
box -12 -8 112 252
use NOR2X1  _1342_
timestamp 1728305106
transform -1 0 2310 0 -1 5050
box -12 -8 92 252
use NAND3X1  _1343_
timestamp 1728305047
transform -1 0 2610 0 -1 4570
box -12 -8 112 252
use INVX1  _1344_
timestamp 1749781103
transform 1 0 2530 0 -1 4090
box -12 -8 72 252
use OAI21X1  _1345_
timestamp 1728305162
transform 1 0 2230 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1346_
timestamp 1728304996
transform 1 0 2330 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1347_
timestamp 1728305106
transform 1 0 2450 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1348_
timestamp 1728305106
transform -1 0 1350 0 1 250
box -12 -8 92 252
use NOR2X1  _1349_
timestamp 1728305106
transform -1 0 210 0 1 1210
box -12 -8 92 252
use NAND2X1  _1350_
timestamp 1728304996
transform -1 0 1430 0 1 250
box -12 -8 92 252
use INVX2  _1351_
timestamp 1749781103
transform 1 0 3270 0 1 250
box -12 -8 72 252
use INVX2  _1352_
timestamp 1749781103
transform 1 0 2590 0 -1 250
box -12 -8 72 252
use NOR2X1  _1353_
timestamp 1728305106
transform 1 0 2390 0 -1 250
box -12 -8 92 252
use AND2X2  _1354_
timestamp 1728304163
transform 1 0 2230 0 -1 730
box -12 -8 112 252
use AOI21X1  _1355_
timestamp 1728304211
transform 1 0 1470 0 1 250
box -12 -8 112 252
use NOR2X1  _1356_
timestamp 1728305106
transform -1 0 2230 0 -1 730
box -12 -8 92 252
use OAI21X1  _1357_
timestamp 1728305162
transform -1 0 2310 0 1 730
box -12 -8 112 252
use INVX1  _1358_
timestamp 1749781103
transform 1 0 2170 0 -1 1210
box -12 -8 72 252
use NAND3X1  _1359_
timestamp 1728305047
transform 1 0 1590 0 1 250
box -12 -8 112 252
use INVX1  _1360_
timestamp 1749781103
transform 1 0 1990 0 1 250
box -12 -8 72 252
use OAI21X1  _1361_
timestamp 1728305162
transform 1 0 2050 0 -1 730
box -12 -8 112 252
use INVX1  _1362_
timestamp 1749781103
transform 1 0 2110 0 1 730
box -12 -8 72 252
use INVX2  _1363_
timestamp 1749781103
transform 1 0 610 0 1 1690
box -12 -8 72 252
use INVX2  _1364_
timestamp 1749781103
transform -1 0 90 0 1 1210
box -12 -8 72 252
use INVX2  _1365_
timestamp 1749781103
transform -1 0 90 0 -1 1690
box -12 -8 72 252
use NAND3X1  _1366_
timestamp 1728305047
transform -1 0 450 0 -1 730
box -12 -8 112 252
use OAI21X1  _1367_
timestamp 1728305162
transform 1 0 1930 0 -1 730
box -12 -8 112 252
use INVX1  _1368_
timestamp 1749781103
transform -1 0 1770 0 1 250
box -12 -8 72 252
use NAND2X1  _1369_
timestamp 1728304996
transform 1 0 1790 0 1 250
box -12 -8 92 252
use NAND3X1  _1370_
timestamp 1728305047
transform -1 0 2470 0 -1 1210
box -12 -8 112 252
use AOI21X1  _1371_
timestamp 1728304211
transform 1 0 2250 0 -1 1210
box -12 -8 112 252
use AND2X2  _1372_
timestamp 1728304163
transform -1 0 2210 0 1 1210
box -12 -8 112 252
use NAND2X1  _1373_
timestamp 1728304996
transform -1 0 110 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1374_
timestamp 1728304996
transform -1 0 110 0 -1 2650
box -12 -8 92 252
use INVX1  _1375_
timestamp 1749781103
transform 1 0 130 0 -1 2650
box -12 -8 72 252
use NAND2X1  _1376_
timestamp 1728304996
transform -1 0 230 0 1 2170
box -12 -8 92 252
use OR2X2  _1377_
timestamp 1728305284
transform -1 0 130 0 1 2170
box -12 -8 112 252
use AOI22X1  _1378_
timestamp 1728304278
transform -1 0 150 0 -1 2170
box -14 -8 132 252
use OAI21X1  _1379_
timestamp 1728305162
transform 1 0 890 0 1 730
box -12 -8 112 252
use NAND2X1  _1380_
timestamp 1728304996
transform -1 0 1470 0 1 730
box -12 -8 92 252
use NAND2X1  _1381_
timestamp 1728304996
transform -1 0 950 0 -1 2170
box -12 -8 92 252
use INVX2  _1382_
timestamp 1749781103
transform -1 0 1210 0 -1 730
box -12 -8 72 252
use OAI21X1  _1383_
timestamp 1728305162
transform 1 0 770 0 1 730
box -12 -8 112 252
use NAND3X1  _1384_
timestamp 1728305047
transform -1 0 470 0 -1 1210
box -12 -8 112 252
use NAND2X1  _1385_
timestamp 1728304996
transform 1 0 830 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1386_
timestamp 1728304996
transform -1 0 1350 0 1 1690
box -12 -8 92 252
use OAI21X1  _1387_
timestamp 1728305162
transform 1 0 250 0 -1 1690
box -12 -8 112 252
use AOI21X1  _1388_
timestamp 1728304211
transform 1 0 610 0 -1 1690
box -12 -8 112 252
use NAND2X1  _1389_
timestamp 1728304996
transform -1 0 490 0 1 1210
box -12 -8 92 252
use NOR2X1  _1390_
timestamp 1728305106
transform -1 0 790 0 1 1690
box -12 -8 92 252
use NOR2X1  _1391_
timestamp 1728305106
transform 1 0 790 0 1 1690
box -12 -8 92 252
use NAND3X1  _1392_
timestamp 1728305047
transform -1 0 1010 0 1 1690
box -12 -8 112 252
use NOR2X1  _1393_
timestamp 1728305106
transform 1 0 770 0 -1 2170
box -12 -8 92 252
use AOI21X1  _1394_
timestamp 1728304211
transform -1 0 770 0 -1 2170
box -12 -8 112 252
use OAI21X1  _1395_
timestamp 1728305162
transform 1 0 450 0 -1 2170
box -12 -8 112 252
use OAI21X1  _1396_
timestamp 1728305162
transform -1 0 1350 0 -1 730
box -12 -8 112 252
use NAND3X1  _1397_
timestamp 1728305047
transform -1 0 1710 0 -1 730
box -12 -8 112 252
use NAND2X1  _1398_
timestamp 1728304996
transform -1 0 1610 0 -1 730
box -12 -8 92 252
use NAND2X1  _1399_
timestamp 1728304996
transform -1 0 1950 0 1 730
box -12 -8 92 252
use AND2X2  _1400_
timestamp 1728304163
transform 1 0 1990 0 1 730
box -12 -8 112 252
use NAND3X1  _1401_
timestamp 1728305047
transform -1 0 2090 0 1 1210
box -12 -8 112 252
use INVX2  _1402_
timestamp 1749781103
transform -1 0 2970 0 1 730
box -12 -8 72 252
use NOR2X1  _1403_
timestamp 1728305106
transform 1 0 2830 0 1 1210
box -12 -8 92 252
use NOR2X1  _1404_
timestamp 1728305106
transform 1 0 2790 0 1 730
box -12 -8 92 252
use OR2X2  _1405_
timestamp 1728305284
transform -1 0 2830 0 1 1210
box -12 -8 112 252
use NAND3X1  _1406_
timestamp 1728305047
transform 1 0 2250 0 1 1210
box -12 -8 112 252
use NOR2X1  _1407_
timestamp 1728305106
transform 1 0 570 0 1 2170
box -12 -8 92 252
use NOR2X1  _1408_
timestamp 1728305106
transform -1 0 570 0 1 2170
box -12 -8 92 252
use NAND2X1  _1409_
timestamp 1728304996
transform -1 0 290 0 1 1210
box -12 -8 92 252
use INVX1  _1410_
timestamp 1749781103
transform -1 0 870 0 -1 730
box -12 -8 72 252
use OAI21X1  _1411_
timestamp 1728305162
transform -1 0 450 0 -1 1690
box -12 -8 112 252
use NAND2X1  _1412_
timestamp 1728304996
transform -1 0 610 0 1 730
box -12 -8 92 252
use INVX1  _1413_
timestamp 1749781103
transform 1 0 610 0 1 730
box -12 -8 72 252
use NAND2X1  _1414_
timestamp 1728304996
transform 1 0 270 0 -1 2170
box -12 -8 92 252
use AOI21X1  _1415_
timestamp 1728304211
transform 1 0 350 0 -1 2170
box -12 -8 112 252
use AND2X2  _1416_
timestamp 1728304163
transform -1 0 1250 0 1 1690
box -12 -8 112 252
use NAND3X1  _1417_
timestamp 1728305047
transform 1 0 1010 0 1 1690
box -12 -8 112 252
use OAI22X1  _1418_
timestamp 1728305200
transform -1 0 2710 0 -1 1690
box -12 -8 132 252
use AOI21X1  _1419_
timestamp 1728304211
transform 1 0 2350 0 1 1210
box -12 -8 112 252
use NOR2X1  _1420_
timestamp 1728305106
transform -1 0 2730 0 1 1210
box -12 -8 92 252
use NAND2X1  _1421_
timestamp 1728304996
transform 1 0 2870 0 1 250
box -12 -8 92 252
use INVX2  _1422_
timestamp 1749781103
transform -1 0 3430 0 1 250
box -12 -8 72 252
use OAI21X1  _1423_
timestamp 1728305162
transform 1 0 3230 0 -1 730
box -12 -8 112 252
use OAI21X1  _1424_
timestamp 1728305162
transform 1 0 3110 0 -1 730
box -12 -8 112 252
use INVX1  _1425_
timestamp 1749781103
transform 1 0 2930 0 1 1210
box -12 -8 72 252
use OAI22X1  _1426_
timestamp 1728305200
transform 1 0 2870 0 -1 2170
box -12 -8 132 252
use INVX2  _1427_
timestamp 1749781103
transform -1 0 2250 0 1 2170
box -12 -8 72 252
use OAI21X1  _1428_
timestamp 1728305162
transform 1 0 3130 0 1 730
box -12 -8 112 252
use NAND3X1  _1429_
timestamp 1728305047
transform 1 0 2830 0 -1 1690
box -12 -8 112 252
use NAND2X1  _1430_
timestamp 1728304996
transform 1 0 3410 0 -1 1690
box -12 -8 92 252
use INVX1  _1431_
timestamp 1749781103
transform -1 0 3390 0 -1 1690
box -12 -8 72 252
use AOI22X1  _1432_
timestamp 1728304278
transform -1 0 2850 0 -1 2170
box -14 -8 132 252
use OAI21X1  _1433_
timestamp 1728305162
transform -1 0 2710 0 -1 2170
box -12 -8 112 252
use NAND2X1  _1434_
timestamp 1728304996
transform -1 0 3090 0 1 1690
box -12 -8 92 252
use NAND2X1  _1435_
timestamp 1728304996
transform 1 0 3210 0 1 1690
box -12 -8 92 252
use NAND2X1  _1436_
timestamp 1728304996
transform 1 0 3110 0 1 1690
box -12 -8 92 252
use OAI21X1  _1437_
timestamp 1728305162
transform 1 0 2650 0 1 1690
box -12 -8 112 252
use AOI21X1  _1438_
timestamp 1728304211
transform -1 0 2630 0 1 1690
box -12 -8 112 252
use NAND2X1  _1439_
timestamp 1728304996
transform -1 0 1870 0 1 730
box -12 -8 92 252
use NAND2X1  _1440_
timestamp 1728304996
transform -1 0 2150 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1441_
timestamp 1728304996
transform 1 0 1830 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1442_
timestamp 1728304996
transform 1 0 1690 0 1 730
box -12 -8 92 252
use NAND2X1  _1443_
timestamp 1728304996
transform 1 0 1730 0 -1 730
box -12 -8 92 252
use NAND2X1  _1444_
timestamp 1728304996
transform -1 0 1670 0 1 730
box -12 -8 92 252
use NOR2X1  _1445_
timestamp 1728305106
transform -1 0 1810 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1446_
timestamp 1728304996
transform 1 0 1910 0 1 1690
box -12 -8 92 252
use NAND2X1  _1447_
timestamp 1728304996
transform -1 0 950 0 1 2170
box -12 -8 92 252
use NAND2X1  _1448_
timestamp 1728304996
transform 1 0 1070 0 1 2170
box -12 -8 92 252
use NAND2X1  _1449_
timestamp 1728304996
transform -1 0 1050 0 1 2170
box -12 -8 92 252
use OAI21X1  _1450_
timestamp 1728305162
transform 1 0 1490 0 1 1690
box -12 -8 112 252
use AOI21X1  _1451_
timestamp 1728304211
transform -1 0 1470 0 1 1690
box -12 -8 112 252
use NOR2X1  _1452_
timestamp 1728305106
transform -1 0 330 0 1 2170
box -12 -8 92 252
use AOI21X1  _1453_
timestamp 1728304211
transform 1 0 350 0 1 2170
box -12 -8 112 252
use NAND3X1  _1454_
timestamp 1728305047
transform -1 0 1070 0 -1 2170
box -12 -8 112 252
use OAI21X1  _1455_
timestamp 1728305162
transform -1 0 1210 0 -1 2170
box -12 -8 112 252
use AOI21X1  _1456_
timestamp 1728304211
transform -1 0 1250 0 1 2170
box -12 -8 112 252
use OAI21X1  _1457_
timestamp 1728305162
transform 1 0 1950 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1458_
timestamp 1728305047
transform -1 0 2990 0 1 1690
box -12 -8 112 252
use OAI21X1  _1459_
timestamp 1728305162
transform 1 0 2790 0 1 1690
box -12 -8 112 252
use AOI21X1  _1460_
timestamp 1728304211
transform 1 0 1990 0 1 1690
box -12 -8 112 252
use OAI21X1  _1461_
timestamp 1728305162
transform 1 0 1510 0 1 2170
box -12 -8 112 252
use INVX1  _1462_
timestamp 1749781103
transform 1 0 650 0 1 2170
box -12 -8 72 252
use OAI21X1  _1463_
timestamp 1728305162
transform 1 0 1290 0 1 2170
box -12 -8 112 252
use NOR2X1  _1464_
timestamp 1728305106
transform -1 0 1470 0 1 2170
box -12 -8 92 252
use NAND3X1  _1465_
timestamp 1728305047
transform 1 0 750 0 1 2170
box -12 -8 112 252
use NAND2X1  _1466_
timestamp 1728304996
transform 1 0 1450 0 -1 2650
box -12 -8 92 252
use AND2X2  _1467_
timestamp 1728304163
transform 1 0 1350 0 -1 2650
box -12 -8 112 252
use NAND2X1  _1468_
timestamp 1728304996
transform -1 0 2550 0 1 4570
box -12 -8 92 252
use AOI21X1  _1469_
timestamp 1728304211
transform -1 0 2630 0 -1 3610
box -12 -8 112 252
use OAI21X1  _1470_
timestamp 1728305162
transform 1 0 1750 0 1 3610
box -12 -8 112 252
use NOR2X1  _1471_
timestamp 1728305106
transform 1 0 2390 0 1 4570
box -12 -8 92 252
use NOR2X1  _1472_
timestamp 1728305106
transform 1 0 2390 0 -1 4570
box -12 -8 92 252
use NAND3X1  _1473_
timestamp 1728305047
transform -1 0 2250 0 -1 4570
box -12 -8 112 252
use NOR2X1  _1474_
timestamp 1728305106
transform 1 0 1850 0 1 3610
box -12 -8 92 252
use OAI21X1  _1475_
timestamp 1728305162
transform -1 0 2030 0 -1 2650
box -12 -8 112 252
use AOI21X1  _1476_
timestamp 1728304211
transform 1 0 1530 0 -1 2650
box -12 -8 112 252
use AOI21X1  _1477_
timestamp 1728304211
transform -1 0 2550 0 -1 2650
box -12 -8 112 252
use AOI21X1  _1478_
timestamp 1728304211
transform 1 0 3550 0 1 2650
box -12 -8 112 252
use INVX8  _1479_
timestamp 1728304916
transform 1 0 2510 0 1 5050
box -12 -8 133 252
use INVX1  _1480_
timestamp 1749781103
transform -1 0 5170 0 -1 3130
box -12 -8 72 252
use NOR2X1  _1481_
timestamp 1728305106
transform -1 0 1970 0 1 3130
box -12 -8 92 252
use NOR2X1  _1482_
timestamp 1728305106
transform -1 0 2290 0 -1 2650
box -12 -8 92 252
use AND2X2  _1483_
timestamp 1728304163
transform 1 0 2050 0 -1 3610
box -12 -8 112 252
use NOR2X1  _1484_
timestamp 1728305106
transform -1 0 1270 0 1 3610
box -12 -8 92 252
use NOR2X1  _1485_
timestamp 1728305106
transform 1 0 1710 0 -1 3610
box -12 -8 92 252
use NAND3X1  _1486_
timestamp 1728305047
transform -1 0 1670 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1487_
timestamp 1728304996
transform 1 0 930 0 -1 2650
box -12 -8 92 252
use NOR2X1  _1488_
timestamp 1728305106
transform -1 0 1190 0 1 3610
box -12 -8 92 252
use NAND3X1  _1489_
timestamp 1728305047
transform 1 0 1310 0 1 3130
box -12 -8 112 252
use NOR2X1  _1490_
timestamp 1728305106
transform 1 0 1430 0 1 3130
box -12 -8 92 252
use NAND2X1  _1491_
timestamp 1728304996
transform -1 0 1470 0 -1 3610
box -12 -8 92 252
use NOR2X1  _1492_
timestamp 1728305106
transform -1 0 1570 0 -1 3610
box -12 -8 92 252
use INVX1  _1493_
timestamp 1749781103
transform 1 0 5230 0 -1 4570
box -12 -8 72 252
use OAI21X1  _1494_
timestamp 1728305162
transform 1 0 5050 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1495_
timestamp 1728305047
transform 1 0 5090 0 1 3130
box -12 -8 112 252
use NAND2X1  _1496_
timestamp 1728304996
transform 1 0 5170 0 -1 3610
box -12 -8 92 252
use NOR2X1  _1497_
timestamp 1728305106
transform -1 0 1790 0 -1 3130
box -12 -8 92 252
use NOR2X1  _1498_
timestamp 1728305106
transform -1 0 1850 0 1 3130
box -12 -8 92 252
use AND2X2  _1499_
timestamp 1728304163
transform 1 0 1810 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1500_
timestamp 1728305047
transform 1 0 2170 0 -1 3610
box -12 -8 112 252
use AND2X2  _1501_
timestamp 1728304163
transform 1 0 1270 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1502_
timestamp 1728305047
transform 1 0 2490 0 1 3610
box -12 -8 112 252
use NOR2X1  _1503_
timestamp 1728305106
transform 1 0 5350 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1504_
timestamp 1728305106
transform 1 0 4990 0 1 3130
box -12 -8 92 252
use INVX1  _1505_
timestamp 1749781103
transform -1 0 5190 0 1 2650
box -12 -8 72 252
use NAND2X1  _1506_
timestamp 1728304996
transform 1 0 4710 0 1 2650
box -12 -8 92 252
use NAND2X1  _1507_
timestamp 1728304996
transform -1 0 4990 0 1 2650
box -12 -8 92 252
use NAND2X1  _1508_
timestamp 1728304996
transform 1 0 4810 0 1 2650
box -12 -8 92 252
use NAND2X1  _1509_
timestamp 1728304996
transform -1 0 5010 0 -1 3130
box -12 -8 92 252
use OR2X2  _1510_
timestamp 1728305284
transform -1 0 4910 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1511_
timestamp 1728305047
transform -1 0 4790 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1512_
timestamp 1728305162
transform 1 0 4570 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1513_
timestamp 1728305162
transform 1 0 5010 0 1 2650
box -12 -8 112 252
use NOR2X1  _1514_
timestamp 1728305106
transform -1 0 5570 0 1 2170
box -12 -8 92 252
use INVX2  _1515_
timestamp 1749781103
transform 1 0 5650 0 1 5050
box -12 -8 72 252
use NOR2X1  _1516_
timestamp 1728305106
transform 1 0 5650 0 -1 2170
box -12 -8 92 252
use NOR2X1  _1517_
timestamp 1728305106
transform 1 0 5590 0 1 2170
box -12 -8 92 252
use NAND2X1  _1518_
timestamp 1728304996
transform 1 0 5510 0 -1 2650
box -12 -8 92 252
use OR2X2  _1519_
timestamp 1728305284
transform -1 0 5730 0 -1 2650
box -12 -8 112 252
use NAND3X1  _1520_
timestamp 1728305047
transform -1 0 5410 0 -1 2650
box -12 -8 112 252
use OAI21X1  _1521_
timestamp 1728305162
transform 1 0 5210 0 -1 2650
box -12 -8 112 252
use NAND3X1  _1522_
timestamp 1728305047
transform 1 0 1910 0 -1 3610
box -12 -8 112 252
use NOR2X1  _1523_
timestamp 1728305106
transform 1 0 2290 0 1 3610
box -12 -8 92 252
use NAND3X1  _1524_
timestamp 1728305047
transform -1 0 2250 0 1 3610
box -12 -8 112 252
use NAND3X1  _1525_
timestamp 1728305047
transform 1 0 1970 0 1 3610
box -12 -8 112 252
use NOR2X1  _1526_
timestamp 1728305106
transform -1 0 2150 0 1 3610
box -12 -8 92 252
use NAND2X1  _1527_
timestamp 1728304996
transform -1 0 2390 0 -1 3610
box -12 -8 92 252
use OR2X2  _1528_
timestamp 1728305284
transform 1 0 2390 0 -1 3610
box -12 -8 112 252
use INVX1  _1529_
timestamp 1749781103
transform -1 0 4970 0 -1 2170
box -12 -8 72 252
use OAI21X1  _1530_
timestamp 1728305162
transform -1 0 5470 0 1 2170
box -12 -8 112 252
use NOR2X1  _1531_
timestamp 1728305106
transform -1 0 5110 0 1 2170
box -12 -8 92 252
use NOR2X1  _1532_
timestamp 1728305106
transform -1 0 5170 0 -1 2170
box -12 -8 92 252
use NOR2X1  _1533_
timestamp 1728305106
transform 1 0 5150 0 1 2170
box -12 -8 92 252
use OR2X2  _1534_
timestamp 1728305284
transform -1 0 5510 0 -1 2170
box -12 -8 112 252
use NAND2X1  _1535_
timestamp 1728304996
transform 1 0 5550 0 -1 2170
box -12 -8 92 252
use NAND3X1  _1536_
timestamp 1728305047
transform -1 0 5410 0 -1 2170
box -12 -8 112 252
use OAI21X1  _1537_
timestamp 1728305162
transform 1 0 5210 0 -1 2170
box -12 -8 112 252
use NOR2X1  _1538_
timestamp 1728305106
transform 1 0 5390 0 1 730
box -12 -8 92 252
use NOR2X1  _1539_
timestamp 1728305106
transform -1 0 5110 0 1 730
box -12 -8 92 252
use OR2X2  _1540_
timestamp 1728305284
transform 1 0 5470 0 1 730
box -12 -8 112 252
use INVX1  _1541_
timestamp 1749781103
transform 1 0 5610 0 1 730
box -12 -8 72 252
use OAI21X1  _1542_
timestamp 1728305162
transform 1 0 5630 0 -1 5050
box -12 -8 112 252
use NAND3X1  _1543_
timestamp 1728305047
transform 1 0 5270 0 1 2170
box -12 -8 112 252
use NAND2X1  _1544_
timestamp 1728304996
transform -1 0 5690 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1545_
timestamp 1728304996
transform 1 0 5650 0 1 4090
box -12 -8 92 252
use OR2X2  _1546_
timestamp 1728305284
transform -1 0 5750 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1547_
timestamp 1728305047
transform -1 0 5390 0 1 730
box -12 -8 112 252
use OAI21X1  _1548_
timestamp 1728305162
transform 1 0 5170 0 -1 730
box -12 -8 112 252
use OAI21X1  _1549_
timestamp 1728305162
transform 1 0 5150 0 1 730
box -12 -8 112 252
use NAND2X1  _1550_
timestamp 1728304996
transform -1 0 4770 0 1 730
box -12 -8 92 252
use NAND2X1  _1551_
timestamp 1728304996
transform 1 0 4910 0 1 730
box -12 -8 92 252
use NAND2X1  _1552_
timestamp 1728304996
transform -1 0 4870 0 1 730
box -12 -8 92 252
use AND2X2  _1553_
timestamp 1728304163
transform 1 0 5510 0 -1 730
box -12 -8 112 252
use NOR2X1  _1554_
timestamp 1728305106
transform 1 0 5410 0 -1 730
box -12 -8 92 252
use OAI21X1  _1555_
timestamp 1728305162
transform -1 0 5390 0 -1 730
box -12 -8 112 252
use OAI21X1  _1556_
timestamp 1728305162
transform 1 0 5070 0 -1 730
box -12 -8 112 252
use NOR2X1  _1557_
timestamp 1728305106
transform 1 0 5630 0 -1 730
box -12 -8 92 252
use NOR2X1  _1558_
timestamp 1728305106
transform -1 0 4670 0 1 1210
box -12 -8 92 252
use INVX1  _1559_
timestamp 1749781103
transform 1 0 4690 0 1 1210
box -12 -8 72 252
use AOI22X1  _1560_
timestamp 1728304278
transform 1 0 5590 0 1 1210
box -14 -8 132 252
use NOR2X1  _1561_
timestamp 1728305106
transform -1 0 5170 0 -1 1210
box -12 -8 92 252
use NOR2X1  _1562_
timestamp 1728305106
transform -1 0 5070 0 -1 1210
box -12 -8 92 252
use NOR2X1  _1563_
timestamp 1728305106
transform 1 0 5130 0 1 1210
box -12 -8 92 252
use INVX1  _1564_
timestamp 1749781103
transform -1 0 5690 0 1 4570
box -12 -8 72 252
use OR2X2  _1565_
timestamp 1728305284
transform -1 0 5330 0 1 1210
box -12 -8 112 252
use OAI21X1  _1566_
timestamp 1728305162
transform -1 0 5110 0 1 1210
box -12 -8 112 252
use NAND3X1  _1567_
timestamp 1728305047
transform -1 0 4990 0 1 1210
box -12 -8 112 252
use OAI21X1  _1568_
timestamp 1728305162
transform 1 0 4770 0 1 1210
box -12 -8 112 252
use OAI21X1  _1569_
timestamp 1728305162
transform 1 0 5110 0 -1 1690
box -12 -8 112 252
use NOR2X1  _1570_
timestamp 1728305106
transform -1 0 4990 0 -1 1690
box -12 -8 92 252
use NOR2X1  _1571_
timestamp 1728305106
transform 1 0 5010 0 -1 1690
box -12 -8 92 252
use NOR2X1  _1572_
timestamp 1728305106
transform 1 0 5350 0 -1 1690
box -12 -8 92 252
use INVX1  _1573_
timestamp 1749781103
transform 1 0 5430 0 -1 2650
box -12 -8 72 252
use OR2X2  _1574_
timestamp 1728305284
transform -1 0 5450 0 1 1210
box -12 -8 112 252
use OAI21X1  _1575_
timestamp 1728305162
transform -1 0 5330 0 -1 1690
box -12 -8 112 252
use NAND3X1  _1576_
timestamp 1728305047
transform -1 0 5090 0 -1 2170
box -12 -8 112 252
use OAI21X1  _1577_
timestamp 1728305162
transform 1 0 4310 0 -1 2170
box -12 -8 112 252
use NAND3X1  _1578_
timestamp 1728305047
transform -1 0 5570 0 1 1210
box -12 -8 112 252
use NAND2X1  _1579_
timestamp 1728304996
transform -1 0 4790 0 -1 1690
box -12 -8 92 252
use NOR2X1  _1580_
timestamp 1728305106
transform 1 0 4810 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1581_
timestamp 1728304996
transform -1 0 4970 0 1 1690
box -12 -8 92 252
use AOI21X1  _1582_
timestamp 1728304211
transform -1 0 5090 0 1 1690
box -12 -8 112 252
use OAI21X1  _1583_
timestamp 1728305162
transform -1 0 5210 0 1 1690
box -12 -8 112 252
use OR2X2  _1584_
timestamp 1728305284
transform -1 0 4090 0 -1 2170
box -12 -8 112 252
use NAND2X1  _1585_
timestamp 1728304996
transform 1 0 4090 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1586_
timestamp 1728304996
transform -1 0 3950 0 -1 2170
box -12 -8 92 252
use NOR2X1  _1587_
timestamp 1728305106
transform 1 0 3410 0 -1 250
box -12 -8 92 252
use NAND3X1  _1588_
timestamp 1728305047
transform -1 0 3090 0 1 250
box -12 -8 112 252
use NAND3X1  _1589_
timestamp 1728305047
transform 1 0 1810 0 -1 730
box -12 -8 112 252
use OAI21X1  _1590_
timestamp 1728305162
transform 1 0 2990 0 -1 730
box -12 -8 112 252
use NAND2X1  _1591_
timestamp 1728304996
transform -1 0 790 0 1 250
box -12 -8 92 252
use AOI21X1  _1592_
timestamp 1728304211
transform 1 0 1390 0 -1 730
box -12 -8 112 252
use NAND3X1  _1593_
timestamp 1728305047
transform 1 0 1470 0 1 730
box -12 -8 112 252
use AND2X2  _1594_
timestamp 1728304163
transform 1 0 3250 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1595_
timestamp 1728305047
transform 1 0 3110 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1596_
timestamp 1728305162
transform -1 0 3110 0 1 730
box -12 -8 112 252
use NAND2X1  _1597_
timestamp 1728304996
transform -1 0 3670 0 -1 730
box -12 -8 92 252
use NAND2X1  _1598_
timestamp 1728304996
transform 1 0 250 0 -1 730
box -12 -8 92 252
use INVX2  _1599_
timestamp 1749781103
transform 1 0 490 0 -1 250
box -12 -8 72 252
use NAND2X1  _1600_
timestamp 1728304996
transform -1 0 130 0 -1 730
box -12 -8 92 252
use NAND2X1  _1601_
timestamp 1728304996
transform -1 0 210 0 -1 730
box -12 -8 92 252
use AND2X2  _1602_
timestamp 1728304163
transform 1 0 3790 0 1 730
box -12 -8 112 252
use NOR2X1  _1603_
timestamp 1728305106
transform 1 0 670 0 1 730
box -12 -8 92 252
use INVX1  _1604_
timestamp 1749781103
transform 1 0 1150 0 -1 250
box -12 -8 72 252
use NOR2X1  _1605_
timestamp 1728305106
transform 1 0 550 0 -1 730
box -12 -8 92 252
use OAI21X1  _1606_
timestamp 1728305162
transform 1 0 670 0 -1 730
box -12 -8 112 252
use OAI21X1  _1607_
timestamp 1728305162
transform 1 0 450 0 -1 730
box -12 -8 112 252
use INVX1  _1608_
timestamp 1749781103
transform -1 0 1110 0 -1 250
box -12 -8 72 252
use NOR2X1  _1609_
timestamp 1728305106
transform -1 0 870 0 1 250
box -12 -8 92 252
use OAI21X1  _1610_
timestamp 1728305162
transform 1 0 910 0 -1 250
box -12 -8 112 252
use OAI21X1  _1611_
timestamp 1728305162
transform 1 0 770 0 -1 250
box -12 -8 112 252
use NAND2X1  _1612_
timestamp 1728304996
transform 1 0 590 0 -1 250
box -12 -8 92 252
use OAI21X1  _1613_
timestamp 1728305162
transform -1 0 770 0 -1 250
box -12 -8 112 252
use NOR2X1  _1614_
timestamp 1728305106
transform -1 0 990 0 1 250
box -12 -8 92 252
use INVX1  _1615_
timestamp 1749781103
transform 1 0 1110 0 1 250
box -12 -8 72 252
use OAI21X1  _1616_
timestamp 1728305162
transform 1 0 1030 0 -1 730
box -12 -8 112 252
use NAND3X1  _1617_
timestamp 1728305047
transform -1 0 1110 0 1 250
box -12 -8 112 252
use OAI21X1  _1618_
timestamp 1728305162
transform 1 0 890 0 -1 730
box -12 -8 112 252
use NAND2X1  _1619_
timestamp 1728304996
transform -1 0 710 0 1 250
box -12 -8 92 252
use OAI21X1  _1620_
timestamp 1728305162
transform -1 0 610 0 1 250
box -12 -8 112 252
use NOR2X1  _1621_
timestamp 1728305106
transform -1 0 1270 0 1 250
box -12 -8 92 252
use NOR2X1  _1622_
timestamp 1728305106
transform -1 0 2010 0 -1 250
box -12 -8 92 252
use OAI21X1  _1623_
timestamp 1728305162
transform -1 0 2250 0 -1 250
box -12 -8 112 252
use OAI21X1  _1624_
timestamp 1728305162
transform 1 0 2030 0 -1 250
box -12 -8 112 252
use NAND2X1  _1625_
timestamp 1728304996
transform -1 0 1910 0 -1 250
box -12 -8 92 252
use OAI21X1  _1626_
timestamp 1728305162
transform 1 0 1710 0 -1 250
box -12 -8 112 252
use AOI21X1  _1627_
timestamp 1728304211
transform 1 0 2490 0 -1 250
box -12 -8 112 252
use NAND2X1  _1628_
timestamp 1728304996
transform -1 0 3590 0 -1 250
box -12 -8 92 252
use NAND2X1  _1629_
timestamp 1728304996
transform -1 0 3810 0 -1 250
box -12 -8 92 252
use NAND3X1  _1630_
timestamp 1728305047
transform 1 0 3610 0 -1 250
box -12 -8 112 252
use NAND2X1  _1631_
timestamp 1728304996
transform 1 0 3830 0 -1 250
box -12 -8 92 252
use NAND2X1  _1632_
timestamp 1728304996
transform -1 0 2350 0 -1 250
box -12 -8 92 252
use NOR2X1  _1633_
timestamp 1728305106
transform -1 0 2970 0 -1 250
box -12 -8 92 252
use NAND2X1  _1634_
timestamp 1728304996
transform -1 0 2870 0 -1 250
box -12 -8 92 252
use OAI21X1  _1635_
timestamp 1728305162
transform 1 0 2670 0 -1 250
box -12 -8 112 252
use NAND2X1  _1636_
timestamp 1728304996
transform 1 0 4730 0 -1 250
box -12 -8 92 252
use NOR2X1  _1637_
timestamp 1728305106
transform 1 0 4630 0 -1 250
box -12 -8 92 252
use AOI21X1  _1638_
timestamp 1728304211
transform 1 0 4410 0 -1 250
box -12 -8 112 252
use NOR2X1  _1639_
timestamp 1728305106
transform 1 0 4530 0 -1 250
box -12 -8 92 252
use NOR2X1  _1640_
timestamp 1728305106
transform 1 0 2210 0 1 250
box -12 -8 92 252
use NOR2X1  _1641_
timestamp 1728305106
transform 1 0 2310 0 1 250
box -12 -8 92 252
use INVX1  _1642_
timestamp 1749781103
transform 1 0 3230 0 -1 250
box -12 -8 72 252
use OAI21X1  _1643_
timestamp 1728305162
transform 1 0 3310 0 -1 250
box -12 -8 112 252
use OAI21X1  _1644_
timestamp 1728305162
transform -1 0 2870 0 1 250
box -12 -8 112 252
use OAI21X1  _1645_
timestamp 1728305162
transform 1 0 2650 0 1 250
box -12 -8 112 252
use AOI22X1  _1646_
timestamp 1728304278
transform -1 0 3110 0 -1 250
box -14 -8 132 252
use NAND2X1  _1647_
timestamp 1728304996
transform 1 0 3130 0 -1 250
box -12 -8 92 252
use OAI21X1  _1648_
timestamp 1728305162
transform -1 0 3230 0 1 250
box -12 -8 112 252
use OR2X2  _1649_
timestamp 1728305284
transform -1 0 2630 0 1 250
box -12 -8 112 252
use AOI21X1  _1650_
timestamp 1728304211
transform -1 0 2530 0 1 250
box -12 -8 112 252
use AOI21X1  _1651_
timestamp 1728304211
transform 1 0 2330 0 -1 730
box -12 -8 112 252
use INVX1  _1652_
timestamp 1749781103
transform -1 0 4330 0 1 3130
box -12 -8 72 252
use OAI21X1  _1653_
timestamp 1728305162
transform 1 0 4470 0 -1 1690
box -12 -8 112 252
use NOR2X1  _1654_
timestamp 1728305106
transform -1 0 4530 0 -1 2170
box -12 -8 92 252
use INVX1  _1655_
timestamp 1749781103
transform 1 0 4670 0 1 1690
box -12 -8 72 252
use NAND3X1  _1656_
timestamp 1728305047
transform 1 0 4770 0 1 1690
box -12 -8 112 252
use NAND2X1  _1657_
timestamp 1728304996
transform -1 0 4610 0 -1 2170
box -12 -8 92 252
use NOR2X1  _1658_
timestamp 1728305106
transform -1 0 4390 0 1 5050
box -12 -8 92 252
use NOR2X1  _1659_
timestamp 1728305106
transform -1 0 4050 0 -1 5050
box -12 -8 92 252
use NAND2X1  _1660_
timestamp 1728304996
transform -1 0 4190 0 1 5050
box -12 -8 92 252
use NOR2X1  _1661_
timestamp 1728305106
transform -1 0 3610 0 -1 4090
box -12 -8 92 252
use INVX1  _1662_
timestamp 1749781103
transform 1 0 3650 0 -1 4090
box -12 -8 72 252
use NAND2X1  _1663_
timestamp 1728304996
transform 1 0 3010 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1664_
timestamp 1728305162
transform 1 0 3430 0 1 3610
box -12 -8 112 252
use NOR2X1  _1665_
timestamp 1728305106
transform -1 0 3610 0 1 3610
box -12 -8 92 252
use OAI21X1  _1666_
timestamp 1728305162
transform -1 0 4130 0 1 1210
box -12 -8 112 252
use OAI21X1  _1667_
timestamp 1728305162
transform 1 0 4150 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1668_
timestamp 1728305047
transform 1 0 3930 0 1 730
box -12 -8 112 252
use NAND2X1  _1669_
timestamp 1728304996
transform -1 0 4110 0 1 730
box -12 -8 92 252
use NAND3X1  _1670_
timestamp 1728305047
transform -1 0 4850 0 1 250
box -12 -8 112 252
use NAND2X1  _1671_
timestamp 1728304996
transform -1 0 4970 0 -1 730
box -12 -8 92 252
use NAND2X1  _1672_
timestamp 1728304996
transform -1 0 4710 0 1 250
box -12 -8 92 252
use NOR2X1  _1673_
timestamp 1728305106
transform 1 0 4610 0 -1 730
box -12 -8 92 252
use OAI21X1  _1674_
timestamp 1728305162
transform -1 0 4150 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1675_
timestamp 1728305162
transform -1 0 3330 0 1 730
box -12 -8 112 252
use NAND3X1  _1676_
timestamp 1728305047
transform 1 0 3490 0 -1 730
box -12 -8 112 252
use NAND3X1  _1677_
timestamp 1728305047
transform 1 0 3650 0 1 730
box -12 -8 112 252
use NAND3X1  _1678_
timestamp 1728305047
transform 1 0 3830 0 -1 730
box -12 -8 112 252
use AOI21X1  _1679_
timestamp 1728304211
transform -1 0 4030 0 -1 730
box -12 -8 112 252
use AOI22X1  _1680_
timestamp 1728304278
transform 1 0 1330 0 -1 2170
box -14 -8 132 252
use INVX1  _1681_
timestamp 1749781103
transform 1 0 1810 0 -1 1690
box -12 -8 72 252
use NAND2X1  _1682_
timestamp 1728304996
transform 1 0 1590 0 -1 1690
box -12 -8 92 252
use INVX1  _1683_
timestamp 1749781103
transform -1 0 1590 0 1 1210
box -12 -8 72 252
use NAND2X1  _1684_
timestamp 1728304996
transform 1 0 1610 0 1 1690
box -12 -8 92 252
use NAND3X1  _1685_
timestamp 1728305047
transform 1 0 1610 0 1 1210
box -12 -8 112 252
use NAND2X1  _1686_
timestamp 1728304996
transform 1 0 1810 0 1 1690
box -12 -8 92 252
use NAND2X1  _1687_
timestamp 1728304996
transform -1 0 1790 0 1 1690
box -12 -8 92 252
use NAND2X1  _1688_
timestamp 1728304996
transform 1 0 1490 0 -1 1690
box -12 -8 92 252
use NOR2X1  _1689_
timestamp 1728305106
transform 1 0 970 0 -1 1690
box -12 -8 92 252
use INVX1  _1690_
timestamp 1749781103
transform 1 0 1170 0 -1 1690
box -12 -8 72 252
use NAND3X1  _1691_
timestamp 1728305047
transform 1 0 730 0 1 1210
box -12 -8 112 252
use INVX1  _1692_
timestamp 1749781103
transform 1 0 1310 0 1 1210
box -12 -8 72 252
use OAI21X1  _1693_
timestamp 1728305162
transform 1 0 1250 0 -1 1690
box -12 -8 112 252
use OAI22X1  _1694_
timestamp 1728305200
transform -1 0 1510 0 1 1210
box -12 -8 132 252
use NAND3X1  _1695_
timestamp 1728305047
transform 1 0 4610 0 -1 1210
box -12 -8 112 252
use AND2X2  _1696_
timestamp 1728304163
transform 1 0 4130 0 1 730
box -12 -8 112 252
use NAND3X1  _1697_
timestamp 1728305047
transform 1 0 5010 0 -1 250
box -12 -8 112 252
use NAND2X1  _1698_
timestamp 1728304996
transform 1 0 4830 0 -1 250
box -12 -8 92 252
use NAND2X1  _1699_
timestamp 1728304996
transform 1 0 5130 0 -1 250
box -12 -8 92 252
use AOI21X1  _1700_
timestamp 1728304211
transform -1 0 3450 0 -1 730
box -12 -8 112 252
use NAND2X1  _1701_
timestamp 1728304996
transform 1 0 3450 0 1 730
box -12 -8 92 252
use OAI21X1  _1702_
timestamp 1728305162
transform -1 0 3650 0 1 730
box -12 -8 112 252
use NAND3X1  _1703_
timestamp 1728305047
transform 1 0 4370 0 1 730
box -12 -8 112 252
use AOI21X1  _1704_
timestamp 1728304211
transform 1 0 4270 0 -1 730
box -12 -8 112 252
use OAI21X1  _1705_
timestamp 1728305162
transform -1 0 4490 0 -1 730
box -12 -8 112 252
use AND2X2  _1706_
timestamp 1728304163
transform 1 0 4510 0 -1 730
box -12 -8 112 252
use NAND3X1  _1707_
timestamp 1728305047
transform 1 0 4730 0 -1 1210
box -12 -8 112 252
use NOR2X1  _1708_
timestamp 1728305106
transform 1 0 730 0 -1 1690
box -12 -8 92 252
use NOR2X1  _1709_
timestamp 1728305106
transform -1 0 1150 0 -1 1690
box -12 -8 92 252
use AND2X2  _1710_
timestamp 1728304163
transform 1 0 1370 0 -1 1690
box -12 -8 112 252
use OAI21X1  _1711_
timestamp 1728305162
transform -1 0 1790 0 -1 1690
box -12 -8 112 252
use NOR2X1  _1712_
timestamp 1728305106
transform -1 0 1810 0 1 1210
box -12 -8 92 252
use NAND3X1  _1713_
timestamp 1728305047
transform 1 0 4490 0 -1 1210
box -12 -8 112 252
use NAND2X1  _1714_
timestamp 1728304996
transform 1 0 4110 0 1 1690
box -12 -8 92 252
use NAND3X1  _1715_
timestamp 1728305047
transform 1 0 4570 0 1 1690
box -12 -8 112 252
use NAND3X1  _1716_
timestamp 1728305047
transform -1 0 2750 0 1 730
box -12 -8 112 252
use OAI21X1  _1717_
timestamp 1728305162
transform -1 0 2550 0 1 730
box -12 -8 112 252
use OAI21X1  _1718_
timestamp 1728305162
transform 1 0 2310 0 1 730
box -12 -8 112 252
use NAND3X1  _1719_
timestamp 1728305047
transform -1 0 710 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1720_
timestamp 1728305047
transform -1 0 390 0 1 1210
box -12 -8 112 252
use OAI21X1  _1721_
timestamp 1728305162
transform 1 0 130 0 -1 1690
box -12 -8 112 252
use NAND3X1  _1722_
timestamp 1728305047
transform -1 0 590 0 1 1690
box -12 -8 112 252
use NAND3X1  _1723_
timestamp 1728305047
transform 1 0 490 0 -1 1690
box -12 -8 112 252
use AND2X2  _1724_
timestamp 1728304163
transform 1 0 610 0 1 1210
box -12 -8 112 252
use NAND3X1  _1725_
timestamp 1728305047
transform -1 0 1370 0 1 730
box -12 -8 112 252
use NAND3X1  _1726_
timestamp 1728305047
transform 1 0 710 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1727_
timestamp 1728305162
transform 1 0 850 0 -1 1690
box -12 -8 112 252
use OAI21X1  _1728_
timestamp 1728305162
transform -1 0 1290 0 1 1210
box -12 -8 112 252
use INVX1  _1729_
timestamp 1749781103
transform -1 0 210 0 -1 1210
box -12 -8 72 252
use AOI21X1  _1730_
timestamp 1728304211
transform -1 0 570 0 -1 1210
box -12 -8 112 252
use AOI21X1  _1731_
timestamp 1728304211
transform 1 0 250 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1732_
timestamp 1728305162
transform 1 0 1350 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1733_
timestamp 1728305047
transform 1 0 2850 0 -1 730
box -12 -8 112 252
use OAI21X1  _1734_
timestamp 1728305162
transform 1 0 2710 0 -1 730
box -12 -8 112 252
use OAI21X1  _1735_
timestamp 1728305162
transform 1 0 2090 0 1 250
box -12 -8 112 252
use NAND3X1  _1736_
timestamp 1728305047
transform -1 0 1970 0 1 250
box -12 -8 112 252
use AOI22X1  _1737_
timestamp 1728304278
transform 1 0 2590 0 -1 730
box -14 -8 132 252
use AOI22X1  _1738_
timestamp 1728304278
transform -1 0 2590 0 -1 1210
box -14 -8 132 252
use NAND2X1  _1739_
timestamp 1728304996
transform -1 0 2550 0 -1 730
box -12 -8 92 252
use NAND3X1  _1740_
timestamp 1728305047
transform 1 0 2550 0 1 730
box -12 -8 112 252
use NAND2X1  _1741_
timestamp 1728304996
transform -1 0 610 0 1 1210
box -12 -8 92 252
use NAND3X1  _1742_
timestamp 1728305047
transform 1 0 910 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1743_
timestamp 1728305047
transform -1 0 1130 0 1 730
box -12 -8 112 252
use AOI21X1  _1744_
timestamp 1728304211
transform 1 0 1010 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1745_
timestamp 1728305047
transform 1 0 1090 0 1 1210
box -12 -8 112 252
use INVX1  _1746_
timestamp 1749781103
transform 1 0 1550 0 -1 1210
box -12 -8 72 252
use NAND2X1  _1747_
timestamp 1728304996
transform -1 0 1710 0 -1 1210
box -12 -8 92 252
use OAI22X1  _1748_
timestamp 1728305200
transform -1 0 2990 0 -1 1210
box -12 -8 132 252
use AOI22X1  _1749_
timestamp 1728304278
transform -1 0 3130 0 1 1210
box -14 -8 132 252
use OAI21X1  _1750_
timestamp 1728305162
transform 1 0 3010 0 -1 1210
box -12 -8 112 252
use AOI22X1  _1751_
timestamp 1728304278
transform -1 0 3770 0 1 1690
box -14 -8 132 252
use OR2X2  _1752_
timestamp 1728305284
transform -1 0 3830 0 -1 2170
box -12 -8 112 252
use NAND2X1  _1753_
timestamp 1728304996
transform 1 0 3370 0 1 4090
box -12 -8 92 252
use AOI21X1  _1754_
timestamp 1728304211
transform -1 0 3030 0 1 4090
box -12 -8 112 252
use NAND2X1  _1755_
timestamp 1728304996
transform -1 0 2910 0 1 4090
box -12 -8 92 252
use NOR3X1  _1756_
timestamp 1728303224
transform 1 0 3050 0 1 4090
box -12 -8 192 252
use AOI21X1  _1757_
timestamp 1728304211
transform 1 0 3510 0 -1 1690
box -12 -8 112 252
use INVX1  _1758_
timestamp 1749781103
transform 1 0 3430 0 -1 2170
box -12 -8 72 252
use NAND3X1  _1759_
timestamp 1728305047
transform -1 0 3410 0 -1 2170
box -12 -8 112 252
use AOI21X1  _1760_
timestamp 1728304211
transform 1 0 3790 0 1 1690
box -12 -8 112 252
use AOI21X1  _1761_
timestamp 1728304211
transform -1 0 4290 0 -1 2170
box -12 -8 112 252
use OAI21X1  _1762_
timestamp 1728305162
transform -1 0 4210 0 1 2650
box -12 -8 112 252
use INVX1  _1763_
timestamp 1749781103
transform 1 0 4210 0 -1 3130
box -12 -8 72 252
use INVX1  _1764_
timestamp 1749781103
transform 1 0 4130 0 -1 2650
box -12 -8 72 252
use NAND2X1  _1765_
timestamp 1728304996
transform 1 0 4050 0 -1 730
box -12 -8 92 252
use AND2X2  _1766_
timestamp 1728304163
transform 1 0 3690 0 -1 730
box -12 -8 112 252
use NAND3X1  _1767_
timestamp 1728305047
transform 1 0 4150 0 -1 730
box -12 -8 112 252
use NOR3X1  _1768_
timestamp 1728303224
transform 1 0 4710 0 -1 730
box -12 -8 192 252
use NAND2X1  _1769_
timestamp 1728304996
transform 1 0 4610 0 1 730
box -12 -8 92 252
use AOI21X1  _1770_
timestamp 1728304211
transform -1 0 4590 0 1 730
box -12 -8 112 252
use NAND3X1  _1771_
timestamp 1728305047
transform -1 0 4350 0 1 730
box -12 -8 112 252
use INVX1  _1772_
timestamp 1749781103
transform -1 0 3990 0 1 1210
box -12 -8 72 252
use OAI21X1  _1773_
timestamp 1728305162
transform 1 0 4250 0 1 1210
box -12 -8 112 252
use OAI21X1  _1774_
timestamp 1728305162
transform -1 0 4370 0 -1 1690
box -12 -8 112 252
use AOI21X1  _1775_
timestamp 1728304211
transform -1 0 4310 0 -1 2650
box -12 -8 112 252
use INVX1  _1776_
timestamp 1749781103
transform -1 0 4490 0 -1 2650
box -12 -8 72 252
use AND2X2  _1777_
timestamp 1728304163
transform -1 0 4530 0 1 1690
box -12 -8 112 252
use NAND2X1  _1778_
timestamp 1728304996
transform -1 0 2710 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1779_
timestamp 1728304996
transform -1 0 910 0 1 1210
box -12 -8 92 252
use OAI21X1  _1780_
timestamp 1728305162
transform -1 0 1050 0 1 1210
box -12 -8 112 252
use AOI21X1  _1781_
timestamp 1728304211
transform -1 0 1230 0 1 730
box -12 -8 112 252
use OAI21X1  _1782_
timestamp 1728305162
transform 1 0 1150 0 -1 1210
box -12 -8 112 252
use AOI21X1  _1783_
timestamp 1728304211
transform 1 0 1250 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1784_
timestamp 1728305162
transform -1 0 2850 0 -1 1210
box -12 -8 112 252
use NOR2X1  _1785_
timestamp 1728305106
transform -1 0 1530 0 -1 1210
box -12 -8 92 252
use AOI22X1  _1786_
timestamp 1728304278
transform -1 0 2610 0 1 1210
box -14 -8 132 252
use OAI22X1  _1787_
timestamp 1728305200
transform 1 0 3070 0 -1 1690
box -12 -8 132 252
use AOI21X1  _1788_
timestamp 1728304211
transform 1 0 2970 0 -1 1690
box -12 -8 112 252
use INVX1  _1789_
timestamp 1749781103
transform -1 0 3950 0 1 1690
box -12 -8 72 252
use NOR2X1  _1790_
timestamp 1728305106
transform -1 0 3530 0 1 2170
box -12 -8 92 252
use INVX1  _1791_
timestamp 1749781103
transform -1 0 3250 0 -1 4090
box -12 -8 72 252
use INVX1  _1792_
timestamp 1749781103
transform 1 0 3130 0 -1 4090
box -12 -8 72 252
use NAND3X1  _1793_
timestamp 1728305047
transform 1 0 3250 0 -1 4090
box -12 -8 112 252
use NOR3X1  _1794_
timestamp 1728303224
transform 1 0 3530 0 -1 2170
box -12 -8 192 252
use OAI21X1  _1795_
timestamp 1728305162
transform 1 0 3950 0 1 1690
box -12 -8 112 252
use AOI21X1  _1796_
timestamp 1728304211
transform -1 0 4410 0 1 1690
box -12 -8 112 252
use NAND3X1  _1797_
timestamp 1728305047
transform -1 0 4410 0 -1 2650
box -12 -8 112 252
use OAI21X1  _1798_
timestamp 1728305162
transform 1 0 4310 0 -1 3130
box -12 -8 112 252
use INVX2  _1799_
timestamp 1749781103
transform 1 0 4270 0 -1 5530
box -12 -8 72 252
use OAI21X1  _1800_
timestamp 1728305162
transform 1 0 4450 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1801_
timestamp 1728305162
transform 1 0 4250 0 1 3610
box -12 -8 112 252
use NAND2X1  _1802_
timestamp 1728304996
transform 1 0 3830 0 -1 5050
box -12 -8 92 252
use NAND2X1  _1803_
timestamp 1728304996
transform 1 0 3590 0 -1 5050
box -12 -8 92 252
use NAND2X1  _1804_
timestamp 1728304996
transform -1 0 3790 0 -1 5050
box -12 -8 92 252
use NAND2X1  _1805_
timestamp 1728304996
transform -1 0 4370 0 1 4570
box -12 -8 92 252
use INVX1  _1806_
timestamp 1749781103
transform 1 0 4730 0 -1 5050
box -12 -8 72 252
use NOR2X1  _1807_
timestamp 1728305106
transform 1 0 5070 0 -1 5050
box -12 -8 92 252
use OR2X2  _1808_
timestamp 1728305284
transform -1 0 4930 0 -1 5050
box -12 -8 112 252
use NOR2X1  _1809_
timestamp 1728305106
transform 1 0 4530 0 1 5050
box -12 -8 92 252
use OAI21X1  _1810_
timestamp 1728305162
transform 1 0 4090 0 1 4570
box -12 -8 112 252
use NAND2X1  _1811_
timestamp 1728304996
transform -1 0 3970 0 -1 3610
box -12 -8 92 252
use NAND2X1  _1812_
timestamp 1728304996
transform -1 0 4550 0 -1 3610
box -12 -8 92 252
use NOR2X1  _1813_
timestamp 1728305106
transform 1 0 4090 0 -1 3610
box -12 -8 92 252
use OAI21X1  _1814_
timestamp 1728305162
transform -1 0 4030 0 1 3610
box -12 -8 112 252
use NOR2X1  _1815_
timestamp 1728305106
transform 1 0 3470 0 1 4090
box -12 -8 92 252
use NOR2X1  _1816_
timestamp 1728305106
transform 1 0 3730 0 1 4090
box -12 -8 92 252
use NOR2X1  _1817_
timestamp 1728305106
transform -1 0 3810 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1818_
timestamp 1728305106
transform 1 0 3790 0 -1 4570
box -12 -8 92 252
use NOR2X1  _1819_
timestamp 1728305106
transform 1 0 3990 0 -1 4570
box -12 -8 92 252
use NOR2X1  _1820_
timestamp 1728305106
transform -1 0 3970 0 -1 4570
box -12 -8 92 252
use NAND3X1  _1821_
timestamp 1728305047
transform 1 0 4050 0 1 4090
box -12 -8 112 252
use NAND2X1  _1822_
timestamp 1728304996
transform 1 0 4210 0 1 4570
box -12 -8 92 252
use NAND2X1  _1823_
timestamp 1728304996
transform 1 0 4670 0 -1 5530
box -12 -8 92 252
use NAND2X1  _1824_
timestamp 1728304996
transform -1 0 4430 0 -1 5530
box -12 -8 92 252
use NAND2X1  _1825_
timestamp 1728304996
transform -1 0 4650 0 -1 5530
box -12 -8 92 252
use INVX1  _1826_
timestamp 1749781103
transform -1 0 5050 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1827_
timestamp 1728304996
transform 1 0 5570 0 -1 5530
box -12 -8 92 252
use INVX1  _1828_
timestamp 1749781103
transform -1 0 5550 0 -1 5530
box -12 -8 72 252
use NOR2X1  _1829_
timestamp 1728305106
transform 1 0 5550 0 1 5050
box -12 -8 92 252
use NOR2X1  _1830_
timestamp 1728305106
transform -1 0 5530 0 1 5050
box -12 -8 92 252
use AND2X2  _1831_
timestamp 1728304163
transform -1 0 4970 0 -1 5530
box -12 -8 112 252
use NAND3X1  _1832_
timestamp 1728305047
transform -1 0 4550 0 -1 5530
box -12 -8 112 252
use INVX1  _1833_
timestamp 1749781103
transform 1 0 4210 0 1 5050
box -12 -8 72 252
use NAND3X1  _1834_
timestamp 1728305047
transform -1 0 4270 0 -1 5530
box -12 -8 112 252
use OAI21X1  _1835_
timestamp 1728305162
transform -1 0 4150 0 -1 5530
box -12 -8 112 252
use OR2X2  _1836_
timestamp 1728305284
transform 1 0 3850 0 1 4570
box -12 -8 112 252
use NAND2X1  _1837_
timestamp 1728304996
transform 1 0 3750 0 1 4570
box -12 -8 92 252
use NAND2X1  _1838_
timestamp 1728304996
transform 1 0 3970 0 1 4570
box -12 -8 92 252
use INVX1  _1839_
timestamp 1749781103
transform 1 0 4290 0 -1 5050
box -12 -8 72 252
use INVX1  _1840_
timestamp 1749781103
transform -1 0 4770 0 1 5050
box -12 -8 72 252
use NAND2X1  _1841_
timestamp 1728304996
transform 1 0 4770 0 -1 5530
box -12 -8 92 252
use OAI21X1  _1842_
timestamp 1728305162
transform 1 0 4430 0 1 5050
box -12 -8 112 252
use NAND2X1  _1843_
timestamp 1728304996
transform 1 0 4610 0 1 5050
box -12 -8 92 252
use NAND3X1  _1844_
timestamp 1728305047
transform 1 0 4390 0 -1 5050
box -12 -8 112 252
use OAI21X1  _1845_
timestamp 1728305162
transform 1 0 4050 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1846_
timestamp 1728304996
transform -1 0 4270 0 -1 5050
box -12 -8 92 252
use AND2X2  _1847_
timestamp 1728304163
transform 1 0 4590 0 -1 5050
box -12 -8 112 252
use OAI21X1  _1848_
timestamp 1728305162
transform 1 0 4970 0 -1 5050
box -12 -8 112 252
use OAI21X1  _1849_
timestamp 1728305162
transform -1 0 5090 0 1 5050
box -12 -8 112 252
use NAND3X1  _1850_
timestamp 1728305047
transform 1 0 4810 0 1 5050
box -12 -8 112 252
use NAND2X1  _1851_
timestamp 1728304996
transform 1 0 4910 0 1 5050
box -12 -8 92 252
use NAND2X1  _1852_
timestamp 1728304996
transform -1 0 5170 0 -1 5530
box -12 -8 92 252
use NAND3X1  _1853_
timestamp 1728305047
transform 1 0 5170 0 -1 5530
box -12 -8 112 252
use INVX1  _1854_
timestamp 1749781103
transform 1 0 5410 0 -1 5530
box -12 -8 72 252
use OAI21X1  _1855_
timestamp 1728305162
transform -1 0 5370 0 -1 5530
box -12 -8 112 252
use NAND2X1  _1856_
timestamp 1728304996
transform 1 0 5250 0 1 5050
box -12 -8 92 252
use INVX1  _1857_
timestamp 1749781103
transform -1 0 3610 0 1 4090
box -12 -8 72 252
use INVX1  _1858_
timestamp 1749781103
transform -1 0 4010 0 -1 4090
box -12 -8 72 252
use OAI21X1  _1859_
timestamp 1728305162
transform -1 0 3710 0 1 4090
box -12 -8 112 252
use OR2X2  _1860_
timestamp 1728305284
transform 1 0 3930 0 1 4090
box -12 -8 112 252
use NAND2X1  _1861_
timestamp 1728304996
transform -1 0 3890 0 1 4090
box -12 -8 92 252
use INVX1  _1862_
timestamp 1749781103
transform -1 0 3910 0 1 3610
box -12 -8 72 252
use NOR2X1  _1863_
timestamp 1728305106
transform 1 0 4370 0 -1 3610
box -12 -8 92 252
use OR2X2  _1864_
timestamp 1728305284
transform 1 0 4070 0 1 3610
box -12 -8 112 252
use INVX1  _1865_
timestamp 1749781103
transform -1 0 3670 0 1 3610
box -12 -8 72 252
use NAND3X1  _1866_
timestamp 1728305047
transform 1 0 3710 0 1 3610
box -12 -8 112 252
use INVX1  _1867_
timestamp 1749781103
transform 1 0 4170 0 -1 3610
box -12 -8 72 252
use OAI21X1  _1868_
timestamp 1728305162
transform 1 0 4270 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1869_
timestamp 1728304996
transform -1 0 4250 0 1 3610
box -12 -8 92 252
use NAND2X1  _1870_
timestamp 1728304996
transform 1 0 4050 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1871_
timestamp 1728305162
transform 1 0 3810 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1872_
timestamp 1728304996
transform 1 0 4170 0 -1 4090
box -12 -8 92 252
use NAND3X1  _1873_
timestamp 1728305047
transform 1 0 4250 0 -1 4090
box -12 -8 112 252
use AOI21X1  _1874_
timestamp 1728304211
transform 1 0 4310 0 1 4090
box -12 -8 112 252
use OR2X2  _1875_
timestamp 1728305284
transform 1 0 5110 0 1 5050
box -12 -8 112 252
use NAND2X1  _1876_
timestamp 1728304996
transform 1 0 5350 0 1 5050
box -12 -8 92 252
use NAND2X1  _1877_
timestamp 1728304996
transform 1 0 4810 0 -1 4570
box -12 -8 92 252
use NOR3X1  _1878_
timestamp 1728303224
transform -1 0 4910 0 1 4570
box -12 -8 192 252
use OAI21X1  _1879_
timestamp 1728305162
transform -1 0 4710 0 1 4570
box -12 -8 112 252
use OR2X2  _1880_
timestamp 1728305284
transform -1 0 4590 0 1 3610
box -12 -8 112 252
use OAI21X1  _1881_
timestamp 1728305162
transform -1 0 4470 0 1 3610
box -12 -8 112 252
use NAND2X1  _1882_
timestamp 1728304996
transform -1 0 4590 0 1 4570
box -12 -8 92 252
use OR2X2  _1883_
timestamp 1728305284
transform 1 0 4370 0 -1 4090
box -12 -8 112 252
use OAI22X1  _1884_
timestamp 1728305200
transform 1 0 4490 0 -1 4090
box -12 -8 132 252
use OAI21X1  _1885_
timestamp 1728305162
transform 1 0 5570 0 -1 4090
box -12 -8 112 252
use OR2X2  _1886_
timestamp 1728305284
transform 1 0 5230 0 -1 4090
box -12 -8 112 252
use OAI21X1  _1887_
timestamp 1728305162
transform 1 0 5450 0 -1 4090
box -12 -8 112 252
use OAI21X1  _1888_
timestamp 1728305162
transform -1 0 4650 0 1 4090
box -12 -8 112 252
use NAND3X1  _1889_
timestamp 1728305047
transform -1 0 4270 0 1 4090
box -12 -8 112 252
use OAI21X1  _1890_
timestamp 1728305162
transform 1 0 4430 0 1 4090
box -12 -8 112 252
use OAI21X1  _1891_
timestamp 1728305162
transform 1 0 5550 0 -1 4570
box -12 -8 112 252
use OR2X2  _1892_
timestamp 1728305284
transform 1 0 5310 0 -1 4570
box -12 -8 112 252
use OAI21X1  _1893_
timestamp 1728305162
transform 1 0 5430 0 -1 4570
box -12 -8 112 252
use OAI21X1  _1894_
timestamp 1728305162
transform -1 0 5210 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1895_
timestamp 1728304996
transform -1 0 5010 0 1 4570
box -12 -8 92 252
use OAI21X1  _1896_
timestamp 1728305162
transform 1 0 5030 0 1 4570
box -12 -8 112 252
use OAI21X1  _1897_
timestamp 1728305162
transform -1 0 5170 0 1 3610
box -12 -8 112 252
use NAND2X1  _1898_
timestamp 1728304996
transform -1 0 4930 0 1 3610
box -12 -8 92 252
use OAI21X1  _1899_
timestamp 1728305162
transform 1 0 4950 0 1 3610
box -12 -8 112 252
use NAND2X1  _1900_
timestamp 1728304996
transform 1 0 4510 0 -1 5050
box -12 -8 92 252
use NAND3X1  _1901_
timestamp 1728305047
transform -1 0 4490 0 1 4570
box -12 -8 112 252
use OAI21X1  _1902_
timestamp 1728305162
transform -1 0 4190 0 -1 4570
box -12 -8 112 252
use OAI21X1  _1903_
timestamp 1728305162
transform -1 0 4310 0 -1 4570
box -12 -8 112 252
use NOR2X1  _1904_
timestamp 1728305106
transform 1 0 3990 0 -1 3610
box -12 -8 92 252
use NAND2X1  _1905_
timestamp 1728304996
transform -1 0 5110 0 -1 3130
box -12 -8 92 252
use OAI21X1  _1906_
timestamp 1728305162
transform -1 0 4690 0 -1 2650
box -12 -8 112 252
use OAI21X1  _1907_
timestamp 1728305162
transform -1 0 4750 0 -1 2170
box -12 -8 112 252
use DFFSR  _1908_
timestamp 1728387359
transform -1 0 5730 0 -1 3610
box -12 -8 492 252
use DFFSR  _1909_
timestamp 1728387359
transform -1 0 4690 0 1 2650
box -12 -8 492 252
use DFFSR  _1910_
timestamp 1728387359
transform 1 0 4690 0 -1 2650
box -12 -8 492 252
use DFFSR  _1911_
timestamp 1728387359
transform 1 0 5210 0 1 1690
box -12 -8 492 252
use DFFSR  _1912_
timestamp 1728387359
transform -1 0 5690 0 -1 250
box -12 -8 492 252
use DFFSR  _1913_
timestamp 1728387359
transform -1 0 5650 0 1 250
box -12 -8 492 252
use DFFSR  _1914_
timestamp 1728387359
transform -1 0 5650 0 -1 1210
box -12 -8 492 252
use DFFSR  _1915_
timestamp 1728387359
transform -1 0 4510 0 1 2170
box -12 -8 492 252
use DFFSR  _1916_
timestamp 1728387359
transform -1 0 4110 0 -1 2650
box -12 -8 492 252
use DFFSR  _1917_
timestamp 1728387359
transform 1 0 10 0 1 730
box -12 -8 492 252
use DFFSR  _1918_
timestamp 1728387359
transform 1 0 10 0 1 1690
box -12 -8 492 252
use DFFSR  _1919_
timestamp 1728387359
transform 1 0 10 0 -1 250
box -12 -8 492 252
use DFFSR  _1920_
timestamp 1728387359
transform 1 0 10 0 1 250
box -12 -8 492 252
use DFFSR  _1921_
timestamp 1728387359
transform 1 0 1210 0 -1 250
box -12 -8 492 252
use DFFSR  _1922_
timestamp 1728387359
transform -1 0 4390 0 -1 250
box -12 -8 492 252
use DFFSR  _1923_
timestamp 1728387359
transform -1 0 4590 0 1 250
box -12 -8 492 252
use DFFSR  _1924_
timestamp 1728387359
transform -1 0 4110 0 1 250
box -12 -8 492 252
use DFFSR  _1925_
timestamp 1728387359
transform 1 0 2070 0 -1 1690
box -12 -8 492 252
use DFFSR  _1926_
timestamp 1728387359
transform -1 0 4810 0 1 3130
box -12 -8 492 252
use DFFSR  _1927_
timestamp 1728387359
transform -1 0 4190 0 -1 3130
box -12 -8 492 252
use DFFSR  _1928_
timestamp 1728387359
transform -1 0 5670 0 1 3130
box -12 -8 492 252
use DFFSR  _1929_
timestamp 1728387359
transform -1 0 5030 0 -1 3610
box -12 -8 492 252
use DFFSR  _1930_
timestamp 1728387359
transform -1 0 5090 0 -1 4090
box -12 -8 492 252
use DFFSR  _1931_
timestamp 1728387359
transform -1 0 5610 0 1 4090
box -12 -8 492 252
use DFFSR  _1932_
timestamp 1728387359
transform -1 0 5130 0 1 4090
box -12 -8 492 252
use DFFSR  _1933_
timestamp 1728387359
transform -1 0 5610 0 1 4570
box -12 -8 492 252
use DFFSR  _1934_
timestamp 1728387359
transform -1 0 5630 0 -1 5050
box -12 -8 492 252
use DFFSR  _1935_
timestamp 1728387359
transform -1 0 5650 0 1 3610
box -12 -8 492 252
use DFFSR  _1936_
timestamp 1728387359
transform -1 0 4790 0 -1 4570
box -12 -8 492 252
use DFFSR  _1937_
timestamp 1728387359
transform -1 0 4230 0 1 3130
box -12 -8 492 252
use DFFSR  _1938_
timestamp 1728387359
transform -1 0 5650 0 -1 3130
box -12 -8 492 252
use DFFSR  _1939_
timestamp 1728387359
transform -1 0 5670 0 1 2650
box -12 -8 492 252
use DFFSR  _1940_
timestamp 1728387359
transform 1 0 4510 0 1 2170
box -12 -8 492 252
use BUFX2  _1941_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304320
transform 1 0 3610 0 1 2170
box -12 -8 92 252
use BUFX2  _1942_
timestamp 1728304320
transform 1 0 3810 0 1 2650
box -12 -8 92 252
use BUFX2  _1943_
timestamp 1728304320
transform 1 0 3530 0 1 2170
box -12 -8 92 252
use BUFX2  _1944_
timestamp 1728304320
transform 1 0 3410 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert0
timestamp 1728304320
transform -1 0 750 0 -1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert1
timestamp 1728304320
transform 1 0 1470 0 1 3610
box -12 -8 92 252
use BUFX2  BUFX2_insert2
timestamp 1728304320
transform -1 0 1430 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert3
timestamp 1728304320
transform 1 0 2310 0 -1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert11
timestamp 1728304320
transform 1 0 5130 0 -1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert12
timestamp 1728304320
transform 1 0 4890 0 1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert13
timestamp 1728304320
transform 1 0 4790 0 -1 2170
box -12 -8 92 252
use BUFX2  BUFX2_insert14
timestamp 1728304320
transform -1 0 4570 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert15
timestamp 1728304320
transform -1 0 1850 0 1 2170
box -12 -8 92 252
use CLKBUF1  CLKBUF1_insert4 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304421
transform 1 0 3430 0 1 250
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert5
timestamp 1728304421
transform -1 0 4830 0 1 3610
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert6
timestamp 1728304421
transform -1 0 1090 0 1 3610
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert7
timestamp 1728304421
transform -1 0 2790 0 -1 5530
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert8
timestamp 1728304421
transform -1 0 4090 0 1 2650
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert9
timestamp 1728304421
transform 1 0 4890 0 1 250
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert10
timestamp 1728304421
transform 1 0 4890 0 -1 4570
box -12 -8 212 252
use FILL  FILL84750x3750 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728341909
transform 1 0 5650 0 1 250
box -12 -8 32 252
use FILL  FILL84750x43350
timestamp 1728341909
transform -1 0 5670 0 -1 3130
box -12 -8 32 252
use FILL  FILL84750x54150
timestamp 1728341909
transform 1 0 5650 0 1 3610
box -12 -8 32 252
use FILL  FILL84750x64950
timestamp 1728341909
transform -1 0 5670 0 -1 4570
box -12 -8 32 252
use FILL  FILL84750x79350
timestamp 1728341909
transform -1 0 5670 0 -1 5530
box -12 -8 32 252
use FILL  FILL85050x3750
timestamp 1728341909
transform 1 0 5670 0 1 250
box -12 -8 32 252
use FILL  FILL85050x10950
timestamp 1728341909
transform 1 0 5670 0 1 730
box -12 -8 32 252
use FILL  FILL85050x32550
timestamp 1728341909
transform 1 0 5670 0 1 2170
box -12 -8 32 252
use FILL  FILL85050x39750
timestamp 1728341909
transform 1 0 5670 0 1 2650
box -12 -8 32 252
use FILL  FILL85050x43350
timestamp 1728341909
transform -1 0 5690 0 -1 3130
box -12 -8 32 252
use FILL  FILL85050x46950
timestamp 1728341909
transform 1 0 5670 0 1 3130
box -12 -8 32 252
use FILL  FILL85050x54150
timestamp 1728341909
transform 1 0 5670 0 1 3610
box -12 -8 32 252
use FILL  FILL85050x57750
timestamp 1728341909
transform -1 0 5690 0 -1 4090
box -12 -8 32 252
use FILL  FILL85050x64950
timestamp 1728341909
transform -1 0 5690 0 -1 4570
box -12 -8 32 252
use FILL  FILL85050x79350
timestamp 1728341909
transform -1 0 5690 0 -1 5530
box -12 -8 32 252
use FILL  FILL85350x150
timestamp 1728341909
transform -1 0 5710 0 -1 250
box -12 -8 32 252
use FILL  FILL85350x3750
timestamp 1728341909
transform 1 0 5690 0 1 250
box -12 -8 32 252
use FILL  FILL85350x10950
timestamp 1728341909
transform 1 0 5690 0 1 730
box -12 -8 32 252
use FILL  FILL85350x21750
timestamp 1728341909
transform -1 0 5710 0 -1 1690
box -12 -8 32 252
use FILL  FILL85350x25350
timestamp 1728341909
transform 1 0 5690 0 1 1690
box -12 -8 32 252
use FILL  FILL85350x32550
timestamp 1728341909
transform 1 0 5690 0 1 2170
box -12 -8 32 252
use FILL  FILL85350x39750
timestamp 1728341909
transform 1 0 5690 0 1 2650
box -12 -8 32 252
use FILL  FILL85350x43350
timestamp 1728341909
transform -1 0 5710 0 -1 3130
box -12 -8 32 252
use FILL  FILL85350x46950
timestamp 1728341909
transform 1 0 5690 0 1 3130
box -12 -8 32 252
use FILL  FILL85350x54150
timestamp 1728341909
transform 1 0 5690 0 1 3610
box -12 -8 32 252
use FILL  FILL85350x57750
timestamp 1728341909
transform -1 0 5710 0 -1 4090
box -12 -8 32 252
use FILL  FILL85350x64950
timestamp 1728341909
transform -1 0 5710 0 -1 4570
box -12 -8 32 252
use FILL  FILL85350x68550
timestamp 1728341909
transform 1 0 5690 0 1 4570
box -12 -8 32 252
use FILL  FILL85350x79350
timestamp 1728341909
transform -1 0 5710 0 -1 5530
box -12 -8 32 252
use FILL  FILL85650x150
timestamp 1728341909
transform -1 0 5730 0 -1 250
box -12 -8 32 252
use FILL  FILL85650x3750
timestamp 1728341909
transform 1 0 5710 0 1 250
box -12 -8 32 252
use FILL  FILL85650x7350
timestamp 1728341909
transform -1 0 5730 0 -1 730
box -12 -8 32 252
use FILL  FILL85650x10950
timestamp 1728341909
transform 1 0 5710 0 1 730
box -12 -8 32 252
use FILL  FILL85650x18150
timestamp 1728341909
transform 1 0 5710 0 1 1210
box -12 -8 32 252
use FILL  FILL85650x21750
timestamp 1728341909
transform -1 0 5730 0 -1 1690
box -12 -8 32 252
use FILL  FILL85650x25350
timestamp 1728341909
transform 1 0 5710 0 1 1690
box -12 -8 32 252
use FILL  FILL85650x32550
timestamp 1728341909
transform 1 0 5710 0 1 2170
box -12 -8 32 252
use FILL  FILL85650x39750
timestamp 1728341909
transform 1 0 5710 0 1 2650
box -12 -8 32 252
use FILL  FILL85650x43350
timestamp 1728341909
transform -1 0 5730 0 -1 3130
box -12 -8 32 252
use FILL  FILL85650x46950
timestamp 1728341909
transform 1 0 5710 0 1 3130
box -12 -8 32 252
use FILL  FILL85650x54150
timestamp 1728341909
transform 1 0 5710 0 1 3610
box -12 -8 32 252
use FILL  FILL85650x57750
timestamp 1728341909
transform -1 0 5730 0 -1 4090
box -12 -8 32 252
use FILL  FILL85650x64950
timestamp 1728341909
transform -1 0 5730 0 -1 4570
box -12 -8 32 252
use FILL  FILL85650x68550
timestamp 1728341909
transform 1 0 5710 0 1 4570
box -12 -8 32 252
use FILL  FILL85650x75750
timestamp 1728341909
transform 1 0 5710 0 1 5050
box -12 -8 32 252
use FILL  FILL85650x79350
timestamp 1728341909
transform -1 0 5730 0 -1 5530
box -12 -8 32 252
use FILL  FILL85950x150
timestamp 1728341909
transform -1 0 5750 0 -1 250
box -12 -8 32 252
use FILL  FILL85950x3750
timestamp 1728341909
transform 1 0 5730 0 1 250
box -12 -8 32 252
use FILL  FILL85950x7350
timestamp 1728341909
transform -1 0 5750 0 -1 730
box -12 -8 32 252
use FILL  FILL85950x10950
timestamp 1728341909
transform 1 0 5730 0 1 730
box -12 -8 32 252
use FILL  FILL85950x18150
timestamp 1728341909
transform 1 0 5730 0 1 1210
box -12 -8 32 252
use FILL  FILL85950x21750
timestamp 1728341909
transform -1 0 5750 0 -1 1690
box -12 -8 32 252
use FILL  FILL85950x25350
timestamp 1728341909
transform 1 0 5730 0 1 1690
box -12 -8 32 252
use FILL  FILL85950x28950
timestamp 1728341909
transform -1 0 5750 0 -1 2170
box -12 -8 32 252
use FILL  FILL85950x32550
timestamp 1728341909
transform 1 0 5730 0 1 2170
box -12 -8 32 252
use FILL  FILL85950x36150
timestamp 1728341909
transform -1 0 5750 0 -1 2650
box -12 -8 32 252
use FILL  FILL85950x39750
timestamp 1728341909
transform 1 0 5730 0 1 2650
box -12 -8 32 252
use FILL  FILL85950x43350
timestamp 1728341909
transform -1 0 5750 0 -1 3130
box -12 -8 32 252
use FILL  FILL85950x46950
timestamp 1728341909
transform 1 0 5730 0 1 3130
box -12 -8 32 252
use FILL  FILL85950x50550
timestamp 1728341909
transform -1 0 5750 0 -1 3610
box -12 -8 32 252
use FILL  FILL85950x54150
timestamp 1728341909
transform 1 0 5730 0 1 3610
box -12 -8 32 252
use FILL  FILL85950x57750
timestamp 1728341909
transform -1 0 5750 0 -1 4090
box -12 -8 32 252
use FILL  FILL85950x61350
timestamp 1728341909
transform 1 0 5730 0 1 4090
box -12 -8 32 252
use FILL  FILL85950x64950
timestamp 1728341909
transform -1 0 5750 0 -1 4570
box -12 -8 32 252
use FILL  FILL85950x68550
timestamp 1728341909
transform 1 0 5730 0 1 4570
box -12 -8 32 252
use FILL  FILL85950x72150
timestamp 1728341909
transform -1 0 5750 0 -1 5050
box -12 -8 32 252
use FILL  FILL85950x75750
timestamp 1728341909
transform 1 0 5730 0 1 5050
box -12 -8 32 252
use FILL  FILL85950x79350
timestamp 1728341909
transform -1 0 5750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__945_
timestamp 1728341909
transform 1 0 1570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__947_
timestamp 1728341909
transform 1 0 1890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__949_
timestamp 1728341909
transform 1 0 3130 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__951_
timestamp 1728341909
transform 1 0 2550 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__953_
timestamp 1728341909
transform 1 0 3150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__955_
timestamp 1728341909
transform 1 0 2410 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__957_
timestamp 1728341909
transform -1 0 2310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__959_
timestamp 1728341909
transform 1 0 2030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__961_
timestamp 1728341909
transform 1 0 2410 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__963_
timestamp 1728341909
transform 1 0 3470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__965_
timestamp 1728341909
transform -1 0 1710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__967_
timestamp 1728341909
transform 1 0 3430 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__969_
timestamp 1728341909
transform -1 0 2410 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__971_
timestamp 1728341909
transform -1 0 1370 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__972_
timestamp 1728341909
transform 1 0 1250 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__973_
timestamp 1728341909
transform -1 0 1030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__974_
timestamp 1728341909
transform -1 0 1130 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__975_
timestamp 1728341909
transform 1 0 2110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__976_
timestamp 1728341909
transform -1 0 2150 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__977_
timestamp 1728341909
transform -1 0 1250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__978_
timestamp 1728341909
transform -1 0 1090 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__979_
timestamp 1728341909
transform 1 0 2870 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__980_
timestamp 1728341909
transform -1 0 2650 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__981_
timestamp 1728341909
transform -1 0 2770 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__982_
timestamp 1728341909
transform 1 0 2210 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__983_
timestamp 1728341909
transform 1 0 1970 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__984_
timestamp 1728341909
transform 1 0 2210 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__985_
timestamp 1728341909
transform -1 0 2110 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__986_
timestamp 1728341909
transform 1 0 1630 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__987_
timestamp 1728341909
transform -1 0 1530 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__988_
timestamp 1728341909
transform 1 0 1670 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__989_
timestamp 1728341909
transform 1 0 1910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__990_
timestamp 1728341909
transform -1 0 2110 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__991_
timestamp 1728341909
transform -1 0 1990 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__992_
timestamp 1728341909
transform -1 0 1810 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__993_
timestamp 1728341909
transform 1 0 2750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__994_
timestamp 1728341909
transform 1 0 1790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__995_
timestamp 1728341909
transform -1 0 2190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__996_
timestamp 1728341909
transform 1 0 2290 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__997_
timestamp 1728341909
transform 1 0 2510 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__998_
timestamp 1728341909
transform 1 0 2630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__999_
timestamp 1728341909
transform -1 0 1590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1000_
timestamp 1728341909
transform 1 0 2030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1002_
timestamp 1728341909
transform 1 0 2370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1004_
timestamp 1728341909
transform -1 0 1450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1006_
timestamp 1728341909
transform -1 0 2590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1008_
timestamp 1728341909
transform 1 0 3130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1010_
timestamp 1728341909
transform 1 0 3330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1012_
timestamp 1728341909
transform 1 0 3190 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1014_
timestamp 1728341909
transform 1 0 2790 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1016_
timestamp 1728341909
transform 1 0 2930 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1017_
timestamp 1728341909
transform 1 0 3070 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1018_
timestamp 1728341909
transform 1 0 590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1019_
timestamp 1728341909
transform 1 0 2030 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1020_
timestamp 1728341909
transform -1 0 1930 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1021_
timestamp 1728341909
transform -1 0 510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1022_
timestamp 1728341909
transform -1 0 610 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1023_
timestamp 1728341909
transform -1 0 510 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1024_
timestamp 1728341909
transform 1 0 910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1025_
timestamp 1728341909
transform -1 0 690 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1026_
timestamp 1728341909
transform -1 0 710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1027_
timestamp 1728341909
transform 1 0 790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1028_
timestamp 1728341909
transform -1 0 510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1029_
timestamp 1728341909
transform -1 0 590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1030_
timestamp 1728341909
transform -1 0 790 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1031_
timestamp 1728341909
transform -1 0 30 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1032_
timestamp 1728341909
transform 1 0 110 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1033_
timestamp 1728341909
transform -1 0 710 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1034_
timestamp 1728341909
transform -1 0 30 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1035_
timestamp 1728341909
transform 1 0 110 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1036_
timestamp 1728341909
transform -1 0 250 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1037_
timestamp 1728341909
transform 1 0 330 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1038_
timestamp 1728341909
transform -1 0 830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1039_
timestamp 1728341909
transform -1 0 30 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1040_
timestamp 1728341909
transform -1 0 1150 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1041_
timestamp 1728341909
transform 1 0 890 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1042_
timestamp 1728341909
transform -1 0 1030 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1043_
timestamp 1728341909
transform -1 0 150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1044_
timestamp 1728341909
transform 1 0 230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1045_
timestamp 1728341909
transform 1 0 1590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1046_
timestamp 1728341909
transform 1 0 1290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1047_
timestamp 1728341909
transform 1 0 890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1048_
timestamp 1728341909
transform -1 0 1110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1050_
timestamp 1728341909
transform 1 0 1670 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1052_
timestamp 1728341909
transform 1 0 1390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1054_
timestamp 1728341909
transform 1 0 1190 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1056_
timestamp 1728341909
transform 1 0 910 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1058_
timestamp 1728341909
transform -1 0 810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1060_
timestamp 1728341909
transform -1 0 590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1062_
timestamp 1728341909
transform -1 0 910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1064_
timestamp 1728341909
transform -1 0 1510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1085_
timestamp 1728341909
transform -1 0 2750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1087_
timestamp 1728341909
transform -1 0 2930 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1089_
timestamp 1728341909
transform -1 0 2610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1091_
timestamp 1728341909
transform 1 0 3170 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1093_
timestamp 1728341909
transform -1 0 3510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1095_
timestamp 1728341909
transform 1 0 3650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1097_
timestamp 1728341909
transform -1 0 3310 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1099_
timestamp 1728341909
transform -1 0 3450 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1100_
timestamp 1728341909
transform -1 0 3470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1101_
timestamp 1728341909
transform 1 0 3770 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1102_
timestamp 1728341909
transform 1 0 3950 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1103_
timestamp 1728341909
transform -1 0 3870 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1104_
timestamp 1728341909
transform -1 0 3390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1105_
timestamp 1728341909
transform 1 0 3230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1106_
timestamp 1728341909
transform 1 0 3950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1107_
timestamp 1728341909
transform -1 0 3810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1108_
timestamp 1728341909
transform 1 0 3670 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1109_
timestamp 1728341909
transform -1 0 3570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1110_
timestamp 1728341909
transform 1 0 2790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1111_
timestamp 1728341909
transform -1 0 3330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1112_
timestamp 1728341909
transform -1 0 2890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1113_
timestamp 1728341909
transform -1 0 2750 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1114_
timestamp 1728341909
transform 1 0 3090 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1115_
timestamp 1728341909
transform -1 0 3010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1116_
timestamp 1728341909
transform -1 0 2910 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1117_
timestamp 1728341909
transform -1 0 3010 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1118_
timestamp 1728341909
transform 1 0 2970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1119_
timestamp 1728341909
transform -1 0 3110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1120_
timestamp 1728341909
transform 1 0 2870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1121_
timestamp 1728341909
transform -1 0 3230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1122_
timestamp 1728341909
transform -1 0 2790 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1123_
timestamp 1728341909
transform 1 0 2990 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1124_
timestamp 1728341909
transform 1 0 2890 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1125_
timestamp 1728341909
transform -1 0 1690 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1126_
timestamp 1728341909
transform 1 0 2790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1127_
timestamp 1728341909
transform -1 0 2650 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1128_
timestamp 1728341909
transform 1 0 2530 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1129_
timestamp 1728341909
transform -1 0 2630 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1130_
timestamp 1728341909
transform 1 0 2030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1131_
timestamp 1728341909
transform -1 0 1970 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1132_
timestamp 1728341909
transform 1 0 1910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1134_
timestamp 1728341909
transform -1 0 830 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1136_
timestamp 1728341909
transform -1 0 1770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1138_
timestamp 1728341909
transform -1 0 1830 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1140_
timestamp 1728341909
transform 1 0 2370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1142_
timestamp 1728341909
transform 1 0 2650 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1144_
timestamp 1728341909
transform -1 0 2650 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1146_
timestamp 1728341909
transform -1 0 2850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1148_
timestamp 1728341909
transform -1 0 1290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1150_
timestamp 1728341909
transform -1 0 1490 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1152_
timestamp 1728341909
transform 1 0 1550 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1154_
timestamp 1728341909
transform 1 0 930 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1156_
timestamp 1728341909
transform 1 0 2250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1158_
timestamp 1728341909
transform -1 0 2530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1160_
timestamp 1728341909
transform -1 0 2390 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1162_
timestamp 1728341909
transform 1 0 3770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1164_
timestamp 1728341909
transform -1 0 3250 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1165_
timestamp 1728341909
transform 1 0 3090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1166_
timestamp 1728341909
transform -1 0 2990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1167_
timestamp 1728341909
transform 1 0 990 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1168_
timestamp 1728341909
transform -1 0 770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1169_
timestamp 1728341909
transform 1 0 5530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1170_
timestamp 1728341909
transform -1 0 310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1171_
timestamp 1728341909
transform 1 0 790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1172_
timestamp 1728341909
transform 1 0 390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1173_
timestamp 1728341909
transform -1 0 210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1174_
timestamp 1728341909
transform -1 0 30 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1175_
timestamp 1728341909
transform 1 0 990 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1176_
timestamp 1728341909
transform -1 0 30 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1177_
timestamp 1728341909
transform -1 0 4830 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1178_
timestamp 1728341909
transform 1 0 450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1179_
timestamp 1728341909
transform -1 0 130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1180_
timestamp 1728341909
transform -1 0 230 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1181_
timestamp 1728341909
transform 1 0 90 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1182_
timestamp 1728341909
transform -1 0 30 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1183_
timestamp 1728341909
transform 1 0 150 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1184_
timestamp 1728341909
transform -1 0 250 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1185_
timestamp 1728341909
transform 1 0 210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1186_
timestamp 1728341909
transform -1 0 350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1187_
timestamp 1728341909
transform 1 0 870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1188_
timestamp 1728341909
transform -1 0 910 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1189_
timestamp 1728341909
transform 1 0 450 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1190_
timestamp 1728341909
transform -1 0 30 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1191_
timestamp 1728341909
transform 1 0 330 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1192_
timestamp 1728341909
transform 1 0 570 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1193_
timestamp 1728341909
transform 1 0 570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1194_
timestamp 1728341909
transform 1 0 470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1195_
timestamp 1728341909
transform 1 0 690 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1196_
timestamp 1728341909
transform 1 0 790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1198_
timestamp 1728341909
transform -1 0 230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1200_
timestamp 1728341909
transform -1 0 350 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1202_
timestamp 1728341909
transform -1 0 2430 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1204_
timestamp 1728341909
transform -1 0 1710 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1206_
timestamp 1728341909
transform -1 0 1410 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1208_
timestamp 1728341909
transform 1 0 1250 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1210_
timestamp 1728341909
transform -1 0 770 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1212_
timestamp 1728341909
transform 1 0 550 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1214_
timestamp 1728341909
transform 1 0 70 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1216_
timestamp 1728341909
transform -1 0 430 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1218_
timestamp 1728341909
transform -1 0 1030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1220_
timestamp 1728341909
transform -1 0 5450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1222_
timestamp 1728341909
transform 1 0 690 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1224_
timestamp 1728341909
transform 1 0 90 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1226_
timestamp 1728341909
transform 1 0 570 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1228_
timestamp 1728341909
transform 1 0 430 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1229_
timestamp 1728341909
transform 1 0 4470 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1230_
timestamp 1728341909
transform -1 0 3970 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1231_
timestamp 1728341909
transform 1 0 3010 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1232_
timestamp 1728341909
transform -1 0 3010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1233_
timestamp 1728341909
transform -1 0 2930 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1234_
timestamp 1728341909
transform 1 0 2810 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1235_
timestamp 1728341909
transform 1 0 2370 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1236_
timestamp 1728341909
transform -1 0 2270 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1237_
timestamp 1728341909
transform -1 0 2450 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1238_
timestamp 1728341909
transform -1 0 2290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1239_
timestamp 1728341909
transform -1 0 4990 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1240_
timestamp 1728341909
transform 1 0 2710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1241_
timestamp 1728341909
transform -1 0 2190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1242_
timestamp 1728341909
transform -1 0 1830 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1243_
timestamp 1728341909
transform -1 0 1910 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1244_
timestamp 1728341909
transform 1 0 5090 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1245_
timestamp 1728341909
transform 1 0 1970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1246_
timestamp 1728341909
transform -1 0 1890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1247_
timestamp 1728341909
transform -1 0 1870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1248_
timestamp 1728341909
transform -1 0 1950 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1249_
timestamp 1728341909
transform -1 0 3130 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1250_
timestamp 1728341909
transform -1 0 2510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1251_
timestamp 1728341909
transform -1 0 2510 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1252_
timestamp 1728341909
transform -1 0 2390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1253_
timestamp 1728341909
transform 1 0 1950 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1254_
timestamp 1728341909
transform -1 0 2070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1255_
timestamp 1728341909
transform 1 0 2710 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1256_
timestamp 1728341909
transform -1 0 2630 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1257_
timestamp 1728341909
transform 1 0 2050 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1258_
timestamp 1728341909
transform 1 0 1610 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1259_
timestamp 1728341909
transform 1 0 2130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1260_
timestamp 1728341909
transform -1 0 570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1261_
timestamp 1728341909
transform 1 0 650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1263_
timestamp 1728341909
transform -1 0 1750 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1265_
timestamp 1728341909
transform 1 0 3910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1267_
timestamp 1728341909
transform -1 0 3830 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1269_
timestamp 1728341909
transform -1 0 3830 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1271_
timestamp 1728341909
transform 1 0 4330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1273_
timestamp 1728341909
transform -1 0 4390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1275_
timestamp 1728341909
transform 1 0 3490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1277_
timestamp 1728341909
transform 1 0 3610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1279_
timestamp 1728341909
transform -1 0 3630 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1281_
timestamp 1728341909
transform 1 0 1030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1283_
timestamp 1728341909
transform 1 0 3090 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1285_
timestamp 1728341909
transform -1 0 1910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1287_
timestamp 1728341909
transform -1 0 1630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1289_
timestamp 1728341909
transform -1 0 1110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1291_
timestamp 1728341909
transform -1 0 3290 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1293_
timestamp 1728341909
transform 1 0 3430 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1294_
timestamp 1728341909
transform -1 0 3570 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1295_
timestamp 1728341909
transform 1 0 3390 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1296_
timestamp 1728341909
transform -1 0 3290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1297_
timestamp 1728341909
transform -1 0 3190 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1298_
timestamp 1728341909
transform -1 0 3270 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1299_
timestamp 1728341909
transform 1 0 1210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1300_
timestamp 1728341909
transform 1 0 650 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1301_
timestamp 1728341909
transform -1 0 790 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1302_
timestamp 1728341909
transform -1 0 3210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1303_
timestamp 1728341909
transform 1 0 2210 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1304_
timestamp 1728341909
transform 1 0 2330 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1305_
timestamp 1728341909
transform 1 0 1110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1306_
timestamp 1728341909
transform 1 0 1070 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1307_
timestamp 1728341909
transform 1 0 1210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1308_
timestamp 1728341909
transform 1 0 2090 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1309_
timestamp 1728341909
transform -1 0 3730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1310_
timestamp 1728341909
transform -1 0 3630 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1311_
timestamp 1728341909
transform 1 0 1450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1312_
timestamp 1728341909
transform 1 0 3370 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1313_
timestamp 1728341909
transform 1 0 3490 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1314_
timestamp 1728341909
transform -1 0 3590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1315_
timestamp 1728341909
transform 1 0 3470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1316_
timestamp 1728341909
transform 1 0 1710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1317_
timestamp 1728341909
transform 1 0 1590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1318_
timestamp 1728341909
transform -1 0 3710 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1319_
timestamp 1728341909
transform 1 0 3330 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1320_
timestamp 1728341909
transform -1 0 3910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1321_
timestamp 1728341909
transform -1 0 3710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1322_
timestamp 1728341909
transform 1 0 3130 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1323_
timestamp 1728341909
transform 1 0 3350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1324_
timestamp 1728341909
transform 1 0 3250 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1325_
timestamp 1728341909
transform -1 0 4370 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1327_
timestamp 1728341909
transform 1 0 4570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1329_
timestamp 1728341909
transform 1 0 3070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1331_
timestamp 1728341909
transform 1 0 4830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1333_
timestamp 1728341909
transform 1 0 3410 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1335_
timestamp 1728341909
transform -1 0 3710 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1337_
timestamp 1728341909
transform 1 0 3190 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1339_
timestamp 1728341909
transform 1 0 3470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1341_
timestamp 1728341909
transform 1 0 2190 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1343_
timestamp 1728341909
transform -1 0 2490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1345_
timestamp 1728341909
transform 1 0 2190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1347_
timestamp 1728341909
transform 1 0 2410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1349_
timestamp 1728341909
transform -1 0 110 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1351_
timestamp 1728341909
transform 1 0 3230 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1353_
timestamp 1728341909
transform 1 0 2350 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1355_
timestamp 1728341909
transform 1 0 1430 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1357_
timestamp 1728341909
transform -1 0 2190 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1358_
timestamp 1728341909
transform 1 0 2150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1359_
timestamp 1728341909
transform 1 0 1570 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1360_
timestamp 1728341909
transform 1 0 1970 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1361_
timestamp 1728341909
transform 1 0 2030 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1362_
timestamp 1728341909
transform 1 0 2090 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1363_
timestamp 1728341909
transform 1 0 590 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1364_
timestamp 1728341909
transform -1 0 30 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1365_
timestamp 1728341909
transform -1 0 30 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1366_
timestamp 1728341909
transform -1 0 350 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1367_
timestamp 1728341909
transform 1 0 1910 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1368_
timestamp 1728341909
transform -1 0 1710 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1369_
timestamp 1728341909
transform 1 0 1770 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1370_
timestamp 1728341909
transform -1 0 2370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1371_
timestamp 1728341909
transform 1 0 2230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1372_
timestamp 1728341909
transform -1 0 2110 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1373_
timestamp 1728341909
transform -1 0 30 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1374_
timestamp 1728341909
transform -1 0 30 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1375_
timestamp 1728341909
transform 1 0 110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1376_
timestamp 1728341909
transform -1 0 150 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1377_
timestamp 1728341909
transform -1 0 30 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1378_
timestamp 1728341909
transform -1 0 30 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1379_
timestamp 1728341909
transform 1 0 870 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1380_
timestamp 1728341909
transform -1 0 1390 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1381_
timestamp 1728341909
transform -1 0 870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1382_
timestamp 1728341909
transform -1 0 1150 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1383_
timestamp 1728341909
transform 1 0 750 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1384_
timestamp 1728341909
transform -1 0 370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1385_
timestamp 1728341909
transform 1 0 810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1386_
timestamp 1728341909
transform -1 0 1270 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1387_
timestamp 1728341909
transform 1 0 230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1388_
timestamp 1728341909
transform 1 0 590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1389_
timestamp 1728341909
transform -1 0 410 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1390_
timestamp 1728341909
transform -1 0 690 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1392_
timestamp 1728341909
transform -1 0 890 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1394_
timestamp 1728341909
transform -1 0 650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1396_
timestamp 1728341909
transform -1 0 1230 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1398_
timestamp 1728341909
transform -1 0 1510 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1400_
timestamp 1728341909
transform 1 0 1950 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1402_
timestamp 1728341909
transform -1 0 2890 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1404_
timestamp 1728341909
transform 1 0 2750 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1406_
timestamp 1728341909
transform 1 0 2210 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1408_
timestamp 1728341909
transform -1 0 470 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1410_
timestamp 1728341909
transform -1 0 790 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1412_
timestamp 1728341909
transform -1 0 510 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1414_
timestamp 1728341909
transform 1 0 230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1416_
timestamp 1728341909
transform -1 0 1130 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1418_
timestamp 1728341909
transform -1 0 2570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1420_
timestamp 1728341909
transform -1 0 2630 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1422_
timestamp 1728341909
transform -1 0 3350 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1423_
timestamp 1728341909
transform 1 0 3210 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1424_
timestamp 1728341909
transform 1 0 3090 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1425_
timestamp 1728341909
transform 1 0 2910 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1426_
timestamp 1728341909
transform 1 0 2850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1427_
timestamp 1728341909
transform -1 0 2190 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1428_
timestamp 1728341909
transform 1 0 3110 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1429_
timestamp 1728341909
transform 1 0 2810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1430_
timestamp 1728341909
transform 1 0 3390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1431_
timestamp 1728341909
transform -1 0 3330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1432_
timestamp 1728341909
transform -1 0 2730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1433_
timestamp 1728341909
transform -1 0 2610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1434_
timestamp 1728341909
transform -1 0 3010 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1435_
timestamp 1728341909
transform 1 0 3190 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1436_
timestamp 1728341909
transform 1 0 3090 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1437_
timestamp 1728341909
transform 1 0 2630 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1438_
timestamp 1728341909
transform -1 0 2530 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1439_
timestamp 1728341909
transform -1 0 1790 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1440_
timestamp 1728341909
transform -1 0 2070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1441_
timestamp 1728341909
transform 1 0 1810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1442_
timestamp 1728341909
transform 1 0 1670 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1443_
timestamp 1728341909
transform 1 0 1710 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1444_
timestamp 1728341909
transform -1 0 1590 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1445_
timestamp 1728341909
transform -1 0 1730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1446_
timestamp 1728341909
transform 1 0 1890 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1447_
timestamp 1728341909
transform -1 0 870 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1448_
timestamp 1728341909
transform 1 0 1050 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1449_
timestamp 1728341909
transform -1 0 970 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1450_
timestamp 1728341909
transform 1 0 1470 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1451_
timestamp 1728341909
transform -1 0 1370 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1452_
timestamp 1728341909
transform -1 0 250 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1453_
timestamp 1728341909
transform 1 0 330 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1454_
timestamp 1728341909
transform -1 0 970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1455_
timestamp 1728341909
transform -1 0 1090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1457_
timestamp 1728341909
transform 1 0 1910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1459_
timestamp 1728341909
transform 1 0 2750 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1461_
timestamp 1728341909
transform 1 0 1470 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1463_
timestamp 1728341909
transform 1 0 1250 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1465_
timestamp 1728341909
transform 1 0 710 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1467_
timestamp 1728341909
transform 1 0 1310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1469_
timestamp 1728341909
transform -1 0 2510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1471_
timestamp 1728341909
transform 1 0 2350 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1473_
timestamp 1728341909
transform -1 0 2130 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1475_
timestamp 1728341909
transform -1 0 1910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1477_
timestamp 1728341909
transform -1 0 2430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1479_
timestamp 1728341909
transform 1 0 2470 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1481_
timestamp 1728341909
transform -1 0 1870 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1483_
timestamp 1728341909
transform 1 0 2010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1485_
timestamp 1728341909
transform 1 0 1670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1487_
timestamp 1728341909
transform 1 0 890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1488_
timestamp 1728341909
transform -1 0 1110 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1489_
timestamp 1728341909
transform 1 0 1290 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1490_
timestamp 1728341909
transform 1 0 1410 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1491_
timestamp 1728341909
transform -1 0 1390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1492_
timestamp 1728341909
transform -1 0 1490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1493_
timestamp 1728341909
transform 1 0 5210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1494_
timestamp 1728341909
transform 1 0 5030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1495_
timestamp 1728341909
transform 1 0 5070 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1496_
timestamp 1728341909
transform 1 0 5150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1497_
timestamp 1728341909
transform -1 0 1710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1498_
timestamp 1728341909
transform -1 0 1770 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1499_
timestamp 1728341909
transform 1 0 1790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1500_
timestamp 1728341909
transform 1 0 2150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1501_
timestamp 1728341909
transform 1 0 1250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1502_
timestamp 1728341909
transform 1 0 2470 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1503_
timestamp 1728341909
transform 1 0 5330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1504_
timestamp 1728341909
transform 1 0 4970 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1505_
timestamp 1728341909
transform -1 0 5130 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1506_
timestamp 1728341909
transform 1 0 4690 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1507_
timestamp 1728341909
transform -1 0 4910 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1508_
timestamp 1728341909
transform 1 0 4790 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1509_
timestamp 1728341909
transform -1 0 4930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1510_
timestamp 1728341909
transform -1 0 4810 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1511_
timestamp 1728341909
transform -1 0 4690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1512_
timestamp 1728341909
transform 1 0 4550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1513_
timestamp 1728341909
transform 1 0 4990 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1514_
timestamp 1728341909
transform -1 0 5490 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1515_
timestamp 1728341909
transform 1 0 5630 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1516_
timestamp 1728341909
transform 1 0 5630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1517_
timestamp 1728341909
transform 1 0 5570 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1518_
timestamp 1728341909
transform 1 0 5490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1519_
timestamp 1728341909
transform -1 0 5610 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1521_
timestamp 1728341909
transform 1 0 5170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1523_
timestamp 1728341909
transform 1 0 2250 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1525_
timestamp 1728341909
transform 1 0 1930 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1527_
timestamp 1728341909
transform -1 0 2290 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1529_
timestamp 1728341909
transform -1 0 4890 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1531_
timestamp 1728341909
transform -1 0 5010 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1533_
timestamp 1728341909
transform 1 0 5110 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1535_
timestamp 1728341909
transform 1 0 5510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1537_
timestamp 1728341909
transform 1 0 5170 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1539_
timestamp 1728341909
transform -1 0 5010 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1541_
timestamp 1728341909
transform 1 0 5570 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1543_
timestamp 1728341909
transform 1 0 5230 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1545_
timestamp 1728341909
transform 1 0 5610 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1547_
timestamp 1728341909
transform -1 0 5270 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1549_
timestamp 1728341909
transform 1 0 5110 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1551_
timestamp 1728341909
transform 1 0 4870 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1552_
timestamp 1728341909
transform -1 0 4790 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1553_
timestamp 1728341909
transform 1 0 5490 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1554_
timestamp 1728341909
transform 1 0 5390 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1555_
timestamp 1728341909
transform -1 0 5290 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1556_
timestamp 1728341909
transform 1 0 5050 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1557_
timestamp 1728341909
transform 1 0 5610 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1558_
timestamp 1728341909
transform -1 0 4590 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1559_
timestamp 1728341909
transform 1 0 4670 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1560_
timestamp 1728341909
transform 1 0 5570 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1561_
timestamp 1728341909
transform -1 0 5090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1562_
timestamp 1728341909
transform -1 0 4990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1563_
timestamp 1728341909
transform 1 0 5110 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1564_
timestamp 1728341909
transform -1 0 5630 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1565_
timestamp 1728341909
transform -1 0 5230 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1566_
timestamp 1728341909
transform -1 0 5010 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1567_
timestamp 1728341909
transform -1 0 4890 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1568_
timestamp 1728341909
transform 1 0 4750 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1569_
timestamp 1728341909
transform 1 0 5090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1570_
timestamp 1728341909
transform -1 0 4910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1571_
timestamp 1728341909
transform 1 0 4990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1572_
timestamp 1728341909
transform 1 0 5330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1573_
timestamp 1728341909
transform 1 0 5410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1574_
timestamp 1728341909
transform -1 0 5350 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1575_
timestamp 1728341909
transform -1 0 5230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1576_
timestamp 1728341909
transform -1 0 4990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1577_
timestamp 1728341909
transform 1 0 4290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1578_
timestamp 1728341909
transform -1 0 5470 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1579_
timestamp 1728341909
transform -1 0 4710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1580_
timestamp 1728341909
transform 1 0 4790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1581_
timestamp 1728341909
transform -1 0 4890 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1582_
timestamp 1728341909
transform -1 0 4990 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1583_
timestamp 1728341909
transform -1 0 5110 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1584_
timestamp 1728341909
transform -1 0 3970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1586_
timestamp 1728341909
transform -1 0 3850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1588_
timestamp 1728341909
transform -1 0 2970 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1590_
timestamp 1728341909
transform 1 0 2950 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1592_
timestamp 1728341909
transform 1 0 1350 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1594_
timestamp 1728341909
transform 1 0 3210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1596_
timestamp 1728341909
transform -1 0 2990 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1598_
timestamp 1728341909
transform 1 0 210 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1600_
timestamp 1728341909
transform -1 0 30 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1602_
timestamp 1728341909
transform 1 0 3750 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1604_
timestamp 1728341909
transform 1 0 1110 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1606_
timestamp 1728341909
transform 1 0 630 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1608_
timestamp 1728341909
transform -1 0 1030 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1610_
timestamp 1728341909
transform 1 0 870 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1612_
timestamp 1728341909
transform 1 0 550 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1614_
timestamp 1728341909
transform -1 0 890 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1616_
timestamp 1728341909
transform 1 0 990 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1617_
timestamp 1728341909
transform -1 0 1010 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1618_
timestamp 1728341909
transform 1 0 870 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1619_
timestamp 1728341909
transform -1 0 630 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1620_
timestamp 1728341909
transform -1 0 510 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1621_
timestamp 1728341909
transform -1 0 1190 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1622_
timestamp 1728341909
transform -1 0 1930 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1623_
timestamp 1728341909
transform -1 0 2150 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1624_
timestamp 1728341909
transform 1 0 2010 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1625_
timestamp 1728341909
transform -1 0 1830 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1626_
timestamp 1728341909
transform 1 0 1690 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1627_
timestamp 1728341909
transform 1 0 2470 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1628_
timestamp 1728341909
transform -1 0 3510 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1629_
timestamp 1728341909
transform -1 0 3730 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1630_
timestamp 1728341909
transform 1 0 3590 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1631_
timestamp 1728341909
transform 1 0 3810 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1632_
timestamp 1728341909
transform -1 0 2270 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1633_
timestamp 1728341909
transform -1 0 2890 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1634_
timestamp 1728341909
transform -1 0 2790 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1635_
timestamp 1728341909
transform 1 0 2650 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1636_
timestamp 1728341909
transform 1 0 4710 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1637_
timestamp 1728341909
transform 1 0 4610 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1638_
timestamp 1728341909
transform 1 0 4390 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1639_
timestamp 1728341909
transform 1 0 4510 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1640_
timestamp 1728341909
transform 1 0 2190 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1641_
timestamp 1728341909
transform 1 0 2290 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1642_
timestamp 1728341909
transform 1 0 3210 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1643_
timestamp 1728341909
transform 1 0 3290 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1644_
timestamp 1728341909
transform -1 0 2770 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1645_
timestamp 1728341909
transform 1 0 2630 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1646_
timestamp 1728341909
transform -1 0 2990 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1647_
timestamp 1728341909
transform 1 0 3110 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1648_
timestamp 1728341909
transform -1 0 3110 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1650_
timestamp 1728341909
transform -1 0 2410 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1652_
timestamp 1728341909
transform -1 0 4250 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1654_
timestamp 1728341909
transform -1 0 4430 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1656_
timestamp 1728341909
transform 1 0 4730 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1658_
timestamp 1728341909
transform -1 0 4290 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1660_
timestamp 1728341909
transform -1 0 4090 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1662_
timestamp 1728341909
transform 1 0 3610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1664_
timestamp 1728341909
transform 1 0 3390 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1666_
timestamp 1728341909
transform -1 0 4010 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1668_
timestamp 1728341909
transform 1 0 3890 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1670_
timestamp 1728341909
transform -1 0 4730 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1672_
timestamp 1728341909
transform -1 0 4610 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1674_
timestamp 1728341909
transform -1 0 4030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1676_
timestamp 1728341909
transform 1 0 3450 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1678_
timestamp 1728341909
transform 1 0 3790 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1680_
timestamp 1728341909
transform 1 0 1290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1681_
timestamp 1728341909
transform 1 0 1790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1682_
timestamp 1728341909
transform 1 0 1570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1683_
timestamp 1728341909
transform -1 0 1530 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1684_
timestamp 1728341909
transform 1 0 1590 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1685_
timestamp 1728341909
transform 1 0 1590 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1686_
timestamp 1728341909
transform 1 0 1790 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1687_
timestamp 1728341909
transform -1 0 1710 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1688_
timestamp 1728341909
transform 1 0 1470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1689_
timestamp 1728341909
transform 1 0 950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1690_
timestamp 1728341909
transform 1 0 1150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1691_
timestamp 1728341909
transform 1 0 710 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1692_
timestamp 1728341909
transform 1 0 1290 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1693_
timestamp 1728341909
transform 1 0 1230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1694_
timestamp 1728341909
transform -1 0 1390 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1695_
timestamp 1728341909
transform 1 0 4590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1696_
timestamp 1728341909
transform 1 0 4110 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1697_
timestamp 1728341909
transform 1 0 4990 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1698_
timestamp 1728341909
transform 1 0 4810 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1699_
timestamp 1728341909
transform 1 0 5110 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1700_
timestamp 1728341909
transform -1 0 3350 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1701_
timestamp 1728341909
transform 1 0 3430 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1702_
timestamp 1728341909
transform -1 0 3550 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1703_
timestamp 1728341909
transform 1 0 4350 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1704_
timestamp 1728341909
transform 1 0 4250 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1705_
timestamp 1728341909
transform -1 0 4390 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1706_
timestamp 1728341909
transform 1 0 4490 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1707_
timestamp 1728341909
transform 1 0 4710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1708_
timestamp 1728341909
transform 1 0 710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1709_
timestamp 1728341909
transform -1 0 1070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1710_
timestamp 1728341909
transform 1 0 1350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1711_
timestamp 1728341909
transform -1 0 1690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1712_
timestamp 1728341909
transform -1 0 1730 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1713_
timestamp 1728341909
transform 1 0 4450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1715_
timestamp 1728341909
transform 1 0 4530 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1717_
timestamp 1728341909
transform -1 0 2430 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1719_
timestamp 1728341909
transform -1 0 590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1721_
timestamp 1728341909
transform 1 0 90 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1723_
timestamp 1728341909
transform 1 0 450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1725_
timestamp 1728341909
transform -1 0 1250 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1727_
timestamp 1728341909
transform 1 0 810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1729_
timestamp 1728341909
transform -1 0 130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1731_
timestamp 1728341909
transform 1 0 210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1733_
timestamp 1728341909
transform 1 0 2810 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1735_
timestamp 1728341909
transform 1 0 2050 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1737_
timestamp 1728341909
transform 1 0 2550 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1739_
timestamp 1728341909
transform -1 0 2450 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1741_
timestamp 1728341909
transform -1 0 510 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1743_
timestamp 1728341909
transform -1 0 1010 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1745_
timestamp 1728341909
transform 1 0 1050 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1746_
timestamp 1728341909
transform 1 0 1530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1747_
timestamp 1728341909
transform -1 0 1630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1748_
timestamp 1728341909
transform -1 0 2870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1749_
timestamp 1728341909
transform -1 0 3010 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1750_
timestamp 1728341909
transform 1 0 2990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1751_
timestamp 1728341909
transform -1 0 3650 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1752_
timestamp 1728341909
transform -1 0 3730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1753_
timestamp 1728341909
transform 1 0 3350 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1754_
timestamp 1728341909
transform -1 0 2930 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1755_
timestamp 1728341909
transform -1 0 2830 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1756_
timestamp 1728341909
transform 1 0 3030 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1757_
timestamp 1728341909
transform 1 0 3490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1758_
timestamp 1728341909
transform 1 0 3410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1759_
timestamp 1728341909
transform -1 0 3310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1760_
timestamp 1728341909
transform 1 0 3770 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1761_
timestamp 1728341909
transform -1 0 4190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1762_
timestamp 1728341909
transform -1 0 4110 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1763_
timestamp 1728341909
transform 1 0 4190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1764_
timestamp 1728341909
transform 1 0 4110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1765_
timestamp 1728341909
transform 1 0 4030 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1766_
timestamp 1728341909
transform 1 0 3670 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1767_
timestamp 1728341909
transform 1 0 4130 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1768_
timestamp 1728341909
transform 1 0 4690 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1769_
timestamp 1728341909
transform 1 0 4590 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1770_
timestamp 1728341909
transform -1 0 4490 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1771_
timestamp 1728341909
transform -1 0 4250 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1772_
timestamp 1728341909
transform -1 0 3930 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1773_
timestamp 1728341909
transform 1 0 4230 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1774_
timestamp 1728341909
transform -1 0 4270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1775_
timestamp 1728341909
transform -1 0 4210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1776_
timestamp 1728341909
transform -1 0 4430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1777_
timestamp 1728341909
transform -1 0 4430 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1778_
timestamp 1728341909
transform -1 0 2610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1780_
timestamp 1728341909
transform -1 0 930 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1782_
timestamp 1728341909
transform 1 0 1110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1784_
timestamp 1728341909
transform -1 0 2730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1786_
timestamp 1728341909
transform -1 0 2470 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1788_
timestamp 1728341909
transform 1 0 2930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1790_
timestamp 1728341909
transform -1 0 3430 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1792_
timestamp 1728341909
transform 1 0 3090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1794_
timestamp 1728341909
transform 1 0 3490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1796_
timestamp 1728341909
transform -1 0 4290 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1798_
timestamp 1728341909
transform 1 0 4270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1800_
timestamp 1728341909
transform 1 0 4410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1802_
timestamp 1728341909
transform 1 0 3790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1804_
timestamp 1728341909
transform -1 0 3690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1806_
timestamp 1728341909
transform 1 0 4690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1808_
timestamp 1728341909
transform -1 0 4810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1810_
timestamp 1728341909
transform 1 0 4050 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1811_
timestamp 1728341909
transform -1 0 3890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1812_
timestamp 1728341909
transform -1 0 4470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1813_
timestamp 1728341909
transform 1 0 4070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1814_
timestamp 1728341909
transform -1 0 3930 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1815_
timestamp 1728341909
transform 1 0 3450 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1816_
timestamp 1728341909
transform 1 0 3710 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1817_
timestamp 1728341909
transform -1 0 3730 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1818_
timestamp 1728341909
transform 1 0 3770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1819_
timestamp 1728341909
transform 1 0 3970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1820_
timestamp 1728341909
transform -1 0 3890 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1821_
timestamp 1728341909
transform 1 0 4030 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1822_
timestamp 1728341909
transform 1 0 4190 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1823_
timestamp 1728341909
transform 1 0 4650 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1824_
timestamp 1728341909
transform -1 0 4350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1825_
timestamp 1728341909
transform -1 0 4570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1826_
timestamp 1728341909
transform -1 0 4990 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1827_
timestamp 1728341909
transform 1 0 5550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1828_
timestamp 1728341909
transform -1 0 5490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1829_
timestamp 1728341909
transform 1 0 5530 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1830_
timestamp 1728341909
transform -1 0 5450 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1831_
timestamp 1728341909
transform -1 0 4870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1832_
timestamp 1728341909
transform -1 0 4450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1833_
timestamp 1728341909
transform 1 0 4190 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1834_
timestamp 1728341909
transform -1 0 4170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1835_
timestamp 1728341909
transform -1 0 4050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1836_
timestamp 1728341909
transform 1 0 3830 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1837_
timestamp 1728341909
transform 1 0 3730 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1838_
timestamp 1728341909
transform 1 0 3950 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1839_
timestamp 1728341909
transform 1 0 4270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1840_
timestamp 1728341909
transform -1 0 4710 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1841_
timestamp 1728341909
transform 1 0 4750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1842_
timestamp 1728341909
transform 1 0 4390 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1844_
timestamp 1728341909
transform 1 0 4350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1846_
timestamp 1728341909
transform -1 0 4170 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1848_
timestamp 1728341909
transform 1 0 4930 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1850_
timestamp 1728341909
transform 1 0 4770 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1852_
timestamp 1728341909
transform -1 0 5070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1854_
timestamp 1728341909
transform 1 0 5370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1856_
timestamp 1728341909
transform 1 0 5210 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1858_
timestamp 1728341909
transform -1 0 3930 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1860_
timestamp 1728341909
transform 1 0 3890 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1862_
timestamp 1728341909
transform -1 0 3830 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1864_
timestamp 1728341909
transform 1 0 4030 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1866_
timestamp 1728341909
transform 1 0 3670 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1868_
timestamp 1728341909
transform 1 0 4230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1870_
timestamp 1728341909
transform 1 0 4010 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1872_
timestamp 1728341909
transform 1 0 4130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1874_
timestamp 1728341909
transform 1 0 4270 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1875_
timestamp 1728341909
transform 1 0 5090 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1876_
timestamp 1728341909
transform 1 0 5330 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1877_
timestamp 1728341909
transform 1 0 4790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1878_
timestamp 1728341909
transform -1 0 4730 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1879_
timestamp 1728341909
transform -1 0 4610 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1880_
timestamp 1728341909
transform -1 0 4490 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1881_
timestamp 1728341909
transform -1 0 4370 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1882_
timestamp 1728341909
transform -1 0 4510 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1883_
timestamp 1728341909
transform 1 0 4350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1884_
timestamp 1728341909
transform 1 0 4470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1885_
timestamp 1728341909
transform 1 0 5550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1886_
timestamp 1728341909
transform 1 0 5210 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1887_
timestamp 1728341909
transform 1 0 5430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1888_
timestamp 1728341909
transform -1 0 4550 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1889_
timestamp 1728341909
transform -1 0 4170 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1890_
timestamp 1728341909
transform 1 0 4410 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1891_
timestamp 1728341909
transform 1 0 5530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1892_
timestamp 1728341909
transform 1 0 5290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1893_
timestamp 1728341909
transform 1 0 5410 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1894_
timestamp 1728341909
transform -1 0 5110 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1895_
timestamp 1728341909
transform -1 0 4930 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1896_
timestamp 1728341909
transform 1 0 5010 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1897_
timestamp 1728341909
transform -1 0 5070 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1898_
timestamp 1728341909
transform -1 0 4850 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1899_
timestamp 1728341909
transform 1 0 4930 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1900_
timestamp 1728341909
transform 1 0 4490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1901_
timestamp 1728341909
transform -1 0 4390 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1902_
timestamp 1728341909
transform -1 0 4090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1903_
timestamp 1728341909
transform -1 0 4210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1904_
timestamp 1728341909
transform 1 0 3970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1905_
timestamp 1728341909
transform -1 0 5030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1906_
timestamp 1728341909
transform -1 0 4590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1907_
timestamp 1728341909
transform -1 0 4630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1942_
timestamp 1728341909
transform 1 0 3770 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1944_
timestamp 1728341909
transform 1 0 3370 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert1
timestamp 1728341909
transform 1 0 1430 0 1 3610
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert3
timestamp 1728341909
transform 1 0 2270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert11
timestamp 1728341909
transform 1 0 5090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert13
timestamp 1728341909
transform 1 0 4750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert15
timestamp 1728341909
transform -1 0 1750 0 1 2170
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert5
timestamp 1728341909
transform -1 0 4610 0 1 3610
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert7
timestamp 1728341909
transform -1 0 2570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1728341909
transform 1 0 4850 0 1 250
box -12 -8 32 252
use FILL  FILL_1__945_
timestamp 1728341909
transform 1 0 1590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__947_
timestamp 1728341909
transform 1 0 1910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__949_
timestamp 1728341909
transform 1 0 3150 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__951_
timestamp 1728341909
transform 1 0 2570 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__953_
timestamp 1728341909
transform 1 0 3170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__955_
timestamp 1728341909
transform 1 0 2430 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__957_
timestamp 1728341909
transform -1 0 2330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__959_
timestamp 1728341909
transform 1 0 2050 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__961_
timestamp 1728341909
transform 1 0 2430 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__963_
timestamp 1728341909
transform 1 0 3490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__965_
timestamp 1728341909
transform -1 0 1730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__967_
timestamp 1728341909
transform 1 0 3450 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__969_
timestamp 1728341909
transform -1 0 2430 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__971_
timestamp 1728341909
transform -1 0 1390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1000_
timestamp 1728341909
transform 1 0 2050 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1002_
timestamp 1728341909
transform 1 0 2390 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1004_
timestamp 1728341909
transform -1 0 1470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1006_
timestamp 1728341909
transform -1 0 2610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1008_
timestamp 1728341909
transform 1 0 3150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1010_
timestamp 1728341909
transform 1 0 3350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1012_
timestamp 1728341909
transform 1 0 3210 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1014_
timestamp 1728341909
transform 1 0 2810 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1016_
timestamp 1728341909
transform 1 0 2950 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1048_
timestamp 1728341909
transform -1 0 1130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1050_
timestamp 1728341909
transform 1 0 1690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1052_
timestamp 1728341909
transform 1 0 1410 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1054_
timestamp 1728341909
transform 1 0 1210 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1056_
timestamp 1728341909
transform 1 0 930 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1058_
timestamp 1728341909
transform -1 0 830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1060_
timestamp 1728341909
transform -1 0 610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1062_
timestamp 1728341909
transform -1 0 930 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1064_
timestamp 1728341909
transform -1 0 1530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1085_
timestamp 1728341909
transform -1 0 2770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1087_
timestamp 1728341909
transform -1 0 2950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1089_
timestamp 1728341909
transform -1 0 2630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1091_
timestamp 1728341909
transform 1 0 3190 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1093_
timestamp 1728341909
transform -1 0 3530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1095_
timestamp 1728341909
transform 1 0 3670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1097_
timestamp 1728341909
transform -1 0 3330 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1099_
timestamp 1728341909
transform -1 0 3470 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1132_
timestamp 1728341909
transform 1 0 1930 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1134_
timestamp 1728341909
transform -1 0 850 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1136_
timestamp 1728341909
transform -1 0 1790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1138_
timestamp 1728341909
transform -1 0 1850 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1140_
timestamp 1728341909
transform 1 0 2390 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1142_
timestamp 1728341909
transform 1 0 2670 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1144_
timestamp 1728341909
transform -1 0 2670 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1146_
timestamp 1728341909
transform -1 0 2870 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1148_
timestamp 1728341909
transform -1 0 1310 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1150_
timestamp 1728341909
transform -1 0 1510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1152_
timestamp 1728341909
transform 1 0 1570 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1154_
timestamp 1728341909
transform 1 0 950 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1156_
timestamp 1728341909
transform 1 0 2270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1158_
timestamp 1728341909
transform -1 0 2550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1160_
timestamp 1728341909
transform -1 0 2410 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1162_
timestamp 1728341909
transform 1 0 3790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1164_
timestamp 1728341909
transform -1 0 3270 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1196_
timestamp 1728341909
transform 1 0 810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1198_
timestamp 1728341909
transform -1 0 250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1200_
timestamp 1728341909
transform -1 0 370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1202_
timestamp 1728341909
transform -1 0 2450 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1204_
timestamp 1728341909
transform -1 0 1730 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1206_
timestamp 1728341909
transform -1 0 1430 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1208_
timestamp 1728341909
transform 1 0 1270 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1210_
timestamp 1728341909
transform -1 0 790 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1212_
timestamp 1728341909
transform 1 0 570 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1214_
timestamp 1728341909
transform 1 0 90 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1216_
timestamp 1728341909
transform -1 0 450 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1218_
timestamp 1728341909
transform -1 0 1050 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1220_
timestamp 1728341909
transform -1 0 5470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1222_
timestamp 1728341909
transform 1 0 710 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1224_
timestamp 1728341909
transform 1 0 110 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1226_
timestamp 1728341909
transform 1 0 590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1228_
timestamp 1728341909
transform 1 0 450 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1261_
timestamp 1728341909
transform 1 0 670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1263_
timestamp 1728341909
transform -1 0 1770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1265_
timestamp 1728341909
transform 1 0 3930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1267_
timestamp 1728341909
transform -1 0 3850 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1269_
timestamp 1728341909
transform -1 0 3850 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1271_
timestamp 1728341909
transform 1 0 4350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1273_
timestamp 1728341909
transform -1 0 4410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1275_
timestamp 1728341909
transform 1 0 3510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1277_
timestamp 1728341909
transform 1 0 3630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1279_
timestamp 1728341909
transform -1 0 3650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1281_
timestamp 1728341909
transform 1 0 1050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1283_
timestamp 1728341909
transform 1 0 3110 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1285_
timestamp 1728341909
transform -1 0 1930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1287_
timestamp 1728341909
transform -1 0 1650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1289_
timestamp 1728341909
transform -1 0 1130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1291_
timestamp 1728341909
transform -1 0 3310 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1293_
timestamp 1728341909
transform 1 0 3450 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1325_
timestamp 1728341909
transform -1 0 4390 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1327_
timestamp 1728341909
transform 1 0 4590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1329_
timestamp 1728341909
transform 1 0 3090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1331_
timestamp 1728341909
transform 1 0 4850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1333_
timestamp 1728341909
transform 1 0 3430 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1335_
timestamp 1728341909
transform -1 0 3730 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1337_
timestamp 1728341909
transform 1 0 3210 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1339_
timestamp 1728341909
transform 1 0 3490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1341_
timestamp 1728341909
transform 1 0 2210 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1343_
timestamp 1728341909
transform -1 0 2510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1345_
timestamp 1728341909
transform 1 0 2210 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1347_
timestamp 1728341909
transform 1 0 2430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1349_
timestamp 1728341909
transform -1 0 130 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1351_
timestamp 1728341909
transform 1 0 3250 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1353_
timestamp 1728341909
transform 1 0 2370 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1355_
timestamp 1728341909
transform 1 0 1450 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1357_
timestamp 1728341909
transform -1 0 2210 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1390_
timestamp 1728341909
transform -1 0 710 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1392_
timestamp 1728341909
transform -1 0 910 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1394_
timestamp 1728341909
transform -1 0 670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1396_
timestamp 1728341909
transform -1 0 1250 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1398_
timestamp 1728341909
transform -1 0 1530 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1400_
timestamp 1728341909
transform 1 0 1970 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1402_
timestamp 1728341909
transform -1 0 2910 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1404_
timestamp 1728341909
transform 1 0 2770 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1406_
timestamp 1728341909
transform 1 0 2230 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1408_
timestamp 1728341909
transform -1 0 490 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1410_
timestamp 1728341909
transform -1 0 810 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1412_
timestamp 1728341909
transform -1 0 530 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1414_
timestamp 1728341909
transform 1 0 250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1416_
timestamp 1728341909
transform -1 0 1150 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1418_
timestamp 1728341909
transform -1 0 2590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1420_
timestamp 1728341909
transform -1 0 2650 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1422_
timestamp 1728341909
transform -1 0 3370 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1455_
timestamp 1728341909
transform -1 0 1110 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1457_
timestamp 1728341909
transform 1 0 1930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1459_
timestamp 1728341909
transform 1 0 2770 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1461_
timestamp 1728341909
transform 1 0 1490 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1463_
timestamp 1728341909
transform 1 0 1270 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1465_
timestamp 1728341909
transform 1 0 730 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1467_
timestamp 1728341909
transform 1 0 1330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1469_
timestamp 1728341909
transform -1 0 2530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1471_
timestamp 1728341909
transform 1 0 2370 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1473_
timestamp 1728341909
transform -1 0 2150 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1475_
timestamp 1728341909
transform -1 0 1930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1477_
timestamp 1728341909
transform -1 0 2450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1479_
timestamp 1728341909
transform 1 0 2490 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1481_
timestamp 1728341909
transform -1 0 1890 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1483_
timestamp 1728341909
transform 1 0 2030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1485_
timestamp 1728341909
transform 1 0 1690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1487_
timestamp 1728341909
transform 1 0 910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1519_
timestamp 1728341909
transform -1 0 5630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1521_
timestamp 1728341909
transform 1 0 5190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1523_
timestamp 1728341909
transform 1 0 2270 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1525_
timestamp 1728341909
transform 1 0 1950 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1527_
timestamp 1728341909
transform -1 0 2310 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1529_
timestamp 1728341909
transform -1 0 4910 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1531_
timestamp 1728341909
transform -1 0 5030 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1533_
timestamp 1728341909
transform 1 0 5130 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1535_
timestamp 1728341909
transform 1 0 5530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1537_
timestamp 1728341909
transform 1 0 5190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1539_
timestamp 1728341909
transform -1 0 5030 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1541_
timestamp 1728341909
transform 1 0 5590 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1543_
timestamp 1728341909
transform 1 0 5250 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1545_
timestamp 1728341909
transform 1 0 5630 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1547_
timestamp 1728341909
transform -1 0 5290 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1549_
timestamp 1728341909
transform 1 0 5130 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1551_
timestamp 1728341909
transform 1 0 4890 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1584_
timestamp 1728341909
transform -1 0 3990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1586_
timestamp 1728341909
transform -1 0 3870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1588_
timestamp 1728341909
transform -1 0 2990 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1590_
timestamp 1728341909
transform 1 0 2970 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1592_
timestamp 1728341909
transform 1 0 1370 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1594_
timestamp 1728341909
transform 1 0 3230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1596_
timestamp 1728341909
transform -1 0 3010 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1598_
timestamp 1728341909
transform 1 0 230 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1600_
timestamp 1728341909
transform -1 0 50 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1602_
timestamp 1728341909
transform 1 0 3770 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1604_
timestamp 1728341909
transform 1 0 1130 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1606_
timestamp 1728341909
transform 1 0 650 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1608_
timestamp 1728341909
transform -1 0 1050 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1610_
timestamp 1728341909
transform 1 0 890 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1612_
timestamp 1728341909
transform 1 0 570 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1614_
timestamp 1728341909
transform -1 0 910 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1616_
timestamp 1728341909
transform 1 0 1010 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1648_
timestamp 1728341909
transform -1 0 3130 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1650_
timestamp 1728341909
transform -1 0 2430 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1652_
timestamp 1728341909
transform -1 0 4270 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1654_
timestamp 1728341909
transform -1 0 4450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1656_
timestamp 1728341909
transform 1 0 4750 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1658_
timestamp 1728341909
transform -1 0 4310 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1660_
timestamp 1728341909
transform -1 0 4110 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1662_
timestamp 1728341909
transform 1 0 3630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1664_
timestamp 1728341909
transform 1 0 3410 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1666_
timestamp 1728341909
transform -1 0 4030 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1668_
timestamp 1728341909
transform 1 0 3910 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1670_
timestamp 1728341909
transform -1 0 4750 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1672_
timestamp 1728341909
transform -1 0 4630 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1674_
timestamp 1728341909
transform -1 0 4050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1676_
timestamp 1728341909
transform 1 0 3470 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1678_
timestamp 1728341909
transform 1 0 3810 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1680_
timestamp 1728341909
transform 1 0 1310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1713_
timestamp 1728341909
transform 1 0 4470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1715_
timestamp 1728341909
transform 1 0 4550 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1717_
timestamp 1728341909
transform -1 0 2450 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1719_
timestamp 1728341909
transform -1 0 610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1721_
timestamp 1728341909
transform 1 0 110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1723_
timestamp 1728341909
transform 1 0 470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1725_
timestamp 1728341909
transform -1 0 1270 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1727_
timestamp 1728341909
transform 1 0 830 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1729_
timestamp 1728341909
transform -1 0 150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1731_
timestamp 1728341909
transform 1 0 230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1733_
timestamp 1728341909
transform 1 0 2830 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1735_
timestamp 1728341909
transform 1 0 2070 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1737_
timestamp 1728341909
transform 1 0 2570 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1739_
timestamp 1728341909
transform -1 0 2470 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1741_
timestamp 1728341909
transform -1 0 530 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1743_
timestamp 1728341909
transform -1 0 1030 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1745_
timestamp 1728341909
transform 1 0 1070 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1778_
timestamp 1728341909
transform -1 0 2630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1780_
timestamp 1728341909
transform -1 0 950 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1782_
timestamp 1728341909
transform 1 0 1130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1784_
timestamp 1728341909
transform -1 0 2750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1786_
timestamp 1728341909
transform -1 0 2490 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1788_
timestamp 1728341909
transform 1 0 2950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1790_
timestamp 1728341909
transform -1 0 3450 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1792_
timestamp 1728341909
transform 1 0 3110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1794_
timestamp 1728341909
transform 1 0 3510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1796_
timestamp 1728341909
transform -1 0 4310 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1798_
timestamp 1728341909
transform 1 0 4290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1800_
timestamp 1728341909
transform 1 0 4430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1802_
timestamp 1728341909
transform 1 0 3810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1804_
timestamp 1728341909
transform -1 0 3710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1806_
timestamp 1728341909
transform 1 0 4710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1808_
timestamp 1728341909
transform -1 0 4830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1810_
timestamp 1728341909
transform 1 0 4070 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1842_
timestamp 1728341909
transform 1 0 4410 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1844_
timestamp 1728341909
transform 1 0 4370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1846_
timestamp 1728341909
transform -1 0 4190 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1848_
timestamp 1728341909
transform 1 0 4950 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1850_
timestamp 1728341909
transform 1 0 4790 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1852_
timestamp 1728341909
transform -1 0 5090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1854_
timestamp 1728341909
transform 1 0 5390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1856_
timestamp 1728341909
transform 1 0 5230 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1858_
timestamp 1728341909
transform -1 0 3950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1860_
timestamp 1728341909
transform 1 0 3910 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1862_
timestamp 1728341909
transform -1 0 3850 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1864_
timestamp 1728341909
transform 1 0 4050 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1866_
timestamp 1728341909
transform 1 0 3690 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1868_
timestamp 1728341909
transform 1 0 4250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1870_
timestamp 1728341909
transform 1 0 4030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1872_
timestamp 1728341909
transform 1 0 4150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1874_
timestamp 1728341909
transform 1 0 4290 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1907_
timestamp 1728341909
transform -1 0 4650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1942_
timestamp 1728341909
transform 1 0 3790 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1944_
timestamp 1728341909
transform 1 0 3390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert1
timestamp 1728341909
transform 1 0 1450 0 1 3610
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert3
timestamp 1728341909
transform 1 0 2290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert11
timestamp 1728341909
transform 1 0 5110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert13
timestamp 1728341909
transform 1 0 4770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert15
timestamp 1728341909
transform -1 0 1770 0 1 2170
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert5
timestamp 1728341909
transform -1 0 4630 0 1 3610
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert7
timestamp 1728341909
transform -1 0 2590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1728341909
transform 1 0 4870 0 1 250
box -12 -8 32 252
<< labels >>
flabel metal1 s 5762 2 5822 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 2737 5577 2743 5583 3 FreeSans 16 90 0 0 clk
port 2 nsew
flabel metal2 s 3097 5577 3103 5583 3 FreeSans 16 90 0 0 down
port 3 nsew
flabel metal2 s 2777 5577 2783 5583 3 FreeSans 16 90 0 0 enable
port 4 nsew
flabel metal2 s 3637 -23 3643 -17 7 FreeSans 16 270 0 0 hsync
port 5 nsew
flabel metal2 s 3837 -23 3843 -17 7 FreeSans 16 270 0 0 p_tick
port 6 nsew
flabel metal2 s 2817 5577 2823 5583 3 FreeSans 16 90 0 0 reset
port 7 nsew
flabel metal2 s 3557 -23 3563 -17 7 FreeSans 16 270 0 0 rgb
port 8 nsew
flabel metal2 s 3137 5577 3143 5583 3 FreeSans 16 90 0 0 up
port 9 nsew
flabel metal2 s 3597 -23 3603 -17 7 FreeSans 16 270 0 0 vsync
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 5760 5580
<< end >>
