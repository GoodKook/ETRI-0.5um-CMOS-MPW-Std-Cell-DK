magic
tech scmos
magscale 1 2
timestamp 1727733579
<< nwell >>
rect -12 134 92 252
<< ntransistor >>
rect 22 14 26 54
rect 32 14 36 54
<< ptransistor >>
rect 20 186 24 226
rect 40 186 44 226
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 32 54
rect 36 14 38 54
<< pdiffusion >>
rect 18 186 20 226
rect 24 186 26 226
rect 38 186 40 226
rect 44 186 46 226
<< ndcontact >>
rect 8 14 20 54
rect 38 14 50 54
<< pdcontact >>
rect 6 186 18 226
rect 26 186 38 226
rect 46 186 58 226
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 234 86 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 20 123 24 186
rect 16 111 24 123
rect 18 80 24 111
rect 40 111 44 186
rect 40 80 46 111
rect 18 74 26 80
rect 22 54 26 74
rect 32 74 46 80
rect 32 54 36 74
rect 22 10 26 14
rect 32 10 36 14
<< polycontact >>
rect 4 111 16 123
rect 44 111 56 123
<< metal1 >>
rect -6 246 86 248
rect -6 232 86 234
rect 6 226 18 232
rect 46 226 58 232
rect 3 123 17 137
rect 26 117 34 186
rect 43 123 57 137
rect 23 103 37 117
rect 26 68 34 103
rect 26 62 50 68
rect 38 54 50 62
rect 8 8 20 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
<< labels >>
rlabel metal1 23 103 37 117 0 Y
port 2 nsew signal output
rlabel metal1 -6 -8 86 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 86 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal1 43 123 57 137 0 B
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
