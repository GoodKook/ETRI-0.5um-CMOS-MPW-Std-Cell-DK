magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -56 -56 84 354
<< diffusion >>
rect 5 5 23 293
<< metal1 >>
rect 4 4 24 294
<< end >>
