magic
tech scmos
magscale 1 3
timestamp 1723010240
<< checkpaint >>
rect -58 -58 202 182
use pipcap_CDNS_723012252914  pipcap_CDNS_723012252914_0
timestamp 1723012252
transform 1 0 0 0 1 0
box 2 2 142 122
<< end >>
