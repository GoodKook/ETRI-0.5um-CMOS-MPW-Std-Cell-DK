MACRO khu_etri050_stdcells
  CLASS BLOCK ;
  FOREIGN khu_etri050_stdcells ;
  ORIGIN 14.550 8.550 ;
  SIZE 290.700 BY 151.500 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -14.550 130.200 -5.550 142.950 ;
        RECT -14.550 127.800 252.900 130.200 ;
        RECT -14.550 85.200 -5.550 127.800 ;
        RECT 0.900 120.900 2.700 127.800 ;
        RECT 6.900 114.900 8.700 127.800 ;
        RECT 12.900 114.900 14.700 127.800 ;
        RECT 18.900 114.900 20.700 127.800 ;
        RECT 21.900 114.900 23.700 127.800 ;
        RECT 27.900 114.900 29.700 127.800 ;
        RECT 33.900 114.900 35.700 127.800 ;
        RECT 40.200 114.900 42.000 127.800 ;
        RECT 51.000 114.900 52.800 127.800 ;
        RECT 60.900 119.700 62.700 127.800 ;
        RECT 69.900 114.900 71.700 127.800 ;
        RECT 72.900 120.900 74.700 127.800 ;
        RECT 78.900 120.900 80.700 127.800 ;
        RECT 81.900 120.900 83.700 127.800 ;
        RECT 87.900 121.500 89.700 127.800 ;
        RECT 93.900 114.900 95.700 127.800 ;
        RECT 105.900 117.900 107.700 127.800 ;
        RECT 127.200 114.900 129.000 127.800 ;
        RECT 135.300 120.900 137.100 127.800 ;
        RECT 138.900 114.900 140.700 127.800 ;
        RECT 149.400 114.900 151.200 127.800 ;
        RECT 158.400 114.900 160.200 127.800 ;
        RECT 170.400 114.900 172.200 127.800 ;
        RECT 178.200 120.900 180.000 127.800 ;
        RECT 189.000 114.900 190.800 127.800 ;
        RECT 192.600 114.900 194.400 127.800 ;
        RECT 207.600 117.000 209.400 127.800 ;
        RECT 216.900 117.000 218.700 127.800 ;
        RECT 225.600 117.000 227.700 127.800 ;
        RECT 234.900 117.000 236.700 127.800 ;
        RECT 243.900 117.000 245.700 127.800 ;
        RECT -14.550 82.800 262.950 85.200 ;
        RECT -14.550 40.200 -5.550 82.800 ;
        RECT 3.900 75.900 5.700 82.800 ;
        RECT 13.500 75.900 15.300 82.800 ;
        RECT 20.100 75.900 21.900 82.800 ;
        RECT 29.100 78.900 30.900 82.800 ;
        RECT 37.650 75.900 39.450 82.800 ;
        RECT 47.850 75.900 49.650 82.800 ;
        RECT 54.450 75.900 56.250 82.800 ;
        RECT 63.150 78.900 64.950 82.800 ;
        RECT 70.200 75.900 72.000 82.800 ;
        RECT 76.200 75.900 78.000 82.800 ;
        RECT 82.200 77.100 84.000 82.800 ;
        RECT 94.800 75.900 96.600 82.800 ;
        RECT 101.700 75.900 103.500 82.800 ;
        RECT 117.900 75.900 119.700 82.800 ;
        RECT 123.900 75.900 125.700 82.800 ;
        RECT 129.900 75.900 131.700 82.800 ;
        RECT 136.500 75.900 138.300 82.800 ;
        RECT 141.900 72.000 143.700 82.800 ;
        RECT 152.400 69.900 154.200 82.800 ;
        RECT 158.400 72.900 160.200 82.800 ;
        RECT 170.700 75.900 172.500 82.800 ;
        RECT 177.300 75.900 179.100 82.800 ;
        RECT 234.900 76.500 236.700 82.800 ;
        RECT 244.500 75.900 246.300 82.800 ;
        RECT 251.700 75.900 253.500 82.800 ;
        RECT -14.550 37.800 204.600 40.200 ;
        RECT -14.550 -7.050 -5.550 37.800 ;
        RECT 0.900 30.900 2.700 37.800 ;
        RECT 6.900 30.900 8.700 37.800 ;
        RECT 14.700 30.900 16.500 37.800 ;
        RECT 20.700 30.900 22.500 37.800 ;
        RECT 31.500 26.700 33.300 37.800 ;
        RECT 45.300 27.000 47.100 37.800 ;
        RECT 62.100 30.900 63.900 37.800 ;
        RECT 72.900 27.900 74.700 37.800 ;
        RECT 78.900 24.900 80.700 37.800 ;
        RECT 83.700 24.900 85.500 37.800 ;
        RECT 89.700 24.900 91.500 37.800 ;
        RECT 95.700 24.900 97.500 37.800 ;
        RECT 101.700 24.900 103.500 37.800 ;
        RECT 107.700 24.900 109.500 37.800 ;
        RECT 111.600 24.900 113.400 37.800 ;
        RECT 117.600 24.900 119.400 37.800 ;
        RECT 123.600 24.900 125.400 37.800 ;
        RECT 129.600 24.900 131.400 37.800 ;
        RECT 135.600 24.900 137.400 37.800 ;
        RECT 141.600 24.900 143.400 37.800 ;
        RECT 147.600 24.900 149.400 37.800 ;
        RECT 150.600 24.900 152.400 37.800 ;
        RECT 156.600 24.900 158.400 37.800 ;
        RECT 162.600 24.900 164.400 37.800 ;
        RECT 168.600 24.900 170.400 37.800 ;
        RECT 174.600 24.900 176.400 37.800 ;
        RECT 180.600 24.900 182.400 37.800 ;
        RECT 186.600 24.900 188.400 37.800 ;
        RECT 192.600 24.900 194.400 37.800 ;
        RECT 198.600 24.900 200.400 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 91.200 2.700 95.100 ;
        RECT 6.900 91.200 8.700 98.100 ;
        RECT 12.900 91.200 14.700 98.100 ;
        RECT 18.900 91.200 20.700 98.100 ;
        RECT 21.900 91.200 23.700 98.100 ;
        RECT 27.900 91.200 29.700 98.100 ;
        RECT 33.900 91.200 35.700 98.100 ;
        RECT 40.200 91.200 42.000 95.100 ;
        RECT 51.000 91.200 52.800 98.100 ;
        RECT 60.900 91.200 62.700 96.300 ;
        RECT 69.900 91.200 71.700 99.300 ;
        RECT 73.200 91.200 75.000 98.100 ;
        RECT 81.900 91.200 83.700 101.100 ;
        RECT 93.900 91.200 95.700 95.100 ;
        RECT 99.900 91.200 101.700 95.100 ;
        RECT 105.600 91.200 107.700 95.100 ;
        RECT 111.900 91.200 113.700 95.100 ;
        RECT 129.900 91.200 131.700 96.300 ;
        RECT 141.900 91.200 143.700 96.600 ;
        RECT 153.900 91.200 155.700 95.100 ;
        RECT 159.900 91.200 161.700 95.100 ;
        RECT 165.900 92.100 167.700 95.100 ;
        RECT 165.900 91.200 167.100 92.100 ;
        RECT 171.900 91.200 173.700 95.100 ;
        RECT 178.200 91.200 180.000 95.100 ;
        RECT 189.000 91.200 190.800 98.100 ;
        RECT 192.600 91.200 194.400 98.100 ;
        RECT 207.600 91.200 209.400 97.200 ;
        RECT 216.900 91.200 218.700 97.200 ;
        RECT 225.600 91.200 227.400 97.200 ;
        RECT 234.900 91.200 236.700 97.200 ;
        RECT 243.900 91.200 245.700 97.200 ;
        RECT 267.150 91.200 276.150 141.450 ;
        RECT -0.900 88.800 276.150 91.200 ;
        RECT 3.900 46.200 5.700 50.100 ;
        RECT 13.200 46.200 15.000 50.100 ;
        RECT 20.100 46.200 21.900 50.100 ;
        RECT 29.100 46.200 30.900 50.100 ;
        RECT 37.650 46.200 39.450 50.100 ;
        RECT 46.950 46.200 48.750 50.100 ;
        RECT 53.850 46.200 55.650 50.100 ;
        RECT 62.850 46.200 64.650 50.100 ;
        RECT 75.600 46.200 77.400 53.100 ;
        RECT 94.200 46.200 96.000 50.100 ;
        RECT 101.700 46.200 103.500 50.100 ;
        RECT 124.200 46.200 126.000 53.100 ;
        RECT 136.500 46.200 138.300 50.100 ;
        RECT 141.900 46.200 143.700 51.300 ;
        RECT 152.400 46.200 154.200 52.500 ;
        RECT 158.400 46.200 160.200 51.000 ;
        RECT 170.700 47.100 172.500 50.100 ;
        RECT 170.700 46.200 171.900 47.100 ;
        RECT 180.300 46.200 182.100 50.100 ;
        RECT 231.900 46.200 233.700 53.100 ;
        RECT 242.700 46.200 244.500 50.100 ;
        RECT 255.300 46.200 257.100 50.100 ;
        RECT 267.150 46.200 276.150 88.800 ;
        RECT -0.900 43.800 276.150 46.200 ;
        RECT 5.400 1.200 7.200 5.100 ;
        RECT 19.200 1.200 21.000 8.100 ;
        RECT 29.100 1.200 30.900 8.100 ;
        RECT 36.600 1.200 38.400 5.100 ;
        RECT 42.600 1.200 44.400 8.100 ;
        RECT 51.600 1.200 53.400 8.100 ;
        RECT 62.100 1.200 63.900 5.100 ;
        RECT 72.900 1.200 74.700 6.600 ;
        RECT 78.900 1.200 80.700 8.100 ;
        RECT 83.700 1.200 85.500 8.100 ;
        RECT 89.700 1.200 91.500 8.100 ;
        RECT 95.700 1.200 97.500 8.100 ;
        RECT 101.700 1.200 103.500 8.100 ;
        RECT 107.700 1.200 109.500 8.100 ;
        RECT 111.600 1.200 113.400 8.100 ;
        RECT 117.600 1.200 119.400 8.100 ;
        RECT 123.600 1.200 125.400 8.100 ;
        RECT 129.600 1.200 131.400 8.100 ;
        RECT 135.600 1.200 137.400 8.100 ;
        RECT 141.600 1.200 143.400 8.100 ;
        RECT 147.600 1.200 149.400 8.100 ;
        RECT 150.600 1.200 152.400 8.100 ;
        RECT 156.600 1.200 158.400 8.100 ;
        RECT 162.600 1.200 164.400 8.100 ;
        RECT 168.600 1.200 170.400 8.100 ;
        RECT 174.600 1.200 176.400 8.100 ;
        RECT 180.600 1.200 182.400 8.100 ;
        RECT 186.600 1.200 188.400 8.100 ;
        RECT 192.600 1.200 194.400 8.100 ;
        RECT 198.600 1.200 200.400 8.100 ;
        RECT 267.150 1.200 276.150 43.800 ;
        RECT -0.900 -1.200 276.150 1.200 ;
        RECT 267.150 -8.550 276.150 -1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 120.900 5.700 126.900 ;
        RECT 0.600 107.550 2.400 109.350 ;
        RECT 3.900 107.550 5.100 120.900 ;
        RECT 9.900 114.900 11.700 126.900 ;
        RECT 15.900 114.900 17.700 126.900 ;
        RECT 0.450 105.450 2.550 107.550 ;
        RECT 3.450 105.450 5.550 107.550 ;
        RECT 9.900 107.400 11.100 114.900 ;
        RECT 16.200 107.550 17.250 114.900 ;
        RECT 24.900 114.000 26.700 126.900 ;
        RECT 30.900 114.900 32.700 126.900 ;
        RECT 37.200 114.900 39.000 126.900 ;
        RECT 45.300 120.900 47.250 126.900 ;
        RECT 45.450 118.800 47.550 120.900 ;
        RECT 54.000 114.900 55.800 126.900 ;
        RECT 30.900 114.000 32.100 114.900 ;
        RECT 24.900 113.100 32.100 114.000 ;
        RECT 3.900 95.100 5.100 105.450 ;
        RECT 6.450 105.300 8.550 107.400 ;
        RECT 9.450 105.300 11.550 107.400 ;
        RECT 12.450 105.450 14.550 107.550 ;
        RECT 16.200 105.450 20.550 107.550 ;
        RECT 24.600 107.400 26.400 109.200 ;
        RECT 30.900 107.400 32.100 113.100 ;
        RECT 37.200 111.300 38.400 114.900 ;
        RECT 45.450 114.000 47.550 114.900 ;
        RECT 45.450 112.800 53.400 114.000 ;
        RECT 51.600 112.200 53.400 112.800 ;
        RECT 37.200 110.400 45.900 111.300 ;
        RECT 6.600 103.500 8.400 105.300 ;
        RECT 9.900 98.100 11.100 105.300 ;
        RECT 12.600 103.650 14.400 105.450 ;
        RECT 16.200 98.100 17.250 105.450 ;
        RECT 24.450 105.300 26.550 107.400 ;
        RECT 30.450 105.300 32.550 107.400 ;
        RECT 30.900 100.200 32.100 105.300 ;
        RECT 24.900 99.000 32.100 100.200 ;
        RECT 24.900 98.100 26.100 99.000 ;
        RECT 30.900 98.100 32.100 99.000 ;
        RECT 37.200 98.100 38.400 110.400 ;
        RECT 44.100 109.500 45.900 110.400 ;
        RECT 41.100 108.450 42.900 109.350 ;
        RECT 47.700 108.750 50.550 110.850 ;
        RECT 47.700 108.450 48.750 108.750 ;
        RECT 41.100 107.550 48.750 108.450 ;
        RECT 54.600 107.550 55.800 114.900 ;
        RECT 57.900 119.700 59.700 125.700 ;
        RECT 57.900 114.600 58.800 119.700 ;
        RECT 65.400 116.400 67.200 125.700 ;
        RECT 75.900 120.900 77.700 126.900 ;
        RECT 84.900 120.900 86.700 126.900 ;
        RECT 65.400 115.500 67.500 116.400 ;
        RECT 57.900 113.700 65.250 114.600 ;
        RECT 64.050 109.200 65.250 113.700 ;
        RECT 51.450 107.250 55.800 107.550 ;
        RECT 60.600 107.400 62.400 109.200 ;
        RECT 63.750 107.400 65.550 109.200 ;
        RECT 66.600 107.400 67.500 115.500 ;
        RECT 69.600 107.400 71.400 109.200 ;
        RECT 75.900 107.400 77.100 120.900 ;
        RECT 85.200 120.600 86.700 120.900 ;
        RECT 90.900 120.900 92.700 126.900 ;
        RECT 90.900 120.600 91.800 120.900 ;
        RECT 85.200 119.700 91.800 120.600 ;
        RECT 84.600 107.400 86.400 109.200 ;
        RECT 90.900 107.400 91.800 119.700 ;
        RECT 99.000 116.100 100.800 126.900 ;
        RECT 102.900 117.000 104.700 126.900 ;
        RECT 108.900 126.000 116.700 126.900 ;
        RECT 108.900 117.000 110.700 126.000 ;
        RECT 102.900 116.100 110.700 117.000 ;
        RECT 111.900 117.300 113.700 125.100 ;
        RECT 114.900 118.200 116.700 126.000 ;
        RECT 118.500 126.000 126.300 126.900 ;
        RECT 118.500 117.300 120.300 126.000 ;
        RECT 111.900 116.400 120.300 117.300 ;
        RECT 121.500 117.300 123.300 125.100 ;
        RECT 97.200 114.900 100.800 116.100 ;
        RECT 121.500 114.900 122.700 117.300 ;
        RECT 124.500 116.700 126.300 126.000 ;
        RECT 132.300 120.900 134.100 126.900 ;
        RECT 93.600 107.550 95.400 109.350 ;
        RECT 97.200 107.550 98.100 114.900 ;
        RECT 119.250 113.700 122.700 114.900 ;
        RECT 99.600 107.550 101.400 109.350 ;
        RECT 49.650 105.450 55.800 107.250 ;
        RECT 45.900 104.550 47.700 104.850 ;
        RECT 39.450 103.050 47.700 104.550 ;
        RECT 39.450 102.450 41.550 103.050 ;
        RECT 39.300 100.650 41.100 102.450 ;
        RECT 44.550 99.900 45.600 103.050 ;
        RECT 44.550 98.100 46.350 99.900 ;
        RECT 54.600 98.100 55.800 105.450 ;
        RECT 57.450 105.300 59.550 107.400 ;
        RECT 60.450 105.300 62.550 107.400 ;
        RECT 57.600 103.500 59.400 105.300 ;
        RECT 63.900 100.500 65.100 107.400 ;
        RECT 66.450 105.300 68.550 107.400 ;
        RECT 69.450 105.300 71.550 107.400 ;
        RECT 72.450 105.300 74.550 107.400 ;
        RECT 75.450 105.300 77.550 107.400 ;
        RECT 78.450 105.300 80.550 107.400 ;
        RECT 81.450 105.300 83.550 107.400 ;
        RECT 84.450 105.300 86.550 107.400 ;
        RECT 87.450 105.300 89.550 107.400 ;
        RECT 90.450 105.300 92.550 107.400 ;
        RECT 93.450 105.450 95.550 107.550 ;
        RECT 96.450 105.450 98.550 107.550 ;
        RECT 99.450 105.450 101.550 107.550 ;
        RECT 105.600 107.400 107.400 109.200 ;
        RECT 114.600 107.400 116.400 109.200 ;
        RECT 119.250 107.400 120.450 113.700 ;
        RECT 126.600 107.550 128.400 109.350 ;
        RECT 132.450 107.550 133.650 120.900 ;
        RECT 143.400 114.900 146.700 126.900 ;
        RECT 3.900 92.100 5.700 95.100 ;
        RECT 9.900 92.100 11.700 98.100 ;
        RECT 15.900 92.100 17.700 98.100 ;
        RECT 24.900 92.100 26.700 98.100 ;
        RECT 30.900 92.100 32.700 98.100 ;
        RECT 37.200 92.100 39.000 98.100 ;
        RECT 45.450 95.100 47.550 97.200 ;
        RECT 45.300 92.100 47.400 95.100 ;
        RECT 54.000 92.100 55.800 98.100 ;
        RECT 57.900 99.600 65.100 100.500 ;
        RECT 57.900 96.300 58.800 99.600 ;
        RECT 66.600 98.700 67.500 105.300 ;
        RECT 72.600 103.500 74.400 105.300 ;
        RECT 75.900 100.200 77.100 105.300 ;
        RECT 78.600 103.500 80.400 105.300 ;
        RECT 81.600 103.500 83.400 105.300 ;
        RECT 87.600 103.500 89.400 105.300 ;
        RECT 90.900 101.700 91.800 105.300 ;
        RECT 88.500 100.500 91.800 101.700 ;
        RECT 75.900 99.300 80.100 100.200 ;
        RECT 65.400 97.800 67.500 98.700 ;
        RECT 57.900 93.300 59.700 96.300 ;
        RECT 65.400 93.300 67.200 97.800 ;
        RECT 78.300 92.100 80.100 99.300 ;
        RECT 88.500 92.100 90.300 100.500 ;
        RECT 97.200 95.100 98.100 105.450 ;
        RECT 105.450 105.300 107.550 107.400 ;
        RECT 111.450 105.300 113.550 107.400 ;
        RECT 114.450 105.300 116.550 107.400 ;
        RECT 119.250 105.300 122.550 107.400 ;
        RECT 126.450 105.450 128.550 107.550 ;
        RECT 129.450 105.450 131.550 107.550 ;
        RECT 132.450 105.450 134.550 107.550 ;
        RECT 135.450 105.450 137.550 107.550 ;
        RECT 138.600 107.400 140.400 109.200 ;
        RECT 144.600 107.400 145.800 114.900 ;
        RECT 153.900 114.000 155.700 126.900 ;
        RECT 162.000 120.900 163.800 126.900 ;
        RECT 162.300 120.000 164.400 120.900 ;
        RECT 153.900 113.100 162.600 114.000 ;
        RECT 160.650 112.200 162.600 113.100 ;
        RECT 150.600 107.400 152.400 109.200 ;
        RECT 153.600 107.550 155.400 109.350 ;
        RECT 111.600 103.500 113.400 105.300 ;
        RECT 119.250 96.900 120.450 105.300 ;
        RECT 129.600 103.650 131.400 105.450 ;
        RECT 133.350 101.250 134.550 105.450 ;
        RECT 135.600 103.650 137.400 105.450 ;
        RECT 138.450 105.300 140.550 107.400 ;
        RECT 141.450 105.300 143.550 107.400 ;
        RECT 144.450 105.300 146.550 107.400 ;
        RECT 147.450 105.300 149.550 107.400 ;
        RECT 150.450 105.300 152.550 107.400 ;
        RECT 153.450 105.450 155.550 107.550 ;
        RECT 156.450 105.450 158.550 107.550 ;
        RECT 141.600 103.500 143.400 105.300 ;
        RECT 144.450 102.900 145.500 105.300 ;
        RECT 147.600 103.500 149.400 105.300 ;
        RECT 156.600 103.650 158.400 105.450 ;
        RECT 133.350 100.200 137.100 101.250 ;
        RECT 109.650 96.000 120.450 96.900 ;
        RECT 126.900 97.200 134.700 98.550 ;
        RECT 109.650 95.100 110.700 96.000 ;
        RECT 115.650 95.100 116.700 96.000 ;
        RECT 96.900 92.100 98.700 95.100 ;
        RECT 108.900 92.100 110.700 95.100 ;
        RECT 114.900 92.100 116.700 95.100 ;
        RECT 126.900 92.100 128.700 97.200 ;
        RECT 132.900 92.100 134.700 97.200 ;
        RECT 135.900 98.100 137.100 100.200 ;
        RECT 144.600 100.800 145.800 102.900 ;
        RECT 144.600 99.600 149.100 100.800 ;
        RECT 135.900 92.100 137.700 98.100 ;
        RECT 138.900 97.500 146.700 98.400 ;
        RECT 148.200 98.100 149.100 99.600 ;
        RECT 160.650 98.400 161.550 112.200 ;
        RECT 163.500 107.550 164.400 120.000 ;
        RECT 165.900 114.900 167.700 126.900 ;
        RECT 173.400 116.400 175.200 126.900 ;
        RECT 181.200 120.900 183.000 126.900 ;
        RECT 173.400 114.900 175.800 116.400 ;
        RECT 165.900 113.400 167.100 114.900 ;
        RECT 165.900 112.200 173.100 113.400 ;
        RECT 171.300 111.600 173.100 112.200 ;
        RECT 168.600 107.550 170.400 109.350 ;
        RECT 162.450 105.450 164.550 107.550 ;
        RECT 165.450 105.450 167.550 107.550 ;
        RECT 168.450 105.450 170.550 107.550 ;
        RECT 138.900 92.100 140.700 97.500 ;
        RECT 144.900 93.000 146.700 97.500 ;
        RECT 147.900 93.900 149.700 98.100 ;
        RECT 150.900 93.000 152.700 98.100 ;
        RECT 160.650 97.500 162.600 98.400 ;
        RECT 157.200 96.600 162.600 97.500 ;
        RECT 157.200 95.100 158.100 96.600 ;
        RECT 163.500 95.100 164.400 105.450 ;
        RECT 165.600 103.650 167.400 105.450 ;
        RECT 172.200 101.100 173.100 111.600 ;
        RECT 174.450 107.550 175.800 114.900 ;
        RECT 182.100 113.550 183.000 120.900 ;
        RECT 184.500 114.900 186.300 126.900 ;
        RECT 195.600 114.900 197.400 126.900 ;
        RECT 198.600 126.000 206.400 126.900 ;
        RECT 198.600 114.900 200.400 126.000 ;
        RECT 201.600 114.900 203.400 125.100 ;
        RECT 204.600 116.100 206.400 126.000 ;
        RECT 210.600 116.100 212.400 126.900 ;
        RECT 204.600 114.900 212.400 116.100 ;
        RECT 213.900 115.800 215.700 126.900 ;
        RECT 221.400 115.800 223.200 126.900 ;
        RECT 228.900 116.100 230.700 126.900 ;
        RECT 182.100 111.750 183.900 113.550 ;
        RECT 178.200 107.550 180.000 109.200 ;
        RECT 174.450 105.450 176.550 107.550 ;
        RECT 177.900 105.450 180.000 107.550 ;
        RECT 171.300 100.200 173.100 101.100 ;
        RECT 169.800 99.300 173.100 100.200 ;
        RECT 169.800 95.100 170.700 99.300 ;
        RECT 175.500 98.100 176.550 105.450 ;
        RECT 144.900 92.100 152.700 93.000 ;
        RECT 156.900 92.100 158.700 95.100 ;
        RECT 162.900 92.100 164.700 95.100 ;
        RECT 168.900 92.100 170.700 95.100 ;
        RECT 174.900 92.100 176.700 98.100 ;
        RECT 182.100 95.100 183.000 111.750 ;
        RECT 184.950 107.550 186.000 114.900 ;
        RECT 196.500 112.950 197.400 114.900 ;
        RECT 196.500 111.150 198.300 112.950 ;
        RECT 187.800 107.550 189.600 109.200 ;
        RECT 183.900 105.450 186.000 107.550 ;
        RECT 187.500 105.450 189.600 107.550 ;
        RECT 192.900 105.450 195.000 107.550 ;
        RECT 184.950 98.100 186.000 105.450 ;
        RECT 193.500 103.650 195.300 105.450 ;
        RECT 196.500 98.100 197.400 111.150 ;
        RECT 201.600 107.550 202.500 114.900 ;
        RECT 213.900 114.600 218.700 115.800 ;
        RECT 221.400 114.900 224.700 115.800 ;
        RECT 216.600 113.700 218.700 114.600 ;
        RECT 216.600 112.800 221.850 113.700 ;
        RECT 220.050 110.700 221.850 112.800 ;
        RECT 223.500 110.400 224.700 114.900 ;
        RECT 225.600 114.900 230.700 116.100 ;
        RECT 231.900 115.800 233.700 126.900 ;
        RECT 231.900 114.900 236.400 115.800 ;
        RECT 239.400 114.900 241.200 126.900 ;
        RECT 246.900 116.100 248.700 126.900 ;
        RECT 225.600 114.000 227.700 114.900 ;
        RECT 234.300 112.800 236.400 114.900 ;
        RECT 240.000 113.400 241.200 114.900 ;
        RECT 243.900 114.900 248.700 116.100 ;
        RECT 243.900 114.000 246.000 114.900 ;
        RECT 240.000 112.500 241.500 113.400 ;
        RECT 237.450 111.000 239.550 111.300 ;
        RECT 222.750 109.800 224.850 110.400 ;
        RECT 218.700 107.700 220.500 109.500 ;
        RECT 221.850 108.300 224.850 109.800 ;
        RECT 235.800 109.200 239.550 111.000 ;
        RECT 240.600 110.400 241.500 112.500 ;
        RECT 201.600 105.450 203.700 107.550 ;
        RECT 207.600 105.450 209.700 107.550 ;
        RECT 201.600 98.100 202.500 105.450 ;
        RECT 207.900 103.650 209.700 105.450 ;
        RECT 213.450 105.300 215.550 107.400 ;
        RECT 218.700 105.600 220.800 107.700 ;
        RECT 213.750 104.700 215.550 105.300 ;
        RECT 213.750 103.500 220.800 104.700 ;
        RECT 218.700 102.600 220.800 103.500 ;
        RECT 216.150 100.500 218.250 101.100 ;
        RECT 219.150 100.800 220.950 102.600 ;
        RECT 221.850 101.700 222.750 108.300 ;
        RECT 228.600 107.400 230.400 109.200 ;
        RECT 240.450 108.300 242.550 110.400 ;
        RECT 237.000 107.400 238.800 108.000 ;
        RECT 223.800 105.600 225.600 107.400 ;
        RECT 223.650 103.500 225.750 105.600 ;
        RECT 228.450 105.300 230.550 107.400 ;
        RECT 231.450 106.200 238.800 107.400 ;
        RECT 239.700 107.400 242.100 108.300 ;
        RECT 246.600 107.400 248.400 109.200 ;
        RECT 231.450 105.300 233.550 106.200 ;
        RECT 231.750 103.500 233.550 105.300 ;
        RECT 237.000 102.900 238.800 104.700 ;
        RECT 213.900 99.000 218.250 100.500 ;
        RECT 221.850 99.600 224.850 101.700 ;
        RECT 204.600 98.100 211.800 99.000 ;
        RECT 213.900 98.100 215.400 99.000 ;
        RECT 181.200 92.100 183.000 95.100 ;
        RECT 184.500 92.100 186.300 98.100 ;
        RECT 195.600 92.100 197.400 98.100 ;
        RECT 198.600 93.000 200.400 98.100 ;
        RECT 201.600 93.900 203.400 98.100 ;
        RECT 204.600 93.000 206.400 98.100 ;
        RECT 198.600 92.100 206.400 93.000 ;
        RECT 210.600 92.100 212.400 98.100 ;
        RECT 213.900 92.100 215.700 98.100 ;
        RECT 221.850 97.500 222.750 99.600 ;
        RECT 226.200 99.000 228.300 101.400 ;
        RECT 236.700 100.800 238.800 102.900 ;
        RECT 232.500 99.900 238.800 100.800 ;
        RECT 239.700 101.700 240.750 107.400 ;
        RECT 242.100 104.700 243.900 106.500 ;
        RECT 246.450 105.300 248.550 107.400 ;
        RECT 241.650 102.600 243.750 104.700 ;
        RECT 226.200 98.100 230.700 99.000 ;
        RECT 232.500 98.100 233.700 99.900 ;
        RECT 239.700 99.600 242.550 101.700 ;
        RECT 239.700 98.100 240.900 99.600 ;
        RECT 243.900 99.000 246.000 100.200 ;
        RECT 243.900 98.100 248.700 99.000 ;
        RECT 221.100 92.100 222.900 97.500 ;
        RECT 228.900 92.100 230.700 98.100 ;
        RECT 231.900 92.100 233.700 98.100 ;
        RECT 239.400 92.100 241.200 98.100 ;
        RECT 246.900 92.100 248.700 98.100 ;
        RECT 0.900 69.300 2.700 81.900 ;
        RECT 8.700 77.100 10.500 81.900 ;
        RECT 6.900 75.900 10.500 77.100 ;
        RECT 6.900 75.300 8.550 75.900 ;
        RECT 6.450 73.200 8.550 75.300 ;
        RECT 16.500 75.000 18.300 81.900 ;
        RECT 24.600 75.900 26.400 81.900 ;
        RECT 9.600 72.300 11.400 75.000 ;
        RECT 12.600 73.800 19.200 75.000 ;
        RECT 24.300 73.800 26.400 75.900 ;
        RECT 12.600 73.200 14.400 73.800 ;
        RECT 17.400 73.200 19.200 73.800 ;
        RECT 9.450 70.200 11.550 72.300 ;
        RECT 25.200 72.000 27.000 72.600 ;
        RECT 20.100 70.800 27.000 72.000 ;
        RECT 20.100 70.200 21.900 70.800 ;
        RECT 20.100 69.300 21.000 70.200 ;
        RECT 0.900 68.100 21.000 69.300 ;
        RECT 32.100 69.900 33.900 81.900 ;
        RECT 34.650 69.900 36.450 81.900 ;
        RECT 43.050 75.900 44.850 81.900 ;
        RECT 43.050 75.000 44.250 75.900 ;
        RECT 50.850 75.000 52.650 81.900 ;
        RECT 58.650 75.900 60.450 81.900 ;
        RECT 39.450 72.900 44.250 75.000 ;
        RECT 46.950 73.950 53.550 75.000 ;
        RECT 46.950 73.200 48.750 73.950 ;
        RECT 51.750 73.200 53.550 73.950 ;
        RECT 58.650 73.800 62.550 75.900 ;
        RECT 43.050 72.000 44.250 72.900 ;
        RECT 55.950 72.300 57.750 72.900 ;
        RECT 43.050 70.800 50.550 72.000 ;
        RECT 48.750 70.200 50.550 70.800 ;
        RECT 51.450 71.400 57.750 72.300 ;
        RECT 0.900 53.100 1.800 68.100 ;
        RECT 7.800 67.500 9.600 68.100 ;
        RECT 14.400 66.600 16.200 67.200 ;
        RECT 6.450 65.400 16.200 66.600 ;
        RECT 24.300 66.000 26.400 66.600 ;
        RECT 29.400 66.000 31.200 66.600 ;
        RECT 6.450 64.500 8.550 65.400 ;
        RECT 24.300 64.800 31.200 66.000 ;
        RECT 24.300 64.500 26.400 64.800 ;
        RECT 3.600 62.550 5.400 64.350 ;
        RECT 32.100 62.550 33.300 69.900 ;
        RECT 3.450 60.450 5.550 62.550 ;
        RECT 30.450 62.250 33.300 62.550 ;
        RECT 27.000 60.450 33.300 62.250 ;
        RECT 9.450 56.400 11.550 58.200 ;
        RECT 15.450 56.400 17.550 59.550 ;
        RECT 2.850 55.200 23.700 56.400 ;
        RECT 2.850 54.600 4.650 55.200 ;
        RECT 7.800 54.000 9.600 55.200 ;
        RECT 21.900 54.600 23.700 55.200 ;
        RECT 32.100 53.100 33.300 60.450 ;
        RECT 34.650 69.000 35.550 69.900 ;
        RECT 51.450 69.300 52.350 71.400 ;
        RECT 55.950 71.100 57.750 71.400 ;
        RECT 58.650 71.100 61.350 72.900 ;
        RECT 58.650 70.200 59.550 71.100 ;
        RECT 43.950 69.000 52.350 69.300 ;
        RECT 34.650 68.400 52.350 69.000 ;
        RECT 54.450 69.300 59.550 70.200 ;
        RECT 60.450 69.300 62.550 70.200 ;
        RECT 66.150 69.900 67.950 81.900 ;
        RECT 73.200 75.900 75.000 81.900 ;
        RECT 73.200 75.000 74.250 75.900 ;
        RECT 34.650 67.800 45.750 68.400 ;
        RECT 34.650 53.100 35.550 67.800 ;
        RECT 43.950 67.500 45.750 67.800 ;
        RECT 36.450 60.450 38.550 62.550 ;
        RECT 45.450 60.900 47.550 62.550 ;
        RECT 36.600 58.650 38.400 60.450 ;
        RECT 39.600 59.700 47.550 60.900 ;
        RECT 39.600 59.100 41.400 59.700 ;
        RECT 37.500 57.900 38.400 58.650 ;
        RECT 42.600 57.900 44.400 58.500 ;
        RECT 37.500 56.700 44.400 57.900 ;
        RECT 54.450 56.700 55.350 69.300 ;
        RECT 60.450 68.100 64.650 69.300 ;
        RECT 63.750 66.300 65.550 68.100 ;
        RECT 66.750 62.550 67.950 69.900 ;
        RECT 63.450 62.250 67.950 62.550 ;
        RECT 61.650 60.450 67.950 62.250 ;
        RECT 43.350 55.500 55.350 56.700 ;
        RECT 43.350 53.700 44.400 55.500 ;
        RECT 53.550 54.900 55.350 55.500 ;
        RECT 0.900 47.100 2.700 53.100 ;
        RECT 6.450 51.000 8.550 53.100 ;
        RECT 12.600 52.200 14.400 52.800 ;
        RECT 12.600 51.000 17.700 52.200 ;
        RECT 6.900 50.100 8.550 51.000 ;
        RECT 16.500 50.100 17.700 51.000 ;
        RECT 6.900 49.050 10.500 50.100 ;
        RECT 8.700 47.100 10.500 49.050 ;
        RECT 16.500 47.100 18.300 50.100 ;
        RECT 24.300 49.200 26.400 52.200 ;
        RECT 24.600 47.100 26.400 49.200 ;
        RECT 32.100 47.100 33.900 53.100 ;
        RECT 34.650 47.100 36.450 53.100 ;
        RECT 39.450 51.000 41.550 53.100 ;
        RECT 43.050 51.900 44.850 53.700 ;
        RECT 66.750 53.100 67.950 60.450 ;
        RECT 46.350 52.050 48.150 52.800 ;
        RECT 60.450 52.200 62.550 53.100 ;
        RECT 46.350 51.000 51.300 52.050 ;
        RECT 40.500 50.100 41.550 51.000 ;
        RECT 50.250 50.100 51.300 51.000 ;
        RECT 58.800 51.000 62.550 52.200 ;
        RECT 58.800 50.100 59.850 51.000 ;
        RECT 40.500 49.200 44.250 50.100 ;
        RECT 42.450 47.100 44.250 49.200 ;
        RECT 50.250 47.100 52.050 50.100 ;
        RECT 58.050 47.100 59.850 50.100 ;
        RECT 66.150 47.100 67.950 53.100 ;
        RECT 70.200 74.100 74.250 75.000 ;
        RECT 70.200 57.900 71.400 74.100 ;
        RECT 74.700 72.900 76.500 73.200 ;
        RECT 79.200 72.900 81.000 81.900 ;
        RECT 85.500 78.900 87.600 81.900 ;
        RECT 88.500 78.900 90.600 81.900 ;
        RECT 91.650 78.900 93.600 81.900 ;
        RECT 85.500 76.200 86.550 78.900 ;
        RECT 88.500 76.200 89.550 78.900 ;
        RECT 91.650 76.200 92.850 78.900 ;
        RECT 84.450 74.100 86.550 76.200 ;
        RECT 87.450 74.100 89.550 76.200 ;
        RECT 90.450 74.100 92.850 76.200 ;
        RECT 98.700 74.400 100.500 81.900 ;
        RECT 104.700 75.900 106.500 81.900 ;
        RECT 108.300 78.900 110.100 81.900 ;
        RECT 111.300 78.900 113.100 81.900 ;
        RECT 114.300 78.900 116.100 81.900 ;
        RECT 108.300 76.800 110.400 78.900 ;
        RECT 111.300 76.800 113.400 78.900 ;
        RECT 114.450 76.800 116.550 78.900 ;
        RECT 74.700 71.700 93.900 72.900 ;
        RECT 98.700 72.300 101.550 74.400 ;
        RECT 104.700 73.800 107.550 75.900 ;
        RECT 112.350 75.000 113.400 76.800 ;
        RECT 120.900 75.000 122.700 81.900 ;
        RECT 126.900 75.900 128.700 81.900 ;
        RECT 112.350 73.800 120.000 75.000 ;
        RECT 120.900 73.800 126.600 75.000 ;
        RECT 104.700 72.000 107.400 73.800 ;
        RECT 118.200 73.200 120.000 73.800 ;
        RECT 124.800 73.200 126.600 73.800 ;
        RECT 74.700 71.400 76.500 71.700 ;
        RECT 92.700 71.100 93.900 71.700 ;
        RECT 108.450 71.100 110.550 72.000 ;
        RECT 78.000 70.200 79.800 70.800 ;
        RECT 87.450 70.200 89.550 70.800 ;
        RECT 78.000 69.000 89.550 70.200 ;
        RECT 92.700 69.900 110.550 71.100 ;
        RECT 114.450 70.800 116.550 72.000 ;
        RECT 127.500 70.800 128.700 75.900 ;
        RECT 133.500 75.900 135.300 81.900 ;
        RECT 114.450 69.900 131.400 70.800 ;
        RECT 87.450 68.700 89.550 69.000 ;
        RECT 92.700 67.800 129.600 69.000 ;
        RECT 92.700 67.200 93.900 67.800 ;
        RECT 127.800 67.200 129.600 67.800 ;
        RECT 80.550 66.300 93.900 67.200 ;
        RECT 80.550 65.400 82.350 66.300 ;
        RECT 72.450 63.300 74.550 65.400 ;
        RECT 78.450 63.600 82.350 65.400 ;
        RECT 99.450 64.800 101.550 66.900 ;
        RECT 105.450 66.600 107.550 66.900 ;
        RECT 103.650 64.800 107.550 66.600 ;
        RECT 112.200 64.800 114.000 66.600 ;
        RECT 78.450 63.300 80.550 63.600 ;
        RECT 83.250 63.300 90.000 64.350 ;
        RECT 72.600 61.800 74.400 63.300 ;
        RECT 83.250 61.800 84.450 63.300 ;
        RECT 72.600 60.600 84.450 61.800 ;
        RECT 86.250 60.600 88.050 62.400 ;
        RECT 88.950 61.800 90.000 63.300 ;
        RECT 90.900 63.600 101.550 64.800 ;
        RECT 113.100 63.600 114.000 64.800 ;
        RECT 90.900 63.000 92.700 63.600 ;
        RECT 99.450 62.700 114.000 63.600 ;
        RECT 117.300 63.300 122.400 65.100 ;
        RECT 125.100 63.300 128.550 65.400 ;
        RECT 117.300 61.800 118.200 63.300 ;
        RECT 88.950 60.600 118.200 61.800 ;
        RECT 125.100 60.600 126.300 63.300 ;
        RECT 70.200 56.700 85.500 57.900 ;
        RECT 70.200 53.100 71.400 56.700 ;
        RECT 74.400 55.200 76.200 55.800 ;
        RECT 74.400 54.000 82.800 55.200 ;
        RECT 81.300 53.100 82.800 54.000 ;
        RECT 70.200 47.100 72.000 53.100 ;
        RECT 81.000 47.100 82.800 53.100 ;
        RECT 84.450 53.100 85.500 56.700 ;
        RECT 87.000 55.500 88.050 60.600 ;
        RECT 119.400 59.400 126.300 60.600 ;
        RECT 96.300 58.500 98.400 59.400 ;
        RECT 119.400 59.100 120.900 59.400 ;
        RECT 93.300 57.300 98.400 58.500 ;
        RECT 102.600 57.600 120.900 59.100 ;
        RECT 123.000 58.200 124.800 58.500 ;
        RECT 127.800 58.200 129.600 58.500 ;
        RECT 90.300 55.500 92.100 57.300 ;
        RECT 93.300 56.700 95.100 57.300 ;
        RECT 87.000 54.300 96.900 55.500 ;
        RECT 102.600 55.200 104.400 57.600 ;
        RECT 121.800 56.700 129.600 58.200 ;
        RECT 110.400 54.900 117.000 56.700 ;
        RECT 96.000 53.100 96.900 54.300 ;
        RECT 121.800 53.100 123.300 56.700 ;
        RECT 130.500 53.100 131.400 69.900 ;
        RECT 84.450 51.000 86.550 53.100 ;
        RECT 87.450 51.000 89.550 53.100 ;
        RECT 90.450 51.000 92.550 53.100 ;
        RECT 96.000 51.300 97.800 53.100 ;
        RECT 85.200 50.100 86.550 51.000 ;
        RECT 88.200 50.100 89.550 51.000 ;
        RECT 91.200 50.100 92.550 51.000 ;
        RECT 99.450 51.000 101.550 53.100 ;
        RECT 105.450 51.000 107.550 53.100 ;
        RECT 108.450 51.000 110.550 53.100 ;
        RECT 111.450 51.000 113.550 53.100 ;
        RECT 114.450 51.000 116.550 53.100 ;
        RECT 119.100 51.900 123.300 53.100 ;
        RECT 99.450 50.100 100.500 51.000 ;
        RECT 105.450 50.100 106.500 51.000 ;
        RECT 108.450 50.100 110.100 51.000 ;
        RECT 111.450 50.100 113.100 51.000 ;
        RECT 114.450 50.100 116.100 51.000 ;
        RECT 85.200 47.100 87.000 50.100 ;
        RECT 88.200 47.100 90.000 50.100 ;
        RECT 91.200 47.100 93.000 50.100 ;
        RECT 98.700 47.100 100.500 50.100 ;
        RECT 104.700 47.100 106.500 50.100 ;
        RECT 108.300 47.100 110.100 50.100 ;
        RECT 111.300 47.100 113.100 50.100 ;
        RECT 114.300 47.100 116.100 50.100 ;
        RECT 119.100 47.100 120.900 51.900 ;
        RECT 129.600 47.100 131.400 53.100 ;
        RECT 133.500 65.400 135.000 75.900 ;
        RECT 138.900 70.800 140.700 81.900 ;
        RECT 144.900 72.000 146.700 81.900 ;
        RECT 144.900 70.800 146.250 72.000 ;
        RECT 147.900 71.100 149.700 81.900 ;
        RECT 155.400 72.000 157.200 81.900 ;
        RECT 161.400 72.000 163.200 81.900 ;
        RECT 155.400 71.100 163.200 72.000 ;
        RECT 138.900 69.900 146.250 70.800 ;
        RECT 147.450 69.000 149.550 71.100 ;
        RECT 164.400 69.000 166.350 81.900 ;
        RECT 173.700 77.250 175.500 81.900 ;
        RECT 159.450 66.900 161.550 69.000 ;
        RECT 162.450 66.900 166.350 69.000 ;
        RECT 173.400 75.900 175.500 77.250 ;
        RECT 180.300 75.900 182.100 81.900 ;
        RECT 231.900 75.900 233.700 81.900 ;
        RECT 173.400 68.400 174.300 75.900 ;
        RECT 175.500 71.400 177.600 71.550 ;
        RECT 175.500 69.600 179.400 71.400 ;
        RECT 175.500 69.450 177.600 69.600 ;
        RECT 180.300 68.400 181.500 75.900 ;
        RECT 232.200 75.600 233.700 75.900 ;
        RECT 237.900 75.900 239.700 81.900 ;
        RECT 241.500 75.900 243.300 81.900 ;
        RECT 237.900 75.600 239.100 75.900 ;
        RECT 232.200 74.700 239.100 75.600 ;
        RECT 173.400 67.500 176.250 68.400 ;
        RECT 159.900 66.300 161.550 66.900 ;
        RECT 133.500 63.300 137.550 65.400 ;
        RECT 159.900 64.500 161.700 66.300 ;
        RECT 165.450 66.150 166.350 66.900 ;
        RECT 165.450 65.250 174.300 66.150 ;
        RECT 172.500 64.350 174.300 65.250 ;
        RECT 133.500 50.100 135.000 63.300 ;
        RECT 141.000 62.550 142.800 64.350 ;
        RECT 157.800 62.700 159.600 63.300 ;
        RECT 163.800 62.700 165.600 63.450 ;
        RECT 157.800 62.550 165.600 62.700 ;
        RECT 141.450 60.450 143.550 62.550 ;
        RECT 144.450 61.500 165.600 62.550 ;
        RECT 166.800 62.550 168.600 63.450 ;
        RECT 175.350 62.550 176.250 67.500 ;
        RECT 177.450 67.200 181.500 68.400 ;
        RECT 177.450 62.550 178.650 67.200 ;
        RECT 238.050 62.850 239.100 74.700 ;
        RECT 144.450 60.750 148.350 61.500 ;
        RECT 144.450 60.450 146.550 60.750 ;
        RECT 166.800 60.600 170.550 62.550 ;
        RECT 141.600 56.700 143.100 60.450 ;
        RECT 155.400 59.550 170.550 60.600 ;
        RECT 174.450 60.450 176.550 62.550 ;
        RECT 177.450 60.450 179.550 62.550 ;
        RECT 231.450 62.400 233.550 62.550 ;
        RECT 231.450 60.450 235.350 62.400 ;
        RECT 237.450 60.750 239.550 62.850 ;
        RECT 241.500 62.550 242.550 75.900 ;
        RECT 247.500 69.900 249.300 81.900 ;
        RECT 254.700 75.900 256.500 81.900 ;
        RECT 247.650 67.950 248.550 69.900 ;
        RECT 247.650 67.050 250.950 67.950 ;
        RECT 240.450 60.450 242.550 62.550 ;
        RECT 246.450 60.450 248.550 62.550 ;
        RECT 144.000 58.650 145.800 59.550 ;
        RECT 149.400 58.650 151.200 59.550 ;
        RECT 155.400 58.650 157.200 59.550 ;
        RECT 144.000 57.600 157.200 58.650 ;
        RECT 160.050 56.700 167.700 57.600 ;
        RECT 141.600 55.800 161.250 56.700 ;
        RECT 166.500 55.800 171.900 56.700 ;
        RECT 152.400 54.900 154.200 55.800 ;
        RECT 138.900 52.200 146.100 53.100 ;
        RECT 147.450 52.800 149.550 54.900 ;
        RECT 162.450 53.700 165.450 55.800 ;
        RECT 170.100 54.750 171.900 55.800 ;
        RECT 133.500 47.100 135.300 50.100 ;
        RECT 138.900 47.100 140.700 52.200 ;
        RECT 144.900 47.100 146.700 52.200 ;
        RECT 147.900 51.900 149.550 52.800 ;
        RECT 155.400 51.900 163.200 52.800 ;
        RECT 147.900 47.100 149.700 51.900 ;
        RECT 155.400 47.100 157.200 51.900 ;
        RECT 161.400 47.100 163.200 51.900 ;
        RECT 164.400 51.600 165.450 53.700 ;
        RECT 175.350 52.200 176.250 60.450 ;
        RECT 164.400 47.100 166.350 51.600 ;
        RECT 174.000 51.000 176.250 52.200 ;
        RECT 174.000 50.100 174.900 51.000 ;
        RECT 177.450 50.100 178.500 60.450 ;
        RECT 233.850 57.150 235.200 60.450 ;
        RECT 237.000 59.550 238.800 59.850 ;
        RECT 246.600 59.550 248.400 60.450 ;
        RECT 237.000 58.650 248.400 59.550 ;
        RECT 249.600 59.250 250.950 67.050 ;
        RECT 254.700 62.550 255.600 75.900 ;
        RECT 252.450 60.450 255.600 62.550 ;
        RECT 237.000 58.050 238.800 58.650 ;
        RECT 249.600 58.350 253.200 59.250 ;
        RECT 249.600 57.150 251.400 57.450 ;
        RECT 233.850 56.100 251.400 57.150 ;
        RECT 249.600 55.650 251.400 56.100 ;
        RECT 252.300 55.650 253.200 58.350 ;
        RECT 254.700 57.450 255.600 60.450 ;
        RECT 254.700 56.550 259.200 57.450 ;
        RECT 236.100 54.900 239.550 55.200 ;
        RECT 236.100 53.100 242.550 54.900 ;
        RECT 252.300 54.750 254.400 55.650 ;
        RECT 248.850 53.850 254.400 54.750 ;
        RECT 248.850 53.100 250.650 53.850 ;
        RECT 173.700 47.100 175.500 50.100 ;
        RECT 177.300 47.100 179.100 50.100 ;
        RECT 236.100 47.100 237.900 53.100 ;
        RECT 239.700 49.950 241.800 52.200 ;
        RECT 239.700 47.100 241.500 49.950 ;
        RECT 245.700 48.000 247.500 53.100 ;
        RECT 248.700 48.900 250.500 53.100 ;
        RECT 251.700 48.000 253.500 52.500 ;
        RECT 245.700 47.100 253.500 48.000 ;
        RECT 258.300 50.100 259.200 56.550 ;
        RECT 258.300 47.100 260.100 50.100 ;
        RECT 3.900 30.900 5.700 36.900 ;
        RECT 9.900 30.900 11.700 36.900 ;
        RECT 17.700 30.900 19.500 36.900 ;
        RECT 0.450 15.450 2.550 17.550 ;
        RECT 0.600 13.650 2.400 15.450 ;
        RECT 4.050 10.800 5.100 30.900 ;
        RECT 6.600 17.550 8.400 19.350 ;
        RECT 9.900 17.550 11.100 30.900 ;
        RECT 6.450 15.450 8.550 17.550 ;
        RECT 9.450 15.450 11.550 17.550 ;
        RECT 0.900 9.600 8.400 10.800 ;
        RECT 0.900 2.100 2.700 9.600 ;
        RECT 6.600 9.000 8.400 9.600 ;
        RECT 9.450 5.850 10.500 15.450 ;
        RECT 14.250 15.300 16.350 17.400 ;
        RECT 14.400 13.500 16.200 15.300 ;
        RECT 17.700 10.800 18.600 30.900 ;
        RECT 23.700 24.900 25.500 36.900 ;
        RECT 28.500 25.800 30.300 36.900 ;
        RECT 34.500 25.800 36.300 36.900 ;
        RECT 28.500 24.900 36.300 25.800 ;
        RECT 37.500 24.900 39.300 36.900 ;
        RECT 42.300 26.100 44.100 36.900 ;
        RECT 48.300 36.000 56.100 36.900 ;
        RECT 48.300 26.100 50.100 36.000 ;
        RECT 42.300 25.200 50.100 26.100 ;
        RECT 20.400 17.400 22.200 19.200 ;
        RECT 24.000 17.400 24.900 24.900 ;
        RECT 31.200 17.400 33.000 19.200 ;
        RECT 37.800 17.400 38.700 24.900 ;
        RECT 51.300 24.000 53.100 35.100 ;
        RECT 54.300 24.900 56.100 36.000 ;
        RECT 59.100 30.900 60.900 36.900 ;
        RECT 48.000 23.100 53.100 24.000 ;
        RECT 59.100 24.000 60.300 30.900 ;
        RECT 65.100 24.900 66.900 36.900 ;
        RECT 59.100 23.100 64.800 24.000 ;
        RECT 45.000 17.400 46.800 19.200 ;
        RECT 48.000 17.400 48.900 23.100 ;
        RECT 62.850 22.200 64.800 23.100 ;
        RECT 51.000 17.400 52.800 19.200 ;
        RECT 58.800 17.550 60.600 19.350 ;
        RECT 20.250 15.300 22.350 17.400 ;
        RECT 23.250 15.300 25.350 17.400 ;
        RECT 28.050 15.300 30.150 17.400 ;
        RECT 31.050 15.300 33.150 17.400 ;
        RECT 34.050 15.300 36.150 17.400 ;
        RECT 37.050 15.300 39.150 17.400 ;
        RECT 41.850 15.300 43.950 17.400 ;
        RECT 44.850 15.300 46.950 17.400 ;
        RECT 47.850 15.300 49.950 17.400 ;
        RECT 50.850 15.300 52.950 17.400 ;
        RECT 53.850 15.300 55.950 17.400 ;
        RECT 58.650 15.450 60.750 17.550 ;
        RECT 8.400 5.100 10.500 5.850 ;
        RECT 14.700 9.900 22.200 10.800 ;
        RECT 8.400 2.100 10.200 5.100 ;
        RECT 14.700 2.100 16.500 9.900 ;
        RECT 20.400 9.000 22.200 9.900 ;
        RECT 24.000 8.100 24.900 15.300 ;
        RECT 28.200 13.500 30.000 15.300 ;
        RECT 34.200 13.500 36.000 15.300 ;
        RECT 37.800 8.100 38.700 15.300 ;
        RECT 42.000 13.500 43.800 15.300 ;
        RECT 47.850 8.100 48.900 15.300 ;
        RECT 54.000 13.500 55.800 15.300 ;
        RECT 62.850 10.800 63.750 22.200 ;
        RECT 65.700 17.550 66.900 24.900 ;
        RECT 69.900 27.900 71.700 36.900 ;
        RECT 69.900 24.300 71.100 27.900 ;
        RECT 75.900 25.200 77.700 36.900 ;
        RECT 69.900 23.400 75.750 24.300 ;
        RECT 73.950 22.500 75.750 23.400 ;
        RECT 69.600 17.550 71.400 19.350 ;
        RECT 64.650 15.450 66.900 17.550 ;
        RECT 69.450 15.450 71.550 17.550 ;
        RECT 62.850 9.900 64.800 10.800 ;
        RECT 22.200 6.300 24.900 8.100 ;
        RECT 33.600 6.900 38.700 8.100 ;
        RECT 22.200 2.100 24.000 6.300 ;
        RECT 33.600 2.100 35.400 6.900 ;
        RECT 47.100 2.100 48.900 8.100 ;
        RECT 59.100 9.000 64.800 9.900 ;
        RECT 59.100 5.100 60.300 9.000 ;
        RECT 65.700 8.100 66.900 15.450 ;
        RECT 73.950 10.800 75.150 22.500 ;
        RECT 76.650 17.550 77.700 25.200 ;
        RECT 86.700 24.000 88.500 36.900 ;
        RECT 92.700 24.000 94.500 36.900 ;
        RECT 98.700 24.000 100.500 36.900 ;
        RECT 104.700 24.000 106.500 36.900 ;
        RECT 114.600 24.000 116.400 36.900 ;
        RECT 120.600 24.000 122.400 36.900 ;
        RECT 126.600 24.000 128.400 36.900 ;
        RECT 132.600 24.000 134.400 36.900 ;
        RECT 138.600 24.000 140.400 36.900 ;
        RECT 144.600 24.000 146.400 36.900 ;
        RECT 153.600 24.000 155.400 36.900 ;
        RECT 159.600 24.000 161.400 36.900 ;
        RECT 165.600 24.000 167.400 36.900 ;
        RECT 171.600 24.000 173.400 36.900 ;
        RECT 177.600 24.000 179.400 36.900 ;
        RECT 183.600 24.000 185.400 36.900 ;
        RECT 189.600 24.000 191.400 36.900 ;
        RECT 195.600 24.000 197.400 36.900 ;
        RECT 86.700 22.800 90.600 24.000 ;
        RECT 92.700 22.800 96.600 24.000 ;
        RECT 98.700 22.800 102.600 24.000 ;
        RECT 104.700 22.800 107.400 24.000 ;
        RECT 114.600 22.800 118.650 24.000 ;
        RECT 120.600 22.800 124.500 24.000 ;
        RECT 126.600 22.800 130.500 24.000 ;
        RECT 132.600 22.800 136.800 24.000 ;
        RECT 138.600 22.800 141.900 24.000 ;
        RECT 144.600 22.800 147.900 24.000 ;
        RECT 153.600 22.800 157.500 24.000 ;
        RECT 159.600 22.800 163.500 24.000 ;
        RECT 165.600 22.800 169.500 24.000 ;
        RECT 171.600 22.800 175.800 24.000 ;
        RECT 177.600 22.800 180.900 24.000 ;
        RECT 183.600 22.800 187.500 24.000 ;
        RECT 189.600 22.800 192.600 24.000 ;
        RECT 195.600 22.800 198.750 24.000 ;
        RECT 76.650 15.450 80.550 17.550 ;
        RECT 73.950 9.900 75.750 10.800 ;
        RECT 59.100 2.100 60.900 5.100 ;
        RECT 65.100 2.100 66.900 8.100 ;
        RECT 69.900 9.000 75.750 9.900 ;
        RECT 69.900 6.600 71.100 9.000 ;
        RECT 76.650 8.100 77.700 15.450 ;
        RECT 86.250 15.300 88.350 17.400 ;
        RECT 86.400 13.500 88.200 15.300 ;
        RECT 89.400 12.300 90.600 22.800 ;
        RECT 91.800 12.300 93.600 12.900 ;
        RECT 89.400 11.100 93.600 12.300 ;
        RECT 95.400 12.300 96.600 22.800 ;
        RECT 97.800 12.300 99.600 12.900 ;
        RECT 95.400 11.100 99.600 12.300 ;
        RECT 101.400 12.300 102.600 22.800 ;
        RECT 106.500 17.400 107.400 22.800 ;
        RECT 106.500 15.300 109.350 17.400 ;
        RECT 114.150 15.450 116.250 17.550 ;
        RECT 103.800 12.300 105.600 12.900 ;
        RECT 101.400 11.100 105.600 12.300 ;
        RECT 89.400 10.200 90.600 11.100 ;
        RECT 95.400 10.200 96.600 11.100 ;
        RECT 101.400 10.200 102.600 11.100 ;
        RECT 106.500 10.200 107.400 15.300 ;
        RECT 114.300 13.650 116.100 15.450 ;
        RECT 117.450 12.300 118.650 22.800 ;
        RECT 119.700 12.300 121.500 12.900 ;
        RECT 117.450 11.100 121.500 12.300 ;
        RECT 123.300 12.300 124.500 22.800 ;
        RECT 125.700 12.300 127.500 12.900 ;
        RECT 123.300 11.100 127.500 12.300 ;
        RECT 129.300 12.300 130.500 22.800 ;
        RECT 131.700 12.300 133.500 12.900 ;
        RECT 129.300 11.100 133.500 12.300 ;
        RECT 135.600 12.300 136.800 22.800 ;
        RECT 137.700 12.300 139.500 12.900 ;
        RECT 135.600 11.100 139.500 12.300 ;
        RECT 140.700 12.300 141.900 22.800 ;
        RECT 146.700 17.550 147.900 22.800 ;
        RECT 146.700 15.450 149.250 17.550 ;
        RECT 153.150 15.450 155.250 17.550 ;
        RECT 143.700 12.300 145.500 12.900 ;
        RECT 140.700 11.100 145.500 12.300 ;
        RECT 117.450 10.200 118.650 11.100 ;
        RECT 123.300 10.200 124.500 11.100 ;
        RECT 129.300 10.200 130.500 11.100 ;
        RECT 135.600 10.200 136.800 11.100 ;
        RECT 140.700 10.200 141.900 11.100 ;
        RECT 146.700 10.200 147.900 15.450 ;
        RECT 153.300 13.650 155.100 15.450 ;
        RECT 156.450 12.300 157.500 22.800 ;
        RECT 158.700 12.300 160.500 12.900 ;
        RECT 156.450 11.100 160.500 12.300 ;
        RECT 162.300 12.300 163.500 22.800 ;
        RECT 164.700 12.300 166.500 12.900 ;
        RECT 162.300 11.100 166.500 12.300 ;
        RECT 168.300 12.300 169.500 22.800 ;
        RECT 170.700 12.300 172.500 12.900 ;
        RECT 168.300 11.100 172.500 12.300 ;
        RECT 174.600 12.300 175.800 22.800 ;
        RECT 176.700 12.300 178.500 12.900 ;
        RECT 174.600 11.100 178.500 12.300 ;
        RECT 179.700 12.300 180.900 22.800 ;
        RECT 182.700 12.300 184.500 12.900 ;
        RECT 179.700 11.100 184.500 12.300 ;
        RECT 186.300 12.300 187.500 22.800 ;
        RECT 188.700 12.300 190.500 12.900 ;
        RECT 186.300 11.100 190.500 12.300 ;
        RECT 191.400 12.300 192.600 22.800 ;
        RECT 197.550 17.550 198.750 22.800 ;
        RECT 197.550 15.450 200.250 17.550 ;
        RECT 194.700 12.300 196.500 12.900 ;
        RECT 191.400 11.100 196.500 12.300 ;
        RECT 156.450 10.200 157.500 11.100 ;
        RECT 162.300 10.200 163.500 11.100 ;
        RECT 168.300 10.200 169.500 11.100 ;
        RECT 174.600 10.200 175.800 11.100 ;
        RECT 179.700 10.200 180.900 11.100 ;
        RECT 186.300 10.200 187.500 11.100 ;
        RECT 191.400 10.200 192.600 11.100 ;
        RECT 197.550 10.200 198.750 15.450 ;
        RECT 69.900 2.100 71.700 6.600 ;
        RECT 75.900 2.100 77.700 8.100 ;
        RECT 86.700 9.000 90.600 10.200 ;
        RECT 92.700 9.000 96.600 10.200 ;
        RECT 98.700 9.000 102.600 10.200 ;
        RECT 104.700 9.000 107.400 10.200 ;
        RECT 114.600 9.000 118.650 10.200 ;
        RECT 120.600 9.000 124.500 10.200 ;
        RECT 126.600 9.000 130.500 10.200 ;
        RECT 132.600 9.000 136.800 10.200 ;
        RECT 138.600 9.000 141.900 10.200 ;
        RECT 144.600 9.000 147.900 10.200 ;
        RECT 153.600 9.000 157.500 10.200 ;
        RECT 159.600 9.000 163.500 10.200 ;
        RECT 165.600 9.000 169.500 10.200 ;
        RECT 171.600 9.000 175.800 10.200 ;
        RECT 177.600 9.000 180.900 10.200 ;
        RECT 183.600 9.000 187.500 10.200 ;
        RECT 189.600 9.000 192.600 10.200 ;
        RECT 195.600 9.000 198.750 10.200 ;
        RECT 86.700 2.100 88.500 9.000 ;
        RECT 92.700 2.100 94.500 9.000 ;
        RECT 98.700 2.100 100.500 9.000 ;
        RECT 104.700 2.100 106.500 9.000 ;
        RECT 114.600 2.100 116.400 9.000 ;
        RECT 120.600 2.100 122.400 9.000 ;
        RECT 126.600 2.100 128.400 9.000 ;
        RECT 132.600 2.100 134.400 9.000 ;
        RECT 138.600 2.100 140.400 9.000 ;
        RECT 144.600 2.100 146.400 9.000 ;
        RECT 153.600 2.100 155.400 9.000 ;
        RECT 159.600 2.100 161.400 9.000 ;
        RECT 165.600 2.100 167.400 9.000 ;
        RECT 171.600 2.100 173.400 9.000 ;
        RECT 177.600 2.100 179.400 9.000 ;
        RECT 183.600 2.100 185.400 9.000 ;
        RECT 189.600 2.100 191.400 9.000 ;
        RECT 195.600 2.100 197.400 9.000 ;
      LAYER metal2 ;
        RECT 45.450 118.800 47.550 120.900 ;
        RECT 45.600 114.900 46.800 118.800 ;
        RECT 45.450 112.800 47.550 114.900 ;
        RECT 216.600 113.700 218.700 115.800 ;
        RECT 225.600 114.000 227.700 116.100 ;
        RECT 3.900 107.550 5.100 110.100 ;
        RECT 0.450 105.450 2.550 107.550 ;
        RECT 3.450 105.450 5.550 107.550 ;
        RECT 6.900 107.400 8.100 110.100 ;
        RECT 12.900 107.550 14.100 110.100 ;
        RECT 0.900 102.900 2.100 105.450 ;
        RECT 6.450 105.300 8.550 107.400 ;
        RECT 9.450 105.300 11.550 107.400 ;
        RECT 12.450 105.450 14.550 107.550 ;
        RECT 18.450 105.450 20.550 107.550 ;
        RECT 30.900 107.400 32.100 110.100 ;
        RECT 9.900 102.900 11.100 105.300 ;
        RECT 18.900 102.900 20.100 105.450 ;
        RECT 24.450 105.300 26.550 107.400 ;
        RECT 30.450 105.300 32.550 107.400 ;
        RECT 24.900 102.900 26.100 105.300 ;
        RECT 39.900 104.550 41.100 107.100 ;
        RECT 39.450 102.450 41.550 104.550 ;
        RECT 45.600 97.200 46.800 112.800 ;
        RECT 48.900 110.850 50.100 113.100 ;
        RECT 48.450 108.750 50.550 110.850 ;
        RECT 51.450 105.450 53.550 107.550 ;
        RECT 57.900 107.400 59.100 110.100 ;
        RECT 66.900 107.400 68.100 110.100 ;
        RECT 72.900 107.400 74.100 110.100 ;
        RECT 78.900 107.400 80.100 110.100 ;
        RECT 81.900 107.400 83.100 110.100 ;
        RECT 87.900 107.400 89.100 110.100 ;
        RECT 96.900 107.550 98.100 110.100 ;
        RECT 51.900 102.900 53.100 105.450 ;
        RECT 57.450 105.300 59.550 107.400 ;
        RECT 60.450 105.300 62.550 107.400 ;
        RECT 66.450 105.300 68.550 107.400 ;
        RECT 69.450 105.300 71.550 107.400 ;
        RECT 72.450 105.300 74.550 107.400 ;
        RECT 75.450 105.300 77.550 107.400 ;
        RECT 78.450 105.300 80.550 107.400 ;
        RECT 81.450 105.300 83.550 107.400 ;
        RECT 84.450 105.300 86.550 107.400 ;
        RECT 87.450 105.300 89.550 107.400 ;
        RECT 90.450 105.300 92.550 107.400 ;
        RECT 93.450 105.450 95.550 107.550 ;
        RECT 96.450 105.450 98.550 107.550 ;
        RECT 99.450 105.450 101.550 107.550 ;
        RECT 111.900 107.400 113.100 110.100 ;
        RECT 120.900 107.400 122.100 110.100 ;
        RECT 129.900 107.550 131.100 110.100 ;
        RECT 135.900 107.550 137.100 110.100 ;
        RECT 60.900 102.900 62.100 105.300 ;
        RECT 69.900 102.900 71.100 105.300 ;
        RECT 75.900 102.900 77.100 105.300 ;
        RECT 84.900 102.900 86.100 105.300 ;
        RECT 90.900 102.900 92.100 105.300 ;
        RECT 93.900 102.900 95.100 105.450 ;
        RECT 99.900 102.900 101.100 105.450 ;
        RECT 105.450 105.300 107.550 107.400 ;
        RECT 111.450 105.300 113.550 107.400 ;
        RECT 114.450 105.300 116.550 107.400 ;
        RECT 120.450 105.300 122.550 107.400 ;
        RECT 126.450 105.450 128.550 107.550 ;
        RECT 129.450 105.450 131.550 107.550 ;
        RECT 132.450 105.450 134.550 107.550 ;
        RECT 135.450 105.450 137.550 107.550 ;
        RECT 141.900 107.400 143.100 110.100 ;
        RECT 147.900 107.400 149.100 110.100 ;
        RECT 156.900 107.550 158.100 110.100 ;
        RECT 165.900 107.550 167.100 110.100 ;
        RECT 174.900 107.550 176.100 110.100 ;
        RECT 177.900 107.550 179.100 110.100 ;
        RECT 183.900 107.550 185.100 110.100 ;
        RECT 188.400 107.550 189.600 110.100 ;
        RECT 105.900 102.900 107.100 105.300 ;
        RECT 114.900 102.900 116.100 105.300 ;
        RECT 126.900 102.900 128.100 105.450 ;
        RECT 132.900 102.900 134.100 105.450 ;
        RECT 138.450 105.300 140.550 107.400 ;
        RECT 141.450 105.300 143.550 107.400 ;
        RECT 144.450 105.300 146.550 107.400 ;
        RECT 147.450 105.300 149.550 107.400 ;
        RECT 150.450 105.300 152.550 107.400 ;
        RECT 153.450 105.450 155.550 107.550 ;
        RECT 156.450 105.450 158.550 107.550 ;
        RECT 162.450 105.450 164.550 107.550 ;
        RECT 165.450 105.450 167.550 107.550 ;
        RECT 168.450 105.450 170.550 107.550 ;
        RECT 174.450 105.450 176.550 107.550 ;
        RECT 177.900 105.450 180.000 107.550 ;
        RECT 183.900 105.450 186.000 107.550 ;
        RECT 187.500 105.450 189.600 107.550 ;
        RECT 192.900 107.550 194.100 110.100 ;
        RECT 201.900 107.550 203.100 110.100 ;
        RECT 207.900 107.550 209.100 110.100 ;
        RECT 192.900 105.450 195.000 107.550 ;
        RECT 201.600 105.450 203.700 107.550 ;
        RECT 207.600 105.450 209.700 107.550 ;
        RECT 213.900 107.400 215.100 110.100 ;
        RECT 138.900 102.900 140.100 105.300 ;
        RECT 144.900 102.900 146.100 105.300 ;
        RECT 150.900 102.900 152.100 105.300 ;
        RECT 153.900 102.900 155.100 105.450 ;
        RECT 162.900 102.900 164.100 105.450 ;
        RECT 168.900 102.900 170.100 105.450 ;
        RECT 213.450 105.300 215.550 107.400 ;
        RECT 216.900 101.100 217.800 113.700 ;
        RECT 222.900 110.400 224.100 113.100 ;
        RECT 222.750 108.300 224.850 110.400 ;
        RECT 218.700 107.400 220.800 107.700 ;
        RECT 226.650 107.400 227.550 114.000 ;
        RECT 234.300 112.800 236.400 114.900 ;
        RECT 243.900 114.000 246.000 116.100 ;
        RECT 231.900 107.400 233.100 110.100 ;
        RECT 218.700 106.500 227.550 107.400 ;
        RECT 218.700 105.600 220.800 106.500 ;
        RECT 223.650 104.700 225.750 105.600 ;
        RECT 218.700 103.500 225.750 104.700 ;
        RECT 218.700 102.600 220.800 103.500 ;
        RECT 216.150 99.000 218.250 101.100 ;
        RECT 222.750 99.600 224.850 101.700 ;
        RECT 226.650 101.400 227.550 106.500 ;
        RECT 228.450 105.300 230.550 107.400 ;
        RECT 231.450 105.300 233.550 107.400 ;
        RECT 228.900 102.900 230.100 105.300 ;
        RECT 235.200 103.800 236.100 112.800 ;
        RECT 237.450 109.200 239.550 111.300 ;
        RECT 240.900 110.400 242.100 113.100 ;
        RECT 238.650 106.800 239.550 109.200 ;
        RECT 240.450 108.300 242.550 110.400 ;
        RECT 244.350 106.800 245.550 114.000 ;
        RECT 238.650 105.600 245.550 106.800 ;
        RECT 241.650 103.800 243.750 104.700 ;
        RECT 235.200 102.600 243.750 103.800 ;
        RECT 45.450 95.100 47.550 97.200 ;
        RECT 222.900 96.900 224.100 99.600 ;
        RECT 226.200 99.300 228.300 101.400 ;
        RECT 236.700 100.800 238.800 102.600 ;
        RECT 240.450 99.600 242.550 101.700 ;
        RECT 244.650 100.200 245.550 105.600 ;
        RECT 246.450 105.300 248.550 107.400 ;
        RECT 246.900 102.900 248.100 105.300 ;
        RECT 240.900 96.900 242.100 99.600 ;
        RECT 243.900 98.100 246.000 100.200 ;
        RECT 108.300 76.800 110.400 78.900 ;
        RECT 111.300 76.800 113.400 78.900 ;
        RECT 6.450 73.200 8.550 75.300 ;
        RECT 24.300 73.800 26.400 75.900 ;
        RECT 7.050 66.600 8.100 73.200 ;
        RECT 9.450 70.200 11.550 72.300 ;
        RECT 6.450 64.500 8.550 66.600 ;
        RECT 3.450 60.450 5.550 62.550 ;
        RECT 3.900 57.900 5.100 60.450 ;
        RECT 7.050 53.100 8.100 64.500 ;
        RECT 10.050 58.200 11.400 70.200 ;
        RECT 24.300 66.600 25.500 73.800 ;
        RECT 39.450 72.900 41.550 75.000 ;
        RECT 60.450 73.800 62.550 75.900 ;
        RECT 84.450 74.100 86.550 76.200 ;
        RECT 87.450 74.100 89.550 76.200 ;
        RECT 90.450 74.100 92.550 76.200 ;
        RECT 24.300 64.500 26.400 66.600 ;
        RECT 15.900 59.550 17.100 62.100 ;
        RECT 9.450 56.100 11.550 58.200 ;
        RECT 15.450 57.450 17.550 59.550 ;
        RECT 6.450 51.000 8.550 53.100 ;
        RECT 24.300 52.200 25.500 64.500 ;
        RECT 36.900 62.550 38.100 65.100 ;
        RECT 30.450 60.450 32.550 62.550 ;
        RECT 36.450 60.450 38.550 62.550 ;
        RECT 30.900 57.900 32.100 60.450 ;
        RECT 40.200 53.100 41.400 72.900 ;
        RECT 60.450 70.200 61.650 73.800 ;
        RECT 60.450 68.100 62.550 70.200 ;
        RECT 45.900 62.550 47.100 65.100 ;
        RECT 45.450 60.450 47.550 62.550 ;
        RECT 60.450 53.100 61.650 68.100 ;
        RECT 72.900 65.400 74.100 68.100 ;
        RECT 72.450 63.300 74.550 65.400 ;
        RECT 78.450 63.300 80.550 65.400 ;
        RECT 63.450 60.450 65.550 62.550 ;
        RECT 78.900 60.900 80.100 63.300 ;
        RECT 63.900 57.900 65.100 60.450 ;
        RECT 84.900 53.100 86.100 74.100 ;
        RECT 87.900 70.800 89.100 74.100 ;
        RECT 87.450 68.700 89.550 70.800 ;
        RECT 88.350 53.100 89.550 68.700 ;
        RECT 91.350 53.100 92.550 74.100 ;
        RECT 99.450 72.300 101.550 74.400 ;
        RECT 105.450 73.800 107.550 75.900 ;
        RECT 99.450 66.900 100.650 72.300 ;
        RECT 105.450 66.900 106.650 73.800 ;
        RECT 109.200 72.000 110.400 76.800 ;
        RECT 112.350 73.800 113.400 76.800 ;
        RECT 114.450 76.800 116.550 78.900 ;
        RECT 108.450 69.900 110.550 72.000 ;
        RECT 99.450 64.800 101.550 66.900 ;
        RECT 105.450 64.800 107.550 66.900 ;
        RECT 96.900 59.400 98.100 62.100 ;
        RECT 96.300 57.300 98.400 59.400 ;
        RECT 100.050 53.100 101.250 64.800 ;
        RECT 105.450 53.100 106.650 64.800 ;
        RECT 109.050 53.100 110.550 69.900 ;
        RECT 112.350 53.100 113.550 73.800 ;
        RECT 24.300 50.100 26.400 52.200 ;
        RECT 39.450 51.000 41.550 53.100 ;
        RECT 60.450 51.000 62.550 53.100 ;
        RECT 84.450 51.000 86.550 53.100 ;
        RECT 87.450 51.000 89.550 53.100 ;
        RECT 90.450 51.000 92.550 53.100 ;
        RECT 99.450 51.000 101.550 53.100 ;
        RECT 105.450 51.000 107.550 53.100 ;
        RECT 108.450 51.000 110.550 53.100 ;
        RECT 111.450 51.000 113.550 53.100 ;
        RECT 114.450 72.000 115.650 76.800 ;
        RECT 114.450 69.900 116.550 72.000 ;
        RECT 175.500 71.100 177.600 71.550 ;
        RECT 147.450 70.200 177.600 71.100 ;
        RECT 114.450 53.100 115.650 69.900 ;
        RECT 147.450 69.000 149.550 70.200 ;
        RECT 126.450 63.300 128.550 65.400 ;
        RECT 135.450 63.300 137.550 65.400 ;
        RECT 126.900 60.900 128.100 63.300 ;
        RECT 135.900 60.900 137.100 63.300 ;
        RECT 144.900 62.550 146.100 65.100 ;
        RECT 141.450 60.450 143.550 62.550 ;
        RECT 144.450 60.450 146.550 62.550 ;
        RECT 141.900 57.900 143.100 60.450 ;
        RECT 148.050 54.900 148.950 69.000 ;
        RECT 159.450 66.900 161.550 70.200 ;
        RECT 175.500 69.450 177.600 70.200 ;
        RECT 162.450 66.900 164.550 69.000 ;
        RECT 163.050 55.800 164.250 66.900 ;
        RECT 177.900 62.550 179.100 65.100 ;
        RECT 168.450 60.450 170.550 62.550 ;
        RECT 174.450 60.450 176.550 62.550 ;
        RECT 177.450 60.450 179.550 62.550 ;
        RECT 231.450 60.450 233.550 62.550 ;
        RECT 237.450 60.750 239.550 62.850 ;
        RECT 240.900 62.550 242.100 65.100 ;
        RECT 246.900 62.550 248.100 65.100 ;
        RECT 168.900 57.900 170.100 60.450 ;
        RECT 174.900 57.900 176.100 60.450 ;
        RECT 231.900 57.900 233.100 60.450 ;
        RECT 114.450 51.000 116.550 53.100 ;
        RECT 147.450 52.800 149.550 54.900 ;
        RECT 162.450 53.700 164.550 55.800 ;
        RECT 237.900 55.200 238.950 60.750 ;
        RECT 240.450 60.450 242.550 62.550 ;
        RECT 246.450 60.450 248.550 62.550 ;
        RECT 252.450 60.450 254.550 62.550 ;
        RECT 237.450 53.100 239.550 55.200 ;
        RECT 241.200 52.200 242.400 60.450 ;
        RECT 252.900 57.900 254.100 60.450 ;
        RECT 239.700 50.100 242.400 52.200 ;
        RECT 0.900 17.550 2.100 20.100 ;
        RECT 9.900 17.550 11.100 20.100 ;
        RECT 0.450 15.450 2.550 17.550 ;
        RECT 6.450 15.450 8.550 17.550 ;
        RECT 9.450 15.450 11.550 17.550 ;
        RECT 14.700 17.400 15.900 20.100 ;
        RECT 23.700 17.400 24.900 20.100 ;
        RECT 28.500 17.400 29.700 20.100 ;
        RECT 34.500 17.400 35.700 20.100 ;
        RECT 42.300 17.400 43.500 20.100 ;
        RECT 48.300 17.400 49.500 20.100 ;
        RECT 54.300 17.400 55.500 20.100 ;
        RECT 65.100 17.550 66.300 20.100 ;
        RECT 78.900 17.550 80.100 20.100 ;
        RECT 6.900 12.900 8.100 15.450 ;
        RECT 14.250 15.300 16.350 17.400 ;
        RECT 20.250 15.300 22.350 17.400 ;
        RECT 23.250 15.300 25.350 17.400 ;
        RECT 28.050 15.300 30.150 17.400 ;
        RECT 31.050 15.300 33.150 17.400 ;
        RECT 34.050 15.300 36.150 17.400 ;
        RECT 37.050 15.300 39.150 17.400 ;
        RECT 41.850 15.300 43.950 17.400 ;
        RECT 44.850 15.300 46.950 17.400 ;
        RECT 47.850 15.300 49.950 17.400 ;
        RECT 50.850 15.300 52.950 17.400 ;
        RECT 53.850 15.300 55.950 17.400 ;
        RECT 58.650 15.450 60.750 17.550 ;
        RECT 64.650 15.450 66.750 17.550 ;
        RECT 69.450 15.450 71.550 17.550 ;
        RECT 78.450 15.450 80.550 17.550 ;
        RECT 86.700 17.400 87.900 20.100 ;
        RECT 107.700 17.400 108.900 20.100 ;
        RECT 114.600 17.550 115.800 20.100 ;
        RECT 147.600 17.550 148.800 20.100 ;
        RECT 153.600 17.550 154.800 20.100 ;
        RECT 198.600 17.550 199.800 20.100 ;
        RECT 20.700 12.900 21.900 15.300 ;
        RECT 31.500 12.900 32.700 15.300 ;
        RECT 37.500 12.900 38.700 15.300 ;
        RECT 45.300 12.900 46.500 15.300 ;
        RECT 51.300 12.900 52.500 15.300 ;
        RECT 59.100 12.900 60.300 15.450 ;
        RECT 69.900 12.900 71.100 15.450 ;
        RECT 86.250 15.300 88.350 17.400 ;
        RECT 107.250 15.300 109.350 17.400 ;
        RECT 114.150 15.450 116.250 17.550 ;
        RECT 147.150 15.450 149.250 17.550 ;
        RECT 153.150 15.450 155.250 17.550 ;
        RECT 198.150 15.450 200.250 17.550 ;
  END
END khu_etri050_stdcells
