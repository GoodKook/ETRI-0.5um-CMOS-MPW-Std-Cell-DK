magic
tech scmos
magscale 1 2
timestamp 1727422155
<< nwell >>
rect -13 154 112 272
<< ntransistor >>
rect 20 14 24 54
rect 28 14 32 54
rect 50 14 54 34
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 60 206 64 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 28 54
rect 32 14 34 54
rect 46 14 50 34
rect 54 14 56 34
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 206 46 246
rect 58 206 60 246
rect 64 206 66 246
<< ndcontact >>
rect 6 14 18 54
rect 34 14 46 54
rect 56 14 68 34
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 46 206 58 246
rect 66 206 78 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 123 24 206
rect 16 111 24 123
rect 20 54 24 111
rect 40 87 44 206
rect 60 202 64 206
rect 60 198 68 202
rect 28 80 44 87
rect 28 54 32 80
rect 64 72 68 198
rect 56 60 68 72
rect 50 34 54 60
rect 20 10 24 14
rect 28 10 32 14
rect 50 10 54 14
<< polycontact >>
rect 4 111 16 123
rect 44 157 56 169
rect 44 60 56 72
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 6 246 18 252
rect 46 246 58 252
rect 3 123 17 137
rect 27 72 34 206
rect 43 143 57 157
rect 66 117 74 206
rect 63 103 77 117
rect 6 64 44 72
rect 6 54 18 64
rect 63 39 70 103
rect 56 34 70 39
rect 34 8 46 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 43 143 57 157
rect 3 123 17 137
rect 63 103 77 117
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 43 143 57 157 0 B
port 1 nsew signal input
rlabel metal1 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal1 63 103 77 117 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
