magic
tech scmos
magscale 1 3
timestamp 1725342160
<< polysilicon >>
rect 2 104 142 122
rect 2 20 123 104
rect 135 20 142 104
rect 2 2 142 20
<< polycontact >>
rect 123 20 135 104
<< genericcontact >>
rect 23 95 29 101
rect 35 95 41 101
rect 47 95 53 101
rect 59 95 65 101
rect 71 95 77 101
rect 83 95 89 101
rect 95 95 101 101
rect 23 83 29 89
rect 35 83 41 89
rect 47 83 53 89
rect 59 83 65 89
rect 71 83 77 89
rect 83 83 89 89
rect 95 83 101 89
rect 23 71 29 77
rect 35 71 41 77
rect 47 71 53 77
rect 59 71 65 77
rect 71 71 77 77
rect 83 71 89 77
rect 95 71 101 77
rect 23 59 29 65
rect 35 59 41 65
rect 47 59 53 65
rect 59 59 65 65
rect 71 59 77 65
rect 83 59 89 65
rect 95 59 101 65
rect 23 47 29 53
rect 35 47 41 53
rect 47 47 53 53
rect 59 47 65 53
rect 71 47 77 53
rect 83 47 89 53
rect 95 47 101 53
rect 23 35 29 41
rect 35 35 41 41
rect 47 35 53 41
rect 59 35 65 41
rect 71 35 77 41
rect 83 35 89 41
rect 95 35 101 41
rect 23 23 29 29
rect 35 23 41 29
rect 47 23 53 29
rect 59 23 65 29
rect 71 23 77 29
rect 83 23 89 29
rect 95 23 101 29
<< metal1 >>
rect 16 16 108 108
rect 120 104 138 108
rect 120 20 123 104
rect 135 20 138 104
rect 120 16 138 20
<< pseudo_rpoly2 >>
rect 12 12 112 112
<< end >>
