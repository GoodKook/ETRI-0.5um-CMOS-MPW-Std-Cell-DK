magic
tech scmos
magscale 1 3
timestamp 1725338064
<< checkpaint >>
rect -15 430 430 455
rect -15 10 455 430
rect 16 -14 424 10
<< nwell >>
rect 110 110 330 330
<< psubstratepdiff >>
rect 45 375 395 395
rect 45 65 65 375
rect 195 195 245 245
rect 375 65 395 375
rect 45 45 395 65
<< nsubstratendiff >>
rect 130 290 310 310
rect 130 150 150 290
rect 290 150 310 290
rect 130 130 310 150
<< genericcontact >>
rect 70 375 370 395
rect 45 70 65 370
rect 150 290 290 310
rect 130 150 150 290
rect 195 195 245 245
rect 290 150 310 290
rect 150 130 290 150
rect 375 70 395 370
rect 70 45 370 65
<< metal1 >>
rect 45 375 395 395
rect 45 65 65 375
rect 130 290 310 310
rect 130 150 150 290
rect 195 195 245 245
rect 290 150 310 290
rect 130 130 310 150
rect 375 65 395 375
rect 45 45 395 65
<< end >>
