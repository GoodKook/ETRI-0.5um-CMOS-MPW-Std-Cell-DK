magic
tech scmos
magscale 1 2
timestamp 1702314024
<< checkpaint >>
rect 26 180 114 181
rect -18 83 117 180
rect -18 81 114 83
rect -18 65 77 81
<< nwell >>
rect -13 154 114 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
rect 78 14 82 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 58 166 62 246
rect 78 166 82 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 36 14 38 54
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
rect 76 14 78 54
rect 82 14 84 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
rect 36 166 38 246
rect 42 166 44 246
rect 56 166 58 246
rect 62 166 64 246
rect 76 166 78 246
rect 82 166 84 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
rect 64 14 76 54
rect 84 14 96 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
rect 44 166 56 246
rect 64 166 76 246
rect 84 166 96 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 78 246 82 250
rect 18 164 22 166
rect 38 164 42 166
rect 58 164 62 166
rect 78 164 82 166
rect 18 160 82 164
rect 18 117 22 160
rect 18 105 24 117
rect 18 62 22 105
rect 18 58 82 62
rect 18 54 22 58
rect 38 54 42 58
rect 58 54 62 58
rect 78 54 82 58
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
rect 78 10 82 14
<< polycontact >>
rect 24 105 36 117
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 4 246 16 252
rect 44 246 56 252
rect 84 246 96 252
rect 24 160 36 166
rect 64 160 74 166
rect 24 154 74 160
rect 66 137 74 154
rect 23 123 37 137
rect 63 123 77 137
rect 24 117 36 123
rect 66 68 74 123
rect 24 60 74 68
rect 24 54 32 60
rect 64 54 74 60
rect 4 8 16 14
rect 44 8 56 14
rect 84 8 96 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect -6 252 106 268
rect 23 123 37 137
rect 63 123 77 137
rect -6 -8 106 8
<< labels >>
rlabel nsubstratencontact 50 260 50 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 50 0 50 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 70 130 70 130 0 Y
port 2 nsew signal output
rlabel metal1 30 127 30 127 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
