magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 154 132 272
<< ntransistor >>
rect 22 14 26 54
rect 32 14 36 54
rect 52 14 56 54
rect 62 14 66 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 32 54
rect 36 14 38 54
rect 50 14 52 54
rect 56 14 62 54
rect 66 14 68 54
<< pdiffusion >>
rect 18 168 20 246
rect 6 166 20 168
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 168 46 246
rect 58 168 60 246
rect 44 166 60 168
rect 64 234 80 246
rect 64 166 66 234
rect 78 166 80 234
rect 84 166 86 246
<< ndcontact >>
rect 8 14 20 54
rect 38 14 50 54
rect 68 14 80 54
<< pdcontact >>
rect 6 168 18 246
rect 26 180 38 246
rect 46 168 58 246
rect 66 166 78 234
rect 86 166 98 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 20 144 24 166
rect 40 144 44 166
rect 6 138 24 144
rect 32 138 44 144
rect 60 144 64 166
rect 80 144 84 166
rect 60 138 68 144
rect 80 138 90 144
rect 6 103 12 138
rect 32 109 36 138
rect 6 64 12 91
rect 6 60 26 64
rect 22 54 26 60
rect 32 54 36 97
rect 62 109 68 138
rect 62 97 64 109
rect 84 103 90 138
rect 62 76 68 97
rect 52 72 68 76
rect 52 54 56 72
rect 84 64 90 91
rect 62 60 90 64
rect 62 54 66 60
rect 22 10 26 14
rect 32 10 36 14
rect 52 10 56 14
rect 62 10 66 14
<< polycontact >>
rect 4 91 16 103
rect 24 97 36 109
rect 64 97 76 109
rect 84 91 96 103
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 26 246 38 252
rect 18 168 46 174
rect 58 240 86 246
rect 66 160 78 166
rect 44 154 78 160
rect 44 117 50 154
rect 43 54 50 103
rect 8 8 20 14
rect 68 8 80 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 103 17 117
rect 43 103 57 117
rect 23 83 37 97
rect 83 103 97 117
rect 63 83 77 97
<< metal2 >>
rect 3 117 17 137
rect 43 117 57 137
rect 83 117 97 137
rect 23 63 37 83
rect 63 63 77 83
<< m2p >>
rect 3 123 17 137
rect 43 123 57 137
rect 83 123 97 137
rect 23 63 37 77
rect 63 63 77 77
<< labels >>
rlabel metal2 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal2 23 63 37 77 0 B
port 1 nsew signal input
rlabel metal2 83 123 97 137 0 C
port 2 nsew signal input
rlabel metal2 63 63 77 77 0 D
port 3 nsew signal input
rlabel metal2 43 123 57 137 0 Y
port 4 nsew signal output
rlabel metal1 -6 252 126 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 126 8 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
