magic
tech scmos
magscale 1 2
timestamp 1727045892
<< metal1 >>
rect -63 11978 -3 12238
rect 12310 12222 12403 12238
rect 2127 12157 2313 12163
rect 8487 12157 8673 12163
rect 3647 12097 3793 12103
rect 11017 12100 11073 12103
rect 11013 12097 11073 12100
rect 11013 12087 11027 12097
rect 487 12077 733 12083
rect 1587 12077 1773 12083
rect 3587 12077 3753 12083
rect 6727 12057 6763 12063
rect 3340 12023 3353 12027
rect 3337 12017 3353 12023
rect 3340 12013 3353 12017
rect 5160 12023 5173 12027
rect 5157 12017 5173 12023
rect 5160 12013 5173 12017
rect 8440 12023 8453 12027
rect 8437 12017 8453 12023
rect 8440 12013 8453 12017
rect -63 11962 30 11978
rect -63 11458 -3 11962
rect 5207 11917 5243 11923
rect 1967 11857 1993 11863
rect 7607 11857 7713 11863
rect 10567 11857 10753 11863
rect 307 11837 333 11843
rect 2267 11837 2433 11843
rect 5067 11777 5233 11783
rect 9287 11777 9473 11783
rect 12343 11718 12403 12222
rect 12310 11702 12403 11718
rect 1187 11637 1313 11643
rect 6907 11617 7033 11623
rect 5387 11597 5453 11603
rect 847 11577 893 11583
rect 2467 11577 2613 11583
rect 527 11557 733 11563
rect 2507 11557 2673 11563
rect 3447 11557 3493 11563
rect 4747 11557 4833 11563
rect 5847 11557 5873 11563
rect 7687 11557 7733 11563
rect 4407 11517 4453 11523
rect 2437 11497 2473 11503
rect 4597 11497 4673 11503
rect 4787 11497 4843 11503
rect 9947 11497 10003 11503
rect 4433 11483 4447 11493
rect 4367 11480 4447 11483
rect 4367 11477 4443 11480
rect -63 11442 30 11458
rect -63 10938 -3 11442
rect 4207 11417 4243 11423
rect 5080 11403 5093 11407
rect 5077 11397 5093 11403
rect 5080 11393 5093 11397
rect 7657 11397 7693 11403
rect 9240 11403 9253 11407
rect 9237 11397 9253 11403
rect 9240 11393 9253 11397
rect 747 11337 833 11343
rect 2967 11337 3033 11343
rect 3747 11337 3813 11343
rect 6687 11317 6833 11323
rect 10707 11277 10813 11283
rect 6307 11257 6333 11263
rect 6487 11217 6553 11223
rect 12343 11198 12403 11702
rect 12310 11182 12403 11198
rect 9547 11117 9693 11123
rect 11687 11117 11773 11123
rect 3987 11097 4133 11103
rect 2467 11077 2593 11083
rect 4487 11037 4633 11043
rect 4647 11037 4693 11043
rect 4887 11037 4973 11043
rect 6267 11037 6373 11043
rect 2487 11017 2573 11023
rect 3660 10983 3673 10987
rect 3657 10977 3673 10983
rect 3660 10973 3673 10977
rect 6900 10983 6913 10987
rect 6897 10977 6913 10983
rect 6900 10973 6913 10977
rect 8940 10983 8953 10987
rect 8937 10977 8953 10983
rect 8940 10973 8953 10977
rect -63 10922 30 10938
rect -63 10418 -3 10922
rect 3260 10883 3273 10887
rect 3257 10877 3273 10883
rect 3260 10873 3273 10877
rect 1367 10837 1573 10843
rect 1507 10817 1613 10823
rect 3527 10817 3553 10823
rect 8147 10817 8213 10823
rect 8727 10817 8873 10823
rect 11580 10803 11593 10807
rect 11577 10793 11593 10803
rect 5407 10777 5473 10783
rect 11577 10767 11583 10793
rect 627 10757 653 10763
rect 9787 10757 9813 10763
rect 11577 10757 11593 10767
rect 11580 10753 11593 10757
rect 10907 10717 11053 10723
rect 11227 10717 11333 10723
rect 4187 10697 4253 10703
rect 12343 10678 12403 11182
rect 12310 10662 12403 10678
rect 4367 10597 4413 10603
rect 4307 10577 4393 10583
rect 4847 10577 4953 10583
rect 6007 10577 6133 10583
rect 4627 10537 4733 10543
rect 4547 10517 4713 10523
rect 4967 10517 5013 10523
rect 8447 10517 8513 10523
rect 11227 10517 11413 10523
rect 11767 10517 11953 10523
rect 1597 10497 1733 10503
rect 2527 10497 2613 10503
rect 4367 10497 4463 10503
rect 7647 10497 7693 10503
rect 10947 10497 11093 10503
rect 2407 10477 2513 10483
rect 11047 10477 11153 10483
rect 5657 10457 5713 10463
rect 5937 10457 5973 10463
rect 7147 10457 7183 10463
rect -63 10402 30 10418
rect -63 9898 -3 10402
rect 3787 10377 3933 10383
rect 3187 10357 3223 10363
rect 4847 10357 4973 10363
rect 3807 10337 3973 10343
rect 4967 10317 5023 10323
rect 827 10297 1013 10303
rect 3847 10297 3973 10303
rect 5747 10297 5773 10303
rect 9987 10297 10073 10303
rect 10087 10297 10133 10303
rect 2327 10277 2413 10283
rect 7080 10283 7093 10287
rect 7077 10273 7093 10283
rect 3767 10257 3793 10263
rect 7077 10247 7083 10273
rect 7077 10237 7093 10247
rect 7080 10233 7093 10237
rect 9727 10237 9833 10243
rect 2247 10217 2353 10223
rect 3087 10217 3193 10223
rect 3827 10217 3933 10223
rect 5667 10217 5813 10223
rect 8707 10217 8733 10223
rect 3027 10197 3153 10203
rect 8967 10177 9013 10183
rect 12343 10158 12403 10662
rect 12310 10142 12403 10158
rect 7847 10117 7933 10123
rect 5667 10077 5833 10083
rect 3887 10057 3913 10063
rect 7007 10057 7153 10063
rect 2407 10017 2513 10023
rect 7033 10023 7047 10033
rect 7007 10017 7193 10023
rect 1067 9997 1253 10003
rect 5887 9997 6033 10003
rect 7267 9997 7373 10003
rect 7387 9997 7433 10003
rect 11167 9997 11233 10003
rect 6607 9977 6643 9983
rect 3577 9937 3613 9943
rect 4147 9943 4160 9947
rect 4147 9937 4163 9943
rect 4147 9933 4160 9937
rect 8247 9937 8283 9943
rect -63 9882 30 9898
rect -63 9378 -3 9882
rect 3867 9857 3893 9863
rect 7067 9857 7113 9863
rect 7567 9860 7703 9863
rect 7567 9857 7707 9860
rect 7693 9847 7707 9857
rect 7287 9817 7453 9823
rect 7247 9797 7453 9803
rect 9607 9797 9813 9803
rect 1207 9777 1253 9783
rect 1327 9777 1433 9783
rect 3827 9777 3913 9783
rect 8567 9777 8733 9783
rect 11647 9777 11693 9783
rect 2547 9757 2633 9763
rect 3880 9763 3893 9767
rect 3877 9753 3893 9763
rect 4587 9757 4653 9763
rect 7367 9757 7413 9763
rect 10987 9763 11000 9767
rect 10987 9753 11003 9763
rect 2287 9717 2333 9723
rect 3877 9706 3883 9753
rect 10997 9727 11003 9753
rect 10047 9717 10093 9723
rect 10987 9717 11003 9727
rect 10987 9713 11000 9717
rect 12167 9717 12193 9723
rect 6667 9697 6773 9703
rect 6947 9697 7093 9703
rect 4787 9657 4913 9663
rect 12343 9638 12403 10142
rect 12310 9622 12403 9638
rect 3047 9597 3173 9603
rect 247 9557 273 9563
rect 10087 9557 10173 9563
rect 2187 9537 2353 9543
rect 7587 9537 7693 9543
rect 9447 9537 9593 9543
rect 8627 9497 8693 9503
rect 487 9477 693 9483
rect 3047 9477 3093 9483
rect 3747 9477 3913 9483
rect 7247 9477 7473 9483
rect 2787 9457 2903 9463
rect 5987 9457 6153 9463
rect 8487 9457 8543 9463
rect 9787 9457 9833 9463
rect 9947 9457 9993 9463
rect 3147 9437 3193 9443
rect 3977 9417 4073 9423
rect 7687 9397 7723 9403
rect -63 9362 30 9378
rect -63 8858 -3 9362
rect 5127 9337 5253 9343
rect 4257 9317 4293 9323
rect 4427 9297 4463 9303
rect 6747 9297 6893 9303
rect 10927 9297 11013 9303
rect 10967 9277 11133 9283
rect 11247 9277 11313 9283
rect 1687 9257 1753 9263
rect 2167 9257 2333 9263
rect 6967 9257 7173 9263
rect 8787 9257 8913 9263
rect 11787 9257 11833 9263
rect 5107 9237 5133 9243
rect 8927 9237 8993 9243
rect 4607 9197 4733 9203
rect 5627 9197 5753 9203
rect 7067 9197 7113 9203
rect 7127 9197 7153 9203
rect 7247 9197 7373 9203
rect 1887 9177 1933 9183
rect 8587 9177 8733 9183
rect 11267 9177 11353 9183
rect 11367 9177 11433 9183
rect 8567 9157 8693 9163
rect 12343 9118 12403 9622
rect 12310 9102 12403 9118
rect 6127 9077 6213 9083
rect 8647 9037 8813 9043
rect 5127 9023 5140 9027
rect 5127 9013 5143 9023
rect 10807 9017 10893 9023
rect 3793 8987 3807 8993
rect 5137 8987 5143 9013
rect 3793 8980 3813 8987
rect 3797 8977 3813 8980
rect 3800 8973 3813 8977
rect 5127 8977 5143 8987
rect 5127 8973 5140 8977
rect 1067 8957 1233 8963
rect 2367 8957 2453 8963
rect 3087 8957 3133 8963
rect 3747 8957 3773 8963
rect 5387 8957 5533 8963
rect 11347 8957 11453 8963
rect 12167 8957 12193 8963
rect 3727 8937 3833 8943
rect 3767 8917 3843 8923
rect 3407 8897 3513 8903
rect 3837 8897 3843 8917
rect 5247 8917 5273 8923
rect 3080 8883 3093 8887
rect 3077 8877 3093 8883
rect 3080 8873 3093 8877
rect -63 8842 30 8858
rect -63 8338 -3 8842
rect 2007 8817 2053 8823
rect 6127 8817 6253 8823
rect 8587 8817 8673 8823
rect 8687 8817 8713 8823
rect 8827 8817 8953 8823
rect 3787 8777 3993 8783
rect 1427 8737 1573 8743
rect 3407 8737 3433 8743
rect 3787 8737 3893 8743
rect 4847 8737 4953 8743
rect 7507 8737 7613 8743
rect 7987 8737 8053 8743
rect 8847 8737 8893 8743
rect 9207 8737 9293 8743
rect 11087 8737 11193 8743
rect 6227 8717 6293 8723
rect 9907 8717 10013 8723
rect 2507 8697 2533 8703
rect 5167 8697 5253 8703
rect 2707 8677 2873 8683
rect 6187 8677 6293 8683
rect 807 8657 1033 8663
rect 2487 8657 2613 8663
rect 6427 8657 6573 8663
rect 12343 8598 12403 9102
rect 12310 8582 12403 8598
rect 4567 8537 4653 8543
rect 3747 8517 3933 8523
rect 6467 8517 6613 8523
rect 10927 8517 11013 8523
rect 11027 8517 11053 8523
rect 12067 8517 12213 8523
rect 12267 8517 12313 8523
rect 347 8497 413 8503
rect 6967 8457 7093 8463
rect 2787 8437 2973 8443
rect 3887 8437 3953 8443
rect 4507 8437 4613 8443
rect 8253 8443 8267 8453
rect 8253 8440 8453 8443
rect 8257 8437 8453 8440
rect 9607 8437 9733 8443
rect 10367 8437 10593 8443
rect 5857 8377 5893 8383
rect 2387 8357 2423 8363
rect 5307 8357 5453 8363
rect 5887 8357 5933 8363
rect -63 8322 30 8338
rect -63 7818 -3 8322
rect 8060 8283 8073 8287
rect 8057 8277 8073 8283
rect 8060 8273 8073 8277
rect 9427 8277 9493 8283
rect 1677 8237 1713 8243
rect 9397 8237 9433 8243
rect 11527 8237 11553 8243
rect 1107 8217 1133 8223
rect 1387 8217 1493 8223
rect 2267 8217 2433 8223
rect 4207 8217 4253 8223
rect 4747 8217 4833 8223
rect 9787 8217 9893 8223
rect 11467 8217 11493 8223
rect 11507 8217 11633 8223
rect 2400 8203 2413 8207
rect 2397 8193 2413 8203
rect 6827 8197 6933 8203
rect 2397 8167 2403 8193
rect 2397 8157 2413 8167
rect 2400 8153 2413 8157
rect 4347 8157 4373 8163
rect 4907 8157 4933 8163
rect 11587 8137 11693 8143
rect 2267 8097 2333 8103
rect 9167 8097 9233 8103
rect 12343 8078 12403 8582
rect 12310 8062 12403 8078
rect 5527 8037 5613 8043
rect 8627 8037 8653 8043
rect 2127 7997 2253 8003
rect 2947 7997 3053 8003
rect 3687 7997 3833 8003
rect 6787 7997 6853 8003
rect 8307 7997 8373 8003
rect 2247 7977 2273 7983
rect 7107 7977 7253 7983
rect 8960 7983 8973 7987
rect 8957 7973 8973 7983
rect 10507 7977 10613 7983
rect 11327 7977 11473 7983
rect 11567 7977 11693 7983
rect 8957 7947 8963 7973
rect 2127 7937 2273 7943
rect 8957 7937 8973 7947
rect 8960 7933 8973 7937
rect 2107 7917 2253 7923
rect 3347 7917 3493 7923
rect 3507 7917 3573 7923
rect 2147 7897 2233 7903
rect 2287 7903 2300 7907
rect 2287 7897 2303 7903
rect 2287 7893 2300 7897
rect 5467 7897 5593 7903
rect 10387 7897 10443 7903
rect 10240 7863 10253 7867
rect 10237 7857 10253 7863
rect 10240 7853 10253 7857
rect -63 7802 30 7818
rect -63 7298 -3 7802
rect 4767 7777 4813 7783
rect 5400 7763 5413 7767
rect 5397 7757 5413 7763
rect 5400 7753 5413 7757
rect 9597 7757 9653 7763
rect 5977 7717 6053 7723
rect 5667 7697 5853 7703
rect 867 7677 1013 7683
rect 3007 7677 3093 7683
rect 9387 7677 9513 7683
rect 5707 7637 5873 7643
rect 7307 7637 7393 7643
rect 367 7617 493 7623
rect 5687 7617 5713 7623
rect 7047 7577 7193 7583
rect 12343 7558 12403 8062
rect 12310 7542 12403 7558
rect 7207 7517 7293 7523
rect 11107 7497 11233 7503
rect 6427 7477 6533 7483
rect 7367 7477 7573 7483
rect 2787 7463 2800 7467
rect 2787 7453 2803 7463
rect 3607 7457 3713 7463
rect 10660 7463 10673 7467
rect 10657 7453 10673 7463
rect 12087 7457 12113 7463
rect 2797 7427 2803 7453
rect 7127 7437 7293 7443
rect 7447 7437 7573 7443
rect 10657 7427 10663 7453
rect 627 7417 713 7423
rect 2787 7417 2803 7427
rect 2787 7413 2800 7417
rect 3527 7417 3713 7423
rect 10657 7417 10673 7427
rect 10660 7413 10673 7417
rect 547 7397 753 7403
rect 1707 7397 1733 7403
rect 3667 7397 3733 7403
rect 6467 7397 6533 7403
rect 7447 7397 7533 7403
rect 9807 7397 9933 7403
rect 6127 7377 6213 7383
rect 1947 7357 2033 7363
rect 7427 7357 7593 7363
rect -63 7282 30 7298
rect -63 6778 -3 7282
rect 5687 7257 5813 7263
rect 6787 7257 6873 7263
rect 7087 7257 7233 7263
rect 9920 7243 9933 7247
rect 9917 7237 9933 7243
rect 9920 7233 9933 7237
rect 3847 7217 3933 7223
rect 5407 7217 5593 7223
rect 4627 7197 4763 7203
rect 5307 7197 5343 7203
rect 1787 7177 1833 7183
rect 4827 7177 4993 7183
rect 7227 7177 7273 7183
rect 8267 7177 8293 7183
rect 4407 7157 4453 7163
rect 4847 7157 4893 7163
rect 5427 7157 5573 7163
rect 307 7117 433 7123
rect 3327 7117 3393 7123
rect 3507 7117 3613 7123
rect 4927 7117 5033 7123
rect 907 7097 933 7103
rect 3727 7097 3893 7103
rect 4847 7097 4933 7103
rect 5507 7097 5533 7103
rect 7887 7097 7993 7103
rect 8187 7097 8293 7103
rect 9987 7097 10113 7103
rect 10427 7097 10533 7103
rect 10547 7097 10613 7103
rect 11787 7097 12053 7103
rect 5487 7077 5613 7083
rect 7147 7077 7233 7083
rect 12343 7038 12403 7542
rect 12310 7022 12403 7038
rect 11067 6977 11093 6983
rect 847 6957 953 6963
rect 10607 6957 10753 6963
rect 11787 6957 11833 6963
rect 11887 6957 11913 6963
rect 3627 6937 3713 6943
rect 6747 6937 6893 6943
rect 8387 6917 8473 6923
rect 6207 6897 6233 6903
rect 9487 6897 9553 6903
rect 1967 6877 2013 6883
rect 4067 6877 4113 6883
rect 5967 6877 6033 6883
rect 7007 6877 7213 6883
rect 7487 6877 7513 6883
rect 1917 6857 1973 6863
rect 7367 6857 7513 6863
rect 11907 6837 12073 6843
rect 8037 6817 8113 6823
rect -63 6762 30 6778
rect -63 6258 -3 6762
rect 9253 6723 9267 6733
rect 9147 6720 9267 6723
rect 9147 6717 9263 6720
rect 4167 6697 4193 6703
rect 10207 6697 10253 6703
rect 10267 6697 10293 6703
rect 1417 6677 1533 6683
rect 9337 6677 9373 6683
rect 2727 6657 2793 6663
rect 4347 6657 4533 6663
rect 5587 6657 5633 6663
rect 7327 6663 7340 6667
rect 7327 6653 7343 6663
rect 10907 6657 11073 6663
rect 11707 6657 11933 6663
rect 3787 6637 3973 6643
rect 6140 6643 6153 6647
rect 6007 6637 6153 6643
rect 6137 6633 6153 6637
rect 6137 6607 6143 6633
rect 7337 6627 7343 6653
rect 7627 6637 7733 6643
rect 11367 6637 11393 6643
rect 11567 6637 11633 6643
rect 12027 6637 12133 6643
rect 7327 6617 7343 6627
rect 7327 6613 7340 6617
rect 12157 6607 12163 6653
rect 2627 6597 2653 6603
rect 3807 6597 3933 6603
rect 6137 6597 6153 6607
rect 6140 6593 6153 6597
rect 12157 6597 12173 6607
rect 12160 6593 12173 6597
rect 2727 6577 2873 6583
rect 5427 6577 5573 6583
rect 6067 6577 6093 6583
rect 7607 6577 7713 6583
rect 1187 6557 1293 6563
rect 4147 6557 4273 6563
rect 5467 6537 5573 6543
rect 12343 6518 12403 7022
rect 12310 6502 12403 6518
rect 7367 6477 7473 6483
rect 9527 6457 9613 6463
rect 927 6437 1013 6443
rect 2287 6437 2313 6443
rect 2567 6437 2593 6443
rect 10867 6437 11073 6443
rect 11207 6437 11233 6443
rect 11327 6437 11373 6443
rect 4587 6417 4613 6423
rect 6007 6417 6033 6423
rect 7927 6417 8033 6423
rect 8147 6417 8293 6423
rect 10067 6417 10233 6423
rect 11787 6417 11893 6423
rect 12127 6417 12253 6423
rect 4713 6387 4727 6393
rect 4707 6380 4727 6387
rect 4707 6377 4723 6380
rect 4707 6373 4720 6377
rect 4787 6377 4873 6383
rect 6927 6377 6953 6383
rect 12067 6377 12213 6383
rect 1887 6357 1913 6363
rect 1927 6357 2073 6363
rect 2767 6357 2813 6363
rect 3327 6357 3493 6363
rect 4407 6357 4453 6363
rect 6747 6357 6893 6363
rect 8907 6357 9133 6363
rect 8097 6337 8133 6343
rect 2867 6317 2933 6323
rect 3627 6297 3653 6303
rect 5980 6303 5993 6307
rect 5977 6297 5993 6303
rect 5980 6293 5993 6297
rect 8937 6297 9013 6303
rect 8427 6277 8553 6283
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 3007 6217 3073 6223
rect 5127 6217 5293 6223
rect 11527 6177 11593 6183
rect 1687 6157 1753 6163
rect 1827 6157 2053 6163
rect 3867 6157 3893 6163
rect 1647 6140 1763 6143
rect 1647 6137 1767 6140
rect 1753 6127 1767 6137
rect 3227 6137 3453 6143
rect 3887 6137 3973 6143
rect 7087 6137 7273 6143
rect 7587 6137 7653 6143
rect 10187 6137 10233 6143
rect 10947 6137 11053 6143
rect 11527 6137 11653 6143
rect 3807 6117 3893 6123
rect 4307 6117 4353 6123
rect 11207 6117 11323 6123
rect 11317 6087 11323 6117
rect 11447 6117 11533 6123
rect 11587 6117 11613 6123
rect 3907 6077 3973 6083
rect 4407 6077 4473 6083
rect 7327 6077 7393 6083
rect 11317 6077 11333 6087
rect 11320 6073 11333 6077
rect 2007 6057 2033 6063
rect 2387 6057 2433 6063
rect 2947 6057 3013 6063
rect 4947 6057 5053 6063
rect 5107 6057 5173 6063
rect 6007 6057 6153 6063
rect 6587 6057 6753 6063
rect 8647 6057 8813 6063
rect 12127 6057 12173 6063
rect 4887 6037 4953 6043
rect 10387 6037 10513 6043
rect 3553 6023 3567 6033
rect 3527 6020 3567 6023
rect 3527 6017 3563 6020
rect 3827 6017 3933 6023
rect 5687 6017 5753 6023
rect 12343 5998 12403 6502
rect 12310 5982 12403 5998
rect 1427 5957 1533 5963
rect 3267 5917 3433 5923
rect 4107 5917 4273 5923
rect 4427 5917 4573 5923
rect 5747 5917 5933 5923
rect 3307 5897 3413 5903
rect 3847 5897 3933 5903
rect 4447 5897 4533 5903
rect 7147 5897 7253 5903
rect 10187 5897 10233 5903
rect 11227 5897 11373 5903
rect 4147 5857 4213 5863
rect 4953 5863 4967 5873
rect 4927 5860 4967 5863
rect 4927 5857 4963 5860
rect 4987 5857 5093 5863
rect 587 5837 733 5843
rect 4167 5837 4293 5843
rect 5467 5837 5693 5843
rect 5747 5837 5773 5843
rect 7747 5837 7853 5843
rect 8707 5837 8893 5843
rect 11587 5837 11713 5843
rect 1357 5817 1473 5823
rect 3547 5817 3593 5823
rect 3007 5797 3053 5803
rect 4073 5803 4087 5813
rect 5467 5817 5633 5823
rect 4073 5800 4273 5803
rect 4077 5797 4273 5800
rect 6537 5777 6593 5783
rect 4947 5757 5073 5763
rect 5507 5757 5593 5763
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 7687 5697 7793 5703
rect 2137 5677 2233 5683
rect 6627 5677 6693 5683
rect 2707 5657 2733 5663
rect 777 5637 853 5643
rect 3087 5637 3133 5643
rect 4367 5637 4393 5643
rect 8267 5637 8353 5643
rect 1607 5617 1653 5623
rect 1847 5617 1893 5623
rect 1907 5617 2013 5623
rect 2647 5617 2813 5623
rect 680 5603 693 5607
rect 677 5593 693 5603
rect 3267 5597 3353 5603
rect 3513 5603 3527 5613
rect 4807 5617 5033 5623
rect 6567 5617 6673 5623
rect 6807 5617 7033 5623
rect 8287 5617 8413 5623
rect 8547 5617 8693 5623
rect 10807 5617 10933 5623
rect 10987 5617 11033 5623
rect 11947 5617 12053 5623
rect 3513 5600 3653 5603
rect 3517 5597 3653 5600
rect 4253 5603 4267 5612
rect 4253 5600 4293 5603
rect 4257 5597 4293 5600
rect 677 5567 683 5593
rect 5313 5603 5327 5613
rect 8920 5603 8933 5607
rect 5313 5600 5423 5603
rect 5317 5597 5423 5600
rect 5417 5587 5423 5597
rect 8917 5593 8933 5603
rect 11107 5597 11133 5603
rect 12160 5603 12173 5607
rect 12157 5593 12173 5603
rect 2187 5577 2253 5583
rect 5367 5577 5413 5583
rect 8917 5567 8923 5593
rect 677 5557 693 5567
rect 680 5553 693 5557
rect 2987 5557 3153 5563
rect 3767 5557 3933 5563
rect 8917 5557 8933 5567
rect 8920 5553 8933 5557
rect 12157 5563 12163 5593
rect 12007 5557 12163 5563
rect 2187 5537 2233 5543
rect 2947 5537 3133 5543
rect 4287 5537 4333 5543
rect 11767 5537 11833 5543
rect 3027 5517 3113 5523
rect 11647 5517 11693 5523
rect 3587 5497 3633 5503
rect 12343 5478 12403 5982
rect 12310 5462 12403 5478
rect 4067 5437 4133 5443
rect 6767 5437 6913 5443
rect 4487 5417 4613 5423
rect 5147 5397 5313 5403
rect 8447 5397 8573 5403
rect 11087 5397 11153 5403
rect 3187 5377 3233 5383
rect 3727 5377 3853 5383
rect 10813 5383 10827 5393
rect 10813 5380 10933 5383
rect 10817 5377 10933 5380
rect 2947 5337 3073 5343
rect 6887 5337 6933 5343
rect 7407 5337 7513 5343
rect 8767 5337 8873 5343
rect 4227 5317 4273 5323
rect 7427 5317 7553 5323
rect 10807 5317 10873 5323
rect 12027 5317 12193 5323
rect 1587 5297 1693 5303
rect 3727 5297 3813 5303
rect 7347 5297 7513 5303
rect 10307 5297 10413 5303
rect 1813 5243 1827 5253
rect 1813 5240 1973 5243
rect 1817 5237 1973 5240
rect 4007 5237 4133 5243
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 10967 5177 11053 5183
rect 2027 5137 2173 5143
rect 2687 5137 2793 5143
rect 3507 5137 3533 5143
rect 3467 5117 3493 5123
rect 4207 5117 4313 5123
rect 8587 5097 8653 5103
rect 9807 5097 10033 5103
rect 10447 5097 10553 5103
rect 11507 5097 11653 5103
rect 12027 5097 12253 5103
rect 2873 5083 2887 5093
rect 2873 5080 2903 5083
rect 2877 5077 2903 5080
rect 2897 5047 2903 5077
rect 5237 5077 5373 5083
rect 4967 5057 5123 5063
rect 5117 5047 5123 5057
rect 5237 5047 5243 5077
rect 10967 5077 11113 5083
rect 11787 5083 11800 5087
rect 11787 5073 11803 5083
rect 11797 5047 11803 5073
rect 2887 5037 2903 5047
rect 2887 5033 2900 5037
rect 4967 5037 5093 5043
rect 5117 5037 5133 5047
rect 5120 5033 5133 5037
rect 5227 5037 5243 5047
rect 5227 5033 5240 5037
rect 5267 5037 5373 5043
rect 8247 5037 8373 5043
rect 11307 5037 11413 5043
rect 11787 5037 11803 5047
rect 11787 5033 11800 5037
rect 3107 5017 3333 5023
rect 7487 5017 7553 5023
rect 7967 5017 8073 5023
rect 10467 5017 10593 5023
rect 10947 5017 11013 5023
rect 1347 4977 1433 4983
rect 5607 4977 5633 4983
rect 8747 4977 8793 4983
rect 12343 4958 12403 5462
rect 12310 4942 12403 4958
rect 3227 4917 3253 4923
rect 5427 4917 5533 4923
rect 5927 4917 6053 4923
rect 7207 4917 7293 4923
rect 4947 4877 4973 4883
rect 7067 4877 7113 4883
rect 8367 4877 8453 4883
rect 9507 4877 9593 4883
rect 11367 4877 11453 4883
rect 11507 4877 11613 4883
rect 11667 4877 11693 4883
rect 1807 4857 1893 4863
rect 3407 4863 3420 4867
rect 3407 4853 3423 4863
rect 4527 4857 4613 4863
rect 6187 4857 6333 4863
rect 10387 4857 10413 4863
rect 10667 4857 10693 4863
rect 12097 4860 12133 4863
rect 12093 4857 12133 4860
rect 3417 4823 3423 4853
rect 12093 4847 12107 4857
rect 12106 4840 12107 4847
rect 12113 4827 12127 4833
rect 3417 4817 3573 4823
rect 3687 4817 3793 4823
rect 4247 4817 4393 4823
rect 5427 4817 5533 4823
rect 6187 4817 6253 4823
rect 6727 4817 6793 4823
rect 6807 4817 6833 4823
rect 8087 4817 8193 4823
rect 8857 4820 8973 4823
rect 8853 4817 8973 4820
rect 8853 4807 8867 4817
rect 9147 4817 9253 4823
rect 10847 4817 10993 4823
rect 11167 4817 11273 4823
rect 12113 4820 12133 4827
rect 12117 4817 12133 4820
rect 12120 4813 12133 4817
rect 1567 4797 1613 4803
rect 3667 4797 3773 4803
rect 4247 4797 4413 4803
rect 4587 4797 4693 4803
rect 5107 4797 5273 4803
rect 857 4777 913 4783
rect 3937 4777 4013 4783
rect 11727 4777 11873 4783
rect 3107 4757 3153 4763
rect 3427 4757 3593 4763
rect 3853 4763 3867 4773
rect 3727 4760 3867 4763
rect 3727 4757 3863 4760
rect 5627 4757 5793 4763
rect 1677 4737 1733 4743
rect 4907 4737 5023 4743
rect 5907 4717 6073 4723
rect 8867 4717 8993 4723
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 6637 4637 6673 4643
rect 5627 4617 5733 4623
rect 5887 4617 6073 4623
rect 10367 4617 10413 4623
rect 797 4597 833 4603
rect 5647 4597 5773 4603
rect 3807 4577 3953 4583
rect 4007 4577 4113 4583
rect 4567 4577 4773 4583
rect 5627 4577 5813 4583
rect 6987 4577 7173 4583
rect 8527 4577 8653 4583
rect 9107 4577 9253 4583
rect 10667 4577 10793 4583
rect 11767 4577 11913 4583
rect 2607 4557 2773 4563
rect 11247 4563 11260 4567
rect 11247 4553 11263 4563
rect 11787 4557 11853 4563
rect 11257 4527 11263 4553
rect 1647 4517 1673 4523
rect 2597 4520 2803 4523
rect 2593 4517 2807 4520
rect 2593 4507 2607 4517
rect 2793 4507 2807 4517
rect 4127 4517 4213 4523
rect 5987 4517 6073 4523
rect 10707 4517 10833 4523
rect 11247 4517 11263 4527
rect 11247 4513 11260 4517
rect 2907 4497 3093 4503
rect 3267 4497 3413 4503
rect 5907 4503 5920 4507
rect 5907 4493 5923 4503
rect 6007 4497 6073 4503
rect 4947 4477 4993 4483
rect 5917 4483 5923 4493
rect 9947 4497 10053 4503
rect 5917 4477 6033 4483
rect 9867 4477 9973 4483
rect 9987 4477 10013 4483
rect 2927 4457 3093 4463
rect 4387 4457 4493 4463
rect 11567 4457 11593 4463
rect 12343 4438 12403 4942
rect 12310 4422 12403 4438
rect 1507 4397 1633 4403
rect 6907 4397 7013 4403
rect 7467 4397 7593 4403
rect 6113 4383 6127 4393
rect 6113 4380 6253 4383
rect 6117 4377 6253 4380
rect 11767 4377 11913 4383
rect 2647 4357 2773 4363
rect 2907 4357 3053 4363
rect 3187 4357 3273 4363
rect 5207 4357 5313 4363
rect 5387 4357 5473 4363
rect 8767 4357 8953 4363
rect 9647 4357 9753 4363
rect 1747 4343 1760 4347
rect 1747 4333 1763 4343
rect 2327 4343 2340 4347
rect 2327 4333 2343 4343
rect 2607 4337 2653 4343
rect 5247 4337 5273 4343
rect 1757 4307 1763 4333
rect 2337 4307 2343 4333
rect 1747 4297 1763 4307
rect 1747 4293 1760 4297
rect 2327 4297 2343 4307
rect 2327 4293 2340 4297
rect 3707 4297 3873 4303
rect 3947 4297 4013 4303
rect 5947 4297 5993 4303
rect 6077 4300 6173 4303
rect 6073 4297 6173 4300
rect 6073 4287 6087 4297
rect 6907 4297 7053 4303
rect 12167 4297 12213 4303
rect 1527 4277 1653 4283
rect 2827 4277 2993 4283
rect 4227 4277 4373 4283
rect 5007 4277 5133 4283
rect 5347 4277 5473 4283
rect 7987 4277 8193 4283
rect 11487 4277 11633 4283
rect 1847 4257 1943 4263
rect 2367 4257 2453 4263
rect 6607 4257 6793 4263
rect 3527 4237 3613 4243
rect 4507 4237 4613 4243
rect 1220 4223 1233 4227
rect 1217 4217 1233 4223
rect 1220 4213 1233 4217
rect 6607 4217 6633 4223
rect 10487 4197 10533 4203
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 3007 4137 3053 4143
rect 9257 4140 9433 4143
rect 9253 4137 9433 4140
rect 9253 4127 9267 4137
rect 8447 4117 8593 4123
rect 667 4077 703 4083
rect 4127 4077 4233 4083
rect 9007 4077 9093 4083
rect 10407 4077 10553 4083
rect 2287 4063 2300 4067
rect 2287 4053 2303 4063
rect 2787 4057 2873 4063
rect 3287 4057 3333 4063
rect 6587 4057 6693 4063
rect 8467 4057 8633 4063
rect 2297 4027 2303 4053
rect 8987 4057 9173 4063
rect 2367 4037 2423 4043
rect 2287 4017 2303 4027
rect 2287 4013 2300 4017
rect 2417 3983 2423 4037
rect 6127 4037 6253 4043
rect 9077 4007 9083 4033
rect 6707 3997 6733 4003
rect 6887 3997 7013 4003
rect 8167 3997 8233 4003
rect 9067 3997 9083 4007
rect 9097 4003 9103 4057
rect 9973 4043 9987 4053
rect 9887 4040 9987 4043
rect 9887 4037 9983 4040
rect 9097 3997 9173 4003
rect 9067 3993 9080 3997
rect 9787 3997 9853 4003
rect 2417 3977 2453 3983
rect 3607 3977 3713 3983
rect 9107 3977 9193 3983
rect 1547 3957 1633 3963
rect 4307 3957 4353 3963
rect 4367 3957 4513 3963
rect 4567 3957 4713 3963
rect 7707 3957 7793 3963
rect 2967 3937 3053 3943
rect 6427 3937 6453 3943
rect 6647 3937 6713 3943
rect 12343 3918 12403 4422
rect 12310 3902 12403 3918
rect 6147 3877 6253 3883
rect 7247 3877 7333 3883
rect 5360 3866 5380 3867
rect 5307 3857 5353 3863
rect 5367 3863 5380 3866
rect 10353 3863 10367 3873
rect 5367 3857 5383 3863
rect 10353 3860 10513 3863
rect 10357 3857 10513 3860
rect 5367 3853 5380 3857
rect 4727 3837 4793 3843
rect 5007 3837 5193 3843
rect 8227 3837 8253 3843
rect 8767 3837 8933 3843
rect 2807 3817 2913 3823
rect 4187 3817 4313 3823
rect 4747 3817 4893 3823
rect 4877 3787 4883 3817
rect 6147 3817 6313 3823
rect 6667 3817 6813 3823
rect 9847 3817 9953 3823
rect 4877 3777 4893 3787
rect 4880 3773 4893 3777
rect 5887 3777 5933 3783
rect 8507 3777 8593 3783
rect 3307 3757 3513 3763
rect 4707 3757 4773 3763
rect 5267 3757 5453 3763
rect 5787 3757 5853 3763
rect 6367 3757 6493 3763
rect 10107 3757 10193 3763
rect 10947 3757 11113 3763
rect 11487 3757 11593 3763
rect 5607 3737 5633 3743
rect 5607 3717 5693 3723
rect 9307 3717 9393 3723
rect 9407 3717 9493 3723
rect 10127 3717 10273 3723
rect 11707 3717 11853 3723
rect 6687 3697 6813 3703
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 1867 3623 1880 3627
rect 1867 3617 1883 3623
rect 1867 3613 1880 3617
rect 5167 3617 5203 3623
rect 10427 3617 10553 3623
rect 3407 3597 3433 3603
rect 7807 3597 7853 3603
rect 11787 3577 11813 3583
rect 1127 3537 1273 3543
rect 2467 3537 2693 3543
rect 3287 3537 3413 3543
rect 3587 3537 3653 3543
rect 5807 3537 5933 3543
rect 8527 3537 8593 3543
rect 10407 3537 10493 3543
rect 11887 3537 11953 3543
rect 6387 3517 6513 3523
rect 10007 3517 10033 3523
rect 10147 3523 10160 3527
rect 10147 3513 10163 3523
rect 10967 3517 11033 3523
rect 11667 3517 11693 3523
rect 12220 3523 12233 3527
rect 12217 3513 12233 3523
rect 10157 3487 10163 3513
rect 12217 3487 12223 3513
rect 4207 3477 4313 3483
rect 5827 3477 5893 3483
rect 7447 3477 7493 3483
rect 9367 3477 9493 3483
rect 10147 3477 10163 3487
rect 10147 3473 10160 3477
rect 10787 3477 10833 3483
rect 11487 3477 11613 3483
rect 12217 3477 12233 3487
rect 12220 3473 12233 3477
rect 4247 3457 4273 3463
rect 4427 3457 4653 3463
rect 5867 3457 5953 3463
rect 6867 3457 6953 3463
rect 7687 3457 7833 3463
rect 11347 3457 11413 3463
rect 11887 3457 11933 3463
rect 5547 3437 5633 3443
rect 9027 3437 9153 3443
rect 6987 3417 7033 3423
rect 7967 3417 8113 3423
rect 9367 3417 9393 3423
rect 12343 3398 12403 3902
rect 12310 3382 12403 3398
rect 4967 3357 4993 3363
rect 9527 3357 9573 3363
rect 5247 3317 5373 3323
rect 5467 3317 5513 3323
rect 9567 3297 9693 3303
rect 12067 3303 12080 3307
rect 12067 3293 12083 3303
rect 4187 3257 4273 3263
rect 7647 3257 7793 3263
rect 8507 3257 8653 3263
rect 12077 3263 12083 3293
rect 12057 3257 12083 3263
rect 6847 3237 7033 3243
rect 9747 3237 9893 3243
rect 10167 3237 10253 3243
rect 10667 3237 10813 3243
rect 11187 3237 11273 3243
rect 11747 3237 11773 3243
rect 12057 3243 12063 3257
rect 12007 3237 12063 3243
rect 7727 3217 7873 3223
rect 10067 3217 10133 3223
rect 5487 3197 5653 3203
rect 9887 3197 9933 3203
rect 11807 3197 11853 3203
rect 10907 3157 11093 3163
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 7047 3097 7133 3103
rect 9767 3097 9853 3103
rect 10027 3097 10133 3103
rect 647 3057 673 3063
rect 5213 3063 5227 3073
rect 5213 3060 5353 3063
rect 5217 3057 5353 3060
rect 8927 3057 9013 3063
rect 8607 3037 8693 3043
rect 687 3017 713 3023
rect 2287 3017 2333 3023
rect 4747 3017 4853 3023
rect 7287 3017 7393 3023
rect 8607 3017 8733 3023
rect 10747 3017 10773 3023
rect 11287 3017 11453 3023
rect 11667 3017 11693 3023
rect 4127 2997 4173 3003
rect 5767 2997 5933 3003
rect 11027 2997 11093 3003
rect 11667 2997 11713 3003
rect 6327 2977 6373 2983
rect 4727 2957 4813 2963
rect 6767 2957 6793 2963
rect 10247 2957 10293 2963
rect 11607 2957 11673 2963
rect 4107 2937 4213 2943
rect 4787 2937 4833 2943
rect 9167 2937 9333 2943
rect 11267 2937 11413 2943
rect 11587 2937 11613 2943
rect 3847 2897 3933 2903
rect 6827 2897 6873 2903
rect 12343 2878 12403 3382
rect 12310 2862 12403 2878
rect 307 2837 433 2843
rect 447 2837 473 2843
rect 2727 2817 2793 2823
rect 4887 2817 4973 2823
rect 12107 2817 12193 2823
rect 2107 2797 2253 2803
rect 2707 2797 2873 2803
rect 4267 2797 4353 2803
rect 5607 2797 5793 2803
rect 6147 2797 6173 2803
rect 6407 2797 6493 2803
rect 6927 2797 7013 2803
rect 8847 2797 8913 2803
rect 3467 2777 3613 2783
rect 4547 2777 4613 2783
rect 4907 2777 4993 2783
rect 5387 2777 5493 2783
rect 4567 2757 4633 2763
rect 2167 2737 2313 2743
rect 947 2717 1013 2723
rect 2087 2717 2173 2723
rect 3707 2717 3893 2723
rect 5867 2717 5973 2723
rect 6167 2717 6353 2723
rect 9367 2717 9593 2723
rect 10167 2717 10193 2723
rect 10207 2717 10313 2723
rect 12027 2717 12213 2723
rect 12267 2717 12293 2723
rect 2397 2697 2473 2703
rect 1327 2677 1393 2683
rect 5927 2637 5993 2643
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 4647 2577 4773 2583
rect 1227 2557 1263 2563
rect 4667 2537 4733 2543
rect 907 2497 953 2503
rect 3767 2497 3833 2503
rect 4587 2497 4833 2503
rect 6447 2497 6673 2503
rect 8307 2497 8453 2503
rect 9407 2497 9453 2503
rect 10727 2497 10893 2503
rect 5907 2477 6013 2483
rect 12087 2477 12193 2483
rect 7027 2437 7153 2443
rect 9707 2417 9753 2423
rect 9927 2397 10113 2403
rect 10167 2397 10333 2403
rect 12343 2358 12403 2862
rect 12310 2342 12403 2358
rect 10547 2320 10643 2323
rect 10547 2317 10647 2320
rect 10633 2307 10647 2317
rect 8647 2297 8733 2303
rect 12087 2297 12193 2303
rect 1387 2277 1473 2283
rect 2167 2277 2333 2283
rect 2647 2277 2853 2283
rect 3747 2277 3933 2283
rect 6107 2277 6213 2283
rect 11807 2277 11913 2283
rect 12027 2277 12073 2283
rect 4033 2263 4047 2273
rect 4033 2260 4193 2263
rect 4037 2257 4193 2260
rect 11567 2257 11633 2263
rect 11787 2263 11800 2267
rect 11787 2253 11803 2263
rect 11797 2227 11803 2253
rect 607 2217 773 2223
rect 8347 2217 8373 2223
rect 9147 2217 9293 2223
rect 9927 2217 10033 2223
rect 11787 2217 11803 2227
rect 11787 2213 11800 2217
rect 2667 2197 2773 2203
rect 3987 2197 4113 2203
rect 5607 2197 5773 2203
rect 6547 2197 6633 2203
rect 9167 2197 9193 2203
rect 9407 2197 9593 2203
rect 11507 2197 11633 2203
rect 2937 2177 3073 2183
rect 7387 2177 7413 2183
rect 8867 2177 9073 2183
rect 9387 2177 9553 2183
rect 10747 2177 10793 2183
rect 6987 2157 7053 2163
rect 1667 2143 1680 2147
rect 1667 2137 1683 2143
rect 1667 2133 1680 2137
rect 2307 2137 2343 2143
rect 5647 2117 5713 2123
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 5157 2057 5233 2063
rect 9347 2057 9453 2063
rect 10187 2057 10253 2063
rect 3527 2037 3633 2043
rect 3477 2020 3653 2023
rect 3473 2017 3653 2020
rect 3473 2007 3487 2017
rect 5727 2017 5813 2023
rect 6567 2017 6713 2023
rect 10087 2017 10253 2023
rect 1687 1977 1733 1983
rect 3427 1977 3593 1983
rect 4587 1977 4713 1983
rect 5827 1977 5913 1983
rect 5987 1977 6073 1983
rect 7907 1977 7993 1983
rect 8747 1977 8913 1983
rect 9327 1977 9413 1983
rect 10907 1977 10993 1983
rect 11987 1977 12073 1983
rect 2787 1957 2813 1963
rect 3767 1957 3793 1963
rect 7107 1957 7173 1963
rect 7247 1957 7273 1963
rect 7287 1957 7313 1963
rect 7967 1957 8013 1963
rect 9107 1917 9233 1923
rect 10657 1917 10853 1923
rect 2107 1897 2213 1903
rect 6247 1897 6333 1903
rect 6347 1897 6433 1903
rect 9067 1897 9173 1903
rect 10657 1903 10663 1917
rect 10627 1897 10663 1903
rect 10147 1877 10233 1883
rect 12343 1838 12403 2342
rect 12310 1822 12403 1838
rect 2427 1757 2533 1763
rect 4667 1757 4713 1763
rect 7067 1757 7293 1763
rect 11167 1757 11233 1763
rect 2047 1737 2093 1743
rect 6647 1737 6713 1743
rect 6867 1737 6993 1743
rect 8847 1737 8933 1743
rect 12160 1743 12173 1747
rect 9993 1723 10007 1733
rect 9907 1720 10007 1723
rect 12157 1733 12173 1743
rect 9907 1717 10003 1720
rect 12157 1707 12163 1733
rect 1427 1697 1493 1703
rect 5167 1697 5213 1703
rect 6287 1697 6353 1703
rect 12157 1697 12173 1707
rect 12160 1693 12173 1697
rect 687 1677 733 1683
rect 6267 1677 6473 1683
rect 6527 1677 6573 1683
rect 7087 1677 7113 1683
rect 8767 1677 8933 1683
rect 11387 1677 11613 1683
rect 11947 1677 12233 1683
rect 887 1657 1003 1663
rect 11227 1657 11333 1663
rect 9047 1637 9193 1643
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 7367 1537 7413 1543
rect 9167 1537 9233 1543
rect 3520 1523 3533 1527
rect 3517 1517 3533 1523
rect 3520 1513 3533 1517
rect 887 1477 1063 1483
rect 5027 1477 5083 1483
rect 6847 1477 6873 1483
rect 547 1457 573 1463
rect 1967 1457 2153 1463
rect 6827 1457 6893 1463
rect 7827 1457 7973 1463
rect 11787 1443 11800 1447
rect 11787 1440 11803 1443
rect 11787 1433 11807 1440
rect 11793 1426 11807 1433
rect 4887 1397 4993 1403
rect 4627 1377 4833 1383
rect 7787 1377 7893 1383
rect 7907 1377 7933 1383
rect 10707 1377 10873 1383
rect 11487 1377 11653 1383
rect 1467 1357 1513 1363
rect 12343 1318 12403 1822
rect 12310 1302 12403 1318
rect 387 1277 413 1283
rect 2327 1257 2433 1263
rect 5387 1237 5553 1243
rect 6567 1237 6653 1243
rect 7087 1237 7153 1243
rect 6447 1217 6533 1223
rect 2607 1177 2653 1183
rect 7837 1180 7933 1183
rect 7833 1177 7933 1180
rect 7833 1167 7847 1177
rect 8647 1177 8753 1183
rect 10287 1177 10373 1183
rect 12027 1177 12073 1183
rect 3067 1157 3233 1163
rect 4527 1157 4553 1163
rect 7087 1157 7233 1163
rect 7727 1157 7753 1163
rect 267 1137 393 1143
rect 7647 1137 7773 1143
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 8437 997 8493 1003
rect 10827 957 10893 963
rect 1327 937 1533 943
rect 4747 937 4813 943
rect 5047 937 5273 943
rect 7527 937 7653 943
rect 11507 937 11553 943
rect 3187 877 3273 883
rect 12127 877 12213 883
rect 11247 857 11353 863
rect 12343 798 12403 1302
rect 12310 782 12403 798
rect 8507 757 8573 763
rect 11907 737 12013 743
rect 4387 717 4413 723
rect 6607 717 6793 723
rect 3587 697 3673 703
rect 6467 697 6493 703
rect 11887 697 11913 703
rect 4667 657 4853 663
rect 727 637 753 643
rect 8667 637 8833 643
rect 10847 637 10993 643
rect 2707 617 2913 623
rect 6687 617 6753 623
rect 11987 617 12063 623
rect 10967 577 11013 583
rect -63 522 30 538
rect -63 18 -3 522
rect 480 483 493 487
rect 477 477 493 483
rect 480 473 493 477
rect 5140 483 5153 487
rect 5137 477 5153 483
rect 5140 473 5153 477
rect 11760 483 11773 487
rect 11757 477 11773 483
rect 11760 473 11773 477
rect 2097 437 2213 443
rect 2847 417 2973 423
rect 4427 417 4593 423
rect 5947 417 6033 423
rect 9227 417 9233 423
rect 9247 417 9413 423
rect 12187 417 12213 423
rect 5707 397 5753 403
rect 6087 377 6113 383
rect 727 337 793 343
rect 807 337 913 343
rect 10287 337 10393 343
rect 10407 337 10473 343
rect 11887 337 11913 343
rect 11033 323 11047 333
rect 11033 320 11233 323
rect 11037 317 11233 320
rect 12343 278 12403 782
rect 12310 262 12403 278
rect 1227 197 1293 203
rect 5467 197 5493 203
rect 1257 147 1263 173
rect 1257 137 1273 147
rect 1260 133 1273 137
rect 1247 117 1313 123
rect 4047 117 4113 123
rect 10967 117 11073 123
rect 1267 97 1303 103
rect 4067 57 4123 63
rect 8040 63 8053 67
rect 6327 57 6503 63
rect 8037 57 8053 63
rect 8040 53 8053 57
rect 8297 57 8393 63
rect 10840 63 10853 67
rect 10837 57 10853 63
rect 10840 53 10853 57
rect -63 2 30 18
rect 12343 2 12403 262
<< m2contact >>
rect 2113 12153 2127 12167
rect 2313 12153 2327 12167
rect 8473 12153 8487 12167
rect 8673 12153 8687 12167
rect 3633 12093 3647 12107
rect 3793 12093 3807 12107
rect 11073 12093 11087 12107
rect 473 12073 487 12087
rect 733 12073 747 12087
rect 1573 12073 1587 12087
rect 1773 12073 1787 12087
rect 3573 12073 3587 12087
rect 3753 12073 3767 12087
rect 11013 12073 11027 12087
rect 6713 12053 6727 12067
rect 3353 12013 3367 12027
rect 5173 12013 5187 12027
rect 8453 12013 8467 12027
rect 9389 12013 9403 12027
rect 9497 12013 9511 12027
rect 2233 11953 2247 11967
rect 8373 11953 8387 11967
rect 5193 11913 5207 11927
rect 1953 11853 1967 11867
rect 1993 11853 2007 11867
rect 7593 11853 7607 11867
rect 7713 11853 7727 11867
rect 10553 11853 10567 11867
rect 10753 11853 10767 11867
rect 293 11833 307 11847
rect 333 11833 347 11847
rect 2253 11833 2267 11847
rect 2433 11833 2447 11847
rect 5053 11773 5067 11787
rect 5233 11773 5247 11787
rect 9273 11773 9287 11787
rect 9473 11773 9487 11787
rect 1173 11633 1187 11647
rect 1313 11633 1327 11647
rect 6893 11613 6907 11627
rect 7033 11613 7047 11627
rect 5373 11593 5387 11607
rect 5453 11593 5467 11607
rect 833 11573 847 11587
rect 893 11573 907 11587
rect 2453 11573 2467 11587
rect 2613 11573 2627 11587
rect 513 11553 527 11567
rect 733 11553 747 11567
rect 2493 11553 2507 11567
rect 2673 11553 2687 11567
rect 3433 11553 3447 11567
rect 3493 11553 3507 11567
rect 4733 11553 4747 11567
rect 4833 11553 4847 11567
rect 5833 11553 5847 11567
rect 5873 11553 5887 11567
rect 7673 11553 7687 11567
rect 7733 11553 7747 11567
rect 4393 11513 4407 11527
rect 4453 11513 4467 11527
rect 6191 11513 6205 11527
rect 2473 11493 2487 11507
rect 4433 11493 4447 11507
rect 4673 11493 4687 11507
rect 4773 11493 4787 11507
rect 9933 11493 9947 11507
rect 4353 11473 4367 11487
rect 2773 11433 2787 11447
rect 3133 11433 3147 11447
rect 4193 11413 4207 11427
rect 5093 11393 5107 11407
rect 7693 11393 7707 11407
rect 9253 11393 9267 11407
rect 733 11333 747 11347
rect 833 11333 847 11347
rect 2953 11333 2967 11347
rect 3033 11333 3047 11347
rect 3733 11333 3747 11347
rect 3813 11333 3827 11347
rect 6673 11313 6687 11327
rect 6833 11313 6847 11327
rect 10693 11273 10707 11287
rect 10813 11273 10827 11287
rect 6293 11253 6307 11267
rect 6333 11253 6347 11267
rect 6473 11213 6487 11227
rect 6553 11213 6567 11227
rect 9533 11113 9547 11127
rect 9693 11113 9707 11127
rect 11673 11113 11687 11127
rect 11773 11113 11787 11127
rect 3973 11093 3987 11107
rect 4133 11093 4147 11107
rect 2453 11073 2467 11087
rect 2593 11073 2607 11087
rect 4473 11033 4487 11047
rect 4633 11033 4647 11047
rect 4693 11033 4707 11047
rect 4873 11033 4887 11047
rect 4973 11033 4987 11047
rect 6253 11033 6267 11047
rect 6373 11033 6387 11047
rect 2473 11012 2487 11026
rect 2573 11013 2587 11027
rect 3673 10973 3687 10987
rect 6913 10973 6927 10987
rect 8953 10973 8967 10987
rect 6633 10913 6647 10927
rect 3273 10873 3287 10887
rect 1353 10833 1367 10847
rect 1573 10833 1587 10847
rect 1493 10813 1507 10827
rect 1613 10813 1627 10827
rect 3513 10813 3527 10827
rect 3553 10813 3567 10827
rect 8133 10813 8147 10827
rect 8213 10813 8227 10827
rect 8713 10813 8727 10827
rect 8873 10813 8887 10827
rect 11593 10793 11607 10807
rect 5393 10773 5407 10787
rect 5473 10772 5487 10786
rect 613 10753 627 10767
rect 653 10753 667 10767
rect 9773 10753 9787 10767
rect 9813 10753 9827 10767
rect 11593 10753 11607 10767
rect 10893 10713 10907 10727
rect 11053 10713 11067 10727
rect 11213 10713 11227 10727
rect 11333 10713 11347 10727
rect 4173 10693 4187 10707
rect 4253 10693 4267 10707
rect 4353 10593 4367 10607
rect 4413 10593 4427 10607
rect 4293 10573 4307 10587
rect 4393 10573 4407 10587
rect 4833 10573 4847 10587
rect 4953 10572 4967 10586
rect 5993 10572 6007 10586
rect 6133 10573 6147 10587
rect 4613 10533 4627 10547
rect 4733 10533 4747 10547
rect 4533 10513 4547 10527
rect 4713 10513 4727 10527
rect 4953 10513 4967 10527
rect 5013 10513 5027 10527
rect 8433 10513 8447 10527
rect 8513 10513 8527 10527
rect 11213 10513 11227 10527
rect 11413 10513 11427 10527
rect 11753 10513 11767 10527
rect 11953 10513 11967 10527
rect 1733 10493 1747 10507
rect 2513 10493 2527 10507
rect 2613 10493 2627 10507
rect 4353 10493 4367 10507
rect 7633 10493 7647 10507
rect 7693 10493 7707 10507
rect 10933 10493 10947 10507
rect 11093 10493 11107 10507
rect 2393 10473 2407 10487
rect 2513 10472 2527 10486
rect 11033 10473 11047 10487
rect 11153 10473 11167 10487
rect 5713 10453 5727 10467
rect 5973 10453 5987 10467
rect 7133 10453 7147 10467
rect 3773 10373 3787 10387
rect 3933 10373 3947 10387
rect 3173 10353 3187 10367
rect 4097 10353 4111 10367
rect 4833 10353 4847 10367
rect 4973 10353 4987 10367
rect 3793 10333 3807 10347
rect 3973 10333 3987 10347
rect 4953 10313 4967 10327
rect 813 10293 827 10307
rect 1013 10293 1027 10307
rect 3833 10293 3847 10307
rect 3973 10293 3987 10307
rect 5733 10293 5747 10307
rect 5773 10293 5787 10307
rect 9973 10293 9987 10307
rect 10073 10293 10087 10307
rect 10133 10293 10147 10307
rect 2313 10273 2327 10287
rect 2413 10273 2427 10287
rect 7093 10273 7107 10287
rect 3753 10253 3767 10267
rect 3793 10253 3807 10267
rect 7093 10233 7107 10247
rect 9713 10233 9727 10247
rect 9833 10233 9847 10247
rect 2233 10213 2247 10227
rect 2353 10213 2367 10227
rect 3073 10213 3087 10227
rect 3193 10213 3207 10227
rect 3813 10213 3827 10227
rect 3933 10212 3947 10226
rect 5653 10213 5667 10227
rect 5813 10213 5827 10227
rect 8693 10212 8707 10226
rect 8733 10213 8747 10227
rect 3013 10193 3027 10207
rect 3153 10193 3167 10207
rect 8953 10173 8967 10187
rect 9013 10173 9027 10187
rect 7833 10113 7847 10127
rect 7933 10113 7947 10127
rect 5653 10073 5667 10087
rect 5833 10073 5847 10087
rect 3873 10053 3887 10067
rect 3913 10053 3927 10067
rect 6993 10053 7007 10067
rect 7153 10053 7167 10067
rect 7033 10033 7047 10047
rect 2393 10013 2407 10027
rect 2513 10013 2527 10027
rect 6993 10013 7007 10027
rect 7193 10013 7207 10027
rect 1053 9993 1067 10007
rect 1253 9993 1267 10007
rect 5873 9993 5887 10007
rect 6033 9993 6047 10007
rect 7253 9993 7267 10007
rect 7373 9993 7387 10007
rect 7433 9993 7447 10007
rect 11153 9993 11167 10007
rect 11233 9993 11247 10007
rect 6593 9973 6607 9987
rect 3613 9933 3627 9947
rect 4133 9933 4147 9947
rect 8233 9933 8247 9947
rect 3313 9873 3327 9887
rect 3853 9853 3867 9867
rect 3893 9853 3907 9867
rect 7053 9852 7067 9866
rect 7113 9853 7127 9867
rect 7553 9853 7567 9867
rect 7693 9833 7707 9847
rect 7273 9813 7287 9827
rect 7453 9813 7467 9827
rect 7233 9793 7247 9807
rect 7453 9792 7467 9806
rect 9593 9793 9607 9807
rect 9813 9793 9827 9807
rect 1193 9773 1207 9787
rect 1253 9773 1267 9787
rect 1313 9773 1327 9787
rect 1433 9773 1447 9787
rect 3813 9773 3827 9787
rect 3913 9773 3927 9787
rect 8553 9773 8567 9787
rect 8733 9773 8747 9787
rect 11633 9772 11647 9786
rect 11693 9773 11707 9787
rect 2533 9753 2547 9767
rect 2633 9753 2647 9767
rect 3893 9753 3907 9767
rect 4573 9753 4587 9767
rect 4653 9753 4667 9767
rect 7353 9753 7367 9767
rect 7413 9753 7427 9767
rect 10973 9753 10987 9767
rect 2273 9713 2287 9727
rect 2333 9713 2347 9727
rect 10033 9713 10047 9727
rect 10093 9713 10107 9727
rect 10973 9713 10987 9727
rect 12153 9713 12167 9727
rect 12193 9713 12207 9727
rect 3873 9692 3887 9706
rect 6653 9693 6667 9707
rect 6773 9693 6787 9707
rect 6933 9693 6947 9707
rect 7093 9693 7107 9707
rect 4773 9653 4787 9667
rect 4913 9653 4927 9667
rect 3033 9593 3047 9607
rect 3173 9593 3187 9607
rect 233 9553 247 9567
rect 273 9553 287 9567
rect 10073 9553 10087 9567
rect 10173 9556 10187 9570
rect 2173 9533 2187 9547
rect 2353 9533 2367 9547
rect 7573 9533 7587 9547
rect 7693 9533 7707 9547
rect 9433 9533 9447 9547
rect 9593 9533 9607 9547
rect 8613 9493 8627 9507
rect 8693 9493 8707 9507
rect 473 9473 487 9487
rect 693 9473 707 9487
rect 3033 9473 3047 9487
rect 3093 9472 3107 9486
rect 3733 9473 3747 9487
rect 3913 9473 3927 9487
rect 7233 9473 7247 9487
rect 7473 9473 7487 9487
rect 2773 9453 2787 9467
rect 5973 9453 5987 9467
rect 6153 9453 6167 9467
rect 8473 9453 8487 9467
rect 9773 9453 9787 9467
rect 9833 9453 9847 9467
rect 9933 9453 9947 9467
rect 9993 9453 10007 9467
rect 3133 9433 3147 9447
rect 3193 9433 3207 9447
rect 4073 9413 4087 9427
rect 7673 9393 7687 9407
rect 4813 9353 4827 9367
rect 8293 9353 8307 9367
rect 9353 9353 9367 9367
rect 5113 9333 5127 9347
rect 5253 9333 5267 9347
rect 4293 9313 4307 9327
rect 4413 9292 4427 9306
rect 6733 9293 6747 9307
rect 6893 9293 6907 9307
rect 10913 9293 10927 9307
rect 11013 9293 11027 9307
rect 10953 9273 10967 9287
rect 11133 9273 11147 9287
rect 11233 9273 11247 9287
rect 11313 9273 11327 9287
rect 1673 9253 1687 9267
rect 1753 9252 1767 9266
rect 2153 9253 2167 9267
rect 2333 9253 2347 9267
rect 6953 9253 6967 9267
rect 7173 9253 7187 9267
rect 8773 9253 8787 9267
rect 8913 9253 8927 9267
rect 11773 9253 11787 9267
rect 11833 9253 11847 9267
rect 5093 9233 5107 9247
rect 5133 9233 5147 9247
rect 8913 9232 8927 9246
rect 8993 9233 9007 9247
rect 4593 9193 4607 9207
rect 4733 9193 4747 9207
rect 5613 9193 5627 9207
rect 5753 9193 5767 9207
rect 7053 9193 7067 9207
rect 7113 9193 7127 9207
rect 7153 9193 7167 9207
rect 7233 9193 7247 9207
rect 7373 9193 7387 9207
rect 1873 9173 1887 9187
rect 1933 9173 1947 9187
rect 8573 9173 8587 9187
rect 8733 9173 8747 9187
rect 11253 9173 11267 9187
rect 11353 9173 11367 9187
rect 11433 9173 11447 9187
rect 8553 9153 8567 9167
rect 8693 9153 8707 9167
rect 6113 9073 6127 9087
rect 6213 9073 6227 9087
rect 8633 9033 8647 9047
rect 8813 9032 8827 9046
rect 5113 9013 5127 9027
rect 10793 9013 10807 9027
rect 10893 9013 10907 9027
rect 3793 8993 3807 9007
rect 3813 8973 3827 8987
rect 5113 8973 5127 8987
rect 1053 8953 1067 8967
rect 1233 8953 1247 8967
rect 2353 8953 2367 8967
rect 2453 8953 2467 8967
rect 3073 8953 3087 8967
rect 3133 8953 3147 8967
rect 3733 8953 3747 8967
rect 3773 8953 3787 8967
rect 5373 8953 5387 8967
rect 5533 8953 5547 8967
rect 11333 8953 11347 8967
rect 11453 8953 11467 8967
rect 12153 8952 12167 8966
rect 12193 8953 12207 8967
rect 3713 8933 3727 8947
rect 3833 8933 3847 8947
rect 3753 8913 3767 8927
rect 3393 8893 3407 8907
rect 3513 8893 3527 8907
rect 5233 8913 5247 8927
rect 5273 8913 5287 8927
rect 3093 8873 3107 8887
rect 4093 8833 4107 8847
rect 8173 8833 8187 8847
rect 1993 8813 2007 8827
rect 2053 8813 2067 8827
rect 6113 8813 6127 8827
rect 6253 8813 6267 8827
rect 8573 8813 8587 8827
rect 8673 8813 8687 8827
rect 8713 8813 8727 8827
rect 8813 8813 8827 8827
rect 8953 8813 8967 8827
rect 3773 8773 3787 8787
rect 3993 8773 4007 8787
rect 1413 8733 1427 8747
rect 1573 8732 1587 8746
rect 3393 8733 3407 8747
rect 3433 8736 3447 8750
rect 3773 8733 3787 8747
rect 3893 8733 3907 8747
rect 4833 8733 4847 8747
rect 4953 8733 4967 8747
rect 7493 8733 7507 8747
rect 7613 8733 7627 8747
rect 7973 8733 7987 8747
rect 8053 8733 8067 8747
rect 8833 8733 8847 8747
rect 8893 8732 8907 8746
rect 9193 8733 9207 8747
rect 9293 8733 9307 8747
rect 11073 8733 11087 8747
rect 11193 8733 11207 8747
rect 6213 8713 6227 8727
rect 6293 8713 6307 8727
rect 9893 8713 9907 8727
rect 10013 8713 10027 8727
rect 2493 8693 2507 8707
rect 2533 8693 2547 8707
rect 5153 8692 5167 8706
rect 5253 8693 5267 8707
rect 2693 8673 2707 8687
rect 2873 8673 2887 8687
rect 6173 8673 6187 8687
rect 6293 8673 6307 8687
rect 793 8653 807 8667
rect 1033 8653 1047 8667
rect 2473 8653 2487 8667
rect 2613 8653 2627 8667
rect 6413 8653 6427 8667
rect 6573 8653 6587 8667
rect 4553 8533 4567 8547
rect 4653 8533 4667 8547
rect 3733 8513 3747 8527
rect 3933 8513 3947 8527
rect 6453 8513 6467 8527
rect 6613 8513 6627 8527
rect 10913 8513 10927 8527
rect 11013 8513 11027 8527
rect 11053 8513 11067 8527
rect 12053 8513 12067 8527
rect 12213 8516 12227 8530
rect 12253 8513 12267 8527
rect 12313 8513 12327 8527
rect 333 8493 347 8507
rect 413 8493 427 8507
rect 6953 8453 6967 8467
rect 7093 8453 7107 8467
rect 8253 8453 8267 8467
rect 2773 8433 2787 8447
rect 2973 8433 2987 8447
rect 3873 8433 3887 8447
rect 3953 8433 3967 8447
rect 4493 8433 4507 8447
rect 4613 8433 4627 8447
rect 8453 8433 8467 8447
rect 9593 8433 9607 8447
rect 9733 8433 9747 8447
rect 10353 8433 10367 8447
rect 10593 8433 10607 8447
rect 5893 8373 5907 8387
rect 2373 8353 2387 8367
rect 5293 8353 5307 8367
rect 5453 8353 5467 8367
rect 5873 8353 5887 8367
rect 5933 8353 5947 8367
rect 4933 8313 4947 8327
rect 5233 8313 5247 8327
rect 8073 8273 8087 8287
rect 8417 8273 8431 8287
rect 9413 8273 9427 8287
rect 9493 8272 9507 8286
rect 1713 8233 1727 8247
rect 9433 8233 9447 8247
rect 11513 8233 11527 8247
rect 11553 8233 11567 8247
rect 1093 8213 1107 8227
rect 1133 8216 1147 8230
rect 1373 8213 1387 8227
rect 1493 8213 1507 8227
rect 2253 8213 2267 8227
rect 2433 8213 2447 8227
rect 4193 8213 4207 8227
rect 4253 8216 4267 8230
rect 4733 8213 4747 8227
rect 4833 8213 4847 8227
rect 9773 8213 9787 8227
rect 9893 8213 9907 8227
rect 11453 8213 11467 8227
rect 11493 8213 11507 8227
rect 11633 8213 11647 8227
rect 2413 8193 2427 8207
rect 6813 8193 6827 8207
rect 6933 8193 6947 8207
rect 2413 8153 2427 8167
rect 4333 8153 4347 8167
rect 4373 8153 4387 8167
rect 4893 8153 4907 8167
rect 4933 8153 4947 8167
rect 11573 8133 11587 8147
rect 11693 8133 11707 8147
rect 2253 8093 2267 8107
rect 2333 8093 2347 8107
rect 9153 8093 9167 8107
rect 9233 8093 9247 8107
rect 5513 8033 5527 8047
rect 5613 8033 5627 8047
rect 8613 8033 8627 8047
rect 8653 8033 8667 8047
rect 2113 7993 2127 8007
rect 2253 7993 2267 8007
rect 2933 7993 2947 8007
rect 3053 7993 3067 8007
rect 3673 7993 3687 8007
rect 3833 7993 3847 8007
rect 6773 7993 6787 8007
rect 6853 7993 6867 8007
rect 8293 7993 8307 8007
rect 8373 7996 8387 8010
rect 2233 7973 2247 7987
rect 2273 7973 2287 7987
rect 7093 7973 7107 7987
rect 7253 7973 7267 7987
rect 8973 7973 8987 7987
rect 10493 7973 10507 7987
rect 10613 7973 10627 7987
rect 11313 7973 11327 7987
rect 11473 7973 11487 7987
rect 11553 7973 11567 7987
rect 11693 7973 11707 7987
rect 2113 7933 2127 7947
rect 2273 7933 2287 7947
rect 8973 7933 8987 7947
rect 2093 7913 2107 7927
rect 2253 7913 2267 7927
rect 3333 7913 3347 7927
rect 3493 7913 3507 7927
rect 3573 7913 3587 7927
rect 2133 7893 2147 7907
rect 2233 7893 2247 7907
rect 2273 7893 2287 7907
rect 5453 7893 5467 7907
rect 5593 7893 5607 7907
rect 10373 7893 10387 7907
rect 10253 7853 10267 7867
rect 6753 7793 6767 7807
rect 8053 7793 8067 7807
rect 10433 7793 10447 7807
rect 4753 7773 4767 7787
rect 4813 7773 4827 7787
rect 5413 7753 5427 7767
rect 9653 7753 9667 7767
rect 6053 7713 6067 7727
rect 5653 7693 5667 7707
rect 5853 7693 5867 7707
rect 853 7673 867 7687
rect 1013 7673 1027 7687
rect 2993 7673 3007 7687
rect 3093 7673 3107 7687
rect 9373 7673 9387 7687
rect 9513 7673 9527 7687
rect 5693 7633 5707 7647
rect 5873 7633 5887 7647
rect 7293 7633 7307 7647
rect 7393 7633 7407 7647
rect 353 7613 367 7627
rect 493 7613 507 7627
rect 5673 7609 5687 7623
rect 5713 7613 5727 7627
rect 7033 7573 7047 7587
rect 7193 7573 7207 7587
rect 7193 7513 7207 7527
rect 7293 7513 7307 7527
rect 11093 7493 11107 7507
rect 11233 7493 11247 7507
rect 6413 7473 6427 7487
rect 6533 7473 6547 7487
rect 7353 7473 7367 7487
rect 7573 7473 7587 7487
rect 2773 7453 2787 7467
rect 3593 7453 3607 7467
rect 3713 7453 3727 7467
rect 10673 7453 10687 7467
rect 12073 7453 12087 7467
rect 12113 7453 12127 7467
rect 7113 7433 7127 7447
rect 7293 7433 7307 7447
rect 7433 7433 7447 7447
rect 7573 7433 7587 7447
rect 613 7413 627 7427
rect 713 7413 727 7427
rect 2773 7413 2787 7427
rect 3513 7413 3527 7427
rect 3713 7413 3727 7427
rect 10673 7413 10687 7427
rect 533 7393 547 7407
rect 753 7393 767 7407
rect 1693 7393 1707 7407
rect 1733 7393 1747 7407
rect 3653 7393 3667 7407
rect 3733 7393 3747 7407
rect 6453 7393 6467 7407
rect 6533 7393 6547 7407
rect 7433 7393 7447 7407
rect 7533 7393 7547 7407
rect 9793 7393 9807 7407
rect 9933 7393 9947 7407
rect 6113 7373 6127 7387
rect 6213 7373 6227 7387
rect 1933 7353 1947 7367
rect 2033 7353 2047 7367
rect 7413 7353 7427 7367
rect 7593 7353 7607 7367
rect 7853 7273 7867 7287
rect 5673 7253 5687 7267
rect 5813 7253 5827 7267
rect 6773 7253 6787 7267
rect 6873 7253 6887 7267
rect 7073 7253 7087 7267
rect 7233 7253 7247 7267
rect 9933 7233 9947 7247
rect 3833 7213 3847 7227
rect 3933 7213 3947 7227
rect 5393 7213 5407 7227
rect 5593 7213 5607 7227
rect 4613 7193 4627 7207
rect 5293 7193 5307 7207
rect 1773 7173 1787 7187
rect 1833 7173 1847 7187
rect 4813 7173 4827 7187
rect 4993 7173 5007 7187
rect 7213 7173 7227 7187
rect 7273 7173 7287 7187
rect 8253 7173 8267 7187
rect 8293 7173 8307 7187
rect 4393 7153 4407 7167
rect 4453 7153 4467 7167
rect 4833 7153 4847 7167
rect 4893 7153 4907 7167
rect 5413 7153 5427 7167
rect 5573 7153 5587 7167
rect 293 7113 307 7127
rect 433 7113 447 7127
rect 3313 7113 3327 7127
rect 3393 7113 3407 7127
rect 3493 7113 3507 7127
rect 3613 7113 3627 7127
rect 4913 7113 4927 7127
rect 5033 7113 5047 7127
rect 893 7092 907 7106
rect 933 7093 947 7107
rect 3713 7093 3727 7107
rect 3893 7093 3907 7107
rect 4833 7093 4847 7107
rect 4933 7093 4947 7107
rect 5493 7093 5507 7107
rect 5533 7092 5547 7106
rect 7873 7093 7887 7107
rect 7993 7093 8007 7107
rect 8173 7093 8187 7107
rect 8293 7093 8307 7107
rect 9973 7093 9987 7107
rect 10113 7093 10127 7107
rect 10413 7093 10427 7107
rect 10533 7093 10547 7107
rect 10613 7093 10627 7107
rect 11773 7093 11787 7107
rect 12053 7093 12067 7107
rect 5473 7073 5487 7087
rect 5613 7073 5627 7087
rect 7133 7073 7147 7087
rect 7233 7072 7247 7086
rect 11053 6973 11067 6987
rect 11093 6973 11107 6987
rect 833 6953 847 6967
rect 953 6953 967 6967
rect 10593 6953 10607 6967
rect 10753 6956 10767 6970
rect 11773 6953 11787 6967
rect 11833 6956 11847 6970
rect 11873 6956 11887 6970
rect 11913 6953 11927 6967
rect 3613 6933 3627 6947
rect 3713 6933 3727 6947
rect 6733 6933 6747 6947
rect 6893 6933 6907 6947
rect 8373 6912 8387 6926
rect 8473 6913 8487 6927
rect 6193 6893 6207 6907
rect 6233 6893 6247 6907
rect 9473 6893 9487 6907
rect 9553 6893 9567 6907
rect 1953 6873 1967 6887
rect 2013 6873 2027 6887
rect 4053 6873 4067 6887
rect 4113 6873 4127 6887
rect 5953 6873 5967 6887
rect 6033 6873 6047 6887
rect 6993 6873 7007 6887
rect 7213 6873 7227 6887
rect 7473 6872 7487 6886
rect 7513 6873 7527 6887
rect 1973 6853 1987 6867
rect 7353 6853 7367 6867
rect 7513 6852 7527 6866
rect 11893 6833 11907 6847
rect 12073 6833 12087 6847
rect 8113 6813 8127 6827
rect 9253 6733 9267 6747
rect 9133 6713 9147 6727
rect 4153 6693 4167 6707
rect 4193 6693 4207 6707
rect 10193 6693 10207 6707
rect 10253 6693 10267 6707
rect 10293 6693 10307 6707
rect 1533 6673 1547 6687
rect 9373 6673 9387 6687
rect 2713 6653 2727 6667
rect 2793 6653 2807 6667
rect 4333 6653 4347 6667
rect 4533 6653 4547 6667
rect 5573 6653 5587 6667
rect 5633 6653 5647 6667
rect 7313 6653 7327 6667
rect 10893 6656 10907 6670
rect 11073 6653 11087 6667
rect 11693 6653 11707 6667
rect 11933 6653 11947 6667
rect 12153 6653 12167 6667
rect 3773 6632 3787 6646
rect 3973 6633 3987 6647
rect 5993 6633 6007 6647
rect 6153 6633 6167 6647
rect 7613 6633 7627 6647
rect 7733 6633 7747 6647
rect 11353 6633 11367 6647
rect 11393 6633 11407 6647
rect 11553 6633 11567 6647
rect 11633 6633 11647 6647
rect 12013 6633 12027 6647
rect 12133 6633 12147 6647
rect 7313 6613 7327 6627
rect 2613 6593 2627 6607
rect 2653 6593 2667 6607
rect 3793 6593 3807 6607
rect 3933 6592 3947 6606
rect 6153 6593 6167 6607
rect 12173 6593 12187 6607
rect 2713 6573 2727 6587
rect 2873 6573 2887 6587
rect 5413 6573 5427 6587
rect 5573 6573 5587 6587
rect 6053 6572 6067 6586
rect 6093 6573 6107 6587
rect 7593 6573 7607 6587
rect 7713 6573 7727 6587
rect 1173 6553 1187 6567
rect 1293 6553 1307 6567
rect 4133 6553 4147 6567
rect 4273 6553 4287 6567
rect 5453 6532 5467 6546
rect 5573 6533 5587 6547
rect 7353 6473 7367 6487
rect 7473 6473 7487 6487
rect 9513 6453 9527 6467
rect 9613 6453 9627 6467
rect 913 6433 927 6447
rect 1013 6433 1027 6447
rect 2273 6433 2287 6447
rect 2313 6433 2327 6447
rect 2553 6433 2567 6447
rect 2593 6433 2607 6447
rect 10853 6433 10867 6447
rect 11073 6433 11087 6447
rect 11193 6433 11207 6447
rect 11233 6433 11247 6447
rect 11313 6433 11327 6447
rect 11373 6437 11387 6451
rect 4573 6413 4587 6427
rect 4613 6413 4627 6427
rect 5993 6413 6007 6427
rect 6033 6413 6047 6427
rect 7913 6413 7927 6427
rect 8033 6413 8047 6427
rect 8133 6413 8147 6427
rect 8293 6413 8307 6427
rect 10053 6413 10067 6427
rect 10233 6413 10247 6427
rect 11773 6413 11787 6427
rect 11893 6413 11907 6427
rect 12113 6413 12127 6427
rect 12253 6413 12267 6427
rect 4713 6393 4727 6407
rect 4693 6373 4707 6387
rect 4773 6373 4787 6387
rect 4873 6373 4887 6387
rect 6913 6373 6927 6387
rect 6953 6373 6967 6387
rect 12053 6373 12067 6387
rect 12213 6373 12227 6387
rect 1873 6353 1887 6367
rect 1913 6353 1927 6367
rect 2073 6353 2087 6367
rect 2753 6353 2767 6367
rect 2813 6353 2827 6367
rect 3313 6353 3327 6367
rect 3493 6353 3507 6367
rect 4393 6353 4407 6367
rect 4453 6353 4467 6367
rect 6733 6353 6747 6367
rect 6893 6353 6907 6367
rect 8893 6353 8907 6367
rect 9133 6353 9147 6367
rect 8133 6333 8147 6347
rect 2853 6313 2867 6327
rect 2933 6313 2947 6327
rect 3613 6293 3627 6307
rect 3653 6293 3667 6307
rect 5993 6293 6007 6307
rect 9013 6293 9027 6307
rect 8413 6273 8427 6287
rect 8553 6273 8567 6287
rect 6953 6233 6967 6247
rect 2993 6213 3007 6227
rect 3073 6213 3087 6227
rect 5113 6213 5127 6227
rect 5293 6213 5307 6227
rect 11513 6173 11527 6187
rect 11593 6173 11607 6187
rect 1673 6153 1687 6167
rect 1753 6153 1767 6167
rect 1813 6153 1827 6167
rect 2053 6153 2067 6167
rect 3853 6153 3867 6167
rect 3893 6153 3907 6167
rect 1633 6133 1647 6147
rect 3213 6133 3227 6147
rect 3453 6133 3467 6147
rect 3873 6133 3887 6147
rect 3973 6133 3987 6147
rect 7073 6133 7087 6147
rect 7273 6133 7287 6147
rect 7573 6133 7587 6147
rect 7653 6133 7667 6147
rect 10173 6133 10187 6147
rect 10233 6133 10247 6147
rect 10933 6133 10947 6147
rect 11053 6133 11067 6147
rect 11513 6133 11527 6147
rect 11653 6133 11667 6147
rect 1753 6113 1767 6127
rect 3793 6113 3807 6127
rect 3893 6113 3907 6127
rect 4293 6113 4307 6127
rect 4353 6113 4367 6127
rect 11193 6113 11207 6127
rect 11433 6113 11447 6127
rect 11533 6113 11547 6127
rect 11573 6113 11587 6127
rect 11613 6113 11627 6127
rect 3893 6073 3907 6087
rect 3973 6073 3987 6087
rect 4393 6073 4407 6087
rect 4473 6073 4487 6087
rect 7313 6073 7327 6087
rect 7393 6073 7407 6087
rect 11333 6073 11347 6087
rect 1993 6053 2007 6067
rect 2033 6053 2047 6067
rect 2373 6053 2387 6067
rect 2433 6053 2447 6067
rect 2933 6053 2947 6067
rect 3013 6053 3027 6067
rect 4933 6053 4947 6067
rect 5053 6053 5067 6067
rect 5093 6053 5107 6067
rect 5173 6053 5187 6067
rect 5993 6053 6007 6067
rect 6153 6053 6167 6067
rect 6573 6053 6587 6067
rect 6753 6053 6767 6067
rect 8633 6053 8647 6067
rect 8813 6053 8827 6067
rect 12113 6052 12127 6066
rect 12173 6053 12187 6067
rect 3553 6033 3567 6047
rect 4873 6033 4887 6047
rect 4953 6033 4967 6047
rect 10373 6033 10387 6047
rect 3513 6013 3527 6027
rect 10513 6032 10527 6046
rect 3813 6012 3827 6026
rect 3933 6013 3947 6027
rect 5673 6013 5687 6027
rect 5753 6013 5767 6027
rect 1413 5953 1427 5967
rect 1533 5953 1547 5967
rect 3253 5913 3267 5927
rect 3433 5913 3447 5927
rect 4093 5913 4107 5927
rect 4273 5913 4287 5927
rect 4413 5913 4427 5927
rect 4573 5913 4587 5927
rect 5733 5913 5747 5927
rect 5933 5913 5947 5927
rect 3293 5893 3307 5907
rect 3413 5893 3427 5907
rect 3833 5893 3847 5907
rect 3933 5893 3947 5907
rect 4433 5893 4447 5907
rect 4533 5893 4547 5907
rect 7133 5893 7147 5907
rect 7253 5893 7267 5907
rect 10173 5892 10187 5906
rect 10233 5893 10247 5907
rect 11213 5893 11227 5907
rect 11373 5893 11387 5907
rect 4953 5873 4967 5887
rect 4133 5852 4147 5866
rect 4213 5853 4227 5867
rect 4913 5853 4927 5867
rect 4973 5853 4987 5867
rect 5093 5853 5107 5867
rect 573 5833 587 5847
rect 733 5833 747 5847
rect 4153 5833 4167 5847
rect 4293 5833 4307 5847
rect 5453 5833 5467 5847
rect 5693 5833 5707 5847
rect 5733 5833 5747 5847
rect 5773 5833 5787 5847
rect 7733 5833 7747 5847
rect 7853 5833 7867 5847
rect 8693 5833 8707 5847
rect 8893 5833 8907 5847
rect 11573 5833 11587 5847
rect 11713 5833 11727 5847
rect 1473 5813 1487 5827
rect 3533 5813 3547 5827
rect 3593 5813 3607 5827
rect 4073 5813 4087 5827
rect 2993 5793 3007 5807
rect 3053 5793 3067 5807
rect 5453 5812 5467 5826
rect 5633 5813 5647 5827
rect 4273 5793 4287 5807
rect 6593 5773 6607 5787
rect 4933 5753 4947 5767
rect 5073 5753 5087 5767
rect 5493 5752 5507 5766
rect 5593 5753 5607 5767
rect 9473 5733 9487 5747
rect 7673 5693 7687 5707
rect 7793 5693 7807 5707
rect 2233 5673 2247 5687
rect 6613 5673 6627 5687
rect 6693 5672 6707 5686
rect 2693 5653 2707 5667
rect 2733 5653 2747 5667
rect 853 5633 867 5647
rect 3073 5633 3087 5647
rect 3133 5633 3147 5647
rect 4353 5633 4367 5647
rect 4393 5633 4407 5647
rect 8253 5633 8267 5647
rect 8353 5633 8367 5647
rect 1593 5613 1607 5627
rect 1653 5613 1667 5627
rect 1833 5613 1847 5627
rect 1893 5613 1907 5627
rect 2013 5613 2027 5627
rect 2633 5613 2647 5627
rect 2813 5613 2827 5627
rect 3513 5613 3527 5627
rect 693 5593 707 5607
rect 3253 5593 3267 5607
rect 3353 5593 3367 5607
rect 4253 5612 4267 5626
rect 4793 5613 4807 5627
rect 5033 5613 5047 5627
rect 5313 5613 5327 5627
rect 6553 5613 6567 5627
rect 6673 5613 6687 5627
rect 6793 5613 6807 5627
rect 7033 5613 7047 5627
rect 8273 5613 8287 5627
rect 8413 5613 8427 5627
rect 8533 5613 8547 5627
rect 8693 5613 8707 5627
rect 10793 5613 10807 5627
rect 10933 5613 10947 5627
rect 10973 5613 10987 5627
rect 11033 5613 11047 5627
rect 11933 5613 11947 5627
rect 12053 5613 12067 5627
rect 3653 5593 3667 5607
rect 4293 5592 4307 5606
rect 8933 5593 8947 5607
rect 11093 5593 11107 5607
rect 11133 5593 11147 5607
rect 12173 5593 12187 5607
rect 2173 5573 2187 5587
rect 2253 5573 2267 5587
rect 5353 5572 5367 5586
rect 5413 5573 5427 5587
rect 693 5553 707 5567
rect 2973 5553 2987 5567
rect 3153 5553 3167 5567
rect 3753 5553 3767 5567
rect 3933 5553 3947 5567
rect 8933 5553 8947 5567
rect 11993 5553 12007 5567
rect 2173 5533 2187 5547
rect 2233 5533 2247 5547
rect 2933 5533 2947 5547
rect 3133 5533 3147 5547
rect 4273 5532 4287 5546
rect 4333 5533 4347 5547
rect 11753 5533 11767 5547
rect 11833 5533 11847 5547
rect 3013 5513 3027 5527
rect 3113 5512 3127 5526
rect 11633 5513 11647 5527
rect 11693 5513 11707 5527
rect 3573 5493 3587 5507
rect 3633 5492 3647 5506
rect 4053 5432 4067 5446
rect 4133 5433 4147 5447
rect 6753 5433 6767 5447
rect 6913 5433 6927 5447
rect 4473 5413 4487 5427
rect 4613 5413 4627 5427
rect 5133 5393 5147 5407
rect 5313 5393 5327 5407
rect 8433 5393 8447 5407
rect 8573 5393 8587 5407
rect 10813 5393 10827 5407
rect 11073 5393 11087 5407
rect 11153 5393 11167 5407
rect 3173 5373 3187 5387
rect 3233 5373 3247 5387
rect 3713 5373 3727 5387
rect 3853 5373 3867 5387
rect 10933 5373 10947 5387
rect 2933 5333 2947 5347
rect 3073 5333 3087 5347
rect 6873 5333 6887 5347
rect 6933 5333 6947 5347
rect 7393 5333 7407 5347
rect 7513 5333 7527 5347
rect 8753 5333 8767 5347
rect 8873 5333 8887 5347
rect 4213 5313 4227 5327
rect 4273 5313 4287 5327
rect 7413 5313 7427 5327
rect 7553 5313 7567 5327
rect 10793 5313 10807 5327
rect 10873 5313 10887 5327
rect 12013 5313 12027 5327
rect 12193 5313 12207 5327
rect 1573 5293 1587 5307
rect 1693 5293 1707 5307
rect 3713 5293 3727 5307
rect 3813 5293 3827 5307
rect 7333 5293 7347 5307
rect 7513 5292 7527 5306
rect 10293 5293 10307 5307
rect 10413 5293 10427 5307
rect 1813 5253 1827 5267
rect 1973 5233 1987 5247
rect 3993 5233 4007 5247
rect 4133 5233 4147 5247
rect 10953 5173 10967 5187
rect 11053 5173 11067 5187
rect 2013 5133 2027 5147
rect 2173 5133 2187 5147
rect 2673 5133 2687 5147
rect 2793 5133 2807 5147
rect 3493 5133 3507 5147
rect 3533 5132 3547 5146
rect 3453 5113 3467 5127
rect 3493 5112 3507 5126
rect 4193 5113 4207 5127
rect 4313 5113 4327 5127
rect 5773 5113 5787 5127
rect 2873 5093 2887 5107
rect 8573 5093 8587 5107
rect 8653 5093 8667 5107
rect 9793 5093 9807 5107
rect 10033 5093 10047 5107
rect 10433 5093 10447 5107
rect 10553 5093 10567 5107
rect 11493 5096 11507 5110
rect 11653 5093 11667 5107
rect 12013 5093 12027 5107
rect 12253 5093 12267 5107
rect 4953 5053 4967 5067
rect 5373 5073 5387 5087
rect 10953 5073 10967 5087
rect 11113 5073 11127 5087
rect 11773 5073 11787 5087
rect 2873 5033 2887 5047
rect 4953 5032 4967 5046
rect 5093 5033 5107 5047
rect 5133 5033 5147 5047
rect 5213 5033 5227 5047
rect 5253 5033 5267 5047
rect 5373 5033 5387 5047
rect 8233 5033 8247 5047
rect 8373 5033 8387 5047
rect 11293 5033 11307 5047
rect 11413 5033 11427 5047
rect 11773 5033 11787 5047
rect 3093 5013 3107 5027
rect 3333 5013 3347 5027
rect 7473 5013 7487 5027
rect 7553 5009 7567 5023
rect 7953 5013 7967 5027
rect 8073 5012 8087 5026
rect 10453 5013 10467 5027
rect 10593 5013 10607 5027
rect 10933 5013 10947 5027
rect 11013 5013 11027 5027
rect 1333 4973 1347 4987
rect 1433 4972 1447 4986
rect 5593 4973 5607 4987
rect 5633 4973 5647 4987
rect 8733 4973 8747 4987
rect 8793 4973 8807 4987
rect 3213 4913 3227 4927
rect 3253 4912 3267 4926
rect 5413 4913 5427 4927
rect 5533 4913 5547 4927
rect 5913 4913 5927 4927
rect 6053 4913 6067 4927
rect 7193 4913 7207 4927
rect 7293 4913 7307 4927
rect 4933 4873 4947 4887
rect 4973 4873 4987 4887
rect 7053 4872 7067 4886
rect 7113 4873 7127 4887
rect 8353 4873 8367 4887
rect 8453 4873 8467 4887
rect 9493 4873 9507 4887
rect 9593 4873 9607 4887
rect 11353 4873 11367 4887
rect 11453 4873 11467 4887
rect 11493 4873 11507 4887
rect 11613 4873 11627 4887
rect 11653 4876 11667 4890
rect 11693 4873 11707 4887
rect 1793 4853 1807 4867
rect 1893 4853 1907 4867
rect 3393 4853 3407 4867
rect 4513 4853 4527 4867
rect 4613 4853 4627 4867
rect 6173 4853 6187 4867
rect 6333 4853 6347 4867
rect 10373 4853 10387 4867
rect 10413 4853 10427 4867
rect 10653 4853 10667 4867
rect 10693 4853 10707 4867
rect 12133 4853 12147 4867
rect 12092 4833 12106 4847
rect 12113 4833 12127 4847
rect 3573 4813 3587 4827
rect 3673 4813 3687 4827
rect 3793 4813 3807 4827
rect 4233 4813 4247 4827
rect 4393 4813 4407 4827
rect 5413 4813 5427 4827
rect 5533 4813 5547 4827
rect 6173 4813 6187 4827
rect 6253 4813 6267 4827
rect 6713 4813 6727 4827
rect 6793 4813 6807 4827
rect 6833 4813 6847 4827
rect 8073 4813 8087 4827
rect 8193 4813 8207 4827
rect 8973 4813 8987 4827
rect 9133 4813 9147 4827
rect 9253 4813 9267 4827
rect 10833 4813 10847 4827
rect 10993 4813 11007 4827
rect 11153 4813 11167 4827
rect 11273 4813 11287 4827
rect 12133 4813 12147 4827
rect 1553 4793 1567 4807
rect 1613 4793 1627 4807
rect 3653 4793 3667 4807
rect 3773 4793 3787 4807
rect 4233 4792 4247 4806
rect 4413 4792 4427 4806
rect 4573 4793 4587 4807
rect 4693 4793 4707 4807
rect 5093 4793 5107 4807
rect 5273 4793 5287 4807
rect 8853 4793 8867 4807
rect 913 4773 927 4787
rect 3853 4773 3867 4787
rect 4013 4773 4027 4787
rect 11713 4773 11727 4787
rect 3093 4753 3107 4767
rect 3153 4753 3167 4767
rect 3413 4753 3427 4767
rect 3593 4753 3607 4767
rect 3713 4753 3727 4767
rect 11873 4772 11887 4786
rect 5613 4752 5627 4766
rect 5793 4753 5807 4767
rect 1733 4733 1747 4747
rect 4893 4733 4907 4747
rect 5893 4713 5907 4727
rect 6073 4713 6087 4727
rect 8853 4713 8867 4727
rect 8993 4713 9007 4727
rect 6673 4633 6687 4647
rect 5613 4613 5627 4627
rect 5733 4613 5747 4627
rect 5873 4613 5887 4627
rect 6073 4613 6087 4627
rect 10353 4613 10367 4627
rect 10413 4613 10427 4627
rect 833 4593 847 4607
rect 5633 4593 5647 4607
rect 5773 4593 5787 4607
rect 3793 4573 3807 4587
rect 3953 4573 3967 4587
rect 3993 4573 4007 4587
rect 4113 4573 4127 4587
rect 4553 4573 4567 4587
rect 4773 4573 4787 4587
rect 5613 4573 5627 4587
rect 5813 4573 5827 4587
rect 6973 4573 6987 4587
rect 7173 4573 7187 4587
rect 8513 4573 8527 4587
rect 8653 4573 8667 4587
rect 9093 4573 9107 4587
rect 9253 4573 9267 4587
rect 10653 4573 10667 4587
rect 10793 4573 10807 4587
rect 11753 4573 11767 4587
rect 11913 4572 11927 4586
rect 2593 4553 2607 4567
rect 2773 4553 2787 4567
rect 11233 4553 11247 4567
rect 11773 4553 11787 4567
rect 11853 4553 11867 4567
rect 1633 4512 1647 4526
rect 1673 4513 1687 4527
rect 2593 4493 2607 4507
rect 4113 4513 4127 4527
rect 4213 4513 4227 4527
rect 5973 4513 5987 4527
rect 6073 4513 6087 4527
rect 10693 4513 10707 4527
rect 10833 4513 10847 4527
rect 11233 4513 11247 4527
rect 2793 4493 2807 4507
rect 2893 4493 2907 4507
rect 3093 4493 3107 4507
rect 3253 4493 3267 4507
rect 3413 4493 3427 4507
rect 5893 4493 5907 4507
rect 5993 4493 6007 4507
rect 4933 4473 4947 4487
rect 4993 4473 5007 4487
rect 6073 4492 6087 4506
rect 9933 4493 9947 4507
rect 10053 4493 10067 4507
rect 6033 4472 6047 4486
rect 9853 4473 9867 4487
rect 9973 4473 9987 4487
rect 10013 4473 10027 4487
rect 2913 4453 2927 4467
rect 3093 4453 3107 4467
rect 4373 4453 4387 4467
rect 4493 4453 4507 4467
rect 11553 4453 11567 4467
rect 11593 4453 11607 4467
rect 1493 4393 1507 4407
rect 1633 4393 1647 4407
rect 6113 4393 6127 4407
rect 6893 4393 6907 4407
rect 7013 4393 7027 4407
rect 7453 4393 7467 4407
rect 7593 4393 7607 4407
rect 6253 4373 6267 4387
rect 11753 4372 11767 4386
rect 11913 4373 11927 4387
rect 2633 4353 2647 4367
rect 2773 4353 2787 4367
rect 2893 4353 2907 4367
rect 3053 4353 3067 4367
rect 3173 4353 3187 4367
rect 3273 4353 3287 4367
rect 5193 4353 5207 4367
rect 5313 4352 5327 4366
rect 5373 4353 5387 4367
rect 5473 4353 5487 4367
rect 8753 4353 8767 4367
rect 8953 4353 8967 4367
rect 9633 4353 9647 4367
rect 9753 4353 9767 4367
rect 1733 4333 1747 4347
rect 2313 4333 2327 4347
rect 2593 4333 2607 4347
rect 2653 4333 2667 4347
rect 5233 4333 5247 4347
rect 5273 4333 5287 4347
rect 1733 4293 1747 4307
rect 2313 4293 2327 4307
rect 3693 4293 3707 4307
rect 3873 4293 3887 4307
rect 3933 4293 3947 4307
rect 4013 4293 4027 4307
rect 5933 4293 5947 4307
rect 5993 4293 6007 4307
rect 6173 4293 6187 4307
rect 6893 4293 6907 4307
rect 7053 4293 7067 4307
rect 12153 4293 12167 4307
rect 12213 4293 12227 4307
rect 1513 4273 1527 4287
rect 1653 4273 1667 4287
rect 2813 4273 2827 4287
rect 2993 4273 3007 4287
rect 4213 4273 4227 4287
rect 4373 4273 4387 4287
rect 4993 4273 5007 4287
rect 5133 4273 5147 4287
rect 5333 4273 5347 4287
rect 5473 4273 5487 4287
rect 6073 4273 6087 4287
rect 7973 4273 7987 4287
rect 8193 4273 8207 4287
rect 11473 4273 11487 4287
rect 11633 4273 11647 4287
rect 1833 4253 1847 4267
rect 2353 4252 2367 4266
rect 2453 4253 2467 4267
rect 6593 4253 6607 4267
rect 6793 4253 6807 4267
rect 3513 4232 3527 4246
rect 3613 4233 3627 4247
rect 4493 4233 4507 4247
rect 4613 4233 4627 4247
rect 1233 4213 1247 4227
rect 6593 4213 6607 4227
rect 6633 4213 6647 4227
rect 10473 4192 10487 4206
rect 10533 4193 10547 4207
rect 2993 4133 3007 4147
rect 3053 4133 3067 4147
rect 9433 4133 9447 4147
rect 8433 4113 8447 4127
rect 8593 4112 8607 4126
rect 9253 4113 9267 4127
rect 653 4073 667 4087
rect 4113 4073 4127 4087
rect 4233 4073 4247 4087
rect 8993 4073 9007 4087
rect 9093 4073 9107 4087
rect 10393 4073 10407 4087
rect 10553 4073 10567 4087
rect 2273 4053 2287 4067
rect 2773 4053 2787 4067
rect 2873 4053 2887 4067
rect 3273 4053 3287 4067
rect 3333 4053 3347 4067
rect 6573 4053 6587 4067
rect 6693 4053 6707 4067
rect 8453 4053 8467 4067
rect 8633 4053 8647 4067
rect 8973 4052 8987 4066
rect 2353 4033 2367 4047
rect 2273 4013 2287 4027
rect 6113 4033 6127 4047
rect 6253 4033 6267 4047
rect 9073 4033 9087 4047
rect 6693 3993 6707 4007
rect 6733 3993 6747 4007
rect 6873 3993 6887 4007
rect 7013 3993 7027 4007
rect 8153 3993 8167 4007
rect 8233 3993 8247 4007
rect 9053 3993 9067 4007
rect 9173 4053 9187 4067
rect 9973 4053 9987 4067
rect 9873 4033 9887 4047
rect 9173 3993 9187 4007
rect 9773 3993 9787 4007
rect 9853 3993 9867 4007
rect 2453 3973 2467 3987
rect 3593 3973 3607 3987
rect 3713 3973 3727 3987
rect 9093 3973 9107 3987
rect 9193 3969 9207 3983
rect 1533 3952 1547 3966
rect 1633 3953 1647 3967
rect 4293 3953 4307 3967
rect 4353 3953 4367 3967
rect 4513 3953 4527 3967
rect 4553 3953 4567 3967
rect 4713 3953 4727 3967
rect 7693 3953 7707 3967
rect 7793 3953 7807 3967
rect 2953 3933 2967 3947
rect 3053 3933 3067 3947
rect 6413 3933 6427 3947
rect 6453 3933 6467 3947
rect 6633 3933 6647 3947
rect 6713 3932 6727 3946
rect 6133 3873 6147 3887
rect 6253 3873 6267 3887
rect 7233 3873 7247 3887
rect 7333 3873 7347 3887
rect 10353 3873 10367 3887
rect 5293 3853 5307 3867
rect 5353 3852 5367 3866
rect 10513 3853 10527 3867
rect 4713 3833 4727 3847
rect 4793 3833 4807 3847
rect 4993 3833 5007 3847
rect 5193 3833 5207 3847
rect 8213 3833 8227 3847
rect 8253 3833 8267 3847
rect 8753 3833 8767 3847
rect 8933 3833 8947 3847
rect 2793 3813 2807 3827
rect 2913 3813 2927 3827
rect 4173 3813 4187 3827
rect 4313 3813 4327 3827
rect 4733 3813 4747 3827
rect 4893 3813 4907 3827
rect 6133 3813 6147 3827
rect 6313 3813 6327 3827
rect 6653 3813 6667 3827
rect 6813 3813 6827 3827
rect 9833 3813 9847 3827
rect 9953 3812 9967 3826
rect 4893 3773 4907 3787
rect 5873 3773 5887 3787
rect 5933 3773 5947 3787
rect 8493 3773 8507 3787
rect 8593 3773 8607 3787
rect 3293 3749 3307 3763
rect 3513 3753 3527 3767
rect 4693 3753 4707 3767
rect 4773 3753 4787 3767
rect 5253 3753 5267 3767
rect 5453 3753 5467 3767
rect 5773 3753 5787 3767
rect 5853 3753 5867 3767
rect 6353 3749 6367 3763
rect 6493 3753 6507 3767
rect 10093 3753 10107 3767
rect 10193 3753 10207 3767
rect 10933 3753 10947 3767
rect 11113 3753 11127 3767
rect 11473 3753 11487 3767
rect 11593 3752 11607 3766
rect 5593 3733 5607 3747
rect 5633 3733 5647 3747
rect 5593 3712 5607 3726
rect 5693 3713 5707 3727
rect 9293 3713 9307 3727
rect 9393 3713 9407 3727
rect 9493 3713 9507 3727
rect 10113 3713 10127 3727
rect 10273 3713 10287 3727
rect 11693 3713 11707 3727
rect 11853 3713 11867 3727
rect 969 3693 983 3707
rect 1077 3693 1091 3707
rect 6673 3692 6687 3706
rect 6813 3693 6827 3707
rect 1853 3613 1867 3627
rect 5153 3613 5167 3627
rect 10413 3613 10427 3627
rect 10553 3613 10567 3627
rect 3393 3593 3407 3607
rect 3433 3593 3447 3607
rect 7793 3593 7807 3607
rect 7853 3593 7867 3607
rect 11773 3573 11787 3587
rect 11813 3572 11827 3586
rect 1113 3533 1127 3547
rect 1273 3533 1287 3547
rect 2453 3533 2467 3547
rect 2693 3533 2707 3547
rect 3273 3533 3287 3547
rect 3413 3533 3427 3547
rect 3573 3533 3587 3547
rect 3653 3533 3667 3547
rect 5793 3533 5807 3547
rect 5933 3532 5947 3546
rect 8513 3533 8527 3547
rect 8593 3533 8607 3547
rect 10393 3533 10407 3547
rect 10493 3533 10507 3547
rect 11873 3532 11887 3546
rect 11953 3533 11967 3547
rect 6373 3513 6387 3527
rect 6513 3513 6527 3527
rect 9993 3513 10007 3527
rect 10033 3513 10047 3527
rect 10133 3513 10147 3527
rect 10953 3513 10967 3527
rect 11033 3513 11047 3527
rect 11653 3513 11667 3527
rect 11693 3513 11707 3527
rect 12233 3513 12247 3527
rect 4193 3473 4207 3487
rect 4313 3473 4327 3487
rect 5813 3473 5827 3487
rect 5893 3473 5907 3487
rect 7433 3473 7447 3487
rect 7493 3473 7507 3487
rect 9353 3473 9367 3487
rect 9493 3473 9507 3487
rect 10133 3473 10147 3487
rect 10773 3473 10787 3487
rect 10833 3473 10847 3487
rect 11473 3473 11487 3487
rect 11613 3473 11627 3487
rect 12233 3473 12247 3487
rect 4233 3452 4247 3466
rect 4273 3453 4287 3467
rect 4413 3453 4427 3467
rect 4653 3453 4667 3467
rect 5853 3453 5867 3467
rect 5953 3453 5967 3467
rect 6853 3453 6867 3467
rect 6953 3452 6967 3466
rect 7673 3453 7687 3467
rect 7833 3453 7847 3467
rect 11333 3453 11347 3467
rect 11413 3453 11427 3467
rect 11873 3452 11887 3466
rect 11933 3453 11947 3467
rect 5533 3433 5547 3447
rect 5633 3433 5647 3447
rect 9013 3433 9027 3447
rect 9153 3433 9167 3447
rect 6973 3413 6987 3427
rect 7033 3413 7047 3427
rect 7953 3413 7967 3427
rect 8113 3413 8127 3427
rect 9353 3413 9367 3427
rect 9393 3413 9407 3427
rect 4953 3353 4967 3367
rect 4993 3353 5007 3367
rect 9513 3353 9527 3367
rect 9573 3353 9587 3367
rect 5233 3313 5247 3327
rect 5373 3313 5387 3327
rect 5453 3313 5467 3327
rect 5513 3313 5527 3327
rect 9553 3293 9567 3307
rect 9693 3293 9707 3307
rect 12053 3293 12067 3307
rect 4173 3253 4187 3267
rect 4273 3253 4287 3267
rect 7633 3253 7647 3267
rect 7793 3253 7807 3267
rect 8493 3253 8507 3267
rect 8653 3253 8667 3267
rect 6833 3233 6847 3247
rect 7033 3233 7047 3247
rect 9733 3233 9747 3247
rect 9893 3233 9907 3247
rect 10153 3233 10167 3247
rect 10253 3233 10267 3247
rect 10653 3233 10667 3247
rect 10813 3233 10827 3247
rect 11173 3233 11187 3247
rect 11273 3233 11287 3247
rect 11733 3233 11747 3247
rect 11773 3233 11787 3247
rect 11993 3233 12007 3247
rect 7713 3213 7727 3227
rect 7873 3213 7887 3227
rect 10053 3212 10067 3226
rect 10133 3213 10147 3227
rect 5473 3192 5487 3206
rect 5653 3193 5667 3207
rect 9873 3193 9887 3207
rect 9933 3193 9947 3207
rect 11793 3193 11807 3207
rect 11853 3193 11867 3207
rect 10893 3153 10907 3167
rect 11093 3153 11107 3167
rect 7033 3093 7047 3107
rect 7133 3093 7147 3107
rect 9753 3093 9767 3107
rect 9853 3093 9867 3107
rect 10013 3093 10027 3107
rect 10133 3093 10147 3107
rect 5213 3073 5227 3087
rect 633 3053 647 3067
rect 673 3053 687 3067
rect 5353 3053 5367 3067
rect 8913 3053 8927 3067
rect 9013 3053 9027 3067
rect 8593 3033 8607 3047
rect 8693 3033 8707 3047
rect 673 3013 687 3027
rect 713 3013 727 3027
rect 2273 3013 2287 3027
rect 2333 3013 2347 3027
rect 4733 3013 4747 3027
rect 4853 3013 4867 3027
rect 7273 3013 7287 3027
rect 7393 3013 7407 3027
rect 8593 3012 8607 3026
rect 8733 3013 8747 3027
rect 10733 3013 10747 3027
rect 10773 3013 10787 3027
rect 11273 3013 11287 3027
rect 11453 3013 11467 3027
rect 11653 3013 11667 3027
rect 11693 3013 11707 3027
rect 4113 2993 4127 3007
rect 4173 2993 4187 3007
rect 5753 2992 5767 3006
rect 5933 2993 5947 3007
rect 11013 2993 11027 3007
rect 11093 2993 11107 3007
rect 11653 2992 11667 3006
rect 11713 2993 11727 3007
rect 6313 2973 6327 2987
rect 6373 2973 6387 2987
rect 4713 2953 4727 2967
rect 4813 2953 4827 2967
rect 6753 2953 6767 2967
rect 6793 2953 6807 2967
rect 10233 2953 10247 2967
rect 10293 2953 10307 2967
rect 11593 2953 11607 2967
rect 11673 2953 11687 2967
rect 4093 2933 4107 2947
rect 4213 2933 4227 2947
rect 4773 2933 4787 2947
rect 4833 2933 4847 2947
rect 9153 2933 9167 2947
rect 9333 2933 9347 2947
rect 11253 2933 11267 2947
rect 11413 2933 11427 2947
rect 11573 2933 11587 2947
rect 11613 2933 11627 2947
rect 3833 2893 3847 2907
rect 3933 2893 3947 2907
rect 6813 2893 6827 2907
rect 6873 2893 6887 2907
rect 293 2833 307 2847
rect 433 2833 447 2847
rect 473 2833 487 2847
rect 2713 2813 2727 2827
rect 2793 2813 2807 2827
rect 4873 2813 4887 2827
rect 4973 2813 4987 2827
rect 12093 2812 12107 2826
rect 12193 2813 12207 2827
rect 2093 2793 2107 2807
rect 2253 2793 2267 2807
rect 2693 2793 2707 2807
rect 2873 2793 2887 2807
rect 4253 2793 4267 2807
rect 4353 2793 4367 2807
rect 5593 2793 5607 2807
rect 5793 2793 5807 2807
rect 6133 2793 6147 2807
rect 6173 2793 6187 2807
rect 6393 2793 6407 2807
rect 6493 2793 6507 2807
rect 6913 2796 6927 2810
rect 7013 2793 7027 2807
rect 8833 2793 8847 2807
rect 8913 2793 8927 2807
rect 3453 2773 3467 2787
rect 3613 2773 3627 2787
rect 4533 2773 4547 2787
rect 4613 2773 4627 2787
rect 4893 2773 4907 2787
rect 4993 2773 5007 2787
rect 5373 2773 5387 2787
rect 5493 2773 5507 2787
rect 4553 2753 4567 2767
rect 4633 2753 4647 2767
rect 2153 2733 2167 2747
rect 2313 2733 2327 2747
rect 933 2713 947 2727
rect 1013 2713 1027 2727
rect 2073 2713 2087 2727
rect 2173 2713 2187 2727
rect 3693 2713 3707 2727
rect 3893 2713 3907 2727
rect 5853 2713 5867 2727
rect 5973 2713 5987 2727
rect 6153 2713 6167 2727
rect 6353 2713 6367 2727
rect 9353 2713 9367 2727
rect 9593 2713 9607 2727
rect 10153 2713 10167 2727
rect 10193 2713 10207 2727
rect 10313 2713 10327 2727
rect 12013 2713 12027 2727
rect 12213 2713 12227 2727
rect 12253 2709 12267 2723
rect 12293 2713 12307 2727
rect 2473 2693 2487 2707
rect 1313 2673 1327 2687
rect 1393 2673 1407 2687
rect 3413 2649 3427 2663
rect 5913 2633 5927 2647
rect 5993 2633 6007 2647
rect 4633 2573 4647 2587
rect 4773 2573 4787 2587
rect 1213 2553 1227 2567
rect 1857 2553 1871 2567
rect 4653 2533 4667 2547
rect 4733 2533 4747 2547
rect 893 2493 907 2507
rect 953 2493 967 2507
rect 3753 2493 3767 2507
rect 3833 2493 3847 2507
rect 4573 2492 4587 2506
rect 4833 2493 4847 2507
rect 6433 2493 6447 2507
rect 6673 2493 6687 2507
rect 8293 2493 8307 2507
rect 8453 2493 8467 2507
rect 9393 2493 9407 2507
rect 9453 2493 9467 2507
rect 10713 2493 10727 2507
rect 10893 2493 10907 2507
rect 5893 2473 5907 2487
rect 6013 2473 6027 2487
rect 12073 2473 12087 2487
rect 12193 2473 12207 2487
rect 7013 2433 7027 2447
rect 7153 2433 7167 2447
rect 9693 2412 9707 2426
rect 9753 2413 9767 2427
rect 9913 2393 9927 2407
rect 10113 2393 10127 2407
rect 10153 2393 10167 2407
rect 10333 2393 10347 2407
rect 10533 2313 10547 2327
rect 8633 2293 8647 2307
rect 8733 2293 8747 2307
rect 10633 2293 10647 2307
rect 12073 2293 12087 2307
rect 12193 2293 12207 2307
rect 1373 2273 1387 2287
rect 1473 2273 1487 2287
rect 2153 2273 2167 2287
rect 2333 2273 2347 2287
rect 2633 2272 2647 2286
rect 2853 2273 2867 2287
rect 3733 2273 3747 2287
rect 3933 2273 3947 2287
rect 4033 2273 4047 2287
rect 6093 2273 6107 2287
rect 6213 2273 6227 2287
rect 11793 2273 11807 2287
rect 11913 2273 11927 2287
rect 12013 2276 12027 2290
rect 12073 2272 12087 2286
rect 4193 2253 4207 2267
rect 11553 2253 11567 2267
rect 11633 2253 11647 2267
rect 11773 2253 11787 2267
rect 593 2213 607 2227
rect 773 2213 787 2227
rect 8333 2213 8347 2227
rect 8373 2213 8387 2227
rect 9133 2213 9147 2227
rect 9293 2213 9307 2227
rect 9913 2213 9927 2227
rect 10033 2213 10047 2227
rect 11773 2213 11787 2227
rect 2653 2193 2667 2207
rect 2773 2193 2787 2207
rect 3973 2193 3987 2207
rect 4113 2193 4127 2207
rect 5593 2193 5607 2207
rect 5773 2193 5787 2207
rect 6533 2193 6547 2207
rect 6633 2193 6647 2207
rect 9153 2193 9167 2207
rect 9193 2193 9207 2207
rect 9393 2193 9407 2207
rect 9593 2189 9607 2203
rect 11493 2193 11507 2207
rect 11633 2193 11647 2207
rect 3073 2173 3087 2187
rect 7373 2173 7387 2187
rect 7413 2173 7427 2187
rect 8853 2172 8867 2186
rect 9073 2173 9087 2187
rect 9373 2173 9387 2187
rect 9553 2173 9567 2187
rect 10733 2173 10747 2187
rect 10793 2173 10807 2187
rect 6973 2153 6987 2167
rect 7053 2153 7067 2167
rect 1653 2133 1667 2147
rect 2293 2133 2307 2147
rect 5633 2113 5647 2127
rect 5713 2113 5727 2127
rect 5233 2053 5247 2067
rect 9333 2053 9347 2067
rect 9453 2053 9467 2067
rect 10173 2053 10187 2067
rect 10253 2053 10267 2067
rect 3513 2033 3527 2047
rect 3633 2033 3647 2047
rect 3653 2012 3667 2026
rect 5713 2013 5727 2027
rect 5813 2013 5827 2027
rect 6553 2013 6567 2027
rect 6713 2013 6727 2027
rect 10073 2013 10087 2027
rect 10253 2013 10267 2027
rect 3473 1993 3487 2007
rect 1673 1973 1687 1987
rect 1733 1973 1747 1987
rect 3413 1973 3427 1987
rect 3593 1973 3607 1987
rect 4573 1973 4587 1987
rect 4713 1973 4727 1987
rect 5813 1973 5827 1987
rect 5913 1973 5927 1987
rect 5973 1973 5987 1987
rect 6073 1973 6087 1987
rect 7893 1973 7907 1987
rect 7993 1973 8007 1987
rect 8733 1973 8747 1987
rect 8913 1973 8927 1987
rect 9313 1973 9327 1987
rect 9413 1973 9427 1987
rect 10893 1976 10907 1990
rect 10993 1973 11007 1987
rect 11973 1973 11987 1987
rect 12073 1973 12087 1987
rect 2773 1953 2787 1967
rect 2813 1953 2827 1967
rect 3753 1953 3767 1967
rect 3793 1953 3807 1967
rect 7093 1953 7107 1967
rect 7173 1953 7187 1967
rect 7233 1953 7247 1967
rect 7273 1953 7287 1967
rect 7313 1953 7327 1967
rect 7953 1953 7967 1967
rect 8013 1953 8027 1967
rect 9093 1913 9107 1927
rect 9233 1913 9247 1927
rect 2093 1893 2107 1907
rect 2213 1893 2227 1907
rect 6233 1893 6247 1907
rect 6333 1893 6347 1907
rect 6433 1893 6447 1907
rect 9053 1893 9067 1907
rect 9173 1893 9187 1907
rect 10853 1913 10867 1927
rect 10613 1889 10627 1903
rect 10133 1873 10147 1887
rect 10233 1873 10247 1887
rect 2413 1753 2427 1767
rect 2533 1753 2547 1767
rect 4653 1753 4667 1767
rect 4713 1753 4727 1767
rect 7053 1753 7067 1767
rect 7293 1753 7307 1767
rect 11153 1753 11167 1767
rect 11233 1753 11247 1767
rect 2033 1733 2047 1747
rect 2093 1733 2107 1747
rect 6633 1733 6647 1747
rect 6713 1733 6727 1747
rect 6853 1733 6867 1747
rect 6993 1733 7007 1747
rect 8833 1733 8847 1747
rect 8933 1733 8947 1747
rect 9993 1733 10007 1747
rect 9893 1713 9907 1727
rect 12173 1733 12187 1747
rect 1413 1693 1427 1707
rect 1493 1693 1507 1707
rect 5153 1693 5167 1707
rect 5213 1693 5227 1707
rect 6273 1693 6287 1707
rect 6353 1693 6367 1707
rect 12173 1693 12187 1707
rect 673 1673 687 1687
rect 733 1673 747 1687
rect 6253 1673 6267 1687
rect 6473 1673 6487 1687
rect 6513 1673 6527 1687
rect 6573 1673 6587 1687
rect 7073 1673 7087 1687
rect 7113 1673 7127 1687
rect 8753 1673 8767 1687
rect 8933 1673 8947 1687
rect 11373 1673 11387 1687
rect 11613 1673 11627 1687
rect 11933 1673 11947 1687
rect 12233 1673 12247 1687
rect 873 1653 887 1667
rect 11213 1652 11227 1666
rect 11333 1653 11347 1667
rect 9033 1633 9047 1647
rect 9193 1633 9207 1647
rect 1593 1553 1607 1567
rect 7353 1533 7367 1547
rect 7413 1533 7427 1547
rect 9153 1533 9167 1547
rect 9233 1533 9247 1547
rect 3533 1513 3547 1527
rect 873 1473 887 1487
rect 5013 1473 5027 1487
rect 6833 1473 6847 1487
rect 6873 1473 6887 1487
rect 533 1453 547 1467
rect 573 1453 587 1467
rect 1953 1453 1967 1467
rect 2153 1453 2167 1467
rect 6813 1453 6827 1467
rect 6893 1453 6907 1467
rect 7813 1453 7827 1467
rect 7973 1453 7987 1467
rect 11773 1433 11787 1447
rect 11793 1412 11807 1426
rect 4873 1393 4887 1407
rect 4993 1393 5007 1407
rect 4613 1373 4627 1387
rect 4833 1373 4847 1387
rect 7773 1373 7787 1387
rect 7893 1373 7907 1387
rect 7933 1373 7947 1387
rect 10693 1373 10707 1387
rect 10873 1373 10887 1387
rect 11473 1373 11487 1387
rect 11653 1373 11667 1387
rect 1453 1353 1467 1367
rect 1513 1353 1527 1367
rect 373 1273 387 1287
rect 413 1273 427 1287
rect 2313 1253 2327 1267
rect 2433 1253 2447 1267
rect 5373 1233 5387 1247
rect 5553 1233 5567 1247
rect 6553 1233 6567 1247
rect 6653 1233 6667 1247
rect 7073 1233 7087 1247
rect 7153 1233 7167 1247
rect 6433 1213 6447 1227
rect 6533 1213 6547 1227
rect 2593 1173 2607 1187
rect 2653 1173 2667 1187
rect 7933 1173 7947 1187
rect 8633 1173 8647 1187
rect 8753 1173 8767 1187
rect 10273 1173 10287 1187
rect 10373 1173 10387 1187
rect 12013 1173 12027 1187
rect 12073 1173 12087 1187
rect 3053 1153 3067 1167
rect 3233 1153 3247 1167
rect 4513 1153 4527 1167
rect 4553 1153 4567 1167
rect 7073 1153 7087 1167
rect 7233 1153 7247 1167
rect 7713 1153 7727 1167
rect 7753 1153 7767 1167
rect 7833 1153 7847 1167
rect 253 1133 267 1147
rect 393 1133 407 1147
rect 7633 1133 7647 1147
rect 7773 1133 7787 1147
rect 57 993 71 1007
rect 8493 993 8507 1007
rect 10813 953 10827 967
rect 10893 953 10907 967
rect 1313 933 1327 947
rect 1533 933 1547 947
rect 4733 933 4747 947
rect 4813 933 4827 947
rect 5033 933 5047 947
rect 5273 933 5287 947
rect 7513 933 7527 947
rect 7653 933 7667 947
rect 11493 933 11507 947
rect 11553 933 11567 947
rect 3173 873 3187 887
rect 3273 873 3287 887
rect 12113 873 12127 887
rect 12213 873 12227 887
rect 11233 853 11247 867
rect 11353 853 11367 867
rect 8493 753 8507 767
rect 8573 753 8587 767
rect 11893 733 11907 747
rect 12013 733 12027 747
rect 4373 717 4387 731
rect 4413 713 4427 727
rect 6593 713 6607 727
rect 6793 713 6807 727
rect 3573 693 3587 707
rect 3673 693 3687 707
rect 6453 693 6467 707
rect 6493 693 6507 707
rect 11873 693 11887 707
rect 11913 693 11927 707
rect 4653 653 4667 667
rect 4853 653 4867 667
rect 713 633 727 647
rect 753 633 767 647
rect 8653 633 8667 647
rect 8833 633 8847 647
rect 10833 633 10847 647
rect 10993 633 11007 647
rect 2693 613 2707 627
rect 2913 613 2927 627
rect 6673 613 6687 627
rect 6753 612 6767 626
rect 11973 613 11987 627
rect 57 573 71 587
rect 10953 573 10967 587
rect 11013 573 11027 587
rect 6873 513 6887 527
rect 493 473 507 487
rect 5153 473 5167 487
rect 11773 473 11787 487
rect 2213 433 2227 447
rect 2833 413 2847 427
rect 2973 413 2987 427
rect 4413 413 4427 427
rect 4593 413 4607 427
rect 5933 416 5947 430
rect 6033 413 6047 427
rect 9213 413 9227 427
rect 9233 413 9247 427
rect 9413 413 9427 427
rect 12173 412 12187 426
rect 12213 413 12227 427
rect 5693 393 5707 407
rect 5753 393 5767 407
rect 6073 373 6087 387
rect 6113 373 6127 387
rect 713 333 727 347
rect 793 333 807 347
rect 913 333 927 347
rect 10273 333 10287 347
rect 10393 333 10407 347
rect 10473 333 10487 347
rect 11033 333 11047 347
rect 11873 333 11887 347
rect 11913 332 11927 346
rect 11233 313 11247 327
rect 1213 193 1227 207
rect 1293 193 1307 207
rect 5453 193 5467 207
rect 5493 193 5507 207
rect 1253 173 1267 187
rect 1273 133 1287 147
rect 1233 113 1247 127
rect 1313 113 1327 127
rect 4033 113 4047 127
rect 4113 113 4127 127
rect 10953 113 10967 127
rect 11073 113 11087 127
rect 1253 93 1267 107
rect 4053 53 4067 67
rect 6313 53 6327 67
rect 8053 53 8067 67
rect 8393 53 8407 67
rect 10853 53 10867 67
rect 2515 33 2529 47
<< metal2 >>
rect 4096 12247 4103 12283
rect 316 11767 323 12136
rect 396 12107 403 12173
rect 496 12136 503 12173
rect 2113 12147 2127 12153
rect 336 11807 343 11833
rect 236 11687 243 11763
rect 256 11663 263 11753
rect 396 11747 403 12093
rect 416 11887 423 12133
rect 476 12100 483 12103
rect 473 12087 487 12100
rect 516 11927 523 12103
rect 836 12104 843 12133
rect 736 12100 743 12103
rect 456 11767 463 11836
rect 516 11800 523 11803
rect 513 11787 527 11800
rect 576 11787 583 11836
rect 236 11656 263 11663
rect 236 11616 243 11656
rect 273 11620 287 11633
rect 276 11616 283 11620
rect 336 11584 343 11633
rect 596 11587 603 11813
rect 676 11687 683 11933
rect 716 11804 723 12093
rect 733 12087 747 12100
rect 796 11836 803 11873
rect 916 11850 923 11913
rect 776 11687 783 11790
rect 256 11527 263 11583
rect 216 11316 223 11513
rect 176 10763 183 11096
rect 316 10803 323 10833
rect 296 10796 323 10803
rect 176 10756 193 10763
rect 236 10627 243 10723
rect 216 10327 223 10543
rect 316 10327 323 10796
rect 276 10276 283 10313
rect 256 10107 263 10243
rect 196 10016 223 10023
rect 196 9767 203 10016
rect 216 9756 223 9973
rect 256 9907 263 10023
rect 196 9547 203 9713
rect 236 9687 243 9723
rect 233 9540 247 9553
rect 236 9536 243 9540
rect 276 9507 283 9553
rect 213 9240 227 9253
rect 216 9236 223 9240
rect 256 9236 263 9273
rect 296 9247 303 9893
rect 196 9167 203 9193
rect 236 9183 243 9203
rect 236 9176 263 9183
rect 236 9016 243 9153
rect 256 9147 263 9176
rect 216 8767 223 8983
rect 216 8716 223 8753
rect 256 8716 263 8793
rect 236 8510 243 8683
rect 276 8567 283 8683
rect 296 8467 303 8613
rect 316 8507 323 9016
rect 336 8647 343 11570
rect 476 11427 483 11583
rect 513 11567 527 11570
rect 456 11316 463 11413
rect 676 11387 683 11673
rect 796 11616 803 11733
rect 816 11647 823 11803
rect 696 11427 703 11616
rect 820 11584 833 11587
rect 736 11580 743 11583
rect 733 11567 747 11580
rect 776 11347 783 11583
rect 827 11573 833 11584
rect 416 11096 443 11103
rect 416 11067 423 11096
rect 556 11063 563 11333
rect 733 11320 747 11333
rect 796 11323 803 11373
rect 736 11316 743 11320
rect 776 11316 803 11323
rect 536 11056 563 11063
rect 556 10847 563 11056
rect 576 10947 583 11133
rect 616 11107 623 11316
rect 576 10796 583 10933
rect 496 10667 503 10796
rect 600 10763 613 10767
rect 556 10707 563 10763
rect 596 10756 613 10763
rect 600 10753 613 10756
rect 667 10753 673 10767
rect 456 10427 463 10543
rect 496 10467 503 10543
rect 556 10527 563 10653
rect 556 10290 563 10413
rect 356 10207 363 10276
rect 396 10244 403 10276
rect 356 8984 363 9573
rect 396 9407 403 10230
rect 536 10207 543 10243
rect 536 10056 543 10093
rect 456 9987 463 10053
rect 496 9783 503 9993
rect 516 9987 523 10023
rect 496 9776 523 9783
rect 516 9756 523 9776
rect 436 9723 443 9756
rect 436 9716 463 9723
rect 456 9536 463 9716
rect 476 9500 483 9503
rect 376 9204 383 9236
rect 356 8567 363 8733
rect 336 8464 343 8493
rect 236 8196 243 8233
rect 216 8143 223 8163
rect 216 8136 243 8143
rect 236 7976 243 8136
rect 316 8107 323 8196
rect 276 7976 283 8013
rect 216 7887 223 7943
rect 316 7907 323 8013
rect 256 7676 263 7713
rect 176 7587 183 7676
rect 236 7607 243 7643
rect 236 7456 243 7572
rect 216 7367 223 7423
rect 256 7420 263 7423
rect 253 7407 267 7420
rect 316 7367 323 7893
rect 216 7156 223 7193
rect 276 7116 293 7123
rect 236 6936 243 7089
rect 216 6867 223 6903
rect 256 6787 263 6903
rect 296 6787 303 7113
rect 316 6867 323 7156
rect 336 7127 343 7630
rect 356 7627 363 8553
rect 376 7607 383 9190
rect 396 8167 403 9393
rect 436 9147 443 9490
rect 473 9487 487 9500
rect 556 9467 563 10023
rect 576 9647 583 9756
rect 496 9236 503 9273
rect 516 9167 523 9203
rect 416 8507 423 8973
rect 496 8807 503 8983
rect 436 8687 443 8753
rect 493 8720 507 8733
rect 496 8716 503 8720
rect 536 8716 543 8933
rect 596 8807 603 10693
rect 616 10590 623 10653
rect 616 9907 623 10576
rect 636 10207 643 10733
rect 696 10667 703 11096
rect 716 10583 723 11283
rect 756 11110 763 11133
rect 836 10987 843 11333
rect 856 10827 863 11633
rect 876 11284 883 11673
rect 896 11587 903 11613
rect 916 11584 923 11836
rect 916 11287 923 11570
rect 976 11507 983 12103
rect 1016 11807 1023 12103
rect 1056 12087 1063 12133
rect 1116 11767 1123 11803
rect 1176 11647 1183 11836
rect 1196 11767 1203 11853
rect 1276 11787 1283 12103
rect 1356 11836 1363 12090
rect 1413 11840 1427 11853
rect 1416 11836 1423 11840
rect 1516 11804 1523 12103
rect 1576 12087 1583 12136
rect 1696 12047 1703 12136
rect 2156 12104 2163 12133
rect 1736 12100 1743 12103
rect 1733 12087 1747 12100
rect 1776 12087 1783 12103
rect 1636 11836 1643 11873
rect 1336 11767 1343 11803
rect 1396 11783 1403 11803
rect 1656 11800 1663 11803
rect 1653 11787 1667 11800
rect 1396 11776 1423 11783
rect 1113 11620 1127 11633
rect 1116 11616 1123 11620
rect 1156 11587 1163 11633
rect 1096 11507 1103 11583
rect 813 10800 827 10813
rect 816 10796 823 10800
rect 856 10796 903 10803
rect 896 10707 903 10796
rect 936 10627 943 11413
rect 1033 11320 1047 11333
rect 1036 11316 1043 11320
rect 976 11227 983 11283
rect 1076 11247 1083 11316
rect 1176 11247 1183 11633
rect 1196 11630 1203 11753
rect 1316 11647 1323 11693
rect 1313 11620 1327 11633
rect 1316 11616 1323 11620
rect 1196 11347 1203 11616
rect 976 11067 983 11213
rect 1036 11096 1043 11153
rect 1016 10667 1023 11063
rect 1056 11007 1063 11063
rect 1116 10987 1123 11096
rect 1156 11064 1163 11153
rect 1076 10827 1083 10973
rect 1076 10796 1083 10813
rect 1096 10707 1103 10763
rect 696 10576 723 10583
rect 776 10576 783 10613
rect 656 9587 663 10573
rect 696 10544 703 10576
rect 756 10407 763 10543
rect 856 10407 863 10576
rect 1016 10540 1023 10543
rect 1013 10527 1027 10540
rect 776 10276 783 10313
rect 813 10280 827 10293
rect 816 10276 823 10280
rect 856 10247 863 10393
rect 756 10207 763 10243
rect 756 10056 763 10093
rect 696 9727 703 9833
rect 776 9770 783 10023
rect 736 9550 743 9693
rect 756 9647 763 9723
rect 876 9550 883 9753
rect 656 9507 663 9536
rect 716 9483 723 9503
rect 707 9476 723 9483
rect 676 9267 683 9453
rect 676 9207 683 9253
rect 676 8684 683 8933
rect 696 8847 703 9473
rect 756 9467 763 9503
rect 836 9487 843 9533
rect 776 9236 783 9293
rect 836 9167 843 9193
rect 796 9016 803 9073
rect 736 8947 743 8983
rect 776 8887 783 8983
rect 836 8947 843 9033
rect 733 8720 747 8733
rect 736 8716 743 8720
rect 776 8716 783 8833
rect 816 8716 823 8793
rect 796 8667 803 8683
rect 756 8496 763 8633
rect 796 8627 803 8653
rect 796 8496 803 8533
rect 496 8460 503 8463
rect 456 8287 463 8450
rect 493 8447 507 8460
rect 776 8460 783 8463
rect 556 8196 563 8233
rect 596 8196 603 8313
rect 576 8160 583 8163
rect 573 8147 587 8160
rect 516 7976 523 8133
rect 536 7907 543 7943
rect 536 7767 543 7893
rect 636 7747 643 8313
rect 656 7827 663 8433
rect 536 7676 543 7713
rect 576 7690 583 7733
rect 416 7107 423 7676
rect 516 7640 523 7643
rect 513 7627 527 7640
rect 496 7456 503 7613
rect 456 7416 483 7423
rect 436 7127 443 7156
rect 456 7127 463 7416
rect 516 7407 523 7423
rect 516 7396 533 7407
rect 520 7393 533 7396
rect 493 7160 507 7173
rect 496 7156 503 7160
rect 556 7167 563 7413
rect 576 7127 583 7456
rect 596 7447 603 7630
rect 616 7427 623 7673
rect 656 7407 663 7673
rect 656 7187 663 7393
rect 676 7207 683 7873
rect 696 7607 703 8450
rect 773 8447 787 8460
rect 856 8427 863 8593
rect 716 7690 723 8193
rect 756 8143 763 8353
rect 796 8210 803 8413
rect 836 8196 843 8233
rect 756 8136 773 8143
rect 776 7990 783 8133
rect 816 8107 823 8163
rect 816 7940 823 7943
rect 813 7927 827 7940
rect 840 7683 853 7687
rect 836 7676 853 7683
rect 840 7673 853 7676
rect 796 7487 803 7613
rect 816 7607 823 7643
rect 876 7487 883 8153
rect 896 7607 903 10010
rect 936 9587 943 10276
rect 976 9770 983 10453
rect 1096 10407 1103 10693
rect 1013 10290 1027 10293
rect 1016 10243 1023 10276
rect 1016 10236 1043 10243
rect 1036 10056 1043 10236
rect 1076 10207 1083 10243
rect 1116 10027 1123 10243
rect 1156 10027 1163 10276
rect 1056 10020 1063 10023
rect 1053 10007 1067 10020
rect 996 9756 1003 9893
rect 996 9536 1003 9573
rect 916 8164 923 8613
rect 793 7460 807 7473
rect 796 7456 803 7460
rect 727 7423 740 7427
rect 727 7420 743 7423
rect 727 7413 747 7420
rect 733 7407 747 7413
rect 776 7407 783 7423
rect 767 7396 783 7407
rect 767 7393 780 7396
rect 676 7170 683 7193
rect 596 6943 603 7153
rect 587 6936 603 6943
rect 476 6867 483 6903
rect 207 6643 220 6647
rect 207 6636 223 6643
rect 207 6633 220 6636
rect 256 6600 263 6603
rect 253 6587 267 6600
rect 296 6587 303 6713
rect 256 6416 263 6473
rect 207 6383 220 6387
rect 207 6376 223 6383
rect 207 6373 220 6376
rect 16 5827 23 6153
rect 216 6116 223 6193
rect 256 6007 263 6083
rect 36 5787 43 5933
rect 76 5867 83 5893
rect 56 5807 63 5853
rect 256 5827 263 5863
rect 16 5607 23 5633
rect 256 5527 263 5563
rect 256 5376 303 5383
rect 296 5347 303 5376
rect 207 5343 220 5347
rect 207 5336 223 5343
rect 207 5333 220 5336
rect 396 5287 403 6813
rect 436 6387 443 6653
rect 473 6640 487 6653
rect 476 6636 483 6640
rect 516 6636 523 6673
rect 456 6567 463 6593
rect 576 6507 583 6936
rect 516 6416 523 6453
rect 636 6430 643 6590
rect 676 6567 683 6973
rect 696 6607 703 7273
rect 836 6904 843 6953
rect 796 6867 803 6903
rect 876 6867 883 7156
rect 896 7127 903 7410
rect 896 6950 903 7092
rect 776 6636 783 6753
rect 796 6600 803 6603
rect 756 6583 763 6590
rect 793 6587 807 6600
rect 756 6576 783 6583
rect 776 6416 783 6576
rect 576 6387 583 6413
rect 207 5083 220 5087
rect 207 5076 223 5083
rect 207 5073 220 5076
rect 296 5043 303 5073
rect 256 5036 303 5043
rect 236 4856 243 4993
rect 187 4556 223 4563
rect 296 4147 303 4856
rect 296 4003 303 4033
rect 256 3996 303 4003
rect 256 3856 263 3933
rect 296 3816 323 3823
rect 16 3627 23 3773
rect 236 3563 243 3733
rect 227 3556 243 3563
rect 216 3516 223 3553
rect 196 3407 203 3483
rect 176 3007 183 3073
rect 276 3007 283 3393
rect 296 3310 303 3553
rect 316 3387 323 3816
rect 336 3530 343 4553
rect 396 3903 403 5273
rect 416 4867 423 5493
rect 436 5007 443 6193
rect 536 6127 543 6383
rect 516 6047 523 6083
rect 536 5896 583 5903
rect 456 5863 463 5896
rect 456 5856 483 5863
rect 476 5596 483 5856
rect 576 5847 583 5896
rect 496 5487 503 5563
rect 496 5376 503 5433
rect 616 5107 623 6173
rect 636 5507 643 6416
rect 796 6347 803 6383
rect 756 6116 763 6333
rect 836 6247 843 6603
rect 876 6287 883 6753
rect 856 6047 863 6213
rect 656 5567 663 5933
rect 716 5707 723 5853
rect 756 5847 763 5863
rect 747 5836 763 5847
rect 747 5833 760 5836
rect 776 5807 783 5853
rect 796 5807 803 5993
rect 896 5907 903 6936
rect 916 6587 923 7976
rect 936 7667 943 9113
rect 956 8367 963 9433
rect 976 9407 983 9503
rect 1016 9347 1023 9503
rect 996 9236 1003 9293
rect 1096 9204 1103 9893
rect 1196 9803 1203 11333
rect 1316 11316 1323 11373
rect 1256 11147 1263 11283
rect 1336 11096 1343 11233
rect 1276 10987 1283 11063
rect 1376 10987 1383 11316
rect 1396 11287 1403 11753
rect 1416 11387 1423 11776
rect 1576 11616 1583 11693
rect 1596 11387 1603 11583
rect 1593 11320 1607 11333
rect 1596 11316 1603 11320
rect 1736 11327 1743 12033
rect 1756 11587 1763 11836
rect 1396 11007 1403 11096
rect 1216 9867 1223 10813
rect 1356 10796 1363 10833
rect 1296 10687 1303 10763
rect 1376 10583 1383 10673
rect 1367 10577 1383 10583
rect 1356 10576 1383 10577
rect 1236 10536 1263 10543
rect 1236 10487 1243 10536
rect 1336 10276 1343 10473
rect 1316 10207 1323 10243
rect 1256 10007 1263 10023
rect 1196 9796 1223 9803
rect 1116 9250 1123 9753
rect 1196 9687 1203 9773
rect 1176 9627 1183 9653
rect 1156 9447 1163 9536
rect 1056 9087 1063 9190
rect 1033 9020 1047 9033
rect 1036 9016 1043 9020
rect 1056 8980 1063 8983
rect 1053 8967 1067 8980
rect 1116 8887 1123 9236
rect 996 8684 1003 8793
rect 1036 8680 1043 8683
rect 1033 8667 1047 8680
rect 1036 8496 1043 8613
rect 1076 8496 1083 8573
rect 1116 8510 1123 8713
rect 976 8407 983 8493
rect 956 7927 963 8193
rect 996 8123 1003 8413
rect 1016 8167 1023 8463
rect 1056 8460 1063 8463
rect 1053 8447 1067 8460
rect 1136 8230 1143 9253
rect 1156 9207 1163 9293
rect 1176 8984 1183 9233
rect 1196 9127 1203 9273
rect 1216 9087 1223 9796
rect 1256 9787 1263 9993
rect 1313 9760 1327 9773
rect 1316 9756 1323 9760
rect 1256 9720 1263 9723
rect 1236 9504 1243 9713
rect 1253 9707 1267 9720
rect 1296 9687 1303 9723
rect 1376 9707 1383 9793
rect 1316 9536 1323 9573
rect 1336 9500 1343 9503
rect 1296 9263 1303 9490
rect 1333 9487 1347 9500
rect 1376 9487 1383 9573
rect 1276 9256 1303 9263
rect 1276 9250 1283 9256
rect 1256 9127 1263 9203
rect 1376 9167 1383 9236
rect 1396 9207 1403 10993
rect 1416 10547 1423 10773
rect 1436 10087 1443 11213
rect 1456 10527 1463 10973
rect 1496 10707 1503 10813
rect 1516 10767 1523 11316
rect 1616 11147 1623 11283
rect 1576 10847 1583 11063
rect 1613 10800 1627 10813
rect 1656 10807 1663 11316
rect 1776 11247 1783 12073
rect 1796 11887 1803 12073
rect 1796 11547 1803 11873
rect 1953 11840 1967 11853
rect 1956 11836 1963 11840
rect 1996 11707 2003 11853
rect 2056 11807 2063 12103
rect 2236 11967 2243 12213
rect 2313 12167 2327 12173
rect 2436 12124 2443 12173
rect 2456 12116 2463 12213
rect 2773 12120 2787 12133
rect 2836 12130 2843 12193
rect 2776 12116 2783 12120
rect 2953 12120 2967 12133
rect 2956 12116 2963 12120
rect 2196 11836 2203 11933
rect 2336 11847 2343 12103
rect 2416 12047 2423 12083
rect 2416 11947 2423 12033
rect 2916 12007 2923 12073
rect 2240 11843 2253 11847
rect 2236 11836 2253 11843
rect 1853 11620 1867 11633
rect 1856 11616 1863 11620
rect 2136 11616 2143 11836
rect 2240 11833 2253 11836
rect 2376 11804 2383 11836
rect 2216 11767 2223 11803
rect 1936 11507 1943 11616
rect 1876 11316 1883 11493
rect 2036 11330 2043 11616
rect 1856 11247 1863 11283
rect 1716 11064 1723 11133
rect 1836 11110 1843 11133
rect 1916 10987 1923 11096
rect 1956 11064 1963 11093
rect 1996 11064 2003 11133
rect 1616 10796 1623 10800
rect 1456 10467 1463 10513
rect 1416 10027 1423 10056
rect 1436 9727 1443 9773
rect 1236 8967 1243 9053
rect 1316 9016 1323 9053
rect 1353 9020 1367 9033
rect 1356 9016 1363 9020
rect 1256 8984 1263 9016
rect 1296 8980 1303 8983
rect 1156 8327 1163 8573
rect 1176 8327 1183 8450
rect 1256 8427 1263 8970
rect 1293 8967 1307 8980
rect 1296 8716 1303 8753
rect 1416 8747 1423 9016
rect 1376 8687 1383 8716
rect 1316 8547 1323 8683
rect 1316 8407 1323 8463
rect 1356 8387 1363 8463
rect 1093 8210 1107 8213
rect 1176 8203 1183 8313
rect 1176 8196 1193 8203
rect 976 8116 1003 8123
rect 936 7107 943 7456
rect 956 6967 963 7913
rect 976 7883 983 8116
rect 1053 7980 1067 7993
rect 1116 7987 1123 8163
rect 1056 7976 1063 7980
rect 1016 7940 1023 7943
rect 1013 7927 1027 7940
rect 976 7876 1003 7883
rect 996 7467 1003 7876
rect 1056 7787 1063 7873
rect 1027 7673 1033 7687
rect 1056 7676 1063 7773
rect 1076 7703 1083 7943
rect 1093 7703 1107 7713
rect 1076 7700 1107 7703
rect 1076 7696 1103 7700
rect 1096 7676 1103 7696
rect 1156 7644 1163 7673
rect 1036 7456 1043 7633
rect 1076 7456 1083 7593
rect 1056 7387 1063 7423
rect 1136 7127 1143 7410
rect 1056 6936 1063 7073
rect 1176 6987 1183 7613
rect 1196 7087 1203 8195
rect 1216 7067 1223 7976
rect 1116 6943 1123 6973
rect 1096 6936 1123 6943
rect 936 6827 943 6936
rect 1036 6827 1043 6903
rect 1076 6767 1083 6903
rect 956 6607 963 6713
rect 1076 6636 1083 6753
rect 1116 6650 1123 6813
rect 916 6187 923 6433
rect 976 6384 983 6633
rect 1056 6547 1063 6603
rect 1096 6600 1103 6603
rect 1093 6587 1107 6600
rect 1013 6420 1027 6433
rect 1016 6416 1023 6420
rect 1056 6416 1063 6493
rect 1096 6430 1103 6513
rect 1136 6427 1143 6603
rect 1236 6587 1243 8333
rect 1256 8210 1263 8233
rect 1373 8200 1387 8213
rect 1376 8196 1383 8200
rect 1256 8127 1263 8196
rect 1356 8160 1363 8163
rect 1353 8147 1367 8160
rect 1256 7367 1263 8113
rect 1356 7676 1363 7713
rect 1336 7483 1343 7643
rect 1316 7480 1343 7483
rect 1313 7476 1343 7480
rect 1313 7467 1327 7476
rect 1353 7460 1367 7473
rect 1396 7470 1403 7993
rect 1416 7947 1423 8733
rect 1436 7787 1443 8193
rect 1456 8007 1463 9793
rect 1496 9770 1503 10573
rect 1536 10367 1543 10796
rect 1596 10760 1603 10763
rect 1593 10747 1607 10760
rect 1596 10540 1603 10543
rect 1593 10527 1607 10540
rect 1736 10507 1743 10783
rect 1836 10576 1843 10613
rect 1816 10467 1823 10530
rect 1916 10467 1923 10493
rect 1656 10244 1663 10276
rect 1533 10060 1547 10073
rect 1536 10056 1543 10060
rect 1616 9907 1623 10243
rect 1596 9756 1603 9793
rect 1636 9770 1643 9833
rect 1656 9827 1663 10230
rect 1476 9187 1483 9553
rect 1496 9487 1503 9756
rect 1656 9724 1663 9813
rect 1553 9540 1567 9553
rect 1556 9536 1563 9540
rect 1596 9536 1603 9573
rect 1616 9567 1623 9710
rect 1476 9047 1483 9173
rect 1496 8967 1503 9473
rect 1576 9447 1583 9503
rect 1616 9500 1623 9503
rect 1613 9487 1627 9500
rect 1556 9236 1563 9273
rect 1596 9236 1603 9473
rect 1616 9447 1623 9473
rect 1676 9267 1683 10393
rect 1536 9200 1543 9203
rect 1533 9187 1547 9200
rect 1576 9167 1583 9203
rect 1596 9016 1603 9073
rect 1636 9016 1643 9233
rect 1676 8984 1683 9013
rect 1576 8980 1583 8983
rect 1573 8967 1587 8980
rect 1576 8767 1583 8953
rect 1476 8027 1483 8493
rect 1496 8187 1503 8213
rect 1496 7947 1503 8173
rect 1516 7990 1523 8496
rect 1536 8210 1543 8753
rect 1573 8720 1587 8732
rect 1576 8716 1583 8720
rect 1636 8680 1643 8683
rect 1633 8667 1647 8680
rect 1616 8547 1623 8613
rect 1616 8496 1623 8533
rect 1656 8510 1663 8613
rect 1696 8547 1703 9113
rect 1736 8687 1743 10193
rect 1756 9287 1763 10073
rect 1776 10067 1783 10093
rect 1816 10056 1823 10413
rect 1916 10276 1923 10453
rect 1976 10247 1983 10276
rect 1896 10107 1903 10243
rect 1836 10020 1843 10023
rect 1833 10007 1847 10020
rect 1876 10007 1883 10053
rect 1796 9567 1803 9893
rect 1916 9863 1923 10193
rect 1936 9887 1943 10243
rect 1916 9856 1943 9863
rect 1856 9756 1863 9853
rect 1836 9720 1843 9723
rect 1833 9707 1847 9720
rect 1876 9627 1883 9723
rect 1936 9547 1943 9856
rect 1836 9467 1843 9503
rect 1876 9327 1883 9503
rect 1756 8567 1763 9252
rect 1816 9243 1823 9293
rect 1776 9236 1823 9243
rect 1776 8587 1783 9236
rect 1876 9200 1883 9203
rect 1776 8464 1783 8573
rect 1596 8283 1603 8463
rect 1636 8460 1643 8463
rect 1633 8447 1647 8460
rect 1576 8276 1603 8283
rect 1576 8147 1583 8276
rect 1716 8163 1723 8233
rect 1756 8167 1763 8373
rect 1796 8347 1803 9190
rect 1873 9187 1887 9200
rect 1936 9187 1943 9353
rect 1876 9127 1883 9173
rect 1956 9107 1963 10053
rect 1816 8967 1823 9093
rect 1836 8887 1843 9053
rect 1876 8980 1883 8983
rect 1873 8967 1887 8980
rect 1916 8947 1923 8983
rect 1976 8967 1983 9553
rect 1996 8863 2003 10553
rect 2016 9987 2023 11233
rect 2036 11007 2043 11316
rect 2096 11287 2103 11533
rect 2116 11507 2123 11583
rect 2156 11547 2163 11583
rect 2176 11330 2183 11493
rect 2296 11330 2303 11693
rect 2336 11584 2343 11673
rect 2376 11647 2383 11790
rect 2416 11727 2423 11933
rect 2556 11856 2563 11933
rect 2996 11923 3003 12133
rect 2996 11916 3023 11923
rect 2436 11807 2443 11833
rect 2576 11727 2583 11813
rect 2373 11620 2387 11633
rect 2376 11616 2383 11620
rect 2416 11616 2423 11653
rect 2440 11583 2453 11587
rect 2436 11576 2453 11583
rect 2440 11573 2453 11576
rect 2476 11507 2483 11593
rect 2496 11567 2503 11633
rect 2536 11564 2543 11713
rect 2196 11227 2203 11283
rect 2236 11187 2243 11316
rect 2136 11096 2143 11173
rect 2076 10987 2083 11063
rect 2036 10687 2043 10753
rect 2056 10747 2063 10783
rect 2156 10727 2163 10993
rect 2076 10576 2083 10713
rect 2056 10367 2063 10543
rect 2096 10427 2103 10543
rect 2176 10447 2183 10770
rect 2236 10627 2243 11096
rect 2056 10207 2063 10353
rect 2196 10276 2203 10576
rect 2236 10290 2243 10613
rect 2276 10467 2283 10973
rect 2296 10567 2303 11316
rect 2316 10907 2323 11096
rect 2453 11087 2467 11093
rect 2376 10947 2383 11063
rect 2416 11060 2423 11063
rect 2413 11047 2427 11060
rect 2356 10796 2363 10893
rect 2316 10747 2323 10793
rect 2376 10576 2383 10693
rect 2436 10544 2443 10573
rect 2396 10487 2403 10543
rect 2116 10103 2123 10276
rect 2176 10207 2183 10243
rect 2216 10240 2223 10243
rect 2213 10227 2227 10240
rect 2276 10227 2283 10313
rect 2116 10096 2143 10103
rect 2136 10067 2143 10096
rect 2076 10007 2083 10023
rect 2056 9996 2073 10003
rect 2056 9724 2063 9996
rect 2116 9756 2123 9973
rect 2016 8927 2023 9693
rect 1996 8856 2013 8863
rect 1836 8327 1843 8670
rect 1936 8496 1943 8793
rect 1856 8187 1863 8496
rect 1916 8460 1923 8463
rect 1913 8447 1927 8460
rect 1956 8427 1963 8463
rect 1896 8196 1903 8373
rect 1976 8247 1983 8273
rect 1676 8127 1683 8163
rect 1696 8156 1723 8163
rect 1356 7456 1363 7460
rect 1376 7387 1383 7423
rect 1416 7420 1423 7423
rect 1413 7407 1427 7420
rect 1176 6527 1183 6553
rect 1156 6396 1163 6453
rect 1216 6410 1223 6493
rect 936 5727 943 6373
rect 996 5947 1003 6173
rect 1036 6130 1043 6313
rect 1076 6287 1083 6383
rect 1116 6207 1123 6373
rect 1196 6147 1203 6353
rect 1256 6327 1263 7233
rect 1293 7160 1307 7173
rect 1296 7156 1303 7160
rect 1356 6936 1363 7053
rect 1396 6936 1403 6973
rect 1456 6927 1463 7456
rect 1276 6507 1283 6853
rect 1296 6567 1303 6833
rect 1336 6747 1343 6903
rect 1456 6527 1463 6636
rect 1476 6587 1483 7156
rect 1516 7047 1523 7976
rect 1676 7964 1683 8013
rect 1696 7956 1703 8156
rect 1996 8063 2003 8813
rect 2016 8087 2023 8853
rect 2036 8667 2043 9533
rect 2056 9467 2063 9710
rect 2093 9540 2107 9553
rect 2096 9536 2103 9540
rect 2136 9536 2143 9723
rect 2176 9547 2183 9873
rect 2116 9447 2123 9503
rect 2056 9167 2063 9313
rect 2196 9307 2203 9893
rect 2216 9367 2223 10053
rect 2153 9240 2167 9253
rect 2156 9236 2163 9240
rect 2076 9207 2083 9236
rect 2176 9167 2183 9203
rect 2056 9030 2063 9153
rect 2236 9107 2243 10213
rect 2316 10207 2323 10273
rect 2356 10227 2363 10473
rect 2376 10290 2383 10373
rect 2456 10367 2463 11052
rect 2476 11047 2483 11113
rect 2476 10487 2483 11012
rect 2496 10767 2503 11270
rect 2496 10627 2503 10753
rect 2516 10507 2523 11513
rect 2536 11044 2543 11550
rect 2536 10830 2543 11030
rect 2316 10056 2323 10193
rect 2276 10016 2303 10023
rect 2276 9727 2283 10016
rect 2336 9987 2343 10023
rect 2376 9987 2383 10276
rect 2396 10027 2403 10353
rect 2427 10283 2440 10287
rect 2427 10276 2443 10283
rect 2516 10287 2523 10472
rect 2427 10273 2440 10276
rect 2456 10187 2463 10230
rect 2476 10007 2483 10213
rect 2536 10187 2543 10293
rect 2556 10147 2563 11633
rect 2576 11027 2583 11713
rect 2596 11607 2603 11823
rect 2616 11787 2623 11816
rect 2896 11727 2903 11810
rect 2916 11747 2923 11823
rect 3016 11747 3023 11916
rect 3196 11836 3203 11993
rect 3316 11907 3323 12083
rect 3356 12027 3363 12113
rect 3536 12007 3543 12103
rect 3576 12100 3583 12103
rect 3573 12087 3587 12100
rect 3296 11896 3313 11903
rect 3116 11667 3123 11733
rect 2796 11623 2803 11653
rect 2796 11620 2823 11623
rect 2796 11616 2827 11620
rect 2616 11587 2623 11613
rect 2813 11604 2827 11616
rect 2676 11567 2683 11583
rect 2687 11556 2703 11563
rect 2696 11316 2703 11556
rect 2716 11527 2723 11583
rect 2716 11467 2723 11513
rect 2673 11100 2687 11113
rect 2676 11096 2683 11100
rect 2607 11084 2620 11087
rect 2607 11073 2613 11084
rect 2776 11076 2783 11433
rect 2896 11284 2903 11393
rect 2953 11320 2967 11333
rect 2956 11316 2963 11320
rect 2936 11187 2943 11283
rect 3036 11227 3043 11333
rect 2656 10907 2663 11063
rect 2296 9643 2303 9973
rect 2316 9724 2323 9853
rect 2296 9636 2323 9643
rect 2216 9016 2223 9053
rect 2056 8827 2063 9016
rect 2156 8980 2163 8983
rect 2153 8967 2167 8980
rect 2096 8716 2103 8933
rect 2076 8680 2083 8683
rect 2073 8667 2087 8680
rect 2096 8347 2103 8496
rect 2116 8467 2123 8683
rect 2196 8627 2203 8970
rect 2236 8427 2243 8493
rect 2256 8347 2263 9490
rect 2276 8607 2283 9453
rect 2296 8947 2303 9053
rect 1996 8056 2023 8063
rect 1616 7907 1623 7943
rect 1596 7676 1603 7713
rect 1616 7640 1623 7643
rect 1613 7627 1627 7640
rect 1656 7456 1663 7676
rect 1536 6987 1543 7456
rect 1636 7387 1643 7423
rect 1736 7407 1743 7713
rect 1616 7327 1623 7353
rect 1576 7170 1583 7233
rect 1616 7156 1623 7313
rect 1656 6947 1663 7253
rect 1636 6936 1653 6943
rect 1496 6604 1503 6633
rect 1496 6567 1503 6590
rect 1276 6367 1283 6413
rect 1536 6396 1543 6673
rect 1656 6596 1683 6603
rect 1576 6356 1603 6363
rect 1116 6100 1123 6103
rect 1113 6087 1127 6100
rect 1036 5896 1043 5993
rect 996 5787 1003 5863
rect 1056 5787 1063 5853
rect 707 5603 720 5607
rect 707 5596 723 5603
rect 756 5596 763 5633
rect 707 5593 720 5596
rect 676 5327 683 5593
rect 696 5387 703 5553
rect 776 5507 783 5563
rect 816 5447 823 5653
rect 836 5527 843 5633
rect 756 5376 763 5413
rect 856 5356 863 5633
rect 1076 5627 1083 6083
rect 1076 5564 1083 5613
rect 776 5340 783 5343
rect 773 5327 787 5340
rect 456 4787 463 5033
rect 496 4967 503 5043
rect 536 4856 543 5063
rect 516 4556 523 4593
rect 556 4570 563 4810
rect 576 4747 583 4773
rect 416 4307 423 4336
rect 436 4303 443 4510
rect 556 4507 563 4556
rect 436 4296 483 4303
rect 536 4187 543 4336
rect 496 4000 503 4003
rect 493 3987 507 4000
rect 376 3896 403 3903
rect 336 3447 343 3516
rect 296 2847 303 3296
rect 336 2790 343 3153
rect 176 2743 183 2773
rect 176 2736 203 2743
rect 176 1970 183 2713
rect 196 2487 203 2736
rect 216 2707 223 2743
rect 256 2740 263 2743
rect 253 2727 267 2740
rect 216 2476 223 2533
rect 253 2480 267 2493
rect 256 2476 263 2480
rect 196 2267 203 2433
rect 236 2343 243 2443
rect 216 2336 243 2343
rect 216 2256 223 2336
rect 256 2256 263 2313
rect 296 2256 303 2493
rect 336 2227 343 2776
rect 196 2007 203 2213
rect 236 1987 243 2223
rect 196 1867 203 1923
rect 236 1767 243 1923
rect 236 1736 243 1753
rect 276 1736 283 1913
rect 296 1747 303 1993
rect 156 1187 163 1690
rect 316 1403 323 1753
rect 336 1449 343 1793
rect 356 1667 363 3893
rect 376 1867 383 3896
rect 516 3830 523 3993
rect 556 3947 563 4053
rect 576 4007 583 4733
rect 596 4327 603 5063
rect 596 3967 603 4133
rect 616 3847 623 4973
rect 636 4824 643 5313
rect 816 5247 823 5323
rect 956 5110 963 5233
rect 656 5047 663 5093
rect 676 4827 683 4953
rect 816 4856 823 4893
rect 856 4856 863 4933
rect 796 4787 803 4823
rect 896 4787 903 4853
rect 916 4787 923 5063
rect 996 4627 1003 5093
rect 1016 5070 1023 5153
rect 1136 4987 1143 5553
rect 1176 5356 1183 6090
rect 1216 5864 1223 6273
rect 1476 6067 1483 6096
rect 1276 5896 1283 5933
rect 1356 5896 1403 5903
rect 1396 5863 1403 5896
rect 1256 5707 1263 5733
rect 1336 5727 1343 5863
rect 1376 5856 1403 5863
rect 1256 5596 1263 5693
rect 1236 5560 1243 5563
rect 1196 5364 1203 5553
rect 1233 5547 1247 5560
rect 1196 5076 1203 5113
rect 1176 4947 1183 5043
rect 1276 4947 1283 5529
rect 1016 4667 1023 4893
rect 1056 4863 1063 4893
rect 1036 4856 1063 4863
rect 1036 4824 1043 4856
rect 1076 4783 1083 4823
rect 1076 4776 1103 4783
rect 636 3907 643 4313
rect 656 4167 663 4613
rect 773 4560 787 4573
rect 776 4556 783 4560
rect 696 4527 703 4556
rect 836 4547 843 4593
rect 1076 4576 1083 4613
rect 1096 4587 1103 4776
rect 1116 4767 1123 4823
rect 1176 4707 1183 4933
rect 1116 4607 1123 4653
rect 1256 4647 1263 4856
rect 1296 4727 1303 5393
rect 1316 5127 1323 5493
rect 1316 4967 1323 5076
rect 1336 4987 1343 5356
rect 1356 5023 1363 5596
rect 1376 5327 1383 5856
rect 1376 5047 1383 5173
rect 1356 5016 1383 5023
rect 1376 4856 1383 5016
rect 1396 4947 1403 5753
rect 1416 4987 1423 5953
rect 1436 5287 1443 5453
rect 1456 5407 1463 5933
rect 1496 5883 1503 6103
rect 1476 5876 1503 5883
rect 1476 5827 1483 5876
rect 1516 5863 1523 6093
rect 1536 5967 1543 6053
rect 1576 5947 1583 6313
rect 1596 6147 1603 6356
rect 1676 6287 1683 6596
rect 1696 6404 1703 7393
rect 1636 6107 1643 6133
rect 1656 6087 1663 6213
rect 1616 5896 1623 5973
rect 1676 5963 1683 6153
rect 1656 5956 1683 5963
rect 1496 5856 1523 5863
rect 1576 5860 1583 5863
rect 1496 5376 1503 5856
rect 1573 5847 1587 5860
rect 1656 5687 1663 5956
rect 1676 5807 1683 5933
rect 1696 5847 1703 6136
rect 1676 5707 1683 5733
rect 1656 5627 1663 5673
rect 1593 5600 1607 5613
rect 1596 5596 1603 5600
rect 1536 5507 1543 5563
rect 1576 5560 1583 5563
rect 1573 5547 1587 5560
rect 1436 5007 1443 5113
rect 1456 5087 1463 5313
rect 1476 5307 1483 5343
rect 1516 5287 1523 5343
rect 1496 5076 1503 5113
rect 1536 5076 1543 5233
rect 1576 5110 1583 5293
rect 1616 5223 1623 5513
rect 1636 5507 1643 5596
rect 1676 5587 1683 5613
rect 1696 5307 1703 5833
rect 1716 5767 1723 6613
rect 1716 5427 1723 5453
rect 1736 5447 1743 7372
rect 1776 7127 1783 7173
rect 1796 7147 1803 7813
rect 1896 7644 1903 7733
rect 1816 7287 1823 7353
rect 1836 7307 1843 7613
rect 1856 7207 1863 7630
rect 1936 7456 1943 7493
rect 1816 7167 1823 7193
rect 1833 7160 1847 7173
rect 1836 7156 1843 7160
rect 1876 7156 1883 7213
rect 1936 7176 1943 7353
rect 1976 7267 1983 8033
rect 2016 8007 2023 8056
rect 2036 7963 2043 8293
rect 2196 8196 2203 8233
rect 2076 7970 2083 8196
rect 2116 8127 2123 8196
rect 2256 8163 2263 8213
rect 2176 8107 2183 8163
rect 2216 8156 2263 8163
rect 2016 7956 2043 7963
rect 2116 7947 2123 7993
rect 1996 7287 2003 7753
rect 2036 7367 2043 7913
rect 2096 7676 2103 7913
rect 2136 7907 2143 7956
rect 2156 7827 2163 8073
rect 2056 7424 2063 7673
rect 2176 7456 2183 7993
rect 2196 7507 2203 7953
rect 2216 7887 2223 8073
rect 2256 8007 2263 8093
rect 2276 7987 2283 8533
rect 2296 8047 2303 8753
rect 2316 8087 2323 9636
rect 2336 9547 2343 9713
rect 2356 9607 2363 9710
rect 2396 9687 2403 9723
rect 2476 9687 2483 9793
rect 2336 9267 2343 9533
rect 2356 9504 2363 9533
rect 2476 9287 2483 9536
rect 2416 9236 2423 9273
rect 2336 8807 2343 9232
rect 2396 9147 2403 9203
rect 2436 9167 2443 9203
rect 2476 9016 2483 9133
rect 2496 9023 2503 10113
rect 2576 10087 2583 10813
rect 2656 10707 2663 10893
rect 2716 10807 2723 10993
rect 3056 10887 3063 11173
rect 3076 11083 3083 11653
rect 3116 11596 3123 11653
rect 3136 11247 3143 11433
rect 3216 11407 3223 11803
rect 3236 11467 3243 11596
rect 3176 11167 3183 11333
rect 3216 11316 3223 11353
rect 3296 11350 3303 11896
rect 3436 11767 3443 11836
rect 3496 11630 3503 11803
rect 3576 11727 3583 12073
rect 3516 11583 3523 11613
rect 3436 11580 3443 11583
rect 3433 11567 3447 11580
rect 3476 11576 3523 11583
rect 3507 11553 3513 11567
rect 3616 11447 3623 12193
rect 3636 12107 3643 12133
rect 3676 12047 3683 12133
rect 3756 12087 3763 12153
rect 3836 12136 3843 12173
rect 3873 12140 3887 12153
rect 3876 12136 3883 12140
rect 3807 12103 3820 12107
rect 3807 12096 3823 12103
rect 3807 12093 3820 12096
rect 3756 11836 3763 12073
rect 3916 12067 3923 12090
rect 3916 11827 3923 12053
rect 4136 11967 4143 12103
rect 4176 11967 4183 12233
rect 4536 12107 4543 12173
rect 4356 12027 4363 12103
rect 4556 12104 4563 12133
rect 4236 11856 4243 11893
rect 3736 11647 3743 11803
rect 3776 11584 3783 11633
rect 3696 11547 3703 11583
rect 3696 11367 3703 11533
rect 3736 11347 3743 11583
rect 3253 11320 3267 11333
rect 3256 11316 3263 11320
rect 3336 11247 3343 11303
rect 3596 11267 3603 11296
rect 3176 11107 3183 11153
rect 3596 11107 3603 11173
rect 3616 11127 3623 11333
rect 3756 11304 3763 11353
rect 3656 11247 3663 11303
rect 3076 11076 3103 11083
rect 3213 11080 3227 11093
rect 3587 11096 3603 11107
rect 3587 11093 3600 11096
rect 3273 11080 3287 11093
rect 3216 11076 3223 11080
rect 3276 11076 3283 11080
rect 2753 10800 2767 10813
rect 2756 10796 2763 10800
rect 2716 10767 2723 10793
rect 2676 10687 2683 10713
rect 2816 10667 2823 10783
rect 2876 10780 2883 10783
rect 2873 10767 2887 10780
rect 2876 10647 2883 10753
rect 2916 10687 2923 10873
rect 3236 10816 3243 11033
rect 3316 11007 3323 11093
rect 3316 10947 3323 10993
rect 3676 10987 3683 11073
rect 3696 11044 3703 11113
rect 3796 11043 3803 11713
rect 3776 11036 3803 11043
rect 3776 10907 3783 11036
rect 3276 10787 3283 10873
rect 2516 9427 2523 10013
rect 2536 9887 2543 10023
rect 2576 9907 2583 10010
rect 2496 9016 2523 9023
rect 2356 8967 2363 9013
rect 2376 8987 2383 9016
rect 2416 8947 2423 8983
rect 2456 8980 2463 8983
rect 2453 8967 2467 8980
rect 2356 8716 2363 8773
rect 2396 8680 2403 8683
rect 2393 8667 2407 8680
rect 2476 8667 2483 8893
rect 2376 8464 2383 8593
rect 2456 8407 2463 8463
rect 2333 8087 2347 8093
rect 2356 8027 2363 8313
rect 2376 8187 2383 8353
rect 2236 7944 2243 7973
rect 2333 7980 2347 7993
rect 2336 7976 2343 7980
rect 2256 7927 2263 7972
rect 2396 7967 2403 8273
rect 2436 8227 2443 8353
rect 2456 8347 2463 8393
rect 2496 8287 2503 8693
rect 2516 8667 2523 9016
rect 2536 8707 2543 9753
rect 2556 9467 2563 9633
rect 2576 9484 2583 9773
rect 2596 9667 2603 9973
rect 2616 9587 2623 10493
rect 2656 10247 2663 10543
rect 2756 10507 2763 10576
rect 2716 10276 2723 10373
rect 2756 10276 2763 10313
rect 2636 9767 2643 10133
rect 2696 10024 2703 10053
rect 2656 9756 2663 9853
rect 2716 9807 2723 9833
rect 2736 9790 2743 10073
rect 2756 9787 2763 10213
rect 2796 10127 2803 10613
rect 2900 10544 2920 10547
rect 2856 10523 2863 10543
rect 2907 10543 2920 10544
rect 2907 10536 2923 10543
rect 2907 10533 2920 10536
rect 2856 10516 2883 10523
rect 2796 10056 2803 10113
rect 2836 9867 2843 10023
rect 2876 9887 2883 10516
rect 2916 10447 2923 10493
rect 2916 9987 2923 10433
rect 2936 9867 2943 10273
rect 2956 10227 2963 10530
rect 2976 10287 2983 10673
rect 2993 10280 3007 10293
rect 3036 10287 3043 10576
rect 2996 10276 3003 10280
rect 3056 10247 3063 10313
rect 3016 10207 3023 10243
rect 3076 10227 3083 10633
rect 3156 10576 3163 10673
rect 3196 10576 3203 10713
rect 3256 10543 3263 10573
rect 3216 10536 3263 10543
rect 3296 10447 3303 10813
rect 3476 10796 3483 10833
rect 3513 10800 3527 10813
rect 3516 10796 3523 10800
rect 3336 10707 3343 10793
rect 3316 10544 3323 10673
rect 3376 10667 3383 10793
rect 3496 10583 3503 10763
rect 3556 10727 3563 10813
rect 3496 10576 3523 10583
rect 3516 10544 3523 10576
rect 3436 10507 3443 10543
rect 3596 10487 3603 10833
rect 3636 10463 3643 10893
rect 3636 10456 3663 10463
rect 3016 9987 3023 10193
rect 3136 10167 3143 10276
rect 3156 10207 3163 10333
rect 3176 10227 3183 10353
rect 3256 10276 3263 10333
rect 3316 10296 3323 10413
rect 3656 10307 3663 10456
rect 3676 10327 3683 10833
rect 3756 10796 3763 10833
rect 3796 10796 3803 11013
rect 3816 10803 3823 11333
rect 3836 11247 3843 11653
rect 3856 11110 3863 11813
rect 3876 11667 3883 11823
rect 3896 11407 3903 11753
rect 3996 11616 4003 11693
rect 4036 11616 4043 11713
rect 3956 11316 3963 11433
rect 3896 11096 3903 11173
rect 3936 11107 3943 11283
rect 4036 11247 4043 11533
rect 4116 11527 4123 11570
rect 3920 11063 3933 11067
rect 3816 10796 3843 10803
rect 3776 10727 3783 10763
rect 3736 10576 3743 10633
rect 3776 10627 3783 10713
rect 3816 10556 3823 10613
rect 3836 10567 3843 10796
rect 3856 10563 3863 10933
rect 3876 10707 3883 11063
rect 3916 11056 3933 11063
rect 3920 11053 3933 11056
rect 3896 10587 3903 10633
rect 3856 10556 3883 10563
rect 3756 10487 3763 10543
rect 3776 10387 3783 10413
rect 3796 10347 3803 10513
rect 3356 10227 3363 10263
rect 3616 10227 3623 10293
rect 3796 10267 3803 10333
rect 3036 10024 3043 10153
rect 3196 10107 3203 10213
rect 3636 10207 3643 10256
rect 3676 10107 3683 10263
rect 3196 10036 3203 10093
rect 2776 9807 2783 9833
rect 2756 9687 2763 9733
rect 2676 9536 2683 9673
rect 2556 9247 2563 9393
rect 2556 9204 2563 9233
rect 2576 8723 2583 9470
rect 2616 9407 2623 9503
rect 2596 8887 2603 9033
rect 2616 8985 2623 9333
rect 2656 9247 2663 9503
rect 2776 9467 2783 9743
rect 3036 9703 3043 9773
rect 3056 9744 3063 9893
rect 3076 9787 3083 9853
rect 3196 9743 3203 9973
rect 3236 9767 3243 10036
rect 3156 9740 3163 9743
rect 3153 9727 3167 9740
rect 3176 9736 3203 9743
rect 3036 9696 3063 9703
rect 2636 9147 2643 9236
rect 2776 9167 2783 9236
rect 2676 8923 2683 9093
rect 2676 8916 2703 8923
rect 2556 8716 2583 8723
rect 2596 8716 2603 8873
rect 2636 8716 2643 8773
rect 2536 8547 2543 8672
rect 2536 8367 2543 8493
rect 2556 8444 2563 8716
rect 2696 8687 2703 8916
rect 2616 8680 2623 8683
rect 2613 8667 2627 8680
rect 2656 8464 2663 8683
rect 2716 8496 2723 8613
rect 2736 8527 2743 8773
rect 2816 8647 2823 9633
rect 2856 9503 2863 9573
rect 2896 9536 2903 9593
rect 2856 9496 2883 9503
rect 2836 9067 2843 9193
rect 2836 8767 2843 9013
rect 2776 8460 2783 8463
rect 2773 8447 2787 8460
rect 2556 8327 2563 8430
rect 2556 8247 2563 8313
rect 2836 8287 2843 8533
rect 2513 8220 2527 8233
rect 2516 8216 2523 8220
rect 2413 8207 2427 8213
rect 2436 8196 2443 8213
rect 2573 8163 2587 8176
rect 2416 8047 2423 8153
rect 2456 8127 2463 8163
rect 2556 8160 2587 8163
rect 2556 8156 2583 8160
rect 2556 8107 2563 8156
rect 2836 8147 2843 8273
rect 2856 8227 2863 9273
rect 2876 8847 2883 9496
rect 2916 9467 2923 9503
rect 2916 8967 2923 9253
rect 2976 9236 2983 9333
rect 2996 9267 3003 9633
rect 3016 9504 3023 9553
rect 3036 9487 3043 9593
rect 3056 9287 3063 9696
rect 3076 9347 3083 9713
rect 3096 9507 3103 9593
rect 2996 9023 3003 9203
rect 2976 9016 3003 9023
rect 3056 9016 3063 9153
rect 3096 9087 3103 9472
rect 2896 8716 2903 8873
rect 2936 8716 2943 8853
rect 2976 8729 2983 9016
rect 3036 8980 3043 8983
rect 3076 8980 3083 8983
rect 3033 8967 3047 8980
rect 3073 8967 3087 8980
rect 3116 8947 3123 9613
rect 3176 9607 3183 9736
rect 3296 9607 3303 9756
rect 3136 9447 3143 9533
rect 3156 9467 3163 9593
rect 3316 9516 3323 9873
rect 3416 9756 3423 9833
rect 3516 9627 3523 9773
rect 3536 9707 3543 9993
rect 3556 9967 3563 10003
rect 3556 9647 3563 9953
rect 3616 9947 3623 10033
rect 3676 9907 3683 10093
rect 3596 9727 3603 9756
rect 3616 9607 3623 9893
rect 3696 9847 3703 10213
rect 3756 10023 3763 10253
rect 3816 10227 3823 10473
rect 3836 10307 3843 10513
rect 3836 10264 3843 10293
rect 3816 10056 3823 10192
rect 3876 10067 3883 10473
rect 3916 10347 3923 10993
rect 3956 10907 3963 11096
rect 3976 10967 3983 11093
rect 3996 11067 4003 11093
rect 4076 11064 4083 11153
rect 3976 10767 3983 10953
rect 4016 10810 4023 10933
rect 4116 10727 4123 11513
rect 4196 11427 4203 11823
rect 4276 11816 4303 11823
rect 4276 11767 4283 11816
rect 4276 11616 4283 11753
rect 4316 11616 4323 11693
rect 4356 11667 4363 11823
rect 4256 11547 4263 11583
rect 4296 11580 4303 11583
rect 4293 11567 4307 11580
rect 4376 11503 4383 11693
rect 4396 11527 4403 12090
rect 4576 12067 4583 12193
rect 4676 12136 4683 12193
rect 4716 12116 4723 12173
rect 4776 12116 4823 12123
rect 4656 12027 4663 12103
rect 4816 12083 4823 12116
rect 4796 12076 4823 12083
rect 4716 11870 4723 11893
rect 4656 11787 4663 11816
rect 4376 11496 4403 11503
rect 4236 11316 4243 11353
rect 4276 11330 4283 11493
rect 4356 11447 4363 11473
rect 4136 11107 4143 11316
rect 4296 11247 4303 11283
rect 4196 11007 4203 11063
rect 4256 11047 4263 11233
rect 4296 11110 4303 11233
rect 4336 11227 4343 11353
rect 4296 10987 4303 11096
rect 4176 10667 4183 10693
rect 4196 10647 4203 10893
rect 4336 10796 4343 11093
rect 4376 10816 4383 11453
rect 4396 11287 4403 11496
rect 4416 11247 4423 11616
rect 4496 11587 4503 11693
rect 4433 11487 4447 11493
rect 4456 11247 4463 11513
rect 4556 11507 4563 11583
rect 4493 11320 4507 11333
rect 4496 11316 4503 11320
rect 4536 11316 4543 11353
rect 4576 11330 4583 11533
rect 4676 11507 4683 11823
rect 4676 11387 4683 11413
rect 4696 11407 4703 11473
rect 4716 11343 4723 11653
rect 4736 11567 4743 11613
rect 4756 11467 4763 11856
rect 4776 11727 4783 11953
rect 4796 11667 4803 12076
rect 4976 11927 4983 12013
rect 5136 11987 5143 12083
rect 5176 12027 5183 12113
rect 4976 11836 4983 11913
rect 5136 11867 5143 11973
rect 4856 11616 4863 11733
rect 4896 11630 4903 11790
rect 4996 11783 5003 11803
rect 5056 11787 5063 11836
rect 4947 11776 5003 11783
rect 5156 11747 5163 11793
rect 5176 11767 5183 11836
rect 5196 11787 5203 11913
rect 5276 11850 5283 11913
rect 5336 11856 5343 11973
rect 5376 11887 5383 12103
rect 5436 12047 5443 12283
rect 9056 12187 9063 12213
rect 6036 12136 6043 12173
rect 6216 12147 6223 12173
rect 6216 12136 6233 12147
rect 5896 12104 5903 12133
rect 5516 12047 5523 12103
rect 5756 12100 5763 12103
rect 5753 12087 5767 12100
rect 5756 11927 5763 12073
rect 5796 11987 5803 12103
rect 5256 11787 5263 11803
rect 5247 11776 5263 11787
rect 5247 11773 5260 11776
rect 5356 11687 5363 11813
rect 5376 11787 5383 11823
rect 5656 11824 5663 11873
rect 5836 11867 5843 12033
rect 5916 11927 5923 12136
rect 6220 12133 6233 12136
rect 6056 12087 6063 12103
rect 6216 12087 6223 12116
rect 6536 12080 6543 12083
rect 6056 12027 6063 12073
rect 6136 11987 6143 12073
rect 6216 12007 6223 12073
rect 6533 12067 6547 12080
rect 4776 11507 4783 11593
rect 4796 11527 4803 11616
rect 5296 11596 5303 11653
rect 5360 11603 5373 11607
rect 5356 11596 5373 11603
rect 5360 11593 5373 11596
rect 4836 11580 4843 11583
rect 4833 11567 4847 11580
rect 4876 11407 4883 11583
rect 4936 11467 4943 11563
rect 5056 11350 5063 11453
rect 5256 11427 5263 11590
rect 4716 11336 4743 11343
rect 4736 11304 4743 11336
rect 4436 11047 4443 11063
rect 4476 11060 4483 11063
rect 4473 11047 4487 11060
rect 4436 10907 4443 11033
rect 4496 11007 4503 11053
rect 4516 10947 4523 11270
rect 4556 11247 4563 11283
rect 4616 11207 4623 11293
rect 4536 11027 4543 11193
rect 4636 11047 4643 11303
rect 5096 11307 5103 11393
rect 5016 11203 5023 11253
rect 4996 11196 5023 11203
rect 4716 11096 4723 11133
rect 4696 11060 4703 11063
rect 4693 11047 4707 11060
rect 4796 10987 4803 11096
rect 4876 11047 4883 11133
rect 4256 10607 4263 10693
rect 4236 10427 4243 10523
rect 4276 10487 4283 10763
rect 4396 10727 4403 10773
rect 4296 10587 4303 10713
rect 4416 10607 4423 10783
rect 4696 10764 4703 10913
rect 4716 10776 4743 10783
rect 4356 10567 4363 10593
rect 4356 10507 4363 10553
rect 3936 10387 3943 10413
rect 3756 10016 3783 10023
rect 3796 10020 3803 10023
rect 3693 9760 3707 9773
rect 3696 9756 3703 9760
rect 3676 9720 3683 9723
rect 3716 9720 3723 9723
rect 3673 9707 3687 9720
rect 3713 9707 3727 9720
rect 3756 9707 3763 9833
rect 3616 9523 3623 9593
rect 3616 9516 3643 9523
rect 3236 9483 3243 9503
rect 3736 9487 3743 9516
rect 3236 9476 3263 9483
rect 3193 9427 3207 9433
rect 3136 8967 3143 9013
rect 2876 8347 2883 8673
rect 3056 8667 3063 8933
rect 2896 8327 2903 8413
rect 2916 8407 2923 8633
rect 2936 8387 2943 8653
rect 3036 8527 3043 8573
rect 3096 8476 3103 8873
rect 3156 8787 3163 9413
rect 3176 8827 3183 9333
rect 3196 8867 3203 9373
rect 3236 9236 3243 9453
rect 3256 9347 3263 9476
rect 3316 9427 3323 9453
rect 3416 9267 3423 9393
rect 3256 9167 3263 9203
rect 3336 9167 3343 9223
rect 3276 8987 3283 9153
rect 3316 8887 3323 8983
rect 3396 8907 3403 9223
rect 3416 8947 3423 9213
rect 3436 8750 3443 9353
rect 3716 9287 3723 9413
rect 3736 9347 3743 9473
rect 3756 9327 3763 9633
rect 3776 9467 3783 10016
rect 3793 10007 3807 10020
rect 3836 10003 3843 10023
rect 3836 9996 3863 10003
rect 3796 9687 3803 9773
rect 3796 9427 3803 9533
rect 3816 9367 3823 9773
rect 3756 9267 3763 9313
rect 3836 9267 3843 9893
rect 3856 9867 3863 9996
rect 3896 9907 3903 10313
rect 3956 10283 3963 10373
rect 3976 10347 3983 10393
rect 3936 10276 3963 10283
rect 3973 10280 3987 10293
rect 3976 10276 3983 10280
rect 4016 10276 4023 10333
rect 4076 10310 4083 10413
rect 4100 10327 4107 10353
rect 3936 10247 3943 10276
rect 3876 9727 3883 9853
rect 3896 9767 3903 9853
rect 3916 9787 3923 10053
rect 3936 9927 3943 10212
rect 3956 9967 3963 10133
rect 3976 10070 3983 10193
rect 3956 9783 3963 9853
rect 3976 9847 3983 10056
rect 3996 10007 4003 10243
rect 4096 10147 4103 10253
rect 4396 10207 4403 10573
rect 4496 10576 4503 10673
rect 4416 10407 4423 10572
rect 4556 10544 4563 10573
rect 4616 10547 4623 10593
rect 4476 10387 4483 10543
rect 4416 10187 4423 10256
rect 4436 10227 4443 10263
rect 4496 10127 4503 10263
rect 4536 10227 4543 10513
rect 4093 10060 4107 10073
rect 4096 10056 4103 10060
rect 3956 9776 3983 9783
rect 3976 9756 3983 9776
rect 3996 9770 4003 9853
rect 4016 9807 4023 10056
rect 4076 9967 4083 10023
rect 4036 9776 4043 9953
rect 4076 9927 4083 9953
rect 4116 9907 4123 10023
rect 4136 9947 4143 10013
rect 4176 9947 4183 10003
rect 4496 9867 4503 10073
rect 4536 10050 4543 10213
rect 4556 10087 4563 10373
rect 4596 10247 4603 10433
rect 3876 9367 3883 9692
rect 3916 9687 3923 9723
rect 3956 9687 3963 9723
rect 4056 9687 4063 9736
rect 3916 9536 3923 9673
rect 4016 9504 4023 9533
rect 3747 9256 3763 9267
rect 3747 9253 3760 9256
rect 3456 9187 3463 9253
rect 3716 9216 3743 9223
rect 3196 8640 3203 8643
rect 3193 8627 3207 8640
rect 3376 8607 3383 8715
rect 3376 8567 3383 8593
rect 2996 8447 3003 8463
rect 3356 8447 3363 8513
rect 3396 8483 3403 8733
rect 3476 8730 3483 9073
rect 3516 8967 3523 9016
rect 3516 8587 3523 8893
rect 3416 8547 3423 8573
rect 3376 8476 3403 8483
rect 3416 8476 3423 8533
rect 3473 8480 3487 8493
rect 3476 8476 3483 8480
rect 2987 8436 3003 8447
rect 2987 8433 3000 8436
rect 2876 8147 2883 8183
rect 2436 7967 2443 8013
rect 2456 7956 2463 8073
rect 2836 8027 2843 8133
rect 2476 7964 2483 7993
rect 2776 7956 2783 8013
rect 2276 7907 2283 7933
rect 2236 7347 2243 7893
rect 2316 7827 2323 7943
rect 2436 7643 2443 7793
rect 2416 7636 2443 7643
rect 2376 7471 2383 7603
rect 2376 7456 2383 7457
rect 1856 7087 1863 7123
rect 1916 6936 1923 6993
rect 1756 6167 1763 6933
rect 1776 6447 1783 6936
rect 1856 6900 1863 6903
rect 1853 6887 1867 6900
rect 1856 6827 1863 6873
rect 1896 6767 1903 6890
rect 1956 6887 1963 7133
rect 1976 6867 1983 7143
rect 1996 7107 2003 7136
rect 1876 6636 1883 6673
rect 1776 6327 1783 6433
rect 1836 6416 1843 6573
rect 1856 6567 1863 6603
rect 1876 6416 1883 6573
rect 1896 6487 1903 6603
rect 1816 6347 1823 6383
rect 1856 6367 1863 6383
rect 1916 6367 1923 6513
rect 1856 6356 1873 6367
rect 1860 6353 1873 6356
rect 1813 6167 1827 6173
rect 1753 6127 1767 6132
rect 1836 6116 1843 6153
rect 1816 6047 1823 6083
rect 1756 5563 1763 5813
rect 1796 5727 1803 5973
rect 1876 5967 1883 6332
rect 1896 6087 1903 6116
rect 1916 6067 1923 6233
rect 1896 5896 1903 5973
rect 1856 5787 1863 5863
rect 1793 5600 1807 5613
rect 1833 5600 1847 5613
rect 1796 5596 1803 5600
rect 1836 5596 1843 5600
rect 1876 5567 1883 5850
rect 1756 5556 1783 5563
rect 1776 5376 1783 5556
rect 1596 5216 1623 5223
rect 1596 5167 1603 5216
rect 1696 5207 1703 5293
rect 1756 5287 1763 5330
rect 1796 5267 1803 5343
rect 1813 5247 1827 5253
rect 1836 5247 1843 5376
rect 1856 5344 1863 5413
rect 1826 5240 1827 5247
rect 1616 5127 1623 5173
rect 1356 4767 1363 4823
rect 1396 4820 1403 4823
rect 1393 4807 1407 4820
rect 1436 4807 1443 4972
rect 1476 4907 1483 5043
rect 1416 4587 1423 4633
rect 1496 4627 1503 4973
rect 1516 4783 1523 5043
rect 1556 4807 1563 5033
rect 1576 4823 1583 4933
rect 1616 4887 1623 5063
rect 1607 4863 1620 4867
rect 1607 4856 1623 4863
rect 1656 4856 1663 4953
rect 1607 4853 1620 4856
rect 1576 4816 1603 4823
rect 1516 4776 1543 4783
rect 1516 4667 1523 4733
rect 1013 4560 1027 4573
rect 1016 4556 1023 4560
rect 696 4336 703 4413
rect 756 4387 763 4523
rect 796 4520 803 4523
rect 793 4507 807 4520
rect 776 4316 783 4433
rect 836 4330 843 4493
rect 1036 4447 1043 4523
rect 1436 4507 1443 4543
rect 1496 4527 1503 4543
rect 1436 4447 1443 4493
rect 1496 4467 1503 4513
rect 1493 4387 1507 4393
rect 876 4324 883 4373
rect 656 4027 663 4073
rect 713 4040 727 4053
rect 716 4036 723 4040
rect 756 4036 763 4093
rect 816 4056 823 4153
rect 873 4003 887 4016
rect 696 3967 703 4003
rect 736 3967 743 4003
rect 856 4000 887 4003
rect 856 3996 883 4000
rect 856 3967 863 3996
rect 696 3907 703 3953
rect 1136 3907 1143 4193
rect 1196 4167 1203 4283
rect 1236 4227 1243 4313
rect 1376 4067 1383 4333
rect 1376 4024 1383 4053
rect 1176 3927 1183 4023
rect 456 3547 463 3813
rect 636 3796 643 3893
rect 1376 3887 1383 4010
rect 1396 4007 1403 4093
rect 1436 4043 1443 4290
rect 1516 4287 1523 4533
rect 1536 4387 1543 4776
rect 1416 4036 1443 4043
rect 1453 4040 1467 4053
rect 1456 4036 1463 4040
rect 1496 4036 1503 4193
rect 1416 3947 1423 4036
rect 1536 3987 1543 4053
rect 1556 3967 1563 4713
rect 1376 3873 1393 3887
rect 536 3587 543 3770
rect 553 3520 567 3533
rect 556 3516 563 3520
rect 656 3487 663 3753
rect 476 3296 483 3373
rect 516 3296 523 3453
rect 576 3447 583 3483
rect 556 3264 563 3293
rect 576 3010 583 3433
rect 676 3067 683 3833
rect 696 3767 703 3790
rect 972 3707 979 3733
rect 736 3296 743 3533
rect 776 3516 783 3573
rect 836 3264 843 3393
rect 996 3367 1003 3750
rect 1080 3707 1087 3733
rect 1376 3587 1383 3873
rect 1416 3796 1423 3893
rect 1436 3804 1443 3853
rect 1480 3803 1493 3807
rect 1476 3796 1493 3803
rect 1480 3793 1493 3796
rect 1100 3543 1113 3547
rect 1096 3533 1113 3543
rect 1096 3516 1103 3533
rect 1016 3487 1023 3516
rect 1176 3487 1183 3516
rect 1076 3407 1083 3483
rect 1116 3447 1123 3483
rect 756 3227 763 3263
rect 396 2964 403 2993
rect 436 2547 443 2833
rect 456 2744 463 2893
rect 476 2847 483 2963
rect 516 2907 523 2973
rect 556 2667 563 2693
rect 476 2263 483 2443
rect 536 2283 543 2633
rect 516 2276 543 2283
rect 516 2270 523 2276
rect 456 2256 483 2263
rect 556 2256 563 2653
rect 396 1970 403 2253
rect 456 2224 463 2256
rect 496 2107 503 2223
rect 536 2187 543 2223
rect 596 2187 603 2213
rect 616 2207 623 2473
rect 496 1956 503 1993
rect 536 1956 543 2133
rect 516 1807 523 1923
rect 493 1740 507 1753
rect 496 1736 503 1740
rect 556 1707 563 1853
rect 576 1807 583 1993
rect 596 1887 603 2093
rect 636 1924 643 3053
rect 676 2787 683 3013
rect 713 3000 727 3013
rect 716 2996 723 3000
rect 876 2967 883 3033
rect 896 2947 903 2993
rect 936 2964 943 3333
rect 1076 3296 1083 3333
rect 1056 3227 1063 3263
rect 1096 3127 1103 3263
rect 916 2956 933 2963
rect 776 2776 783 2813
rect 716 2476 723 2773
rect 756 2476 763 2743
rect 296 1396 323 1403
rect 256 1147 263 1363
rect 336 1230 343 1435
rect 336 1167 343 1216
rect 36 936 43 1073
rect 60 947 67 993
rect 356 887 363 1653
rect 496 1436 503 1493
rect 533 1440 547 1453
rect 536 1436 543 1440
rect 427 1276 483 1283
rect 376 947 383 1273
rect 436 1227 443 1253
rect 476 1216 483 1276
rect 516 1267 523 1403
rect 576 1223 583 1453
rect 567 1216 583 1223
rect 496 1147 503 1183
rect 407 1133 413 1147
rect 396 900 403 903
rect 393 887 407 900
rect 36 607 43 643
rect 60 587 67 633
rect 356 507 363 873
rect 376 707 383 733
rect 396 676 403 873
rect 453 680 467 693
rect 456 676 463 680
rect 516 607 523 1073
rect 556 847 563 1216
rect 616 904 623 1493
rect 636 707 643 1033
rect 656 807 663 2253
rect 676 1807 683 2293
rect 816 2270 823 2533
rect 896 2507 903 2933
rect 916 2744 923 2956
rect 976 2907 983 2963
rect 936 2727 943 2893
rect 996 2776 1003 2813
rect 1016 2740 1023 2743
rect 1013 2727 1027 2740
rect 953 2480 967 2493
rect 956 2476 963 2480
rect 916 2447 923 2476
rect 1056 2447 1063 2476
rect 976 2440 983 2443
rect 973 2427 987 2440
rect 1076 2427 1083 2773
rect 856 2256 863 2293
rect 787 2224 800 2227
rect 787 2213 793 2224
rect 876 2147 883 2223
rect 976 2067 983 2413
rect 1136 2287 1143 2713
rect 1156 2627 1163 3353
rect 1236 2996 1243 3293
rect 1276 3067 1283 3533
rect 1336 3516 1343 3573
rect 1296 3264 1303 3433
rect 1356 3296 1363 3373
rect 1396 3296 1403 3333
rect 1436 3267 1443 3516
rect 1516 3347 1523 3933
rect 1536 3467 1543 3952
rect 1576 3943 1583 4633
rect 1596 4527 1603 4816
rect 1616 4607 1623 4793
rect 1636 4767 1643 4823
rect 1596 4030 1603 4393
rect 1616 4307 1623 4593
rect 1636 4547 1643 4753
rect 1656 4747 1663 4793
rect 1676 4787 1683 4823
rect 1736 4747 1743 4873
rect 1636 4407 1643 4512
rect 1656 4367 1663 4693
rect 1676 4527 1683 4673
rect 1776 4583 1783 4933
rect 1756 4576 1783 4583
rect 1756 4556 1763 4576
rect 1796 4556 1803 4853
rect 1836 4576 1843 4893
rect 1876 4607 1883 4913
rect 1896 4867 1903 5613
rect 1916 5567 1923 5633
rect 1936 5167 1943 6593
rect 1956 5787 1963 6373
rect 1976 6247 1983 6636
rect 1996 6547 2003 6773
rect 1996 6130 2003 6273
rect 1996 6067 2003 6116
rect 1956 5347 1963 5773
rect 1976 5247 1983 6013
rect 1996 5247 2003 5633
rect 2016 5627 2023 6873
rect 2036 6587 2043 6973
rect 2176 6936 2183 7033
rect 2096 6827 2103 6936
rect 2156 6887 2163 6903
rect 2096 6607 2103 6813
rect 2156 6727 2163 6873
rect 2156 6650 2163 6673
rect 2193 6640 2207 6653
rect 2196 6636 2203 6640
rect 2133 6587 2147 6590
rect 2176 6547 2183 6603
rect 2116 6416 2123 6453
rect 2096 6367 2103 6383
rect 2087 6356 2103 6367
rect 2087 6353 2100 6356
rect 2053 6167 2067 6173
rect 2036 5627 2043 6053
rect 2156 6027 2163 6453
rect 2176 6007 2183 6393
rect 2236 6247 2243 6890
rect 2256 6527 2263 7410
rect 2296 7136 2323 7143
rect 2356 7136 2383 7143
rect 2296 6907 2303 6993
rect 2276 6507 2283 6653
rect 2276 6287 2283 6433
rect 2116 5896 2123 5993
rect 2176 5827 2183 5863
rect 2176 5647 2183 5713
rect 2136 5596 2143 5633
rect 2173 5587 2187 5596
rect 2036 5390 2043 5473
rect 2076 5376 2083 5493
rect 2116 5487 2123 5563
rect 2176 5363 2183 5533
rect 2196 5387 2203 5793
rect 2276 5787 2283 6070
rect 2296 5847 2303 6893
rect 2316 6867 2323 7136
rect 2376 7107 2383 7136
rect 2316 6447 2323 6853
rect 2336 6604 2343 6673
rect 2356 6467 2363 7073
rect 2336 6287 2343 6383
rect 2376 6143 2383 6453
rect 2396 6383 2403 7493
rect 2516 7416 2543 7423
rect 2436 7027 2443 7333
rect 2476 6936 2483 7153
rect 2536 7047 2543 7416
rect 2556 7247 2563 7753
rect 2616 7676 2623 7713
rect 2656 7676 2663 7813
rect 2636 7567 2643 7643
rect 2636 7470 2643 7553
rect 2776 7467 2783 7676
rect 2556 7167 2563 7233
rect 2596 7156 2603 7213
rect 2576 7120 2583 7123
rect 2573 7107 2587 7120
rect 2456 6900 2463 6903
rect 2453 6887 2467 6900
rect 2496 6607 2503 6733
rect 2456 6600 2463 6603
rect 2453 6587 2467 6600
rect 2516 6587 2523 6773
rect 2396 6376 2423 6383
rect 2356 6136 2383 6143
rect 2356 6116 2363 6136
rect 2396 6116 2403 6353
rect 2416 6130 2423 6376
rect 2476 6347 2483 6383
rect 2536 6347 2543 6793
rect 2336 6047 2343 6083
rect 2376 6080 2383 6083
rect 2373 6067 2387 6080
rect 2436 5910 2443 6053
rect 2476 6047 2483 6333
rect 2496 5863 2503 6153
rect 2316 5687 2323 5773
rect 2456 5747 2463 5863
rect 2476 5856 2503 5863
rect 2216 5507 2223 5573
rect 2236 5547 2243 5673
rect 2356 5596 2363 5673
rect 2393 5600 2407 5613
rect 2396 5596 2403 5600
rect 2253 5567 2267 5573
rect 2456 5567 2463 5693
rect 2476 5427 2483 5856
rect 2456 5364 2463 5393
rect 2176 5356 2203 5363
rect 2016 5147 2023 5333
rect 2056 5323 2063 5330
rect 2056 5316 2083 5323
rect 2036 5064 2043 5113
rect 1996 5027 2003 5063
rect 2007 5016 2023 5023
rect 1936 4856 1943 4993
rect 1976 4856 1983 4913
rect 1916 4767 1923 4823
rect 2016 4787 2023 5016
rect 2056 4687 2063 5293
rect 2076 4824 2083 5316
rect 2096 5187 2103 5343
rect 2456 5327 2463 5350
rect 2136 5316 2163 5323
rect 2096 4727 2103 5152
rect 2116 4967 2123 5213
rect 2136 5207 2143 5316
rect 2136 4907 2143 5193
rect 2156 5047 2163 5233
rect 2176 4907 2183 5133
rect 2276 5076 2283 5193
rect 2176 4856 2183 4893
rect 2196 4887 2203 5073
rect 2296 4967 2303 5043
rect 2216 4856 2223 4933
rect 1876 4536 1903 4543
rect 1736 4427 1743 4523
rect 1653 4340 1667 4353
rect 1656 4336 1663 4340
rect 1696 4336 1703 4393
rect 1736 4347 1743 4413
rect 1776 4387 1783 4523
rect 1636 3967 1643 4036
rect 1556 3936 1583 3943
rect 1556 3307 1563 3936
rect 1576 3527 1583 3793
rect 1636 3707 1643 3816
rect 1656 3787 1663 4273
rect 1716 4267 1723 4303
rect 1733 4287 1747 4293
rect 1676 3947 1683 4253
rect 1756 4247 1763 4353
rect 1836 4267 1843 4473
rect 1856 4427 1863 4536
rect 1696 4007 1703 4233
rect 1816 4067 1823 4113
rect 1836 4056 1843 4153
rect 1876 4107 1883 4513
rect 1896 4507 1903 4536
rect 1976 4336 1983 4413
rect 1956 4267 1963 4303
rect 2036 4267 2043 4333
rect 1956 4187 1963 4253
rect 2136 4167 2143 4413
rect 1773 4040 1787 4053
rect 1776 4036 1783 4040
rect 1736 3816 1743 3933
rect 1756 3867 1763 4003
rect 1820 4003 1833 4007
rect 1816 3993 1833 4003
rect 1876 4003 1883 4023
rect 2136 4007 2143 4053
rect 1856 3996 1883 4003
rect 1716 3607 1723 3770
rect 1616 3516 1623 3593
rect 1696 3487 1703 3516
rect 1596 3387 1603 3483
rect 1636 3480 1643 3483
rect 1633 3467 1647 3480
rect 1376 3227 1383 3263
rect 1636 3227 1643 3263
rect 1276 2996 1283 3032
rect 1216 2960 1223 2963
rect 1213 2947 1227 2960
rect 1076 2220 1083 2223
rect 1116 2220 1123 2223
rect 1073 2207 1087 2220
rect 1113 2207 1127 2220
rect 676 1687 683 1753
rect 676 1507 683 1673
rect 696 1327 703 1993
rect 776 1956 783 1993
rect 1156 1950 1163 2313
rect 1176 2207 1183 2673
rect 1196 2007 1203 2893
rect 1256 2887 1263 2963
rect 1247 2816 1303 2823
rect 1253 2780 1267 2793
rect 1256 2776 1263 2780
rect 1296 2776 1303 2816
rect 1356 2744 1363 2833
rect 1276 2740 1283 2743
rect 1273 2727 1287 2740
rect 1376 2727 1383 3213
rect 1516 2996 1523 3053
rect 1536 2907 1543 2963
rect 1396 2687 1403 2793
rect 1553 2780 1567 2793
rect 1556 2776 1563 2780
rect 1656 2687 1663 3250
rect 1216 2467 1223 2553
rect 1316 2503 1323 2673
rect 1296 2496 1323 2503
rect 1356 2496 1363 2613
rect 1656 2607 1663 2673
rect 1296 2476 1303 2496
rect 1387 2463 1400 2467
rect 1387 2456 1403 2463
rect 1387 2453 1400 2456
rect 1276 2387 1283 2443
rect 1316 2440 1323 2443
rect 1313 2427 1327 2440
rect 1376 2287 1383 2413
rect 1396 2387 1403 2433
rect 1656 2427 1663 2493
rect 1353 2260 1367 2273
rect 1356 2256 1363 2260
rect 1376 2207 1383 2223
rect 756 1736 763 1873
rect 736 1700 743 1703
rect 776 1700 783 1703
rect 733 1687 747 1700
rect 773 1687 787 1700
rect 816 1687 823 1853
rect 876 1667 883 1943
rect 696 1127 703 1313
rect 776 1216 783 1353
rect 816 1227 823 1363
rect 716 943 723 1213
rect 876 1196 883 1473
rect 896 1403 903 1493
rect 916 1449 923 1753
rect 996 1736 1003 1833
rect 1036 1736 1043 1793
rect 976 1367 983 1473
rect 996 1327 1003 1373
rect 1016 1363 1023 1703
rect 1196 1667 1203 1943
rect 1296 1847 1303 2133
rect 1316 1944 1323 2173
rect 1376 2087 1383 2193
rect 1387 2076 1403 2083
rect 1293 1740 1307 1753
rect 1296 1736 1303 1740
rect 1316 1683 1323 1690
rect 1296 1676 1323 1683
rect 1107 1496 1133 1503
rect 1116 1436 1123 1473
rect 1056 1400 1063 1403
rect 1053 1387 1067 1400
rect 1016 1356 1073 1363
rect 1096 1307 1103 1403
rect 1136 1367 1143 1403
rect 1176 1347 1183 1436
rect 1196 1196 1203 1653
rect 1216 1367 1223 1493
rect 1276 1387 1283 1473
rect 756 1180 763 1183
rect 753 1167 767 1180
rect 796 1127 803 1183
rect 836 1087 843 1163
rect 1296 1127 1303 1676
rect 716 936 743 943
rect 736 916 743 936
rect 996 916 1003 953
rect 1256 916 1263 1113
rect 1316 947 1323 1493
rect 1356 1443 1363 2053
rect 1376 1507 1383 1993
rect 1396 1867 1403 2076
rect 1416 1707 1423 2256
rect 1436 2224 1443 2273
rect 1476 2007 1483 2273
rect 1516 2147 1523 2293
rect 1616 2256 1623 2293
rect 1676 2267 1683 3413
rect 1736 3387 1743 3693
rect 1736 3127 1743 3333
rect 1756 3167 1763 3733
rect 1796 3587 1803 3990
rect 1816 3427 1823 3993
rect 1856 3627 1863 3996
rect 1876 3747 1883 3953
rect 2016 3816 2023 3913
rect 1916 3647 1923 3733
rect 1896 3516 1903 3613
rect 1736 2964 1743 3113
rect 1776 2996 1783 3293
rect 1896 3227 1903 3263
rect 1896 3167 1903 3213
rect 1796 2776 1803 2913
rect 1836 2907 1843 2963
rect 1836 2847 1843 2893
rect 1756 2736 1773 2743
rect 1696 2507 1703 2673
rect 1756 2507 1763 2736
rect 1816 2607 1823 2743
rect 1896 2667 1903 3093
rect 1956 2807 1963 3816
rect 1836 2496 1843 2613
rect 1976 2607 1983 3773
rect 1996 3484 2003 3783
rect 1996 2647 2003 2773
rect 2016 2567 2023 3633
rect 2076 2996 2083 3653
rect 2156 3647 2163 4673
rect 2196 4607 2203 4810
rect 2236 4787 2243 4823
rect 2176 4067 2183 4533
rect 2196 4447 2203 4543
rect 2256 4507 2263 4543
rect 2196 4087 2203 4433
rect 2296 4427 2303 4873
rect 2276 4336 2283 4373
rect 2316 4347 2323 4713
rect 2256 4283 2263 4303
rect 2256 4276 2283 4283
rect 2276 4067 2283 4276
rect 2296 4267 2303 4303
rect 2273 4003 2287 4013
rect 2256 4000 2287 4003
rect 2256 3996 2283 4000
rect 2176 3547 2183 3893
rect 2213 3830 2227 3833
rect 2256 3816 2263 3996
rect 2296 3907 2303 4153
rect 2316 3847 2323 4293
rect 2276 3780 2283 3783
rect 2273 3767 2287 3780
rect 2196 3516 2203 3693
rect 2136 3447 2143 3483
rect 2176 3367 2183 3483
rect 2113 3300 2127 3313
rect 2116 3296 2123 3300
rect 2156 3296 2163 3353
rect 2216 3264 2223 3433
rect 2176 3187 2183 3263
rect 2096 2847 2103 2963
rect 2093 2780 2107 2793
rect 2096 2776 2103 2780
rect 2156 2747 2163 2833
rect 2176 2827 2183 2893
rect 2076 2740 2083 2743
rect 2116 2740 2123 2743
rect 2073 2727 2087 2740
rect 2113 2727 2127 2740
rect 2176 2727 2183 2773
rect 2196 2727 2203 3193
rect 1860 2507 1867 2553
rect 2216 2547 2223 3053
rect 2236 2507 2243 3533
rect 2256 3427 2263 3516
rect 2256 2807 2263 3353
rect 2276 2507 2283 3013
rect 2296 2623 2303 3016
rect 2316 3003 2323 3793
rect 2336 3027 2343 5253
rect 2356 4547 2363 4893
rect 2356 4287 2363 4493
rect 2376 4487 2383 5013
rect 2416 4647 2423 5213
rect 2476 5207 2483 5413
rect 2516 5370 2523 6273
rect 2536 5387 2543 6113
rect 2556 5827 2563 6433
rect 2576 6327 2583 6936
rect 2596 6447 2603 7013
rect 2616 6607 2623 6636
rect 2616 6116 2623 6373
rect 2636 6167 2643 7456
rect 2736 7420 2743 7423
rect 2733 7407 2747 7420
rect 2773 7407 2787 7413
rect 2656 7107 2663 7153
rect 2676 7087 2683 7193
rect 2676 6936 2683 6973
rect 2716 6936 2723 7313
rect 2696 6900 2703 6903
rect 2693 6887 2707 6900
rect 2736 6747 2743 6903
rect 2716 6667 2723 6713
rect 2756 6643 2763 6713
rect 2736 6636 2763 6643
rect 2776 6627 2783 7233
rect 2796 6707 2803 7873
rect 2876 7667 2883 7956
rect 2916 7807 2923 8153
rect 2936 8047 2943 8183
rect 2936 7690 2943 7993
rect 2976 7767 2983 8213
rect 2996 7827 3003 8373
rect 3016 7787 3023 8313
rect 3036 8167 3043 8393
rect 3056 8007 3063 8053
rect 3056 7976 3063 7993
rect 2980 7683 2993 7687
rect 2976 7676 2993 7683
rect 2980 7673 2993 7676
rect 2876 7607 2883 7653
rect 2936 7087 2943 7593
rect 3016 7456 3023 7673
rect 2996 7387 3003 7410
rect 2876 7047 2883 7083
rect 2856 6687 2863 6973
rect 2796 6607 2803 6653
rect 2656 6267 2663 6593
rect 2716 6600 2723 6603
rect 2713 6587 2727 6600
rect 2876 6587 2883 6953
rect 2916 6603 2923 7013
rect 2936 6907 2943 7033
rect 2976 7027 2983 7313
rect 2996 6976 3003 7213
rect 3016 7007 3023 7133
rect 3036 7127 3043 7273
rect 3056 6967 3063 7629
rect 3096 7470 3103 7673
rect 3116 7647 3123 8333
rect 3096 7427 3103 7456
rect 3136 7327 3143 8253
rect 3176 8196 3183 8293
rect 3196 8067 3203 8163
rect 3156 7567 3163 7976
rect 3176 7947 3183 8013
rect 3336 7976 3343 8013
rect 3316 7907 3323 7943
rect 3236 7456 3243 7603
rect 2996 6636 3003 6753
rect 2916 6596 2943 6603
rect 2693 6420 2707 6433
rect 2696 6416 2703 6420
rect 2736 6416 2743 6453
rect 2756 6380 2763 6383
rect 2753 6367 2767 6380
rect 2656 6116 2663 6153
rect 2676 6147 2683 6213
rect 2756 6107 2763 6313
rect 2796 6307 2803 6553
rect 2816 6367 2823 6533
rect 2816 6187 2823 6213
rect 2576 5727 2583 5896
rect 2636 5864 2643 6083
rect 2716 5927 2723 5993
rect 2676 5787 2683 5863
rect 2716 5856 2743 5863
rect 2633 5600 2647 5613
rect 2676 5610 2683 5673
rect 2696 5667 2703 5813
rect 2636 5596 2643 5600
rect 2656 5547 2663 5563
rect 2576 5356 2583 5453
rect 2656 5387 2663 5533
rect 2496 5087 2503 5313
rect 2516 5076 2523 5173
rect 2376 4304 2383 4333
rect 2356 4047 2363 4252
rect 2396 4147 2403 4593
rect 2436 4587 2443 5073
rect 2476 4767 2483 4823
rect 2516 4783 2523 4813
rect 2516 4776 2543 4783
rect 2476 4563 2483 4713
rect 2456 4556 2483 4563
rect 2493 4560 2507 4573
rect 2496 4556 2503 4560
rect 2536 4556 2543 4776
rect 2576 4707 2583 4993
rect 2596 4827 2603 5030
rect 2580 4563 2593 4567
rect 2576 4556 2593 4563
rect 2436 4507 2443 4533
rect 2356 3807 2363 4012
rect 2376 3947 2383 4113
rect 2376 3727 2383 3912
rect 2396 3784 2403 4133
rect 2416 3667 2423 4473
rect 2436 3907 2443 4453
rect 2456 4267 2463 4556
rect 2580 4553 2593 4556
rect 2556 4467 2563 4523
rect 2593 4507 2607 4510
rect 2476 4087 2483 4393
rect 2580 4343 2593 4347
rect 2576 4336 2593 4343
rect 2580 4333 2593 4336
rect 2516 4300 2523 4303
rect 2513 4287 2527 4300
rect 2556 4283 2563 4303
rect 2556 4276 2583 4283
rect 2456 3707 2463 3973
rect 2536 3867 2543 4193
rect 2556 4024 2563 4173
rect 2516 3780 2523 3783
rect 2513 3767 2527 3780
rect 2356 3303 2363 3613
rect 2476 3587 2483 3673
rect 2576 3607 2583 4276
rect 2453 3520 2467 3533
rect 2456 3516 2463 3520
rect 2436 3427 2443 3483
rect 2356 3296 2383 3303
rect 2413 3300 2427 3313
rect 2416 3296 2423 3300
rect 2436 3087 2443 3263
rect 2476 3107 2483 3293
rect 2496 3264 2503 3513
rect 2516 3187 2523 3553
rect 2596 3207 2603 4193
rect 2616 4050 2623 5373
rect 2636 5127 2643 5353
rect 2636 4407 2643 4873
rect 2656 4387 2663 5373
rect 2676 5227 2683 5413
rect 2676 5007 2683 5133
rect 2696 5007 2703 5553
rect 2636 4287 2643 4353
rect 2656 4307 2663 4333
rect 2676 4267 2683 4893
rect 2696 4667 2703 4993
rect 2696 4307 2703 4493
rect 2636 4036 2643 4073
rect 2616 3727 2623 3816
rect 2676 3567 2683 4113
rect 2696 3927 2703 4293
rect 2716 4167 2723 5833
rect 2736 5827 2743 5856
rect 2736 5167 2743 5653
rect 2736 4927 2743 5113
rect 2756 4887 2763 6033
rect 2776 5610 2783 5993
rect 2796 5864 2803 5893
rect 2796 5627 2803 5813
rect 2816 5687 2823 6173
rect 2836 6067 2843 6416
rect 2796 5376 2803 5413
rect 2816 5403 2823 5613
rect 2836 5427 2843 6053
rect 2856 5767 2863 6313
rect 2876 6187 2883 6573
rect 2916 6467 2923 6493
rect 2936 6327 2943 6596
rect 2976 6547 2983 6603
rect 3036 6507 3043 6636
rect 2996 6327 3003 6370
rect 2987 6213 2993 6227
rect 2913 6120 2927 6133
rect 2916 6116 2923 6120
rect 2856 5647 2863 5753
rect 2876 5603 2883 5913
rect 2896 5787 2903 6083
rect 2936 6080 2943 6083
rect 2933 6067 2947 6080
rect 3016 6067 3023 6333
rect 2936 5896 2943 5933
rect 3036 5864 3043 6173
rect 3056 6007 3063 6273
rect 3076 6227 3083 7273
rect 3133 7160 3147 7173
rect 3136 7156 3143 7160
rect 3116 6687 3123 7123
rect 3216 7107 3223 7156
rect 3316 7127 3323 7713
rect 3336 7689 3343 7913
rect 3336 7647 3343 7675
rect 3336 7424 3343 7633
rect 3356 7387 3363 7456
rect 3136 6927 3143 7073
rect 3076 5963 3083 6173
rect 3056 5956 3083 5963
rect 2996 5856 3023 5863
rect 2856 5596 2883 5603
rect 2956 5596 2963 5633
rect 2856 5427 2863 5596
rect 2896 5487 2903 5563
rect 2936 5560 2943 5563
rect 2933 5547 2947 5560
rect 2973 5547 2987 5553
rect 2936 5487 2943 5512
rect 2816 5396 2843 5403
rect 2836 5376 2843 5396
rect 2856 5340 2863 5343
rect 2853 5327 2867 5340
rect 2816 5207 2823 5233
rect 2796 5147 2803 5173
rect 2793 5080 2807 5093
rect 2873 5090 2887 5093
rect 2796 5076 2803 5080
rect 2856 4870 2863 5030
rect 2756 4767 2763 4823
rect 2736 4647 2743 4733
rect 2756 4727 2763 4753
rect 2796 4727 2803 4823
rect 2696 3547 2703 3653
rect 2716 3587 2723 4073
rect 2736 3830 2743 4633
rect 2756 4407 2763 4613
rect 2856 4556 2863 4813
rect 2876 4727 2883 5033
rect 2896 4570 2903 5413
rect 2936 5347 2943 5373
rect 2916 4627 2923 5093
rect 2936 5027 2943 5312
rect 2976 5267 2983 5330
rect 2956 5067 2963 5133
rect 2936 4807 2943 4913
rect 2956 4767 2963 5053
rect 2776 4507 2783 4553
rect 2793 4507 2807 4513
rect 2836 4487 2843 4523
rect 2893 4483 2907 4493
rect 2876 4480 2907 4483
rect 2876 4476 2903 4480
rect 2876 4403 2883 4476
rect 2916 4467 2923 4510
rect 2856 4396 2883 4403
rect 2773 4340 2787 4353
rect 2816 4343 2823 4393
rect 2776 4336 2783 4340
rect 2816 4336 2843 4343
rect 2796 4267 2803 4303
rect 2813 4287 2827 4293
rect 2776 4004 2783 4053
rect 2796 3827 2803 4253
rect 2836 4207 2843 4336
rect 2856 4127 2863 4396
rect 2696 3516 2703 3533
rect 2736 3530 2743 3613
rect 2756 3547 2763 3783
rect 2776 3527 2783 3613
rect 2716 3447 2723 3483
rect 2636 3264 2643 3313
rect 2716 3310 2723 3353
rect 2736 3227 2743 3263
rect 2596 3147 2603 3193
rect 2776 3107 2783 3296
rect 2316 2996 2343 3003
rect 2356 2907 2363 2963
rect 2416 2867 2423 2973
rect 2436 2887 2443 2953
rect 2393 2780 2407 2793
rect 2396 2776 2403 2780
rect 2327 2743 2340 2747
rect 2456 2744 2463 2893
rect 2327 2736 2343 2743
rect 2327 2733 2340 2736
rect 2376 2707 2383 2743
rect 2476 2707 2483 2983
rect 2756 2923 2763 3073
rect 2796 3047 2803 3253
rect 2816 3027 2823 4073
rect 2876 4067 2883 4373
rect 2896 4187 2903 4353
rect 2916 4267 2923 4393
rect 2936 4087 2943 4733
rect 2956 4003 2963 4693
rect 2976 4667 2983 5253
rect 2996 4907 3003 5793
rect 3016 5527 3023 5856
rect 3036 5463 3043 5850
rect 3056 5807 3063 5956
rect 3056 5567 3063 5772
rect 3076 5727 3083 5933
rect 3076 5647 3083 5713
rect 3096 5610 3103 6413
rect 3116 6187 3123 6613
rect 3136 6207 3143 6913
rect 3156 6487 3163 6813
rect 3176 6607 3183 7093
rect 3256 6936 3263 6993
rect 3296 6936 3303 6973
rect 3336 6807 3343 7013
rect 3356 6767 3363 7253
rect 3376 6787 3383 8476
rect 3396 7807 3403 8433
rect 3436 8220 3473 8223
rect 3433 8216 3473 8220
rect 3433 8210 3447 8216
rect 3446 8200 3447 8210
rect 3476 8156 3503 8163
rect 3456 7607 3463 8073
rect 3476 7527 3483 8113
rect 3496 7927 3503 8156
rect 3516 7747 3523 8513
rect 3536 8087 3543 8813
rect 3556 8647 3563 8953
rect 3556 8267 3563 8633
rect 3576 8427 3583 8716
rect 3596 8307 3603 8833
rect 3616 8167 3623 8773
rect 3636 8127 3643 9073
rect 3716 8987 3723 9193
rect 3736 9043 3743 9216
rect 3736 9036 3763 9043
rect 3716 8947 3723 8973
rect 3736 8716 3743 8953
rect 3756 8927 3763 9036
rect 3776 8967 3783 9213
rect 3816 9147 3823 9223
rect 3816 9103 3823 9133
rect 3796 9096 3823 9103
rect 3796 9007 3803 9096
rect 3836 9087 3843 9213
rect 3876 9167 3883 9223
rect 3876 9047 3883 9153
rect 3916 9127 3923 9473
rect 3936 9367 3943 9503
rect 4076 9427 4083 9743
rect 4356 9667 4363 9793
rect 4376 9736 4403 9743
rect 4276 9536 4283 9633
rect 4376 9607 4383 9736
rect 4396 9667 4403 9713
rect 4516 9627 4523 9993
rect 4216 9407 4223 9503
rect 4256 9407 4263 9503
rect 4236 9256 4243 9313
rect 3936 9227 3943 9253
rect 4296 9227 4303 9313
rect 3976 8996 3983 9033
rect 3776 8787 3783 8932
rect 3796 8887 3803 8972
rect 3816 8947 3823 8973
rect 3876 8947 3883 8983
rect 3836 8887 3843 8933
rect 3796 8807 3803 8873
rect 3773 8720 3787 8733
rect 3776 8716 3783 8720
rect 3716 8527 3723 8683
rect 3733 8500 3747 8513
rect 3736 8496 3743 8500
rect 3693 8210 3707 8213
rect 3596 7976 3603 8073
rect 3676 8047 3683 8163
rect 3636 7990 3643 8033
rect 3536 7676 3543 7976
rect 3676 7943 3683 7993
rect 3576 7940 3583 7943
rect 3616 7940 3623 7943
rect 3573 7927 3587 7940
rect 3613 7927 3627 7940
rect 3656 7936 3683 7943
rect 3576 7676 3583 7733
rect 3500 7423 3513 7427
rect 3496 7416 3513 7423
rect 3500 7413 3513 7416
rect 3413 7160 3427 7173
rect 3416 7156 3423 7160
rect 3276 6667 3283 6713
rect 3273 6640 3287 6653
rect 3276 6636 3283 6640
rect 3316 6627 3323 6713
rect 3256 6600 3263 6603
rect 3253 6587 3267 6600
rect 3156 6384 3163 6413
rect 3176 6347 3183 6493
rect 3156 6247 3163 6313
rect 3156 6116 3163 6233
rect 3216 6147 3223 6433
rect 3256 6416 3263 6473
rect 3293 6420 3307 6433
rect 3296 6416 3303 6420
rect 3276 6247 3283 6383
rect 3316 6380 3323 6383
rect 3313 6367 3327 6380
rect 3076 5507 3083 5573
rect 3116 5547 3123 6073
rect 3136 5807 3143 6083
rect 3156 5727 3163 6033
rect 3176 5827 3183 6083
rect 3256 6007 3263 6116
rect 3276 6047 3283 6233
rect 3253 5927 3267 5933
rect 3253 5900 3267 5913
rect 3296 5907 3303 6353
rect 3316 5947 3323 6133
rect 3356 6047 3363 6636
rect 3256 5896 3263 5900
rect 3236 5843 3243 5863
rect 3216 5840 3243 5843
rect 3213 5836 3243 5840
rect 3213 5827 3227 5836
rect 3136 5547 3143 5633
rect 3196 5596 3203 5713
rect 3276 5707 3283 5850
rect 3256 5607 3263 5673
rect 3316 5647 3323 5933
rect 3356 5747 3363 5913
rect 3167 5563 3180 5567
rect 3167 5556 3183 5563
rect 3167 5553 3180 5556
rect 3036 5456 3063 5463
rect 3016 4967 3023 5373
rect 3036 5043 3043 5433
rect 3056 5107 3063 5456
rect 3116 5376 3123 5512
rect 3167 5376 3173 5387
rect 3160 5373 3173 5376
rect 3076 5307 3083 5333
rect 3096 5207 3103 5343
rect 3136 5247 3143 5343
rect 3093 5080 3107 5093
rect 3096 5076 3103 5080
rect 3036 5036 3083 5043
rect 3087 5013 3093 5027
rect 3116 4927 3123 5043
rect 2916 3947 2923 4003
rect 2936 3996 2963 4003
rect 2836 3827 2843 3853
rect 2876 3267 2883 3816
rect 2916 3484 2923 3813
rect 2936 3687 2943 3996
rect 2976 3947 2983 4553
rect 2996 4303 3003 4856
rect 3136 4823 3143 4853
rect 3016 4687 3023 4793
rect 3036 4787 3043 4823
rect 3096 4816 3143 4823
rect 3156 4767 3163 4933
rect 3176 4767 3183 5273
rect 3196 5067 3203 5353
rect 3216 4927 3223 5529
rect 3247 5373 3253 5387
rect 3236 5007 3243 5233
rect 3256 4947 3263 5113
rect 3036 4527 3043 4633
rect 3056 4507 3063 4556
rect 3096 4507 3103 4753
rect 3196 4743 3203 4793
rect 3176 4736 3203 4743
rect 3176 4556 3183 4736
rect 3216 4607 3223 4773
rect 3216 4556 3223 4593
rect 3016 4347 3023 4493
rect 3053 4340 3067 4353
rect 3096 4350 3103 4453
rect 3056 4336 3063 4340
rect 2996 4296 3023 4303
rect 2996 4147 3003 4273
rect 3016 4247 3023 4296
rect 3076 4283 3083 4303
rect 3056 4276 3083 4283
rect 3056 4247 3063 4276
rect 2956 3887 2963 3933
rect 3016 3847 3023 4153
rect 3053 4147 3067 4153
rect 3036 4027 3043 4133
rect 3056 4007 3063 4036
rect 3056 3887 3063 3933
rect 3013 3820 3027 3833
rect 3016 3816 3023 3820
rect 2996 3747 3003 3783
rect 3036 3780 3043 3783
rect 3033 3767 3047 3780
rect 2936 3483 2943 3673
rect 2976 3627 2983 3653
rect 2976 3516 2983 3613
rect 2936 3476 2963 3483
rect 2956 3296 2963 3476
rect 2936 3243 2943 3263
rect 2936 3236 2963 3243
rect 2796 2947 2803 2983
rect 2896 2983 2903 3153
rect 2856 2976 2903 2983
rect 2756 2916 2783 2923
rect 2756 2867 2763 2893
rect 2680 2803 2693 2807
rect 2676 2793 2693 2803
rect 2676 2776 2683 2793
rect 2296 2616 2313 2623
rect 2316 2496 2323 2613
rect 2336 2507 2343 2593
rect 2716 2507 2723 2813
rect 2756 2503 2763 2832
rect 2776 2807 2783 2916
rect 2796 2827 2803 2933
rect 2776 2744 2783 2793
rect 2756 2496 2783 2503
rect 1716 2327 1723 2463
rect 2136 2427 2143 2493
rect 2056 2267 2063 2313
rect 2156 2287 2163 2493
rect 2196 2460 2223 2463
rect 2196 2456 2227 2460
rect 2053 2240 2067 2253
rect 2156 2250 2163 2273
rect 2056 2236 2063 2240
rect 1636 2187 1643 2223
rect 1656 2147 1663 2213
rect 1476 1956 1483 1993
rect 1696 1990 1703 2203
rect 2016 2127 2023 2230
rect 1596 1776 1603 1956
rect 1676 1907 1683 1973
rect 1656 1743 1663 1813
rect 1647 1737 1663 1743
rect 1636 1736 1663 1737
rect 1336 1436 1363 1443
rect 1316 916 1323 933
rect 1336 930 1343 1436
rect 1416 1400 1423 1403
rect 1413 1387 1427 1400
rect 1356 1007 1363 1373
rect 1447 1353 1453 1367
rect 1496 1347 1503 1693
rect 1536 1447 1543 1633
rect 1496 1216 1503 1333
rect 1516 1327 1523 1353
rect 1536 1207 1543 1433
rect 1556 1387 1563 1593
rect 1596 1196 1603 1553
rect 1676 1436 1683 1773
rect 1696 1647 1703 1976
rect 1733 1960 1747 1973
rect 1736 1956 1743 1960
rect 1796 1956 1803 2113
rect 2036 2087 2043 2193
rect 1956 1927 1963 1956
rect 1716 1436 1723 1473
rect 1656 1400 1663 1403
rect 1653 1387 1667 1400
rect 1756 1387 1763 1893
rect 1776 1887 1783 1923
rect 1976 1924 1983 1993
rect 2036 1956 2043 2033
rect 2176 1927 2183 2456
rect 2213 2447 2227 2456
rect 1896 1507 1903 1703
rect 1956 1467 1963 1693
rect 1956 1436 1963 1453
rect 1996 1436 2003 1493
rect 2036 1347 2043 1733
rect 2056 1704 2063 1733
rect 2056 1404 2063 1433
rect 2036 1267 2043 1333
rect 1916 1196 1923 1253
rect 2076 1230 2083 1833
rect 2096 1747 2103 1893
rect 2196 1847 2203 2413
rect 2216 2267 2223 2433
rect 2216 1907 2223 2253
rect 2256 2147 2263 2463
rect 2276 1963 2283 2453
rect 2336 2327 2343 2453
rect 2356 2287 2363 2463
rect 2376 2427 2383 2456
rect 2616 2423 2623 2473
rect 2636 2464 2643 2493
rect 2736 2460 2743 2463
rect 2733 2447 2747 2460
rect 2616 2416 2643 2423
rect 2296 2147 2303 2273
rect 2333 2260 2347 2273
rect 2336 2256 2343 2260
rect 2356 2203 2363 2223
rect 2356 2196 2383 2203
rect 2256 1956 2283 1963
rect 2296 1956 2303 2013
rect 2376 1970 2383 2196
rect 2396 2187 2403 2253
rect 2476 1970 2483 2313
rect 2156 1787 2163 1813
rect 2136 1736 2143 1773
rect 2156 1700 2163 1703
rect 2153 1687 2167 1700
rect 2216 1687 2223 1853
rect 2236 1707 2243 1736
rect 2256 1467 2263 1956
rect 2376 1924 2383 1956
rect 2316 1920 2323 1923
rect 2313 1907 2327 1920
rect 1973 1200 1987 1213
rect 1976 1196 1983 1200
rect 1556 1087 1563 1150
rect 696 696 703 853
rect 716 747 723 883
rect 756 847 763 883
rect 1056 884 1063 913
rect 636 664 643 693
rect 716 660 723 663
rect 713 647 727 660
rect 756 647 763 833
rect 516 507 523 593
rect 136 384 143 493
rect 456 416 463 493
rect 36 287 43 383
rect 496 387 503 473
rect 696 396 703 453
rect 396 347 403 376
rect 716 360 723 363
rect 713 347 727 360
rect 796 347 803 873
rect 1016 767 1023 883
rect 1296 807 1303 883
rect 1356 807 1363 883
rect 996 696 1003 733
rect 956 447 963 663
rect 1016 660 1023 663
rect 1013 647 1027 660
rect 1056 647 1063 793
rect 1076 507 1083 753
rect 1296 727 1303 793
rect 1256 696 1303 703
rect 1236 507 1243 663
rect 1296 627 1303 696
rect 896 364 903 433
rect 196 176 203 273
rect 756 247 763 333
rect 456 -24 463 143
rect 496 140 503 143
rect 493 127 507 140
rect 536 127 543 233
rect 716 190 723 233
rect 756 176 763 233
rect 676 107 683 173
rect 776 107 783 143
rect 816 107 823 176
rect 916 144 923 333
rect 1076 176 1083 493
rect 1176 396 1183 453
rect 1213 400 1227 413
rect 1216 396 1223 400
rect 1016 107 1023 143
rect 1116 107 1123 193
rect 1176 47 1183 233
rect 1213 187 1227 193
rect 1236 127 1243 363
rect 1276 327 1283 413
rect 1356 407 1363 433
rect 1456 407 1463 993
rect 1536 747 1543 933
rect 1636 916 1643 993
rect 1876 987 1883 1173
rect 2156 1147 2163 1453
rect 2296 1404 2303 1853
rect 2376 1736 2383 1910
rect 2413 1740 2427 1753
rect 2416 1736 2423 1740
rect 1576 807 1583 883
rect 1836 847 1843 973
rect 1933 920 1947 933
rect 1936 916 1943 920
rect 1996 884 2003 993
rect 2096 887 2103 916
rect 1916 847 1923 883
rect 1493 700 1507 713
rect 1496 696 1503 700
rect 1536 696 1543 733
rect 1467 396 1483 403
rect 1516 396 1523 433
rect 1256 187 1263 253
rect 1293 180 1307 193
rect 1296 176 1303 180
rect 1336 176 1343 213
rect 1376 207 1383 393
rect 1576 364 1583 693
rect 1776 567 1783 650
rect 1756 396 1763 453
rect 1796 396 1803 533
rect 1816 507 1823 663
rect 1496 307 1503 363
rect 1736 267 1743 363
rect 1776 327 1783 363
rect 1376 176 1383 193
rect 1256 107 1263 152
rect 1756 163 1763 293
rect 1796 163 1803 293
rect 1856 183 1863 733
rect 1996 190 2003 870
rect 2076 807 2083 853
rect 2036 696 2043 793
rect 2116 727 2123 993
rect 2156 916 2163 953
rect 2196 916 2203 993
rect 2216 947 2223 1183
rect 2176 827 2183 883
rect 2073 700 2087 713
rect 2076 696 2083 700
rect 2056 627 2063 663
rect 2036 396 2043 493
rect 2156 467 2163 773
rect 2176 664 2183 813
rect 2076 396 2083 453
rect 2096 227 2103 350
rect 2116 247 2123 273
rect 1736 156 1763 163
rect 1776 156 1803 163
rect 1836 176 1863 183
rect 1836 156 1843 176
rect 1316 140 1323 143
rect 1273 127 1287 133
rect 1313 127 1327 140
rect 1736 107 1743 156
rect 2016 144 2023 213
rect 2196 167 2203 413
rect 2216 156 2223 433
rect 2236 364 2243 393
rect 2276 367 2283 1333
rect 2316 1267 2323 1433
rect 2336 696 2343 915
rect 2376 747 2383 1453
rect 2396 1427 2403 1690
rect 2496 1607 2503 2333
rect 2636 2307 2643 2416
rect 2656 2307 2663 2393
rect 2756 2347 2763 2453
rect 2516 2027 2523 2293
rect 2633 2260 2647 2272
rect 2636 2256 2643 2260
rect 2656 2220 2663 2223
rect 2653 2207 2667 2220
rect 2616 1956 2623 2153
rect 2476 1436 2483 1513
rect 2516 1404 2523 1613
rect 2396 1087 2403 1353
rect 2436 1216 2443 1253
rect 2316 567 2323 663
rect 2356 627 2363 650
rect 2336 410 2343 453
rect 2396 430 2403 1073
rect 2516 1047 2523 1390
rect 2536 1127 2543 1753
rect 2676 1736 2683 1813
rect 2716 1747 2723 2273
rect 2776 2207 2783 2496
rect 2796 2224 2803 2773
rect 2776 2127 2783 2193
rect 2816 1967 2823 2973
rect 2916 2927 2923 3113
rect 2856 2847 2863 2913
rect 2873 2780 2887 2793
rect 2876 2776 2883 2780
rect 2916 2776 2923 2833
rect 2836 1990 2843 2773
rect 2956 2767 2963 3236
rect 2996 3010 3003 3483
rect 3036 2947 3043 3053
rect 3076 3003 3083 4253
rect 3096 3923 3103 4113
rect 3116 4087 3123 4303
rect 3176 4127 3183 4353
rect 3196 4350 3203 4523
rect 3196 4207 3203 4336
rect 3136 3967 3143 4003
rect 3236 4003 3243 4513
rect 3256 4507 3263 4912
rect 3276 4527 3283 5596
rect 3296 5090 3303 5613
rect 3316 5564 3323 5633
rect 3356 5507 3363 5593
rect 3316 5347 3323 5413
rect 3356 5376 3363 5493
rect 3376 5467 3383 6773
rect 3396 6367 3403 7113
rect 3536 7124 3543 7513
rect 3396 6123 3403 6193
rect 3416 6147 3423 6573
rect 3436 6287 3443 7110
rect 3476 6767 3483 6853
rect 3496 6807 3503 7113
rect 3556 7027 3563 7453
rect 3576 7107 3583 7593
rect 3616 7547 3623 7653
rect 3596 6987 3603 7453
rect 3636 7207 3643 7753
rect 3656 7407 3663 7936
rect 3676 7207 3683 7513
rect 3696 7467 3703 8113
rect 3716 7927 3723 8163
rect 3716 7587 3723 7913
rect 3756 7847 3763 8413
rect 3716 7467 3723 7573
rect 3756 7456 3763 7812
rect 3796 7727 3803 8149
rect 3816 7690 3823 8493
rect 3836 8007 3843 8852
rect 3896 8747 3903 8953
rect 3936 8767 3943 8953
rect 3956 8647 3963 8953
rect 4016 8867 4023 9113
rect 4036 9007 4043 9033
rect 4296 8996 4303 9213
rect 4316 9007 4323 9190
rect 4336 9167 4343 9333
rect 4356 9047 4363 9553
rect 4376 9207 4383 9453
rect 4396 9267 4403 9513
rect 4416 9327 4423 9413
rect 4476 9307 4483 9353
rect 4496 9347 4503 9503
rect 4536 9347 4543 9833
rect 4556 9487 4563 9993
rect 4636 9987 4643 10633
rect 4576 9527 4583 9753
rect 4416 9203 4423 9292
rect 4476 9236 4483 9293
rect 4496 9287 4503 9333
rect 4576 9207 4583 9236
rect 4596 9207 4603 9973
rect 4656 9767 4663 10593
rect 4716 10527 4723 10776
rect 4756 10627 4763 10776
rect 4836 10687 4843 10770
rect 4816 10576 4823 10633
rect 4836 10587 4843 10673
rect 4747 10543 4760 10547
rect 4856 10544 4863 10953
rect 4747 10536 4763 10543
rect 4747 10533 4760 10536
rect 4676 10127 4683 10213
rect 4676 9847 4683 10113
rect 4696 10027 4703 10493
rect 4716 10427 4723 10513
rect 4876 10387 4883 10793
rect 4756 10276 4763 10373
rect 4827 10353 4833 10367
rect 4716 10007 4723 10233
rect 4736 9947 4743 10243
rect 4776 10187 4783 10243
rect 4876 10167 4883 10313
rect 4716 9756 4723 9793
rect 4756 9787 4763 10013
rect 4776 9907 4783 10053
rect 4896 10047 4903 11096
rect 4916 10507 4923 11193
rect 4996 11096 5003 11196
rect 5036 11096 5043 11173
rect 4976 11060 4983 11063
rect 4973 11047 4987 11060
rect 5016 11027 5023 11063
rect 5056 11007 5063 11050
rect 5076 10967 5083 11213
rect 4936 10367 4943 10873
rect 4956 10607 4963 10813
rect 5036 10796 5043 10873
rect 5096 10827 5103 11193
rect 5116 11067 5123 11336
rect 4956 10527 4963 10572
rect 4976 10367 4983 10633
rect 5033 10580 5047 10593
rect 5036 10576 5043 10580
rect 5016 10540 5023 10543
rect 5013 10527 5027 10540
rect 4936 10227 4943 10276
rect 4956 10036 4963 10313
rect 4976 10244 4983 10353
rect 5036 10276 5043 10513
rect 5056 10487 5063 10543
rect 5096 10507 5103 10543
rect 5136 10487 5143 10713
rect 5156 10607 5163 10933
rect 5156 10147 5163 10572
rect 5176 10507 5183 11413
rect 5196 11063 5203 11393
rect 5316 11387 5323 11433
rect 5316 11316 5323 11373
rect 5356 11316 5363 11353
rect 5396 11283 5403 11616
rect 5236 11110 5243 11253
rect 5196 11056 5223 11063
rect 5196 10707 5203 11013
rect 5216 10807 5223 11056
rect 5256 10764 5263 10953
rect 5336 10927 5343 11283
rect 5376 11276 5403 11283
rect 5356 10967 5363 11133
rect 5376 10987 5383 11276
rect 5396 11007 5403 11050
rect 5296 10796 5303 10833
rect 5356 10823 5363 10913
rect 5336 10816 5363 10823
rect 5336 10810 5343 10816
rect 5396 10787 5403 10993
rect 5196 10387 5203 10693
rect 5216 10167 5223 10413
rect 5236 10307 5243 10533
rect 4753 9760 4767 9773
rect 4756 9756 4763 9760
rect 4636 9687 4643 9753
rect 4816 9727 4823 10010
rect 4856 9967 4863 10023
rect 4636 9487 4643 9503
rect 4636 9367 4643 9473
rect 4696 9287 4703 9433
rect 4776 9427 4783 9653
rect 4796 9607 4803 9633
rect 4796 9507 4803 9593
rect 4416 9196 4443 9203
rect 4436 8996 4443 9196
rect 4496 9200 4503 9203
rect 4493 9187 4507 9200
rect 4556 9107 4563 9153
rect 4696 9107 4703 9273
rect 4796 9250 4803 9393
rect 4816 9367 4823 9513
rect 4836 9243 4843 9693
rect 4856 9667 4863 9713
rect 4876 9687 4883 9756
rect 4896 9567 4903 9993
rect 4916 9667 4923 10003
rect 5236 9907 5243 10293
rect 5256 10247 5263 10750
rect 5276 10590 5283 10633
rect 5336 10627 5343 10673
rect 5356 10667 5363 10763
rect 5416 10647 5423 11433
rect 5436 11207 5443 11453
rect 5456 11367 5463 11593
rect 5456 11187 5463 11316
rect 5476 11227 5483 11570
rect 5496 11187 5503 11673
rect 5656 11667 5663 11810
rect 5696 11787 5703 11810
rect 5516 11267 5523 11493
rect 5676 11467 5683 11753
rect 5756 11707 5763 11823
rect 5816 11727 5823 11823
rect 5876 11787 5883 11823
rect 5816 11584 5823 11713
rect 5896 11616 5903 11816
rect 5916 11723 5923 11913
rect 6236 11856 6243 11933
rect 5936 11807 5943 11853
rect 5916 11716 5943 11723
rect 5936 11630 5943 11716
rect 5836 11567 5843 11613
rect 5876 11580 5883 11583
rect 5873 11567 5887 11580
rect 5856 11447 5863 11473
rect 5656 11287 5663 11413
rect 5836 11316 5843 11353
rect 5696 11287 5703 11316
rect 5916 11287 5923 11583
rect 5556 11280 5563 11283
rect 5553 11267 5567 11280
rect 5436 10887 5443 11096
rect 5276 10487 5283 10576
rect 5416 10544 5423 10612
rect 5336 10276 5343 10473
rect 5256 10044 5263 10093
rect 5276 10036 5283 10153
rect 5296 10047 5303 10230
rect 5336 10147 5343 10173
rect 5336 10036 5343 10133
rect 4996 9756 5003 9893
rect 4916 9536 4923 9613
rect 4976 9607 4983 9723
rect 5076 9627 5083 9753
rect 5196 9647 5203 9793
rect 5216 9724 5223 9853
rect 5256 9756 5263 9833
rect 5296 9756 5303 9793
rect 5336 9787 5343 9833
rect 5336 9756 5343 9773
rect 5276 9543 5283 9633
rect 5296 9587 5303 9613
rect 5316 9567 5323 9710
rect 5256 9536 5283 9543
rect 4876 9383 4883 9490
rect 5256 9487 5263 9536
rect 5356 9523 5363 9553
rect 5376 9547 5383 10373
rect 5396 9587 5403 10353
rect 5356 9516 5383 9523
rect 4956 9427 4963 9483
rect 5276 9447 5283 9516
rect 4876 9376 4903 9383
rect 4836 9236 4863 9243
rect 4716 9147 4723 9236
rect 4707 9096 4723 9103
rect 4173 8883 4187 8893
rect 4173 8880 4203 8883
rect 4176 8876 4203 8880
rect 3996 8730 4003 8773
rect 4036 8716 4043 8753
rect 3876 7976 3883 8433
rect 3896 8047 3903 8613
rect 3916 8467 3923 8593
rect 3947 8513 3953 8527
rect 3973 8500 3987 8513
rect 3976 8496 3983 8500
rect 4016 8496 4023 8533
rect 4096 8476 4103 8833
rect 4156 8730 4163 8813
rect 4156 8607 4163 8716
rect 4176 8627 4183 8773
rect 4196 8647 4203 8876
rect 4316 8827 4323 8953
rect 4336 8887 4343 8963
rect 4376 8956 4403 8963
rect 4336 8687 4343 8716
rect 4236 8680 4243 8683
rect 4233 8667 4247 8680
rect 4276 8647 4283 8683
rect 3956 8460 3963 8463
rect 3953 8447 3967 8460
rect 3916 7990 3923 8293
rect 3996 8267 4003 8463
rect 4056 8407 4063 8443
rect 4376 8407 4383 8956
rect 4716 8907 4723 9096
rect 4736 9007 4743 9193
rect 4776 9127 4783 9153
rect 4756 8996 4763 9093
rect 4813 9000 4827 9013
rect 4816 8996 4823 9000
rect 4856 8967 4863 9236
rect 4416 8587 4423 8893
rect 4516 8716 4523 8753
rect 4596 8683 4603 8813
rect 4576 8676 4603 8683
rect 4416 8507 4423 8573
rect 4416 8476 4423 8493
rect 4436 8484 4443 8573
rect 4476 8476 4483 8593
rect 4036 8207 4043 8253
rect 3956 7944 3963 8073
rect 3996 8007 4003 8123
rect 3856 7907 3863 7943
rect 3856 7676 3863 7733
rect 3796 7527 3803 7643
rect 3836 7567 3843 7643
rect 3796 7456 3843 7463
rect 3727 7423 3740 7427
rect 3727 7416 3743 7423
rect 3727 7413 3740 7416
rect 3676 7183 3683 7193
rect 3656 7176 3683 7183
rect 3656 7156 3663 7176
rect 3627 7123 3640 7127
rect 3627 7116 3643 7123
rect 3676 7120 3683 7123
rect 3627 7113 3640 7116
rect 3673 7107 3687 7120
rect 3616 6947 3623 6993
rect 3636 6951 3643 7093
rect 3600 6943 3613 6947
rect 3596 6936 3613 6943
rect 3600 6933 3613 6936
rect 3516 6667 3523 6893
rect 3536 6867 3543 6903
rect 3456 6367 3463 6653
rect 3536 6636 3543 6773
rect 3516 6583 3523 6603
rect 3496 6576 3523 6583
rect 3496 6367 3503 6576
rect 3576 6567 3583 6793
rect 3596 6727 3603 6793
rect 3516 6247 3523 6553
rect 3596 6507 3603 6613
rect 3616 6567 3623 6693
rect 3636 6587 3643 6937
rect 3656 6904 3663 6973
rect 3656 6727 3663 6833
rect 3556 6347 3563 6383
rect 3396 6116 3423 6123
rect 3453 6120 3467 6133
rect 3456 6116 3463 6120
rect 3436 6027 3443 6083
rect 3476 6080 3483 6083
rect 3473 6067 3487 6080
rect 3507 6013 3513 6027
rect 3436 5927 3443 6013
rect 3496 5896 3503 5973
rect 3536 5896 3543 6053
rect 3553 6027 3567 6033
rect 3396 5383 3403 5733
rect 3416 5687 3423 5893
rect 3556 5856 3583 5863
rect 3416 5487 3423 5673
rect 3536 5647 3543 5813
rect 3556 5767 3563 5793
rect 3476 5596 3483 5633
rect 3513 5607 3527 5613
rect 3396 5376 3423 5383
rect 3396 5187 3403 5213
rect 3416 5167 3423 5376
rect 3436 5127 3443 5553
rect 3456 5447 3463 5513
rect 3456 5127 3463 5433
rect 3476 5263 3483 5473
rect 3476 5256 3503 5263
rect 3436 5083 3443 5113
rect 3416 5076 3443 5083
rect 3316 4907 3323 5076
rect 3356 5027 3363 5043
rect 3347 5016 3363 5027
rect 3347 5013 3360 5016
rect 3396 4867 3403 5030
rect 3456 4967 3463 5092
rect 3376 4856 3393 4863
rect 3296 4816 3313 4823
rect 3296 4483 3303 4816
rect 3276 4476 3303 4483
rect 3276 4367 3283 4476
rect 3276 4067 3283 4332
rect 3216 3996 3243 4003
rect 3096 3916 3123 3923
rect 3096 3727 3103 3893
rect 3096 3367 3103 3516
rect 3116 3127 3123 3916
rect 3136 3167 3143 3913
rect 3216 3687 3223 3996
rect 3256 3847 3263 3973
rect 3276 3947 3283 4032
rect 3276 3816 3283 3893
rect 3296 3847 3303 4453
rect 3316 4347 3323 4753
rect 3356 4727 3363 4823
rect 3416 4787 3423 4833
rect 3476 4824 3483 5153
rect 3496 5147 3503 5256
rect 3413 4767 3427 4773
rect 3456 4747 3463 4773
rect 3416 4556 3423 4713
rect 3496 4567 3503 5112
rect 3336 4336 3343 4393
rect 3376 4336 3383 4556
rect 3416 4387 3423 4493
rect 3416 4336 3423 4373
rect 3356 4187 3363 4303
rect 3316 3827 3323 4073
rect 3256 3627 3263 3783
rect 3287 3763 3300 3767
rect 3287 3753 3293 3763
rect 3156 3567 3163 3613
rect 3273 3520 3287 3533
rect 3276 3516 3283 3520
rect 3156 3207 3163 3513
rect 3316 3487 3323 3613
rect 3056 2996 3083 3003
rect 3156 2996 3163 3193
rect 3196 3007 3203 3093
rect 2976 2807 2983 2853
rect 2976 2756 2983 2793
rect 3016 2767 3023 2873
rect 3036 2756 3043 2933
rect 3056 2787 3063 2996
rect 3096 2863 3103 2963
rect 3136 2960 3143 2963
rect 3133 2947 3147 2960
rect 3196 2947 3203 2993
rect 3276 2887 3283 3293
rect 3336 2927 3343 4053
rect 3356 3784 3363 3813
rect 3356 3127 3363 3573
rect 3376 3530 3383 4213
rect 3396 4127 3403 4290
rect 3456 4036 3463 4173
rect 3476 4087 3483 4523
rect 3496 4227 3503 4513
rect 3516 4267 3523 5193
rect 3536 5167 3543 5633
rect 3576 5507 3583 5856
rect 3596 5827 3603 6233
rect 3616 6067 3623 6293
rect 3616 5864 3623 5893
rect 3636 5607 3643 6313
rect 3656 6307 3663 6713
rect 3696 6687 3703 7073
rect 3716 6947 3723 7093
rect 3736 7087 3743 7393
rect 3756 6905 3763 7193
rect 3716 6867 3723 6893
rect 3736 6807 3743 6833
rect 3776 6667 3783 7353
rect 3836 7327 3843 7456
rect 3676 6604 3683 6653
rect 3760 6646 3780 6647
rect 3760 6643 3773 6646
rect 3756 6636 3773 6643
rect 3760 6633 3773 6636
rect 3676 6347 3683 6493
rect 3696 6384 3703 6613
rect 3796 6607 3803 7293
rect 3827 7213 3833 7227
rect 3816 7127 3823 7156
rect 3856 7067 3863 7456
rect 3876 7107 3883 7213
rect 3896 7107 3903 7676
rect 3916 7367 3923 7833
rect 3936 7347 3943 7773
rect 3976 7307 3983 7976
rect 4036 7470 4043 8033
rect 4076 7767 4083 8253
rect 4156 8127 4163 8273
rect 4176 8167 4183 8233
rect 4267 8216 4303 8223
rect 4153 7980 4167 7993
rect 4196 7987 4203 8213
rect 4296 8196 4303 8216
rect 4156 7976 4163 7980
rect 4116 7887 4123 7943
rect 4116 7827 4123 7873
rect 4116 7676 4123 7733
rect 4096 7587 4103 7643
rect 4176 7427 4183 7893
rect 3933 7227 3947 7233
rect 3936 7156 3943 7192
rect 3876 6976 3883 7033
rect 3896 7027 3903 7093
rect 3916 6767 3923 6873
rect 3816 6430 3823 6673
rect 3856 6416 3863 6453
rect 3793 6367 3807 6370
rect 3836 6363 3843 6383
rect 3816 6356 3843 6363
rect 3716 6207 3723 6333
rect 3676 5864 3683 6173
rect 3756 6116 3763 6173
rect 3796 6127 3803 6253
rect 3696 5987 3703 6073
rect 3736 6047 3743 6083
rect 3816 6047 3823 6356
rect 3896 6287 3903 6653
rect 3936 6627 3943 6913
rect 3956 6787 3963 6933
rect 3996 6887 4003 6993
rect 4016 6867 4023 7410
rect 4196 7387 4203 7456
rect 4216 7387 4223 8073
rect 4236 8047 4243 8163
rect 4236 7907 4243 8033
rect 4276 7456 4283 8113
rect 4316 8107 4323 8163
rect 4336 7947 4343 8153
rect 4356 7927 4363 8333
rect 4376 8167 4383 8195
rect 4476 8167 4483 8413
rect 4496 8127 4503 8433
rect 4536 8347 4543 8613
rect 4556 8287 4563 8533
rect 4576 8427 4583 8676
rect 4616 8447 4623 8833
rect 4656 8547 4663 8753
rect 4696 8667 4703 8713
rect 4636 8387 4643 8533
rect 4696 8496 4703 8653
rect 4736 8627 4743 8953
rect 4833 8720 4847 8733
rect 4856 8730 4863 8953
rect 4876 8767 4883 9353
rect 4896 9204 4903 9376
rect 5113 9347 5127 9353
rect 5136 9347 5143 9373
rect 4916 8827 4923 9333
rect 5080 9243 5093 9247
rect 5076 9236 5093 9243
rect 5080 9233 5093 9236
rect 5007 9203 5020 9207
rect 5007 9196 5023 9203
rect 5007 9193 5020 9196
rect 4836 8716 4843 8720
rect 4916 8707 4923 8733
rect 4936 8683 4943 9153
rect 5116 9147 5123 9236
rect 5073 9020 5087 9033
rect 5113 9027 5127 9033
rect 5136 9027 5143 9233
rect 5076 9016 5083 9020
rect 5016 8787 5023 8993
rect 5136 8987 5143 9013
rect 5056 8947 5063 8983
rect 5056 8807 5063 8933
rect 4816 8583 4823 8683
rect 4796 8576 4823 8583
rect 4916 8676 4943 8683
rect 4736 8496 4743 8573
rect 4796 8507 4803 8576
rect 4656 8447 4663 8493
rect 4667 8436 4683 8443
rect 4576 8267 4583 8293
rect 4636 8163 4643 8373
rect 4393 7980 4407 7993
rect 4396 7976 4403 7980
rect 4436 7976 4443 8093
rect 4536 8087 4543 8150
rect 4576 8107 4583 8163
rect 4616 8156 4643 8163
rect 4496 8007 4503 8033
rect 4576 7956 4583 8053
rect 4596 7967 4603 8133
rect 4416 7887 4423 7943
rect 4416 7644 4423 7673
rect 4376 7567 4383 7643
rect 4256 7307 4263 7423
rect 4296 7407 4303 7423
rect 4056 7124 4063 7193
rect 4056 6887 4063 7110
rect 4076 6887 4083 7293
rect 4116 6987 4123 7293
rect 4136 7047 4143 7156
rect 4136 6936 4143 7033
rect 4176 6936 4183 7073
rect 4216 7063 4223 7123
rect 4256 7087 4263 7113
rect 4196 7056 4223 7063
rect 4196 6987 4203 7056
rect 4216 6947 4223 7033
rect 4236 6930 4243 6953
rect 4276 6927 4283 7373
rect 4296 7187 4303 7393
rect 4296 6916 4303 6993
rect 4116 6887 4123 6903
rect 4056 6787 4063 6833
rect 3976 6647 3983 6673
rect 4056 6636 4063 6773
rect 4116 6607 4123 6873
rect 3807 6026 3820 6027
rect 3807 6013 3813 6026
rect 3656 5607 3663 5773
rect 3736 5596 3743 5973
rect 3836 5907 3843 6193
rect 3896 6167 3903 6273
rect 3936 6247 3943 6592
rect 3856 6084 3863 6153
rect 3876 6007 3883 6133
rect 3896 6087 3903 6113
rect 3896 5910 3903 6052
rect 3816 5827 3823 5863
rect 3636 5527 3643 5593
rect 3576 5427 3583 5472
rect 3556 5416 3573 5423
rect 3536 4927 3543 5132
rect 3536 4747 3543 4913
rect 3516 4147 3523 4232
rect 3496 4036 3503 4113
rect 3536 4047 3543 4553
rect 3556 4167 3563 5416
rect 3636 5376 3643 5492
rect 3576 4947 3583 5376
rect 3716 5344 3723 5373
rect 3616 5287 3623 5343
rect 3596 5087 3603 5153
rect 3636 5076 3643 5253
rect 3656 5247 3663 5330
rect 3713 5287 3727 5293
rect 3736 5247 3743 5353
rect 3673 5080 3687 5093
rect 3696 5087 3703 5193
rect 3756 5107 3763 5553
rect 3776 5287 3783 5653
rect 3796 5327 3803 5753
rect 3876 5647 3883 5673
rect 3896 5667 3903 5896
rect 3916 5767 3923 6116
rect 3936 6084 3943 6233
rect 3933 6007 3947 6013
rect 3936 5567 3943 5893
rect 3956 5767 3963 6590
rect 4036 6567 4043 6603
rect 4076 6487 4083 6603
rect 4136 6567 4143 6853
rect 4156 6707 4163 6903
rect 4096 6416 4103 6513
rect 4176 6427 4183 6873
rect 4196 6567 4203 6693
rect 4056 6287 4063 6413
rect 3976 6147 3983 6193
rect 4036 6147 4043 6173
rect 4033 6120 4047 6133
rect 4036 6116 4043 6120
rect 4016 6080 4023 6083
rect 3973 6067 3987 6073
rect 4013 6067 4027 6080
rect 4116 6047 4123 6383
rect 4056 5896 4063 6033
rect 4096 5927 4103 5953
rect 4076 5856 4103 5863
rect 3996 5643 4003 5773
rect 3996 5636 4023 5643
rect 4016 5607 4023 5636
rect 3836 5487 3843 5550
rect 3816 5447 3823 5473
rect 3816 5307 3823 5376
rect 3836 5343 3843 5452
rect 3856 5387 3863 5413
rect 3836 5336 3883 5343
rect 3676 5076 3683 5080
rect 3616 5040 3623 5043
rect 3613 5027 3627 5040
rect 3616 4856 3623 4893
rect 3656 4856 3663 5009
rect 3596 4820 3603 4823
rect 3576 4467 3583 4813
rect 3593 4807 3607 4820
rect 3636 4807 3643 4823
rect 3636 4796 3653 4807
rect 3640 4793 3653 4796
rect 3576 4387 3583 4413
rect 3396 3607 3403 4033
rect 3396 3310 3403 3572
rect 3416 3547 3423 3833
rect 3436 3647 3443 4003
rect 3476 3967 3483 4003
rect 3516 3927 3523 3990
rect 3556 3987 3563 4053
rect 3596 3987 3603 4753
rect 3636 4527 3643 4753
rect 3676 4687 3683 4813
rect 3696 4587 3703 5013
rect 3716 4767 3723 4993
rect 3736 4767 3743 5063
rect 3756 4807 3763 5053
rect 3776 4847 3783 4993
rect 3796 4927 3803 5063
rect 3796 4827 3803 4913
rect 3736 4687 3743 4753
rect 3727 4663 3740 4667
rect 3727 4653 3743 4663
rect 3656 4547 3663 4573
rect 3716 4556 3723 4613
rect 3736 4607 3743 4653
rect 3680 4303 3693 4307
rect 3636 4283 3643 4303
rect 3676 4296 3693 4303
rect 3680 4293 3693 4296
rect 3636 4276 3653 4283
rect 3627 4233 3633 4247
rect 3656 4227 3663 4273
rect 3576 3816 3583 3853
rect 3536 3767 3543 3783
rect 3527 3756 3543 3767
rect 3527 3753 3540 3756
rect 3596 3707 3603 3783
rect 3636 3747 3643 4093
rect 3656 4004 3663 4113
rect 3716 4036 3723 4333
rect 3756 4127 3763 4733
rect 3776 4287 3783 4793
rect 3796 4304 3803 4573
rect 3816 4263 3823 4953
rect 3836 4287 3843 5313
rect 3916 5207 3923 5343
rect 3996 5247 4003 5550
rect 4016 5287 4023 5373
rect 4036 5347 4043 5850
rect 4056 5467 4063 5813
rect 4073 5807 4087 5813
rect 4076 5564 4083 5653
rect 4096 5527 4103 5856
rect 4056 5227 4063 5432
rect 4076 5390 4083 5493
rect 4116 5427 4123 5973
rect 4136 5887 4143 6133
rect 4136 5507 4143 5852
rect 4156 5847 4163 6370
rect 4196 6347 4203 6513
rect 4176 6147 4183 6193
rect 4176 5927 4183 6093
rect 4196 6084 4203 6253
rect 4216 5867 4223 6873
rect 4336 6727 4343 7293
rect 4356 7123 4363 7233
rect 4436 7227 4443 7913
rect 4456 7407 4463 7930
rect 4496 7747 4503 7913
rect 4556 7587 4563 7913
rect 4616 7827 4623 8156
rect 4656 8147 4663 8196
rect 4676 8083 4683 8436
rect 4716 8427 4723 8463
rect 4880 8463 4893 8467
rect 4816 8460 4823 8463
rect 4813 8447 4827 8460
rect 4876 8456 4893 8463
rect 4880 8453 4893 8456
rect 4916 8427 4923 8676
rect 4733 8227 4747 8233
rect 4776 8167 4783 8233
rect 4796 8107 4803 8353
rect 4833 8200 4847 8213
rect 4836 8196 4843 8200
rect 4656 8080 4683 8083
rect 4653 8076 4683 8080
rect 4653 8067 4667 8076
rect 4896 7956 4903 8153
rect 4916 8147 4923 8413
rect 4936 8407 4943 8653
rect 4956 8647 4963 8733
rect 5116 8716 5123 8973
rect 5156 8727 5163 9393
rect 4956 8607 4963 8633
rect 4936 8363 4943 8393
rect 4936 8356 4963 8363
rect 4936 8167 4943 8313
rect 4956 7967 4963 8356
rect 5056 8307 5063 8683
rect 5156 8367 5163 8692
rect 5176 8463 5183 9353
rect 5256 9347 5263 9373
rect 5196 8947 5203 9253
rect 5256 9207 5263 9236
rect 5276 8927 5283 9433
rect 5296 9427 5303 9473
rect 5356 9307 5363 9473
rect 5356 9236 5363 9293
rect 5336 9127 5343 9203
rect 5376 9167 5383 9203
rect 5416 9087 5423 10493
rect 5436 10447 5443 10833
rect 5456 10627 5463 11173
rect 5496 11096 5503 11133
rect 5536 10987 5543 11063
rect 5476 10807 5483 10873
rect 5296 8967 5303 9033
rect 5336 8980 5343 8983
rect 5376 8980 5383 8983
rect 5333 8967 5347 8980
rect 5373 8967 5387 8980
rect 5196 8510 5203 8773
rect 5216 8647 5223 8713
rect 5236 8547 5243 8913
rect 5376 8907 5383 8953
rect 5436 8947 5443 10193
rect 5456 10070 5463 10613
rect 5476 10247 5483 10772
rect 5496 10544 5503 10913
rect 5516 10707 5523 10813
rect 5576 10796 5583 11173
rect 5756 11110 5763 11153
rect 5856 11063 5863 11213
rect 5816 11056 5863 11063
rect 5616 10796 5623 10853
rect 5676 10816 5683 10953
rect 5916 10927 5923 11273
rect 5936 11267 5943 11316
rect 6016 11110 6023 11616
rect 5996 11064 6003 11093
rect 5516 10207 5523 10653
rect 5536 10427 5543 10753
rect 5556 10667 5563 10763
rect 5596 10707 5603 10763
rect 5676 10667 5683 10733
rect 5596 10576 5603 10613
rect 5633 10580 5647 10593
rect 5696 10590 5703 10773
rect 5636 10576 5643 10580
rect 5556 10507 5563 10573
rect 5656 10507 5663 10543
rect 5556 10407 5563 10453
rect 5576 10276 5583 10373
rect 5596 10307 5603 10473
rect 5716 10467 5723 10783
rect 5976 10747 5983 10813
rect 5556 10207 5563 10243
rect 5596 10167 5603 10243
rect 5656 10227 5663 10276
rect 5696 10247 5703 10273
rect 5596 10056 5603 10093
rect 5256 8707 5263 8793
rect 5276 8647 5283 8892
rect 5353 8720 5367 8733
rect 5376 8727 5383 8853
rect 5416 8787 5423 8893
rect 5436 8847 5443 8912
rect 5456 8867 5463 10056
rect 5476 9567 5483 9933
rect 5496 9767 5503 10033
rect 5656 10024 5663 10073
rect 5696 10024 5703 10173
rect 5576 9967 5583 10023
rect 5496 9667 5503 9753
rect 5516 9727 5523 9813
rect 5576 9756 5583 9953
rect 5676 9847 5683 9893
rect 5716 9867 5723 10093
rect 5616 9756 5663 9763
rect 5656 9727 5663 9756
rect 5556 9567 5563 9723
rect 5596 9627 5603 9723
rect 5476 8987 5483 9013
rect 5476 8807 5483 8952
rect 5496 8747 5503 9493
rect 5516 9167 5523 9553
rect 5516 9007 5523 9053
rect 5536 8967 5543 9433
rect 5576 9267 5583 9573
rect 5636 9536 5643 9653
rect 5676 9536 5683 9653
rect 5736 9504 5743 10293
rect 5756 10207 5763 10653
rect 5776 10307 5783 10633
rect 5776 10183 5783 10272
rect 5796 10244 5803 10573
rect 5816 10447 5823 10613
rect 5916 10576 5923 10613
rect 5896 10487 5903 10543
rect 5936 10536 5953 10543
rect 5827 10223 5840 10227
rect 5827 10220 5843 10223
rect 5827 10213 5847 10220
rect 5833 10207 5847 10213
rect 5876 10207 5883 10243
rect 5756 10176 5783 10183
rect 5616 9347 5623 9503
rect 5656 9367 5663 9503
rect 5576 9236 5583 9253
rect 5600 9203 5613 9207
rect 5596 9193 5613 9203
rect 5596 9147 5603 9193
rect 5736 9127 5743 9373
rect 5756 9207 5763 10176
rect 5573 9020 5587 9033
rect 5576 9016 5583 9020
rect 5736 8984 5743 9113
rect 5596 8980 5603 8983
rect 5593 8967 5607 8980
rect 5776 8927 5783 10056
rect 5796 9387 5803 10193
rect 5936 10187 5943 10276
rect 5847 10083 5860 10087
rect 5847 10073 5863 10083
rect 5856 10056 5863 10073
rect 5956 10027 5963 10533
rect 5976 10467 5983 10673
rect 5996 10607 6003 10873
rect 6016 10827 6023 11096
rect 6036 10867 6043 11553
rect 6156 11547 6163 11583
rect 6196 11527 6203 11823
rect 6216 11567 6223 11793
rect 6276 11727 6283 11833
rect 6296 11580 6303 11583
rect 6293 11567 6307 11580
rect 6336 11547 6343 11993
rect 6376 11807 6383 11873
rect 6416 11807 6423 11973
rect 6536 11947 6543 12053
rect 6676 11987 6683 12153
rect 6753 12140 6767 12153
rect 8467 12153 8473 12167
rect 6793 12140 6807 12153
rect 6756 12136 6763 12140
rect 6796 12136 6803 12140
rect 6936 12124 6943 12153
rect 6716 12067 6723 12113
rect 6496 11836 6503 11913
rect 6476 11647 6483 11803
rect 6376 11427 6383 11633
rect 6536 11616 6543 11773
rect 6076 11276 6103 11283
rect 6076 11167 6083 11276
rect 6096 11096 6103 11133
rect 6116 11027 6123 11063
rect 6116 10827 6123 10933
rect 6156 10907 6163 10953
rect 6176 10947 6183 11413
rect 6156 10816 6163 10893
rect 6196 10847 6203 11353
rect 6256 11047 6263 11373
rect 6376 11316 6383 11413
rect 6296 11267 6303 11313
rect 6316 11027 6323 11093
rect 6336 11064 6343 11253
rect 6456 11076 6463 11213
rect 6476 11147 6483 11213
rect 6496 11167 6503 11533
rect 6516 11227 6523 11583
rect 6556 11387 6563 11570
rect 6636 11447 6643 11836
rect 6593 11320 6607 11333
rect 6596 11316 6603 11320
rect 6636 11316 6643 11433
rect 6696 11367 6703 12013
rect 6776 11907 6783 12103
rect 6816 12047 6823 12103
rect 7196 12087 7203 12116
rect 6876 12067 6883 12083
rect 6796 11836 6803 11913
rect 6716 11787 6723 11836
rect 6856 11807 6863 12033
rect 6876 12007 6883 12053
rect 6816 11767 6823 11803
rect 6673 11327 6687 11333
rect 6696 11287 6703 11353
rect 6716 11247 6723 11733
rect 6776 11616 6783 11673
rect 6816 11616 6823 11713
rect 6496 11087 6503 11153
rect 6556 11087 6563 11213
rect 6796 11187 6803 11570
rect 6896 11487 6903 11613
rect 6847 11323 6860 11327
rect 6847 11316 6863 11323
rect 6896 11316 6903 11473
rect 6936 11327 6943 11993
rect 6956 11850 6963 11973
rect 7336 11967 7343 12116
rect 7680 12103 7693 12107
rect 7296 11850 7303 11953
rect 6847 11313 6860 11316
rect 6876 11280 6883 11283
rect 6873 11267 6887 11280
rect 6556 11084 6580 11087
rect 6507 11076 6523 11083
rect 6556 11076 6573 11084
rect 6560 11073 6573 11076
rect 6376 11060 6383 11063
rect 6373 11047 6387 11060
rect 5876 10020 5883 10023
rect 5873 10007 5887 10020
rect 5876 9967 5883 9993
rect 5836 9756 5843 9813
rect 5876 9756 5883 9953
rect 5916 9587 5923 9933
rect 5976 9907 5983 10273
rect 5996 9507 6003 10572
rect 6016 10247 6023 10773
rect 6036 10747 6043 10783
rect 6036 10527 6043 10693
rect 6036 10007 6043 10513
rect 6096 10507 6103 10783
rect 6076 10327 6083 10453
rect 6116 10343 6123 10773
rect 6176 10707 6183 10773
rect 6196 10687 6203 10783
rect 6476 10784 6483 11033
rect 6466 10776 6467 10780
rect 6453 10763 6467 10776
rect 6453 10760 6483 10763
rect 6456 10756 6483 10760
rect 6476 10727 6483 10756
rect 6516 10747 6523 10770
rect 6516 10667 6523 10733
rect 6136 10587 6143 10613
rect 6173 10580 6187 10593
rect 6176 10576 6183 10580
rect 6316 10556 6323 10653
rect 6636 10556 6643 10913
rect 6876 10907 6883 11030
rect 6916 10987 6923 11073
rect 6936 11044 6943 11313
rect 6956 11267 6963 11836
rect 7256 11767 7263 11813
rect 7316 11800 7323 11803
rect 7313 11787 7327 11800
rect 7016 11547 7023 11673
rect 7056 11627 7063 11753
rect 7047 11616 7063 11627
rect 7096 11616 7103 11693
rect 7047 11613 7060 11616
rect 7156 11584 7163 11733
rect 7296 11627 7303 11653
rect 7336 11616 7343 11753
rect 7076 11547 7083 11583
rect 6976 11284 6983 11513
rect 7356 11507 7363 11583
rect 7396 11487 7403 11583
rect 7476 11547 7483 11593
rect 6656 10784 6663 10833
rect 6156 10507 6163 10543
rect 6196 10540 6203 10543
rect 6193 10527 6207 10540
rect 6096 10336 6123 10343
rect 6096 10107 6103 10336
rect 6156 10290 6163 10333
rect 6196 10276 6203 10492
rect 6296 10407 6303 10433
rect 6356 10427 6363 10550
rect 6676 10427 6683 10523
rect 6656 10416 6673 10423
rect 6656 10296 6663 10416
rect 6716 10383 6723 10653
rect 6736 10427 6743 10893
rect 6696 10376 6723 10383
rect 6696 10287 6703 10376
rect 6776 10327 6783 10793
rect 6816 10687 6823 10763
rect 6856 10647 6863 10763
rect 6796 10347 6803 10533
rect 6816 10507 6823 10633
rect 6936 10627 6943 10893
rect 6956 10576 6963 11053
rect 6976 10847 6983 11093
rect 6707 10276 6723 10283
rect 6096 10083 6103 10093
rect 6096 10076 6123 10083
rect 6116 10056 6123 10076
rect 6156 10056 6163 10173
rect 6176 10087 6183 10243
rect 6236 10187 6243 10263
rect 5936 9447 5943 9503
rect 5876 9236 5883 9273
rect 5816 8947 5823 9203
rect 5916 9107 5923 9236
rect 5356 8716 5363 8720
rect 5213 8500 5227 8513
rect 5216 8496 5223 8500
rect 5176 8456 5203 8463
rect 5236 8460 5243 8463
rect 4996 8047 5003 8196
rect 5036 8167 5043 8196
rect 5056 7956 5063 8253
rect 5096 8247 5103 8273
rect 5136 8196 5143 8333
rect 5116 8160 5123 8163
rect 5113 8147 5127 8160
rect 4616 7676 4623 7792
rect 4596 7607 4603 7643
rect 4536 7456 4543 7495
rect 4576 7456 4623 7463
rect 4556 7420 4563 7423
rect 4553 7407 4567 7420
rect 4616 7247 4623 7456
rect 4396 7167 4403 7213
rect 4616 6916 4623 7193
rect 4636 7127 4643 7593
rect 4636 6924 4643 7053
rect 4656 6947 4663 7573
rect 4696 7467 4703 7573
rect 4676 6927 4683 7393
rect 4696 6907 4703 6953
rect 4656 6867 4663 6883
rect 4320 6663 4333 6667
rect 4316 6653 4333 6663
rect 4316 6636 4323 6653
rect 4236 6227 4243 6636
rect 4256 6347 4263 6473
rect 4276 6187 4283 6553
rect 4296 6387 4303 6590
rect 4336 6567 4343 6603
rect 4356 6416 4363 6453
rect 4396 6430 4403 6673
rect 4280 6123 4293 6127
rect 4276 6116 4293 6123
rect 4280 6113 4293 6116
rect 4316 6107 4323 6413
rect 4456 6367 4463 6713
rect 4336 6087 4343 6133
rect 4356 5987 4363 6113
rect 4376 5987 4383 6333
rect 4396 6087 4403 6353
rect 4256 5827 4263 5973
rect 4416 5927 4423 6273
rect 4273 5907 4287 5913
rect 4313 5900 4327 5913
rect 4316 5896 4323 5900
rect 4296 5847 4303 5863
rect 4136 5447 4143 5493
rect 4176 5407 4183 5693
rect 4216 5687 4223 5753
rect 4216 5596 4223 5673
rect 4256 5647 4263 5693
rect 4253 5607 4267 5612
rect 4276 5567 4283 5793
rect 4296 5667 4303 5833
rect 4296 5627 4303 5653
rect 4236 5507 4243 5563
rect 4236 5427 4243 5493
rect 4216 5340 4223 5343
rect 4213 5327 4227 5340
rect 4096 5207 4103 5233
rect 4136 5127 4143 5233
rect 4156 5096 4163 5213
rect 3856 5027 3863 5093
rect 4116 5043 4123 5063
rect 4116 5036 4143 5043
rect 3936 4887 3943 4933
rect 3933 4860 3947 4873
rect 3936 4856 3943 4860
rect 3876 4787 3883 4823
rect 3853 4767 3867 4773
rect 3916 4767 3923 4823
rect 3976 4787 3983 4853
rect 3816 4256 3843 4263
rect 3776 4127 3783 4233
rect 3796 4047 3803 4153
rect 3676 3967 3683 4036
rect 3607 3696 3623 3703
rect 3556 3667 3563 3693
rect 3436 3303 3443 3593
rect 3573 3520 3587 3533
rect 3576 3516 3583 3520
rect 3416 3296 3443 3303
rect 3496 3296 3503 3433
rect 3516 3407 3523 3483
rect 3536 3367 3543 3413
rect 3376 2996 3383 3053
rect 3076 2856 3103 2863
rect 3076 2827 3083 2856
rect 3356 2770 3363 2953
rect 3416 2887 3423 3296
rect 3436 2947 3443 3153
rect 3456 3067 3463 3263
rect 3436 2787 3443 2853
rect 2896 2707 2903 2743
rect 2856 2287 2863 2553
rect 2876 2287 2883 2533
rect 2896 2347 2903 2473
rect 2896 2256 2903 2293
rect 2916 2287 2923 2713
rect 2996 2487 3003 2653
rect 3036 2496 3043 2613
rect 3076 2547 3083 2733
rect 3396 2663 3403 2723
rect 3396 2656 3413 2663
rect 3436 2627 3443 2752
rect 3456 2687 3463 2773
rect 3476 2667 3483 3033
rect 3516 2996 3523 3113
rect 3556 3007 3563 3483
rect 2956 2407 2963 2430
rect 2936 2256 2943 2333
rect 2976 2227 2983 2273
rect 2876 2087 2883 2223
rect 2916 2103 2923 2210
rect 2896 2096 2923 2103
rect 2896 1983 2903 2096
rect 2876 1976 2903 1983
rect 2596 1187 2603 1493
rect 2616 1404 2623 1733
rect 2656 1667 2663 1703
rect 2696 1627 2703 1703
rect 2736 1647 2743 1953
rect 2736 1436 2743 1473
rect 2616 1187 2623 1253
rect 2536 876 2563 883
rect 2556 827 2563 876
rect 2576 847 2583 993
rect 2636 787 2643 1433
rect 2696 1216 2703 1253
rect 2667 1183 2680 1187
rect 2667 1176 2683 1183
rect 2667 1173 2680 1176
rect 2716 1147 2723 1183
rect 2776 1007 2783 1953
rect 2796 1927 2803 1955
rect 2876 1956 2883 1976
rect 2916 1927 2923 2073
rect 2956 1987 2963 2013
rect 2796 987 2803 1913
rect 2936 1847 2943 1973
rect 2996 1867 3003 2353
rect 3076 2187 3083 2463
rect 3356 2447 3363 2513
rect 3396 2460 3403 2463
rect 3393 2447 3407 2460
rect 3236 2067 3243 2256
rect 3176 1956 3183 1993
rect 3196 1970 3203 2013
rect 2836 1184 2843 1473
rect 2856 1027 2863 1833
rect 2956 1736 2963 1813
rect 2876 1527 2883 1573
rect 2896 1567 2903 1703
rect 2876 1404 2883 1513
rect 2936 1507 2943 1703
rect 3116 1704 3123 1923
rect 3236 1907 3243 2053
rect 2976 1450 2983 1593
rect 3016 1436 3023 1693
rect 3036 1447 3043 1513
rect 3156 1507 3163 1633
rect 2996 1327 3003 1403
rect 3076 1287 3083 1410
rect 3136 1347 3143 1423
rect 3156 1327 3163 1416
rect 2936 1147 2943 1213
rect 2716 867 2723 933
rect 2773 920 2787 933
rect 2776 916 2783 920
rect 2756 807 2763 883
rect 2536 627 2543 696
rect 2576 567 2583 663
rect 2576 507 2583 553
rect 2656 547 2663 663
rect 2696 627 2703 696
rect 2776 664 2783 733
rect 2796 427 2803 883
rect 2856 703 2863 973
rect 2976 930 2983 1170
rect 3056 1167 3063 1213
rect 3076 1184 3083 1273
rect 2876 887 2883 916
rect 2976 807 2983 916
rect 2836 696 2863 703
rect 2896 696 2903 753
rect 2836 427 2843 696
rect 2696 390 2703 413
rect 2356 360 2363 363
rect 2276 307 2283 353
rect 2353 347 2367 360
rect 2356 267 2363 333
rect 2436 287 2443 383
rect 2756 380 2763 383
rect 2816 380 2823 383
rect 2753 367 2767 380
rect 2813 367 2827 380
rect 2756 327 2763 353
rect 2116 107 2123 143
rect 2496 43 2503 273
rect 2596 156 2603 253
rect 2756 170 2763 313
rect 2776 147 2783 233
rect 2856 176 2863 653
rect 2956 623 2963 653
rect 2976 627 2983 693
rect 2927 616 2963 623
rect 2976 190 2983 413
rect 2996 364 3003 1013
rect 3036 916 3043 1013
rect 3116 927 3123 1216
rect 3116 747 3123 773
rect 3116 664 3123 733
rect 3136 627 3143 993
rect 3176 887 3183 1893
rect 3296 1703 3303 2133
rect 3316 1827 3323 2113
rect 3216 1667 3223 1703
rect 3256 1696 3303 1703
rect 3336 1527 3343 2273
rect 3456 2256 3463 2413
rect 3496 2347 3503 2933
rect 3516 2287 3523 2913
rect 3436 2187 3443 2223
rect 3473 2007 3487 2013
rect 3413 1960 3427 1973
rect 3416 1956 3423 1960
rect 3496 1924 3503 2113
rect 3513 2047 3527 2053
rect 3536 2007 3543 2873
rect 3556 2687 3563 2993
rect 3556 2464 3563 2513
rect 3556 2227 3563 2256
rect 3396 1704 3403 1923
rect 3496 1736 3503 1773
rect 3536 1767 3543 1972
rect 3556 1943 3563 2173
rect 3576 1970 3583 2913
rect 3596 2067 3603 3133
rect 3616 2787 3623 3696
rect 3656 3547 3663 3713
rect 3636 3487 3643 3516
rect 3636 3127 3643 3193
rect 3656 2827 3663 3173
rect 3676 2967 3683 3133
rect 3696 2887 3703 3953
rect 3716 3347 3723 3973
rect 3736 3507 3743 3990
rect 3776 3947 3783 4003
rect 3836 3816 3843 4256
rect 3856 3867 3863 4732
rect 3996 4647 4003 4873
rect 4016 4787 4023 4853
rect 3876 4387 3883 4613
rect 3956 4587 3963 4613
rect 3956 4556 3963 4573
rect 3993 4560 4007 4573
rect 4036 4567 4043 4953
rect 3996 4556 4003 4560
rect 3896 4524 3903 4553
rect 3916 4336 3923 4453
rect 3976 4447 3983 4523
rect 4016 4403 4023 4523
rect 3996 4400 4023 4403
rect 3993 4396 4023 4400
rect 3993 4387 4007 4396
rect 4006 4380 4007 4387
rect 3887 4304 3900 4307
rect 3887 4297 3903 4304
rect 3887 4293 3900 4297
rect 3876 3967 3883 4272
rect 3896 4147 3903 4233
rect 3896 3887 3903 3913
rect 3896 3823 3903 3873
rect 3876 3816 3903 3823
rect 3756 3310 3763 3770
rect 3896 3587 3903 3613
rect 3796 3516 3803 3553
rect 3896 3427 3903 3516
rect 3916 3484 3923 4053
rect 3936 3647 3943 4293
rect 3956 3987 3963 4093
rect 3996 4067 4003 4373
rect 4016 4307 4023 4373
rect 4016 4036 4023 4213
rect 3736 3207 3743 3263
rect 3836 3207 3843 3373
rect 3936 3367 3943 3633
rect 3956 3527 3963 3553
rect 3736 2996 3743 3053
rect 3836 2963 3843 3193
rect 3736 2747 3743 2873
rect 3696 2740 3703 2743
rect 3693 2727 3707 2740
rect 3636 2567 3643 2673
rect 3776 2647 3783 2813
rect 3636 2327 3643 2553
rect 3753 2480 3767 2493
rect 3796 2490 3803 2963
rect 3816 2956 3843 2963
rect 3816 2567 3823 2956
rect 3836 2507 3843 2893
rect 3756 2476 3763 2480
rect 3696 2267 3703 2443
rect 3736 2440 3743 2443
rect 3733 2427 3747 2440
rect 3733 2260 3747 2273
rect 3736 2256 3743 2260
rect 3593 1987 3607 1993
rect 3556 1936 3583 1943
rect 3533 1740 3547 1753
rect 3536 1736 3543 1740
rect 3396 1567 3403 1690
rect 3516 1607 3523 1703
rect 3516 1547 3523 1593
rect 3196 1387 3203 1456
rect 3536 1427 3543 1513
rect 3576 1387 3583 1936
rect 3256 1216 3263 1313
rect 3336 1184 3343 1253
rect 3236 1180 3243 1183
rect 3233 1167 3247 1180
rect 3256 884 3263 953
rect 3316 916 3323 1113
rect 3356 916 3363 953
rect 3216 696 3223 753
rect 3276 663 3283 873
rect 3336 847 3343 883
rect 3456 696 3463 1373
rect 3476 1176 3503 1183
rect 3476 1147 3483 1176
rect 3616 967 3623 2253
rect 3776 2127 3783 2413
rect 3796 2167 3803 2253
rect 3836 2107 3843 2193
rect 3647 2033 3653 2047
rect 3660 2026 3680 2027
rect 3667 2023 3680 2026
rect 3667 2013 3683 2023
rect 3676 1956 3683 2013
rect 3740 1963 3753 1967
rect 3736 1956 3753 1963
rect 3740 1953 3753 1956
rect 3716 1920 3723 1923
rect 3713 1907 3727 1920
rect 3756 1763 3763 1893
rect 3776 1787 3783 2053
rect 3796 1867 3803 1953
rect 3756 1756 3783 1763
rect 3656 1707 3663 1753
rect 3776 1736 3783 1756
rect 3696 1587 3703 1736
rect 3756 1587 3763 1703
rect 3836 1627 3843 1813
rect 3676 1327 3683 1493
rect 3696 1404 3703 1573
rect 3756 1436 3763 1493
rect 3636 916 3643 1153
rect 3676 930 3683 1313
rect 3776 987 3783 1403
rect 3856 1223 3863 3093
rect 3876 2964 3883 3293
rect 3896 3047 3903 3353
rect 3976 3327 3983 3993
rect 3996 3387 4003 4003
rect 4036 3947 4043 4003
rect 4076 3927 4083 4933
rect 4096 3847 4103 4893
rect 4136 4867 4143 5036
rect 4176 4947 4183 5053
rect 4196 5007 4203 5113
rect 4216 4967 4223 5113
rect 4236 4907 4243 5333
rect 4220 4823 4233 4827
rect 4156 4820 4163 4823
rect 4116 4527 4123 4573
rect 4136 4507 4143 4813
rect 4153 4807 4167 4820
rect 4216 4816 4233 4823
rect 4220 4813 4233 4816
rect 4256 4807 4263 5513
rect 4276 5387 4283 5532
rect 4296 5527 4303 5592
rect 4276 5067 4283 5313
rect 4316 5307 4323 5813
rect 4336 5547 4343 5863
rect 4396 5647 4403 5913
rect 4316 5127 4323 5293
rect 4296 5047 4303 5073
rect 4316 5023 4323 5092
rect 4296 5016 4323 5023
rect 4136 4350 4143 4472
rect 4156 4447 4163 4556
rect 4156 4300 4163 4303
rect 4153 4287 4167 4300
rect 4156 4187 4163 4273
rect 4116 4007 4123 4073
rect 4016 3784 4023 3833
rect 4176 3827 4183 4033
rect 4056 3667 4063 3816
rect 4096 3747 4103 3783
rect 4147 3783 4160 3787
rect 4147 3776 4163 3783
rect 4147 3773 4160 3776
rect 4016 3587 4023 3653
rect 3916 3227 3923 3293
rect 3916 3027 3923 3213
rect 3936 2907 3943 3313
rect 3996 3296 4003 3373
rect 4036 3310 4043 3493
rect 4116 3447 4123 3483
rect 3956 2927 3963 3153
rect 3976 2947 3983 3250
rect 4016 3067 4023 3263
rect 4056 3207 4063 3250
rect 4096 3107 4103 3293
rect 4116 3087 4123 3433
rect 4013 3000 4027 3013
rect 4016 2996 4023 3000
rect 4100 3003 4113 3007
rect 4096 2996 4113 3003
rect 4100 2993 4113 2996
rect 3987 2936 4003 2943
rect 3836 1216 3863 1223
rect 3816 1180 3823 1183
rect 3813 1167 3827 1180
rect 3876 1147 3883 2733
rect 3896 2167 3903 2713
rect 3916 2490 3923 2743
rect 3976 2667 3983 2833
rect 3996 2527 4003 2936
rect 4036 2847 4043 2963
rect 4073 2947 4087 2950
rect 4136 2947 4143 3413
rect 4016 2547 4023 2776
rect 4076 2683 4083 2873
rect 4096 2707 4103 2933
rect 4156 2923 4163 3753
rect 4176 3267 4183 3773
rect 4196 3767 4203 4793
rect 4233 4787 4247 4792
rect 4236 4556 4243 4673
rect 4276 4667 4283 4953
rect 4296 4767 4303 5016
rect 4316 4747 4323 4993
rect 4216 4287 4223 4513
rect 4236 4087 4243 4473
rect 4256 4307 4263 4523
rect 4296 4520 4303 4523
rect 4293 4507 4307 4520
rect 4196 3487 4203 3693
rect 4216 3627 4223 4073
rect 4276 4036 4283 4273
rect 4316 4167 4323 4193
rect 4236 3487 4243 3573
rect 4216 3476 4233 3483
rect 4136 2916 4163 2923
rect 4116 2787 4123 2833
rect 4116 2727 4123 2773
rect 4076 2676 4103 2683
rect 3916 1723 3923 2333
rect 3936 2287 3943 2513
rect 4036 2476 4043 2593
rect 3976 2367 3983 2443
rect 4033 2270 4047 2273
rect 4056 2224 4063 2333
rect 3976 2220 3983 2223
rect 3973 2207 3987 2220
rect 4076 2207 4083 2553
rect 4096 2267 4103 2676
rect 3973 1960 3987 1973
rect 3976 1956 3983 1960
rect 4036 1956 4083 1963
rect 4076 1927 4083 1956
rect 4016 1920 4023 1923
rect 4013 1907 4027 1920
rect 3916 1716 3943 1723
rect 3896 1407 3903 1690
rect 3936 1427 3943 1716
rect 3236 627 3243 663
rect 3256 656 3283 663
rect 3136 347 3143 613
rect 3256 367 3263 656
rect 3336 396 3343 613
rect 3376 176 3383 653
rect 3476 627 3483 663
rect 3416 364 3423 393
rect 3476 227 3483 613
rect 3576 396 3583 693
rect 3616 664 3623 883
rect 3676 707 3683 916
rect 3716 787 3723 913
rect 3616 396 3623 593
rect 3636 407 3643 696
rect 3736 696 3743 733
rect 3796 687 3803 1053
rect 3816 707 3823 1132
rect 3856 916 3863 1013
rect 3876 847 3883 883
rect 3956 867 3963 1773
rect 3996 1704 4003 1773
rect 4056 1736 4063 1893
rect 4096 1787 4103 2253
rect 4116 2207 4123 2233
rect 4076 1683 4083 1703
rect 4076 1676 4103 1683
rect 4096 1587 4103 1676
rect 4016 1367 4023 1403
rect 4036 1216 4043 1273
rect 4096 1067 4103 1573
rect 4116 1287 4123 1533
rect 4136 1407 4143 2916
rect 4176 2907 4183 2993
rect 4176 2776 4183 2813
rect 4196 2807 4203 3333
rect 4216 2947 4223 3476
rect 4236 2887 4243 3452
rect 4256 3267 4263 4003
rect 4296 3967 4303 4003
rect 4276 3467 4283 3913
rect 4296 3387 4303 3873
rect 4316 3707 4323 3813
rect 4336 3787 4343 5473
rect 4356 5207 4363 5633
rect 4376 5207 4383 5413
rect 4396 5367 4403 5612
rect 4396 5076 4403 5273
rect 4416 5107 4423 5913
rect 4436 5907 4443 6173
rect 4436 5407 4443 5872
rect 4456 5767 4463 6253
rect 4476 6147 4483 6813
rect 4533 6643 4547 6653
rect 4533 6640 4563 6643
rect 4536 6636 4563 6640
rect 4596 6636 4603 6793
rect 4656 6727 4663 6853
rect 4496 6327 4503 6636
rect 4576 6600 4583 6603
rect 4573 6587 4587 6600
rect 4616 6567 4623 6603
rect 4516 6347 4523 6453
rect 4496 6116 4503 6173
rect 4536 6116 4543 6473
rect 4616 6427 4623 6553
rect 4656 6416 4663 6573
rect 4676 6467 4683 6873
rect 4576 6087 4583 6413
rect 4596 6384 4603 6413
rect 4716 6407 4723 7813
rect 4756 7787 4763 7853
rect 4736 7424 4743 7453
rect 4756 7387 4763 7752
rect 4776 7667 4783 7793
rect 4796 7470 4803 7833
rect 4827 7773 4833 7787
rect 4816 7647 4823 7733
rect 4856 7676 4863 7773
rect 4916 7676 4923 7753
rect 4936 7707 4943 7910
rect 4976 7747 4983 7913
rect 5096 7887 5103 8133
rect 5156 8067 5163 8163
rect 5196 8087 5203 8456
rect 5233 8447 5247 8460
rect 5276 8427 5283 8463
rect 5236 8107 5243 8313
rect 5296 8267 5303 8353
rect 5316 8067 5323 8293
rect 5356 8196 5363 8353
rect 5396 8207 5403 8693
rect 5416 8647 5423 8703
rect 5416 8196 5423 8293
rect 5436 8247 5443 8613
rect 5476 8547 5483 8703
rect 5516 8667 5523 8753
rect 5816 8747 5823 8813
rect 5833 8740 5847 8753
rect 5836 8736 5843 8740
rect 5536 8687 5543 8733
rect 5796 8607 5803 8703
rect 5476 8496 5523 8503
rect 5476 8387 5483 8496
rect 5536 8460 5543 8463
rect 5456 8227 5463 8353
rect 5496 8307 5503 8453
rect 5533 8447 5547 8460
rect 5576 8427 5583 8463
rect 5493 8200 5507 8213
rect 5496 8196 5503 8200
rect 5556 8196 5563 8293
rect 5576 8267 5583 8313
rect 5576 8227 5583 8253
rect 5376 8127 5383 8163
rect 5436 8147 5443 8163
rect 5376 7956 5383 8092
rect 5436 8027 5443 8133
rect 5416 7920 5423 7923
rect 5413 7907 5427 7920
rect 5453 7907 5467 7913
rect 5036 7747 5043 7793
rect 4887 7636 4903 7643
rect 4776 7156 4783 7233
rect 4816 7187 4823 7423
rect 4856 7287 4863 7433
rect 4896 7424 4903 7636
rect 4820 7163 4833 7167
rect 4816 7156 4833 7163
rect 4820 7153 4833 7156
rect 4876 7147 4883 7353
rect 4896 7267 4903 7410
rect 4736 6727 4743 7113
rect 4756 7007 4763 7123
rect 4796 7067 4803 7123
rect 4756 6847 4763 6993
rect 4756 6387 4763 6773
rect 4776 6387 4783 6933
rect 4796 6807 4803 6973
rect 4836 6867 4843 7093
rect 4856 6947 4863 7013
rect 4896 6936 4903 7153
rect 4916 7087 4923 7113
rect 4936 7107 4943 7613
rect 4956 7567 4963 7663
rect 5056 7664 5063 7753
rect 5376 7710 5383 7893
rect 5396 7707 5403 7733
rect 4956 6927 4963 7353
rect 4976 7107 4983 7653
rect 5076 7627 5083 7696
rect 5416 7667 5423 7753
rect 4996 7047 5003 7173
rect 4976 7007 4983 7033
rect 4976 6916 4983 6993
rect 5016 6987 5023 7533
rect 5056 7527 5063 7573
rect 5073 7460 5087 7473
rect 5076 7456 5083 7460
rect 5356 7456 5363 7573
rect 5056 7207 5063 7423
rect 5076 7156 5083 7213
rect 5136 7187 5143 7213
rect 5136 7156 5143 7173
rect 5047 7123 5060 7127
rect 5047 7116 5063 7123
rect 5047 7113 5060 7116
rect 5033 7083 5047 7092
rect 5033 7080 5063 7083
rect 5036 7076 5063 7080
rect 5056 6923 5063 7076
rect 5036 6916 5063 6923
rect 4836 6636 4843 6753
rect 4876 6687 4883 6890
rect 4916 6847 4923 6903
rect 4916 6603 4923 6733
rect 4676 6347 4683 6370
rect 4696 6307 4703 6373
rect 4476 5610 4483 6073
rect 4576 5967 4583 6073
rect 4573 5900 4587 5913
rect 4613 5900 4627 5913
rect 4576 5896 4583 5900
rect 4616 5896 4623 5900
rect 4536 5603 4543 5893
rect 4536 5596 4563 5603
rect 4527 5556 4543 5563
rect 4473 5427 4487 5433
rect 4473 5380 4487 5392
rect 4496 5387 4503 5453
rect 4536 5427 4543 5556
rect 4476 5376 4483 5380
rect 4516 5307 4523 5353
rect 4536 5107 4543 5413
rect 4556 5127 4563 5596
rect 4576 5107 4583 5833
rect 4596 5807 4603 5863
rect 4356 4687 4363 4813
rect 4376 4707 4383 5043
rect 4396 4827 4403 4873
rect 4456 4856 4463 5033
rect 4476 4967 4483 5053
rect 4496 5007 4503 5063
rect 4496 4856 4503 4933
rect 4516 4867 4523 5013
rect 4427 4823 4440 4827
rect 4427 4816 4443 4823
rect 4427 4813 4440 4816
rect 4420 4806 4433 4807
rect 4427 4793 4433 4806
rect 4356 4387 4363 4652
rect 4376 4467 4383 4693
rect 4396 4487 4403 4653
rect 4436 4570 4443 4613
rect 4376 4336 4383 4432
rect 4416 4350 4423 4493
rect 4436 4387 4443 4556
rect 4356 3967 4363 4293
rect 4376 3927 4383 4273
rect 4456 3967 4463 4773
rect 4416 3816 4423 3893
rect 4376 3516 4383 3653
rect 4476 3607 4483 4823
rect 4536 4787 4543 5053
rect 4556 4927 4563 5063
rect 4556 4807 4563 4913
rect 4576 4807 4583 4933
rect 4553 4560 4567 4573
rect 4556 4556 4563 4560
rect 4496 4247 4503 4453
rect 4536 4447 4543 4523
rect 4536 4036 4543 4373
rect 4556 4107 4563 4473
rect 4576 4247 4583 4513
rect 4596 4487 4603 5753
rect 4613 5427 4627 5433
rect 4636 5307 4643 5633
rect 4656 5567 4663 6033
rect 4676 5727 4683 6116
rect 4696 5967 4703 6293
rect 4696 5707 4703 5853
rect 4716 5847 4723 6372
rect 4736 6187 4743 6293
rect 4736 5647 4743 6133
rect 4856 6123 4863 6603
rect 4896 6596 4923 6603
rect 4896 6416 4903 6596
rect 4936 6527 4943 6893
rect 4956 6767 4963 6833
rect 5076 6807 5083 7093
rect 5116 7087 5123 7123
rect 5176 7107 5183 7313
rect 5256 7087 5263 7253
rect 5296 7247 5303 7423
rect 5336 7367 5343 7423
rect 5396 7227 5403 7453
rect 5296 7107 5303 7193
rect 5356 7156 5363 7193
rect 5416 7167 5423 7473
rect 5336 7067 5343 7123
rect 5096 6887 5103 6933
rect 5356 6916 5363 7093
rect 5416 7043 5423 7113
rect 5436 7087 5443 7853
rect 5416 7036 5443 7043
rect 5376 7020 5423 7023
rect 5373 7016 5423 7020
rect 5373 7007 5387 7016
rect 5386 7000 5387 7007
rect 5396 6947 5403 6993
rect 5416 6987 5423 7016
rect 5396 6880 5403 6883
rect 5393 6867 5407 6880
rect 5096 6650 5103 6733
rect 4956 6567 4963 6636
rect 4936 6447 4943 6513
rect 4956 6487 4963 6553
rect 4933 6420 4947 6433
rect 4936 6416 4943 6420
rect 4836 6116 4863 6123
rect 4756 5807 4763 6073
rect 4776 5847 4783 5993
rect 4816 5983 4823 6083
rect 4856 5987 4863 6070
rect 4876 6047 4883 6373
rect 4896 6047 4903 6093
rect 4796 5976 4823 5983
rect 4796 5627 4803 5976
rect 4816 5723 4823 5953
rect 4896 5896 4903 6033
rect 4916 6007 4923 6383
rect 4936 6067 4943 6133
rect 4956 6087 4963 6383
rect 4876 5847 4883 5863
rect 4876 5836 4893 5847
rect 4880 5833 4893 5836
rect 4816 5716 4843 5723
rect 4773 5600 4787 5613
rect 4776 5596 4783 5600
rect 4696 5507 4703 5596
rect 4836 5567 4843 5716
rect 4856 5567 4863 5833
rect 4916 5803 4923 5853
rect 4936 5843 4943 5973
rect 4956 5887 4963 6033
rect 4976 5867 4983 6373
rect 4996 6003 5003 6513
rect 5016 6147 5023 6433
rect 5056 6267 5063 6636
rect 5036 6207 5043 6233
rect 5116 6227 5123 6603
rect 5256 6487 5263 6793
rect 5256 6383 5263 6473
rect 5016 6027 5023 6112
rect 5136 6087 5143 6153
rect 5056 6080 5063 6083
rect 4996 5996 5023 6003
rect 4936 5836 4963 5843
rect 4896 5796 4923 5803
rect 4656 5347 4663 5453
rect 4696 5307 4703 5343
rect 4796 5267 4803 5550
rect 4836 5247 4843 5343
rect 4876 5327 4883 5793
rect 4896 5107 4903 5796
rect 4916 5227 4923 5573
rect 4936 5527 4943 5753
rect 4916 5127 4923 5213
rect 4916 5096 4923 5113
rect 4616 5070 4623 5093
rect 4956 5067 4963 5836
rect 5016 5687 5023 5996
rect 5036 5667 5043 6073
rect 5053 6067 5067 6080
rect 5096 6067 5103 6083
rect 5176 6067 5183 6383
rect 5216 6267 5223 6383
rect 5236 6376 5263 6383
rect 5216 6207 5223 6232
rect 5096 5947 5103 6053
rect 5116 5896 5123 5933
rect 5156 5896 5163 6013
rect 5076 5867 5083 5896
rect 5136 5860 5143 5863
rect 5096 5767 5103 5853
rect 5133 5847 5147 5860
rect 5176 5787 5183 5863
rect 5076 5707 5083 5753
rect 5033 5600 5047 5613
rect 5036 5596 5043 5600
rect 4616 5027 4623 5056
rect 4856 5023 4863 5053
rect 4876 5043 4883 5063
rect 4876 5036 4903 5043
rect 4856 5016 4883 5023
rect 4696 4856 4703 4913
rect 4733 4860 4747 4873
rect 4736 4856 4743 4860
rect 4616 4667 4623 4853
rect 4616 4427 4623 4613
rect 4656 4336 4663 4573
rect 4696 4527 4703 4793
rect 4716 4707 4723 4823
rect 4756 4803 4763 4823
rect 4736 4796 4763 4803
rect 4736 4767 4743 4796
rect 4627 4303 4640 4307
rect 4627 4296 4643 4303
rect 4627 4293 4640 4296
rect 4576 4207 4583 4233
rect 4576 4004 4583 4153
rect 4496 3807 4503 3853
rect 4416 3516 4423 3553
rect 4316 3367 4323 3473
rect 4356 3427 4363 3483
rect 4396 3447 4403 3470
rect 4416 3427 4423 3453
rect 4356 3296 4363 3373
rect 4253 2790 4267 2793
rect 4156 2427 4163 2713
rect 4236 2707 4243 2743
rect 4256 2707 4263 2730
rect 4156 1247 4163 2153
rect 4176 1970 4183 2553
rect 4196 2267 4203 2673
rect 4236 2476 4243 2633
rect 4276 2547 4283 3253
rect 4296 3227 4303 3263
rect 4316 2996 4323 3053
rect 4376 2996 4383 3213
rect 4396 3067 4403 3250
rect 4296 2567 4303 2813
rect 4316 2476 4323 2893
rect 4356 2807 4363 2873
rect 4416 2823 4423 3333
rect 4396 2816 4423 2823
rect 4336 2744 4343 2793
rect 4336 2687 4343 2730
rect 4256 2440 4263 2443
rect 4253 2427 4267 2440
rect 4296 2407 4303 2443
rect 4216 2167 4223 2223
rect 4256 2207 4263 2223
rect 4296 2207 4303 2313
rect 4256 2027 4263 2193
rect 4356 2147 4363 2772
rect 4216 1507 4223 2013
rect 4296 1956 4303 2013
rect 4256 1547 4263 1833
rect 4316 1787 4323 1923
rect 4356 1750 4363 2133
rect 4116 1187 4123 1217
rect 4216 1007 4223 1493
rect 4256 1436 4263 1473
rect 4296 1436 4303 1493
rect 4276 1230 4283 1253
rect 4296 1127 4303 1183
rect 3876 767 3883 833
rect 3816 664 3823 693
rect 4056 663 4063 993
rect 4096 667 4103 933
rect 4173 920 4187 933
rect 4213 920 4227 933
rect 4176 916 4183 920
rect 4216 916 4223 920
rect 4156 807 4163 883
rect 4256 703 4263 973
rect 4276 887 4283 933
rect 4296 827 4303 916
rect 4236 696 4263 703
rect 4316 697 4323 733
rect 4376 731 4383 2813
rect 4396 2163 4403 2816
rect 4416 2607 4423 2793
rect 4436 2787 4443 3473
rect 4476 3447 4483 3493
rect 4496 3227 4503 3693
rect 4456 2827 4463 3173
rect 4496 3167 4503 3213
rect 4516 3107 4523 3953
rect 4536 3547 4543 3913
rect 4556 3727 4563 3953
rect 4596 3784 4603 4253
rect 4616 3823 4623 4233
rect 4636 4067 4643 4233
rect 4676 3907 4683 4193
rect 4696 3883 4703 4133
rect 4716 4107 4723 4213
rect 4736 4063 4743 4753
rect 4776 4727 4783 4793
rect 4787 4583 4800 4587
rect 4787 4573 4803 4583
rect 4796 4556 4803 4573
rect 4776 4407 4783 4523
rect 4776 4367 4783 4393
rect 4796 4287 4803 4433
rect 4816 4327 4823 4493
rect 4716 4056 4743 4063
rect 4716 4007 4723 4056
rect 4716 3967 4723 3993
rect 4736 3967 4743 4033
rect 4796 4000 4803 4003
rect 4793 3987 4807 4000
rect 4676 3876 4703 3883
rect 4616 3816 4643 3823
rect 4676 3816 4683 3876
rect 4713 3847 4727 3853
rect 4736 3827 4743 3893
rect 4756 3784 4763 3833
rect 4696 3780 4703 3783
rect 4693 3767 4707 3780
rect 4776 3767 4783 3893
rect 4793 3847 4807 3853
rect 4556 3467 4563 3713
rect 4676 3516 4683 3673
rect 4716 3567 4723 3713
rect 4776 3607 4783 3633
rect 4716 3516 4723 3553
rect 4596 3347 4603 3513
rect 4656 3467 4663 3483
rect 4696 3480 4703 3483
rect 4693 3467 4707 3480
rect 4656 3427 4663 3453
rect 4636 3296 4643 3333
rect 4473 2780 4487 2793
rect 4476 2776 4483 2780
rect 4536 2787 4543 3293
rect 4576 3167 4583 3263
rect 4636 2996 4643 3093
rect 4556 2767 4563 2933
rect 4496 2740 4503 2743
rect 4493 2727 4507 2740
rect 4516 2444 4523 2633
rect 4556 2503 4563 2533
rect 4576 2527 4583 2753
rect 4616 2607 4623 2773
rect 4636 2587 4643 2753
rect 4656 2547 4663 2913
rect 4556 2496 4573 2503
rect 4573 2480 4587 2492
rect 4576 2476 4583 2480
rect 4656 2447 4663 2512
rect 4676 2490 4683 3193
rect 4696 2787 4703 3253
rect 4716 3167 4723 3293
rect 4736 3027 4743 3453
rect 4756 3264 4763 3533
rect 4716 2776 4723 2953
rect 4776 2947 4783 3593
rect 4796 3147 4803 3733
rect 4816 2967 4823 3953
rect 4836 3707 4843 4873
rect 4836 3347 4843 3513
rect 4856 3407 4863 4953
rect 4876 4447 4883 5016
rect 4896 4747 4903 5036
rect 4916 4787 4923 4813
rect 4896 4336 4903 4693
rect 4916 4667 4923 4713
rect 4936 4487 4943 4873
rect 4956 4543 4963 5032
rect 4976 4887 4983 5173
rect 4996 4967 5003 5493
rect 5056 5487 5063 5563
rect 5016 4887 5023 5453
rect 5056 5376 5063 5433
rect 5076 5407 5083 5550
rect 5096 5376 5103 5732
rect 5133 5407 5147 5413
rect 5036 4987 5043 5253
rect 5056 5047 5063 5313
rect 5076 5087 5083 5343
rect 5116 5323 5123 5343
rect 5096 5316 5123 5323
rect 5096 5047 5103 5316
rect 5156 5227 5163 5613
rect 5176 5107 5183 5593
rect 5196 5147 5203 5473
rect 5216 5443 5223 5993
rect 5236 5467 5243 6376
rect 5256 6207 5263 6293
rect 5256 6047 5263 6113
rect 5276 5867 5283 6753
rect 5356 6707 5363 6813
rect 5436 6747 5443 7036
rect 5376 6636 5383 6693
rect 5296 6327 5303 6636
rect 5296 6227 5303 6273
rect 5316 6116 5323 6613
rect 5336 6163 5343 6553
rect 5356 6347 5363 6593
rect 5396 6587 5403 6603
rect 5396 6576 5413 6587
rect 5400 6573 5413 6576
rect 5456 6567 5463 7872
rect 5476 7547 5483 8153
rect 5596 8107 5603 8353
rect 5476 7387 5483 7453
rect 5476 7087 5483 7352
rect 5496 7107 5503 7913
rect 5516 7423 5523 8033
rect 5536 7867 5543 8073
rect 5556 7907 5563 8033
rect 5576 7944 5583 8053
rect 5616 8047 5623 8373
rect 5676 8367 5683 8593
rect 5816 8587 5823 8693
rect 5876 8676 5903 8683
rect 5876 8627 5883 8676
rect 5956 8667 5963 9493
rect 5976 9207 5983 9453
rect 6036 9207 6043 9893
rect 6093 9760 6107 9773
rect 6096 9756 6103 9760
rect 6136 9756 6143 10023
rect 6176 9947 6183 10023
rect 6216 9787 6223 10073
rect 6236 9807 6243 10093
rect 6256 10027 6263 10233
rect 5976 8963 5983 9013
rect 5976 8956 6003 8963
rect 5696 8327 5703 8573
rect 5716 8164 5723 8293
rect 5596 8007 5603 8033
rect 5676 7976 5683 8033
rect 5736 7927 5743 8513
rect 5796 8496 5803 8533
rect 5876 8503 5883 8592
rect 5876 8496 5903 8503
rect 5856 8460 5863 8463
rect 5756 8067 5763 8450
rect 5853 8447 5867 8460
rect 5776 8327 5783 8433
rect 5896 8387 5903 8496
rect 5916 8447 5923 8593
rect 5936 8367 5943 8513
rect 5956 8407 5963 8613
rect 5756 7944 5763 7973
rect 5556 7827 5563 7872
rect 5596 7867 5603 7893
rect 5536 7627 5543 7733
rect 5556 7644 5563 7693
rect 5653 7680 5667 7693
rect 5656 7676 5663 7680
rect 5636 7620 5643 7643
rect 5636 7613 5673 7620
rect 5596 7567 5603 7593
rect 5616 7547 5623 7613
rect 5647 7576 5673 7583
rect 5696 7563 5703 7633
rect 5716 7627 5723 7733
rect 5676 7556 5703 7563
rect 5576 7456 5583 7533
rect 5656 7467 5663 7553
rect 5676 7527 5683 7556
rect 5653 7440 5667 7453
rect 5696 7443 5703 7533
rect 5716 7487 5723 7553
rect 5736 7447 5743 7676
rect 5656 7436 5663 7440
rect 5696 7436 5723 7443
rect 5516 7416 5543 7423
rect 5516 7187 5523 7333
rect 5476 6827 5483 7052
rect 5496 6803 5503 7072
rect 5476 6796 5503 6803
rect 5476 6767 5483 6796
rect 5376 6387 5383 6493
rect 5336 6156 5353 6163
rect 5356 6116 5363 6153
rect 5396 6047 5403 6553
rect 5456 6507 5463 6532
rect 5496 6527 5503 6773
rect 5516 6607 5523 7152
rect 5536 7127 5543 7416
rect 5596 7420 5603 7423
rect 5593 7407 5607 7420
rect 5536 6787 5543 7092
rect 5536 6567 5543 6613
rect 5453 6420 5467 6433
rect 5456 6416 5463 6420
rect 5536 6396 5543 6553
rect 5556 6407 5563 7253
rect 5607 7213 5613 7227
rect 5636 7156 5643 7353
rect 5676 7267 5683 7393
rect 5576 6927 5583 7153
rect 5716 7124 5723 7373
rect 5736 7367 5743 7393
rect 5736 7307 5743 7332
rect 5756 7247 5763 7813
rect 5776 7787 5783 8253
rect 5776 7747 5783 7773
rect 5776 7547 5783 7733
rect 5796 7567 5803 8233
rect 5836 7687 5843 8150
rect 5856 7707 5863 7993
rect 5876 7647 5883 8353
rect 5933 8200 5947 8213
rect 5936 8196 5943 8200
rect 5976 8196 5983 8913
rect 5996 8727 6003 8956
rect 6016 8747 6023 8983
rect 6056 8827 6063 9613
rect 6076 9167 6083 9573
rect 6116 9547 6123 9723
rect 6156 9627 6163 9723
rect 6296 9627 6303 10250
rect 6336 10167 6343 10256
rect 6616 10083 6623 10263
rect 6596 10076 6623 10083
rect 6216 9536 6223 9573
rect 6156 9467 6163 9503
rect 6196 9447 6203 9503
rect 6113 9240 6127 9253
rect 6116 9236 6123 9240
rect 6176 9163 6183 9190
rect 6176 9156 6203 9163
rect 6116 8827 6123 9073
rect 6036 8723 6043 8753
rect 6016 8716 6043 8723
rect 5996 8367 6003 8673
rect 5916 8007 5923 8163
rect 5996 7944 6003 8013
rect 5916 7867 5923 7943
rect 6016 7827 6023 8653
rect 5913 7680 5927 7693
rect 5916 7676 5923 7680
rect 6016 7643 6023 7673
rect 5936 7547 5943 7643
rect 5976 7636 6023 7643
rect 6016 7444 6023 7473
rect 6036 7467 6043 8593
rect 6116 8496 6123 8753
rect 6136 8607 6143 9153
rect 6156 8547 6163 8933
rect 6176 8687 6183 9073
rect 6196 8907 6203 9156
rect 6216 9087 6223 9236
rect 6236 9067 6243 9433
rect 6316 9287 6323 9536
rect 6256 9016 6263 9253
rect 6316 9207 6323 9236
rect 6236 8907 6243 8983
rect 6276 8976 6303 8983
rect 6176 8503 6183 8652
rect 6167 8496 6183 8503
rect 6056 8467 6063 8493
rect 6056 8407 6063 8432
rect 6136 8327 6143 8450
rect 5776 7407 5783 7433
rect 6056 7443 6063 7713
rect 6096 7507 6103 8053
rect 6116 7944 6123 8093
rect 6116 7827 6123 7930
rect 6036 7436 6063 7443
rect 6116 7403 6123 7813
rect 6096 7396 6123 7403
rect 5816 7207 5823 7253
rect 5656 7116 5683 7123
rect 5616 6936 5623 7073
rect 5676 6867 5683 7116
rect 5716 6867 5723 6973
rect 5576 6807 5583 6833
rect 5576 6587 5583 6653
rect 5573 6527 5587 6533
rect 5596 6447 5603 6693
rect 5616 6647 5623 6853
rect 5633 6640 5647 6653
rect 5636 6636 5643 6640
rect 5676 6636 5683 6693
rect 5736 6687 5743 7093
rect 5756 6707 5763 7173
rect 5776 6767 5783 7193
rect 5796 6907 5803 7053
rect 5816 7047 5823 7156
rect 5896 7027 5903 7123
rect 5956 7067 5963 7156
rect 5936 7027 5943 7053
rect 5896 6936 5903 6992
rect 5936 6936 5943 6973
rect 5736 6604 5743 6673
rect 5616 6427 5623 6493
rect 5296 5596 5303 5633
rect 5316 5627 5323 5993
rect 5336 5747 5343 6033
rect 5416 6007 5423 6373
rect 5436 5987 5443 6383
rect 5566 6353 5567 6360
rect 5456 6067 5463 6113
rect 5313 5610 5327 5613
rect 5356 5607 5363 5853
rect 5376 5787 5383 5863
rect 5436 5847 5443 5863
rect 5436 5837 5453 5847
rect 5440 5833 5453 5837
rect 5476 5827 5483 6333
rect 5376 5627 5383 5693
rect 5276 5487 5283 5563
rect 5216 5436 5243 5443
rect 5216 5367 5223 5413
rect 5076 4870 5083 4913
rect 5116 4887 5123 5093
rect 4976 4570 4983 4852
rect 5056 4727 5063 4823
rect 5093 4787 5107 4793
rect 4956 4536 4983 4543
rect 4936 4387 4943 4452
rect 4936 4336 4943 4373
rect 4876 3747 4883 4056
rect 4896 3927 4903 4273
rect 4936 3887 4943 4073
rect 4956 3967 4963 4193
rect 4976 4047 4983 4536
rect 4996 4287 5003 4473
rect 5036 4247 5043 4493
rect 5056 4307 5063 4523
rect 5116 4387 5123 4852
rect 5136 4487 5143 5033
rect 5156 4847 5163 4873
rect 5156 4687 5163 4833
rect 5176 4767 5183 4973
rect 5216 4507 5223 5033
rect 5236 5027 5243 5436
rect 5316 5407 5323 5433
rect 5356 5376 5363 5572
rect 5396 5376 5403 5813
rect 5416 5587 5423 5773
rect 5256 5047 5263 5373
rect 5436 5347 5443 5653
rect 5376 5323 5383 5343
rect 5356 5316 5383 5323
rect 5276 4907 5283 5233
rect 5193 4340 5207 4353
rect 5236 4347 5243 4893
rect 5296 4856 5303 5133
rect 5316 5090 5323 5153
rect 5316 4947 5323 5076
rect 5356 4987 5363 5316
rect 5456 5307 5463 5812
rect 5496 5787 5503 6353
rect 5553 6343 5567 6353
rect 5536 6340 5567 6343
rect 5536 6336 5563 6340
rect 5516 6087 5523 6293
rect 5487 5766 5500 5767
rect 5487 5753 5493 5766
rect 5536 5647 5543 6336
rect 5556 5767 5563 6313
rect 5576 6127 5583 6353
rect 5616 6327 5623 6353
rect 5596 6116 5603 6273
rect 5636 6187 5643 6573
rect 5656 6507 5663 6603
rect 5836 6587 5843 6913
rect 5976 6904 5983 7033
rect 5947 6873 5953 6887
rect 5876 6547 5883 6833
rect 5996 6807 6003 7253
rect 6016 7107 6023 7313
rect 6076 7063 6083 7333
rect 6056 7056 6083 7063
rect 6036 6887 6043 6913
rect 6056 6847 6063 7056
rect 6076 6867 6083 6893
rect 5980 6643 5993 6647
rect 5976 6636 5993 6643
rect 5980 6633 5993 6636
rect 5936 6567 5943 6603
rect 5976 6447 5983 6473
rect 5656 6367 5663 6433
rect 5996 6427 6003 6573
rect 5956 6267 5963 6313
rect 5996 6307 6003 6392
rect 6016 6327 6023 6733
rect 6036 6487 6043 6653
rect 6056 6607 6063 6633
rect 5616 5827 5623 6083
rect 5696 6047 5703 6173
rect 5636 5827 5643 5993
rect 5596 5687 5603 5753
rect 5476 5247 5483 5633
rect 5556 5603 5563 5673
rect 5556 5596 5583 5603
rect 5376 5087 5383 5193
rect 5416 5076 5423 5213
rect 5376 4827 5383 5033
rect 5396 5023 5403 5043
rect 5436 5040 5443 5043
rect 5433 5027 5447 5040
rect 5396 5016 5423 5023
rect 5416 4927 5423 5016
rect 5496 4947 5503 5076
rect 5276 4820 5283 4823
rect 5316 4820 5323 4823
rect 5273 4807 5287 4820
rect 5313 4807 5327 4820
rect 5313 4560 5327 4573
rect 5316 4556 5323 4560
rect 5296 4487 5303 4523
rect 5196 4336 5203 4340
rect 5136 4300 5143 4303
rect 5133 4287 5147 4300
rect 5136 4247 5143 4273
rect 5256 4167 5263 4336
rect 5056 4036 5063 4073
rect 5076 4047 5083 4133
rect 5276 4127 5283 4333
rect 5296 4207 5303 4473
rect 5316 4387 5323 4453
rect 5316 4147 5323 4352
rect 5336 4287 5343 4523
rect 5376 4304 5383 4353
rect 5396 4187 5403 4853
rect 5416 4827 5423 4913
rect 5436 4807 5443 4853
rect 5416 4507 5423 4533
rect 5456 4427 5463 4933
rect 5496 4787 5503 4873
rect 5476 4776 5493 4783
rect 5476 4367 5483 4776
rect 5496 4407 5503 4673
rect 5516 4607 5523 5563
rect 5536 5487 5543 5533
rect 5536 4927 5543 5473
rect 5556 4887 5563 5373
rect 5576 4907 5583 5596
rect 5596 5587 5603 5613
rect 5616 5376 5623 5473
rect 5656 5376 5663 6033
rect 5676 5987 5683 6013
rect 5696 5896 5703 5933
rect 5716 5927 5723 5953
rect 5736 5927 5743 6153
rect 5756 6130 5763 6173
rect 5796 6167 5803 6233
rect 5756 5987 5763 6013
rect 5736 5896 5783 5903
rect 5776 5847 5783 5896
rect 5707 5836 5733 5843
rect 5696 5387 5703 5613
rect 5596 4987 5603 5330
rect 5636 5323 5643 5343
rect 5616 5316 5643 5323
rect 5616 4967 5623 5316
rect 5636 5027 5643 5293
rect 5536 4627 5543 4813
rect 5556 4687 5563 4810
rect 5596 4787 5603 4823
rect 5600 4766 5620 4767
rect 5607 4753 5613 4766
rect 5616 4627 5623 4653
rect 5453 4340 5467 4353
rect 5456 4336 5463 4340
rect 5496 4336 5503 4372
rect 5516 4347 5523 4453
rect 5536 4307 5543 4613
rect 5636 4607 5643 4973
rect 5656 4824 5663 5213
rect 5600 4583 5613 4587
rect 5596 4573 5613 4583
rect 5596 4556 5603 4573
rect 5656 4527 5663 4733
rect 5476 4300 5483 4303
rect 5473 4287 5487 4300
rect 4976 3907 4983 3993
rect 4996 3983 5003 4003
rect 4996 3976 5023 3983
rect 4907 3823 4920 3827
rect 4907 3816 4923 3823
rect 4956 3816 4963 3893
rect 4996 3847 5003 3953
rect 4907 3813 4920 3816
rect 4896 3567 4903 3773
rect 4936 3647 4943 3783
rect 4976 3780 4983 3783
rect 4973 3767 4987 3780
rect 5016 3447 5023 3976
rect 5036 3927 5043 4003
rect 5056 3623 5063 3933
rect 5056 3616 5073 3623
rect 4947 3353 4953 3367
rect 4856 3227 4863 3263
rect 4896 3260 4903 3263
rect 4893 3247 4907 3260
rect 4956 3207 4963 3313
rect 4896 3107 4903 3133
rect 4853 3000 4867 3013
rect 4856 2996 4863 3000
rect 4753 2780 4767 2793
rect 4756 2776 4763 2780
rect 4476 2307 4483 2393
rect 4476 2256 4483 2293
rect 4556 2263 4563 2443
rect 4556 2256 4583 2263
rect 4576 2224 4583 2256
rect 4396 2156 4423 2163
rect 4396 2107 4403 2133
rect 4396 1184 4403 1933
rect 4416 1827 4423 2156
rect 4496 2087 4503 2223
rect 4456 1987 4463 2053
rect 4536 2027 4543 2093
rect 4556 2047 4563 2133
rect 4536 1956 4543 2013
rect 4616 2007 4623 2193
rect 4636 2107 4643 2273
rect 4573 1960 4587 1973
rect 4576 1956 4583 1960
rect 4516 1920 4523 1923
rect 4513 1907 4527 1920
rect 4496 1847 4503 1873
rect 4556 1847 4563 1923
rect 4416 1527 4423 1773
rect 4476 1763 4483 1813
rect 4616 1787 4623 1993
rect 4456 1756 4483 1763
rect 4416 1167 4423 1513
rect 4436 930 4443 1413
rect 4456 943 4463 1756
rect 4556 1736 4563 1773
rect 4476 1007 4483 1473
rect 4516 1467 4523 1693
rect 4576 1647 4583 1703
rect 4536 1436 4543 1573
rect 4516 1167 4523 1390
rect 4556 1367 4563 1403
rect 4616 1387 4623 1436
rect 4636 1407 4643 1893
rect 4656 1767 4663 2333
rect 4676 2167 4683 2476
rect 4696 2207 4703 2713
rect 4656 1627 4663 1732
rect 4676 1587 4683 2073
rect 4696 1347 4703 2133
rect 4716 1987 4723 2473
rect 4736 2347 4743 2533
rect 4756 2307 4763 2673
rect 4756 2263 4763 2293
rect 4776 2287 4783 2573
rect 4816 2487 4823 2932
rect 4836 2687 4843 2933
rect 4876 2887 4883 2963
rect 4916 2960 4923 2963
rect 4913 2947 4927 2960
rect 4856 2744 4863 2853
rect 4876 2707 4883 2813
rect 4847 2503 4860 2507
rect 4847 2493 4863 2503
rect 4856 2476 4863 2493
rect 4896 2487 4903 2773
rect 4916 2667 4923 2833
rect 4936 2647 4943 2873
rect 4796 2283 4803 2453
rect 4836 2423 4843 2443
rect 4836 2416 4863 2423
rect 4796 2276 4823 2283
rect 4756 2256 4783 2263
rect 4816 2256 4823 2276
rect 4796 2203 4803 2223
rect 4776 2196 4803 2203
rect 4636 1230 4643 1333
rect 4636 1196 4643 1216
rect 4696 1210 4703 1293
rect 4716 1203 4723 1753
rect 4736 1227 4743 1973
rect 4756 1947 4763 2053
rect 4776 1987 4783 2196
rect 4856 2147 4863 2416
rect 4876 2407 4883 2443
rect 4796 1956 4803 2133
rect 4896 2027 4903 2433
rect 4816 1887 4823 1923
rect 4856 1763 4863 1923
rect 4856 1760 4883 1763
rect 4856 1756 4887 1760
rect 4833 1740 4847 1753
rect 4873 1747 4887 1756
rect 4836 1736 4843 1740
rect 4756 1567 4763 1736
rect 4816 1667 4823 1703
rect 4816 1587 4823 1653
rect 4756 1527 4763 1553
rect 4896 1487 4903 1873
rect 4756 1347 4763 1453
rect 4796 1436 4803 1473
rect 4856 1387 4863 1403
rect 4896 1404 4903 1473
rect 4847 1376 4863 1387
rect 4847 1373 4860 1376
rect 4876 1327 4883 1393
rect 4916 1307 4923 2313
rect 4936 1970 4943 2593
rect 4936 1367 4943 1613
rect 4956 1307 4963 3153
rect 4976 3010 4983 3333
rect 4976 2827 4983 2996
rect 4996 2887 5003 3353
rect 5036 3143 5043 3553
rect 5076 3227 5083 3613
rect 5096 3487 5103 3893
rect 5116 3387 5123 3953
rect 5136 3647 5143 4013
rect 5156 3627 5163 4023
rect 5436 4007 5443 4133
rect 5516 4127 5523 4253
rect 5456 4067 5463 4113
rect 5556 4063 5563 4373
rect 5576 4083 5583 4393
rect 5576 4076 5603 4083
rect 5556 4056 5583 4063
rect 5467 4023 5480 4027
rect 5467 4016 5483 4023
rect 5536 4020 5543 4023
rect 5467 4013 5480 4016
rect 5196 3607 5203 3833
rect 5256 3816 5263 3913
rect 5356 3887 5363 3913
rect 5287 3853 5293 3867
rect 5360 3866 5380 3867
rect 5367 3853 5373 3866
rect 5236 3767 5243 3783
rect 5236 3756 5253 3767
rect 5240 3753 5253 3756
rect 5236 3547 5243 3633
rect 5233 3520 5247 3533
rect 5236 3516 5243 3520
rect 5296 3484 5303 3653
rect 5256 3447 5263 3483
rect 5016 3136 5043 3143
rect 5056 3216 5073 3223
rect 5016 2803 5023 3136
rect 5036 2827 5043 3073
rect 5056 2927 5063 3216
rect 5076 3147 5083 3192
rect 4996 2800 5023 2803
rect 4993 2796 5023 2800
rect 4976 1450 4983 2792
rect 4993 2787 5007 2796
rect 5076 2776 5083 3073
rect 5096 2803 5103 3233
rect 5136 3227 5143 3263
rect 5196 3260 5223 3263
rect 5193 3256 5223 3260
rect 5193 3247 5207 3256
rect 5216 3147 5223 3256
rect 5156 3047 5163 3113
rect 5096 2796 5123 2803
rect 5116 2744 5123 2796
rect 4996 2327 5003 2613
rect 5156 2587 5163 2963
rect 5076 2476 5083 2553
rect 5176 2507 5183 2773
rect 5196 2567 5203 3093
rect 5213 3067 5227 3073
rect 5216 2927 5223 2973
rect 5216 2627 5223 2793
rect 5216 2587 5223 2613
rect 5236 2527 5243 3313
rect 5256 2687 5263 3433
rect 5276 3087 5283 3296
rect 5296 2807 5303 3373
rect 5316 2947 5323 3593
rect 5336 3047 5343 3753
rect 5356 3267 5363 3633
rect 5376 3327 5383 3733
rect 5396 3327 5403 3873
rect 5436 3767 5443 3993
rect 5456 3967 5463 4013
rect 5533 4007 5547 4020
rect 5516 3816 5523 3893
rect 5576 3847 5583 4056
rect 5596 3967 5603 4076
rect 5453 3767 5467 3770
rect 5476 3703 5483 3783
rect 5456 3696 5483 3703
rect 5416 3347 5423 3653
rect 5436 3547 5443 3673
rect 5456 3587 5463 3696
rect 5496 3516 5503 3733
rect 5556 3627 5563 3770
rect 5456 3327 5463 3470
rect 5556 3467 5563 3573
rect 5380 3306 5400 3307
rect 5387 3303 5400 3306
rect 5387 3296 5403 3303
rect 5387 3293 5400 3296
rect 5356 3067 5363 3253
rect 5476 3227 5483 3393
rect 5467 3206 5480 3207
rect 5467 3193 5473 3206
rect 5496 3147 5503 3296
rect 5336 2964 5343 3033
rect 5436 2996 5483 3003
rect 5436 2787 5443 2933
rect 5476 2803 5483 2996
rect 5456 2796 5483 2803
rect 5360 2783 5373 2787
rect 5356 2776 5373 2783
rect 5360 2773 5373 2776
rect 5456 2744 5463 2796
rect 5296 2740 5303 2743
rect 5293 2727 5307 2740
rect 5476 2707 5483 2776
rect 5496 2747 5503 2773
rect 5516 2723 5523 3313
rect 5536 2947 5543 3433
rect 5576 2867 5583 3833
rect 5596 3747 5603 3953
rect 5596 3023 5603 3712
rect 5616 3167 5623 4173
rect 5636 3947 5643 4253
rect 5656 4007 5663 4492
rect 5636 3447 5643 3733
rect 5656 3307 5663 3813
rect 5676 3487 5683 5233
rect 5696 5083 5703 5193
rect 5716 5167 5723 5793
rect 5736 5547 5743 5733
rect 5776 5596 5783 5693
rect 5796 5627 5803 6033
rect 5816 5747 5823 6233
rect 5836 5807 5843 6133
rect 5896 6116 5903 6173
rect 5956 6116 5963 6253
rect 5876 6080 5883 6083
rect 5856 5947 5863 6070
rect 5873 6067 5887 6080
rect 5876 5927 5883 5973
rect 5896 5827 5903 5896
rect 5796 5407 5803 5563
rect 5876 5347 5883 5596
rect 5896 5467 5903 5653
rect 5916 5567 5923 5973
rect 5936 5967 5943 6083
rect 5996 6067 6003 6093
rect 6036 6047 6043 6413
rect 6056 5967 6063 6572
rect 6076 6147 6083 6753
rect 6096 6587 6103 7396
rect 6116 7087 6123 7373
rect 6136 7347 6143 8273
rect 6176 8203 6183 8313
rect 6196 8227 6203 8733
rect 6216 8407 6223 8713
rect 6256 8703 6263 8813
rect 6236 8696 6263 8703
rect 6236 8667 6243 8696
rect 6236 8447 6243 8573
rect 6256 8464 6263 8673
rect 6156 8196 6183 8203
rect 6156 8147 6163 8196
rect 6236 8160 6243 8163
rect 6233 8147 6247 8160
rect 6236 7940 6243 7943
rect 6233 7927 6247 7940
rect 6196 7690 6203 7773
rect 6176 7607 6183 7643
rect 6156 7547 6163 7573
rect 6156 7387 6163 7533
rect 6176 7347 6183 7493
rect 6216 7387 6223 7633
rect 6236 7367 6243 7833
rect 6276 7647 6283 8953
rect 6296 8727 6303 8976
rect 6316 8947 6323 9113
rect 6316 8787 6323 8873
rect 6316 8716 6323 8773
rect 6336 8747 6343 9813
rect 6396 9687 6403 9723
rect 6476 9627 6483 9993
rect 6516 9687 6523 10010
rect 6476 9504 6483 9613
rect 6456 9496 6473 9503
rect 6356 8967 6363 9413
rect 6396 9236 6403 9273
rect 6456 9243 6463 9496
rect 6516 9487 6523 9673
rect 6536 9587 6543 10053
rect 6596 9987 6603 10076
rect 6627 10063 6640 10067
rect 6627 10056 6643 10063
rect 6676 10056 6683 10253
rect 6627 10053 6640 10056
rect 6696 9987 6703 10023
rect 6516 9447 6523 9473
rect 6536 9467 6543 9573
rect 6456 9236 6483 9243
rect 6576 9207 6583 9853
rect 6616 9627 6623 9723
rect 6656 9720 6663 9723
rect 6653 9707 6667 9720
rect 6716 9667 6723 9753
rect 6756 9627 6763 10113
rect 6776 9707 6783 10013
rect 6816 9647 6823 10493
rect 6836 9827 6843 10313
rect 6916 10056 6923 10113
rect 6936 10107 6943 10543
rect 6956 10387 6963 10433
rect 6996 10067 7003 11173
rect 7016 10547 7023 11433
rect 7076 11387 7083 11433
rect 7516 11427 7523 11993
rect 7536 11887 7543 12103
rect 7676 12096 7693 12103
rect 7680 12093 7693 12096
rect 7593 11840 7607 11853
rect 7596 11836 7603 11840
rect 7576 11667 7583 11803
rect 7616 11747 7623 11803
rect 7676 11707 7683 11836
rect 7716 11787 7723 11853
rect 7616 11616 7623 11693
rect 7576 11487 7583 11616
rect 7636 11580 7643 11583
rect 7676 11580 7683 11583
rect 7633 11567 7647 11580
rect 7673 11567 7687 11580
rect 7736 11567 7743 11873
rect 7756 11487 7763 12136
rect 7993 12120 8007 12133
rect 7996 12116 8003 12120
rect 8356 12124 8363 12153
rect 7136 11330 7143 11413
rect 7636 11350 7643 11413
rect 7176 11207 7183 11270
rect 7216 11187 7223 11303
rect 7276 11147 7283 11303
rect 7576 11267 7583 11296
rect 7336 11096 7343 11173
rect 7616 11096 7623 11253
rect 7536 11067 7543 11096
rect 7116 10943 7123 11063
rect 7640 11063 7653 11067
rect 7596 10947 7603 11063
rect 7636 11056 7653 11063
rect 7640 11053 7653 11056
rect 7116 10936 7143 10943
rect 7016 10083 7023 10230
rect 7036 10107 7043 10853
rect 7116 10827 7123 10913
rect 7136 10810 7143 10936
rect 7056 10756 7083 10763
rect 7056 10727 7063 10756
rect 7056 10547 7063 10576
rect 7076 10447 7083 10733
rect 7096 10287 7103 10573
rect 7136 10467 7143 10693
rect 7156 10587 7163 10753
rect 7216 10707 7223 10783
rect 7496 10783 7503 10833
rect 7496 10776 7523 10783
rect 7256 10583 7263 10653
rect 7496 10647 7503 10753
rect 7516 10667 7523 10776
rect 7536 10747 7543 10783
rect 7596 10707 7603 10783
rect 7236 10576 7263 10583
rect 7176 10523 7183 10543
rect 7176 10516 7203 10523
rect 7196 10467 7203 10516
rect 7016 10076 7043 10083
rect 6980 10023 6993 10027
rect 6976 10016 6993 10023
rect 6980 10013 6993 10016
rect 7016 9987 7023 10053
rect 7036 10047 7043 10076
rect 7036 9987 7043 10012
rect 6896 9667 6903 9723
rect 6936 9720 6943 9723
rect 6933 9707 6947 9720
rect 6596 9427 6603 9536
rect 6596 9387 6603 9413
rect 6616 9347 6623 9613
rect 6676 9500 6683 9503
rect 6673 9487 6687 9500
rect 6596 9187 6603 9236
rect 6376 8847 6383 9093
rect 6416 9067 6423 9093
rect 6416 8984 6423 9053
rect 6456 9047 6463 9133
rect 6536 9016 6543 9173
rect 6427 8976 6443 8983
rect 6296 8287 6303 8673
rect 6336 8627 6343 8683
rect 6376 8647 6383 8683
rect 6416 8667 6423 8773
rect 6436 8687 6443 8976
rect 6456 8687 6463 9012
rect 6616 8984 6623 9053
rect 6476 8730 6483 8833
rect 6376 8547 6383 8633
rect 6316 8167 6323 8333
rect 6336 8307 6343 8493
rect 6456 8467 6463 8513
rect 6476 8447 6483 8716
rect 6296 7907 6303 8133
rect 6356 8067 6363 8433
rect 6296 7470 6303 7893
rect 6156 7156 6163 7213
rect 6196 7170 6203 7233
rect 6216 7087 6223 7123
rect 6153 6940 6167 6953
rect 6156 6936 6163 6940
rect 6180 6903 6193 6907
rect 6176 6896 6193 6903
rect 6180 6893 6193 6896
rect 6096 6307 6103 6350
rect 6116 6247 6123 6833
rect 6156 6647 6163 6853
rect 6216 6847 6223 7073
rect 6256 7007 6263 7453
rect 6316 7387 6323 7423
rect 6236 6907 6243 6973
rect 6136 6387 6143 6636
rect 6236 6636 6243 6793
rect 6156 6443 6163 6593
rect 6216 6547 6223 6603
rect 6156 6436 6183 6443
rect 6176 6416 6183 6436
rect 6096 6130 6103 6193
rect 6196 6116 6203 6193
rect 5936 5376 5943 5913
rect 6036 5896 6043 5953
rect 6096 5890 6103 6116
rect 6156 5907 6163 6053
rect 6153 5880 6167 5893
rect 6156 5876 6163 5880
rect 5996 5767 6003 5863
rect 6056 5860 6063 5863
rect 5976 5390 5983 5593
rect 5736 5087 5743 5330
rect 5916 5267 5923 5343
rect 5956 5323 5963 5330
rect 5956 5316 5983 5323
rect 5976 5167 5983 5316
rect 6016 5307 6023 5853
rect 6053 5847 6067 5860
rect 6056 5610 6063 5793
rect 6116 5707 6123 5833
rect 6116 5347 6123 5693
rect 6136 5427 6143 5753
rect 5776 5087 5783 5113
rect 5813 5100 5827 5113
rect 5816 5096 5823 5100
rect 5696 5076 5723 5083
rect 5696 3727 5703 4893
rect 5716 4507 5723 5013
rect 5736 4627 5743 4993
rect 5756 4687 5763 5030
rect 6116 5023 6123 5093
rect 6136 5070 6143 5233
rect 6156 5107 6163 5813
rect 6176 5547 6183 5713
rect 6196 5487 6203 6053
rect 6256 5987 6263 6453
rect 6276 6067 6283 7156
rect 6316 7083 6323 7333
rect 6296 7076 6323 7083
rect 6296 6567 6303 7076
rect 6336 7063 6343 7413
rect 6356 7327 6363 7513
rect 6376 7427 6383 8353
rect 6516 8267 6523 8853
rect 6536 8427 6543 8933
rect 6596 8716 6603 8753
rect 6576 8680 6583 8683
rect 6476 7976 6483 8013
rect 6496 8007 6503 8163
rect 6516 7976 6523 8073
rect 6416 7907 6423 7973
rect 6396 7387 6403 7793
rect 6436 7676 6443 7913
rect 6456 7807 6463 7943
rect 6316 7056 6343 7063
rect 6296 6387 6303 6416
rect 6316 6047 6323 7056
rect 6336 6747 6343 6993
rect 6356 6723 6363 7292
rect 6416 7227 6423 7473
rect 6436 7307 6443 7613
rect 6456 7407 6463 7643
rect 6496 7423 6503 7676
rect 6556 7627 6563 8673
rect 6573 8667 6587 8680
rect 6636 8567 6643 9113
rect 6613 8500 6627 8513
rect 6616 8496 6623 8500
rect 6656 8496 6663 8773
rect 6636 8367 6643 8463
rect 6656 7990 6663 8253
rect 6696 8163 6703 9453
rect 6716 9407 6723 9503
rect 6876 9427 6883 9633
rect 6716 9204 6723 9273
rect 6716 9027 6723 9133
rect 6736 8987 6743 9293
rect 6836 9016 6843 9413
rect 6856 9204 6863 9333
rect 6896 9307 6903 9653
rect 6976 9587 6983 9793
rect 7036 9707 7043 9973
rect 7056 9887 7063 10193
rect 7056 9683 7063 9852
rect 7036 9676 7063 9683
rect 6996 9507 7003 9536
rect 6976 9387 6983 9453
rect 6896 9236 6903 9272
rect 6953 9267 6967 9273
rect 6916 9103 6923 9203
rect 6896 9096 6923 9103
rect 6896 9067 6903 9096
rect 6756 8907 6763 9013
rect 6716 8464 6723 8593
rect 6736 8367 6743 8716
rect 6756 8684 6763 8893
rect 6776 8267 6783 8973
rect 6816 8867 6823 8983
rect 6816 8716 6823 8753
rect 6856 8730 6863 8753
rect 6896 8727 6903 8970
rect 6876 8496 6883 8593
rect 6916 8496 6923 9073
rect 6936 8947 6943 9016
rect 6956 8667 6963 9190
rect 6976 8623 6983 8716
rect 6956 8616 6983 8623
rect 6956 8507 6963 8616
rect 6940 8463 6953 8467
rect 6796 8164 6803 8353
rect 6896 8327 6903 8463
rect 6936 8456 6953 8463
rect 6940 8453 6953 8456
rect 6976 8287 6983 8513
rect 7016 8267 7023 9553
rect 7036 8983 7043 9676
rect 7056 9407 7063 9613
rect 7056 9207 7063 9236
rect 7076 9127 7083 10273
rect 7107 10243 7120 10247
rect 7107 10236 7123 10243
rect 7156 10236 7173 10243
rect 7107 10233 7120 10236
rect 7096 9723 7103 10093
rect 7116 9867 7123 10213
rect 7136 10047 7143 10113
rect 7156 9947 7163 10053
rect 7156 9756 7163 9933
rect 7176 9887 7183 10233
rect 7196 10227 7203 10453
rect 7216 10327 7223 10530
rect 7276 10487 7283 10573
rect 7396 10527 7403 10576
rect 7447 10516 7473 10523
rect 7216 10247 7223 10313
rect 7256 10247 7263 10373
rect 7207 10023 7220 10027
rect 7207 10016 7223 10023
rect 7256 10020 7263 10023
rect 7207 10013 7220 10016
rect 7253 10007 7267 10020
rect 7236 9807 7243 9833
rect 7273 9807 7287 9813
rect 7096 9720 7143 9723
rect 7093 9716 7143 9720
rect 7093 9707 7107 9716
rect 7116 9407 7123 9693
rect 7176 9567 7183 9723
rect 7236 9687 7243 9756
rect 7136 9536 7183 9543
rect 7216 9536 7223 9613
rect 7116 9207 7123 9393
rect 7136 9347 7143 9536
rect 7196 9407 7203 9503
rect 7233 9487 7247 9490
rect 7136 9207 7143 9273
rect 7173 9240 7187 9253
rect 7176 9236 7183 9240
rect 7216 9236 7223 9313
rect 7036 8976 7063 8983
rect 7036 8387 7043 8793
rect 7056 8347 7063 8976
rect 7116 8947 7123 8983
rect 7156 8847 7163 9193
rect 7156 8716 7163 8833
rect 7136 8587 7143 8683
rect 7176 8680 7183 8683
rect 7173 8667 7187 8680
rect 7076 8227 7083 8533
rect 7096 8467 7103 8553
rect 6947 8203 6960 8207
rect 6947 8196 6963 8203
rect 6993 8200 7007 8213
rect 6996 8196 7003 8200
rect 6947 8193 6960 8196
rect 6676 8156 6703 8163
rect 6656 7927 6663 7976
rect 6676 7847 6683 8156
rect 6756 8127 6763 8163
rect 6696 7827 6703 8033
rect 6773 7980 6787 7993
rect 6776 7976 6783 7980
rect 6756 7887 6763 7943
rect 6696 7767 6703 7813
rect 6636 7607 6643 7733
rect 6676 7676 6683 7713
rect 6756 7567 6763 7793
rect 6816 7787 6823 8193
rect 6896 8087 6903 8193
rect 6976 8143 6983 8163
rect 6956 8136 6983 8143
rect 6867 8083 6880 8087
rect 6867 8073 6883 8083
rect 6876 8027 6883 8073
rect 6856 7867 6863 7993
rect 6956 7847 6963 8136
rect 7076 7976 7083 8033
rect 7096 7987 7103 8413
rect 7156 8407 7163 8463
rect 7196 8456 7223 8463
rect 6976 7676 6983 7973
rect 7016 7907 7023 7943
rect 7036 7687 7043 7713
rect 6896 7647 6903 7676
rect 7036 7644 7043 7673
rect 6956 7567 6963 7643
rect 7033 7587 7047 7593
rect 6533 7460 6547 7473
rect 6536 7456 6543 7460
rect 6576 7456 6583 7513
rect 6616 7456 6623 7513
rect 6716 7436 6723 7553
rect 6996 7424 7003 7493
rect 7016 7467 7023 7553
rect 7036 7436 7043 7573
rect 7056 7447 7063 7893
rect 7096 7463 7103 7753
rect 7116 7507 7123 8253
rect 7156 8167 7163 8372
rect 7136 7644 7143 7973
rect 7096 7460 7123 7463
rect 7096 7456 7127 7460
rect 7113 7447 7127 7456
rect 6496 7416 6523 7423
rect 6496 7327 6503 7390
rect 6516 7307 6523 7416
rect 6516 7267 6523 7293
rect 6376 7127 6383 7156
rect 6416 7087 6423 7110
rect 6336 6716 6363 6723
rect 6336 6167 6343 6716
rect 6356 6247 6363 6693
rect 6376 5987 6383 7073
rect 6456 7047 6463 7123
rect 6436 6687 6443 6903
rect 6496 6650 6503 7093
rect 6516 7067 6523 7173
rect 6536 7107 6543 7393
rect 6556 7387 6563 7423
rect 6616 7243 6623 7333
rect 6596 7236 6623 7243
rect 6556 7087 6563 7156
rect 6536 6687 6543 7033
rect 6536 6636 6543 6673
rect 6576 6603 6583 6773
rect 6596 6707 6603 7236
rect 6616 7170 6623 7213
rect 6616 7127 6623 7156
rect 6636 6943 6643 7373
rect 6676 7347 6683 7403
rect 6776 7267 6783 7293
rect 6656 7007 6663 7233
rect 6696 7120 6703 7123
rect 6693 7107 6707 7120
rect 6736 7087 6743 7123
rect 6627 6936 6643 6943
rect 6656 6936 6663 6993
rect 6436 6416 6443 6473
rect 6496 6387 6503 6553
rect 6516 6347 6523 6603
rect 6556 6596 6583 6603
rect 6416 6084 6423 6193
rect 6476 5903 6483 6083
rect 6456 5900 6483 5903
rect 6453 5896 6483 5900
rect 6216 5847 6223 5893
rect 6453 5884 6467 5896
rect 6466 5880 6467 5884
rect 6556 5807 6563 6596
rect 6596 6307 6603 6693
rect 6576 6067 6583 6116
rect 6596 5787 6603 5873
rect 6276 5667 6283 5713
rect 6616 5687 6623 6936
rect 6736 6904 6743 6933
rect 6776 6927 6783 7053
rect 6796 7027 6803 7156
rect 6856 6950 6863 7333
rect 6876 7267 6883 7313
rect 6876 7007 6883 7253
rect 6936 7127 6943 7213
rect 6996 7156 7003 7410
rect 7076 7227 7083 7253
rect 7096 7207 7103 7253
rect 7033 7170 7047 7173
rect 7116 7163 7123 7393
rect 7156 7347 7163 8013
rect 7116 7156 7143 7163
rect 6893 6947 6907 6953
rect 6996 6936 7003 6993
rect 7016 6987 7023 7123
rect 7096 7087 7103 7156
rect 6676 6650 6683 6903
rect 6636 6130 6643 6473
rect 6696 6467 6703 6753
rect 6816 6650 6823 6873
rect 6916 6867 6923 6903
rect 6976 6887 6983 6903
rect 7056 6887 7063 6953
rect 6976 6876 6993 6887
rect 6980 6873 6993 6876
rect 7096 6767 7103 6913
rect 7116 6847 7123 7133
rect 7136 7087 7143 7156
rect 7133 7067 7147 7073
rect 7136 6807 7143 6973
rect 7156 6767 7163 7213
rect 7176 6863 7183 8433
rect 7196 7907 7203 8393
rect 7216 8387 7223 8456
rect 7236 8447 7243 9193
rect 7256 9167 7263 9473
rect 7276 8907 7283 9772
rect 7296 9483 7303 10473
rect 7496 10467 7503 10543
rect 7316 9507 7323 10373
rect 7476 10347 7483 10433
rect 7456 10276 7463 10313
rect 7336 9787 7343 10276
rect 7516 10243 7523 10413
rect 7476 10236 7523 10243
rect 7536 10207 7543 10573
rect 7556 10547 7563 10673
rect 7436 10063 7443 10153
rect 7416 10056 7443 10063
rect 7496 10056 7503 10093
rect 7556 10070 7563 10273
rect 7596 10207 7603 10576
rect 7627 10493 7633 10507
rect 7656 10387 7663 11013
rect 7676 10487 7683 11473
rect 7696 11307 7703 11393
rect 7776 10747 7783 12093
rect 7936 12047 7943 12103
rect 7796 11387 7803 11833
rect 7916 11804 7923 11833
rect 7836 11800 7843 11803
rect 7833 11787 7847 11800
rect 7876 11727 7883 11790
rect 7836 11547 7843 11616
rect 7996 11596 8003 11713
rect 8076 11627 8083 12073
rect 8416 12007 8423 12083
rect 8456 12027 8463 12113
rect 8196 11850 8203 11873
rect 8116 11767 8123 11803
rect 8176 11727 8183 11803
rect 8236 11747 8243 11853
rect 8076 11603 8083 11613
rect 8056 11596 8083 11603
rect 8376 11596 8383 11953
rect 8413 11840 8427 11853
rect 8416 11836 8423 11840
rect 8456 11727 8463 11803
rect 8396 11604 8403 11693
rect 7896 11580 7903 11583
rect 7893 11567 7907 11580
rect 7816 10907 7823 11316
rect 7836 11287 7843 11533
rect 7956 11507 7963 11583
rect 8416 11560 8423 11563
rect 8413 11547 8427 11560
rect 7916 11316 7923 11473
rect 7956 11407 7963 11493
rect 7956 11027 7963 11393
rect 7996 11027 8003 11096
rect 7707 10493 7713 10507
rect 7816 10307 7823 10733
rect 7856 10487 7863 10763
rect 7856 10347 7863 10473
rect 7876 10467 7883 10633
rect 7956 10576 7963 10693
rect 7973 10527 7987 10530
rect 8016 10447 8023 11313
rect 8036 10407 8043 11453
rect 8096 11207 8103 11316
rect 8136 11247 8143 11283
rect 8136 11147 8143 11233
rect 8316 11227 8323 11473
rect 8456 11316 8463 11393
rect 8493 11320 8507 11333
rect 8496 11316 8503 11320
rect 8056 10687 8063 10793
rect 7776 10260 7783 10263
rect 7773 10247 7787 10260
rect 7876 10263 7883 10393
rect 8076 10387 8083 11133
rect 8156 11123 8163 11153
rect 8136 11116 8163 11123
rect 8136 11096 8143 11116
rect 8116 10847 8123 11050
rect 8216 10927 8223 11093
rect 8256 10927 8263 11013
rect 8216 10827 8223 10913
rect 8133 10800 8147 10813
rect 8136 10796 8143 10800
rect 8116 10667 8123 10763
rect 8216 10590 8223 10813
rect 8236 10647 8243 10796
rect 8256 10667 8263 10913
rect 8276 10764 8283 10793
rect 8256 10576 8263 10653
rect 8316 10627 8323 11213
rect 8376 11110 8383 11293
rect 8436 11280 8443 11283
rect 8433 11267 8447 11280
rect 8476 11227 8483 11283
rect 8536 11267 8543 11836
rect 8556 11824 8563 12173
rect 8687 12163 8700 12167
rect 8687 12153 8703 12163
rect 8696 12136 8703 12153
rect 8956 12136 9003 12143
rect 8636 12047 8643 12103
rect 8736 12007 8743 12136
rect 8996 12116 9003 12136
rect 9056 12116 9063 12173
rect 9096 12104 9103 12153
rect 9376 12147 9383 12193
rect 9367 12136 9383 12147
rect 9367 12133 9380 12136
rect 8556 11627 8563 11810
rect 8556 11247 8563 11613
rect 8576 11307 8583 11993
rect 8936 11967 8943 12103
rect 9416 12076 9443 12083
rect 9476 12080 9483 12083
rect 9392 12027 9399 12073
rect 9436 12067 9443 12076
rect 9473 12067 9487 12080
rect 8696 11836 8703 11873
rect 8616 11584 8623 11713
rect 8716 11687 8723 11803
rect 8756 11800 8763 11803
rect 8753 11787 8767 11800
rect 8816 11787 8823 11893
rect 8936 11847 8943 11953
rect 9436 11887 9443 12053
rect 9500 12027 9507 12073
rect 9796 12047 9803 12153
rect 9836 12116 9843 12213
rect 10416 12136 10423 12193
rect 9893 12120 9907 12133
rect 9896 12116 9903 12120
rect 9936 12027 9943 12110
rect 10456 12104 10463 12173
rect 10996 12136 11043 12143
rect 10136 12100 10143 12103
rect 10133 12087 10147 12100
rect 8976 11836 8983 11873
rect 8956 11787 8963 11803
rect 8676 11636 8743 11643
rect 8676 11616 8683 11636
rect 8736 11623 8743 11636
rect 8736 11616 8763 11623
rect 8956 11616 8963 11773
rect 9016 11623 9023 11833
rect 8996 11616 9023 11623
rect 8696 11580 8703 11583
rect 8693 11567 8707 11580
rect 8756 11567 8763 11616
rect 8596 11347 8603 11553
rect 8696 11527 8703 11553
rect 8736 11350 8743 11533
rect 8496 11076 8503 11153
rect 8556 11076 8563 11233
rect 8396 11027 8403 11063
rect 8436 10927 8443 11063
rect 8456 10987 8463 11053
rect 8596 10847 8603 11333
rect 8733 11320 8747 11336
rect 8736 11316 8743 11320
rect 8656 11284 8663 11313
rect 8796 11300 8803 11303
rect 8793 11287 8807 11300
rect 8856 11247 8863 11303
rect 8876 11167 8883 11273
rect 8896 11207 8903 11616
rect 8936 11487 8943 11583
rect 8976 11527 8983 11583
rect 9156 11467 9163 11836
rect 9216 11783 9223 11803
rect 9296 11787 9303 11836
rect 9216 11776 9273 11783
rect 9236 11616 9243 11693
rect 9276 11616 9283 11693
rect 9216 11580 9223 11583
rect 9213 11567 9227 11580
rect 9216 11350 9223 11373
rect 9256 11307 9263 11393
rect 9016 11110 9023 11193
rect 8616 11047 8623 11070
rect 8916 11007 8923 11043
rect 8636 10796 8643 10933
rect 8736 10927 8743 10973
rect 8707 10816 8713 10827
rect 8700 10813 8713 10816
rect 8416 10760 8423 10763
rect 8413 10747 8427 10760
rect 8236 10467 8243 10543
rect 8276 10540 8283 10543
rect 8273 10527 8287 10540
rect 8176 10307 8183 10373
rect 8196 10327 8203 10433
rect 8416 10367 8423 10533
rect 8436 10527 8443 10553
rect 8456 10387 8463 10793
rect 8556 10576 8563 10673
rect 8496 10487 8503 10543
rect 8476 10407 8483 10473
rect 8496 10427 8503 10473
rect 8516 10447 8523 10513
rect 8616 10387 8623 10733
rect 8196 10296 8203 10313
rect 8253 10300 8267 10313
rect 8256 10296 8263 10300
rect 7856 10256 7883 10263
rect 7676 10167 7683 10230
rect 7356 10024 7363 10053
rect 7376 10007 7383 10053
rect 7296 9476 7323 9483
rect 7296 9204 7303 9313
rect 7316 9183 7323 9476
rect 7356 9243 7363 9753
rect 7296 9176 7323 9183
rect 7336 9236 7363 9243
rect 7296 8967 7303 9176
rect 7336 9167 7343 9236
rect 7336 9030 7343 9153
rect 7356 9127 7363 9213
rect 7376 9207 7383 9873
rect 7396 9827 7403 9953
rect 7416 9767 7423 10056
rect 7436 9947 7443 9993
rect 7436 9807 7443 9933
rect 7476 9883 7483 10023
rect 7576 10020 7583 10023
rect 7573 10007 7587 10020
rect 7456 9876 7483 9883
rect 7456 9827 7463 9876
rect 7556 9867 7563 9973
rect 7456 9756 7463 9792
rect 7416 9607 7423 9732
rect 7556 9724 7563 9793
rect 7476 9627 7483 9723
rect 7476 9500 7483 9503
rect 7473 9487 7487 9500
rect 7516 9387 7523 9503
rect 7516 9327 7523 9373
rect 7476 9236 7483 9273
rect 7296 8607 7303 8713
rect 7316 8464 7323 8493
rect 7256 8196 7263 8253
rect 7216 7944 7223 8033
rect 7276 7987 7283 8163
rect 7256 7944 7263 7973
rect 7193 7567 7207 7573
rect 7196 7147 7203 7513
rect 7216 7450 7223 7493
rect 7216 7327 7223 7436
rect 7236 7267 7243 7456
rect 7216 7047 7223 7173
rect 7236 7107 7243 7193
rect 7256 7167 7263 7613
rect 7276 7407 7283 7593
rect 7296 7527 7303 7633
rect 7316 7603 7323 7676
rect 7336 7627 7343 8953
rect 7356 7607 7363 8893
rect 7376 8730 7383 8983
rect 7456 8887 7463 9203
rect 7416 8716 7423 8753
rect 7496 8684 7503 8733
rect 7396 8567 7403 8683
rect 7436 8527 7443 8573
rect 7376 8047 7383 8493
rect 7476 8443 7483 8463
rect 7456 8436 7483 8443
rect 7456 8407 7463 8436
rect 7396 7647 7403 8333
rect 7456 8067 7463 8333
rect 7476 7943 7483 8413
rect 7456 7936 7483 7943
rect 7316 7596 7343 7603
rect 7336 7456 7343 7596
rect 7416 7567 7423 7733
rect 7353 7487 7367 7493
rect 7416 7467 7423 7513
rect 7436 7447 7443 7893
rect 7293 7424 7307 7433
rect 7273 7160 7287 7173
rect 7276 7156 7283 7160
rect 7316 7156 7323 7213
rect 7336 7187 7343 7393
rect 7416 7207 7423 7353
rect 7436 7227 7443 7393
rect 7456 7187 7463 7936
rect 7496 7907 7503 8433
rect 7516 8387 7523 8453
rect 7536 8447 7543 9493
rect 7556 8427 7563 9593
rect 7576 9387 7583 9533
rect 7596 9016 7603 9793
rect 7616 9047 7623 9913
rect 7636 9867 7643 10023
rect 7696 9927 7703 10193
rect 7836 10127 7843 10250
rect 7807 10063 7820 10067
rect 7807 10056 7823 10063
rect 7800 10053 7823 10056
rect 7636 9107 7643 9756
rect 7676 9727 7683 9853
rect 7693 9847 7707 9853
rect 7816 9807 7823 10053
rect 7836 9770 7843 10092
rect 7716 9647 7723 9723
rect 7656 9487 7663 9633
rect 7856 9607 7863 10256
rect 8156 10127 8163 10263
rect 7916 9827 7923 10073
rect 7876 9687 7883 9753
rect 7936 9707 7943 10113
rect 8016 10056 8023 10093
rect 8176 10070 8183 10253
rect 7996 10007 8003 10023
rect 7996 9867 8003 9993
rect 8036 9927 8043 10023
rect 8216 9967 8223 10173
rect 8236 9947 8243 10113
rect 8276 10103 8283 10233
rect 8296 10127 8303 10263
rect 8276 10096 8303 10103
rect 8296 10056 8303 10096
rect 8276 10020 8283 10023
rect 8316 10020 8323 10023
rect 8273 10007 8287 10020
rect 8313 10007 8327 10020
rect 8376 10007 8383 10113
rect 8576 10063 8583 10373
rect 8656 10307 8663 10763
rect 8716 10523 8723 10613
rect 8736 10544 8743 10873
rect 8716 10516 8743 10523
rect 8576 10056 8603 10063
rect 8396 10027 8403 10056
rect 8496 9947 8503 10056
rect 8036 9807 8043 9913
rect 8116 9787 8123 9873
rect 8556 9787 8563 10010
rect 8216 9747 8223 9773
rect 8093 9724 8107 9730
rect 8016 9667 8023 9723
rect 7707 9543 7720 9547
rect 7707 9536 7723 9543
rect 7707 9533 7720 9536
rect 8033 9540 8047 9553
rect 8036 9536 8043 9540
rect 7676 9504 7683 9533
rect 7976 9504 7983 9533
rect 7656 9407 7663 9473
rect 7736 9467 7743 9503
rect 8056 9500 8063 9503
rect 8053 9487 8067 9500
rect 7676 9227 7683 9393
rect 7716 9236 7723 9373
rect 7756 9147 7763 9203
rect 8096 9187 8103 9216
rect 7616 8747 7623 8983
rect 7676 8716 7683 8793
rect 7716 8716 7723 8773
rect 7616 8684 7623 8712
rect 7756 8687 7763 9033
rect 7576 8267 7583 8553
rect 7596 8367 7603 8473
rect 7616 8347 7623 8513
rect 7656 8227 7663 8533
rect 7756 8496 7763 8613
rect 7796 8547 7803 9133
rect 8116 9107 8123 9433
rect 8136 9270 8143 9733
rect 8156 9707 8163 9743
rect 8156 9287 8163 9693
rect 8196 9504 8203 9613
rect 8216 9347 8223 9553
rect 8296 9536 8303 9633
rect 8316 9500 8323 9503
rect 8313 9487 8327 9500
rect 8256 9224 8263 9273
rect 8216 9107 8223 9223
rect 7913 9000 7927 9013
rect 7916 8996 7923 9000
rect 8296 8996 8303 9353
rect 8336 9147 8343 9413
rect 8316 9004 8323 9053
rect 8356 9003 8363 9333
rect 8356 8996 8383 9003
rect 7836 8523 7843 8973
rect 7856 8767 7863 8983
rect 8376 8903 8383 8996
rect 8396 8964 8403 9253
rect 8336 8896 8383 8903
rect 7973 8720 7987 8733
rect 7976 8716 7983 8720
rect 8053 8727 8067 8733
rect 7876 8587 7883 8670
rect 7956 8607 7963 8683
rect 7836 8516 7853 8523
rect 7856 8476 7863 8513
rect 7716 8267 7723 8463
rect 7896 8407 7903 8593
rect 7916 8447 7923 8476
rect 8176 8476 8183 8833
rect 8216 8716 8223 8753
rect 8196 8484 8203 8573
rect 8236 8547 8243 8683
rect 8253 8447 8267 8453
rect 8196 8436 8223 8443
rect 7536 8160 7543 8163
rect 7533 8147 7547 8160
rect 7536 8027 7543 8133
rect 7556 7847 7563 8053
rect 7496 7787 7503 7833
rect 7496 7676 7503 7773
rect 7556 7747 7563 7833
rect 7576 7827 7583 8163
rect 7596 7947 7603 8153
rect 7616 8107 7623 8183
rect 7676 8180 7683 8183
rect 7673 8167 7687 8180
rect 7716 8147 7723 8253
rect 8036 8216 8043 8293
rect 8176 8283 8183 8393
rect 8196 8327 8203 8436
rect 8276 8387 8283 8673
rect 8156 8276 8183 8283
rect 8076 8187 8083 8273
rect 8000 8183 8013 8187
rect 7996 8176 8013 8183
rect 7973 8167 7987 8176
rect 8000 8173 8013 8176
rect 7973 8160 7993 8167
rect 7976 8156 7993 8160
rect 7980 8153 7993 8156
rect 7596 7727 7603 7933
rect 7636 7707 7643 8013
rect 7733 7960 7747 7973
rect 7736 7956 7743 7960
rect 7676 7907 7683 7943
rect 7656 7896 7673 7903
rect 7516 7607 7523 7643
rect 7556 7607 7563 7663
rect 7296 7087 7303 7123
rect 7336 7120 7343 7123
rect 7333 7107 7347 7120
rect 7236 7027 7243 7072
rect 7216 6936 7223 6973
rect 7256 6936 7263 6973
rect 7236 6887 7243 6903
rect 7227 6876 7243 6887
rect 7227 6873 7240 6876
rect 7176 6856 7203 6863
rect 6876 6656 6883 6693
rect 6716 6607 6723 6636
rect 6756 6507 6763 6603
rect 6767 6496 6783 6503
rect 6653 6423 6667 6433
rect 6653 6420 6683 6423
rect 6656 6416 6683 6420
rect 6716 6416 6723 6473
rect 6696 6380 6703 6383
rect 6736 6380 6743 6383
rect 6693 6367 6707 6380
rect 6733 6367 6747 6380
rect 6776 6367 6783 6496
rect 6296 5596 6303 5633
rect 6540 5623 6553 5627
rect 6536 5613 6553 5623
rect 6536 5596 6543 5613
rect 6316 5527 6323 5563
rect 6216 5376 6223 5433
rect 6196 5127 6203 5330
rect 6116 5016 6133 5023
rect 6136 4987 6143 5013
rect 6176 4987 6183 5063
rect 6187 4976 6203 4983
rect 5776 4767 5783 4953
rect 5816 4856 5823 4893
rect 5856 4856 5863 4973
rect 5913 4927 5927 4933
rect 5756 4507 5763 4673
rect 5776 4647 5783 4753
rect 5796 4667 5803 4753
rect 5896 4687 5903 4713
rect 5876 4627 5883 4653
rect 5776 4467 5783 4593
rect 5856 4587 5863 4613
rect 5827 4583 5840 4587
rect 5827 4573 5843 4583
rect 5836 4556 5843 4573
rect 5816 4520 5823 4523
rect 5813 4507 5827 4520
rect 5893 4507 5907 4513
rect 5867 4477 5893 4484
rect 5916 4467 5923 4653
rect 5736 4336 5743 4373
rect 5796 4336 5803 4433
rect 5716 4187 5723 4213
rect 5756 4087 5763 4233
rect 5776 4050 5783 4213
rect 5796 4187 5803 4273
rect 5856 4207 5863 4452
rect 5916 4247 5923 4373
rect 5936 4307 5943 4873
rect 5956 4447 5963 4893
rect 5976 4527 5983 4913
rect 5996 4507 6003 4733
rect 6016 4547 6023 4613
rect 6036 4507 6043 4810
rect 5896 4236 5913 4243
rect 5813 4040 5827 4053
rect 5816 4036 5823 4040
rect 5696 3407 5703 3692
rect 5716 3527 5723 4033
rect 5756 4000 5763 4003
rect 5753 3987 5767 4000
rect 5756 3927 5763 3973
rect 5796 3907 5803 4003
rect 5876 3987 5883 4033
rect 5776 3780 5783 3783
rect 5773 3767 5787 3780
rect 5856 3767 5863 3893
rect 5876 3787 5883 3933
rect 5736 3516 5743 3593
rect 5776 3516 5783 3553
rect 5796 3547 5803 3713
rect 5876 3707 5883 3733
rect 5896 3503 5903 4236
rect 5916 4067 5923 4173
rect 5916 3747 5923 4053
rect 5936 3830 5943 4073
rect 5936 3567 5943 3773
rect 5896 3496 5923 3503
rect 5800 3483 5813 3487
rect 5756 3447 5763 3483
rect 5796 3476 5813 3483
rect 5800 3473 5813 3476
rect 5676 3296 5683 3353
rect 5716 3296 5723 3373
rect 5656 3167 5663 3193
rect 5776 3187 5783 3313
rect 5796 3167 5803 3293
rect 5816 3264 5823 3333
rect 5816 3187 5823 3213
rect 5596 3016 5623 3023
rect 5596 2807 5603 2996
rect 5593 2780 5607 2793
rect 5616 2787 5623 3016
rect 5656 2996 5663 3033
rect 5756 3027 5763 3073
rect 5740 3006 5760 3007
rect 5740 3003 5753 3006
rect 5736 2996 5753 3003
rect 5740 2993 5753 2996
rect 5596 2776 5603 2780
rect 5496 2716 5523 2723
rect 5496 2627 5503 2716
rect 5193 2500 5207 2513
rect 5196 2496 5203 2500
rect 5036 2427 5043 2476
rect 5007 2296 5033 2303
rect 4996 1807 5003 2093
rect 5016 1587 5023 2153
rect 5076 2107 5083 2256
rect 5096 2127 5103 2443
rect 5136 2067 5143 2443
rect 4993 1407 5007 1413
rect 4716 1196 4743 1203
rect 4576 1180 4583 1183
rect 4573 1167 4587 1180
rect 4456 936 4483 943
rect 4476 916 4483 936
rect 4536 884 4543 973
rect 4556 863 4563 1153
rect 4536 856 4563 863
rect 3976 507 3983 663
rect 4016 656 4063 663
rect 3776 384 3783 493
rect 4096 416 4103 573
rect 4116 547 4123 673
rect 3596 207 3603 363
rect 3736 307 3743 383
rect 3633 180 3647 193
rect 3636 176 3643 180
rect 3676 144 3683 193
rect 3916 144 3923 213
rect 2836 107 2843 130
rect 2496 36 2515 43
rect 3096 -17 3103 143
rect 3076 -24 3103 -17
rect 3336 -24 3343 143
rect 3596 -24 3603 143
rect 3876 136 3913 143
rect 4036 127 4043 173
rect 4056 67 4063 383
rect 4076 107 4083 213
rect 4136 176 4143 376
rect 4176 176 4183 393
rect 4236 190 4243 696
rect 4416 665 4423 713
rect 4436 667 4443 696
rect 4296 507 4303 533
rect 4296 364 4303 493
rect 4416 176 4423 413
rect 4116 140 4123 143
rect 4113 127 4127 140
rect 4236 107 4243 176
rect 4496 167 4503 453
rect 4516 407 4523 733
rect 4536 647 4543 856
rect 4596 710 4603 993
rect 4656 884 4663 913
rect 4536 307 4543 453
rect 4556 327 4563 693
rect 4616 647 4623 663
rect 4647 653 4653 667
rect 4616 447 4623 633
rect 4576 407 4583 433
rect 4676 427 4683 1153
rect 4736 1047 4743 1196
rect 5016 1196 5023 1473
rect 5036 1407 5043 1956
rect 5196 1924 5203 2433
rect 5096 1787 5103 1923
rect 5216 1707 5223 2153
rect 5236 2067 5243 2463
rect 5496 2464 5503 2493
rect 5516 2367 5523 2693
rect 5536 2507 5543 2573
rect 5636 2507 5643 2953
rect 5436 2224 5443 2253
rect 5140 1703 5153 1707
rect 5096 1647 5103 1703
rect 5136 1696 5153 1703
rect 5140 1693 5153 1696
rect 5076 1436 5083 1633
rect 5036 1287 5043 1393
rect 5076 1204 5083 1273
rect 5056 1143 5063 1163
rect 5056 1136 5083 1143
rect 4733 920 4747 933
rect 4776 930 4783 1033
rect 4736 916 4743 920
rect 4816 887 4823 933
rect 4996 916 5003 1073
rect 5016 1047 5023 1113
rect 5033 920 5047 933
rect 5036 916 5043 920
rect 4716 607 4723 883
rect 4836 647 4843 913
rect 4976 747 4983 883
rect 4976 697 4983 733
rect 4867 663 4880 667
rect 5016 665 5023 713
rect 5036 667 5043 833
rect 4867 656 4883 663
rect 4867 653 4880 656
rect 4856 567 4863 613
rect 5076 587 5083 1136
rect 5116 1027 5123 1213
rect 5116 747 5123 1013
rect 5136 987 5143 1473
rect 5156 1087 5163 1653
rect 5176 1147 5183 1573
rect 5236 1404 5243 1753
rect 5256 1383 5263 2013
rect 5296 1807 5303 2193
rect 5316 2187 5323 2223
rect 5336 1924 5343 2193
rect 5376 2007 5383 2073
rect 5376 1956 5383 1993
rect 5456 1970 5463 2313
rect 5476 2167 5483 2353
rect 5576 2256 5583 2433
rect 5616 2327 5623 2463
rect 5613 2260 5627 2273
rect 5616 2256 5623 2260
rect 5316 1916 5333 1923
rect 5276 1704 5283 1773
rect 5236 1376 5263 1383
rect 4593 400 4607 413
rect 4596 396 4603 400
rect 4796 390 4803 453
rect 5116 416 5123 573
rect 5176 547 5183 916
rect 5216 723 5223 1353
rect 5236 1007 5243 1376
rect 5276 1216 5283 1553
rect 5316 1507 5323 1916
rect 5496 1767 5503 2256
rect 5596 2220 5603 2223
rect 5593 2207 5607 2220
rect 5656 2207 5663 2933
rect 5676 2927 5683 2963
rect 5716 2960 5723 2963
rect 5713 2947 5727 2960
rect 5676 2707 5683 2913
rect 5696 2827 5703 2893
rect 5676 2327 5683 2633
rect 5696 2407 5703 2773
rect 5716 2527 5723 2853
rect 5596 2167 5603 2193
rect 5516 1727 5523 2093
rect 5576 1924 5583 2093
rect 5596 1704 5603 1773
rect 5636 1763 5643 2113
rect 5676 2107 5683 2313
rect 5716 2127 5723 2492
rect 5676 1956 5683 2013
rect 5716 1970 5723 2013
rect 5736 1963 5743 2793
rect 5756 2647 5763 2873
rect 5836 2807 5843 3353
rect 5856 3264 5863 3453
rect 5876 3167 5883 3473
rect 5893 3467 5907 3473
rect 5756 2287 5763 2633
rect 5776 2490 5783 2773
rect 5796 2667 5803 2793
rect 5856 2790 5863 3033
rect 5836 2727 5843 2743
rect 5896 2727 5903 3353
rect 5836 2717 5853 2727
rect 5840 2713 5853 2717
rect 5856 2567 5863 2692
rect 5856 2476 5863 2553
rect 5896 2487 5903 2713
rect 5916 2647 5923 3496
rect 5936 3447 5943 3532
rect 5956 3467 5963 4353
rect 5956 3296 5963 3373
rect 5976 3367 5983 4453
rect 6016 4387 6023 4453
rect 6036 4336 6043 4472
rect 6056 4447 6063 4913
rect 6136 4887 6143 4952
rect 6160 4863 6173 4867
rect 6156 4856 6173 4863
rect 6160 4853 6173 4856
rect 6116 4787 6123 4823
rect 6176 4787 6183 4813
rect 6076 4727 6083 4773
rect 6176 4707 6183 4752
rect 6076 4567 6083 4613
rect 6196 4607 6203 4976
rect 6236 4907 6243 5063
rect 6256 4827 6263 4973
rect 6216 4627 6223 4713
rect 6116 4556 6123 4593
rect 6236 4587 6243 4810
rect 6256 4687 6263 4753
rect 6276 4667 6283 5473
rect 6087 4523 6100 4527
rect 6087 4516 6103 4523
rect 6087 4513 6100 4516
rect 6073 4487 6087 4492
rect 5996 3827 6003 4293
rect 6056 4247 6063 4303
rect 6073 4287 6087 4290
rect 6016 3947 6023 4073
rect 6076 4067 6083 4213
rect 6096 4187 6103 4493
rect 6113 4387 6127 4393
rect 6116 4123 6123 4333
rect 6136 4327 6143 4523
rect 6176 4467 6183 4533
rect 6196 4487 6203 4543
rect 6116 4116 6143 4123
rect 6076 3967 6083 4003
rect 6116 3907 6123 4033
rect 6016 3816 6023 3893
rect 6136 3887 6143 4116
rect 6056 3816 6063 3853
rect 6076 3780 6083 3783
rect 5996 3727 6003 3770
rect 6073 3767 6087 3780
rect 5996 3527 6003 3593
rect 6013 3520 6027 3533
rect 6016 3516 6023 3520
rect 6056 3516 6063 3613
rect 6076 3607 6083 3713
rect 6036 3327 6043 3483
rect 6076 3407 6083 3483
rect 6096 3387 6103 3473
rect 6016 3227 6023 3263
rect 6056 3247 6063 3333
rect 5976 3107 5983 3153
rect 5976 2996 5983 3093
rect 6016 2996 6023 3133
rect 5936 2827 5943 2993
rect 6096 2964 6103 3033
rect 5796 2307 5803 2453
rect 5916 2444 5923 2573
rect 5836 2387 5843 2443
rect 5756 2187 5763 2273
rect 5776 2207 5783 2253
rect 5816 2027 5823 2223
rect 5736 1956 5763 1963
rect 5696 1787 5703 1923
rect 5636 1756 5663 1763
rect 5656 1736 5663 1756
rect 5376 1607 5383 1703
rect 5336 1436 5343 1473
rect 5316 1216 5323 1273
rect 5376 1184 5383 1233
rect 5456 1227 5463 1513
rect 5616 1436 5623 1473
rect 5556 1347 5563 1403
rect 5296 1107 5303 1183
rect 5287 943 5300 947
rect 5287 933 5303 943
rect 5296 916 5303 933
rect 5336 916 5343 1133
rect 5276 787 5283 883
rect 5396 787 5403 973
rect 5216 716 5243 723
rect 5236 696 5243 716
rect 5276 567 5283 673
rect 4616 307 4623 363
rect 4696 327 4703 383
rect 4716 287 4723 373
rect 5156 387 5163 473
rect 4436 107 4443 143
rect 4676 -17 4683 143
rect 4756 67 4763 370
rect 5196 190 5203 453
rect 5216 176 5223 433
rect 5296 364 5303 733
rect 5456 727 5463 1213
rect 5516 1184 5523 1233
rect 5536 1230 5543 1253
rect 5596 1247 5603 1403
rect 5567 1243 5580 1247
rect 5567 1233 5583 1243
rect 5576 1216 5583 1233
rect 5496 1176 5513 1183
rect 5496 696 5503 1176
rect 5596 1127 5603 1183
rect 5596 983 5603 1033
rect 5616 1007 5623 1073
rect 5596 976 5623 983
rect 5616 916 5623 976
rect 5656 916 5663 953
rect 5536 827 5543 916
rect 5416 190 5423 513
rect 5456 207 5463 663
rect 5556 307 5563 393
rect 5460 183 5473 187
rect 5456 176 5473 183
rect 5460 173 5473 176
rect 4656 -24 4683 -17
rect 4916 -24 4923 143
rect 5176 -24 5183 143
rect 5496 27 5503 193
rect 5516 107 5523 173
rect 5576 47 5583 733
rect 5596 667 5603 883
rect 5636 711 5643 870
rect 5636 696 5643 697
rect 5696 696 5703 1293
rect 5736 1167 5743 1433
rect 5756 767 5763 1956
rect 5776 1667 5783 1953
rect 5776 884 5783 1433
rect 5796 1404 5803 1773
rect 5816 1447 5823 1973
rect 5836 1567 5843 1736
rect 5856 1470 5863 1993
rect 5876 1527 5883 2373
rect 5916 1987 5923 2430
rect 5936 2047 5943 2513
rect 5956 2227 5963 2913
rect 5976 2727 5983 2776
rect 5996 2707 6003 2963
rect 6116 2927 6123 3733
rect 6136 2807 6143 3813
rect 6156 2967 6163 3993
rect 6176 3487 6183 4293
rect 6196 3463 6203 4433
rect 6216 4227 6223 4533
rect 6216 3887 6223 4036
rect 6216 3667 6223 3793
rect 6236 3527 6243 4413
rect 6253 4387 6267 4393
rect 6276 4387 6283 4453
rect 6256 4047 6263 4352
rect 6276 4343 6283 4373
rect 6296 4367 6303 5373
rect 6316 4827 6323 5273
rect 6336 4967 6343 5153
rect 6356 4863 6363 5573
rect 6560 5563 6573 5567
rect 6556 5556 6573 5563
rect 6560 5553 6573 5556
rect 6436 5376 6443 5473
rect 6347 4856 6363 4863
rect 6376 4856 6383 4893
rect 6336 4727 6343 4853
rect 6476 4767 6483 5043
rect 6436 4647 6443 4753
rect 6556 4687 6563 5533
rect 6636 5447 6643 5973
rect 6676 5847 6683 6293
rect 6796 6207 6803 6603
rect 6836 6467 6843 6603
rect 6896 6367 6903 6613
rect 6916 6387 6923 6623
rect 7176 6627 7183 6653
rect 7196 6423 7203 6856
rect 7216 6667 7223 6833
rect 7276 6767 7283 6903
rect 7316 6667 7323 7013
rect 7187 6416 7203 6423
rect 7216 6416 7223 6613
rect 7236 6527 7243 6623
rect 7296 6467 7303 6610
rect 6816 6087 6823 6116
rect 6776 6067 6783 6083
rect 6767 6056 6783 6067
rect 6767 6053 6780 6056
rect 6696 5707 6703 6033
rect 6773 5900 6787 5913
rect 6776 5896 6783 5900
rect 6716 5767 6723 5850
rect 6736 5747 6743 5773
rect 6756 5767 6763 5829
rect 6796 5787 6803 5863
rect 6673 5610 6687 5613
rect 6576 4827 6583 5433
rect 6696 5376 6703 5672
rect 6736 5383 6743 5733
rect 6793 5600 6807 5613
rect 6796 5596 6803 5600
rect 6756 5447 6763 5553
rect 6776 5487 6783 5563
rect 6816 5560 6823 5563
rect 6813 5547 6827 5560
rect 6736 5376 6763 5383
rect 6616 5087 6623 5376
rect 6756 5344 6763 5376
rect 6796 5347 6803 5513
rect 6876 5347 6883 6233
rect 6916 6167 6923 6253
rect 6956 6247 6963 6373
rect 6996 6363 7003 6383
rect 7176 6384 7183 6413
rect 6976 6356 7003 6363
rect 6936 6007 6943 6193
rect 6976 6047 6983 6356
rect 7016 6167 7023 6333
rect 7036 6247 7043 6373
rect 7016 6116 7023 6153
rect 7060 6143 7073 6147
rect 7056 6133 7073 6143
rect 7056 6130 7063 6133
rect 7116 6083 7123 6253
rect 7316 6187 7323 6613
rect 7336 6587 7343 6893
rect 7356 6867 7363 7113
rect 7376 6867 7383 7143
rect 7436 7136 7463 7143
rect 7396 6847 7403 6973
rect 7356 6567 7363 6753
rect 7376 6624 7383 6713
rect 7347 6473 7353 6487
rect 7076 6076 7123 6083
rect 7076 5896 7083 6033
rect 7120 5903 7133 5907
rect 7116 5896 7133 5903
rect 7016 5727 7023 5896
rect 7120 5893 7133 5896
rect 7056 5727 7063 5863
rect 7156 5863 7163 6013
rect 7147 5856 7163 5863
rect 6896 5547 6903 5633
rect 7047 5623 7060 5627
rect 7047 5613 7063 5623
rect 7056 5596 7063 5613
rect 6916 5391 6923 5433
rect 7076 5387 7083 5563
rect 6676 5287 6683 5343
rect 6656 5087 6663 5133
rect 6656 4856 6663 5073
rect 6316 4507 6323 4573
rect 6547 4443 6560 4447
rect 6547 4433 6563 4443
rect 6276 4336 6303 4343
rect 6316 4300 6323 4303
rect 6313 4287 6327 4300
rect 6307 3996 6323 4003
rect 6176 3456 6203 3463
rect 6176 3143 6183 3456
rect 6256 3296 6263 3873
rect 6296 3830 6303 3953
rect 6316 3827 6323 3996
rect 6276 3647 6283 3713
rect 6296 3587 6303 3816
rect 6336 3816 6343 4193
rect 6356 3967 6363 4213
rect 6376 3987 6383 4273
rect 6436 4267 6443 4393
rect 6396 3947 6403 4253
rect 6456 3947 6463 4373
rect 6556 4336 6563 4433
rect 6476 4227 6483 4336
rect 6416 3823 6423 3933
rect 6416 3816 6443 3823
rect 6340 3763 6360 3767
rect 6340 3760 6353 3763
rect 6336 3753 6353 3760
rect 6336 3707 6343 3753
rect 6296 3547 6303 3573
rect 6376 3563 6383 3693
rect 6396 3647 6403 3783
rect 6436 3763 6443 3816
rect 6416 3756 6443 3763
rect 6356 3556 6383 3563
rect 6293 3520 6307 3533
rect 6356 3527 6363 3556
rect 6296 3516 6303 3520
rect 6196 3167 6203 3293
rect 6236 3260 6243 3263
rect 6233 3247 6247 3260
rect 6176 3136 6203 3143
rect 6116 2707 6123 2743
rect 6156 2727 6163 2833
rect 6176 2744 6183 2793
rect 5976 2307 5983 2673
rect 5996 2007 6003 2633
rect 6016 2567 6023 2593
rect 6136 2476 6143 2553
rect 6176 2476 6183 2593
rect 6196 2507 6203 3136
rect 6236 2996 6243 3153
rect 6276 3127 6283 3263
rect 5973 1960 5987 1973
rect 5976 1956 5983 1960
rect 5916 1920 5923 1923
rect 5913 1907 5927 1920
rect 5956 1787 5963 1923
rect 5896 1607 5903 1733
rect 5936 1667 5943 1690
rect 5976 1567 5983 1703
rect 6016 1683 6023 2473
rect 6116 2327 6123 2443
rect 6093 2260 6107 2273
rect 6096 2256 6103 2260
rect 6036 1867 6043 2013
rect 5996 1676 6023 1683
rect 5836 1180 5843 1183
rect 5876 1180 5883 1183
rect 5833 1167 5847 1180
rect 5873 1167 5887 1180
rect 5916 1167 5923 1433
rect 5616 396 5623 453
rect 5680 403 5693 407
rect 5676 396 5693 403
rect 5680 393 5693 396
rect 5716 364 5723 393
rect 5636 147 5643 313
rect 5676 176 5683 213
rect 5736 207 5743 663
rect 5756 327 5763 393
rect 5776 144 5783 693
rect 5796 223 5803 1153
rect 5816 884 5823 1013
rect 5896 1007 5903 1113
rect 5896 916 5903 993
rect 5816 307 5823 373
rect 5836 227 5843 493
rect 5896 410 5903 753
rect 5916 627 5923 773
rect 5936 430 5943 1453
rect 5996 1267 6003 1676
rect 6056 1443 6063 2033
rect 6076 1987 6083 2223
rect 6096 1467 6103 1910
rect 6116 1587 6123 2213
rect 6136 1647 6143 2373
rect 6156 1607 6163 2443
rect 6216 2287 6223 2773
rect 6236 2667 6243 2773
rect 6236 2263 6243 2430
rect 6227 2256 6243 2263
rect 6216 1956 6223 2252
rect 6256 1970 6263 2963
rect 6276 2267 6283 2813
rect 6276 2087 6283 2253
rect 6236 1920 6243 1923
rect 6233 1907 6247 1920
rect 6236 1736 6243 1853
rect 6276 1747 6283 2073
rect 6036 1436 6063 1443
rect 6096 1436 6103 1453
rect 5996 967 6003 1253
rect 6016 930 6023 1213
rect 6016 696 6023 916
rect 6036 847 6043 1436
rect 6136 1287 6143 1453
rect 6156 1407 6163 1593
rect 6176 1347 6183 1693
rect 6256 1700 6263 1703
rect 6253 1687 6267 1700
rect 6096 1216 6103 1273
rect 6116 1007 6123 1183
rect 6156 1047 6163 1183
rect 6216 1087 6223 1353
rect 6156 916 6163 993
rect 6196 887 6203 1033
rect 6236 747 6243 1633
rect 6276 987 6283 1693
rect 6296 1307 6303 2653
rect 6316 2387 6323 2973
rect 6336 2907 6343 3483
rect 6356 2947 6363 3213
rect 6376 2987 6383 3513
rect 6416 3503 6423 3756
rect 6396 3496 6423 3503
rect 6336 2827 6343 2893
rect 6376 2776 6383 2913
rect 6396 2807 6403 3496
rect 6416 2903 6423 3473
rect 6436 2927 6443 3733
rect 6456 3667 6463 3816
rect 6476 3643 6483 4173
rect 6496 4087 6503 4233
rect 6536 4207 6543 4303
rect 6587 4253 6593 4267
rect 6636 4227 6643 4493
rect 6516 4036 6523 4093
rect 6596 4083 6603 4213
rect 6596 4076 6613 4083
rect 6496 3767 6503 3953
rect 6456 3636 6483 3643
rect 6416 2896 6443 2903
rect 6353 2727 6367 2730
rect 6396 2687 6403 2743
rect 6436 2647 6443 2896
rect 6456 2787 6463 3636
rect 6516 3527 6523 3973
rect 6576 3807 6583 4053
rect 6616 4007 6623 4073
rect 6636 3947 6643 4192
rect 6656 3827 6663 4613
rect 6676 4547 6683 4633
rect 6556 3516 6563 3593
rect 6576 3567 6583 3793
rect 6676 3727 6683 4290
rect 6696 4067 6703 4893
rect 6716 4827 6723 4856
rect 6736 4667 6743 5113
rect 6696 4007 6703 4032
rect 6716 3967 6723 4576
rect 6756 4227 6763 5013
rect 6776 4967 6783 5043
rect 6816 5007 6823 5043
rect 6916 4927 6923 5377
rect 6776 4467 6783 4913
rect 6816 4827 6823 4856
rect 6796 4343 6803 4813
rect 6836 4687 6843 4813
rect 6816 4507 6823 4673
rect 6876 4627 6883 4823
rect 6936 4647 6943 5333
rect 7056 5340 7063 5343
rect 7053 5327 7067 5340
rect 7096 5307 7103 5377
rect 6976 4587 6983 4856
rect 7016 4824 7023 4993
rect 6896 4407 6903 4483
rect 6776 4336 6803 4343
rect 6776 4207 6783 4336
rect 6916 4307 6923 4336
rect 6796 4147 6803 4253
rect 6816 4247 6823 4303
rect 6856 4267 6863 4303
rect 6796 4036 6803 4073
rect 6696 3747 6703 3816
rect 6716 3727 6723 3932
rect 6667 3706 6680 3707
rect 6667 3693 6673 3706
rect 6736 3687 6743 3993
rect 6776 3947 6783 4003
rect 6856 3847 6863 4193
rect 6876 4007 6883 4233
rect 6896 4187 6903 4293
rect 6916 3907 6923 4213
rect 6576 3447 6583 3483
rect 6616 3310 6623 3470
rect 6476 3203 6483 3233
rect 6496 3227 6503 3263
rect 6476 3196 6513 3203
rect 6496 2996 6503 3173
rect 6356 2387 6363 2553
rect 6416 2547 6423 2613
rect 6427 2493 6433 2507
rect 6416 2476 6423 2493
rect 6376 2256 6383 2333
rect 6356 2220 6363 2223
rect 6353 2207 6367 2220
rect 6396 2167 6403 2223
rect 6336 1907 6343 2153
rect 6356 1707 6363 2073
rect 6456 1956 6463 2033
rect 6496 1956 6503 2793
rect 6516 2667 6523 2963
rect 6516 2467 6523 2513
rect 6536 2443 6543 2933
rect 6556 2707 6563 3213
rect 6596 2776 6603 2950
rect 6656 2867 6663 3293
rect 6676 3264 6683 3513
rect 6716 3227 6723 3533
rect 6736 3087 6743 3673
rect 6756 3307 6763 3813
rect 6796 3530 6803 3833
rect 6816 3784 6823 3813
rect 6827 3693 6833 3707
rect 6896 3687 6903 3783
rect 6836 3516 6843 3653
rect 6856 3480 6863 3483
rect 6853 3467 6867 3480
rect 6776 3187 6783 3263
rect 6796 2967 6803 3253
rect 6836 3207 6843 3233
rect 6616 2687 6623 2743
rect 6653 2727 6667 2730
rect 6516 2436 6543 2443
rect 6516 2167 6523 2436
rect 6536 2207 6543 2393
rect 6556 2223 6563 2672
rect 6673 2480 6687 2493
rect 6676 2476 6683 2480
rect 6656 2387 6663 2443
rect 6696 2440 6703 2443
rect 6693 2427 6707 2440
rect 6616 2256 6623 2333
rect 6556 2216 6583 2223
rect 6376 1807 6383 1853
rect 6316 1667 6323 1693
rect 6356 1436 6363 1573
rect 6316 1027 6323 1213
rect 6336 1187 6343 1403
rect 6416 1247 6423 1953
rect 6556 1924 6563 2013
rect 6436 1827 6443 1893
rect 6436 1227 6443 1813
rect 6516 1787 6523 1923
rect 6420 1223 6433 1227
rect 6416 1216 6433 1223
rect 6420 1213 6433 1216
rect 6256 867 6263 893
rect 6296 747 6303 773
rect 6236 696 6243 733
rect 5876 327 5883 363
rect 5916 327 5923 363
rect 5976 247 5983 663
rect 6196 660 6223 663
rect 6193 656 6223 660
rect 6193 647 6207 656
rect 6276 416 6283 573
rect 6316 447 6323 913
rect 6456 887 6463 1773
rect 6496 1687 6503 1703
rect 6576 1687 6583 2216
rect 6596 2207 6603 2223
rect 6636 2220 6643 2223
rect 6633 2207 6647 2220
rect 6596 2047 6603 2193
rect 6487 1676 6503 1687
rect 6487 1673 6500 1676
rect 6376 847 6383 883
rect 6456 527 6463 693
rect 6476 664 6483 1053
rect 6516 807 6523 1673
rect 6596 1647 6603 1956
rect 6616 1927 6623 2113
rect 6556 1247 6563 1533
rect 6596 1487 6603 1513
rect 6596 1436 6603 1473
rect 6636 1450 6643 1733
rect 6676 1627 6683 2153
rect 6656 1347 6663 1403
rect 6696 1287 6703 2253
rect 6716 2187 6723 2333
rect 6716 2027 6723 2173
rect 6736 1963 6743 2473
rect 6756 2087 6763 2953
rect 6836 2927 6843 3033
rect 6776 2444 6783 2813
rect 6796 2067 6803 2853
rect 6816 2407 6823 2893
rect 6816 2107 6823 2313
rect 6836 2127 6843 2653
rect 6856 2227 6863 3432
rect 6876 2907 6883 3296
rect 6896 2964 6903 2993
rect 6916 2810 6923 3473
rect 6936 3447 6943 4453
rect 6956 3487 6963 4293
rect 6976 4007 6983 4573
rect 7016 4407 7023 4810
rect 7036 4569 7043 4933
rect 7056 4907 7063 5043
rect 7116 4887 7123 5693
rect 7136 5027 7143 5850
rect 7176 4947 7183 6173
rect 7287 6143 7300 6147
rect 7287 6133 7303 6143
rect 7196 5787 7203 6133
rect 7296 6116 7303 6133
rect 7396 6087 7403 6673
rect 7276 6080 7283 6083
rect 7273 6067 7287 6080
rect 7196 4927 7203 5713
rect 7216 5487 7223 5993
rect 7276 5967 7283 6053
rect 7316 5910 7323 6073
rect 7216 5090 7223 5173
rect 7216 5047 7223 5076
rect 7216 4887 7223 4973
rect 7036 4427 7043 4555
rect 7016 4187 7023 4393
rect 7056 4307 7063 4872
rect 7076 4407 7083 4773
rect 7096 4767 7103 4853
rect 7216 4824 7223 4873
rect 7096 4607 7103 4732
rect 7096 4527 7103 4593
rect 7136 4556 7143 4593
rect 7173 4560 7187 4573
rect 7176 4556 7183 4560
rect 7236 4527 7243 5813
rect 7256 5667 7263 5893
rect 7356 5767 7363 5850
rect 7376 5727 7383 5793
rect 7396 5727 7403 6052
rect 7416 5827 7423 7133
rect 7436 6347 7443 7113
rect 7456 7067 7463 7136
rect 7456 6787 7463 6993
rect 7476 6907 7483 7493
rect 7516 7424 7523 7593
rect 7536 7527 7543 7553
rect 7536 7407 7543 7513
rect 7556 7347 7563 7533
rect 7576 7487 7583 7553
rect 7656 7467 7663 7896
rect 7836 7847 7843 7956
rect 8116 7956 8123 8173
rect 8136 7964 8143 8033
rect 8156 7983 8163 8276
rect 8176 8087 8183 8213
rect 8156 7980 8183 7983
rect 8156 7976 8187 7980
rect 8173 7967 8187 7976
rect 8196 7927 8203 8313
rect 8136 7916 8153 7923
rect 7956 7707 7963 7833
rect 7973 7700 7987 7713
rect 7976 7696 7983 7700
rect 7676 7627 7683 7693
rect 8056 7667 8063 7793
rect 8136 7727 8143 7916
rect 7736 7436 7743 7513
rect 7576 7307 7583 7433
rect 7616 7367 7623 7423
rect 7607 7353 7623 7367
rect 7616 7327 7623 7353
rect 7776 7287 7783 7453
rect 8056 7436 8063 7653
rect 8076 7567 8083 7673
rect 8116 7444 8123 7513
rect 8096 7367 8103 7403
rect 8136 7367 8143 7713
rect 8156 7643 8163 7813
rect 8216 7747 8223 8373
rect 8276 8196 8283 8333
rect 8316 8210 8323 8893
rect 8336 8407 8343 8896
rect 8356 8247 8363 8793
rect 8376 8267 8383 8450
rect 8416 8367 8423 9573
rect 8456 9236 8463 9533
rect 8476 9467 8483 9743
rect 8496 9487 8503 9653
rect 8596 9587 8603 10056
rect 8616 9707 8623 10263
rect 8676 10260 8703 10263
rect 8676 10256 8707 10260
rect 8693 10247 8707 10256
rect 8533 9540 8547 9553
rect 8536 9536 8543 9540
rect 8636 9507 8643 10193
rect 8696 9507 8703 10212
rect 8716 9790 8723 10273
rect 8736 10227 8743 10516
rect 8756 10127 8763 10933
rect 8776 10847 8783 10893
rect 8776 10207 8783 10833
rect 8876 10827 8883 10993
rect 8956 10987 8963 11073
rect 8796 10764 8803 10793
rect 8816 10540 8823 10543
rect 8813 10527 8827 10540
rect 8876 10287 8883 10813
rect 8976 10796 8983 10953
rect 8936 10687 8943 10763
rect 8916 10276 8923 10473
rect 9016 10187 9023 11096
rect 9056 11047 9063 11153
rect 9176 11096 9183 11253
rect 9156 10907 9163 11063
rect 9196 11043 9203 11063
rect 9187 11036 9203 11043
rect 9116 10590 9123 10813
rect 9176 10747 9183 11033
rect 9256 10927 9263 11093
rect 9276 11007 9283 11373
rect 9296 11267 9303 11316
rect 9416 11284 9423 11693
rect 9436 11387 9443 11873
rect 9496 11867 9503 11893
rect 9973 11860 9987 11873
rect 9976 11856 9983 11860
rect 9496 11836 9503 11853
rect 10016 11847 10023 11993
rect 9556 11820 9563 11823
rect 9553 11807 9567 11820
rect 9473 11787 9487 11790
rect 9513 11620 9527 11633
rect 9516 11616 9523 11620
rect 9496 11316 9503 11413
rect 9656 11284 9663 11553
rect 9736 11547 9743 11583
rect 9776 11507 9783 11583
rect 9773 11320 9787 11333
rect 9776 11316 9783 11320
rect 9476 11280 9483 11283
rect 9473 11267 9487 11280
rect 9476 11060 9483 11063
rect 9473 11047 9487 11060
rect 9476 10967 9483 11033
rect 9427 10836 9453 10843
rect 9216 10796 9223 10833
rect 9433 10800 9447 10813
rect 9473 10800 9487 10813
rect 9436 10796 9443 10800
rect 9476 10796 9483 10800
rect 9536 10767 9543 11113
rect 9556 11110 9563 11133
rect 9056 10487 9063 10543
rect 8736 9787 8743 10056
rect 8733 9760 8747 9773
rect 8736 9756 8743 9760
rect 8776 9756 8783 9993
rect 8796 9927 8803 10023
rect 8836 9767 8843 10023
rect 8476 9200 8483 9203
rect 8473 9187 8487 9200
rect 8436 8687 8443 9033
rect 8456 8767 8463 9016
rect 8516 8767 8523 9203
rect 8556 9167 8563 9490
rect 8576 9187 8583 9236
rect 8596 9107 8603 9503
rect 8596 9016 8603 9053
rect 8616 9047 8623 9493
rect 8756 9407 8763 9723
rect 8776 9527 8783 9633
rect 8796 9547 8803 9723
rect 8836 9667 8843 9753
rect 8876 9750 8883 10053
rect 8896 9927 8903 10113
rect 8816 9536 8823 9573
rect 8856 9536 8863 9593
rect 8633 9020 8647 9033
rect 8656 9027 8663 9273
rect 8736 9250 8743 9273
rect 8836 9263 8843 9503
rect 8896 9467 8903 9573
rect 8916 9267 8923 10093
rect 8956 9567 8963 10173
rect 9036 10024 9043 10293
rect 9096 10244 9103 10373
rect 9156 10276 9163 10473
rect 9096 10107 9103 10230
rect 9116 9927 9123 10023
rect 9056 9756 9063 9813
rect 8773 9240 8787 9253
rect 8816 9256 8843 9263
rect 8776 9236 8783 9240
rect 8696 9183 8703 9236
rect 8696 9176 8723 9183
rect 8636 9016 8643 9020
rect 8576 8827 8583 8983
rect 8636 8827 8643 8873
rect 8676 8843 8683 9093
rect 8696 8947 8703 9153
rect 8656 8836 8683 8843
rect 8456 8716 8503 8723
rect 8536 8716 8543 8793
rect 8456 8683 8463 8716
rect 8596 8687 8603 8753
rect 8456 8676 8483 8683
rect 8476 8496 8483 8676
rect 8516 8587 8523 8683
rect 8516 8496 8523 8533
rect 8556 8527 8563 8670
rect 8656 8647 8663 8836
rect 8716 8827 8723 9176
rect 8736 9107 8743 9173
rect 8736 8984 8743 9093
rect 8616 8567 8623 8613
rect 8676 8467 8683 8813
rect 8756 8787 8763 9203
rect 8816 9067 8823 9256
rect 8776 8887 8783 9053
rect 8796 8867 8803 8996
rect 8816 8907 8823 9032
rect 8816 8827 8823 8893
rect 8836 8747 8843 9233
rect 8876 9016 8883 9073
rect 8916 9016 8923 9232
rect 8956 9147 8963 9553
rect 8976 9327 8983 9533
rect 8996 9247 9003 9713
rect 9036 9504 9043 9613
rect 9076 9407 9083 9503
rect 9156 9407 9163 9756
rect 9176 9587 9183 10230
rect 9176 9507 9183 9573
rect 9196 9427 9203 10013
rect 9016 9236 9023 9353
rect 9056 9236 9063 9273
rect 9013 9000 9027 9013
rect 9016 8996 9023 9000
rect 8896 8927 8903 8983
rect 8456 8460 8463 8463
rect 8453 8447 8467 8460
rect 8696 8463 8703 8670
rect 8796 8647 8803 8683
rect 8776 8496 8783 8553
rect 8696 8456 8723 8463
rect 8656 8327 8663 8353
rect 8676 8347 8683 8453
rect 8396 8216 8403 8313
rect 8420 8227 8427 8273
rect 8256 8107 8263 8163
rect 8236 7847 8243 8013
rect 8376 8010 8383 8173
rect 8696 8143 8703 8213
rect 8716 8187 8723 8456
rect 8816 8427 8823 8513
rect 8796 8416 8813 8423
rect 8796 8227 8803 8416
rect 8736 8176 8763 8183
rect 8696 8140 8723 8143
rect 8696 8136 8727 8140
rect 8713 8127 8727 8136
rect 8236 7676 8243 7773
rect 8156 7636 8183 7643
rect 7496 7127 7503 7173
rect 7736 7107 7743 7136
rect 7656 6916 7663 7033
rect 7836 7027 7843 7273
rect 7856 7147 7863 7273
rect 7893 7203 7907 7213
rect 7893 7200 7923 7203
rect 7896 7196 7923 7200
rect 7867 7093 7873 7107
rect 7896 7047 7903 7176
rect 7916 7067 7923 7196
rect 7956 7067 7963 7293
rect 8116 7267 8123 7313
rect 8076 7170 8083 7253
rect 7993 7107 8007 7113
rect 7516 6900 7523 6903
rect 7556 6900 7563 6903
rect 7513 6887 7527 6900
rect 7553 6887 7567 6900
rect 7696 6887 7703 7013
rect 7976 6947 7983 7093
rect 7996 6923 8003 6953
rect 8036 6927 8043 7033
rect 7976 6916 8003 6923
rect 7476 6587 7483 6872
rect 8056 6883 8063 7053
rect 8036 6876 8063 6883
rect 8036 6863 8043 6876
rect 8016 6856 8043 6863
rect 7476 6487 7483 6573
rect 7496 6487 7503 6733
rect 7516 6607 7523 6852
rect 7576 6650 7583 6753
rect 7616 6647 7623 6793
rect 7556 6507 7563 6603
rect 7596 6600 7603 6603
rect 7593 6587 7607 6600
rect 7436 5867 7443 6273
rect 7416 5687 7423 5753
rect 7276 5207 7283 5563
rect 7356 5547 7363 5653
rect 7356 5376 7363 5433
rect 7380 5343 7393 5347
rect 7336 5323 7343 5343
rect 7376 5336 7393 5343
rect 7380 5333 7393 5336
rect 7336 5316 7363 5323
rect 7327 5293 7333 5307
rect 7356 5247 7363 5316
rect 7296 5076 7303 5133
rect 7356 5083 7363 5113
rect 7336 5076 7363 5083
rect 7276 5007 7283 5043
rect 7156 4503 7163 4523
rect 7256 4503 7263 4933
rect 7156 4496 7183 4503
rect 7136 4336 7143 4393
rect 7116 4147 7123 4253
rect 6996 4007 7003 4093
rect 7076 4067 7083 4133
rect 6953 3447 6967 3452
rect 6976 3387 6983 3413
rect 6976 3187 6983 3373
rect 6996 3267 7003 3953
rect 7016 3707 7023 3993
rect 7036 3907 7043 4003
rect 7016 3387 7023 3633
rect 7036 3427 7043 3893
rect 7056 3547 7063 3833
rect 7116 3816 7123 3873
rect 7136 3847 7143 4273
rect 7156 3947 7163 4073
rect 7176 3967 7183 4496
rect 7236 4496 7263 4503
rect 7196 4127 7203 4393
rect 7236 4247 7243 4496
rect 7276 4247 7283 4713
rect 7296 4287 7303 4913
rect 7316 4267 7323 4810
rect 7376 4487 7383 5273
rect 7396 4947 7403 5233
rect 7416 4887 7423 5313
rect 7436 4967 7443 5813
rect 7456 5327 7463 6433
rect 7456 5044 7463 5133
rect 7476 5027 7483 6416
rect 7533 6130 7547 6133
rect 7573 6120 7587 6133
rect 7576 6116 7583 6120
rect 7516 6027 7523 6083
rect 7556 6080 7563 6083
rect 7553 6067 7567 6080
rect 7616 5987 7623 6573
rect 7636 6567 7643 6813
rect 7656 6727 7663 6793
rect 7676 6687 7683 6773
rect 7636 6467 7643 6513
rect 7636 6267 7643 6416
rect 7656 6147 7663 6633
rect 7696 6507 7703 6636
rect 7516 5347 7523 5896
rect 7553 5600 7567 5613
rect 7556 5596 7563 5600
rect 7616 5596 7623 5653
rect 7576 5427 7583 5563
rect 7656 5507 7663 6112
rect 7676 5747 7683 6373
rect 7696 5787 7703 6493
rect 7676 5707 7683 5733
rect 7576 5383 7583 5413
rect 7676 5407 7683 5593
rect 7556 5376 7583 5383
rect 7676 5383 7683 5393
rect 7656 5376 7683 5383
rect 7513 5327 7527 5333
rect 7556 5327 7563 5376
rect 7516 5043 7523 5292
rect 7576 5076 7583 5293
rect 7596 5187 7603 5343
rect 7636 5307 7643 5343
rect 7636 5267 7643 5293
rect 7696 5287 7703 5433
rect 7516 5036 7543 5043
rect 7413 4860 7427 4873
rect 7416 4856 7423 4860
rect 7456 4856 7463 4913
rect 7496 4887 7503 4953
rect 7493 4860 7507 4873
rect 7496 4856 7503 4860
rect 7476 4767 7483 4823
rect 7496 4627 7503 4693
rect 7433 4560 7447 4573
rect 7436 4556 7443 4560
rect 7416 4427 7423 4523
rect 7393 4340 7407 4353
rect 7396 4336 7403 4340
rect 7376 4283 7383 4303
rect 7356 4276 7383 4283
rect 7156 3867 7163 3912
rect 7196 3907 7203 4013
rect 7236 3887 7243 4053
rect 7176 3776 7193 3783
rect 7076 3516 7083 3573
rect 7116 3547 7123 3713
rect 7196 3627 7203 3773
rect 7113 3520 7127 3533
rect 7116 3516 7123 3520
rect 7096 3447 7103 3483
rect 7036 3296 7043 3333
rect 7056 3247 7063 3263
rect 7047 3236 7063 3247
rect 7047 3233 7060 3236
rect 7033 3107 7047 3113
rect 7016 2996 7023 3033
rect 6996 2947 7003 2963
rect 6896 2740 6903 2743
rect 6893 2727 6907 2740
rect 6996 2587 7003 2933
rect 7016 2607 7023 2793
rect 7036 2587 7043 2693
rect 6916 2270 6923 2430
rect 6936 2256 6943 2393
rect 6716 1956 6743 1963
rect 6756 1956 6763 2033
rect 6796 1970 6803 1993
rect 6716 1747 6723 1956
rect 6816 1920 6823 1923
rect 6813 1907 6827 1920
rect 6836 1867 6843 1913
rect 6856 1827 6863 2013
rect 6856 1707 6863 1733
rect 6536 787 6543 1213
rect 6576 883 6583 1216
rect 6596 930 6603 1233
rect 6653 1220 6667 1233
rect 6656 1216 6663 1220
rect 6636 1147 6643 1183
rect 6676 1147 6683 1183
rect 6696 923 6703 1153
rect 6676 916 6703 923
rect 6576 876 6603 883
rect 6507 703 6520 707
rect 6507 696 6523 703
rect 6556 696 6563 833
rect 6596 727 6603 876
rect 6616 863 6623 883
rect 6616 856 6643 863
rect 6593 700 6607 713
rect 6596 696 6603 700
rect 6507 693 6520 696
rect 6576 660 6583 663
rect 6573 647 6587 660
rect 6636 627 6643 856
rect 6656 687 6663 883
rect 6676 627 6683 793
rect 6716 483 6723 1093
rect 6736 1067 6743 1703
rect 6776 1667 6783 1703
rect 6756 1107 6763 1613
rect 6876 1487 6883 2053
rect 6896 1750 6903 2223
rect 6916 1867 6923 2213
rect 6816 1127 6823 1453
rect 6776 867 6783 973
rect 6736 507 6743 853
rect 6756 647 6763 773
rect 6816 747 6823 913
rect 6836 727 6843 1473
rect 6856 1247 6863 1473
rect 6896 1467 6903 1736
rect 6936 1704 6943 1833
rect 6956 1647 6963 2113
rect 6916 1436 6923 1553
rect 6976 1407 6983 2153
rect 6996 1967 7003 2533
rect 7016 2447 7023 2513
rect 7036 1956 7043 2333
rect 7056 2167 7063 3213
rect 7096 3147 7103 3253
rect 7116 3107 7123 3296
rect 7136 3107 7143 3133
rect 7076 2907 7083 2973
rect 7156 2947 7163 3353
rect 7076 2787 7083 2893
rect 7176 2887 7183 3533
rect 7196 3227 7203 3613
rect 7216 3003 7223 3713
rect 7236 3227 7243 3633
rect 7196 2996 7223 3003
rect 7236 2996 7243 3113
rect 7256 3027 7263 4173
rect 7276 3923 7283 4233
rect 7356 4087 7363 4276
rect 7276 3916 7303 3923
rect 7276 3647 7283 3893
rect 7296 3727 7303 3916
rect 7336 3887 7343 3953
rect 7376 3787 7383 4253
rect 7416 4147 7423 4253
rect 7396 4004 7403 4033
rect 7436 3830 7443 4433
rect 7456 4007 7463 4393
rect 7476 4350 7483 4573
rect 7496 4367 7503 4613
rect 7416 3727 7423 3783
rect 7456 3780 7463 3783
rect 7453 3767 7467 3780
rect 7276 3347 7283 3533
rect 7353 3520 7367 3533
rect 7356 3516 7363 3520
rect 7496 3487 7503 4213
rect 7396 3447 7403 3483
rect 7333 3300 7347 3313
rect 7336 3296 7343 3300
rect 7396 3264 7403 3393
rect 7356 3243 7363 3263
rect 7336 3236 7363 3243
rect 7273 3000 7287 3013
rect 7276 2996 7283 3000
rect 7196 2847 7203 2996
rect 7256 2960 7263 2963
rect 7253 2947 7267 2960
rect 7076 2647 7083 2733
rect 7096 2667 7103 2773
rect 7176 2687 7183 2743
rect 7096 2027 7103 2553
rect 7136 2444 7143 2513
rect 7216 2490 7223 2730
rect 7236 2527 7243 2833
rect 7156 2327 7163 2433
rect 7256 2387 7263 2776
rect 7116 2127 7123 2293
rect 7156 2187 7163 2223
rect 7080 1963 7093 1967
rect 7076 1956 7093 1963
rect 7080 1953 7093 1956
rect 7016 1827 7023 1923
rect 7056 1847 7063 1923
rect 7007 1743 7020 1747
rect 7007 1736 7023 1743
rect 7053 1740 7067 1753
rect 7056 1736 7063 1740
rect 7007 1733 7020 1736
rect 7076 1700 7083 1703
rect 7073 1687 7087 1700
rect 7116 1687 7123 2113
rect 7136 1807 7143 2093
rect 7156 1787 7163 2033
rect 7176 1667 7183 1953
rect 6896 1367 6903 1403
rect 6716 476 6743 483
rect 5796 216 5823 223
rect 5696 107 5703 143
rect 5796 27 5803 193
rect 5816 107 5823 216
rect 5456 -24 5463 13
rect 5716 -24 5723 13
rect 5916 -24 5923 233
rect 5996 -17 6003 143
rect 5976 -24 6003 -17
rect 6036 -24 6043 413
rect 6067 373 6073 387
rect 6096 327 6103 396
rect 6127 373 6133 387
rect 6116 144 6123 173
rect 6136 167 6143 373
rect 6196 327 6203 363
rect 6296 327 6303 376
rect 6316 67 6323 383
rect 6596 364 6603 433
rect 6636 307 6643 383
rect 6696 347 6703 383
rect 6736 347 6743 476
rect 6516 176 6523 253
rect 6556 176 6563 213
rect 6456 144 6463 173
rect 6636 67 6643 293
rect 6676 267 6683 313
rect 6756 287 6763 612
rect 6696 147 6703 273
rect 6776 267 6783 713
rect 6796 663 6803 713
rect 6856 703 6863 873
rect 6876 807 6883 1273
rect 6896 1184 6903 1253
rect 6916 1230 6923 1293
rect 6936 1267 6943 1403
rect 7016 1347 7023 1553
rect 6936 1240 7023 1243
rect 6936 1236 7027 1240
rect 6936 1216 6943 1236
rect 7013 1227 7027 1236
rect 6956 967 6963 1170
rect 6996 1107 7003 1183
rect 7036 1087 7043 1390
rect 7056 1147 7063 1633
rect 7076 1247 7083 1293
rect 7076 1167 7083 1212
rect 7096 1147 7103 1653
rect 7196 1627 7203 2223
rect 7216 1687 7223 1933
rect 7236 1927 7243 1953
rect 7256 1907 7263 2373
rect 7276 2007 7283 2913
rect 7296 2687 7303 2873
rect 7296 2224 7303 2473
rect 7316 2347 7323 3013
rect 7336 2723 7343 3236
rect 7356 2947 7363 3073
rect 7396 3027 7403 3073
rect 7436 2776 7443 3473
rect 7516 3047 7523 4473
rect 7536 3207 7543 5036
rect 7556 4407 7563 5009
rect 7576 4367 7583 4873
rect 7596 4727 7603 5043
rect 7716 4947 7723 6573
rect 7736 6547 7743 6633
rect 7756 6507 7763 6733
rect 7796 6600 7803 6603
rect 7793 6587 7807 6600
rect 7756 6187 7763 6383
rect 7816 6116 7823 6333
rect 7856 6147 7863 6553
rect 7916 6547 7923 6623
rect 7976 6587 7983 6623
rect 7976 6467 7983 6573
rect 7996 6487 8003 6553
rect 8016 6447 8023 6856
rect 8076 6847 8083 7073
rect 8096 6947 8103 7123
rect 8116 6827 8123 6953
rect 8136 6747 8143 7293
rect 8156 6887 8163 7613
rect 8176 7307 8183 7636
rect 8176 7107 8183 7133
rect 8216 7083 8223 7456
rect 8256 7087 8263 7173
rect 8276 7170 8283 7953
rect 8296 7407 8303 7993
rect 8416 7976 8423 8033
rect 8436 8003 8443 8113
rect 8436 7996 8463 8003
rect 8456 7976 8463 7996
rect 8336 7907 8343 7975
rect 8396 7940 8403 7943
rect 8393 7927 8407 7940
rect 8436 7847 8443 7943
rect 8496 7887 8503 8073
rect 8656 8047 8663 8073
rect 8736 8047 8743 8176
rect 8756 8107 8763 8133
rect 8356 7456 8363 7493
rect 8396 7456 8403 7833
rect 8596 7807 8603 7976
rect 8436 7643 8443 7733
rect 8476 7676 8483 7773
rect 8436 7636 8463 7643
rect 8336 7327 8343 7423
rect 8376 7420 8383 7423
rect 8373 7407 8387 7420
rect 8293 7160 8307 7173
rect 8296 7156 8303 7160
rect 8336 7156 8383 7163
rect 8316 7107 8323 7123
rect 8307 7096 8323 7107
rect 8307 7093 8320 7096
rect 8196 7076 8223 7083
rect 8176 6747 8183 6893
rect 8196 6787 8203 7076
rect 8216 6827 8223 7013
rect 8276 6936 8283 7073
rect 8376 6943 8383 7156
rect 8396 7087 8403 7313
rect 8416 6967 8423 7413
rect 8376 6936 8393 6943
rect 8256 6807 8263 6903
rect 8296 6900 8303 6903
rect 8293 6887 8307 6900
rect 8336 6670 8343 6733
rect 8036 6607 8043 6633
rect 8047 6423 8060 6427
rect 8047 6416 8063 6423
rect 8096 6416 8103 6493
rect 8047 6413 8060 6416
rect 7916 6387 7923 6413
rect 7796 6007 7803 6083
rect 7836 6080 7843 6083
rect 7833 6067 7847 6080
rect 7876 5896 7883 6233
rect 7916 5967 7923 6373
rect 7996 6367 8003 6413
rect 8136 6347 8143 6413
rect 8256 6367 8263 6473
rect 8296 6427 8303 6623
rect 8336 6507 8343 6573
rect 8376 6487 8383 6912
rect 8316 6430 8323 6453
rect 8396 6430 8403 6933
rect 8276 6387 8283 6416
rect 7816 5867 7823 5896
rect 7956 5864 7963 5933
rect 7856 5860 7863 5863
rect 7853 5847 7867 5860
rect 7736 5687 7743 5833
rect 7736 5427 7743 5673
rect 7736 5127 7743 5392
rect 7596 4407 7603 4713
rect 7616 4687 7623 4753
rect 7636 4663 7643 4856
rect 7756 4827 7763 5473
rect 7776 5263 7783 5713
rect 7796 5344 7803 5693
rect 7833 5600 7847 5613
rect 7836 5596 7843 5600
rect 7876 5596 7883 5633
rect 7896 5487 7903 5563
rect 7856 5376 7863 5413
rect 7896 5400 7943 5403
rect 7896 5396 7947 5400
rect 7896 5376 7903 5396
rect 7933 5390 7947 5396
rect 7776 5256 7803 5263
rect 7616 4656 7643 4663
rect 7616 4447 7623 4656
rect 7676 4556 7683 4633
rect 7636 4523 7643 4556
rect 7636 4516 7663 4523
rect 7656 4336 7663 4516
rect 7776 4523 7783 4993
rect 7796 4807 7803 5256
rect 7856 5076 7863 5293
rect 7896 5076 7903 5233
rect 7876 4907 7883 5043
rect 7956 5027 7963 5850
rect 7976 5787 7983 6193
rect 7996 6063 8003 6233
rect 8016 6083 8023 6213
rect 8073 6120 8087 6133
rect 8076 6116 8083 6120
rect 8016 6076 8043 6083
rect 7996 6056 8023 6063
rect 7996 5967 8003 6013
rect 7996 5564 8003 5953
rect 7996 5007 8003 5493
rect 7976 4856 7983 4933
rect 7956 4787 7963 4823
rect 7976 4556 7983 4793
rect 8016 4587 8023 6056
rect 7756 4516 7783 4523
rect 7716 4304 7723 4333
rect 7636 4300 7643 4303
rect 7633 4287 7647 4300
rect 7616 3996 7643 4003
rect 7556 3727 7563 3816
rect 7556 3447 7563 3516
rect 7576 3407 7583 3933
rect 7616 3807 7623 3893
rect 7636 3887 7643 3996
rect 7687 3953 7693 3967
rect 7596 3347 7603 3573
rect 7616 3567 7623 3653
rect 7636 3530 7643 3633
rect 7696 3484 7703 3553
rect 7616 3327 7623 3473
rect 7676 3264 7683 3453
rect 7456 2927 7463 3033
rect 7556 3027 7563 3213
rect 7496 2960 7503 2963
rect 7493 2947 7507 2960
rect 7356 2747 7363 2776
rect 7336 2716 7363 2723
rect 7336 2023 7343 2473
rect 7316 2016 7343 2023
rect 7316 1967 7323 2016
rect 7336 1970 7343 1993
rect 7356 1987 7363 2716
rect 7416 2707 7423 2743
rect 7376 2187 7383 2693
rect 7456 2667 7463 2743
rect 7436 2476 7443 2593
rect 7556 2507 7563 3013
rect 7576 2927 7583 3193
rect 7596 2887 7603 3113
rect 7513 2480 7527 2493
rect 7516 2476 7523 2480
rect 7436 2363 7443 2393
rect 7456 2387 7463 2443
rect 7496 2407 7503 2443
rect 7436 2356 7473 2363
rect 7436 2256 7443 2313
rect 7376 1956 7383 2093
rect 7156 1436 7163 1493
rect 7196 1436 7203 1513
rect 7116 1184 7123 1433
rect 7176 1327 7183 1403
rect 7056 1027 7063 1133
rect 7016 987 7023 1013
rect 6976 807 6983 883
rect 7036 847 7043 883
rect 6856 696 6883 703
rect 6936 697 6943 733
rect 6996 665 7003 793
rect 7076 687 7083 1053
rect 7136 929 7143 1233
rect 7156 1107 7163 1233
rect 7216 1216 7223 1403
rect 7256 1327 7263 1613
rect 7253 1220 7267 1233
rect 7276 1223 7283 1953
rect 7296 1767 7303 1953
rect 7336 1736 7343 1893
rect 7356 1887 7363 1923
rect 7296 1587 7303 1633
rect 7316 1507 7323 1703
rect 7336 1367 7343 1673
rect 7356 1607 7363 1703
rect 7396 1563 7403 1813
rect 7353 1547 7367 1553
rect 7376 1556 7403 1563
rect 7256 1216 7263 1220
rect 7276 1216 7303 1223
rect 7236 1180 7243 1183
rect 7233 1167 7247 1180
rect 7236 987 7243 1033
rect 7296 987 7303 1216
rect 7356 1067 7363 1533
rect 7376 1404 7383 1556
rect 7416 1547 7423 2173
rect 7456 2087 7463 2223
rect 7596 2187 7603 2833
rect 7616 2147 7623 2893
rect 7636 2567 7643 3253
rect 7716 3227 7723 3713
rect 7736 3647 7743 4393
rect 7756 3807 7763 4516
rect 7956 4487 7963 4523
rect 7996 4447 8003 4523
rect 7776 4004 7783 4113
rect 7856 4050 7863 4433
rect 7996 4407 8003 4433
rect 7876 4303 7883 4353
rect 7933 4340 7947 4353
rect 7936 4336 7943 4340
rect 7876 4296 7903 4303
rect 7916 4300 7923 4303
rect 7976 4300 7983 4303
rect 7816 3983 7823 3990
rect 7816 3976 7843 3983
rect 7756 3527 7763 3733
rect 7676 2964 7683 2993
rect 7696 2776 7703 3053
rect 7756 3047 7763 3513
rect 7776 3467 7783 3693
rect 7796 3647 7803 3953
rect 7796 3267 7803 3593
rect 7776 2903 7783 2963
rect 7776 2896 7803 2903
rect 7716 2627 7723 2743
rect 7756 2740 7763 2743
rect 7753 2727 7767 2740
rect 7796 2667 7803 2896
rect 7756 2476 7763 2513
rect 7736 2307 7743 2443
rect 7656 2223 7663 2293
rect 7656 2216 7683 2223
rect 7456 1887 7463 1956
rect 7676 1927 7683 2216
rect 7756 2087 7763 2223
rect 7596 1887 7603 1923
rect 7556 1736 7563 1813
rect 7596 1736 7603 1773
rect 7576 1607 7583 1703
rect 7396 1307 7403 1533
rect 7456 1436 7463 1593
rect 7496 1450 7503 1493
rect 7576 1404 7583 1593
rect 7616 1587 7623 1703
rect 7616 1450 7623 1573
rect 7476 1287 7483 1403
rect 7516 1216 7523 1253
rect 7576 1184 7583 1273
rect 7156 827 7163 913
rect 7256 883 7263 973
rect 7356 916 7363 1053
rect 7456 930 7463 1173
rect 7496 1107 7503 1183
rect 7396 879 7403 883
rect 7393 867 7407 879
rect 7216 696 7223 733
rect 7256 696 7263 733
rect 7476 696 7483 1093
rect 7516 696 7523 933
rect 6796 656 6823 663
rect 6796 227 6803 613
rect 6816 447 6823 656
rect 6836 567 6843 663
rect 6876 387 6883 513
rect 6996 447 7003 573
rect 7136 527 7143 696
rect 7236 647 7243 663
rect 7236 547 7243 633
rect 6936 396 6943 433
rect 6993 420 7007 433
rect 6996 416 7003 420
rect 6916 360 6923 363
rect 6913 347 6927 360
rect 7356 307 7363 383
rect 7416 380 7423 383
rect 7413 367 7427 380
rect 7456 367 7463 663
rect 6996 176 7003 253
rect 7356 187 7363 293
rect 7536 176 7543 396
rect 7556 287 7563 1133
rect 7596 1007 7603 1216
rect 7636 1147 7643 1633
rect 7676 1287 7683 1873
rect 7716 1750 7723 1993
rect 7716 1467 7723 1736
rect 7713 1440 7727 1453
rect 7716 1436 7723 1440
rect 7756 1436 7763 1956
rect 7776 1487 7783 2133
rect 7796 1967 7803 2293
rect 7796 1436 7803 1673
rect 7816 1467 7823 3793
rect 7836 3467 7843 3976
rect 7856 3607 7863 3973
rect 7876 3727 7883 3993
rect 7896 3987 7903 4296
rect 7913 4287 7927 4300
rect 7973 4287 7987 4300
rect 7976 3947 7983 4273
rect 7996 4004 8003 4033
rect 8016 3963 8023 4413
rect 8036 3987 8043 6076
rect 8056 5007 8063 6083
rect 8156 5896 8163 5933
rect 8196 5867 8203 6053
rect 8176 5687 8183 5713
rect 8176 5596 8183 5673
rect 8076 5167 8083 5596
rect 8116 5507 8123 5563
rect 8156 5507 8163 5563
rect 8216 5447 8223 5633
rect 8076 5047 8083 5113
rect 8096 5083 8103 5393
rect 8156 5307 8163 5343
rect 8216 5307 8223 5376
rect 8156 5147 8163 5272
rect 8096 5076 8123 5083
rect 8236 5047 8243 6153
rect 8256 5647 8263 6353
rect 8336 6347 8343 6383
rect 8416 6287 8423 6953
rect 8436 6267 8443 7213
rect 8456 6767 8463 7636
rect 8476 6927 8483 7613
rect 8516 7427 8523 7643
rect 8556 7207 8563 7673
rect 8576 7156 8583 7733
rect 8616 7627 8623 8033
rect 8636 7667 8643 8033
rect 8716 7976 8723 8013
rect 8753 7980 8767 7993
rect 8756 7976 8763 7980
rect 8696 7927 8703 7943
rect 8696 7747 8703 7913
rect 8796 7887 8803 8173
rect 8776 7676 8783 7873
rect 8676 7647 8683 7676
rect 8716 7627 8723 7643
rect 8647 7516 8673 7523
rect 8616 7367 8623 7423
rect 8536 6936 8543 6993
rect 8556 6987 8563 7123
rect 8596 7120 8603 7123
rect 8593 7107 8607 7120
rect 8656 7067 8663 7156
rect 8456 6670 8463 6713
rect 8456 6307 8463 6656
rect 8356 6116 8363 6173
rect 8376 6080 8383 6083
rect 8373 6067 8387 6080
rect 8396 5896 8403 5973
rect 8256 5547 8263 5596
rect 8256 5067 8263 5533
rect 8276 5407 8283 5613
rect 8276 5047 8283 5076
rect 8076 4827 8083 5012
rect 8056 4427 8063 4573
rect 8076 4487 8083 4510
rect 8056 4287 8063 4333
rect 8096 4307 8103 5033
rect 8156 4807 8163 4953
rect 8116 4103 8123 4733
rect 8176 4707 8183 5043
rect 8236 4856 8243 4993
rect 8196 4687 8203 4813
rect 8216 4787 8223 4823
rect 8256 4747 8263 4823
rect 8316 4570 8323 5653
rect 8336 5647 8343 5850
rect 8376 5727 8383 5863
rect 8476 5807 8483 6733
rect 8516 6703 8523 6903
rect 8556 6867 8563 6903
rect 8496 6696 8523 6703
rect 8496 6547 8503 6696
rect 8516 6447 8523 6673
rect 8536 6547 8543 6813
rect 8596 6707 8603 7033
rect 8696 6867 8703 6936
rect 8556 6667 8563 6693
rect 8716 6687 8723 7613
rect 8756 7447 8763 7643
rect 8816 7470 8823 8133
rect 8836 7227 8843 8153
rect 8856 7847 8863 8833
rect 8876 7944 8883 8773
rect 8896 8767 8903 8913
rect 8896 7627 8903 8732
rect 8916 7547 8923 8873
rect 8936 8807 8943 8893
rect 8953 8807 8967 8813
rect 9036 8716 9043 8933
rect 9056 8727 9063 9133
rect 9096 9107 9103 9273
rect 9216 9247 9223 10733
rect 9236 10727 9243 10750
rect 9556 10743 9563 11096
rect 9656 10947 9663 11270
rect 9693 11100 9707 11113
rect 9696 11096 9703 11100
rect 9736 11096 9743 11173
rect 9716 11060 9723 11063
rect 9713 11047 9727 11060
rect 9576 10767 9583 10813
rect 9716 10796 9723 10953
rect 9756 10796 9763 10833
rect 9816 10767 9823 11533
rect 9936 11507 9943 11823
rect 10013 11620 10027 11633
rect 10053 11620 10067 11633
rect 10016 11616 10023 11620
rect 10056 11616 10063 11620
rect 9996 11547 10003 11583
rect 9536 10736 9563 10743
rect 9236 9867 9243 10576
rect 9236 9727 9243 9853
rect 9256 9767 9263 10673
rect 9436 10276 9443 10633
rect 9456 10207 9463 10243
rect 9496 10207 9503 10576
rect 9536 10547 9543 10736
rect 9576 10576 9583 10613
rect 9656 10447 9663 10576
rect 9656 10276 9663 10433
rect 9676 10303 9683 10493
rect 9696 10347 9703 10750
rect 9676 10296 9703 10303
rect 9696 10276 9703 10296
rect 9276 9887 9283 10053
rect 9296 9756 9303 9973
rect 9336 9927 9343 9953
rect 9236 9427 9243 9533
rect 9256 9527 9263 9553
rect 9276 9367 9283 9710
rect 9316 9527 9323 9723
rect 9396 9536 9403 9653
rect 9427 9536 9433 9547
rect 9420 9533 9433 9536
rect 9276 9236 9283 9293
rect 9296 9107 9303 9203
rect 9336 9043 9343 9093
rect 9316 9036 9343 9043
rect 9316 9004 9323 9036
rect 9356 9023 9363 9353
rect 9336 9016 9363 9023
rect 9336 8996 9343 9016
rect 9396 9007 9403 9236
rect 9436 9003 9443 9453
rect 9416 8996 9443 9003
rect 9196 8747 9203 8853
rect 9076 8627 9083 8683
rect 9116 8667 9123 8713
rect 9176 8627 9183 8670
rect 9156 8616 9173 8623
rect 8936 8587 8943 8613
rect 9056 8496 9063 8593
rect 8936 7947 8943 8496
rect 8936 7487 8943 7933
rect 8956 7787 8963 8133
rect 8976 7987 8983 8196
rect 8996 8007 9003 8353
rect 9036 8327 9043 8463
rect 9056 8347 9063 8413
rect 9096 8196 9103 8253
rect 9156 8187 9163 8616
rect 9076 8127 9083 8163
rect 9116 8160 9123 8163
rect 9113 8147 9127 8160
rect 9147 8093 9153 8107
rect 9176 8063 9183 8493
rect 9196 8087 9203 8733
rect 9216 8647 9223 8873
rect 9236 8547 9243 8653
rect 9216 8127 9223 8196
rect 9236 8147 9243 8533
rect 9256 8464 9263 8753
rect 9293 8720 9307 8733
rect 9296 8716 9303 8720
rect 9316 8647 9323 8683
rect 9356 8680 9363 8683
rect 9353 8667 9367 8680
rect 9416 8287 9423 8996
rect 9436 8887 9443 8973
rect 9456 8287 9463 9913
rect 9536 9823 9543 10056
rect 9596 9907 9603 10023
rect 9636 10007 9643 10023
rect 9536 9816 9553 9823
rect 9556 9756 9563 9813
rect 9596 9807 9603 9893
rect 9636 9787 9643 9993
rect 9676 9947 9683 10243
rect 9593 9760 9607 9772
rect 9596 9756 9603 9760
rect 9636 9724 9643 9773
rect 9516 9716 9543 9723
rect 9576 9720 9583 9723
rect 9516 9627 9523 9716
rect 9573 9707 9587 9720
rect 9676 9667 9683 9933
rect 9696 9627 9703 10073
rect 9476 8767 9483 9513
rect 9496 8523 9503 9553
rect 9556 9307 9563 9613
rect 9607 9543 9620 9547
rect 9607 9536 9623 9543
rect 9607 9533 9620 9536
rect 9716 9503 9723 10233
rect 9676 9496 9723 9503
rect 9596 9250 9603 9393
rect 9516 8827 9523 9236
rect 9576 9107 9583 9203
rect 9636 9047 9643 9236
rect 9536 8907 9543 9013
rect 9556 8887 9563 9033
rect 9633 9020 9647 9033
rect 9636 9016 9643 9020
rect 9596 8827 9603 8983
rect 9656 8947 9663 8983
rect 9696 8947 9703 9496
rect 9716 9207 9723 9333
rect 9476 8516 9503 8523
rect 9476 8464 9483 8516
rect 9496 8307 9503 8493
rect 9376 8196 9383 8273
rect 9356 8107 9363 8163
rect 9247 8093 9253 8107
rect 9156 8056 9183 8063
rect 9053 7970 9067 7973
rect 9116 7963 9123 8033
rect 9156 7987 9163 8056
rect 9116 7956 9163 7963
rect 8976 7763 8983 7933
rect 8956 7756 8983 7763
rect 8956 7647 8963 7756
rect 8996 7676 9003 7793
rect 9036 7690 9043 7913
rect 9096 7643 9103 7833
rect 8956 7463 8963 7513
rect 8936 7456 8963 7463
rect 8876 7267 8883 7423
rect 8976 7207 8983 7473
rect 8996 7424 9003 7533
rect 8756 7124 8763 7193
rect 8856 7156 8863 7193
rect 8896 7156 8943 7163
rect 8816 6936 8823 7033
rect 8876 6767 8883 7123
rect 8936 7107 8943 7156
rect 8896 6904 8903 6993
rect 8556 6567 8563 6593
rect 8396 5707 8403 5733
rect 8336 4587 8343 5633
rect 8356 4887 8363 5633
rect 8413 5600 8427 5613
rect 8416 5596 8423 5600
rect 8376 5367 8383 5453
rect 8433 5380 8447 5393
rect 8436 5376 8443 5380
rect 8416 5307 8423 5343
rect 8476 5187 8483 5563
rect 8496 5044 8503 5333
rect 8136 4207 8143 4556
rect 8256 4487 8263 4523
rect 8196 4336 8203 4373
rect 8216 4300 8223 4303
rect 8107 4096 8123 4103
rect 8096 4036 8103 4093
rect 8056 3996 8073 4003
rect 8016 3956 8043 3963
rect 7936 3816 7943 3853
rect 8016 3787 8023 3913
rect 7916 3747 7923 3783
rect 7933 3520 7947 3533
rect 7936 3516 7943 3520
rect 7896 3296 7903 3453
rect 7976 3427 7983 3533
rect 7836 3087 7843 3250
rect 7836 2847 7843 3073
rect 7856 2790 7863 3073
rect 7836 2167 7843 2713
rect 7836 1907 7843 2153
rect 7856 2027 7863 2573
rect 7876 2567 7883 3213
rect 7896 2270 7903 3213
rect 7916 3067 7923 3133
rect 7956 3123 7963 3413
rect 7976 3247 7983 3296
rect 7996 3147 8003 3733
rect 8016 3207 8023 3633
rect 8036 3367 8043 3956
rect 8056 3830 8063 3996
rect 8056 3547 8063 3713
rect 7936 3116 7963 3123
rect 7936 3043 7943 3116
rect 7916 3036 7943 3043
rect 7916 2547 7923 3036
rect 7956 2783 7963 3033
rect 8036 2996 8043 3293
rect 8056 3127 8063 3533
rect 8076 3007 8083 3969
rect 8096 3264 8103 3753
rect 8116 3427 8123 3853
rect 8156 3767 8163 3993
rect 8176 3867 8183 4293
rect 8213 4287 8227 4300
rect 8196 3947 8203 4273
rect 8216 3847 8223 4036
rect 8236 4007 8243 4193
rect 8256 4050 8263 4093
rect 8256 3927 8263 4036
rect 8213 3820 8227 3833
rect 8216 3816 8223 3820
rect 8196 3587 8203 3783
rect 8136 3527 8143 3573
rect 8173 3520 8187 3533
rect 8216 3530 8223 3753
rect 8236 3667 8243 3693
rect 8256 3667 8263 3833
rect 8176 3516 8183 3520
rect 8196 3427 8203 3483
rect 8196 3347 8203 3373
rect 8156 3296 8163 3333
rect 8016 2943 8023 2963
rect 8016 2936 8043 2943
rect 7936 2776 7983 2783
rect 8013 2780 8027 2793
rect 8036 2787 8043 2936
rect 8016 2776 8023 2780
rect 7916 2407 7923 2533
rect 7936 2444 7943 2776
rect 8056 2487 8063 2873
rect 8076 2687 8083 2733
rect 7956 2267 7963 2473
rect 8036 2347 8043 2443
rect 7896 1987 7903 2256
rect 7893 1960 7907 1973
rect 7940 1963 7953 1967
rect 7896 1956 7903 1960
rect 7936 1956 7953 1963
rect 7940 1953 7953 1956
rect 7856 1916 7883 1923
rect 7856 1867 7863 1916
rect 7876 1736 7883 1893
rect 7916 1887 7923 1923
rect 7976 1887 7983 2073
rect 7856 1607 7863 1690
rect 7776 1400 7783 1403
rect 7773 1387 7787 1400
rect 7716 1167 7723 1293
rect 7736 1227 7743 1253
rect 7773 1220 7787 1233
rect 7776 1216 7783 1220
rect 7756 1180 7763 1183
rect 7753 1167 7767 1180
rect 7833 1167 7847 1173
rect 7576 664 7583 953
rect 7653 920 7667 933
rect 7656 916 7663 920
rect 7716 884 7723 933
rect 7776 904 7783 1133
rect 7676 827 7683 883
rect 7796 767 7803 1113
rect 7816 1063 7823 1153
rect 7816 1056 7843 1063
rect 7656 627 7663 733
rect 7733 700 7747 713
rect 7736 696 7743 700
rect 7816 667 7823 993
rect 7836 847 7843 1056
rect 7656 396 7663 613
rect 7836 267 7843 833
rect 7856 647 7863 1473
rect 7876 1167 7883 1633
rect 7896 1527 7903 1703
rect 7896 1387 7903 1513
rect 7916 1247 7923 1613
rect 7996 1547 8003 1973
rect 8016 1887 8023 1953
rect 7876 967 7883 1033
rect 7896 947 7903 1213
rect 7936 1187 7943 1373
rect 7976 1307 7983 1453
rect 8056 1436 8063 1690
rect 8076 1647 8083 2633
rect 8096 1967 8103 3250
rect 8116 1927 8123 3173
rect 8136 2127 8143 3263
rect 8176 3247 8183 3263
rect 8176 3207 8183 3233
rect 8156 2587 8163 3193
rect 8176 2523 8183 3113
rect 8156 2516 8183 2523
rect 8156 2047 8163 2516
rect 8176 2167 8183 2476
rect 8196 2187 8203 3253
rect 8216 3027 8223 3353
rect 8256 3267 8263 3516
rect 8276 3187 8283 4510
rect 8236 3067 8243 3113
rect 8296 3047 8303 4433
rect 8356 4407 8363 4852
rect 8376 4807 8383 5033
rect 8416 5023 8423 5043
rect 8416 5016 8443 5023
rect 8316 4007 8323 4336
rect 8396 4067 8403 4510
rect 8416 4267 8423 4993
rect 8436 4987 8443 5016
rect 8516 5007 8523 6253
rect 8536 5867 8543 6533
rect 8556 6427 8563 6553
rect 8596 6547 8603 6603
rect 8636 6567 8643 6623
rect 8696 6620 8703 6623
rect 8693 6607 8707 6620
rect 8573 6420 8587 6433
rect 8576 6416 8583 6420
rect 8656 6416 8663 6553
rect 8696 6507 8703 6593
rect 8636 6380 8643 6383
rect 8633 6367 8647 6380
rect 8536 5567 8543 5613
rect 8536 5344 8543 5393
rect 8556 5207 8563 6273
rect 8576 6027 8583 6070
rect 8576 5607 8583 5913
rect 8536 5027 8543 5133
rect 8456 4787 8463 4873
rect 8516 4856 8523 4933
rect 8556 4870 8563 5153
rect 8576 5107 8583 5393
rect 8576 4907 8583 5093
rect 8596 5087 8603 6083
rect 8636 6080 8643 6083
rect 8633 6067 8647 6080
rect 8636 6007 8643 6053
rect 8693 5900 8707 5913
rect 8696 5896 8703 5900
rect 8616 5527 8623 5896
rect 8693 5827 8707 5833
rect 8716 5787 8723 5833
rect 8636 5427 8643 5753
rect 8656 5487 8663 5733
rect 8736 5667 8743 6753
rect 9016 6747 9023 7110
rect 9036 6947 9043 7533
rect 9056 7170 9063 7643
rect 9076 7636 9103 7643
rect 9076 7087 9083 7636
rect 9096 7347 9103 7573
rect 9116 7567 9123 7873
rect 9116 7247 9123 7553
rect 9136 7463 9143 7673
rect 9156 7507 9163 7956
rect 9436 7956 9443 8233
rect 9496 8164 9503 8272
rect 9516 7944 9523 8553
rect 9576 8496 9583 8593
rect 9556 8460 9563 8463
rect 9596 8460 9603 8463
rect 9553 8447 9567 8460
rect 9593 8447 9607 8460
rect 9636 8447 9643 8813
rect 9556 8367 9563 8433
rect 9176 7547 9183 7793
rect 9296 7690 9303 7733
rect 9476 7727 9483 7923
rect 9516 7687 9523 7930
rect 9536 7867 9543 8193
rect 9556 7847 9563 8233
rect 9616 8196 9623 8273
rect 9656 8247 9663 8873
rect 9676 8287 9683 8493
rect 9596 8160 9603 8163
rect 9593 8147 9607 8160
rect 9576 7807 9583 8013
rect 9596 7990 9603 8133
rect 9636 8127 9643 8163
rect 9716 8027 9723 9073
rect 9736 8447 9743 10173
rect 9756 9707 9763 9833
rect 9756 9504 9763 9573
rect 9776 9467 9783 10753
rect 9856 10576 9863 11353
rect 9996 11096 10003 11433
rect 10036 11330 10043 11570
rect 9876 10727 9883 10913
rect 9916 10687 9923 11093
rect 10056 11064 10063 11113
rect 10076 11067 10083 11096
rect 9976 10803 9983 11063
rect 9956 10796 9983 10803
rect 10016 10796 10023 10873
rect 9836 10527 9843 10543
rect 9836 10247 9843 10513
rect 9876 10267 9883 10543
rect 9956 10387 9963 10796
rect 10016 10507 10023 10613
rect 10096 10607 10103 11313
rect 10116 11284 10123 11313
rect 10136 10867 10143 12073
rect 10356 11967 10363 12103
rect 10196 11856 10233 11863
rect 10196 11843 10203 11856
rect 10176 11840 10203 11843
rect 10173 11836 10203 11840
rect 10516 11836 10523 12053
rect 10547 11853 10553 11867
rect 10173 11830 10187 11836
rect 10256 11800 10263 11803
rect 10253 11787 10267 11800
rect 10156 11267 10163 11493
rect 10216 11347 10223 11773
rect 10253 11620 10267 11633
rect 10256 11616 10263 11620
rect 10296 11616 10303 11713
rect 10356 11627 10363 11753
rect 10356 11584 10363 11613
rect 9960 10303 9973 10307
rect 9956 10293 9973 10303
rect 9956 10276 9963 10293
rect 10016 10244 10023 10493
rect 9976 10236 10003 10243
rect 9936 10107 9943 10173
rect 9893 10060 9907 10073
rect 9896 10056 9903 10060
rect 9936 10056 9943 10093
rect 9996 10087 10003 10236
rect 9836 10024 9843 10053
rect 9816 9807 9823 9913
rect 9816 9756 9823 9793
rect 9956 9707 9963 9853
rect 9856 9547 9863 9613
rect 9856 9504 9863 9533
rect 9836 9387 9843 9453
rect 9756 8887 9763 9313
rect 9796 9236 9803 9313
rect 9836 9236 9843 9373
rect 9756 8684 9763 8873
rect 9816 8867 9823 9203
rect 9936 9107 9943 9453
rect 9916 9047 9923 9073
rect 9956 8984 9963 9373
rect 9836 8716 9843 8933
rect 9876 8907 9883 8983
rect 9880 8723 9893 8727
rect 9876 8716 9893 8723
rect 9880 8713 9893 8716
rect 9776 8507 9783 8713
rect 9936 8687 9943 8793
rect 9856 8627 9863 8683
rect 9956 8647 9963 8970
rect 9976 8567 9983 10056
rect 9996 9467 10003 10073
rect 10036 9727 10043 10253
rect 9787 8496 9803 8503
rect 9836 8496 9883 8503
rect 9876 8367 9883 8496
rect 9736 7976 9743 8273
rect 9776 8127 9783 8213
rect 9796 7956 9803 8193
rect 9836 8007 9843 8293
rect 9996 8247 10003 9233
rect 10016 9207 10023 9673
rect 10016 8984 10023 9193
rect 10016 8467 10023 8713
rect 10036 8527 10043 9692
rect 10056 9247 10063 10593
rect 10176 10544 10183 11313
rect 10336 11284 10343 11413
rect 10256 11280 10263 11283
rect 10253 11267 10267 11280
rect 10296 10796 10303 10873
rect 10256 10544 10263 10573
rect 10136 10307 10143 10543
rect 10076 10024 10083 10293
rect 10096 9867 10103 10293
rect 10216 10276 10223 10393
rect 10156 10056 10163 10230
rect 10216 10027 10223 10193
rect 10236 10187 10243 10243
rect 10276 10187 10283 10713
rect 10376 10576 10383 11790
rect 10496 11727 10503 11803
rect 10396 11587 10403 11633
rect 10576 11616 10583 11893
rect 10596 11707 10603 12136
rect 10756 12107 10763 12136
rect 10636 12100 10643 12103
rect 10633 12087 10647 12100
rect 10676 12027 10683 12103
rect 10716 12067 10723 12103
rect 10916 12103 10923 12136
rect 10916 12096 10943 12103
rect 10736 11836 10743 11873
rect 10767 11863 10780 11867
rect 10767 11853 10783 11863
rect 10776 11836 10783 11853
rect 10516 11327 10523 11616
rect 10556 11580 10563 11583
rect 10553 11567 10567 11580
rect 10596 11407 10603 11570
rect 10696 11547 10703 11836
rect 10856 11804 10863 11873
rect 10756 11707 10763 11803
rect 10396 10727 10403 11096
rect 10416 10887 10423 11316
rect 10556 11316 10563 11353
rect 10636 11307 10643 11393
rect 10476 11096 10483 11270
rect 10576 11247 10583 11283
rect 10456 11027 10463 11063
rect 10536 10796 10543 10833
rect 10436 10627 10443 10796
rect 10136 10020 10143 10023
rect 10133 10007 10147 10020
rect 10176 9927 10183 10023
rect 10196 9927 10203 9953
rect 10236 9887 10243 10173
rect 10076 9767 10083 9793
rect 10236 9767 10243 9873
rect 10076 9724 10083 9753
rect 10073 9567 10087 9573
rect 10076 9504 10083 9553
rect 10076 9236 10083 9273
rect 10096 9247 10103 9713
rect 10156 9720 10163 9723
rect 10153 9707 10167 9720
rect 10116 9467 10123 9633
rect 10176 9570 10183 9713
rect 10296 9687 10303 9756
rect 10196 9327 10203 9490
rect 10216 9347 10223 9413
rect 10136 9236 10143 9273
rect 10256 9250 10263 9433
rect 10096 9047 10103 9193
rect 10116 9147 10123 9203
rect 10096 8947 10103 9033
rect 10156 9030 10163 9133
rect 10176 8947 10183 8983
rect 10156 8716 10163 8773
rect 10276 8647 10283 9613
rect 10296 9204 10303 9533
rect 10316 8723 10323 10576
rect 10456 10544 10463 10753
rect 10576 10707 10583 10763
rect 10636 10576 10643 10873
rect 10676 10764 10683 11293
rect 10696 11287 10703 11533
rect 10836 11447 10843 11583
rect 10896 11316 10903 11353
rect 10716 11096 10723 11153
rect 10756 11096 10763 11316
rect 10827 11283 10840 11287
rect 10827 11276 10843 11283
rect 10827 11273 10840 11276
rect 10876 11247 10883 11283
rect 10816 11064 10823 11213
rect 10736 10847 10743 11063
rect 10776 10967 10783 11050
rect 10836 10867 10843 11173
rect 10816 10796 10823 10833
rect 10356 10244 10363 10333
rect 10476 10276 10483 10453
rect 10356 9807 10363 10230
rect 10496 10187 10503 10243
rect 10436 10056 10443 10093
rect 10396 9987 10403 10023
rect 10396 9756 10403 9793
rect 10376 9549 10383 9723
rect 10456 9536 10463 9833
rect 10373 9240 10387 9253
rect 10376 9236 10383 9240
rect 10436 9204 10443 9503
rect 10496 9387 10503 9793
rect 10516 9507 10523 9973
rect 10536 9487 10543 10533
rect 10556 10087 10563 10153
rect 10436 9016 10443 9190
rect 10516 9067 10523 9253
rect 10316 8716 10333 8723
rect 10416 8723 10423 8983
rect 10556 8767 10563 9753
rect 10576 8907 10583 10393
rect 10596 9247 10603 10276
rect 10616 9847 10623 10543
rect 10656 10407 10663 10530
rect 10716 10367 10723 10796
rect 10836 10760 10843 10763
rect 10833 10747 10847 10760
rect 10896 10727 10903 10796
rect 10936 10747 10943 12096
rect 10976 12047 10983 12103
rect 11013 12087 11027 12093
rect 11036 12087 11043 12136
rect 11056 11836 11063 12136
rect 11087 12093 11093 12107
rect 11216 11867 11223 12103
rect 11376 12087 11383 12136
rect 11376 11863 11383 12073
rect 11396 12067 11403 12173
rect 11476 12136 11483 12173
rect 11993 12140 12007 12153
rect 11996 12136 12003 12140
rect 11456 12067 11463 12103
rect 11656 11907 11663 12136
rect 11776 12103 11783 12136
rect 11756 12096 11783 12103
rect 11376 11856 11403 11863
rect 11116 11803 11123 11836
rect 11016 11796 11043 11803
rect 10956 11630 10963 11733
rect 10956 11330 10963 11616
rect 10956 11147 10963 11316
rect 11016 11287 11023 11796
rect 11076 11767 11083 11803
rect 11096 11796 11123 11803
rect 11096 11616 11103 11796
rect 11036 11243 11043 11533
rect 11076 11527 11083 11583
rect 11056 11516 11073 11523
rect 11056 11267 11063 11516
rect 11116 11367 11123 11583
rect 11036 11236 11063 11243
rect 11056 11096 11063 11236
rect 10956 11027 10963 11096
rect 10696 10290 10703 10333
rect 10716 10127 10723 10243
rect 10776 10167 10783 10276
rect 10796 10067 10803 10353
rect 10836 10127 10843 10673
rect 10896 10576 10903 10613
rect 10856 10107 10863 10413
rect 10876 10387 10883 10530
rect 10927 10493 10933 10507
rect 10956 10307 10963 11013
rect 10996 10687 11003 11063
rect 11036 10987 11043 11063
rect 10976 10544 10983 10573
rect 10953 10280 10967 10293
rect 10956 10276 10963 10280
rect 10976 10240 10983 10243
rect 10973 10227 10987 10240
rect 10716 9927 10723 10023
rect 10696 9720 10703 9723
rect 10693 9707 10707 9720
rect 10756 9707 10763 9913
rect 10776 9727 10783 9756
rect 10696 9647 10703 9693
rect 10656 9536 10663 9613
rect 10756 9503 10763 9653
rect 10716 9500 10723 9503
rect 10616 9236 10623 9353
rect 10676 9287 10683 9490
rect 10713 9487 10727 9500
rect 10736 9496 10763 9503
rect 10636 9147 10643 9203
rect 10696 9016 10703 9313
rect 10676 8827 10683 8983
rect 10416 8716 10443 8723
rect 10656 8716 10663 8753
rect 10056 8407 10063 8463
rect 10096 8460 10103 8463
rect 10093 8447 10107 8460
rect 10136 8387 10143 8493
rect 10156 8447 10163 8633
rect 10336 8523 10343 8713
rect 10396 8647 10403 8683
rect 10336 8516 10363 8523
rect 10313 8500 10327 8513
rect 10316 8496 10323 8500
rect 10356 8496 10363 8516
rect 10336 8447 10343 8463
rect 10336 8436 10353 8447
rect 10340 8433 10353 8436
rect 9893 8200 9907 8213
rect 9896 8196 9903 8200
rect 9936 8196 9943 8233
rect 9856 7967 9863 8170
rect 9847 7956 9863 7967
rect 9876 7964 9883 8053
rect 9847 7953 9860 7956
rect 9716 7807 9723 7930
rect 9596 7676 9603 7753
rect 9376 7643 9383 7673
rect 9336 7636 9383 7643
rect 9536 7640 9543 7643
rect 9533 7627 9547 7640
rect 9136 7456 9163 7463
rect 9276 7436 9283 7553
rect 9336 7436 9343 7493
rect 9356 7444 9363 7593
rect 9156 7120 9163 7123
rect 9153 7107 9167 7120
rect 9056 6936 9063 6973
rect 9136 6903 9143 7073
rect 9056 6656 9063 6713
rect 9076 6663 9083 6893
rect 9096 6867 9103 6903
rect 9116 6896 9143 6903
rect 9076 6656 9103 6663
rect 8916 6416 8923 6453
rect 8756 5747 8763 6353
rect 8836 6147 8843 6413
rect 8896 6380 8903 6383
rect 8856 6167 8863 6373
rect 8893 6367 8907 6380
rect 8976 6247 8983 6473
rect 9016 6307 9023 6623
rect 9096 6607 9103 6656
rect 9036 6347 9043 6416
rect 8916 6116 8923 6153
rect 8796 5987 8803 6116
rect 8693 5627 8707 5633
rect 8693 5600 8707 5613
rect 8696 5596 8703 5600
rect 8676 5267 8683 5343
rect 8716 5167 8723 5513
rect 8736 5247 8743 5533
rect 8756 5347 8763 5473
rect 8756 5207 8763 5233
rect 8653 5080 8667 5093
rect 8656 5076 8663 5080
rect 8496 4747 8503 4823
rect 8436 4487 8443 4613
rect 8496 4587 8503 4613
rect 8516 4587 8523 4773
rect 8536 4767 8543 4823
rect 8496 4556 8503 4573
rect 8516 4520 8523 4523
rect 8513 4507 8527 4520
rect 8476 4336 8483 4373
rect 8516 4336 8523 4393
rect 8416 4036 8423 4193
rect 8436 4127 8443 4273
rect 8456 4147 8463 4303
rect 8556 4303 8563 4793
rect 8536 4296 8563 4303
rect 8336 3996 8363 4003
rect 8336 3887 8343 3996
rect 8316 3687 8323 3853
rect 8336 3787 8343 3873
rect 8336 3507 8343 3773
rect 8316 3267 8323 3293
rect 8356 3227 8363 3973
rect 8396 3823 8403 4003
rect 8456 3947 8463 4053
rect 8376 3816 8403 3823
rect 8456 3816 8463 3853
rect 8476 3847 8483 4253
rect 8376 3767 8383 3816
rect 8516 3787 8523 4053
rect 8536 3987 8543 4296
rect 8576 4163 8583 4553
rect 8556 4156 8583 4163
rect 8556 3963 8563 4156
rect 8596 4143 8603 4933
rect 8616 4787 8623 5076
rect 8756 5047 8763 5172
rect 8676 4987 8683 5043
rect 8776 4987 8783 5793
rect 8816 5767 8823 6053
rect 8896 6047 8903 6083
rect 8933 5900 8947 5913
rect 8936 5896 8943 5900
rect 8796 5507 8803 5596
rect 8816 5487 8823 5753
rect 8856 5567 8863 5896
rect 8876 5503 8883 5813
rect 8896 5687 8903 5833
rect 8896 5547 8903 5633
rect 8856 5496 8883 5503
rect 8816 5327 8823 5373
rect 8796 4987 8803 5193
rect 8816 5027 8823 5253
rect 8836 4987 8843 5413
rect 8856 5344 8863 5496
rect 8916 5407 8923 5863
rect 9056 5827 9063 6533
rect 9116 6487 9123 6896
rect 9133 6727 9147 6733
rect 9156 6547 9163 6936
rect 9176 6587 9183 7073
rect 9216 6827 9223 7423
rect 9236 7170 9243 7413
rect 9256 6907 9263 7133
rect 9076 5967 9083 6453
rect 9196 6416 9203 6733
rect 9236 6630 9243 6773
rect 9253 6727 9267 6733
rect 9136 6367 9143 6383
rect 9176 6380 9183 6383
rect 9173 6367 9187 6380
rect 9136 6307 9143 6353
rect 9096 6083 9103 6133
rect 9156 6116 9163 6173
rect 9096 6076 9143 6083
rect 9176 6080 9183 6083
rect 9173 6067 9187 6080
rect 9116 5864 9123 5913
rect 9136 5863 9143 6053
rect 9216 6047 9223 6116
rect 9256 6027 9263 6673
rect 9276 6647 9283 7293
rect 9356 7144 9363 7393
rect 9376 7287 9383 7613
rect 9576 7547 9583 7643
rect 9396 7407 9403 7473
rect 9656 7436 9663 7753
rect 9676 7447 9683 7673
rect 9696 7367 9703 7403
rect 9416 7156 9423 7273
rect 9736 7247 9743 7533
rect 9756 7367 9763 7713
rect 9776 7487 9783 7913
rect 9816 7507 9823 7643
rect 9796 7407 9803 7433
rect 9816 7387 9823 7493
rect 9836 7307 9843 7613
rect 9856 7467 9863 7513
rect 9576 7150 9583 7233
rect 9876 7227 9883 7833
rect 9896 7627 9903 8133
rect 9916 8067 9923 8163
rect 9956 8107 9963 8163
rect 9996 8147 10003 8183
rect 10096 8107 10103 8373
rect 10436 8247 10443 8716
rect 10476 8547 10483 8593
rect 10456 8327 10463 8513
rect 10496 8407 10503 8716
rect 10736 8684 10743 9496
rect 10756 8827 10763 9233
rect 10096 8067 10103 8093
rect 10216 7907 10223 7923
rect 10216 7727 10223 7893
rect 10256 7867 10263 7953
rect 10056 7607 10063 7643
rect 9916 7456 9923 7573
rect 9956 7456 9963 7593
rect 10056 7436 10063 7493
rect 10096 7444 10103 7643
rect 10116 7436 10123 7513
rect 10156 7424 10163 7673
rect 10296 7647 10303 8073
rect 10316 7687 10323 8033
rect 10376 7907 10383 8183
rect 10396 7907 10403 8173
rect 10476 8087 10483 8353
rect 10433 7980 10447 7993
rect 10480 7983 10493 7987
rect 10436 7976 10443 7980
rect 10476 7976 10493 7983
rect 10480 7973 10493 7976
rect 10516 7967 10523 8670
rect 10636 8567 10643 8683
rect 10536 8167 10543 8553
rect 10656 8496 10663 8593
rect 10596 8460 10603 8463
rect 10636 8460 10643 8463
rect 10593 8447 10607 8460
rect 10633 8447 10647 8460
rect 10456 7847 10463 7943
rect 10336 7676 10343 7733
rect 10373 7680 10387 7693
rect 10376 7676 10383 7680
rect 10436 7436 10443 7793
rect 10536 7767 10543 8013
rect 10496 7443 10503 7673
rect 10516 7607 10523 7733
rect 10516 7563 10523 7593
rect 10516 7556 10543 7563
rect 10496 7436 10523 7443
rect 9936 7420 9943 7423
rect 9933 7407 9947 7420
rect 9436 7087 9443 7123
rect 9476 7087 9483 7143
rect 9936 7147 9943 7233
rect 9496 7067 9503 7093
rect 9536 7067 9543 7130
rect 9956 7047 9963 7176
rect 9976 7107 9983 7410
rect 9376 6767 9383 6973
rect 9316 6636 9323 6673
rect 9376 6627 9383 6673
rect 9296 6547 9303 6603
rect 9416 6547 9423 6853
rect 9436 6467 9443 6993
rect 9476 6907 9483 7013
rect 9476 6467 9483 6713
rect 9496 6527 9503 6636
rect 9516 6467 9523 7013
rect 9616 6976 9623 7013
rect 9656 6943 9663 6944
rect 9676 6943 9683 7013
rect 9656 6936 9683 6943
rect 9796 6907 9803 6936
rect 9816 6727 9823 7033
rect 9913 6940 9927 6953
rect 9916 6936 9923 6940
rect 9856 6867 9863 6903
rect 9896 6807 9903 6903
rect 9556 6636 9563 6673
rect 9656 6656 9663 6713
rect 9556 6447 9563 6573
rect 9596 6447 9603 6603
rect 9956 6587 9963 6653
rect 9976 6624 9983 7053
rect 9996 6904 10003 7213
rect 10016 7027 10023 7373
rect 10036 6667 10043 7273
rect 10156 7247 10163 7410
rect 10516 7407 10523 7436
rect 10476 7367 10483 7403
rect 10116 7120 10123 7123
rect 10113 7107 10127 7120
rect 10216 6967 10223 7033
rect 10216 6936 10223 6953
rect 10096 6707 10103 6753
rect 10076 6616 10103 6623
rect 9493 6420 9507 6433
rect 9496 6416 9503 6420
rect 9433 6367 9447 6370
rect 9236 5896 9243 5933
rect 9136 5856 9163 5863
rect 8933 5607 8947 5613
rect 8973 5600 8987 5613
rect 8976 5596 8983 5600
rect 9156 5583 9163 5856
rect 9216 5807 9223 5863
rect 9276 5827 9283 6353
rect 9476 6207 9483 6383
rect 9416 5947 9423 6083
rect 9496 5896 9503 6153
rect 9536 5896 9543 6033
rect 9576 5910 9583 6353
rect 9616 5864 9623 6453
rect 9476 5616 9483 5733
rect 9516 5607 9523 5713
rect 8936 5427 8943 5553
rect 8956 5507 8963 5563
rect 8996 5560 9003 5563
rect 8993 5547 9007 5560
rect 9056 5547 9063 5583
rect 8936 5376 8943 5413
rect 8636 4427 8643 4473
rect 8616 4347 8623 4393
rect 8636 4287 8643 4373
rect 8656 4267 8663 4573
rect 8587 4136 8603 4143
rect 8536 3956 8563 3963
rect 8480 3783 8493 3787
rect 8436 3780 8443 3783
rect 8433 3767 8447 3780
rect 8476 3776 8493 3783
rect 8480 3773 8493 3776
rect 8416 3587 8423 3633
rect 8536 3587 8543 3956
rect 8556 3727 8563 3816
rect 8456 3516 8463 3573
rect 8500 3543 8513 3547
rect 8496 3533 8513 3543
rect 8496 3516 8503 3533
rect 8556 3484 8563 3513
rect 8476 3387 8483 3483
rect 8416 3296 8423 3373
rect 8496 3267 8503 3296
rect 8576 3247 8583 4133
rect 8596 3967 8603 4112
rect 8616 4047 8623 4153
rect 8636 4067 8643 4133
rect 8656 4036 8663 4173
rect 8676 4167 8683 4673
rect 8696 4387 8703 4856
rect 8716 4336 8723 4613
rect 8736 4567 8743 4973
rect 8816 4907 8823 4953
rect 8856 4947 8863 5330
rect 8793 4860 8807 4873
rect 8796 4856 8803 4860
rect 8816 4803 8823 4823
rect 8796 4800 8823 4803
rect 8793 4796 8823 4800
rect 8853 4807 8867 4810
rect 8793 4787 8807 4796
rect 8876 4787 8883 5333
rect 8956 5340 8963 5343
rect 8953 5327 8967 5340
rect 8996 5167 9003 5353
rect 9016 5147 9023 5253
rect 8756 4556 8763 4773
rect 8816 4387 8823 4733
rect 8753 4340 8767 4353
rect 8756 4336 8763 4340
rect 8696 4123 8703 4290
rect 8736 4283 8743 4303
rect 8716 4276 8743 4283
rect 8716 4147 8723 4276
rect 8696 4120 8723 4123
rect 8696 4116 8727 4120
rect 8713 4107 8727 4116
rect 8696 4036 8703 4073
rect 8596 3787 8603 3873
rect 8636 3787 8643 4003
rect 8596 3387 8603 3533
rect 8656 3307 8663 3833
rect 8716 3830 8723 3953
rect 8736 3887 8743 4253
rect 8756 3847 8763 4273
rect 8796 4247 8803 4273
rect 8836 4187 8843 4773
rect 8896 4747 8903 5053
rect 8916 4947 8923 5033
rect 8916 4807 8923 4933
rect 8936 4870 8943 5043
rect 9036 5007 9043 5076
rect 9096 5047 9103 5376
rect 9116 5027 9123 5583
rect 9136 5576 9163 5583
rect 9136 5343 9143 5576
rect 9176 5376 9183 5413
rect 9136 5336 9163 5343
rect 9096 4907 9103 4973
rect 8936 4827 8943 4856
rect 9113 4860 9127 4873
rect 9116 4856 9123 4860
rect 8976 4827 8983 4853
rect 9056 4787 9063 4810
rect 8856 4667 8863 4713
rect 8876 4647 8883 4713
rect 8796 3967 8803 4153
rect 8753 3820 8767 3833
rect 8756 3816 8763 3820
rect 8736 3747 8743 3783
rect 8256 2867 8263 2996
rect 8316 2927 8323 2963
rect 8253 2780 8267 2793
rect 8256 2776 8263 2780
rect 8236 2707 8243 2743
rect 8293 2480 8307 2493
rect 8296 2476 8303 2480
rect 8276 2367 8283 2443
rect 8356 2367 8363 2893
rect 8276 2256 8283 2293
rect 8216 2207 8223 2256
rect 8376 2227 8383 3033
rect 8396 2407 8403 2776
rect 8416 2744 8423 3033
rect 8436 2787 8443 2853
rect 8436 2707 8443 2773
rect 8320 2223 8333 2227
rect 8256 2220 8263 2223
rect 8253 2207 8267 2220
rect 8316 2216 8333 2223
rect 8320 2213 8333 2216
rect 8416 2187 8423 2573
rect 8456 2507 8463 2853
rect 8436 2387 8443 2493
rect 8436 2247 8443 2352
rect 8196 1956 8203 2113
rect 8096 1647 8103 1873
rect 8156 1736 8163 1873
rect 8196 1787 8203 1813
rect 8196 1736 8203 1773
rect 8236 1707 8243 1773
rect 8136 1487 8143 1703
rect 8176 1607 8183 1703
rect 8156 1230 8163 1353
rect 8216 1347 8223 1553
rect 8256 1527 8263 2033
rect 8276 1687 8283 2153
rect 8296 1787 8303 2173
rect 8456 2107 8463 2493
rect 8476 2443 8483 2996
rect 8516 2967 8523 3233
rect 8596 3047 8603 3293
rect 8667 3263 8680 3267
rect 8667 3256 8683 3263
rect 8667 3253 8680 3256
rect 8616 3023 8623 3193
rect 8607 3016 8623 3023
rect 8593 3000 8607 3012
rect 8596 2996 8603 3000
rect 8636 2843 8643 2996
rect 8636 2836 8653 2843
rect 8576 2776 8583 2833
rect 8516 2687 8523 2743
rect 8536 2476 8543 2533
rect 8476 2436 8503 2443
rect 8456 2047 8463 2093
rect 8316 1607 8323 1956
rect 8496 1927 8503 2436
rect 8516 2407 8523 2443
rect 8556 2347 8563 2443
rect 8576 2256 8583 2413
rect 8596 2270 8603 2353
rect 8556 2187 8563 2223
rect 8616 2127 8623 2730
rect 8436 1847 8443 1923
rect 8436 1736 8443 1773
rect 8316 1436 8323 1593
rect 8356 1404 8363 1573
rect 7956 1087 7963 1213
rect 7976 1067 7983 1113
rect 8056 1047 8063 1170
rect 8216 1047 8223 1073
rect 8336 1047 8343 1183
rect 8376 1087 8383 1736
rect 8396 1407 8403 1673
rect 8416 1567 8423 1690
rect 8456 1607 8463 1703
rect 7916 916 7923 1013
rect 8416 967 8423 1033
rect 8096 927 8103 953
rect 8416 936 8423 953
rect 7876 707 7883 733
rect 7856 364 7863 633
rect 7896 627 7903 883
rect 7936 807 7943 883
rect 7936 547 7943 793
rect 7956 787 7963 853
rect 8056 847 8063 903
rect 8456 887 8463 1170
rect 7996 696 8003 753
rect 8296 696 8303 733
rect 7956 396 7963 693
rect 8016 567 8023 663
rect 8056 660 8063 663
rect 8053 647 8067 660
rect 8316 507 8323 663
rect 8356 627 8363 663
rect 8416 627 8423 873
rect 8436 587 8443 813
rect 8456 667 8463 773
rect 8436 430 8443 573
rect 8476 567 8483 1513
rect 8516 1487 8523 1736
rect 8516 1187 8523 1473
rect 8536 1447 8543 1473
rect 8576 1436 8583 1873
rect 8596 1507 8603 1956
rect 8636 1687 8643 2293
rect 8656 2227 8663 2833
rect 8676 2067 8683 2313
rect 8696 2147 8703 3033
rect 8716 2647 8723 3173
rect 8736 2687 8743 3013
rect 8776 2907 8783 3470
rect 8796 3447 8803 3816
rect 8796 3264 8803 3293
rect 8816 3047 8823 4093
rect 8836 3707 8843 3893
rect 8856 3067 8863 4510
rect 8936 4427 8943 4753
rect 9007 4713 9013 4727
rect 8956 4567 8963 4693
rect 9036 4556 9043 4753
rect 9096 4647 9103 4823
rect 9076 4487 9083 4556
rect 9096 4527 9103 4573
rect 8876 3747 8883 4413
rect 9076 4367 9083 4473
rect 8956 4247 8963 4353
rect 8996 4267 9003 4303
rect 9016 4167 9023 4213
rect 8956 4107 8963 4133
rect 8987 4073 8993 4087
rect 8973 4040 8987 4052
rect 9036 4047 9043 4193
rect 9056 4127 9063 4293
rect 8976 4036 8983 4040
rect 9056 4023 9063 4113
rect 9076 4047 9083 4353
rect 9096 4187 9103 4313
rect 9093 4087 9107 4093
rect 9056 4016 9083 4023
rect 8916 3883 8923 4003
rect 8956 4000 8963 4003
rect 8953 3987 8967 4000
rect 8916 3876 8943 3883
rect 8936 3847 8943 3876
rect 8876 3167 8883 3333
rect 8896 3187 8903 3673
rect 8876 2996 8883 3153
rect 8916 3067 8923 3816
rect 8936 3527 8943 3833
rect 9016 3830 9023 4013
rect 8956 3747 8963 3773
rect 8996 3747 9003 3783
rect 8996 3567 9003 3593
rect 8996 3516 9003 3553
rect 8936 3484 8943 3513
rect 9016 3447 9023 3483
rect 8936 3307 8943 3353
rect 8993 3300 9007 3313
rect 8996 3296 9003 3300
rect 8816 2823 8823 2963
rect 8856 2927 8863 2963
rect 8796 2816 8823 2823
rect 8796 2776 8803 2816
rect 8833 2780 8847 2793
rect 8913 2787 8927 2793
rect 8836 2776 8843 2780
rect 8736 2307 8743 2533
rect 8756 2047 8763 2553
rect 8776 2443 8783 2653
rect 8816 2503 8823 2743
rect 8816 2496 8843 2503
rect 8836 2476 8843 2496
rect 8873 2480 8887 2493
rect 8876 2476 8883 2480
rect 8776 2436 8803 2443
rect 8816 2440 8823 2443
rect 8796 2256 8803 2436
rect 8813 2427 8827 2440
rect 8856 2387 8863 2443
rect 8816 2203 8823 2223
rect 8856 2220 8863 2223
rect 8853 2207 8867 2220
rect 8816 2196 8843 2203
rect 8696 1970 8703 2033
rect 8733 1960 8747 1973
rect 8736 1956 8743 1960
rect 8656 1603 8663 1793
rect 8716 1736 8723 1853
rect 8676 1696 8703 1703
rect 8736 1700 8743 1703
rect 8676 1627 8683 1696
rect 8733 1687 8747 1700
rect 8656 1596 8683 1603
rect 8616 1450 8623 1533
rect 8556 1367 8563 1403
rect 8596 1230 8603 1403
rect 8620 1183 8633 1187
rect 8496 907 8503 993
rect 8516 827 8523 953
rect 8496 767 8503 793
rect 8496 547 8503 696
rect 8016 380 8023 383
rect 8013 367 8027 380
rect 7936 327 7943 363
rect 8076 267 8083 383
rect 8096 327 8103 353
rect 7656 187 7663 253
rect 6716 27 6723 173
rect 7653 160 7667 173
rect 7656 156 7663 160
rect 6776 -24 6783 13
rect 7036 -17 7043 143
rect 7556 27 7563 143
rect 7696 27 7703 150
rect 8056 67 8063 153
rect 8116 124 8123 413
rect 8176 67 8183 253
rect 8276 176 8283 273
rect 8396 67 8403 383
rect 8476 167 8483 433
rect 8536 176 8543 773
rect 8556 707 8563 1173
rect 8576 1087 8583 1183
rect 8616 1176 8633 1183
rect 8620 1173 8633 1176
rect 8656 1087 8663 1436
rect 8576 1007 8583 1073
rect 8587 753 8593 767
rect 8636 697 8643 953
rect 8676 916 8683 1596
rect 8696 1287 8703 1673
rect 8756 1407 8763 1673
rect 8796 1607 8803 2053
rect 8816 1627 8823 1956
rect 8836 1867 8843 2196
rect 8856 1747 8863 2172
rect 8936 2167 8943 3253
rect 8956 3187 8963 3263
rect 8956 2267 8963 3053
rect 8976 2667 8983 3053
rect 8996 2744 9003 2933
rect 9016 2867 9023 3053
rect 9036 2847 9043 3273
rect 9056 2887 9063 3993
rect 9076 3327 9083 4016
rect 9093 3987 9107 3993
rect 9096 3467 9103 3952
rect 9096 3023 9103 3453
rect 9116 3047 9123 4793
rect 9136 3687 9143 4813
rect 9156 3967 9163 5336
rect 9176 5043 9183 5293
rect 9196 5287 9203 5343
rect 9256 5076 9263 5113
rect 9176 5036 9203 5043
rect 9176 4707 9183 4873
rect 9196 4807 9203 5036
rect 9236 5023 9243 5043
rect 9316 5043 9323 5473
rect 9296 5036 9323 5043
rect 9216 5016 9243 5023
rect 9176 4067 9183 4672
rect 9196 4524 9203 4753
rect 9196 4307 9203 4433
rect 9216 4207 9223 5016
rect 9236 4787 9243 4853
rect 9256 4827 9263 5013
rect 9276 4607 9283 4953
rect 9296 4787 9303 5036
rect 9356 4856 9363 5413
rect 9376 5047 9383 5473
rect 9536 5427 9543 5813
rect 9556 5687 9563 5863
rect 9396 5247 9403 5376
rect 9396 4927 9403 4953
rect 9416 4907 9423 5076
rect 9316 4687 9323 4810
rect 9336 4803 9343 4823
rect 9336 4796 9363 4803
rect 9356 4747 9363 4796
rect 9267 4576 9323 4583
rect 9316 4556 9323 4576
rect 9336 4570 9343 4653
rect 9356 4527 9363 4733
rect 9256 4336 9263 4433
rect 9253 4127 9267 4133
rect 9176 3887 9183 3993
rect 9236 3983 9243 4003
rect 9207 3976 9243 3983
rect 9176 3627 9183 3873
rect 9196 3787 9203 3913
rect 9196 3687 9203 3752
rect 9136 3267 9143 3613
rect 9156 3447 9163 3513
rect 9156 3067 9163 3433
rect 9216 3427 9223 3873
rect 9256 3863 9263 3953
rect 9276 3887 9283 4233
rect 9336 4227 9343 4393
rect 9376 4307 9383 4773
rect 9436 4747 9443 5233
rect 9456 4647 9463 5213
rect 9476 5167 9483 5330
rect 9556 5167 9563 5493
rect 9576 5307 9583 5793
rect 9596 5347 9603 5376
rect 9476 4807 9483 5153
rect 9596 5007 9603 5093
rect 9616 4983 9623 5813
rect 9636 5227 9643 6293
rect 9656 5584 9663 6453
rect 9713 6420 9727 6433
rect 9716 6416 9723 6420
rect 9736 6347 9743 6383
rect 9776 6307 9783 6383
rect 9836 6327 9843 6513
rect 9956 6430 9963 6513
rect 9996 6416 10003 6533
rect 9676 5487 9683 6253
rect 9896 6084 9903 6116
rect 9716 5987 9723 6083
rect 9756 6027 9763 6083
rect 9796 5896 9803 5933
rect 9876 5910 9883 5953
rect 9716 5627 9723 5896
rect 9876 5867 9883 5896
rect 9713 5600 9727 5613
rect 9776 5610 9783 5853
rect 9716 5596 9723 5600
rect 9656 5344 9663 5453
rect 9736 5376 9743 5473
rect 9716 5247 9723 5343
rect 9796 5307 9803 5550
rect 9596 4976 9623 4983
rect 9476 4767 9483 4793
rect 9396 4447 9403 4553
rect 9296 4004 9303 4113
rect 9336 4007 9343 4073
rect 9256 3856 9283 3863
rect 9276 3816 9283 3856
rect 9256 3707 9263 3783
rect 9256 3516 9263 3633
rect 9296 3530 9303 3713
rect 9356 3487 9363 4193
rect 9416 3967 9423 4413
rect 9436 4327 9443 4433
rect 9456 4247 9463 4633
rect 9496 4343 9503 4873
rect 9516 4587 9523 4856
rect 9536 4687 9543 4973
rect 9556 4824 9563 4933
rect 9596 4887 9603 4976
rect 9636 4856 9643 5053
rect 9676 5047 9683 5113
rect 9696 5003 9703 5076
rect 9696 4996 9723 5003
rect 9556 4567 9563 4713
rect 9576 4707 9583 4856
rect 9576 4556 9583 4693
rect 9656 4527 9663 4823
rect 9536 4520 9543 4523
rect 9533 4507 9547 4520
rect 9487 4336 9503 4343
rect 9513 4340 9527 4353
rect 9516 4336 9523 4340
rect 9436 4147 9443 4173
rect 9476 4127 9483 4336
rect 9476 4036 9483 4113
rect 9416 3887 9423 3913
rect 9256 3267 9263 3413
rect 9276 3367 9283 3483
rect 9316 3367 9323 3483
rect 9176 3227 9183 3253
rect 9096 3016 9123 3023
rect 9116 2996 9123 3016
rect 8836 1547 8843 1733
rect 8876 1567 8883 2133
rect 8996 1983 9003 2513
rect 9016 2067 9023 2793
rect 9116 2776 9123 2853
rect 9136 2807 9143 2963
rect 9156 2867 9163 2933
rect 9076 2687 9083 2713
rect 9096 2667 9103 2743
rect 9056 2490 9063 2533
rect 9093 2480 9107 2493
rect 9096 2476 9103 2480
rect 9156 2476 9163 2553
rect 9056 2444 9063 2476
rect 9076 2187 9083 2223
rect 9116 2167 9123 2223
rect 8996 1976 9023 1983
rect 8916 1807 8923 1973
rect 9016 1956 9023 1976
rect 9076 1927 9083 2013
rect 9096 1927 9103 2153
rect 8896 1667 8903 1753
rect 8916 1687 8923 1793
rect 8996 1767 9003 1923
rect 9036 1920 9063 1923
rect 9036 1916 9067 1920
rect 9053 1907 9067 1916
rect 8947 1743 8960 1747
rect 8947 1736 8963 1743
rect 8947 1733 8960 1736
rect 8933 1667 8947 1673
rect 8976 1647 8983 1673
rect 8996 1647 9003 1703
rect 9036 1647 9043 1673
rect 9056 1647 9063 1853
rect 9076 1667 9083 1753
rect 8836 1447 8843 1533
rect 8856 1436 8863 1553
rect 8716 1067 8723 1253
rect 8756 1187 8763 1393
rect 8816 1230 8823 1273
rect 8856 1216 8863 1353
rect 8776 1184 8783 1213
rect 8836 1147 8843 1183
rect 8736 1047 8743 1113
rect 8716 879 8723 883
rect 8713 867 8727 879
rect 8776 787 8783 883
rect 8816 707 8823 893
rect 8836 867 8843 1133
rect 8916 947 8923 1293
rect 8936 1147 8943 1216
rect 8956 1187 8963 1613
rect 9136 1503 9143 2213
rect 9196 2207 9203 2873
rect 9156 1547 9163 2193
rect 9176 2107 9183 2133
rect 9176 1907 9183 2033
rect 9216 2027 9223 3033
rect 9236 2447 9243 3213
rect 9256 3067 9263 3153
rect 9256 2587 9263 2996
rect 9276 2927 9283 3313
rect 9316 3187 9323 3353
rect 9336 2947 9343 3473
rect 9356 3387 9363 3413
rect 9376 3207 9383 3770
rect 9396 3727 9403 3816
rect 9456 3487 9463 3990
rect 9536 3867 9543 4290
rect 9476 3747 9483 3816
rect 9516 3780 9523 3783
rect 9513 3767 9527 3780
rect 9507 3713 9513 3727
rect 9476 3467 9483 3533
rect 9536 3527 9543 3633
rect 9556 3516 9563 3673
rect 9516 3480 9523 3483
rect 9496 3443 9503 3473
rect 9513 3467 9527 3480
rect 9496 3436 9523 3443
rect 9407 3413 9413 3427
rect 9496 3367 9503 3393
rect 9516 3367 9523 3436
rect 9536 3367 9543 3433
rect 9596 3427 9603 4513
rect 9616 4407 9623 4473
rect 9376 2996 9383 3153
rect 9476 3127 9483 3263
rect 9536 3227 9543 3296
rect 9496 3147 9503 3193
rect 9276 2427 9283 2913
rect 9416 2907 9423 2963
rect 9336 2776 9343 2853
rect 9316 2727 9323 2743
rect 9356 2740 9363 2743
rect 9353 2727 9367 2740
rect 9316 2323 9323 2713
rect 9476 2587 9483 2713
rect 9356 2476 9363 2573
rect 9393 2480 9407 2493
rect 9396 2476 9403 2480
rect 9296 2316 9323 2323
rect 9296 2227 9303 2316
rect 9356 2256 9363 2413
rect 9176 1667 9183 1872
rect 9196 1867 9203 1956
rect 9216 1847 9223 2013
rect 9256 1970 9263 2073
rect 9336 2067 9343 2223
rect 9376 2187 9383 2223
rect 9393 2207 9407 2213
rect 9416 2207 9423 2273
rect 9373 2167 9387 2173
rect 9313 1987 9327 1993
rect 9236 1736 9243 1913
rect 9207 1633 9213 1647
rect 9256 1627 9263 1703
rect 9356 1627 9363 1956
rect 9376 1727 9383 2093
rect 9436 2047 9443 2493
rect 9456 2347 9463 2493
rect 9456 2067 9463 2333
rect 9476 2107 9483 2573
rect 9496 2387 9503 3133
rect 9536 3107 9543 3133
rect 9556 2627 9563 3293
rect 9576 2927 9583 3353
rect 9596 3247 9603 3413
rect 9616 3327 9623 4393
rect 9633 4350 9647 4353
rect 9636 4267 9643 4336
rect 9656 4287 9663 4373
rect 9676 4107 9683 4593
rect 9716 4427 9723 4996
rect 9696 4187 9703 4273
rect 9716 4167 9723 4413
rect 9736 4387 9743 5293
rect 9816 5207 9823 5863
rect 9856 5147 9863 5193
rect 9793 5080 9807 5093
rect 9796 5076 9803 5080
rect 9876 5044 9883 5433
rect 9896 5007 9903 6070
rect 9916 5887 9923 6393
rect 9976 6347 9983 6383
rect 10056 6327 10063 6413
rect 9936 5983 9943 6233
rect 9996 6116 10003 6193
rect 10096 6187 10103 6616
rect 9936 5976 9963 5983
rect 9936 5387 9943 5933
rect 9956 5807 9963 5976
rect 10016 5767 10023 6013
rect 10076 5896 10083 6153
rect 10096 6047 10103 6093
rect 10116 6027 10123 6936
rect 10276 6904 10283 6953
rect 10156 6867 10163 6903
rect 10136 6347 10143 6793
rect 10196 6707 10203 6903
rect 10036 5627 10043 5733
rect 10033 5600 10047 5613
rect 10056 5607 10063 5850
rect 10096 5747 10103 5863
rect 10136 5827 10143 6153
rect 10036 5596 10043 5600
rect 9956 5556 9983 5563
rect 9956 5527 9963 5556
rect 9776 4467 9783 4993
rect 9956 4987 9963 5053
rect 9896 4927 9903 4953
rect 9836 4556 9843 4893
rect 9896 4627 9903 4823
rect 9936 4820 9943 4823
rect 9933 4807 9947 4820
rect 9976 4787 9983 5533
rect 10096 5527 10103 5693
rect 10116 5564 10123 5593
rect 9996 5336 10023 5343
rect 9996 5247 10003 5336
rect 9996 5067 10003 5113
rect 9816 4503 9823 4523
rect 9816 4496 9843 4503
rect 9753 4340 9767 4353
rect 9796 4350 9803 4433
rect 9756 4336 9763 4340
rect 9776 4247 9783 4303
rect 9693 4040 9707 4053
rect 9696 4036 9703 4040
rect 9656 3784 9663 4033
rect 9636 3107 9643 3753
rect 9656 3467 9663 3553
rect 9656 3027 9663 3453
rect 9676 3267 9683 3653
rect 9696 3307 9703 3853
rect 9716 3647 9723 4003
rect 9776 3816 9783 3993
rect 9816 3983 9823 4093
rect 9836 4007 9843 4496
rect 9856 4487 9863 4523
rect 9856 4007 9863 4452
rect 9876 4167 9883 4336
rect 9816 3976 9843 3983
rect 9836 3827 9843 3976
rect 9796 3780 9803 3783
rect 9793 3767 9807 3780
rect 9856 3587 9863 3816
rect 9876 3727 9883 4033
rect 9896 3784 9903 4553
rect 9793 3520 9807 3533
rect 9796 3516 9803 3520
rect 9820 3483 9833 3487
rect 9776 3407 9783 3483
rect 9816 3476 9833 3483
rect 9820 3473 9833 3476
rect 9753 3300 9767 3313
rect 9756 3296 9763 3300
rect 9736 3260 9743 3263
rect 9733 3247 9747 3260
rect 9816 3263 9823 3393
rect 9796 3256 9823 3263
rect 9716 2964 9723 3013
rect 9616 2776 9623 2893
rect 9596 2727 9603 2743
rect 9636 2740 9643 2743
rect 9633 2727 9647 2740
rect 9516 2187 9523 2210
rect 9556 2203 9563 2613
rect 9596 2487 9603 2713
rect 9636 2476 9643 2553
rect 9696 2447 9703 2813
rect 9616 2440 9623 2443
rect 9613 2427 9627 2440
rect 9616 2256 9623 2293
rect 9536 2196 9563 2203
rect 9116 1496 9143 1503
rect 9116 1436 9123 1496
rect 9067 1403 9080 1407
rect 9067 1396 9083 1403
rect 9067 1393 9080 1396
rect 9156 1347 9163 1433
rect 9156 1216 9163 1253
rect 9107 1183 9120 1187
rect 9107 1176 9123 1183
rect 9107 1173 9120 1176
rect 9196 1147 9203 1593
rect 9036 916 9043 993
rect 9016 863 9023 883
rect 9016 856 9043 863
rect 8656 660 8663 663
rect 8653 647 8667 660
rect 8676 396 8683 433
rect 8736 364 8743 693
rect 8836 647 8843 853
rect 8936 696 8943 753
rect 8976 696 8983 813
rect 9036 711 9043 856
rect 9056 787 9063 883
rect 8956 567 8963 663
rect 8996 627 9003 650
rect 9036 647 9043 697
rect 8756 176 8763 553
rect 8916 447 8923 553
rect 8916 396 8923 433
rect 8956 396 8963 433
rect 9016 176 9023 553
rect 9076 144 9083 433
rect 9096 327 9103 1133
rect 9216 1087 9223 1213
rect 9196 1027 9203 1053
rect 9236 987 9243 1533
rect 9376 1436 9383 1713
rect 9416 1707 9423 1973
rect 9436 1404 9443 1953
rect 9456 1924 9463 2053
rect 9536 1967 9543 2196
rect 9556 1956 9563 2173
rect 9516 1920 9523 1923
rect 9513 1907 9527 1920
rect 9473 1750 9487 1753
rect 9516 1736 9523 1813
rect 9536 1700 9543 1703
rect 9533 1687 9547 1700
rect 9576 1587 9583 1893
rect 9596 1847 9603 2189
rect 9596 1687 9603 1833
rect 9336 1267 9343 1403
rect 9356 1107 9363 1183
rect 9396 1147 9403 1183
rect 9136 367 9143 973
rect 9216 696 9223 933
rect 9296 916 9303 1033
rect 9336 879 9343 883
rect 9333 867 9347 879
rect 9396 787 9403 883
rect 9196 627 9203 663
rect 9196 447 9203 613
rect 9236 427 9243 663
rect 9213 400 9227 413
rect 9216 396 9223 400
rect 9196 327 9203 363
rect 9216 144 9223 193
rect 9276 176 9283 693
rect 9436 664 9443 1093
rect 9476 1067 9483 1493
rect 9473 723 9487 733
rect 9496 723 9503 1553
rect 9616 1436 9623 2193
rect 9636 2087 9643 2223
rect 9656 1927 9663 2133
rect 9636 1607 9643 1736
rect 9676 1704 9683 1793
rect 9696 1607 9703 2412
rect 9716 1967 9723 2473
rect 9736 2247 9743 2993
rect 9756 2427 9763 3093
rect 9776 2907 9783 3250
rect 9796 3167 9803 3256
rect 9796 2964 9803 3153
rect 9836 3067 9843 3153
rect 9856 3107 9863 3573
rect 9876 3487 9883 3713
rect 9876 3207 9883 3473
rect 9896 3247 9903 3633
rect 9916 3207 9923 4773
rect 9933 4487 9947 4493
rect 9936 4007 9943 4290
rect 9956 4107 9963 4493
rect 10016 4487 10023 5313
rect 10096 5267 10103 5376
rect 10036 5187 10043 5233
rect 10033 5087 10047 5093
rect 10056 5076 10063 5173
rect 10116 5076 10123 5153
rect 10156 5043 10163 6553
rect 10176 6247 10183 6673
rect 10236 6604 10243 6733
rect 10216 6384 10223 6453
rect 10256 6447 10263 6693
rect 10296 6636 10303 6693
rect 10336 6687 10343 7133
rect 10496 7124 10503 7233
rect 10336 6507 10343 6533
rect 10356 6527 10363 6573
rect 10247 6423 10260 6427
rect 10247 6416 10263 6423
rect 10293 6420 10307 6433
rect 10296 6416 10303 6420
rect 10247 6413 10260 6416
rect 10316 6376 10343 6383
rect 10176 5927 10183 6133
rect 10176 5327 10183 5892
rect 10196 5847 10203 6253
rect 10236 6147 10243 6333
rect 10233 6120 10247 6133
rect 10236 6116 10243 6120
rect 10276 6116 10283 6193
rect 10256 6063 10263 6083
rect 10236 6056 10263 6063
rect 10236 5907 10243 6056
rect 10296 6027 10303 6083
rect 10196 5167 10203 5833
rect 10256 5747 10263 5913
rect 10336 5910 10343 6376
rect 10356 6047 10363 6513
rect 10376 6047 10383 6370
rect 10416 6347 10423 7093
rect 10516 7047 10523 7393
rect 10536 7107 10543 7556
rect 10556 7170 10563 8233
rect 10596 7990 10603 8433
rect 10676 8196 10683 8393
rect 10576 7427 10583 7953
rect 10616 7887 10623 7973
rect 10636 7807 10643 8163
rect 10716 8027 10723 8553
rect 10756 8464 10763 8493
rect 10696 7644 10703 7793
rect 10596 7470 10603 7573
rect 10716 7507 10723 7943
rect 10676 7467 10683 7493
rect 10576 7287 10583 7413
rect 10656 7307 10663 7456
rect 10476 6936 10483 6993
rect 10516 6936 10523 7033
rect 10576 6904 10583 7193
rect 10676 7156 10683 7413
rect 10616 7120 10623 7123
rect 10613 7107 10627 7120
rect 10656 7047 10663 7123
rect 10456 6867 10463 6903
rect 10436 6547 10443 6633
rect 10373 5900 10387 5913
rect 10376 5896 10383 5900
rect 10076 4947 10083 5043
rect 10136 5036 10163 5043
rect 10076 4556 10083 4653
rect 10056 4520 10063 4523
rect 10053 4507 10067 4520
rect 9976 4207 9983 4473
rect 10056 4336 10063 4433
rect 9956 3847 9963 4093
rect 9996 4067 10003 4336
rect 10076 4283 10083 4303
rect 10056 4276 10083 4283
rect 10056 4247 10063 4276
rect 9973 4050 9987 4053
rect 9993 4040 10007 4053
rect 9996 4036 10003 4040
rect 10076 4043 10083 4253
rect 10076 4036 10103 4043
rect 10096 4004 10103 4036
rect 10116 3967 10123 4193
rect 9996 3867 10003 3953
rect 10036 3816 10043 3953
rect 9936 3047 9943 3193
rect 9956 3147 9963 3812
rect 10136 3783 10143 5036
rect 10196 4856 10203 5093
rect 10216 4887 10223 5593
rect 10276 5527 10283 5563
rect 10276 5376 10283 5413
rect 10256 5287 10263 5343
rect 10156 4524 10163 4793
rect 10176 4587 10183 4823
rect 10156 4207 10163 4373
rect 10176 4347 10183 4573
rect 10096 3776 10123 3783
rect 10136 3776 10153 3783
rect 10056 3747 10063 3770
rect 10116 3763 10123 3776
rect 10116 3756 10143 3763
rect 9996 3296 10003 3513
rect 10016 3487 10023 3673
rect 10096 3530 10103 3753
rect 10113 3707 10127 3713
rect 10047 3523 10060 3527
rect 10047 3516 10063 3523
rect 10136 3527 10143 3756
rect 10047 3513 10060 3516
rect 9896 2996 9903 3033
rect 9936 2996 9943 3033
rect 9856 2776 9863 2913
rect 9916 2827 9923 2963
rect 9996 2887 10003 3233
rect 10016 3107 10023 3263
rect 10056 3260 10063 3263
rect 10053 3247 10067 3260
rect 9636 1367 9643 1403
rect 9616 1267 9623 1293
rect 9616 1216 9623 1253
rect 9656 1107 9663 1183
rect 9636 916 9643 973
rect 9676 916 9683 1013
rect 9616 880 9623 883
rect 9613 867 9627 880
rect 9473 720 9503 723
rect 9476 716 9503 720
rect 9476 696 9483 716
rect 9513 700 9527 713
rect 9516 696 9523 700
rect 9576 687 9583 813
rect 9696 663 9703 713
rect 9716 707 9723 1453
rect 9736 867 9743 2233
rect 9776 2207 9783 2730
rect 9856 2307 9863 2693
rect 9916 2607 9923 2743
rect 9896 2476 9903 2533
rect 9916 2407 9923 2443
rect 9876 2256 9883 2373
rect 9776 1956 9783 2172
rect 9796 2087 9803 2256
rect 9856 2187 9863 2223
rect 9896 2027 9903 2223
rect 9816 1736 9823 1813
rect 9876 1703 9883 1956
rect 9896 1847 9903 2013
rect 9893 1727 9907 1733
rect 9836 1647 9843 1703
rect 9856 1696 9883 1703
rect 9856 1567 9863 1696
rect 9756 696 9763 1313
rect 9816 1167 9823 1553
rect 9876 1436 9883 1533
rect 9916 1467 9923 2213
rect 9936 2187 9943 2273
rect 9956 2227 9963 2353
rect 9976 2347 9983 2430
rect 10016 2427 10023 2973
rect 9936 1727 9943 1873
rect 9956 1647 9963 1736
rect 9856 1400 9863 1403
rect 9853 1387 9867 1400
rect 9896 1367 9903 1403
rect 9916 1216 9923 1273
rect 9836 787 9843 1216
rect 9896 1147 9903 1183
rect 9916 916 9923 1153
rect 9956 1107 9963 1612
rect 9976 1187 9983 2333
rect 10036 2227 10043 2873
rect 10056 2367 10063 3212
rect 9996 1927 10003 2193
rect 10036 1956 10043 2073
rect 10076 2027 10083 3193
rect 10096 2747 10103 3453
rect 10116 3247 10123 3483
rect 10136 3227 10143 3473
rect 10156 3467 10163 3770
rect 10176 3567 10183 3833
rect 10196 3767 10203 4773
rect 10216 3907 10223 4823
rect 10256 4043 10263 4873
rect 10276 4627 10283 5253
rect 10296 5207 10303 5293
rect 10356 5267 10363 5863
rect 10296 4787 10303 5193
rect 10396 5090 10403 5330
rect 10416 5307 10423 5793
rect 10456 5683 10463 6653
rect 10476 6384 10483 6713
rect 10496 6587 10503 6903
rect 10596 6667 10603 6953
rect 10536 6607 10543 6636
rect 10676 6607 10683 6773
rect 10536 6416 10543 6513
rect 10516 6363 10523 6383
rect 10516 6356 10543 6363
rect 10536 6116 10543 6356
rect 10516 6080 10523 6083
rect 10513 6067 10527 6080
rect 10496 5687 10503 5893
rect 10436 5676 10463 5683
rect 10436 5107 10443 5676
rect 10456 5347 10463 5633
rect 10516 5596 10523 6032
rect 10596 5987 10603 6593
rect 10616 6467 10623 6603
rect 10696 6267 10703 6993
rect 10756 6970 10763 7613
rect 10776 6967 10783 9393
rect 10816 9043 10823 9453
rect 10836 9407 10843 9533
rect 10856 9467 10863 9553
rect 10876 9550 10883 10113
rect 10956 10056 10963 10133
rect 10996 10056 11003 10093
rect 11016 10087 11023 10796
rect 11036 10487 11043 10973
rect 11076 10810 11083 10893
rect 11116 10796 11123 11173
rect 11196 10827 11203 11773
rect 11216 11227 11223 11853
rect 11353 11840 11367 11853
rect 11356 11836 11363 11840
rect 11396 11807 11403 11856
rect 11296 11630 11303 11803
rect 11416 11707 11423 11833
rect 11596 11800 11603 11803
rect 11593 11787 11607 11800
rect 11033 10467 11047 10473
rect 10936 9987 10943 10023
rect 10976 9927 10983 10023
rect 10973 9767 10987 9773
rect 10960 9723 10973 9727
rect 10956 9716 10973 9723
rect 10960 9713 10973 9716
rect 10876 9327 10883 9536
rect 10916 9307 10923 9573
rect 10996 9536 11003 9933
rect 11016 9587 11023 9733
rect 10976 9427 10983 9503
rect 10876 9276 10913 9283
rect 10876 9236 10883 9276
rect 10856 9200 10863 9203
rect 10853 9187 10867 9200
rect 10936 9203 10943 9373
rect 10916 9196 10943 9203
rect 10816 9036 10843 9043
rect 10796 7207 10803 9013
rect 10816 7707 10823 8793
rect 10836 7587 10843 9036
rect 10896 9027 10903 9190
rect 10916 9030 10923 9196
rect 10956 9147 10963 9273
rect 10996 9204 11003 9253
rect 10956 9030 10963 9093
rect 10856 8887 10863 9016
rect 10936 8767 10943 8983
rect 10876 8510 10883 8753
rect 11016 8730 11023 9293
rect 10936 8567 10943 8683
rect 10976 8680 10983 8683
rect 10973 8667 10987 8680
rect 10913 8500 10927 8513
rect 10916 8496 10923 8500
rect 10896 8460 10903 8463
rect 10893 8447 10907 8460
rect 10996 8447 11003 8553
rect 10876 7944 10883 8313
rect 10916 8196 10923 8233
rect 10996 8163 11003 8333
rect 10936 8127 10943 8163
rect 10976 8156 11003 8163
rect 10896 8007 10903 8093
rect 10976 7976 10983 8156
rect 11016 7987 11023 8513
rect 10916 7707 10923 7973
rect 10996 7867 11003 7943
rect 10976 7644 10983 7693
rect 10876 7640 10883 7643
rect 10873 7627 10887 7640
rect 10796 6936 10803 7033
rect 10616 5987 10623 6173
rect 10536 5847 10543 5973
rect 10593 5900 10607 5913
rect 10596 5896 10603 5900
rect 10576 5807 10583 5863
rect 10476 5556 10503 5563
rect 10356 4707 10363 5043
rect 10436 5027 10443 5072
rect 10456 5027 10463 5233
rect 10476 5227 10483 5556
rect 10516 5376 10523 5473
rect 10596 5307 10603 5376
rect 10496 5067 10503 5113
rect 10396 4867 10403 4893
rect 10427 4863 10440 4867
rect 10427 4856 10443 4863
rect 10476 4856 10483 5013
rect 10516 4867 10523 5153
rect 10427 4853 10440 4856
rect 10376 4807 10383 4853
rect 10316 4556 10323 4693
rect 10356 4627 10363 4693
rect 10276 4516 10293 4523
rect 10276 4304 10283 4516
rect 10336 4467 10343 4523
rect 10336 4336 10343 4393
rect 10396 4387 10403 4556
rect 10416 4507 10423 4613
rect 10316 4067 10323 4303
rect 10356 4283 10363 4303
rect 10356 4280 10383 4283
rect 10353 4276 10383 4280
rect 10353 4267 10367 4276
rect 10236 4036 10263 4043
rect 10316 4036 10323 4053
rect 10216 3707 10223 3893
rect 10176 3487 10183 3516
rect 10216 3343 10223 3413
rect 10196 3336 10223 3343
rect 10156 3247 10163 3296
rect 10136 3067 10143 3093
rect 10136 2776 10143 3032
rect 10196 2996 10203 3336
rect 10236 3007 10243 4036
rect 10356 4004 10363 4193
rect 10353 3867 10367 3873
rect 10313 3820 10327 3833
rect 10316 3816 10323 3820
rect 10256 3703 10263 3816
rect 10287 3713 10293 3727
rect 10256 3696 10283 3703
rect 10256 3307 10263 3516
rect 10276 3483 10283 3696
rect 10336 3587 10343 3783
rect 10376 3587 10383 4276
rect 10416 4247 10423 4336
rect 10396 3547 10403 4073
rect 10416 3830 10423 3873
rect 10413 3607 10427 3613
rect 10356 3516 10403 3523
rect 10276 3476 10303 3483
rect 10296 3296 10303 3476
rect 10396 3483 10403 3516
rect 10376 3476 10403 3483
rect 10376 3310 10383 3476
rect 10220 2963 10233 2967
rect 10176 2927 10183 2963
rect 10216 2956 10233 2963
rect 10220 2953 10233 2956
rect 10156 2740 10163 2743
rect 10153 2727 10167 2740
rect 10176 2447 10183 2733
rect 10176 2407 10183 2433
rect 10127 2396 10153 2403
rect 10196 2367 10203 2713
rect 10216 2487 10223 2913
rect 10256 2567 10263 3233
rect 10156 2256 10163 2353
rect 10216 2347 10223 2373
rect 10056 1867 10063 1923
rect 9993 1727 10007 1733
rect 10096 1707 10103 1910
rect 10116 1787 10123 1956
rect 10136 1887 10143 2223
rect 10176 2167 10183 2223
rect 10236 2183 10243 2430
rect 10256 2407 10263 2553
rect 10256 2270 10263 2393
rect 10276 2387 10283 3133
rect 10296 2967 10303 3173
rect 10316 2727 10323 3263
rect 10376 3127 10383 3296
rect 10396 3227 10403 3433
rect 10416 3203 10423 3572
rect 10436 3543 10443 4733
rect 10516 4647 10523 4753
rect 10476 4227 10483 4613
rect 10536 4207 10543 5293
rect 10556 4883 10563 5093
rect 10616 5076 10623 5833
rect 10636 5287 10643 5513
rect 10596 5040 10603 5043
rect 10593 5027 10607 5040
rect 10556 4876 10583 4883
rect 10556 4607 10563 4856
rect 10576 4563 10583 4876
rect 10596 4824 10603 4893
rect 10556 4556 10583 4563
rect 10593 4560 10607 4573
rect 10596 4556 10603 4560
rect 10636 4556 10643 4653
rect 10656 4587 10663 4853
rect 10676 4787 10683 6053
rect 10696 4867 10703 6193
rect 10716 5527 10723 6935
rect 10736 6167 10743 6433
rect 10756 6384 10763 6853
rect 10776 6567 10783 6903
rect 10836 6467 10843 7173
rect 10856 6867 10863 7253
rect 10876 7007 10883 7456
rect 10896 7167 10903 7553
rect 11016 7487 11023 7673
rect 11036 7463 11043 10393
rect 11056 9287 11063 10713
rect 11096 10523 11103 10763
rect 11216 10727 11223 11133
rect 11236 11027 11243 11616
rect 11296 11427 11303 11616
rect 11296 11096 11303 11413
rect 11356 11316 11363 11353
rect 11376 11147 11383 11283
rect 11436 11187 11443 11316
rect 11456 11163 11463 11353
rect 11436 11156 11463 11163
rect 11216 10590 11223 10692
rect 11236 10687 11243 10913
rect 11256 10667 11263 10853
rect 11276 10764 11283 11050
rect 11256 10544 11263 10653
rect 11276 10590 11283 10750
rect 11196 10527 11203 10543
rect 11096 10516 11123 10523
rect 11076 9263 11083 10473
rect 11096 10427 11103 10493
rect 11096 9724 11103 10273
rect 11076 9256 11103 9263
rect 11056 8527 11063 9173
rect 11076 8747 11083 9233
rect 11096 8967 11103 9256
rect 11116 9247 11123 10516
rect 11196 10513 11213 10527
rect 11136 9787 11143 10053
rect 11156 10007 11163 10473
rect 11176 10147 11183 10353
rect 11196 10287 11203 10513
rect 11216 10276 11223 10433
rect 11156 9667 11163 9993
rect 11196 9947 11203 10230
rect 11276 10227 11283 10576
rect 11296 10527 11303 11013
rect 11316 10987 11323 11063
rect 11316 10747 11323 10973
rect 11376 10796 11383 10833
rect 11436 10787 11443 11156
rect 11456 11067 11463 11096
rect 11396 10743 11403 10763
rect 11376 10736 11403 10743
rect 11316 10327 11323 10633
rect 11276 10087 11283 10213
rect 11236 10020 11243 10023
rect 11233 10007 11247 10020
rect 11276 9987 11283 10023
rect 11196 9756 11203 9833
rect 11236 9756 11243 9873
rect 11216 9563 11223 9723
rect 11196 9556 11223 9563
rect 11196 9536 11203 9556
rect 11133 9287 11147 9293
rect 11127 9236 11143 9243
rect 11176 9236 11183 9293
rect 11216 9267 11223 9503
rect 11196 9183 11203 9203
rect 11176 9176 11203 9183
rect 11176 9016 11183 9176
rect 11216 9027 11223 9113
rect 11156 8980 11163 8983
rect 11153 8967 11167 8980
rect 11236 8807 11243 9273
rect 11253 9187 11267 9193
rect 11276 9187 11283 9753
rect 11256 9030 11263 9053
rect 11256 8867 11263 9016
rect 11296 8984 11303 9413
rect 11316 9287 11323 10073
rect 11336 9550 11343 10713
rect 11356 10487 11363 10576
rect 11376 10547 11383 10736
rect 11376 10427 11383 10533
rect 11413 10507 11427 10513
rect 11476 10407 11483 11693
rect 11636 11616 11683 11623
rect 11576 11347 11583 11583
rect 11676 11343 11683 11616
rect 11696 11587 11703 11790
rect 11656 11336 11683 11343
rect 11496 10587 11503 11333
rect 11576 11316 11623 11323
rect 11656 11316 11663 11336
rect 11576 11247 11583 11316
rect 11596 11223 11603 11270
rect 11576 11216 11603 11223
rect 11576 11096 11583 11216
rect 11396 10244 11403 10373
rect 11516 10147 11523 10273
rect 11536 10107 11543 10813
rect 11356 9807 11363 10013
rect 11396 9707 11403 10093
rect 11536 10056 11543 10093
rect 11556 10067 11563 11063
rect 11596 11023 11603 11050
rect 11576 11016 11603 11023
rect 11576 10907 11583 11016
rect 11636 10907 11643 11233
rect 11676 11127 11683 11173
rect 11416 9887 11423 10053
rect 11496 9927 11503 10023
rect 11336 9504 11343 9536
rect 11416 9504 11423 9873
rect 11496 9720 11503 9723
rect 11493 9707 11507 9720
rect 11536 9587 11543 9973
rect 11536 9536 11543 9573
rect 11476 9447 11483 9503
rect 11193 8720 11207 8733
rect 11196 8716 11203 8720
rect 11136 8496 11143 8553
rect 11156 8547 11163 8716
rect 11216 8680 11223 8683
rect 11213 8667 11227 8680
rect 11256 8647 11263 8683
rect 11296 8607 11303 8970
rect 11336 8967 11343 9253
rect 11356 8730 11363 9173
rect 11056 7627 11063 8213
rect 11076 7567 11083 8493
rect 11096 8127 11103 8253
rect 11116 8167 11123 8463
rect 11153 8447 11167 8450
rect 11276 8427 11283 8493
rect 11296 8227 11303 8593
rect 11316 8464 11323 8713
rect 11153 8210 11167 8213
rect 11193 8200 11207 8213
rect 11196 8196 11203 8200
rect 11276 8187 11283 8213
rect 11176 7787 11183 8150
rect 11276 8067 11283 8173
rect 11276 7976 11283 8053
rect 11316 7987 11323 8450
rect 11336 8407 11343 8693
rect 11376 8684 11383 9353
rect 11416 9236 11423 9353
rect 11456 9236 11463 9393
rect 11436 9200 11443 9203
rect 11433 9187 11447 9200
rect 11476 9167 11483 9203
rect 11516 9167 11523 9236
rect 11473 9020 11487 9033
rect 11476 9016 11483 9020
rect 11456 8980 11463 8983
rect 11453 8967 11467 8980
rect 11556 8723 11563 8853
rect 11576 8747 11583 10893
rect 11596 10807 11603 10893
rect 11636 10796 11643 10833
rect 11676 10796 11683 11113
rect 11607 10763 11620 10767
rect 11607 10756 11623 10763
rect 11656 10760 11663 10763
rect 11607 10753 11620 10756
rect 11653 10747 11667 10760
rect 11596 9987 11603 10693
rect 11716 10583 11723 11733
rect 11736 11527 11743 11593
rect 11736 10747 11743 11513
rect 11756 11287 11763 12096
rect 11896 11836 11903 11893
rect 11776 11747 11783 11836
rect 11976 11807 11983 12103
rect 11816 11447 11823 11633
rect 11853 11620 11867 11633
rect 11856 11616 11863 11620
rect 11896 11616 11903 11753
rect 12016 11587 12023 12103
rect 11876 11547 11883 11583
rect 11776 11127 11783 11313
rect 11896 11247 11903 11283
rect 11776 11067 11783 11092
rect 11896 11027 11903 11233
rect 11956 11027 11963 11433
rect 11716 10576 11743 10583
rect 11616 10507 11623 10573
rect 11736 10544 11743 10576
rect 11656 10540 11663 10543
rect 11653 10527 11667 10540
rect 11636 10516 11653 10523
rect 11616 10107 11623 10493
rect 11596 8787 11603 9573
rect 11556 8716 11583 8723
rect 11376 8647 11383 8670
rect 11453 8500 11467 8513
rect 11476 8507 11483 8683
rect 11456 8496 11463 8500
rect 11196 7903 11203 7973
rect 11336 7944 11343 8393
rect 11356 8267 11363 8496
rect 11196 7896 11223 7903
rect 11196 7767 11203 7873
rect 11196 7644 11203 7753
rect 11116 7587 11123 7643
rect 11036 7456 11063 7463
rect 10936 7403 10943 7423
rect 10936 7396 10963 7403
rect 10956 7267 10963 7396
rect 10956 7156 10963 7253
rect 10976 7187 10983 7423
rect 10896 6670 10903 7113
rect 10916 6707 10923 7123
rect 10936 6636 10943 6673
rect 10956 6647 10963 6993
rect 11056 6987 11063 7456
rect 11076 7007 11083 7473
rect 11096 7424 11103 7493
rect 11216 7467 11223 7896
rect 11236 7507 11243 7673
rect 11233 7460 11247 7472
rect 11236 7456 11243 7460
rect 10916 6567 10923 6603
rect 10813 6420 10827 6433
rect 10853 6420 10867 6433
rect 10816 6416 10823 6420
rect 10856 6416 10863 6420
rect 10796 6347 10803 6370
rect 10796 6116 10803 6293
rect 10836 6127 10843 6383
rect 10853 6120 10867 6133
rect 10856 6116 10863 6120
rect 10736 5607 10743 6113
rect 10776 5596 10783 5633
rect 10796 5627 10803 6033
rect 10816 5910 10823 6083
rect 10936 6007 10943 6133
rect 10816 5867 10823 5896
rect 10856 5447 10863 5863
rect 10896 5827 10903 5863
rect 10813 5387 10827 5393
rect 10836 5390 10843 5413
rect 10826 5380 10827 5387
rect 10756 5307 10763 5343
rect 10796 5340 10803 5343
rect 10793 5327 10807 5340
rect 10876 5327 10883 5573
rect 10936 5447 10943 5613
rect 10936 5307 10943 5373
rect 10716 5044 10723 5073
rect 10736 4887 10743 4913
rect 10756 4870 10763 4933
rect 10476 3967 10483 4192
rect 10556 4087 10563 4556
rect 10696 4527 10703 4573
rect 10616 4520 10623 4523
rect 10613 4507 10627 4520
rect 10616 4336 10623 4373
rect 10696 4303 10703 4492
rect 10687 4296 10703 4303
rect 10656 4107 10663 4253
rect 10496 3927 10503 4036
rect 10516 3867 10523 4073
rect 10516 3747 10523 3853
rect 10436 3536 10463 3543
rect 10456 3484 10463 3536
rect 10396 3196 10423 3203
rect 10336 2907 10343 3113
rect 10396 2967 10403 3196
rect 10476 3067 10483 3733
rect 10536 3687 10543 3833
rect 10596 3816 10603 3953
rect 10616 3863 10623 4003
rect 10616 3856 10633 3863
rect 10636 3816 10643 3853
rect 10576 3687 10583 3783
rect 10616 3780 10623 3783
rect 10613 3767 10627 3780
rect 10556 3627 10563 3653
rect 10616 3607 10623 3633
rect 10456 3027 10463 3053
rect 10453 3000 10467 3013
rect 10456 2996 10463 3000
rect 10496 2867 10503 3533
rect 10533 3300 10547 3313
rect 10536 3296 10543 3300
rect 10576 3296 10583 3353
rect 10433 2780 10447 2793
rect 10436 2776 10443 2780
rect 10376 2567 10383 2743
rect 10416 2647 10423 2743
rect 10416 2527 10423 2633
rect 10396 2403 10403 2443
rect 10456 2423 10463 2733
rect 10476 2447 10483 2476
rect 10456 2416 10483 2423
rect 10347 2396 10403 2403
rect 10216 2176 10243 2183
rect 10196 2127 10203 2153
rect 10116 1627 10123 1773
rect 10096 1404 10103 1533
rect 10136 1527 10143 1793
rect 10176 1436 10183 2053
rect 10216 1387 10223 2176
rect 10256 2067 10263 2256
rect 10236 1467 10243 1873
rect 10256 1703 10263 2013
rect 10316 1956 10323 2113
rect 10376 1970 10383 2256
rect 10476 2203 10483 2416
rect 10456 2196 10483 2203
rect 10336 1920 10343 1923
rect 10333 1907 10347 1920
rect 10296 1736 10303 1793
rect 10376 1707 10383 1956
rect 10456 1823 10463 2196
rect 10496 2167 10503 2793
rect 10516 2527 10523 3250
rect 10556 3187 10563 3263
rect 10593 3247 10607 3250
rect 10636 3227 10643 3313
rect 10656 3247 10663 3753
rect 10676 3387 10683 4290
rect 10696 3623 10703 4036
rect 10716 4007 10723 4733
rect 10736 4667 10743 4823
rect 10776 4803 10783 4823
rect 10756 4796 10783 4803
rect 10736 4447 10743 4593
rect 10756 4407 10763 4796
rect 10696 3616 10713 3623
rect 10536 2747 10543 3053
rect 10456 1816 10483 1823
rect 10256 1696 10283 1703
rect 10256 1567 10263 1593
rect 10156 1247 10163 1373
rect 10236 1187 10243 1453
rect 10256 1347 10263 1553
rect 10256 1147 10263 1216
rect 10276 1187 10283 1696
rect 10256 1067 10263 1133
rect 9896 787 9903 883
rect 9936 827 9943 883
rect 9976 787 9983 953
rect 10176 916 10183 1053
rect 10156 827 10163 883
rect 10196 876 10223 883
rect 9536 627 9543 663
rect 9696 656 9743 663
rect 9413 427 9427 433
rect 9416 396 9423 413
rect 9476 396 9483 533
rect 9296 287 9303 396
rect 9456 360 9463 363
rect 9453 347 9467 360
rect 9536 347 9543 613
rect 9716 447 9723 656
rect 9716 396 9723 433
rect 9776 410 9783 473
rect 9296 207 9303 273
rect 9576 176 9583 393
rect 9736 327 9743 363
rect 9816 327 9823 453
rect 9896 327 9903 773
rect 10036 696 10043 813
rect 10216 787 10223 876
rect 9936 367 9943 633
rect 9996 410 10003 513
rect 10016 467 10023 663
rect 10056 643 10063 663
rect 10036 636 10063 643
rect 10036 487 10043 636
rect 10036 396 10043 473
rect 9816 176 9823 313
rect 9616 147 9623 176
rect 9956 147 9963 396
rect 10076 176 10083 313
rect 10096 287 10103 393
rect 10116 187 10123 213
rect 8776 107 8783 143
rect 9036 140 9043 143
rect 9033 127 9047 140
rect 10136 143 10143 173
rect 10196 147 10203 613
rect 10236 567 10243 733
rect 10296 696 10303 1053
rect 10336 827 10343 1216
rect 10356 1127 10363 1613
rect 10436 1400 10443 1403
rect 10396 1267 10403 1390
rect 10433 1387 10447 1400
rect 10436 1287 10443 1373
rect 10476 1327 10483 1816
rect 10436 1216 10443 1252
rect 10496 1187 10503 2013
rect 10516 1847 10523 2373
rect 10536 2207 10543 2313
rect 10556 2270 10563 3093
rect 10576 2247 10583 2853
rect 10596 2747 10603 3212
rect 10676 3187 10683 3373
rect 10696 3264 10703 3513
rect 10716 3484 10723 3613
rect 10616 2964 10623 3173
rect 10736 3027 10743 4033
rect 10756 3947 10763 4213
rect 10756 3427 10763 3933
rect 10776 3847 10783 4773
rect 10816 4747 10823 5293
rect 10836 4827 10843 5273
rect 10956 5187 10963 6070
rect 10976 5803 10983 6936
rect 10996 6147 11003 6733
rect 11016 6384 11023 6633
rect 11076 6447 11083 6653
rect 10996 5827 11003 6133
rect 11016 6027 11023 6153
rect 10976 5796 11003 5803
rect 10956 5087 10963 5113
rect 10916 4987 10923 5043
rect 10916 4824 10923 4853
rect 10916 4627 10923 4753
rect 10936 4747 10943 5013
rect 10956 4767 10963 4873
rect 10796 4047 10803 4573
rect 10916 4556 10963 4563
rect 10816 4167 10823 4556
rect 10956 4524 10963 4556
rect 10836 4487 10843 4513
rect 10856 4407 10863 4523
rect 10896 4487 10903 4523
rect 10856 4347 10863 4393
rect 10956 4387 10963 4510
rect 10956 4267 10963 4336
rect 10816 4127 10823 4153
rect 10836 4036 10843 4073
rect 10796 3996 10823 4003
rect 10776 3487 10783 3673
rect 10796 3407 10803 3996
rect 10856 3927 10863 4003
rect 10856 3816 10863 3873
rect 10916 3867 10923 4033
rect 10876 3747 10883 3783
rect 10936 3767 10943 3813
rect 10876 3516 10883 3712
rect 10916 3567 10923 3733
rect 10956 3527 10963 4153
rect 10976 3647 10983 5613
rect 10996 5343 11003 5796
rect 11016 5610 11023 5933
rect 11036 5627 11043 6413
rect 11056 6147 11063 6173
rect 11076 6116 11083 6433
rect 11096 6427 11103 6973
rect 11136 6747 11143 7453
rect 11256 7183 11263 7423
rect 11236 7176 11263 7183
rect 11236 7156 11243 7176
rect 11156 7087 11163 7156
rect 11296 7123 11303 7593
rect 11316 7427 11323 7853
rect 11376 7683 11383 8233
rect 11416 8196 11423 8253
rect 11516 8247 11523 8670
rect 11453 8200 11467 8213
rect 11456 8196 11463 8200
rect 11496 7987 11503 8213
rect 11516 8003 11523 8053
rect 11536 8027 11543 8493
rect 11516 7996 11543 8003
rect 11536 7976 11543 7996
rect 11556 7987 11563 8233
rect 11576 8147 11583 8716
rect 11596 8210 11603 8773
rect 11356 7676 11383 7683
rect 11456 7676 11463 7973
rect 11476 7683 11483 7973
rect 11576 7967 11583 8133
rect 11516 7767 11523 7930
rect 11476 7676 11503 7683
rect 11256 7116 11303 7123
rect 11156 6636 11163 6673
rect 11136 6583 11143 6603
rect 11136 6576 11163 6583
rect 11116 6416 11123 6513
rect 11156 6430 11163 6576
rect 11136 6247 11143 6383
rect 11156 6130 11163 6333
rect 11196 6127 11203 6433
rect 11096 6047 11103 6083
rect 11027 5596 11043 5603
rect 11096 5607 11103 6033
rect 11056 5527 11063 5563
rect 11033 5390 11047 5393
rect 11073 5380 11087 5393
rect 11096 5387 11103 5550
rect 11076 5376 11083 5380
rect 10996 5336 11023 5343
rect 10996 5090 11003 5133
rect 11016 5027 11023 5336
rect 11116 5343 11123 5973
rect 11196 5947 11203 6092
rect 11216 5907 11223 6733
rect 11236 6447 11243 6953
rect 11176 5807 11183 5863
rect 11096 5336 11123 5343
rect 11036 4967 11043 5273
rect 11056 5027 11063 5173
rect 11036 4856 11043 4893
rect 11076 4867 11083 5093
rect 10996 3767 11003 4813
rect 11096 4823 11103 5336
rect 11136 5107 11143 5593
rect 11156 5507 11163 5596
rect 11156 5287 11163 5393
rect 11196 5347 11203 5833
rect 11216 5090 11223 5733
rect 11127 5083 11140 5087
rect 11127 5076 11143 5083
rect 11127 5073 11140 5076
rect 11236 5047 11243 6412
rect 11256 5847 11263 7073
rect 11316 6936 11323 6993
rect 11336 6967 11343 7673
rect 11356 6943 11363 7676
rect 11476 7456 11483 7613
rect 11496 7607 11503 7676
rect 11516 7456 11523 7513
rect 11356 6936 11383 6943
rect 11336 6867 11343 6903
rect 11276 6047 11283 6673
rect 11296 6604 11303 6753
rect 11356 6604 11363 6633
rect 11376 6451 11383 6936
rect 11396 6727 11403 7153
rect 11396 6647 11403 6713
rect 11416 6687 11423 7413
rect 11496 7047 11503 7123
rect 11456 6767 11463 6933
rect 11296 5707 11303 6113
rect 11276 5596 11283 5673
rect 11316 5647 11323 6433
rect 11436 6417 11443 6513
rect 11476 6467 11483 6953
rect 11476 6380 11483 6383
rect 11473 6367 11487 6380
rect 11516 6187 11523 7013
rect 11556 6967 11563 7673
rect 11576 7027 11583 7713
rect 11596 6967 11603 8013
rect 11616 7627 11623 9913
rect 11636 9807 11643 10516
rect 11696 10367 11703 10530
rect 11636 9127 11643 9772
rect 11656 9367 11663 10173
rect 11676 10167 11683 10243
rect 11676 9947 11683 10153
rect 11696 10024 11703 10213
rect 11756 10056 11763 10513
rect 11776 10447 11783 10773
rect 11796 10647 11803 10796
rect 11796 10087 11803 10576
rect 11816 10187 11823 10733
rect 11836 10247 11843 11013
rect 11896 10760 11903 10763
rect 11936 10760 11943 10763
rect 11893 10747 11907 10760
rect 11933 10747 11947 10760
rect 11976 10576 11983 11570
rect 11996 10707 12003 11253
rect 12016 10544 12023 11313
rect 11916 10447 11923 10543
rect 11953 10527 11967 10530
rect 11956 10290 11963 10473
rect 11793 10060 11807 10073
rect 11796 10056 11803 10060
rect 11776 9907 11783 10023
rect 11816 10020 11823 10023
rect 11813 10007 11827 10020
rect 11693 9760 11707 9773
rect 11696 9756 11703 9760
rect 11756 9587 11763 9653
rect 11756 9536 11763 9573
rect 11736 9367 11743 9503
rect 11796 9387 11803 9756
rect 11676 9204 11683 9273
rect 11773 9240 11787 9253
rect 11776 9236 11783 9240
rect 11716 9107 11723 9203
rect 11656 8984 11663 9033
rect 11636 8227 11643 8593
rect 11676 8567 11683 9093
rect 11716 9016 11723 9053
rect 11816 9030 11823 9273
rect 11836 9227 11843 9253
rect 11756 8716 11763 8813
rect 11793 8720 11807 8733
rect 11796 8716 11803 8720
rect 11656 8367 11663 8513
rect 11696 8460 11703 8463
rect 11736 8460 11743 8463
rect 11693 8447 11707 8460
rect 11733 8447 11747 8460
rect 11776 8447 11783 8683
rect 11656 7907 11663 8193
rect 11696 8160 11703 8163
rect 11676 8107 11683 8153
rect 11693 8147 11707 8160
rect 11796 8027 11803 8493
rect 11676 7947 11683 7976
rect 11816 7983 11823 8553
rect 11836 8127 11843 8496
rect 11816 7976 11843 7983
rect 11696 7707 11703 7973
rect 11756 7907 11763 7943
rect 11796 7787 11803 7943
rect 11776 7776 11793 7783
rect 11776 7644 11783 7776
rect 11836 7703 11843 7976
rect 11816 7696 11843 7703
rect 11653 7627 11667 7630
rect 11756 7456 11763 7593
rect 11796 7527 11803 7693
rect 11816 7587 11823 7696
rect 11796 7456 11803 7513
rect 11616 6947 11623 7153
rect 11636 7124 11643 7373
rect 11536 6384 11543 6853
rect 11596 6807 11603 6903
rect 11636 6647 11643 6953
rect 11676 6867 11683 7333
rect 11716 7156 11723 7253
rect 11756 7170 11763 7393
rect 11776 7183 11783 7423
rect 11776 7176 11803 7183
rect 11796 7156 11803 7176
rect 11736 6887 11743 7123
rect 11773 7107 11787 7110
rect 11680 6663 11693 6667
rect 11676 6653 11693 6663
rect 11676 6636 11683 6653
rect 11356 6130 11363 6173
rect 11420 6123 11433 6127
rect 11416 6116 11433 6123
rect 11420 6113 11433 6116
rect 11336 5747 11343 6073
rect 11396 6047 11403 6083
rect 11416 5896 11423 5933
rect 11456 5896 11463 6073
rect 11476 6047 11483 6153
rect 11293 5380 11307 5393
rect 11316 5387 11323 5533
rect 11296 5376 11303 5380
rect 10756 3027 10763 3213
rect 10776 3207 10783 3353
rect 10816 3296 10823 3513
rect 10836 3423 10843 3473
rect 10856 3447 10863 3483
rect 10976 3447 10983 3633
rect 10836 3416 10863 3423
rect 10856 3296 10863 3416
rect 10696 2927 10703 2963
rect 10696 2887 10703 2913
rect 10736 2867 10743 2992
rect 10656 2607 10663 2743
rect 10656 2476 10663 2513
rect 10716 2507 10723 2813
rect 10736 2790 10743 2853
rect 10693 2490 10707 2493
rect 10636 2407 10643 2443
rect 10536 1987 10543 2033
rect 10596 1956 10603 2293
rect 10616 2207 10623 2353
rect 10633 2307 10647 2313
rect 10736 2287 10743 2733
rect 10636 1956 10643 2113
rect 10656 1967 10663 2223
rect 10607 1903 10620 1907
rect 10607 1893 10613 1903
rect 10576 1736 10583 1833
rect 10616 1736 10623 1773
rect 10556 1667 10563 1703
rect 10596 1547 10603 1690
rect 10376 987 10383 1173
rect 10356 887 10363 953
rect 10216 364 10223 473
rect 10256 396 10263 650
rect 10276 527 10283 663
rect 10376 467 10383 973
rect 10476 916 10483 973
rect 10396 667 10403 916
rect 10496 664 10503 853
rect 10556 696 10563 1533
rect 10676 1436 10683 2193
rect 10696 1707 10703 1993
rect 10696 1400 10703 1403
rect 10576 1267 10583 1373
rect 10656 1367 10663 1390
rect 10693 1387 10707 1400
rect 10576 887 10583 1253
rect 10696 1216 10703 1253
rect 10696 916 10703 1113
rect 10736 1087 10743 2173
rect 10756 1750 10763 3013
rect 10716 847 10723 883
rect 10616 687 10623 793
rect 10756 667 10763 1736
rect 10776 707 10783 3013
rect 10796 3010 10803 3113
rect 10796 2490 10803 2996
rect 10816 2827 10823 3233
rect 10876 3207 10883 3263
rect 10816 2527 10823 2593
rect 10796 2187 10803 2476
rect 10816 2147 10823 2513
rect 10836 2407 10843 3173
rect 10896 2790 10903 3153
rect 10996 3127 11003 3553
rect 10996 2996 11003 3053
rect 11016 3007 11023 4453
rect 11036 3787 11043 4733
rect 11056 4427 11063 4823
rect 11076 4816 11103 4823
rect 10936 2776 10943 2893
rect 10976 2827 10983 2963
rect 10976 2744 10983 2813
rect 10876 2707 10883 2743
rect 10916 2667 10923 2743
rect 10836 2224 10843 2293
rect 10856 2107 10863 2613
rect 10896 2444 10903 2493
rect 10956 2476 10963 2573
rect 10996 2547 11003 2776
rect 10976 2423 10983 2443
rect 10956 2416 10983 2423
rect 10796 1867 10803 2073
rect 10816 1969 10823 2013
rect 10876 2007 10883 2273
rect 10916 2256 10923 2333
rect 10956 2307 10963 2416
rect 10856 1976 10893 1983
rect 10856 1963 10863 1976
rect 10836 1956 10863 1963
rect 10836 1924 10843 1956
rect 10933 1960 10947 1973
rect 10936 1956 10943 1960
rect 10867 1924 10880 1927
rect 10867 1917 10883 1924
rect 10916 1920 10923 1923
rect 10867 1913 10880 1917
rect 10913 1907 10927 1920
rect 10796 1707 10803 1773
rect 10856 1736 10863 1892
rect 10876 1700 10883 1703
rect 10873 1687 10887 1700
rect 10936 1587 10943 1753
rect 10796 1387 10803 1513
rect 10936 1436 10943 1573
rect 10976 1527 10983 2393
rect 10996 2087 11003 2373
rect 11036 2283 11043 3513
rect 11016 2276 11043 2283
rect 10996 1887 11003 1973
rect 10807 953 10813 967
rect 10856 887 10863 1353
rect 10876 1267 10883 1373
rect 10916 1367 10923 1403
rect 10956 1400 10963 1403
rect 10953 1387 10967 1400
rect 10876 1147 10883 1253
rect 10956 1216 10963 1253
rect 10996 1167 11003 1673
rect 10907 953 10913 967
rect 10956 916 10963 1073
rect 10816 696 10823 753
rect 10936 727 10943 883
rect 10376 364 10383 453
rect 10496 396 10503 650
rect 10536 627 10543 663
rect 10796 407 10803 663
rect 10836 647 10843 663
rect 10807 396 10823 403
rect 10816 364 10823 396
rect 10476 360 10483 363
rect 10273 347 10287 350
rect 10473 347 10487 360
rect 10296 190 10303 313
rect 10336 176 10343 233
rect 10396 156 10403 333
rect 10736 327 10743 363
rect 10836 327 10843 633
rect 10096 136 10143 143
rect 9293 127 9307 130
rect 10496 67 10503 156
rect 10856 67 10863 153
rect 10876 124 10883 573
rect 10896 207 10903 693
rect 10936 647 10943 713
rect 10996 647 11003 676
rect 11016 587 11023 2276
rect 11036 2227 11043 2256
rect 10956 127 10963 573
rect 11016 410 11023 552
rect 11036 403 11043 1953
rect 11056 1687 11063 3990
rect 11076 2307 11083 4816
rect 11096 4507 11103 4653
rect 11116 4447 11123 4853
rect 11136 4687 11143 5013
rect 11156 5007 11163 5043
rect 11256 5023 11263 5333
rect 11276 5307 11283 5343
rect 11336 5340 11343 5343
rect 11276 5067 11283 5293
rect 11316 5287 11323 5333
rect 11333 5327 11347 5340
rect 11296 5047 11303 5213
rect 11236 5016 11263 5023
rect 11156 4827 11163 4953
rect 11176 4556 11183 4693
rect 11216 4570 11223 4933
rect 11236 4567 11243 5016
rect 11146 4513 11147 4520
rect 11133 4503 11147 4513
rect 11196 4520 11203 4523
rect 11193 4507 11207 4520
rect 11133 4500 11163 4503
rect 11136 4496 11163 4500
rect 11156 4336 11163 4496
rect 11196 4336 11203 4373
rect 11156 4036 11163 4273
rect 11176 4227 11183 4303
rect 11236 4287 11243 4513
rect 11216 4050 11223 4233
rect 11136 3947 11143 4003
rect 11216 3887 11223 3933
rect 11136 3816 11143 3853
rect 11116 3780 11123 3783
rect 11096 3387 11103 3773
rect 11113 3767 11127 3780
rect 11156 3567 11163 3783
rect 11116 3527 11123 3553
rect 11196 3516 11203 3673
rect 11216 3527 11223 3873
rect 11136 3296 11143 3433
rect 11176 3387 11183 3483
rect 11156 3227 11163 3263
rect 11196 3260 11203 3263
rect 11193 3247 11207 3260
rect 11093 3147 11107 3153
rect 11076 1367 11083 2293
rect 11096 1807 11103 2993
rect 11116 1967 11123 3033
rect 11136 2927 11143 3093
rect 11156 2867 11163 2996
rect 11176 2967 11183 3233
rect 11196 3187 11203 3212
rect 11236 3047 11243 3873
rect 11256 3447 11263 4993
rect 11316 4867 11323 5273
rect 11336 4857 11343 5053
rect 11356 4887 11363 5073
rect 11376 4867 11383 5893
rect 11476 5807 11483 5863
rect 11396 5027 11403 5493
rect 11416 5087 11423 5633
rect 11456 5076 11463 5173
rect 11496 5110 11503 5673
rect 11516 5647 11523 6133
rect 11536 5864 11543 6113
rect 11556 6084 11563 6633
rect 11596 6604 11603 6633
rect 11696 6507 11703 6603
rect 11596 6407 11603 6493
rect 11756 6467 11763 6973
rect 11836 6970 11843 7673
rect 11856 6987 11863 10053
rect 11876 9727 11883 10230
rect 11936 10167 11943 10243
rect 11976 9907 11983 10230
rect 12016 9843 12023 10273
rect 12036 10067 12043 11353
rect 12076 11247 12083 12136
rect 12096 11804 12103 11893
rect 12153 11840 12167 11853
rect 12156 11836 12163 11840
rect 12176 11767 12183 11803
rect 12256 11707 12263 12103
rect 12156 11367 12163 11583
rect 12136 11280 12143 11283
rect 12133 11267 12147 11280
rect 12056 10747 12063 10796
rect 12076 10667 12083 11050
rect 12116 11027 12123 11063
rect 12176 10987 12183 11283
rect 12096 10747 12103 10973
rect 12156 10760 12163 10763
rect 12153 10747 12167 10760
rect 12076 10327 12083 10653
rect 12096 10147 12103 10733
rect 12196 10687 12203 10763
rect 12136 10247 12143 10276
rect 12056 10056 12063 10093
rect 12096 10056 12103 10133
rect 12076 10020 12083 10023
rect 12073 10007 12087 10020
rect 12016 9836 12043 9843
rect 11876 7727 11883 9013
rect 11896 7683 11903 9833
rect 11916 8707 11923 9793
rect 11996 9756 12003 9793
rect 12036 9563 12043 9836
rect 12016 9556 12043 9563
rect 12016 9550 12023 9556
rect 12056 9536 12063 9753
rect 12076 9727 12083 9893
rect 11956 9504 11963 9533
rect 12036 9287 12043 9503
rect 11976 9016 11983 9053
rect 12036 8987 12043 9053
rect 11936 8687 11943 8970
rect 12016 8716 12023 8853
rect 11936 8607 11943 8673
rect 12056 8464 12063 8513
rect 12016 8163 12023 8450
rect 12076 8427 12083 8495
rect 12076 8164 12083 8193
rect 11936 8127 11943 8163
rect 11976 8156 12023 8163
rect 12016 7976 12023 8013
rect 11876 7676 11903 7683
rect 11916 7676 11923 7713
rect 11876 6970 11883 7676
rect 11936 7640 11943 7643
rect 11933 7627 11947 7640
rect 12036 7547 12043 7943
rect 11936 7107 11943 7473
rect 11576 5847 11583 6113
rect 11596 5687 11603 6173
rect 11616 6127 11623 6453
rect 11776 6427 11783 6953
rect 11636 6116 11643 6153
rect 11656 6147 11663 6413
rect 11756 6380 11763 6383
rect 11753 6367 11767 6380
rect 11616 5787 11623 6033
rect 11696 6007 11703 6083
rect 11636 5807 11643 5933
rect 11656 5907 11663 5993
rect 11696 5896 11703 5953
rect 11756 5927 11763 6233
rect 11776 6047 11783 6373
rect 11676 5707 11683 5863
rect 11716 5860 11723 5863
rect 11713 5847 11727 5860
rect 11636 5596 11643 5633
rect 11516 5083 11523 5593
rect 11616 5527 11623 5550
rect 11636 5377 11643 5513
rect 11676 5487 11683 5633
rect 11696 5527 11703 5833
rect 11536 5303 11543 5377
rect 11716 5347 11723 5773
rect 11616 5340 11623 5343
rect 11613 5327 11627 5340
rect 11536 5296 11563 5303
rect 11516 5076 11543 5083
rect 11427 5043 11440 5047
rect 11427 5036 11443 5043
rect 11427 5033 11440 5036
rect 11396 4857 11403 4893
rect 11276 4527 11283 4813
rect 11336 4816 11363 4823
rect 11336 4767 11343 4816
rect 11436 4807 11443 5013
rect 11476 4987 11483 5043
rect 11276 4304 11283 4333
rect 11296 4247 11303 4373
rect 11276 4050 11283 4113
rect 11276 3247 11283 4036
rect 11296 3264 11303 4212
rect 11316 3887 11323 4433
rect 11336 3863 11343 4573
rect 11316 3856 11343 3863
rect 11316 3303 11323 3856
rect 11356 3843 11363 4793
rect 11376 3947 11383 4673
rect 11436 4556 11443 4613
rect 11456 4587 11463 4873
rect 11496 4787 11503 4873
rect 11516 4827 11523 5033
rect 11416 4387 11423 4523
rect 11456 4520 11463 4523
rect 11453 4507 11467 4520
rect 11496 4443 11503 4513
rect 11516 4467 11523 4792
rect 11496 4436 11523 4443
rect 11476 4336 11483 4393
rect 11416 4247 11423 4303
rect 11396 4007 11403 4133
rect 11436 4036 11443 4233
rect 11456 4087 11463 4303
rect 11476 4050 11483 4273
rect 11496 4207 11503 4293
rect 11516 4147 11523 4436
rect 11336 3836 11363 3843
rect 11336 3727 11343 3836
rect 11396 3816 11403 3953
rect 11336 3467 11343 3493
rect 11376 3487 11383 3783
rect 11416 3780 11423 3783
rect 11413 3767 11427 3780
rect 11476 3767 11483 3933
rect 11416 3516 11423 3553
rect 11316 3296 11343 3303
rect 11416 3296 11423 3453
rect 11256 3010 11263 3233
rect 11276 3027 11283 3133
rect 11236 2947 11243 2963
rect 11236 2936 11253 2947
rect 11240 2933 11253 2936
rect 11236 2867 11243 2913
rect 11236 2776 11243 2853
rect 11136 2587 11143 2773
rect 11216 2707 11223 2743
rect 11136 2387 11143 2533
rect 11216 2476 11223 2573
rect 11276 2567 11283 2953
rect 11296 2807 11303 3250
rect 11316 2607 11323 3273
rect 11176 2343 11183 2473
rect 11236 2427 11243 2443
rect 11176 2336 11203 2343
rect 11196 2256 11203 2336
rect 11176 2163 11183 2223
rect 11236 2207 11243 2413
rect 11156 2156 11183 2163
rect 11156 2027 11163 2156
rect 11176 1956 11183 2133
rect 11136 1767 11143 1923
rect 11153 1743 11167 1753
rect 11136 1740 11167 1743
rect 11136 1736 11163 1740
rect 11176 1667 11183 1733
rect 11216 1687 11223 2153
rect 11236 1767 11243 1953
rect 11216 1436 11223 1652
rect 11076 767 11083 1216
rect 11136 1187 11143 1413
rect 11176 1307 11183 1403
rect 11173 1230 11187 1233
rect 11216 1216 11223 1313
rect 11216 1107 11223 1133
rect 11216 916 11223 1093
rect 11256 927 11263 2353
rect 11276 1823 11283 2253
rect 11316 2127 11323 2553
rect 11336 2267 11343 3296
rect 11356 2627 11363 3113
rect 11376 2927 11383 3253
rect 11396 3207 11403 3263
rect 11396 3067 11403 3193
rect 11436 3067 11443 3263
rect 11476 3227 11483 3473
rect 11496 3447 11503 4003
rect 11516 3607 11523 3753
rect 11496 3407 11503 3433
rect 11516 3267 11523 3593
rect 11296 1924 11303 2093
rect 11276 1816 11303 1823
rect 11076 696 11083 753
rect 11113 700 11127 713
rect 11116 696 11123 700
rect 11036 396 11063 403
rect 10996 247 11003 350
rect 11033 327 11047 333
rect 11056 176 11063 396
rect 11096 176 11103 293
rect 11136 144 11143 393
rect 11156 190 11163 913
rect 11176 327 11183 813
rect 11196 727 11203 883
rect 11236 880 11243 883
rect 11233 867 11247 880
rect 11233 847 11247 853
rect 11236 447 11243 713
rect 11256 664 11263 773
rect 11196 144 11203 413
rect 11256 396 11263 650
rect 11276 487 11283 1793
rect 11296 427 11303 1816
rect 11336 1807 11343 2232
rect 11356 2167 11363 2533
rect 11376 2224 11383 2273
rect 11396 2167 11403 3053
rect 11467 3023 11480 3027
rect 11467 3013 11483 3023
rect 11476 2996 11483 3013
rect 11536 3003 11543 5076
rect 11556 5047 11563 5296
rect 11556 4467 11563 4853
rect 11556 4167 11563 4432
rect 11576 4287 11583 4973
rect 11596 4947 11603 5076
rect 11636 4947 11643 5133
rect 11656 4890 11663 5093
rect 11696 5090 11703 5153
rect 11736 5127 11743 5693
rect 11756 5547 11763 5853
rect 11776 5727 11783 5953
rect 11756 5103 11763 5393
rect 11736 5096 11763 5103
rect 11736 5090 11743 5096
rect 11776 5087 11783 5593
rect 11613 4860 11627 4873
rect 11616 4856 11623 4860
rect 11556 3027 11563 4073
rect 11596 3883 11603 4453
rect 11616 3947 11623 4413
rect 11636 4287 11643 4510
rect 11656 4427 11663 4673
rect 11696 4563 11703 4873
rect 11716 4787 11723 5043
rect 11756 4587 11763 4953
rect 11676 4556 11703 4563
rect 11776 4567 11783 5033
rect 11676 4467 11683 4556
rect 11756 4407 11763 4523
rect 11656 3887 11663 4193
rect 11696 4047 11703 4293
rect 11716 4247 11723 4303
rect 11736 4036 11743 4273
rect 11756 4207 11763 4372
rect 11776 4087 11783 4453
rect 11576 3876 11603 3883
rect 11536 2996 11563 3003
rect 11416 2947 11423 2996
rect 11476 2776 11483 2913
rect 11496 2907 11503 2963
rect 11536 2743 11543 2793
rect 11456 2490 11463 2743
rect 11496 2707 11503 2743
rect 11516 2736 11543 2743
rect 11496 2527 11503 2693
rect 11516 2476 11523 2736
rect 11456 2427 11463 2476
rect 11496 2347 11503 2443
rect 11496 2256 11503 2293
rect 11556 2283 11563 2996
rect 11576 2947 11583 3876
rect 11596 3787 11603 3853
rect 11676 3816 11683 4013
rect 11716 3967 11723 4003
rect 11756 3996 11773 4003
rect 11596 3530 11603 3752
rect 11596 3107 11603 3516
rect 11616 3487 11623 3713
rect 11636 3487 11643 3733
rect 11656 3727 11663 3783
rect 11736 3747 11743 3913
rect 11756 3727 11763 3873
rect 11616 3243 11623 3452
rect 11656 3303 11663 3513
rect 11676 3347 11683 3713
rect 11696 3527 11703 3713
rect 11716 3516 11723 3633
rect 11776 3587 11783 3990
rect 11796 3647 11803 6935
rect 11816 3607 11823 6793
rect 11836 5563 11843 6873
rect 11856 6683 11863 6903
rect 11856 6676 11883 6683
rect 11856 5607 11863 6653
rect 11876 6647 11883 6676
rect 11896 6636 11903 6833
rect 11916 6667 11923 6953
rect 11956 6747 11963 7533
rect 12033 7460 12047 7473
rect 12076 7467 12083 7753
rect 12036 7456 12043 7460
rect 11996 7420 12003 7423
rect 11993 7407 12007 7420
rect 11976 6807 11983 7153
rect 11996 7023 12003 7313
rect 12036 7156 12043 7373
rect 12056 7347 12063 7423
rect 12096 7327 12103 9236
rect 12116 8730 12123 9533
rect 12116 8684 12123 8716
rect 12136 8663 12143 10173
rect 12156 9727 12163 10633
rect 12216 10576 12223 10713
rect 12256 10647 12263 11570
rect 12276 10727 12283 10796
rect 12196 10487 12203 10543
rect 12216 10276 12223 10313
rect 12196 10240 12203 10243
rect 12193 10227 12207 10240
rect 12236 9847 12243 10243
rect 12156 8987 12163 9233
rect 12116 8656 12143 8663
rect 12116 7567 12123 8656
rect 12136 7647 12143 8613
rect 12116 7387 12123 7453
rect 12116 7156 12123 7253
rect 12056 7120 12063 7123
rect 12053 7107 12067 7120
rect 11996 7016 12023 7023
rect 11933 6640 11947 6653
rect 11936 6636 11943 6640
rect 11916 6567 11923 6603
rect 11876 6387 11883 6553
rect 11876 5867 11883 6313
rect 11896 6287 11903 6413
rect 11916 6187 11923 6453
rect 11936 6267 11943 6573
rect 11956 6467 11963 6603
rect 11976 6443 11983 6593
rect 11996 6587 12003 6936
rect 12016 6647 12023 7016
rect 12036 6587 12043 7093
rect 12096 7087 12103 7123
rect 12056 6447 12063 7072
rect 12076 6896 12103 6903
rect 12076 6847 12083 6896
rect 11976 6436 12003 6443
rect 11996 6416 12003 6436
rect 11976 6380 11983 6383
rect 11973 6367 11987 6380
rect 11913 6120 11927 6133
rect 11916 6116 11923 6120
rect 11976 6116 11983 6193
rect 11896 5843 11903 6053
rect 11936 6047 11943 6083
rect 12016 6067 12023 6383
rect 11876 5836 11903 5843
rect 11876 5667 11883 5836
rect 11916 5823 11923 5873
rect 11896 5816 11923 5823
rect 11876 5596 11883 5653
rect 11896 5647 11903 5816
rect 11916 5607 11923 5793
rect 11936 5627 11943 5993
rect 11976 5896 11983 6033
rect 12036 6007 12043 6173
rect 12056 6047 12063 6373
rect 12013 5900 12027 5913
rect 12016 5896 12023 5900
rect 11996 5767 12003 5863
rect 12036 5860 12043 5863
rect 12033 5847 12047 5860
rect 11940 5603 11953 5607
rect 11936 5596 11953 5603
rect 11940 5593 11953 5596
rect 11836 5556 11863 5563
rect 11836 5007 11843 5533
rect 11856 4983 11863 5556
rect 11976 5527 11983 5563
rect 11876 5344 11883 5433
rect 11936 5427 11943 5473
rect 11936 5376 11943 5413
rect 11976 5376 11983 5473
rect 11996 5407 12003 5553
rect 12016 5487 12023 5573
rect 12016 5327 12023 5413
rect 11836 4976 11863 4983
rect 11836 4567 11843 4976
rect 11876 4967 11883 5076
rect 11916 5044 11923 5153
rect 12036 5127 12043 5653
rect 12056 5344 12063 5613
rect 12076 5207 12083 6812
rect 12096 6487 12103 6873
rect 12156 6667 12163 8952
rect 12176 8207 12183 9013
rect 12196 8967 12203 9713
rect 12216 9667 12223 9723
rect 12296 9504 12303 11093
rect 12316 10187 12323 11616
rect 12276 9016 12283 9053
rect 12256 8963 12263 8983
rect 12236 8956 12263 8963
rect 12216 8530 12223 8713
rect 12236 8527 12243 8956
rect 12336 8627 12343 12136
rect 12253 8500 12267 8513
rect 12256 8496 12263 8500
rect 12316 8367 12323 8513
rect 12216 8196 12223 8233
rect 12196 8107 12203 8163
rect 12236 7767 12243 8150
rect 12216 7676 12223 7713
rect 12176 6827 12183 7633
rect 12196 7587 12203 7643
rect 12196 6887 12203 7552
rect 12236 6727 12243 7643
rect 12096 6327 12103 6433
rect 11936 4870 11943 5113
rect 11876 4820 11883 4823
rect 11873 4807 11887 4820
rect 11836 3663 11843 4553
rect 11856 3727 11863 4553
rect 11876 4350 11883 4772
rect 11916 4607 11923 4823
rect 11876 4267 11883 4336
rect 11876 3907 11883 4033
rect 11896 3867 11903 4573
rect 11916 4387 11923 4572
rect 11936 4567 11943 4753
rect 11956 4587 11963 5113
rect 12013 5080 12027 5093
rect 12016 5076 12023 5080
rect 11996 4947 12003 5043
rect 11976 4556 11983 4673
rect 12016 4556 12023 4853
rect 12036 4787 12043 4953
rect 12056 4827 12063 4993
rect 12096 4863 12103 6273
rect 12116 6147 12123 6413
rect 12116 6087 12123 6133
rect 12116 5327 12123 6052
rect 12076 4856 12103 4863
rect 12036 4567 12043 4653
rect 11956 4407 11963 4523
rect 11996 4336 12003 4433
rect 12056 4304 12063 4613
rect 11936 4283 11943 4303
rect 11936 4276 11963 4283
rect 11916 3987 11923 4013
rect 11936 4003 11943 4253
rect 11956 4227 11963 4276
rect 11936 3996 11963 4003
rect 11976 4000 11983 4003
rect 11956 3816 11963 3996
rect 11973 3987 11987 4000
rect 11836 3656 11863 3663
rect 11756 3516 11763 3553
rect 11796 3483 11803 3553
rect 11636 3296 11663 3303
rect 11696 3296 11703 3473
rect 11736 3383 11743 3483
rect 11716 3376 11743 3383
rect 11776 3476 11803 3483
rect 11716 3327 11723 3376
rect 11776 3367 11783 3476
rect 11736 3296 11743 3353
rect 11636 3263 11643 3296
rect 11636 3256 11663 3263
rect 11616 3236 11643 3243
rect 11636 3027 11643 3236
rect 11656 3027 11663 3256
rect 11716 3167 11723 3263
rect 11776 3247 11783 3332
rect 11576 2867 11583 2912
rect 11536 2276 11563 2283
rect 11416 2216 11443 2223
rect 11416 2187 11423 2216
rect 11356 1750 11363 1993
rect 11416 1956 11423 2173
rect 11336 1667 11343 1703
rect 11376 1687 11383 1703
rect 11336 1607 11343 1653
rect 11316 1027 11323 1513
rect 11336 1227 11343 1436
rect 11376 1427 11383 1673
rect 11416 1503 11423 1853
rect 11456 1647 11463 1793
rect 11476 1607 11483 2153
rect 11396 1496 11423 1503
rect 11376 1184 11383 1293
rect 11396 1127 11403 1496
rect 11496 1447 11503 2193
rect 11516 1507 11523 2213
rect 11476 1400 11483 1403
rect 11473 1387 11487 1400
rect 11436 1287 11443 1353
rect 11436 1216 11443 1273
rect 11473 1230 11487 1233
rect 11316 747 11323 1013
rect 11493 920 11507 933
rect 11496 916 11503 920
rect 11336 767 11343 793
rect 11356 696 11363 853
rect 11396 727 11403 916
rect 11476 676 11483 813
rect 11536 783 11543 2276
rect 11556 1007 11563 2253
rect 11596 2227 11603 2953
rect 11616 2367 11623 2933
rect 11636 2267 11643 2992
rect 11656 2623 11663 2992
rect 11676 2967 11683 3113
rect 11716 3087 11723 3153
rect 11736 3063 11743 3233
rect 11716 3056 11743 3063
rect 11696 2867 11703 3013
rect 11716 3007 11723 3056
rect 11756 2996 11763 3213
rect 11693 2780 11707 2793
rect 11696 2776 11703 2780
rect 11736 2776 11743 2950
rect 11676 2647 11683 2733
rect 11716 2667 11723 2743
rect 11656 2616 11683 2623
rect 11616 2187 11623 2253
rect 11636 2207 11643 2232
rect 11656 2223 11663 2513
rect 11676 2407 11683 2616
rect 11776 2567 11783 2853
rect 11796 2790 11803 3193
rect 11816 2907 11823 3572
rect 11716 2287 11723 2553
rect 11796 2490 11803 2593
rect 11736 2256 11743 2293
rect 11776 2267 11783 2393
rect 11656 2216 11683 2223
rect 11676 1970 11683 2216
rect 11716 2203 11723 2223
rect 11716 2196 11743 2203
rect 11736 2127 11743 2196
rect 11576 987 11583 1913
rect 11636 1736 11643 1793
rect 11696 1747 11703 1923
rect 11616 1700 11623 1703
rect 11613 1687 11627 1700
rect 11656 1687 11663 1703
rect 11716 1687 11723 1910
rect 11736 1867 11743 2113
rect 11756 2087 11763 2223
rect 11756 1907 11763 1993
rect 11596 1487 11603 1553
rect 11596 1367 11603 1473
rect 11616 1147 11623 1436
rect 11636 1404 11643 1593
rect 11656 1387 11663 1673
rect 11736 1487 11743 1736
rect 11756 1704 11763 1793
rect 11776 1447 11783 2213
rect 11796 1447 11803 2273
rect 11656 1184 11663 1273
rect 11716 1216 11723 1353
rect 11756 1227 11763 1403
rect 11796 1147 11803 1412
rect 11556 787 11563 933
rect 11636 827 11643 1113
rect 11816 1047 11823 2273
rect 11756 916 11803 923
rect 11676 867 11683 916
rect 11736 827 11743 883
rect 11796 847 11803 916
rect 11816 867 11823 973
rect 11516 776 11543 783
rect 11516 684 11523 776
rect 11796 767 11803 833
rect 11836 703 11843 3633
rect 11856 3207 11863 3656
rect 11876 3567 11883 3816
rect 11876 3487 11883 3532
rect 11856 727 11863 3172
rect 11876 707 11883 3452
rect 11896 3187 11903 3593
rect 11916 3427 11923 3753
rect 11936 3687 11943 3783
rect 11936 3467 11943 3573
rect 11956 3547 11963 3713
rect 11976 3647 11983 3783
rect 12016 3587 12023 3853
rect 12056 3767 12063 4213
rect 11976 3516 11983 3553
rect 12056 3527 12063 3633
rect 11896 2447 11903 3152
rect 11916 2287 11923 3293
rect 11936 2964 11943 3432
rect 11956 3307 11963 3473
rect 12036 3447 12043 3483
rect 11976 3296 11983 3413
rect 12056 3307 12063 3473
rect 11996 3260 12003 3263
rect 11993 3247 12007 3260
rect 12036 3207 12043 3263
rect 12016 2927 12023 2963
rect 11976 2776 11983 2833
rect 11916 2187 11923 2252
rect 11936 2167 11943 2473
rect 11956 2444 11963 2493
rect 11976 2483 11983 2633
rect 11996 2507 12003 2743
rect 12016 2527 12023 2713
rect 12056 2547 12063 3253
rect 11976 2476 12003 2483
rect 12076 2487 12083 4856
rect 12116 4847 12123 5073
rect 12136 4867 12143 6633
rect 12236 6636 12243 6673
rect 12276 6647 12283 7633
rect 12296 6687 12303 8193
rect 12156 6307 12163 6632
rect 12176 6283 12183 6593
rect 12156 6276 12183 6283
rect 12156 5343 12163 6276
rect 12196 6263 12203 6573
rect 12216 6547 12223 6603
rect 12216 6387 12223 6473
rect 12256 6427 12263 6603
rect 12276 6416 12283 6453
rect 12316 6416 12323 6713
rect 12336 6427 12343 7713
rect 12176 6256 12203 6263
rect 12176 6067 12183 6256
rect 12236 6116 12243 6353
rect 12296 6123 12303 6383
rect 12276 6116 12303 6123
rect 12176 5607 12183 6032
rect 12256 5967 12263 6083
rect 12196 5807 12203 5896
rect 12256 5860 12263 5863
rect 12253 5847 12267 5860
rect 12256 5596 12263 5753
rect 12216 5527 12223 5553
rect 12276 5387 12283 5550
rect 12156 5336 12183 5343
rect 12196 5340 12203 5343
rect 12156 4967 12163 5313
rect 12176 5247 12183 5336
rect 12193 5327 12207 5340
rect 12196 4856 12203 5076
rect 12216 5047 12223 5333
rect 12256 5263 12263 5343
rect 12276 5287 12283 5333
rect 12296 5263 12303 5513
rect 12256 5256 12303 5263
rect 12096 4267 12103 4833
rect 12116 4327 12123 4812
rect 12116 4243 12123 4313
rect 12136 4283 12143 4813
rect 12156 4307 12163 4673
rect 12136 4276 12163 4283
rect 12096 4236 12123 4243
rect 12096 3727 12103 4236
rect 12136 4223 12143 4253
rect 12116 4216 12143 4223
rect 12096 2847 12103 3673
rect 12096 2744 12103 2812
rect 11976 2256 11983 2293
rect 12016 2290 12023 2430
rect 12036 2267 12043 2413
rect 12056 2403 12063 2443
rect 12056 2396 12083 2403
rect 11973 1960 11987 1973
rect 11976 1956 11983 1960
rect 11936 1920 11943 1923
rect 11933 1907 11947 1920
rect 11916 1736 11923 1773
rect 11953 1740 11967 1753
rect 12016 1750 12023 1953
rect 11956 1736 11963 1740
rect 11936 1687 11943 1703
rect 11896 747 11903 1453
rect 11916 1287 11923 1633
rect 11936 1547 11943 1673
rect 12016 1436 12023 1533
rect 12036 1467 12043 1973
rect 12056 1927 12063 2373
rect 12076 2307 12083 2396
rect 12076 1987 12083 2272
rect 12096 1847 12103 2730
rect 12076 1704 12083 1753
rect 11976 1396 12003 1403
rect 11933 1220 11947 1233
rect 11936 1216 11943 1220
rect 11976 1216 11983 1396
rect 11956 1163 11963 1183
rect 12036 1184 12043 1213
rect 12076 1187 12083 1690
rect 12096 1407 12103 1833
rect 11956 1156 11983 1163
rect 11836 696 11863 703
rect 11856 683 11863 696
rect 11856 676 11883 683
rect 11336 567 11343 663
rect 11836 587 11843 643
rect 11236 327 11243 363
rect 11316 347 11323 383
rect 11376 327 11383 383
rect 11416 347 11423 433
rect 11736 416 11743 553
rect 11776 387 11783 473
rect 11796 347 11803 393
rect 11076 140 11083 143
rect 11073 127 11087 140
rect 11296 67 11303 313
rect 11336 176 11343 253
rect 11616 176 11623 273
rect 11676 144 11683 173
rect 11816 144 11823 473
rect 11876 347 11883 676
rect 11896 203 11903 712
rect 11916 367 11923 693
rect 11876 196 11903 203
rect 11876 190 11883 196
rect 11916 176 11923 332
rect 11936 183 11943 993
rect 11956 647 11963 1133
rect 11976 1027 11983 1156
rect 12016 916 12023 1173
rect 12076 884 12083 953
rect 12116 887 12123 4216
rect 12136 1987 12143 4033
rect 12156 1963 12163 4276
rect 12176 2387 12183 4773
rect 12216 4767 12223 4823
rect 12196 4247 12203 4573
rect 12216 4507 12223 4713
rect 12236 4563 12243 4813
rect 12256 4587 12263 5093
rect 12276 4827 12283 5233
rect 12296 4687 12303 5193
rect 12316 4727 12323 6253
rect 12236 4556 12263 4563
rect 12313 4560 12327 4573
rect 12336 4567 12343 6373
rect 12316 4556 12323 4560
rect 12276 4516 12303 4523
rect 12236 4336 12243 4513
rect 12276 4336 12283 4393
rect 12296 4347 12303 4516
rect 12216 4223 12223 4293
rect 12196 4216 12223 4223
rect 12196 3827 12203 4216
rect 12256 4036 12263 4233
rect 12296 4047 12303 4293
rect 12236 3927 12243 4003
rect 12276 3947 12283 4003
rect 12256 3830 12263 3873
rect 12196 3407 12203 3733
rect 12216 3567 12223 3783
rect 12296 3783 12303 3993
rect 12276 3776 12303 3783
rect 12236 3587 12243 3773
rect 12256 3563 12263 3753
rect 12236 3556 12263 3563
rect 12236 3527 12243 3556
rect 12276 3547 12283 3776
rect 12316 3767 12323 4493
rect 12336 3747 12343 4513
rect 12216 3387 12223 3516
rect 12296 3516 12303 3653
rect 12336 3527 12343 3553
rect 12233 3463 12247 3473
rect 12233 3460 12263 3463
rect 12236 3456 12263 3460
rect 12196 3207 12203 3333
rect 12236 3296 12243 3433
rect 12256 3327 12263 3456
rect 12276 3296 12283 3373
rect 12296 3347 12303 3433
rect 12316 3307 12323 3470
rect 12216 3227 12223 3253
rect 12256 3127 12263 3263
rect 12196 2827 12203 3033
rect 12253 3000 12267 3013
rect 12256 2996 12263 3000
rect 12236 2776 12243 2963
rect 12216 2740 12223 2743
rect 12213 2727 12227 2740
rect 12296 2727 12303 3193
rect 12196 2363 12203 2473
rect 12176 2356 12203 2363
rect 12176 2007 12183 2356
rect 12136 1956 12163 1963
rect 12196 1956 12203 2293
rect 12256 2256 12263 2709
rect 12236 2167 12243 2223
rect 11996 880 12003 883
rect 11993 867 12007 880
rect 11976 627 11983 673
rect 11996 447 12003 693
rect 12016 403 12023 733
rect 12076 727 12083 833
rect 12096 696 12103 773
rect 12016 396 12043 403
rect 11936 176 11963 183
rect 11396 140 11403 143
rect 11393 127 11407 140
rect 11596 107 11603 143
rect 11816 107 11823 130
rect 11896 67 11903 143
rect 11956 127 11963 176
rect 12036 107 12043 396
rect 12056 147 12063 633
rect 12136 190 12143 1956
rect 12156 307 12163 1913
rect 12176 1747 12183 1923
rect 12216 1887 12223 1923
rect 12256 1736 12263 1913
rect 12276 1847 12283 2223
rect 12176 1387 12183 1693
rect 12236 1700 12243 1703
rect 12233 1687 12247 1700
rect 12236 1436 12243 1493
rect 12176 447 12183 1273
rect 12236 1216 12243 1373
rect 12196 427 12203 1033
rect 12256 916 12263 1183
rect 12216 427 12223 873
rect 12176 367 12183 412
rect 12196 403 12203 413
rect 12196 396 12223 403
rect 12256 396 12263 433
rect 12216 107 12223 143
rect 12296 67 12303 1993
rect 12316 287 12323 3213
rect 12336 267 12343 3393
rect 7016 -24 7043 -17
rect 7516 -24 7523 13
<< m3contact >>
rect 4093 12233 4107 12247
rect 4173 12233 4187 12247
rect 2233 12213 2247 12227
rect 2453 12213 2467 12227
rect 393 12173 407 12187
rect 493 12173 507 12187
rect 233 12136 247 12150
rect 313 12136 327 12150
rect 213 12090 227 12104
rect 193 11789 207 11803
rect 413 12133 427 12147
rect 453 12136 467 12150
rect 753 12136 767 12150
rect 833 12133 847 12147
rect 993 12136 1007 12150
rect 1053 12133 1067 12147
rect 1253 12136 1267 12150
rect 1533 12136 1547 12150
rect 1573 12136 1587 12150
rect 1693 12136 1707 12150
rect 1753 12136 1767 12150
rect 1793 12136 1807 12150
rect 2033 12136 2047 12150
rect 2073 12136 2087 12150
rect 393 12093 407 12107
rect 333 11793 347 11807
rect 253 11753 267 11767
rect 313 11753 327 11767
rect 233 11673 247 11687
rect 713 12093 727 12107
rect 673 11933 687 11947
rect 513 11913 527 11927
rect 413 11873 427 11887
rect 453 11836 467 11850
rect 493 11836 507 11850
rect 533 11836 547 11850
rect 573 11836 587 11850
rect 593 11813 607 11827
rect 513 11773 527 11787
rect 573 11773 587 11787
rect 453 11753 467 11767
rect 393 11733 407 11747
rect 273 11633 287 11647
rect 333 11633 347 11647
rect 493 11616 507 11630
rect 773 12090 787 12104
rect 833 12090 847 12104
rect 733 12073 747 12087
rect 913 11913 927 11927
rect 793 11873 807 11887
rect 753 11836 767 11850
rect 913 11836 927 11850
rect 713 11790 727 11804
rect 773 11790 787 11804
rect 793 11733 807 11747
rect 673 11673 687 11687
rect 773 11673 787 11687
rect 213 11570 227 11584
rect 333 11570 347 11584
rect 213 11513 227 11527
rect 253 11513 267 11527
rect 233 11270 247 11284
rect 173 11096 187 11110
rect 233 11096 247 11110
rect 213 11050 227 11064
rect 313 10833 327 10847
rect 193 10749 207 10763
rect 233 10613 247 10627
rect 233 10576 247 10590
rect 213 10313 227 10327
rect 273 10313 287 10327
rect 313 10313 327 10327
rect 233 10276 247 10290
rect 293 10230 307 10244
rect 253 10093 267 10107
rect 233 10056 247 10070
rect 213 9973 227 9987
rect 193 9753 207 9767
rect 253 9893 267 9907
rect 293 9893 307 9907
rect 253 9756 267 9770
rect 193 9713 207 9727
rect 233 9673 247 9687
rect 193 9533 207 9547
rect 213 9490 227 9504
rect 273 9493 287 9507
rect 253 9273 267 9287
rect 213 9253 227 9267
rect 293 9233 307 9247
rect 193 9193 207 9207
rect 273 9190 287 9204
rect 193 9153 207 9167
rect 233 9153 247 9167
rect 253 9133 267 9147
rect 273 9016 287 9030
rect 313 9016 327 9030
rect 253 8970 267 8984
rect 253 8793 267 8807
rect 213 8753 227 8767
rect 293 8613 307 8627
rect 273 8553 287 8567
rect 233 8496 247 8510
rect 513 11570 527 11584
rect 593 11573 607 11587
rect 453 11413 467 11427
rect 473 11413 487 11427
rect 693 11616 707 11630
rect 753 11616 767 11630
rect 873 11673 887 11687
rect 813 11633 827 11647
rect 853 11633 867 11647
rect 693 11413 707 11427
rect 673 11373 687 11387
rect 813 11570 827 11584
rect 793 11373 807 11387
rect 553 11333 567 11347
rect 773 11333 787 11347
rect 493 11316 507 11330
rect 473 11270 487 11284
rect 473 11135 487 11149
rect 413 11053 427 11067
rect 613 11316 627 11330
rect 573 11133 587 11147
rect 613 11093 627 11107
rect 693 11096 707 11110
rect 573 10933 587 10947
rect 553 10833 567 10847
rect 493 10796 507 10810
rect 533 10796 547 10810
rect 673 10753 687 10767
rect 633 10733 647 10747
rect 553 10693 567 10707
rect 593 10693 607 10707
rect 493 10653 507 10667
rect 553 10653 567 10667
rect 473 10576 487 10590
rect 513 10576 527 10590
rect 553 10513 567 10527
rect 493 10453 507 10467
rect 453 10413 467 10427
rect 553 10413 567 10427
rect 353 10276 367 10290
rect 393 10276 407 10290
rect 513 10276 527 10290
rect 553 10276 567 10290
rect 393 10230 407 10244
rect 353 10193 367 10207
rect 353 9573 367 9587
rect 533 10193 547 10207
rect 533 10093 547 10107
rect 453 10053 467 10067
rect 493 10056 507 10070
rect 493 9993 507 10007
rect 453 9973 467 9987
rect 513 9973 527 9987
rect 433 9756 447 9770
rect 473 9756 487 9770
rect 493 9710 507 9724
rect 433 9490 447 9504
rect 393 9393 407 9407
rect 373 9236 387 9250
rect 373 9190 387 9204
rect 353 8970 367 8984
rect 353 8733 367 8747
rect 333 8633 347 8647
rect 353 8553 367 8567
rect 313 8493 327 8507
rect 213 8450 227 8464
rect 293 8453 307 8467
rect 333 8450 347 8464
rect 233 8233 247 8247
rect 273 8196 287 8210
rect 313 8196 327 8210
rect 253 8150 267 8164
rect 313 8093 327 8107
rect 273 8013 287 8027
rect 313 8013 327 8027
rect 253 7930 267 7944
rect 313 7893 327 7907
rect 213 7873 227 7887
rect 253 7713 267 7727
rect 173 7676 187 7690
rect 213 7676 227 7690
rect 273 7630 287 7644
rect 233 7593 247 7607
rect 173 7573 187 7587
rect 233 7572 247 7586
rect 253 7393 267 7407
rect 333 7630 347 7644
rect 213 7353 227 7367
rect 313 7353 327 7367
rect 213 7193 227 7207
rect 253 7156 267 7170
rect 313 7156 327 7170
rect 233 7110 247 7124
rect 233 7089 247 7103
rect 213 6853 227 6867
rect 573 9756 587 9770
rect 573 9633 587 9647
rect 553 9453 567 9467
rect 493 9273 507 9287
rect 513 9153 527 9167
rect 433 9133 447 9147
rect 513 9016 527 9030
rect 413 8973 427 8987
rect 533 8933 547 8947
rect 493 8793 507 8807
rect 433 8753 447 8767
rect 493 8733 507 8747
rect 613 10653 627 10667
rect 613 10576 627 10590
rect 693 10653 707 10667
rect 653 10573 667 10587
rect 753 11270 767 11284
rect 753 11133 767 11147
rect 753 11096 767 11110
rect 793 11096 807 11110
rect 773 11050 787 11064
rect 833 10973 847 10987
rect 893 11613 907 11627
rect 913 11570 927 11584
rect 1233 12090 1247 12104
rect 1053 12073 1067 12087
rect 1193 11853 1207 11867
rect 1053 11836 1067 11850
rect 1093 11836 1107 11850
rect 1173 11836 1187 11850
rect 1013 11793 1027 11807
rect 1073 11790 1087 11804
rect 1113 11753 1127 11767
rect 1353 12090 1367 12104
rect 1413 11853 1427 11867
rect 2113 12133 2127 12147
rect 2153 12133 2167 12147
rect 1733 12073 1747 12087
rect 1793 12073 1807 12087
rect 1693 12033 1707 12047
rect 1733 12033 1747 12047
rect 1633 11873 1647 11887
rect 1673 11836 1687 11850
rect 1273 11773 1287 11787
rect 1513 11790 1527 11804
rect 1693 11790 1707 11804
rect 1193 11753 1207 11767
rect 1333 11753 1347 11767
rect 1393 11753 1407 11767
rect 1113 11633 1127 11647
rect 1153 11633 1167 11647
rect 1073 11616 1087 11630
rect 1053 11570 1067 11584
rect 1153 11573 1167 11587
rect 973 11493 987 11507
rect 1093 11493 1107 11507
rect 933 11413 947 11427
rect 873 11270 887 11284
rect 913 11273 927 11287
rect 813 10813 827 10827
rect 853 10813 867 10827
rect 833 10750 847 10764
rect 893 10693 907 10707
rect 1033 11333 1047 11347
rect 993 11316 1007 11330
rect 1073 11316 1087 11330
rect 1013 11270 1027 11284
rect 1313 11693 1327 11707
rect 1193 11616 1207 11630
rect 1353 11616 1367 11630
rect 1333 11570 1347 11584
rect 1313 11373 1327 11387
rect 1193 11333 1207 11347
rect 1073 11233 1087 11247
rect 1173 11233 1187 11247
rect 973 11213 987 11227
rect 1033 11153 1047 11167
rect 1153 11153 1167 11167
rect 1073 11096 1087 11110
rect 1113 11096 1127 11110
rect 973 11053 987 11067
rect 1053 10993 1067 11007
rect 1153 11050 1167 11064
rect 1073 10973 1087 10987
rect 1113 10973 1127 10987
rect 1073 10813 1087 10827
rect 1093 10693 1107 10707
rect 1013 10653 1027 10667
rect 773 10613 787 10627
rect 933 10613 947 10627
rect 733 10576 747 10590
rect 853 10576 867 10590
rect 993 10576 1007 10590
rect 633 10193 647 10207
rect 613 9893 627 9907
rect 693 10530 707 10544
rect 793 10530 807 10544
rect 1013 10513 1027 10527
rect 973 10453 987 10467
rect 753 10393 767 10407
rect 853 10393 867 10407
rect 773 10313 787 10327
rect 933 10276 947 10290
rect 793 10230 807 10244
rect 853 10233 867 10247
rect 753 10193 767 10207
rect 753 10093 767 10107
rect 693 9833 707 9847
rect 893 10010 907 10024
rect 733 9756 747 9770
rect 773 9756 787 9770
rect 873 9753 887 9767
rect 693 9713 707 9727
rect 733 9693 747 9707
rect 653 9573 667 9587
rect 753 9633 767 9647
rect 653 9536 667 9550
rect 693 9536 707 9550
rect 733 9536 747 9550
rect 833 9533 847 9547
rect 873 9536 887 9550
rect 653 9493 667 9507
rect 673 9453 687 9467
rect 673 9253 687 9267
rect 673 9193 687 9207
rect 673 8933 687 8947
rect 593 8793 607 8807
rect 433 8673 447 8687
rect 833 9473 847 9487
rect 753 9453 767 9467
rect 773 9293 787 9307
rect 733 9236 747 9250
rect 753 9190 767 9204
rect 833 9193 847 9207
rect 833 9153 847 9167
rect 793 9073 807 9087
rect 753 9016 767 9030
rect 833 9033 847 9047
rect 733 8933 747 8947
rect 833 8933 847 8947
rect 773 8873 787 8887
rect 693 8833 707 8847
rect 773 8833 787 8847
rect 733 8733 747 8747
rect 813 8793 827 8807
rect 513 8670 527 8684
rect 673 8670 687 8684
rect 753 8670 767 8684
rect 753 8633 767 8647
rect 433 8496 447 8510
rect 473 8496 487 8510
rect 793 8613 807 8627
rect 853 8593 867 8607
rect 793 8533 807 8547
rect 453 8450 467 8464
rect 693 8450 707 8464
rect 733 8450 747 8464
rect 493 8433 507 8447
rect 653 8433 667 8447
rect 593 8313 607 8327
rect 633 8313 647 8327
rect 453 8273 467 8287
rect 553 8233 567 8247
rect 513 8196 527 8210
rect 393 8153 407 8167
rect 533 8150 547 8164
rect 513 8133 527 8147
rect 573 8133 587 8147
rect 493 7930 507 7944
rect 533 7893 547 7907
rect 533 7753 547 7767
rect 673 7873 687 7887
rect 653 7813 667 7827
rect 573 7733 587 7747
rect 633 7733 647 7747
rect 533 7713 547 7727
rect 413 7676 427 7690
rect 493 7676 507 7690
rect 573 7676 587 7690
rect 373 7593 387 7607
rect 333 7113 347 7127
rect 613 7673 627 7687
rect 653 7673 667 7687
rect 553 7630 567 7644
rect 593 7630 607 7644
rect 513 7613 527 7627
rect 533 7456 547 7470
rect 573 7456 587 7470
rect 433 7156 447 7170
rect 553 7413 567 7427
rect 493 7173 507 7187
rect 532 7156 546 7170
rect 553 7153 567 7167
rect 593 7433 607 7447
rect 653 7393 667 7407
rect 773 8433 787 8447
rect 793 8413 807 8427
rect 853 8413 867 8427
rect 753 8353 767 8367
rect 713 8193 727 8207
rect 833 8233 847 8247
rect 793 8196 807 8210
rect 773 8133 787 8147
rect 873 8153 887 8167
rect 813 8093 827 8107
rect 773 7976 787 7990
rect 753 7930 767 7944
rect 813 7913 827 7927
rect 713 7676 727 7690
rect 793 7676 807 7690
rect 793 7613 807 7627
rect 693 7593 707 7607
rect 813 7593 827 7607
rect 1093 10393 1107 10407
rect 1013 10276 1027 10290
rect 1053 10276 1067 10290
rect 1093 10276 1107 10290
rect 1153 10276 1167 10290
rect 1073 10193 1087 10207
rect 1013 10010 1027 10024
rect 1113 10013 1127 10027
rect 1153 10013 1167 10027
rect 993 9893 1007 9907
rect 1093 9893 1107 9907
rect 973 9756 987 9770
rect 1033 9756 1047 9770
rect 1013 9710 1027 9724
rect 933 9573 947 9587
rect 993 9573 1007 9587
rect 1033 9536 1047 9550
rect 953 9433 967 9447
rect 933 9113 947 9127
rect 913 8613 927 8627
rect 913 8150 927 8164
rect 913 7976 927 7990
rect 893 7593 907 7607
rect 793 7473 807 7487
rect 873 7473 887 7487
rect 753 7456 767 7470
rect 813 7410 827 7424
rect 893 7410 907 7424
rect 733 7393 747 7407
rect 693 7273 707 7287
rect 673 7193 687 7207
rect 653 7173 667 7187
rect 593 7153 607 7167
rect 673 7156 687 7170
rect 453 7113 467 7127
rect 513 7110 527 7124
rect 573 7113 587 7127
rect 413 7093 427 7107
rect 493 6936 507 6950
rect 573 6936 587 6950
rect 673 6973 687 6987
rect 533 6890 547 6904
rect 313 6853 327 6867
rect 473 6853 487 6867
rect 393 6813 407 6827
rect 253 6773 267 6787
rect 293 6773 307 6787
rect 293 6713 307 6727
rect 193 6633 207 6647
rect 253 6573 267 6587
rect 293 6573 307 6587
rect 253 6473 267 6487
rect 193 6373 207 6387
rect 213 6193 227 6207
rect 13 6153 27 6167
rect 253 5993 267 6007
rect 33 5933 47 5947
rect 13 5813 27 5827
rect 73 5893 87 5907
rect 213 5896 227 5910
rect 52 5853 66 5867
rect 73 5853 87 5867
rect 253 5813 267 5827
rect 53 5793 67 5807
rect 33 5773 47 5787
rect 13 5633 27 5647
rect 13 5593 27 5607
rect 213 5596 227 5610
rect 253 5513 267 5527
rect 193 5333 207 5347
rect 293 5333 307 5347
rect 513 6673 527 6687
rect 433 6653 447 6667
rect 473 6653 487 6667
rect 453 6593 467 6607
rect 493 6590 507 6604
rect 533 6590 547 6604
rect 453 6553 467 6567
rect 633 6590 647 6604
rect 573 6493 587 6507
rect 513 6453 527 6467
rect 773 7156 787 7170
rect 813 7156 827 7170
rect 873 7156 887 7170
rect 793 7110 807 7124
rect 833 7110 847 7124
rect 773 6936 787 6950
rect 733 6890 747 6904
rect 833 6890 847 6904
rect 893 7113 907 7127
rect 893 6936 907 6950
rect 793 6853 807 6867
rect 873 6853 887 6867
rect 773 6753 787 6767
rect 873 6753 887 6767
rect 813 6636 827 6650
rect 693 6593 707 6607
rect 753 6590 767 6604
rect 673 6553 687 6567
rect 573 6413 587 6427
rect 633 6416 647 6430
rect 733 6416 747 6430
rect 793 6573 807 6587
rect 433 6373 447 6387
rect 473 6370 487 6384
rect 433 6193 447 6207
rect 413 5493 427 5507
rect 393 5273 407 5287
rect 193 5073 207 5087
rect 293 5073 307 5087
rect 233 4993 247 5007
rect 193 4856 207 4870
rect 293 4856 307 4870
rect 213 4810 227 4824
rect 253 4810 267 4824
rect 173 4553 187 4567
rect 253 4510 267 4524
rect 253 4336 267 4350
rect 213 4290 227 4304
rect 333 4553 347 4567
rect 293 4133 307 4147
rect 213 4036 227 4050
rect 293 4033 307 4047
rect 253 3933 267 3947
rect 13 3773 27 3787
rect 193 3771 207 3785
rect 233 3733 247 3747
rect 13 3613 27 3627
rect 213 3553 227 3567
rect 293 3553 307 3567
rect 253 3516 267 3530
rect 233 3470 247 3484
rect 193 3393 207 3407
rect 273 3393 287 3407
rect 213 3296 227 3310
rect 233 3250 247 3264
rect 173 3073 187 3087
rect 173 2993 187 3007
rect 213 2996 227 3010
rect 353 3893 367 3907
rect 473 6116 487 6130
rect 573 6373 587 6387
rect 613 6173 627 6187
rect 533 6113 547 6127
rect 513 6033 527 6047
rect 453 5896 467 5910
rect 493 5850 507 5864
rect 493 5473 507 5487
rect 493 5433 507 5447
rect 473 5330 487 5344
rect 753 6370 767 6384
rect 753 6333 767 6347
rect 793 6333 807 6347
rect 873 6273 887 6287
rect 833 6233 847 6247
rect 853 6213 867 6227
rect 813 6116 827 6130
rect 793 6070 807 6084
rect 853 6033 867 6047
rect 793 5993 807 6007
rect 653 5933 667 5947
rect 733 5896 747 5910
rect 713 5853 727 5867
rect 773 5853 787 5867
rect 973 9393 987 9407
rect 1053 9490 1067 9504
rect 1013 9333 1027 9347
rect 993 9293 1007 9307
rect 1033 9236 1047 9250
rect 1273 11316 1287 11330
rect 1373 11316 1387 11330
rect 1293 11270 1307 11284
rect 1333 11233 1347 11247
rect 1253 11133 1267 11147
rect 1293 11096 1307 11110
rect 1313 11050 1327 11064
rect 1653 11773 1667 11787
rect 1573 11693 1587 11707
rect 1413 11373 1427 11387
rect 1593 11373 1607 11387
rect 1593 11333 1607 11347
rect 1513 11316 1527 11330
rect 1553 11316 1567 11330
rect 1653 11316 1667 11330
rect 1753 11836 1767 11850
rect 1753 11573 1767 11587
rect 1393 11273 1407 11287
rect 1433 11213 1447 11227
rect 1393 11096 1407 11110
rect 1393 10993 1407 11007
rect 1273 10973 1287 10987
rect 1373 10973 1387 10987
rect 1213 10813 1227 10827
rect 1313 10796 1327 10810
rect 1333 10750 1347 10764
rect 1293 10673 1307 10687
rect 1373 10673 1387 10687
rect 1313 10615 1327 10629
rect 1353 10577 1367 10591
rect 1233 10473 1247 10487
rect 1333 10473 1347 10487
rect 1353 10230 1367 10244
rect 1313 10193 1327 10207
rect 1293 10056 1307 10070
rect 1313 10010 1327 10024
rect 1213 9853 1227 9867
rect 1113 9753 1127 9767
rect 1193 9673 1207 9687
rect 1173 9653 1187 9667
rect 1173 9613 1187 9627
rect 1153 9536 1167 9550
rect 1153 9433 1167 9447
rect 1153 9293 1167 9307
rect 1133 9253 1147 9267
rect 1113 9236 1127 9250
rect 1013 9190 1027 9204
rect 1053 9190 1067 9204
rect 1093 9190 1107 9204
rect 1053 9073 1067 9087
rect 1033 9033 1047 9047
rect 993 9016 1007 9030
rect 1013 8970 1027 8984
rect 1113 8873 1127 8887
rect 993 8793 1007 8807
rect 1053 8716 1067 8730
rect 1113 8713 1127 8727
rect 993 8670 1007 8684
rect 1073 8670 1087 8684
rect 1033 8613 1047 8627
rect 973 8493 987 8507
rect 1073 8573 1087 8587
rect 1113 8496 1127 8510
rect 993 8413 1007 8427
rect 973 8393 987 8407
rect 953 8353 967 8367
rect 953 8193 967 8207
rect 1093 8450 1107 8464
rect 1053 8433 1067 8447
rect 1193 9273 1207 9287
rect 1173 9233 1187 9247
rect 1153 9193 1167 9207
rect 1193 9113 1207 9127
rect 1373 9793 1387 9807
rect 1273 9756 1287 9770
rect 1233 9713 1247 9727
rect 1253 9693 1267 9707
rect 1373 9693 1387 9707
rect 1293 9673 1307 9687
rect 1313 9573 1327 9587
rect 1373 9573 1387 9587
rect 1273 9536 1287 9550
rect 1233 9490 1247 9504
rect 1293 9490 1307 9504
rect 1333 9473 1347 9487
rect 1373 9473 1387 9487
rect 1273 9236 1287 9250
rect 1313 9236 1327 9250
rect 1373 9236 1387 9250
rect 1293 9190 1307 9204
rect 1413 10773 1427 10787
rect 1413 10533 1427 10547
rect 1453 10973 1467 10987
rect 1573 11270 1587 11284
rect 1613 11133 1627 11147
rect 1593 11096 1607 11110
rect 1533 10796 1547 10810
rect 1573 10796 1587 10810
rect 1733 11313 1747 11327
rect 1793 11873 1807 11887
rect 1913 11836 1927 11850
rect 1893 11790 1907 11804
rect 1933 11790 1947 11804
rect 2093 12090 2107 12104
rect 2153 12090 2167 12104
rect 2313 12173 2327 12187
rect 2433 12173 2447 12187
rect 2353 12136 2367 12150
rect 2433 12110 2447 12124
rect 2833 12193 2847 12207
rect 3613 12193 3627 12207
rect 2773 12133 2787 12147
rect 2573 12110 2587 12124
rect 2953 12133 2967 12147
rect 2993 12133 3007 12147
rect 3553 12136 3567 12150
rect 2833 12116 2847 12130
rect 2893 12116 2907 12130
rect 2193 11933 2207 11947
rect 2133 11836 2147 11850
rect 2373 12090 2387 12104
rect 2913 12073 2927 12087
rect 2413 12033 2427 12047
rect 2913 11993 2927 12007
rect 2413 11933 2427 11947
rect 2553 11933 2567 11947
rect 2053 11793 2067 11807
rect 1993 11693 2007 11707
rect 1853 11633 1867 11647
rect 1893 11616 1907 11630
rect 1933 11616 1947 11630
rect 2033 11616 2047 11630
rect 2093 11616 2107 11630
rect 2333 11833 2347 11847
rect 2373 11836 2387 11850
rect 2173 11790 2187 11804
rect 2373 11790 2387 11804
rect 2213 11753 2227 11767
rect 2293 11693 2307 11707
rect 1873 11570 1887 11584
rect 1793 11533 1807 11547
rect 1873 11493 1887 11507
rect 1933 11493 1947 11507
rect 1833 11316 1847 11330
rect 2093 11533 2107 11547
rect 1913 11316 1927 11330
rect 2033 11316 2047 11330
rect 1893 11270 1907 11284
rect 1773 11233 1787 11247
rect 1853 11233 1867 11247
rect 2013 11233 2027 11247
rect 1713 11133 1727 11147
rect 1833 11133 1847 11147
rect 1993 11133 2007 11147
rect 1833 11096 1847 11110
rect 1873 11096 1887 11110
rect 1913 11096 1927 11110
rect 1713 11050 1727 11064
rect 1813 11050 1827 11064
rect 1853 11050 1867 11064
rect 1953 11093 1967 11107
rect 1953 11050 1967 11064
rect 1993 11050 2007 11064
rect 1913 10973 1927 10987
rect 1693 10816 1707 10830
rect 1513 10753 1527 10767
rect 1493 10693 1507 10707
rect 1493 10573 1507 10587
rect 1453 10513 1467 10527
rect 1453 10453 1467 10467
rect 1433 10073 1447 10087
rect 1413 10056 1427 10070
rect 1413 10013 1427 10027
rect 1453 9793 1467 9807
rect 1433 9713 1447 9727
rect 1393 9193 1407 9207
rect 1373 9153 1387 9167
rect 1253 9113 1267 9127
rect 1213 9073 1227 9087
rect 1233 9053 1247 9067
rect 1313 9053 1327 9067
rect 1173 8970 1187 8984
rect 1253 9016 1267 9030
rect 1353 9033 1367 9047
rect 1413 9016 1427 9030
rect 1253 8970 1267 8984
rect 1153 8573 1167 8587
rect 1173 8450 1187 8464
rect 1333 8970 1347 8984
rect 1293 8953 1307 8967
rect 1293 8753 1307 8767
rect 1333 8716 1347 8730
rect 1373 8716 1387 8730
rect 1373 8673 1387 8687
rect 1313 8533 1327 8547
rect 1293 8496 1307 8510
rect 1333 8496 1347 8510
rect 1253 8413 1267 8427
rect 1313 8393 1327 8407
rect 1353 8373 1367 8387
rect 1233 8333 1247 8347
rect 1152 8313 1166 8327
rect 1173 8313 1187 8327
rect 1093 8196 1107 8210
rect 1133 8195 1147 8209
rect 1193 8195 1207 8209
rect 1013 8153 1027 8167
rect 1073 8150 1087 8164
rect 953 7913 967 7927
rect 933 7653 947 7667
rect 933 7456 947 7470
rect 1053 7993 1067 8007
rect 1113 7973 1127 7987
rect 1013 7913 1027 7927
rect 1053 7873 1067 7887
rect 1053 7773 1067 7787
rect 1033 7673 1047 7687
rect 1093 7713 1107 7727
rect 1153 7673 1167 7687
rect 1033 7633 1047 7647
rect 993 7453 1007 7467
rect 1073 7630 1087 7644
rect 1113 7630 1127 7644
rect 1153 7630 1167 7644
rect 1173 7613 1187 7627
rect 1073 7593 1087 7607
rect 1093 7410 1107 7424
rect 1133 7410 1147 7424
rect 1053 7373 1067 7387
rect 1053 7156 1067 7170
rect 1093 7156 1107 7170
rect 1073 7110 1087 7124
rect 1133 7113 1147 7127
rect 1053 7073 1067 7087
rect 933 6936 947 6950
rect 1013 6936 1027 6950
rect 1213 7976 1227 7990
rect 1193 7073 1207 7087
rect 1213 7053 1227 7067
rect 1113 6973 1127 6987
rect 1173 6973 1187 6987
rect 933 6813 947 6827
rect 1033 6813 1047 6827
rect 1113 6813 1127 6827
rect 1073 6753 1087 6767
rect 953 6713 967 6727
rect 973 6633 987 6647
rect 1113 6636 1127 6650
rect 953 6593 967 6607
rect 913 6573 927 6587
rect 933 6373 947 6387
rect 1093 6573 1107 6587
rect 1053 6533 1067 6547
rect 1093 6513 1107 6527
rect 1053 6493 1067 6507
rect 1093 6416 1107 6430
rect 1253 8233 1267 8247
rect 1253 8196 1267 8210
rect 1333 8196 1347 8210
rect 1353 8133 1367 8147
rect 1253 8113 1267 8127
rect 1393 7993 1407 8007
rect 1293 7976 1307 7990
rect 1313 7930 1327 7944
rect 1353 7713 1367 7727
rect 1313 7676 1327 7690
rect 1313 7453 1327 7467
rect 1353 7473 1367 7487
rect 1433 8193 1447 8207
rect 1413 7933 1427 7947
rect 1653 10793 1667 10807
rect 1633 10750 1647 10764
rect 1593 10733 1607 10747
rect 1573 10576 1587 10590
rect 1593 10513 1607 10527
rect 1853 10776 1867 10790
rect 1833 10613 1847 10627
rect 1993 10553 2007 10567
rect 1813 10530 1827 10544
rect 1913 10493 1927 10507
rect 1813 10453 1827 10467
rect 1913 10453 1927 10467
rect 1813 10413 1827 10427
rect 1673 10393 1687 10407
rect 1533 10353 1547 10367
rect 1573 10276 1587 10290
rect 1653 10276 1667 10290
rect 1533 10073 1547 10087
rect 1553 10010 1567 10024
rect 1653 10230 1667 10244
rect 1613 9893 1627 9907
rect 1633 9833 1647 9847
rect 1593 9793 1607 9807
rect 1493 9756 1507 9770
rect 1553 9756 1567 9770
rect 1653 9813 1667 9827
rect 1633 9756 1647 9770
rect 1473 9553 1487 9567
rect 1573 9710 1587 9724
rect 1613 9710 1627 9724
rect 1653 9710 1667 9724
rect 1593 9573 1607 9587
rect 1553 9553 1567 9567
rect 1613 9553 1627 9567
rect 1493 9473 1507 9487
rect 1473 9173 1487 9187
rect 1473 9033 1487 9047
rect 1593 9473 1607 9487
rect 1613 9473 1627 9487
rect 1573 9433 1587 9447
rect 1553 9273 1567 9287
rect 1613 9433 1627 9447
rect 1733 10193 1747 10207
rect 1633 9233 1647 9247
rect 1533 9173 1547 9187
rect 1573 9153 1587 9167
rect 1593 9073 1607 9087
rect 1553 9016 1567 9030
rect 1693 9113 1707 9127
rect 1673 9013 1687 9027
rect 1613 8970 1627 8984
rect 1673 8970 1687 8984
rect 1493 8953 1507 8967
rect 1573 8953 1587 8967
rect 1533 8753 1547 8767
rect 1573 8753 1587 8767
rect 1473 8493 1487 8507
rect 1513 8496 1527 8510
rect 1493 8173 1507 8187
rect 1473 8013 1487 8027
rect 1453 7993 1467 8007
rect 1613 8716 1627 8730
rect 1593 8670 1607 8684
rect 1633 8653 1647 8667
rect 1613 8613 1627 8627
rect 1653 8613 1667 8627
rect 1613 8533 1627 8547
rect 1773 10093 1787 10107
rect 1753 10073 1767 10087
rect 1773 10053 1787 10067
rect 1873 10276 1887 10290
rect 1973 10276 1987 10290
rect 1913 10193 1927 10207
rect 1893 10093 1907 10107
rect 1873 10053 1887 10067
rect 1793 10010 1807 10024
rect 1833 9993 1847 10007
rect 1873 9993 1887 10007
rect 1793 9893 1807 9907
rect 1853 9853 1867 9867
rect 1973 10233 1987 10247
rect 1953 10053 1967 10067
rect 1933 9873 1947 9887
rect 1893 9756 1907 9770
rect 1833 9693 1847 9707
rect 1873 9613 1887 9627
rect 1793 9553 1807 9567
rect 1853 9536 1867 9550
rect 1933 9533 1947 9547
rect 1833 9453 1847 9467
rect 1933 9353 1947 9367
rect 1873 9313 1887 9327
rect 1813 9293 1827 9307
rect 1753 9273 1767 9287
rect 1733 8673 1747 8687
rect 1853 9236 1867 9250
rect 1893 9236 1907 9250
rect 1793 9190 1807 9204
rect 1833 9190 1847 9204
rect 1773 8573 1787 8587
rect 1753 8553 1767 8567
rect 1693 8533 1707 8547
rect 1653 8496 1667 8510
rect 1673 8450 1687 8464
rect 1773 8450 1787 8464
rect 1633 8433 1647 8447
rect 1753 8373 1767 8387
rect 1533 8196 1547 8210
rect 1613 8196 1627 8210
rect 1653 8196 1667 8210
rect 1633 8150 1647 8164
rect 1873 9113 1887 9127
rect 1973 9553 1987 9567
rect 1813 9093 1827 9107
rect 1953 9093 1967 9107
rect 1833 9053 1847 9067
rect 1813 8953 1827 8967
rect 1893 9016 1907 9030
rect 1933 9016 1947 9030
rect 1873 8953 1887 8967
rect 1973 8953 1987 8967
rect 1913 8933 1927 8947
rect 1833 8873 1847 8887
rect 2153 11533 2167 11547
rect 2113 11493 2127 11507
rect 2173 11493 2187 11507
rect 2333 11673 2347 11687
rect 3153 12110 3167 12124
rect 3273 12116 3287 12130
rect 3353 12113 3367 12127
rect 3193 11993 3207 12007
rect 2473 11836 2487 11850
rect 2513 11836 2527 11850
rect 2573 11813 2587 11827
rect 2433 11793 2447 11807
rect 2493 11790 2507 11804
rect 2413 11713 2427 11727
rect 2533 11713 2547 11727
rect 2573 11713 2587 11727
rect 2413 11653 2427 11667
rect 2373 11633 2387 11647
rect 2493 11633 2507 11647
rect 2473 11593 2487 11607
rect 2333 11570 2347 11584
rect 2393 11570 2407 11584
rect 2553 11633 2567 11647
rect 2533 11550 2547 11564
rect 2513 11513 2527 11527
rect 2133 11316 2147 11330
rect 2173 11316 2187 11330
rect 2233 11316 2247 11330
rect 2293 11316 2307 11330
rect 2453 11316 2467 11330
rect 2093 11273 2107 11287
rect 2153 11270 2167 11284
rect 2193 11213 2207 11227
rect 2133 11173 2147 11187
rect 2233 11173 2247 11187
rect 2093 11096 2107 11110
rect 2233 11096 2247 11110
rect 2033 10993 2047 11007
rect 2113 11050 2127 11064
rect 2153 10993 2167 11007
rect 2073 10973 2087 10987
rect 2033 10753 2047 10767
rect 2113 10770 2127 10784
rect 2053 10733 2067 10747
rect 2173 10770 2187 10784
rect 2073 10713 2087 10727
rect 2153 10713 2167 10727
rect 2033 10673 2047 10687
rect 2113 10576 2127 10590
rect 2273 10973 2287 10987
rect 2233 10613 2247 10627
rect 2193 10576 2207 10590
rect 2173 10433 2187 10447
rect 2093 10413 2107 10427
rect 2053 10353 2067 10367
rect 2113 10276 2127 10290
rect 2153 10276 2167 10290
rect 2413 11270 2427 11284
rect 2493 11270 2507 11284
rect 2473 11113 2487 11127
rect 2313 11096 2327 11110
rect 2353 11096 2367 11110
rect 2393 11096 2407 11110
rect 2453 11093 2467 11107
rect 2453 11052 2467 11066
rect 2413 11033 2427 11047
rect 2373 10933 2387 10947
rect 2313 10893 2327 10907
rect 2353 10893 2367 10907
rect 2313 10793 2327 10807
rect 2393 10750 2407 10764
rect 2313 10733 2327 10747
rect 2373 10693 2387 10707
rect 2433 10573 2447 10587
rect 2293 10553 2307 10567
rect 2353 10530 2367 10544
rect 2433 10530 2447 10544
rect 2353 10473 2367 10487
rect 2273 10453 2287 10467
rect 2273 10313 2287 10327
rect 2233 10276 2247 10290
rect 2053 10193 2067 10207
rect 2213 10213 2227 10227
rect 2273 10213 2287 10227
rect 2173 10193 2187 10207
rect 2053 10056 2067 10070
rect 2133 10053 2147 10067
rect 2213 10053 2227 10067
rect 2013 9973 2027 9987
rect 2073 9993 2087 10007
rect 2113 9973 2127 9987
rect 2193 9893 2207 9907
rect 2173 9873 2187 9887
rect 2053 9710 2067 9724
rect 2093 9710 2107 9724
rect 2013 9693 2027 9707
rect 2033 9533 2047 9547
rect 2013 8913 2027 8927
rect 2013 8853 2027 8867
rect 1933 8793 1947 8807
rect 1853 8716 1867 8730
rect 1833 8670 1847 8684
rect 1793 8333 1807 8347
rect 1853 8496 1867 8510
rect 1893 8496 1907 8510
rect 1833 8313 1847 8327
rect 1913 8433 1927 8447
rect 1953 8413 1967 8427
rect 1893 8373 1907 8387
rect 1973 8273 1987 8287
rect 1973 8233 1987 8247
rect 1933 8196 1947 8210
rect 1853 8173 1867 8187
rect 1573 8133 1587 8147
rect 1673 8113 1687 8127
rect 1673 8013 1687 8027
rect 1513 7976 1527 7990
rect 1573 7976 1587 7990
rect 1493 7933 1507 7947
rect 1433 7773 1447 7787
rect 1393 7456 1407 7470
rect 1453 7456 1467 7470
rect 1333 7410 1347 7424
rect 1413 7393 1427 7407
rect 1373 7373 1387 7387
rect 1253 7353 1267 7367
rect 1253 7233 1267 7247
rect 1233 6573 1247 6587
rect 1173 6513 1187 6527
rect 1213 6493 1227 6507
rect 1153 6453 1167 6467
rect 1133 6413 1147 6427
rect 1213 6396 1227 6410
rect 913 6173 927 6187
rect 893 5893 907 5907
rect 772 5793 786 5807
rect 793 5793 807 5807
rect 973 6370 987 6384
rect 1033 6370 1047 6384
rect 1033 6313 1047 6327
rect 993 6173 1007 6187
rect 1113 6373 1127 6387
rect 1073 6273 1087 6287
rect 1193 6353 1207 6367
rect 1113 6193 1127 6207
rect 1293 7173 1307 7187
rect 1333 7156 1347 7170
rect 1313 7110 1327 7124
rect 1353 7053 1367 7067
rect 1393 6973 1407 6987
rect 1473 7156 1487 7170
rect 1453 6913 1467 6927
rect 1273 6853 1287 6867
rect 1293 6833 1307 6847
rect 1373 6890 1387 6904
rect 1333 6733 1347 6747
rect 1353 6636 1367 6650
rect 1393 6636 1407 6650
rect 1453 6636 1467 6650
rect 1373 6590 1387 6604
rect 1413 6590 1427 6604
rect 1673 7950 1687 7964
rect 1753 8153 1767 8167
rect 1913 8150 1927 8164
rect 2093 9553 2107 9567
rect 2173 9533 2187 9547
rect 2053 9453 2067 9467
rect 2153 9490 2167 9504
rect 2113 9433 2127 9447
rect 2053 9313 2067 9327
rect 2213 9353 2227 9367
rect 2193 9293 2207 9307
rect 2153 9253 2167 9267
rect 2073 9236 2087 9250
rect 2193 9236 2207 9250
rect 2073 9193 2087 9207
rect 2133 9190 2147 9204
rect 2053 9153 2067 9167
rect 2173 9153 2187 9167
rect 2373 10373 2387 10387
rect 2473 11033 2487 11047
rect 2493 10753 2507 10767
rect 2493 10613 2507 10627
rect 2533 11030 2547 11044
rect 2533 10816 2547 10830
rect 2473 10473 2487 10487
rect 2393 10353 2407 10367
rect 2453 10353 2467 10367
rect 2373 10276 2387 10290
rect 2313 10193 2327 10207
rect 2473 10276 2487 10290
rect 2533 10293 2547 10307
rect 2513 10273 2527 10287
rect 2453 10230 2467 10244
rect 2493 10230 2507 10244
rect 2473 10213 2487 10227
rect 2453 10173 2467 10187
rect 2533 10173 2547 10187
rect 2613 11816 2627 11830
rect 2713 11816 2727 11830
rect 2893 11810 2907 11824
rect 2613 11773 2627 11787
rect 2973 11810 2987 11824
rect 3533 11993 3547 12007
rect 3233 11836 3247 11850
rect 2913 11733 2927 11747
rect 3013 11733 3027 11747
rect 3113 11733 3127 11747
rect 2893 11713 2907 11727
rect 2793 11653 2807 11667
rect 3073 11653 3087 11667
rect 3113 11653 3127 11667
rect 2613 11613 2627 11627
rect 2693 11616 2707 11630
rect 2593 11593 2607 11607
rect 2792 11596 2806 11610
rect 2813 11590 2827 11604
rect 2913 11590 2927 11604
rect 2753 11550 2767 11564
rect 2713 11513 2727 11527
rect 2713 11453 2727 11467
rect 2653 11270 2667 11284
rect 2673 11113 2687 11127
rect 2613 11070 2627 11084
rect 2893 11393 2907 11407
rect 2993 11316 3007 11330
rect 2893 11270 2907 11284
rect 2973 11270 2987 11284
rect 3033 11213 3047 11227
rect 2933 11173 2947 11187
rect 3053 11173 3067 11187
rect 2893 11070 2907 11084
rect 2693 11050 2707 11064
rect 2733 11030 2747 11044
rect 2713 10993 2727 11007
rect 2653 10893 2667 10907
rect 2573 10813 2587 10827
rect 2553 10133 2567 10147
rect 2493 10113 2507 10127
rect 2473 9993 2487 10007
rect 2293 9973 2307 9987
rect 2333 9973 2347 9987
rect 2373 9973 2387 9987
rect 2313 9853 2327 9867
rect 2473 9793 2487 9807
rect 2373 9756 2387 9770
rect 2413 9756 2427 9770
rect 2313 9710 2327 9724
rect 2253 9490 2267 9504
rect 2233 9093 2247 9107
rect 2213 9053 2227 9067
rect 2053 9016 2067 9030
rect 2173 9016 2187 9030
rect 2193 8970 2207 8984
rect 2153 8953 2167 8967
rect 2093 8933 2107 8947
rect 2033 8653 2047 8667
rect 2073 8653 2087 8667
rect 2093 8496 2107 8510
rect 2193 8613 2207 8627
rect 2173 8496 2187 8510
rect 2233 8493 2247 8507
rect 2113 8453 2127 8467
rect 2193 8450 2207 8464
rect 2233 8413 2247 8427
rect 2273 9453 2287 9467
rect 2293 9053 2307 9067
rect 2293 8933 2307 8947
rect 2293 8753 2307 8767
rect 2273 8593 2287 8607
rect 2273 8533 2287 8547
rect 2093 8333 2107 8347
rect 2253 8333 2267 8347
rect 2033 8293 2047 8307
rect 2013 8073 2027 8087
rect 1973 8033 1987 8047
rect 1813 7950 1827 7964
rect 1553 7930 1567 7944
rect 1653 7910 1667 7924
rect 1613 7893 1627 7907
rect 1793 7813 1807 7827
rect 1593 7713 1607 7727
rect 1733 7713 1747 7727
rect 1653 7676 1667 7690
rect 1613 7613 1627 7627
rect 1533 7456 1547 7470
rect 1693 7456 1707 7470
rect 1513 7033 1527 7047
rect 1673 7410 1687 7424
rect 1633 7373 1647 7387
rect 1613 7353 1627 7367
rect 1613 7313 1627 7327
rect 1573 7233 1587 7247
rect 1573 7156 1587 7170
rect 1653 7253 1667 7267
rect 1593 7110 1607 7124
rect 1533 6973 1547 6987
rect 1653 6933 1667 6947
rect 1613 6890 1627 6904
rect 1493 6633 1507 6647
rect 1493 6590 1507 6604
rect 1473 6573 1487 6587
rect 1493 6553 1507 6567
rect 1453 6513 1467 6527
rect 1273 6493 1287 6507
rect 1273 6413 1287 6427
rect 1413 6390 1427 6404
rect 1633 6636 1647 6650
rect 1273 6353 1287 6367
rect 1253 6313 1267 6327
rect 1573 6313 1587 6327
rect 1213 6273 1227 6287
rect 1193 6133 1207 6147
rect 1033 6116 1047 6130
rect 1173 6090 1187 6104
rect 1033 5993 1047 6007
rect 993 5933 1007 5947
rect 1053 5853 1067 5867
rect 993 5773 1007 5787
rect 1053 5773 1067 5787
rect 933 5713 947 5727
rect 713 5693 727 5707
rect 813 5653 827 5667
rect 753 5633 767 5647
rect 673 5593 687 5607
rect 653 5553 667 5567
rect 633 5493 647 5507
rect 733 5550 747 5564
rect 773 5493 787 5507
rect 833 5633 847 5647
rect 833 5513 847 5527
rect 813 5433 827 5447
rect 753 5413 767 5427
rect 693 5373 707 5387
rect 1113 6073 1127 6087
rect 1073 5613 1087 5627
rect 993 5596 1007 5610
rect 1033 5550 1047 5564
rect 1073 5550 1087 5564
rect 1133 5553 1147 5567
rect 973 5350 987 5364
rect 713 5330 727 5344
rect 633 5313 647 5327
rect 673 5313 687 5327
rect 773 5313 787 5327
rect 613 5093 627 5107
rect 473 5076 487 5090
rect 453 5033 467 5047
rect 433 4993 447 5007
rect 413 4853 427 4867
rect 493 4953 507 4967
rect 493 4810 507 4824
rect 553 4810 567 4824
rect 453 4773 467 4787
rect 513 4593 527 4607
rect 473 4556 487 4570
rect 573 4773 587 4787
rect 573 4733 587 4747
rect 553 4556 567 4570
rect 433 4510 447 4524
rect 493 4510 507 4524
rect 413 4336 427 4350
rect 413 4293 427 4307
rect 553 4493 567 4507
rect 493 4336 507 4350
rect 533 4336 547 4350
rect 533 4173 547 4187
rect 553 4053 567 4067
rect 473 4036 487 4050
rect 513 3993 527 4007
rect 493 3973 507 3987
rect 333 3516 347 3530
rect 333 3433 347 3447
rect 313 3373 327 3387
rect 293 3296 307 3310
rect 273 2993 287 3007
rect 193 2950 207 2964
rect 333 3153 347 3167
rect 173 2773 187 2787
rect 233 2776 247 2790
rect 273 2776 287 2790
rect 333 2776 347 2790
rect 173 2713 187 2727
rect 253 2713 267 2727
rect 213 2693 227 2707
rect 213 2533 227 2547
rect 193 2473 207 2487
rect 253 2493 267 2507
rect 293 2493 307 2507
rect 193 2433 207 2447
rect 193 2253 207 2267
rect 253 2313 267 2327
rect 193 2213 207 2227
rect 193 1993 207 2007
rect 273 2210 287 2224
rect 333 2213 347 2227
rect 293 1993 307 2007
rect 233 1973 247 1987
rect 173 1956 187 1970
rect 213 1956 227 1970
rect 253 1956 267 1970
rect 193 1853 207 1867
rect 273 1913 287 1927
rect 233 1753 247 1767
rect 333 1793 347 1807
rect 313 1753 327 1767
rect 293 1733 307 1747
rect 153 1690 167 1704
rect 213 1690 227 1704
rect 253 1690 267 1704
rect 193 1435 207 1449
rect 613 4973 627 4987
rect 593 4313 607 4327
rect 593 4133 607 4147
rect 573 3993 587 4007
rect 593 3953 607 3967
rect 553 3933 567 3947
rect 813 5233 827 5247
rect 953 5233 967 5247
rect 1013 5153 1027 5167
rect 653 5093 667 5107
rect 953 5096 967 5110
rect 993 5093 1007 5107
rect 793 5056 807 5070
rect 653 5033 667 5047
rect 673 4953 687 4967
rect 853 4933 867 4947
rect 813 4893 827 4907
rect 893 4853 907 4867
rect 633 4810 647 4824
rect 673 4813 687 4827
rect 833 4810 847 4824
rect 793 4773 807 4787
rect 893 4773 907 4787
rect 1013 5056 1027 5070
rect 1533 6136 1547 6150
rect 1373 6096 1387 6110
rect 1473 6096 1487 6110
rect 1473 6053 1487 6067
rect 1273 5933 1287 5947
rect 1313 5896 1327 5910
rect 1213 5850 1227 5864
rect 1293 5850 1307 5864
rect 1253 5733 1267 5747
rect 1333 5713 1347 5727
rect 1253 5693 1267 5707
rect 1293 5596 1307 5610
rect 1353 5596 1367 5610
rect 1193 5553 1207 5567
rect 1273 5550 1287 5564
rect 1233 5533 1247 5547
rect 1273 5529 1287 5543
rect 1193 5350 1207 5364
rect 1233 5356 1247 5370
rect 1193 5113 1207 5127
rect 1233 5076 1247 5090
rect 1133 4973 1147 4987
rect 1213 5030 1227 5044
rect 1313 5493 1327 5507
rect 1293 5393 1307 5407
rect 1173 4933 1187 4947
rect 1273 4933 1287 4947
rect 1013 4893 1027 4907
rect 1053 4893 1067 4907
rect 1093 4856 1107 4870
rect 1133 4856 1147 4870
rect 1033 4810 1047 4824
rect 1013 4653 1027 4667
rect 653 4613 667 4627
rect 993 4613 1007 4627
rect 1073 4613 1087 4627
rect 633 4313 647 4327
rect 773 4573 787 4587
rect 693 4556 707 4570
rect 733 4556 747 4570
rect 1013 4573 1027 4587
rect 1113 4753 1127 4767
rect 1253 4856 1267 4870
rect 1173 4693 1187 4707
rect 1113 4653 1127 4667
rect 1333 5356 1347 5370
rect 1313 5113 1327 5127
rect 1313 5076 1327 5090
rect 1393 5753 1407 5767
rect 1373 5313 1387 5327
rect 1373 5173 1387 5187
rect 1373 5033 1387 5047
rect 1313 4953 1327 4967
rect 1333 4856 1347 4870
rect 1453 5933 1467 5947
rect 1433 5453 1447 5467
rect 1513 6093 1527 6107
rect 1533 6053 1547 6067
rect 1733 7372 1747 7386
rect 1713 6613 1727 6627
rect 1693 6390 1707 6404
rect 1673 6273 1687 6287
rect 1653 6213 1667 6227
rect 1593 6133 1607 6147
rect 1633 6093 1647 6107
rect 1653 6073 1667 6087
rect 1613 5973 1627 5987
rect 1573 5933 1587 5947
rect 1693 6136 1707 6150
rect 1453 5393 1467 5407
rect 1573 5833 1587 5847
rect 1673 5933 1687 5947
rect 1693 5833 1707 5847
rect 1673 5793 1687 5807
rect 1673 5733 1687 5747
rect 1673 5693 1687 5707
rect 1653 5673 1667 5687
rect 1673 5613 1687 5627
rect 1553 5596 1567 5610
rect 1633 5596 1647 5610
rect 1573 5533 1587 5547
rect 1613 5513 1627 5527
rect 1533 5493 1547 5507
rect 1533 5376 1547 5390
rect 1453 5313 1467 5327
rect 1433 5273 1447 5287
rect 1433 5113 1447 5127
rect 1473 5293 1487 5307
rect 1513 5273 1527 5287
rect 1533 5233 1547 5247
rect 1493 5113 1507 5127
rect 1453 5073 1467 5087
rect 1673 5573 1687 5587
rect 1633 5493 1647 5507
rect 1713 5753 1727 5767
rect 1713 5453 1727 5467
rect 1893 7733 1907 7747
rect 1833 7676 1847 7690
rect 1853 7630 1867 7644
rect 1893 7630 1907 7644
rect 1833 7613 1847 7627
rect 1813 7353 1827 7367
rect 1833 7293 1847 7307
rect 1813 7273 1827 7287
rect 1933 7493 1947 7507
rect 1913 7410 1927 7424
rect 1873 7213 1887 7227
rect 1813 7193 1827 7207
rect 1853 7193 1867 7207
rect 1813 7153 1827 7167
rect 2013 7993 2027 8007
rect 2193 8233 2207 8247
rect 2073 8196 2087 8210
rect 2113 8196 2127 8210
rect 2153 8196 2167 8210
rect 2113 8113 2127 8127
rect 2173 8093 2187 8107
rect 2153 8073 2167 8087
rect 2213 8073 2227 8087
rect 2073 7956 2087 7970
rect 2133 7956 2147 7970
rect 2033 7913 2047 7927
rect 1993 7753 2007 7767
rect 2053 7673 2067 7687
rect 2173 7993 2187 8007
rect 2153 7813 2167 7827
rect 2113 7630 2127 7644
rect 2133 7456 2147 7470
rect 2193 7953 2207 7967
rect 2353 9710 2367 9724
rect 2393 9673 2407 9687
rect 2473 9673 2487 9687
rect 2353 9593 2367 9607
rect 2333 9533 2347 9547
rect 2393 9536 2407 9550
rect 2473 9536 2487 9550
rect 2353 9490 2367 9504
rect 2413 9490 2427 9504
rect 2413 9273 2427 9287
rect 2473 9273 2487 9287
rect 2333 9232 2347 9246
rect 2453 9236 2467 9250
rect 2433 9153 2447 9167
rect 2393 9133 2407 9147
rect 2473 9133 2487 9147
rect 2352 9013 2366 9027
rect 2373 9016 2387 9030
rect 2433 9016 2447 9030
rect 2613 10796 2627 10810
rect 3173 11596 3187 11610
rect 3233 11596 3247 11610
rect 3233 11453 3247 11467
rect 3213 11393 3227 11407
rect 3213 11353 3227 11367
rect 3173 11333 3187 11347
rect 3133 11233 3147 11247
rect 3313 11893 3327 11907
rect 3433 11836 3447 11850
rect 3473 11836 3487 11850
rect 3513 11836 3527 11850
rect 3433 11753 3447 11767
rect 3573 11713 3587 11727
rect 3413 11616 3427 11630
rect 3453 11616 3467 11630
rect 3492 11616 3506 11630
rect 3513 11613 3527 11627
rect 3513 11553 3527 11567
rect 3833 12173 3847 12187
rect 3753 12153 3767 12167
rect 3633 12133 3647 12147
rect 3673 12133 3687 12147
rect 3873 12153 3887 12167
rect 4093 12136 4107 12150
rect 3853 12090 3867 12104
rect 3913 12090 3927 12104
rect 3673 12033 3687 12047
rect 3713 11836 3727 11850
rect 3913 12053 3927 12067
rect 4573 12193 4587 12207
rect 4673 12193 4687 12207
rect 4533 12173 4547 12187
rect 4373 12136 4387 12150
rect 4553 12133 4567 12147
rect 4393 12090 4407 12104
rect 4532 12093 4546 12107
rect 4553 12090 4567 12104
rect 4353 12013 4367 12027
rect 4133 11953 4147 11967
rect 4173 11953 4187 11967
rect 4233 11893 4247 11907
rect 3813 11810 3827 11824
rect 3853 11813 3867 11827
rect 3793 11713 3807 11727
rect 3733 11633 3747 11647
rect 3773 11633 3787 11647
rect 3713 11616 3727 11630
rect 3693 11533 3707 11547
rect 3613 11433 3627 11447
rect 3693 11353 3707 11367
rect 3253 11333 3267 11347
rect 3293 11336 3307 11350
rect 3773 11570 3787 11584
rect 3753 11353 3767 11367
rect 3613 11333 3627 11347
rect 3233 11270 3247 11284
rect 3453 11296 3467 11310
rect 3593 11296 3607 11310
rect 3593 11253 3607 11267
rect 3333 11233 3347 11247
rect 3593 11173 3607 11187
rect 3173 11153 3187 11167
rect 3713 11290 3727 11304
rect 3753 11290 3767 11304
rect 3653 11233 3667 11247
rect 3613 11113 3627 11127
rect 3693 11113 3707 11127
rect 3173 11093 3187 11107
rect 3213 11093 3227 11107
rect 3153 11076 3167 11090
rect 3273 11093 3287 11107
rect 3313 11093 3327 11107
rect 3573 11093 3587 11107
rect 3233 11033 3247 11047
rect 2913 10873 2927 10887
rect 3053 10873 3067 10887
rect 2753 10813 2767 10827
rect 2713 10793 2727 10807
rect 2713 10753 2727 10767
rect 2673 10713 2687 10727
rect 2653 10693 2667 10707
rect 2673 10673 2687 10687
rect 2873 10753 2887 10767
rect 2813 10653 2827 10667
rect 3473 11070 3487 11084
rect 3593 11076 3607 11090
rect 3673 11073 3687 11087
rect 3633 11030 3647 11044
rect 3313 10993 3327 11007
rect 3693 11030 3707 11044
rect 3833 11653 3847 11667
rect 3313 10933 3327 10947
rect 3793 11013 3807 11027
rect 3633 10893 3647 10907
rect 3773 10893 3787 10907
rect 3073 10776 3087 10790
rect 3473 10833 3487 10847
rect 3593 10833 3607 10847
rect 3293 10813 3307 10827
rect 3193 10770 3207 10784
rect 3273 10773 3287 10787
rect 3193 10713 3207 10727
rect 2913 10673 2927 10687
rect 2973 10673 2987 10687
rect 3153 10673 3167 10687
rect 2873 10633 2887 10647
rect 2793 10613 2807 10627
rect 2633 10576 2647 10590
rect 2753 10576 2767 10590
rect 2613 10530 2627 10544
rect 2573 10073 2587 10087
rect 2553 10056 2567 10070
rect 2573 10010 2587 10024
rect 2593 9973 2607 9987
rect 2573 9893 2587 9907
rect 2533 9873 2547 9887
rect 2573 9773 2587 9787
rect 2513 9413 2527 9427
rect 2373 8973 2387 8987
rect 2413 8933 2427 8947
rect 2473 8893 2487 8907
rect 2333 8793 2347 8807
rect 2353 8773 2367 8787
rect 2393 8653 2407 8667
rect 2373 8593 2387 8607
rect 2433 8496 2447 8510
rect 2373 8450 2387 8464
rect 2413 8450 2427 8464
rect 2453 8393 2467 8407
rect 2433 8353 2447 8367
rect 2353 8313 2367 8327
rect 2312 8073 2326 8087
rect 2333 8073 2347 8087
rect 2293 8033 2307 8047
rect 2393 8273 2407 8287
rect 2373 8173 2387 8187
rect 2353 8013 2367 8027
rect 2333 7993 2347 8007
rect 2253 7972 2267 7986
rect 2293 7976 2307 7990
rect 2233 7930 2247 7944
rect 2453 8333 2467 8347
rect 2553 9633 2567 9647
rect 2593 9653 2607 9667
rect 2753 10493 2767 10507
rect 2713 10373 2727 10387
rect 2753 10313 2767 10327
rect 2653 10233 2667 10247
rect 2733 10230 2747 10244
rect 2753 10213 2767 10227
rect 2633 10133 2647 10147
rect 2733 10073 2747 10087
rect 2693 10053 2707 10067
rect 2693 10010 2707 10024
rect 2653 9853 2667 9867
rect 2713 9833 2727 9847
rect 2713 9793 2727 9807
rect 2732 9776 2746 9790
rect 2873 10576 2887 10590
rect 2933 10576 2947 10590
rect 2893 10530 2907 10544
rect 2953 10530 2967 10544
rect 2793 10113 2807 10127
rect 2913 10493 2927 10507
rect 2913 10433 2927 10447
rect 2933 10273 2947 10287
rect 2913 9973 2927 9987
rect 2873 9873 2887 9887
rect 3073 10633 3087 10647
rect 3033 10576 3047 10590
rect 2993 10293 3007 10307
rect 2973 10273 2987 10287
rect 3053 10313 3067 10327
rect 3033 10273 3047 10287
rect 2953 10213 2967 10227
rect 3053 10233 3067 10247
rect 3253 10573 3267 10587
rect 3173 10530 3187 10544
rect 3333 10793 3347 10807
rect 3373 10793 3387 10807
rect 3333 10693 3347 10707
rect 3313 10673 3327 10687
rect 3373 10653 3387 10667
rect 3453 10576 3467 10590
rect 3553 10713 3567 10727
rect 3313 10530 3327 10544
rect 3473 10530 3487 10544
rect 3513 10530 3527 10544
rect 3433 10493 3447 10507
rect 3593 10473 3607 10487
rect 3673 10833 3687 10847
rect 3753 10833 3767 10847
rect 3293 10433 3307 10447
rect 3313 10413 3327 10427
rect 3153 10333 3167 10347
rect 3133 10276 3147 10290
rect 3253 10333 3267 10347
rect 3213 10276 3227 10290
rect 3713 10796 3727 10810
rect 3833 11233 3847 11247
rect 3913 11813 3927 11827
rect 4073 11816 4087 11830
rect 3893 11753 3907 11767
rect 3873 11653 3887 11667
rect 4033 11713 4047 11727
rect 3993 11693 4007 11707
rect 3973 11570 3987 11584
rect 4013 11570 4027 11584
rect 4113 11570 4127 11584
rect 4033 11533 4047 11547
rect 3953 11433 3967 11447
rect 3893 11393 3907 11407
rect 3993 11316 4007 11330
rect 3893 11173 3907 11187
rect 3853 11096 3867 11110
rect 3973 11270 3987 11284
rect 4113 11513 4127 11527
rect 4033 11233 4047 11247
rect 4073 11153 4087 11167
rect 3933 11093 3947 11107
rect 3953 11096 3967 11110
rect 3853 10933 3867 10947
rect 3733 10750 3747 10764
rect 3773 10713 3787 10727
rect 3733 10633 3747 10647
rect 3773 10613 3787 10627
rect 3813 10613 3827 10627
rect 3773 10576 3787 10590
rect 3833 10553 3847 10567
rect 3933 11053 3947 11067
rect 3913 10993 3927 11007
rect 3873 10693 3887 10707
rect 3893 10633 3907 10647
rect 3893 10573 3907 10587
rect 3713 10530 3727 10544
rect 3793 10513 3807 10527
rect 3833 10513 3847 10527
rect 3753 10473 3767 10487
rect 3773 10413 3787 10427
rect 3813 10473 3827 10487
rect 3673 10313 3687 10327
rect 3613 10293 3627 10307
rect 3653 10293 3667 10307
rect 3233 10230 3247 10244
rect 3473 10256 3487 10270
rect 3633 10256 3647 10270
rect 3173 10213 3187 10227
rect 3353 10213 3367 10227
rect 3613 10213 3627 10227
rect 3033 10153 3047 10167
rect 3133 10153 3147 10167
rect 3633 10193 3647 10207
rect 3733 10250 3747 10264
rect 3693 10213 3707 10227
rect 3193 10093 3207 10107
rect 3673 10093 3687 10107
rect 3073 10056 3087 10070
rect 3133 10036 3147 10050
rect 3233 10036 3247 10050
rect 3033 10010 3047 10024
rect 3093 10010 3107 10024
rect 3013 9973 3027 9987
rect 3193 9973 3207 9987
rect 3053 9893 3067 9907
rect 2833 9853 2847 9867
rect 2933 9853 2947 9867
rect 2773 9833 2787 9847
rect 2773 9793 2787 9807
rect 2753 9773 2767 9787
rect 3033 9773 3047 9787
rect 2693 9756 2707 9770
rect 2753 9733 2767 9747
rect 2673 9710 2687 9724
rect 2673 9673 2687 9687
rect 2753 9673 2767 9687
rect 2613 9573 2627 9587
rect 2633 9536 2647 9550
rect 2573 9470 2587 9484
rect 2553 9453 2567 9467
rect 2553 9393 2567 9407
rect 2553 9233 2567 9247
rect 2553 9190 2567 9204
rect 2613 9393 2627 9407
rect 2613 9333 2627 9347
rect 2593 9033 2607 9047
rect 2633 9236 2647 9250
rect 2893 9736 2907 9750
rect 3073 9853 3087 9867
rect 3073 9773 3087 9787
rect 3053 9730 3067 9744
rect 3093 9730 3107 9744
rect 3393 10030 3407 10044
rect 3513 10036 3527 10050
rect 3613 10033 3627 10047
rect 3533 9993 3547 10007
rect 3233 9753 3247 9767
rect 3293 9756 3307 9770
rect 3073 9713 3087 9727
rect 3153 9713 3167 9727
rect 2813 9633 2827 9647
rect 2993 9633 3007 9647
rect 2653 9233 2667 9247
rect 2693 9236 2707 9250
rect 2733 9236 2747 9250
rect 2773 9236 2787 9250
rect 2673 9190 2687 9204
rect 2713 9190 2727 9204
rect 2773 9153 2787 9167
rect 2633 9133 2647 9147
rect 2673 9093 2687 9107
rect 2613 8971 2627 8985
rect 2753 9055 2767 9069
rect 2793 9017 2807 9031
rect 2693 8971 2707 8985
rect 2593 8873 2607 8887
rect 2633 8773 2647 8787
rect 2533 8672 2547 8686
rect 2513 8653 2527 8667
rect 2533 8533 2547 8547
rect 2533 8493 2547 8507
rect 2733 8773 2747 8787
rect 2713 8613 2727 8627
rect 2893 9593 2907 9607
rect 2853 9573 2867 9587
rect 2933 9536 2947 9550
rect 2853 9273 2867 9287
rect 2833 9193 2847 9207
rect 2833 9053 2847 9067
rect 2833 9013 2847 9027
rect 2833 8753 2847 8767
rect 2813 8633 2827 8647
rect 2833 8533 2847 8547
rect 2733 8513 2747 8527
rect 2753 8496 2767 8510
rect 2653 8450 2667 8464
rect 2693 8450 2707 8464
rect 2733 8450 2747 8464
rect 2553 8430 2567 8444
rect 2533 8353 2547 8367
rect 2553 8313 2567 8327
rect 2493 8273 2507 8287
rect 2833 8273 2847 8287
rect 2513 8233 2527 8247
rect 2553 8233 2567 8247
rect 2413 8213 2427 8227
rect 2473 8196 2487 8210
rect 2552 8170 2566 8184
rect 2573 8176 2587 8190
rect 2673 8176 2687 8190
rect 2453 8113 2467 8127
rect 2953 9490 2967 9504
rect 2913 9453 2927 9467
rect 2973 9333 2987 9347
rect 2913 9253 2927 9267
rect 3013 9553 3027 9567
rect 3013 9490 3027 9504
rect 3113 9613 3127 9627
rect 3093 9593 3107 9607
rect 3093 9493 3107 9507
rect 3073 9333 3087 9347
rect 3053 9273 3067 9287
rect 2993 9253 3007 9267
rect 3013 9236 3027 9250
rect 2953 9190 2967 9204
rect 3053 9153 3067 9167
rect 3013 9016 3027 9030
rect 3093 9073 3107 9087
rect 2913 8953 2927 8967
rect 2893 8873 2907 8887
rect 2873 8833 2887 8847
rect 2933 8853 2947 8867
rect 3033 8953 3047 8967
rect 3153 9593 3167 9607
rect 3293 9593 3307 9607
rect 3133 9533 3147 9547
rect 3213 9536 3227 9550
rect 3413 9833 3427 9847
rect 3373 9756 3387 9770
rect 3513 9773 3527 9787
rect 3393 9710 3407 9724
rect 3553 9953 3567 9967
rect 3533 9693 3547 9707
rect 3613 9893 3627 9907
rect 3673 9893 3687 9907
rect 3593 9756 3607 9770
rect 3593 9713 3607 9727
rect 3553 9633 3567 9647
rect 3513 9613 3527 9627
rect 3873 10473 3887 10487
rect 3833 10250 3847 10264
rect 3813 10192 3827 10206
rect 3853 10056 3867 10070
rect 3993 11093 4007 11107
rect 3993 11053 4007 11067
rect 4073 11050 4087 11064
rect 3973 10953 3987 10967
rect 3953 10893 3967 10907
rect 4013 10933 4027 10947
rect 4013 10796 4027 10810
rect 3973 10753 3987 10767
rect 4033 10750 4047 10764
rect 4273 11753 4287 11767
rect 4313 11693 4327 11707
rect 4373 11693 4387 11707
rect 4353 11653 4367 11667
rect 4333 11570 4347 11584
rect 4293 11553 4307 11567
rect 4253 11533 4267 11547
rect 4273 11493 4287 11507
rect 4633 12136 4647 12150
rect 4713 12173 4727 12187
rect 4613 12090 4627 12104
rect 4573 12053 4587 12067
rect 4973 12110 4987 12124
rect 5093 12116 5107 12130
rect 5173 12113 5187 12127
rect 4653 12013 4667 12027
rect 4773 11953 4787 11967
rect 4713 11893 4727 11907
rect 4713 11856 4727 11870
rect 4753 11856 4767 11870
rect 4553 11816 4567 11830
rect 4653 11816 4667 11830
rect 4653 11773 4667 11787
rect 4493 11693 4507 11707
rect 4413 11616 4427 11630
rect 4233 11353 4247 11367
rect 4133 11316 4147 11330
rect 4373 11453 4387 11467
rect 4353 11433 4367 11447
rect 4333 11353 4347 11367
rect 4273 11316 4287 11330
rect 4253 11270 4267 11284
rect 4253 11233 4267 11247
rect 4293 11233 4307 11247
rect 4173 11096 4187 11110
rect 4213 11096 4227 11110
rect 4153 11050 4167 11064
rect 4333 11213 4347 11227
rect 4293 11096 4307 11110
rect 4253 11033 4267 11047
rect 4193 10993 4207 11007
rect 4333 11093 4347 11107
rect 4293 10973 4307 10987
rect 4193 10893 4207 10907
rect 4113 10713 4127 10727
rect 4173 10653 4187 10667
rect 4293 10796 4307 10810
rect 4393 11273 4407 11287
rect 4533 11616 4547 11630
rect 4573 11616 4587 11630
rect 4493 11573 4507 11587
rect 4433 11473 4447 11487
rect 4593 11570 4607 11584
rect 4573 11533 4587 11547
rect 4553 11493 4567 11507
rect 4533 11353 4547 11367
rect 4493 11333 4507 11347
rect 4713 11653 4727 11667
rect 4693 11473 4707 11487
rect 4673 11413 4687 11427
rect 4693 11393 4707 11407
rect 4673 11373 4687 11387
rect 4733 11613 4747 11627
rect 4773 11713 4787 11727
rect 4973 12013 4987 12027
rect 5133 11973 5147 11987
rect 5333 11973 5347 11987
rect 4973 11913 4987 11927
rect 5273 11913 5287 11927
rect 5133 11853 5147 11867
rect 5013 11836 5027 11850
rect 5053 11836 5067 11850
rect 5173 11836 5187 11850
rect 4893 11790 4907 11804
rect 4953 11790 4967 11804
rect 4853 11733 4867 11747
rect 4793 11653 4807 11667
rect 4793 11616 4807 11630
rect 4933 11773 4947 11787
rect 5153 11793 5167 11807
rect 9053 12213 9067 12227
rect 9833 12213 9847 12227
rect 9373 12193 9387 12207
rect 6033 12173 6047 12187
rect 6213 12173 6227 12187
rect 8553 12173 8567 12187
rect 9053 12173 9067 12187
rect 5773 12136 5787 12150
rect 5892 12133 5906 12147
rect 5913 12136 5927 12150
rect 6073 12136 6087 12150
rect 6673 12153 6687 12167
rect 6753 12153 6767 12167
rect 5753 12073 5767 12087
rect 5433 12033 5447 12047
rect 5513 12033 5527 12047
rect 5893 12090 5907 12104
rect 5833 12033 5847 12047
rect 5793 11973 5807 11987
rect 5753 11913 5767 11927
rect 5373 11873 5387 11887
rect 5653 11873 5667 11887
rect 5233 11836 5247 11850
rect 5273 11836 5287 11850
rect 5353 11813 5367 11827
rect 5193 11773 5207 11787
rect 5173 11753 5187 11767
rect 5153 11733 5167 11747
rect 5493 11816 5507 11830
rect 6233 12133 6247 12147
rect 6113 12116 6127 12130
rect 6173 12116 6187 12130
rect 6213 12116 6227 12130
rect 6013 12090 6027 12104
rect 6373 12110 6387 12124
rect 6493 12116 6507 12130
rect 6053 12073 6067 12087
rect 6133 12073 6147 12087
rect 6213 12073 6227 12087
rect 6053 12013 6067 12027
rect 6533 12053 6547 12067
rect 6213 11993 6227 12007
rect 6333 11993 6347 12007
rect 6133 11973 6147 11987
rect 6233 11933 6247 11947
rect 5913 11913 5927 11927
rect 5833 11853 5847 11867
rect 5653 11810 5667 11824
rect 5693 11810 5707 11824
rect 5373 11773 5387 11787
rect 5353 11673 5367 11687
rect 5493 11673 5507 11687
rect 5293 11653 5307 11667
rect 4893 11616 4907 11630
rect 4773 11593 4787 11607
rect 4973 11596 4987 11610
rect 5093 11590 5107 11604
rect 5253 11590 5267 11604
rect 5393 11616 5407 11630
rect 4793 11513 4807 11527
rect 4753 11453 4767 11467
rect 4933 11453 4947 11467
rect 5053 11453 5067 11467
rect 4873 11393 4887 11407
rect 5313 11433 5327 11447
rect 5173 11413 5187 11427
rect 5253 11413 5267 11427
rect 5053 11336 5067 11350
rect 4573 11316 4587 11330
rect 4613 11293 4627 11307
rect 4513 11270 4527 11284
rect 4413 11233 4427 11247
rect 4453 11233 4467 11247
rect 4453 11096 4467 11110
rect 4493 11053 4507 11067
rect 4433 11033 4447 11047
rect 4493 10993 4507 11007
rect 4553 11233 4567 11247
rect 4533 11193 4547 11207
rect 4613 11193 4627 11207
rect 4693 11290 4707 11304
rect 4733 11290 4747 11304
rect 4893 11296 4907 11310
rect 5113 11336 5127 11350
rect 5013 11290 5027 11304
rect 5093 11293 5107 11307
rect 5013 11253 5027 11267
rect 4913 11193 4927 11207
rect 5073 11213 5087 11227
rect 4713 11133 4727 11147
rect 4873 11133 4887 11147
rect 4753 11096 4767 11110
rect 4793 11096 4807 11110
rect 4733 11050 4747 11064
rect 4533 11013 4547 11027
rect 4893 11096 4907 11110
rect 4793 10973 4807 10987
rect 4853 10953 4867 10967
rect 4513 10933 4527 10947
rect 4693 10913 4707 10927
rect 4433 10893 4447 10907
rect 4393 10773 4407 10787
rect 4193 10633 4207 10647
rect 4253 10593 4267 10607
rect 4073 10550 4087 10564
rect 4193 10556 4207 10570
rect 4313 10750 4327 10764
rect 4293 10713 4307 10727
rect 4393 10713 4407 10727
rect 4533 10776 4547 10790
rect 4753 10776 4767 10790
rect 4693 10750 4707 10764
rect 4493 10673 4507 10687
rect 4353 10553 4367 10567
rect 4273 10473 4287 10487
rect 3933 10413 3947 10427
rect 4073 10413 4087 10427
rect 4233 10413 4247 10427
rect 3973 10393 3987 10407
rect 3953 10373 3967 10387
rect 3913 10333 3927 10347
rect 3893 10313 3907 10327
rect 3693 9833 3707 9847
rect 3753 9833 3767 9847
rect 3693 9773 3707 9787
rect 3653 9756 3667 9770
rect 3673 9693 3687 9707
rect 3713 9693 3727 9707
rect 3753 9693 3767 9707
rect 3753 9633 3767 9647
rect 3613 9593 3627 9607
rect 3433 9510 3447 9524
rect 3693 9516 3707 9530
rect 3733 9516 3747 9530
rect 3193 9490 3207 9504
rect 3153 9453 3167 9467
rect 3233 9453 3247 9467
rect 3153 9413 3167 9427
rect 3193 9413 3207 9427
rect 3133 9013 3147 9027
rect 3053 8933 3067 8947
rect 3113 8933 3127 8947
rect 2973 8715 2987 8729
rect 2913 8670 2927 8684
rect 2933 8653 2947 8667
rect 3053 8653 3067 8667
rect 2913 8633 2927 8647
rect 2893 8413 2907 8427
rect 2873 8333 2887 8347
rect 2913 8393 2927 8407
rect 3033 8573 3047 8587
rect 3033 8513 3047 8527
rect 3013 8496 3027 8510
rect 3193 9373 3207 9387
rect 3173 9333 3187 9347
rect 3273 9470 3287 9484
rect 3313 9453 3327 9467
rect 3313 9413 3327 9427
rect 3713 9413 3727 9427
rect 3413 9393 3427 9407
rect 3253 9333 3267 9347
rect 3433 9353 3447 9367
rect 3413 9253 3427 9267
rect 3273 9236 3287 9250
rect 3252 9153 3266 9167
rect 3273 9153 3287 9167
rect 3333 9153 3347 9167
rect 3333 9016 3347 9030
rect 3273 8973 3287 8987
rect 3353 8970 3367 8984
rect 3413 9213 3427 9227
rect 3413 8933 3427 8947
rect 3313 8873 3327 8887
rect 3193 8853 3207 8867
rect 3173 8813 3187 8827
rect 3153 8773 3167 8787
rect 3733 9333 3747 9347
rect 3793 9993 3807 10007
rect 3833 9893 3847 9907
rect 3793 9773 3807 9787
rect 3793 9673 3807 9687
rect 3793 9533 3807 9547
rect 3773 9453 3787 9467
rect 3793 9413 3807 9427
rect 3813 9353 3827 9367
rect 3753 9313 3767 9327
rect 3713 9273 3727 9287
rect 4013 10333 4027 10347
rect 4097 10313 4111 10327
rect 4073 10296 4087 10310
rect 4092 10253 4106 10267
rect 3933 10233 3947 10247
rect 3893 9893 3907 9907
rect 3873 9853 3887 9867
rect 3973 10193 3987 10207
rect 3953 10133 3967 10147
rect 3973 10056 3987 10070
rect 3953 9953 3967 9967
rect 3933 9913 3947 9927
rect 3953 9853 3967 9867
rect 4033 10230 4047 10244
rect 4113 10250 4127 10264
rect 4233 10256 4247 10270
rect 4413 10572 4427 10586
rect 4453 10576 4467 10590
rect 4633 10633 4647 10647
rect 4613 10593 4627 10607
rect 4553 10573 4567 10587
rect 4413 10393 4427 10407
rect 4513 10530 4527 10544
rect 4553 10530 4567 10544
rect 4473 10373 4487 10387
rect 4413 10256 4427 10270
rect 4393 10193 4407 10207
rect 4433 10213 4447 10227
rect 4413 10173 4427 10187
rect 4093 10133 4107 10147
rect 4593 10433 4607 10447
rect 4553 10373 4567 10387
rect 4533 10213 4547 10227
rect 4493 10113 4507 10127
rect 4093 10073 4107 10087
rect 4493 10073 4507 10087
rect 4013 10056 4027 10070
rect 4053 10056 4067 10070
rect 3993 9993 4007 10007
rect 3993 9853 4007 9867
rect 3973 9833 3987 9847
rect 3933 9756 3947 9770
rect 4213 10036 4227 10050
rect 4333 10030 4347 10044
rect 4033 9953 4047 9967
rect 4073 9953 4087 9967
rect 4013 9793 4027 9807
rect 4073 9913 4087 9927
rect 4133 10013 4147 10027
rect 4173 9933 4187 9947
rect 4113 9893 4127 9907
rect 4593 10233 4607 10247
rect 4553 10073 4567 10087
rect 4533 10036 4547 10050
rect 4593 10036 4607 10050
rect 4513 9993 4527 10007
rect 4553 9993 4567 10007
rect 4493 9853 4507 9867
rect 4353 9793 4367 9807
rect 3993 9756 4007 9770
rect 4053 9736 4067 9750
rect 3873 9713 3887 9727
rect 3913 9673 3927 9687
rect 3953 9673 3967 9687
rect 4053 9673 4067 9687
rect 3953 9536 3967 9550
rect 4013 9533 4027 9547
rect 3873 9353 3887 9367
rect 3453 9253 3467 9267
rect 3733 9253 3747 9267
rect 3833 9253 3847 9267
rect 3593 9216 3607 9230
rect 3713 9193 3727 9207
rect 3453 9173 3467 9187
rect 3473 9073 3487 9087
rect 3633 9073 3647 9087
rect 3133 8715 3147 8729
rect 3373 8715 3387 8729
rect 3233 8669 3247 8683
rect 3193 8613 3207 8627
rect 3373 8593 3387 8607
rect 3373 8553 3387 8567
rect 3353 8513 3367 8527
rect 3213 8470 3227 8484
rect 3513 9016 3527 9030
rect 3553 9016 3567 9030
rect 3593 8970 3607 8984
rect 3513 8953 3527 8967
rect 3553 8953 3567 8967
rect 3433 8715 3447 8729
rect 3473 8716 3487 8730
rect 3453 8670 3467 8684
rect 3533 8813 3547 8827
rect 3413 8573 3427 8587
rect 3513 8573 3527 8587
rect 3413 8533 3427 8547
rect 3513 8513 3527 8527
rect 3473 8493 3487 8507
rect 3053 8430 3067 8444
rect 3353 8433 3367 8447
rect 3033 8393 3047 8407
rect 2933 8373 2947 8387
rect 2993 8373 3007 8387
rect 2893 8313 2907 8327
rect 2853 8213 2867 8227
rect 2973 8213 2987 8227
rect 2913 8153 2927 8167
rect 2833 8133 2847 8147
rect 2873 8133 2887 8147
rect 2553 8093 2567 8107
rect 2453 8073 2467 8087
rect 2413 8033 2427 8047
rect 2433 8013 2447 8027
rect 2393 7953 2407 7967
rect 2433 7953 2447 7967
rect 2773 8013 2787 8027
rect 2833 8013 2847 8027
rect 2473 7993 2487 8007
rect 2473 7950 2487 7964
rect 2573 7950 2587 7964
rect 2833 7956 2847 7970
rect 2873 7956 2887 7970
rect 2213 7873 2227 7887
rect 2193 7493 2207 7507
rect 2053 7410 2067 7424
rect 2153 7410 2167 7424
rect 2193 7410 2207 7424
rect 2353 7930 2367 7944
rect 2413 7910 2427 7924
rect 2793 7873 2807 7887
rect 2313 7813 2327 7827
rect 2653 7813 2667 7827
rect 2433 7793 2447 7807
rect 2313 7675 2327 7689
rect 2553 7753 2567 7767
rect 2393 7493 2407 7507
rect 2453 7495 2467 7509
rect 2373 7457 2387 7471
rect 2253 7410 2267 7424
rect 2233 7333 2247 7347
rect 1993 7273 2007 7287
rect 1973 7253 1987 7267
rect 1793 7133 1807 7147
rect 1953 7133 1967 7147
rect 1773 7113 1787 7127
rect 1893 7110 1907 7124
rect 1853 7073 1867 7087
rect 1913 6993 1927 7007
rect 1752 6933 1766 6947
rect 1773 6936 1787 6950
rect 1833 6936 1847 6950
rect 1873 6936 1887 6950
rect 1893 6890 1907 6904
rect 1853 6873 1867 6887
rect 1853 6813 1867 6827
rect 1993 7136 2007 7150
rect 2093 7136 2107 7150
rect 1993 7093 2007 7107
rect 2173 7033 2187 7047
rect 2033 6973 2047 6987
rect 1993 6773 2007 6787
rect 1893 6753 1907 6767
rect 1873 6673 1887 6687
rect 1913 6636 1927 6650
rect 1973 6636 1987 6650
rect 1833 6573 1847 6587
rect 1773 6433 1787 6447
rect 1873 6573 1887 6587
rect 1853 6553 1867 6567
rect 1933 6593 1947 6607
rect 1913 6513 1927 6527
rect 1893 6473 1907 6487
rect 1813 6333 1827 6347
rect 1873 6332 1887 6346
rect 1773 6313 1787 6327
rect 1813 6173 1827 6187
rect 1833 6153 1847 6167
rect 1753 6132 1767 6146
rect 1793 6116 1807 6130
rect 1773 6070 1787 6084
rect 1813 6033 1827 6047
rect 1793 5973 1807 5987
rect 1753 5813 1767 5827
rect 1913 6233 1927 6247
rect 1893 6116 1907 6130
rect 1893 6073 1907 6087
rect 1913 6053 1927 6067
rect 1893 5973 1907 5987
rect 1873 5953 1887 5967
rect 1873 5850 1887 5864
rect 1853 5773 1867 5787
rect 1793 5713 1807 5727
rect 1793 5613 1807 5627
rect 1913 5633 1927 5647
rect 1733 5433 1747 5447
rect 1713 5413 1727 5427
rect 1733 5376 1747 5390
rect 1813 5550 1827 5564
rect 1873 5553 1887 5567
rect 1853 5413 1867 5427
rect 1833 5376 1847 5390
rect 1753 5330 1767 5344
rect 1753 5273 1767 5287
rect 1793 5253 1807 5267
rect 1853 5330 1867 5344
rect 1812 5233 1826 5247
rect 1833 5233 1847 5247
rect 1693 5193 1707 5207
rect 1613 5173 1627 5187
rect 1593 5153 1607 5167
rect 1613 5113 1627 5127
rect 1573 5096 1587 5110
rect 1433 4993 1447 5007
rect 1413 4973 1427 4987
rect 1393 4933 1407 4947
rect 1493 4973 1507 4987
rect 1473 4893 1487 4907
rect 1393 4793 1407 4807
rect 1433 4793 1447 4807
rect 1353 4753 1367 4767
rect 1293 4713 1307 4727
rect 1253 4633 1267 4647
rect 1413 4633 1427 4647
rect 1113 4593 1127 4607
rect 1553 5033 1567 5047
rect 1573 4933 1587 4947
rect 1733 5056 1747 5070
rect 1653 4953 1667 4967
rect 1613 4873 1627 4887
rect 1593 4853 1607 4867
rect 1773 4933 1787 4947
rect 1733 4873 1747 4887
rect 1513 4733 1527 4747
rect 1513 4653 1527 4667
rect 1493 4613 1507 4627
rect 1093 4573 1107 4587
rect 1413 4573 1427 4587
rect 833 4533 847 4547
rect 1113 4530 1127 4544
rect 1233 4536 1247 4550
rect 693 4513 707 4527
rect 693 4413 707 4427
rect 793 4493 807 4507
rect 833 4493 847 4507
rect 773 4433 787 4447
rect 753 4373 767 4387
rect 1513 4533 1527 4547
rect 1493 4513 1507 4527
rect 1433 4493 1447 4507
rect 1493 4453 1507 4467
rect 1033 4433 1047 4447
rect 1433 4433 1447 4447
rect 873 4373 887 4387
rect 1493 4373 1507 4387
rect 833 4316 847 4330
rect 1373 4333 1387 4347
rect 1413 4336 1427 4350
rect 873 4310 887 4324
rect 1033 4310 1047 4324
rect 1153 4316 1167 4330
rect 1233 4313 1247 4327
rect 713 4290 727 4304
rect 1133 4193 1147 4207
rect 653 4153 667 4167
rect 813 4153 827 4167
rect 753 4093 767 4107
rect 713 4053 727 4067
rect 653 4013 667 4027
rect 852 4010 866 4024
rect 873 4016 887 4030
rect 973 4016 987 4030
rect 693 3953 707 3967
rect 733 3953 747 3967
rect 853 3953 867 3967
rect 1193 4153 1207 4167
rect 1433 4290 1447 4304
rect 1393 4093 1407 4107
rect 1373 4053 1387 4067
rect 1233 4010 1247 4024
rect 1373 4010 1387 4024
rect 1173 3913 1187 3927
rect 633 3893 647 3907
rect 693 3893 707 3907
rect 1133 3893 1147 3907
rect 613 3833 627 3847
rect 453 3813 467 3827
rect 513 3816 527 3830
rect 573 3796 587 3810
rect 1553 4713 1567 4727
rect 1533 4373 1547 4387
rect 1493 4193 1507 4207
rect 1453 4053 1467 4067
rect 1533 4053 1547 4067
rect 1393 3993 1407 4007
rect 1473 3990 1487 4004
rect 1533 3973 1547 3987
rect 1573 4633 1587 4647
rect 1553 3953 1567 3967
rect 1413 3933 1427 3947
rect 1513 3933 1527 3947
rect 1413 3893 1427 3907
rect 1393 3873 1407 3887
rect 673 3833 687 3847
rect 533 3770 547 3784
rect 653 3753 667 3767
rect 533 3573 547 3587
rect 453 3533 467 3547
rect 553 3533 567 3547
rect 513 3516 527 3530
rect 493 3470 507 3484
rect 533 3470 547 3484
rect 513 3453 527 3467
rect 473 3373 487 3387
rect 653 3473 667 3487
rect 573 3433 587 3447
rect 553 3293 567 3307
rect 453 3250 467 3264
rect 493 3250 507 3264
rect 553 3250 567 3264
rect 693 3790 707 3804
rect 833 3790 847 3804
rect 953 3796 967 3810
rect 1093 3796 1107 3810
rect 1213 3790 1227 3804
rect 693 3753 707 3767
rect 993 3750 1007 3764
rect 1053 3750 1067 3764
rect 969 3733 983 3747
rect 773 3573 787 3587
rect 733 3533 747 3547
rect 813 3516 827 3530
rect 793 3470 807 3484
rect 833 3393 847 3407
rect 773 3296 787 3310
rect 1077 3733 1091 3747
rect 1433 3853 1447 3867
rect 1433 3790 1447 3804
rect 1493 3793 1507 3807
rect 1333 3573 1347 3587
rect 1373 3573 1387 3587
rect 1013 3516 1027 3530
rect 1053 3516 1067 3530
rect 1133 3516 1147 3530
rect 1173 3516 1187 3530
rect 1013 3473 1027 3487
rect 1173 3473 1187 3487
rect 1113 3433 1127 3447
rect 1073 3393 1087 3407
rect 993 3353 1007 3367
rect 1153 3353 1167 3367
rect 933 3333 947 3347
rect 1073 3333 1087 3347
rect 793 3250 807 3264
rect 833 3250 847 3264
rect 753 3213 767 3227
rect 393 2993 407 3007
rect 453 2996 467 3010
rect 573 2996 587 3010
rect 513 2973 527 2987
rect 393 2950 407 2964
rect 433 2950 447 2964
rect 453 2893 467 2907
rect 513 2893 527 2907
rect 513 2776 527 2790
rect 453 2730 467 2744
rect 493 2730 507 2744
rect 533 2730 547 2744
rect 553 2693 567 2707
rect 553 2653 567 2667
rect 533 2633 547 2647
rect 433 2533 447 2547
rect 493 2476 507 2490
rect 393 2253 407 2267
rect 513 2256 527 2270
rect 613 2473 627 2487
rect 453 2210 467 2224
rect 573 2210 587 2224
rect 613 2193 627 2207
rect 533 2173 547 2187
rect 593 2173 607 2187
rect 533 2133 547 2147
rect 493 2093 507 2107
rect 493 1993 507 2007
rect 393 1956 407 1970
rect 593 2093 607 2107
rect 573 1993 587 2007
rect 373 1853 387 1867
rect 553 1853 567 1867
rect 513 1793 527 1807
rect 493 1753 507 1767
rect 873 3033 887 3047
rect 753 2996 767 3010
rect 893 2993 907 3007
rect 733 2950 747 2964
rect 873 2953 887 2967
rect 1033 3296 1047 3310
rect 1053 3213 1067 3227
rect 1093 3113 1107 3127
rect 993 2996 1007 3010
rect 893 2933 907 2947
rect 773 2813 787 2827
rect 673 2773 687 2787
rect 713 2773 727 2787
rect 813 2533 827 2547
rect 733 2430 747 2444
rect 673 2293 687 2307
rect 653 2253 667 2267
rect 633 1910 647 1924
rect 593 1873 607 1887
rect 573 1793 587 1807
rect 513 1690 527 1704
rect 553 1693 567 1707
rect 353 1653 367 1667
rect 333 1435 347 1449
rect 193 1216 207 1230
rect 153 1173 167 1187
rect 213 1170 227 1184
rect 333 1216 347 1230
rect 333 1153 347 1167
rect 33 1073 47 1087
rect 57 933 71 947
rect 73 890 87 904
rect 193 896 207 910
rect 493 1493 507 1507
rect 613 1493 627 1507
rect 433 1253 447 1267
rect 433 1213 447 1227
rect 513 1253 527 1267
rect 513 1216 527 1230
rect 553 1216 567 1230
rect 453 1170 467 1184
rect 413 1133 427 1147
rect 493 1133 507 1147
rect 513 1073 527 1087
rect 373 933 387 947
rect 453 890 467 904
rect 353 873 367 887
rect 393 873 407 887
rect 73 676 87 690
rect 193 670 207 684
rect 57 633 71 647
rect 33 593 47 607
rect 373 733 387 747
rect 373 693 387 707
rect 453 693 467 707
rect 633 1033 647 1047
rect 613 890 627 904
rect 553 833 567 847
rect 933 2950 947 2964
rect 1013 2950 1027 2964
rect 933 2893 947 2907
rect 973 2893 987 2907
rect 913 2730 927 2744
rect 993 2813 1007 2827
rect 1033 2776 1047 2790
rect 1073 2773 1087 2787
rect 973 2730 987 2744
rect 893 2493 907 2507
rect 913 2476 927 2490
rect 993 2476 1007 2490
rect 1053 2476 1067 2490
rect 913 2433 927 2447
rect 1013 2430 1027 2444
rect 1053 2433 1067 2447
rect 1133 2713 1147 2727
rect 973 2413 987 2427
rect 1073 2413 1087 2427
rect 853 2293 867 2307
rect 813 2256 827 2270
rect 793 2210 807 2224
rect 833 2210 847 2224
rect 873 2133 887 2147
rect 1233 3293 1247 3307
rect 1373 3516 1387 3530
rect 1433 3516 1447 3530
rect 1353 3470 1367 3484
rect 1293 3433 1307 3447
rect 1353 3373 1367 3387
rect 1393 3333 1407 3347
rect 1653 4793 1667 4807
rect 1633 4753 1647 4767
rect 1613 4593 1627 4607
rect 1593 4513 1607 4527
rect 1593 4393 1607 4407
rect 1673 4773 1687 4787
rect 1653 4733 1667 4747
rect 1653 4693 1667 4707
rect 1633 4533 1647 4547
rect 1673 4673 1687 4687
rect 1873 4913 1887 4927
rect 1833 4893 1847 4907
rect 1913 5553 1927 5567
rect 1953 6373 1967 6387
rect 1993 6533 2007 6547
rect 1993 6273 2007 6287
rect 1973 6233 1987 6247
rect 1993 6116 2007 6130
rect 1973 6013 1987 6027
rect 1953 5773 1967 5787
rect 1953 5333 1967 5347
rect 1993 5633 2007 5647
rect 2093 6936 2107 6950
rect 2133 6936 2147 6950
rect 2213 6936 2227 6950
rect 2193 6890 2207 6904
rect 2233 6890 2247 6904
rect 2153 6873 2167 6887
rect 2093 6813 2107 6827
rect 2153 6713 2167 6727
rect 2153 6673 2167 6687
rect 2193 6653 2207 6667
rect 2153 6636 2167 6650
rect 2093 6593 2107 6607
rect 2133 6590 2147 6604
rect 2033 6573 2047 6587
rect 2133 6573 2147 6587
rect 2173 6533 2187 6547
rect 2113 6453 2127 6467
rect 2153 6453 2167 6467
rect 2053 6173 2067 6187
rect 2053 6116 2067 6130
rect 2093 6116 2107 6130
rect 2073 6070 2087 6084
rect 2173 6393 2187 6407
rect 2153 6013 2167 6027
rect 2293 6993 2307 7007
rect 2293 6893 2307 6907
rect 2273 6653 2287 6667
rect 2253 6513 2267 6527
rect 2273 6493 2287 6507
rect 2273 6273 2287 6287
rect 2233 6233 2247 6247
rect 2273 6070 2287 6084
rect 2113 5993 2127 6007
rect 2173 5993 2187 6007
rect 2153 5896 2167 5910
rect 2133 5850 2147 5864
rect 2173 5813 2187 5827
rect 2193 5793 2207 5807
rect 2173 5713 2187 5727
rect 2133 5633 2147 5647
rect 2173 5633 2187 5647
rect 2033 5613 2047 5627
rect 2093 5596 2107 5610
rect 2173 5596 2187 5610
rect 2073 5550 2087 5564
rect 2073 5493 2087 5507
rect 2033 5473 2047 5487
rect 2033 5376 2047 5390
rect 2113 5473 2127 5487
rect 2373 7093 2387 7107
rect 2353 7073 2367 7087
rect 2313 6853 2327 6867
rect 2333 6673 2347 6687
rect 2333 6590 2347 6604
rect 2352 6453 2366 6467
rect 2373 6453 2387 6467
rect 2333 6273 2347 6287
rect 2413 7457 2427 7471
rect 2433 7333 2447 7347
rect 2473 7153 2487 7167
rect 2433 7013 2447 7027
rect 2613 7713 2627 7727
rect 2693 7676 2707 7690
rect 2773 7676 2787 7690
rect 2673 7630 2687 7644
rect 2633 7553 2647 7567
rect 2633 7456 2647 7470
rect 2713 7456 2727 7470
rect 2753 7456 2767 7470
rect 2553 7233 2567 7247
rect 2593 7213 2607 7227
rect 2553 7153 2567 7167
rect 2573 7093 2587 7107
rect 2533 7033 2547 7047
rect 2593 7013 2607 7027
rect 2573 6936 2587 6950
rect 2453 6873 2467 6887
rect 2533 6793 2547 6807
rect 2513 6773 2527 6787
rect 2493 6733 2507 6747
rect 2433 6636 2447 6650
rect 2493 6593 2507 6607
rect 2453 6573 2467 6587
rect 2513 6573 2527 6587
rect 2393 6353 2407 6367
rect 2473 6333 2487 6347
rect 2533 6333 2547 6347
rect 2413 6116 2427 6130
rect 2333 6033 2347 6047
rect 2513 6273 2527 6287
rect 2493 6153 2507 6167
rect 2473 6033 2487 6047
rect 2393 5896 2407 5910
rect 2433 5896 2447 5910
rect 2413 5850 2427 5864
rect 2293 5833 2307 5847
rect 2273 5773 2287 5787
rect 2313 5773 2327 5787
rect 2453 5733 2467 5747
rect 2453 5693 2467 5707
rect 2313 5673 2327 5687
rect 2353 5673 2367 5687
rect 2213 5573 2227 5587
rect 2393 5613 2407 5627
rect 2253 5553 2267 5567
rect 2373 5550 2387 5564
rect 2453 5553 2467 5567
rect 2213 5493 2227 5507
rect 2473 5413 2487 5427
rect 2453 5393 2467 5407
rect 2193 5373 2207 5387
rect 2313 5350 2327 5364
rect 2453 5350 2467 5364
rect 2013 5333 2027 5347
rect 1993 5233 2007 5247
rect 1933 5153 1947 5167
rect 2053 5330 2067 5344
rect 2053 5293 2067 5307
rect 2033 5113 2047 5127
rect 1933 5050 1947 5064
rect 2033 5050 2047 5064
rect 1993 5013 2007 5027
rect 1933 4993 1947 5007
rect 1973 4913 1987 4927
rect 1953 4810 1967 4824
rect 2013 4773 2027 4787
rect 1913 4753 1927 4767
rect 2113 5213 2127 5227
rect 2093 5173 2107 5187
rect 2093 5152 2107 5166
rect 2073 4810 2087 4824
rect 2453 5313 2467 5327
rect 2333 5253 2347 5267
rect 2153 5233 2167 5247
rect 2133 5193 2147 5207
rect 2113 4953 2127 4967
rect 2273 5193 2287 5207
rect 2153 5033 2167 5047
rect 2193 5073 2207 5087
rect 2233 5076 2247 5090
rect 2133 4893 2147 4907
rect 2173 4893 2187 4907
rect 2253 5030 2267 5044
rect 2293 4953 2307 4967
rect 2213 4933 2227 4947
rect 2193 4873 2207 4887
rect 2293 4873 2307 4887
rect 2193 4810 2207 4824
rect 2093 4713 2107 4727
rect 2053 4673 2067 4687
rect 2153 4673 2167 4687
rect 1873 4593 1887 4607
rect 1853 4536 1867 4550
rect 1993 4536 2007 4550
rect 1733 4413 1747 4427
rect 1693 4393 1707 4407
rect 1653 4353 1667 4367
rect 1833 4473 1847 4487
rect 1773 4373 1787 4387
rect 1753 4353 1767 4367
rect 1613 4293 1627 4307
rect 1673 4290 1687 4304
rect 1633 4036 1647 4050
rect 1593 4016 1607 4030
rect 1533 3453 1547 3467
rect 1513 3333 1527 3347
rect 1633 3816 1647 3830
rect 1573 3793 1587 3807
rect 1733 4273 1747 4287
rect 1673 4253 1687 4267
rect 1713 4253 1727 4267
rect 1873 4513 1887 4527
rect 1853 4413 1867 4427
rect 1693 4233 1707 4247
rect 1753 4233 1767 4247
rect 1833 4153 1847 4167
rect 1813 4113 1827 4127
rect 1773 4053 1787 4067
rect 1813 4053 1827 4067
rect 1893 4493 1907 4507
rect 1973 4413 1987 4427
rect 2133 4413 2147 4427
rect 1933 4336 1947 4350
rect 2033 4333 2047 4347
rect 1993 4290 2007 4304
rect 1953 4253 1967 4267
rect 2033 4253 2047 4267
rect 1953 4173 1967 4187
rect 2133 4153 2147 4167
rect 1873 4093 1887 4107
rect 2133 4053 2147 4067
rect 1733 4036 1747 4050
rect 1693 3993 1707 4007
rect 1673 3933 1687 3947
rect 1733 3933 1747 3947
rect 1693 3816 1707 3830
rect 1793 3990 1807 4004
rect 1833 3993 1847 4007
rect 1993 4016 2007 4030
rect 1753 3853 1767 3867
rect 1653 3773 1667 3787
rect 1713 3770 1727 3784
rect 1753 3770 1767 3784
rect 1633 3693 1647 3707
rect 1753 3733 1767 3747
rect 1733 3693 1747 3707
rect 1613 3593 1627 3607
rect 1713 3593 1727 3607
rect 1573 3513 1587 3527
rect 1653 3516 1667 3530
rect 1693 3516 1707 3530
rect 1693 3473 1707 3487
rect 1633 3453 1647 3467
rect 1673 3413 1687 3427
rect 1593 3373 1607 3387
rect 1553 3293 1567 3307
rect 1613 3296 1627 3310
rect 1293 3250 1307 3264
rect 1333 3250 1347 3264
rect 1433 3253 1447 3267
rect 1653 3250 1667 3264
rect 1373 3213 1387 3227
rect 1633 3213 1647 3227
rect 1273 3053 1287 3067
rect 1273 3032 1287 3046
rect 1213 2933 1227 2947
rect 1193 2893 1207 2907
rect 1173 2673 1187 2687
rect 1153 2613 1167 2627
rect 1153 2313 1167 2327
rect 1133 2273 1147 2287
rect 1093 2256 1107 2270
rect 1073 2193 1087 2207
rect 1113 2193 1127 2207
rect 973 2053 987 2067
rect 693 1993 707 2007
rect 773 1993 787 2007
rect 673 1793 687 1807
rect 673 1753 687 1767
rect 673 1493 687 1507
rect 833 1976 847 1990
rect 1173 2193 1187 2207
rect 1293 2950 1307 2964
rect 1253 2873 1267 2887
rect 1353 2833 1367 2847
rect 1233 2813 1247 2827
rect 1253 2793 1267 2807
rect 1313 2730 1327 2744
rect 1353 2730 1367 2744
rect 1513 3053 1527 3067
rect 1553 2996 1567 3010
rect 1533 2893 1547 2907
rect 1393 2793 1407 2807
rect 1553 2793 1567 2807
rect 1273 2713 1287 2727
rect 1373 2713 1387 2727
rect 1573 2730 1587 2744
rect 1653 2673 1667 2687
rect 1353 2613 1367 2627
rect 1653 2593 1667 2607
rect 1253 2476 1267 2490
rect 1653 2493 1667 2507
rect 1213 2453 1227 2467
rect 1373 2453 1387 2467
rect 1513 2456 1527 2470
rect 1393 2433 1407 2447
rect 1313 2413 1327 2427
rect 1373 2413 1387 2427
rect 1273 2373 1287 2387
rect 1653 2413 1667 2427
rect 1393 2373 1407 2387
rect 1513 2293 1527 2307
rect 1613 2293 1627 2307
rect 1353 2273 1367 2287
rect 1433 2273 1447 2287
rect 1413 2256 1427 2270
rect 1373 2193 1387 2207
rect 1313 2173 1327 2187
rect 1293 2133 1307 2147
rect 1193 1993 1207 2007
rect 733 1910 747 1924
rect 753 1873 767 1887
rect 813 1853 827 1867
rect 773 1673 787 1687
rect 813 1673 827 1687
rect 993 1936 1007 1950
rect 1153 1936 1167 1950
rect 993 1833 1007 1847
rect 913 1753 927 1767
rect 893 1493 907 1507
rect 753 1435 767 1449
rect 853 1389 867 1403
rect 773 1353 787 1367
rect 693 1313 707 1327
rect 713 1213 727 1227
rect 813 1213 827 1227
rect 693 1113 707 1127
rect 1033 1793 1047 1807
rect 973 1473 987 1487
rect 913 1435 927 1449
rect 893 1389 907 1403
rect 993 1373 1007 1387
rect 973 1353 987 1367
rect 1253 1930 1267 1944
rect 1373 2073 1387 2087
rect 1353 2053 1367 2067
rect 1313 1930 1327 1944
rect 1293 1833 1307 1847
rect 1293 1753 1307 1767
rect 1273 1690 1287 1704
rect 1313 1690 1327 1704
rect 1193 1653 1207 1667
rect 1093 1493 1107 1507
rect 1133 1493 1147 1507
rect 1113 1473 1127 1487
rect 1073 1436 1087 1450
rect 1173 1436 1187 1450
rect 1053 1373 1067 1387
rect 1073 1353 1087 1367
rect 993 1313 1007 1327
rect 1133 1353 1147 1367
rect 1173 1333 1187 1347
rect 1093 1293 1107 1307
rect 993 1190 1007 1204
rect 1213 1493 1227 1507
rect 1273 1473 1287 1487
rect 1273 1373 1287 1387
rect 1213 1353 1227 1367
rect 1253 1196 1267 1210
rect 753 1153 767 1167
rect 793 1113 807 1127
rect 1313 1493 1327 1507
rect 1253 1113 1267 1127
rect 1293 1113 1307 1127
rect 833 1073 847 1087
rect 993 953 1007 967
rect 693 916 707 930
rect 1053 913 1067 927
rect 1373 1993 1387 2007
rect 1393 1853 1407 1867
rect 1433 2210 1447 2224
rect 1573 2256 1587 2270
rect 1733 3373 1747 3387
rect 1733 3333 1747 3347
rect 1793 3573 1807 3587
rect 2133 3993 2147 4007
rect 1873 3953 1887 3967
rect 2013 3913 2027 3927
rect 1953 3816 1967 3830
rect 1873 3733 1887 3747
rect 1913 3733 1927 3747
rect 1913 3633 1927 3647
rect 1893 3613 1907 3627
rect 1873 3470 1887 3484
rect 1813 3413 1827 3427
rect 1773 3293 1787 3307
rect 1873 3296 1887 3310
rect 1753 3153 1767 3167
rect 1733 3113 1747 3127
rect 1853 3250 1867 3264
rect 1893 3213 1907 3227
rect 1893 3153 1907 3167
rect 1893 3093 1907 3107
rect 1813 2996 1827 3010
rect 1853 2996 1867 3010
rect 1733 2950 1747 2964
rect 1793 2950 1807 2964
rect 1793 2913 1807 2927
rect 1833 2893 1847 2907
rect 1833 2833 1847 2847
rect 1693 2673 1707 2687
rect 1773 2730 1787 2744
rect 1973 3773 1987 3787
rect 1953 2793 1967 2807
rect 1893 2653 1907 2667
rect 1833 2613 1847 2627
rect 1813 2593 1827 2607
rect 1693 2493 1707 2507
rect 1753 2493 1767 2507
rect 2073 3653 2087 3667
rect 2013 3633 2027 3647
rect 1993 3470 2007 3484
rect 1993 2773 2007 2787
rect 1993 2633 2007 2647
rect 1973 2593 1987 2607
rect 2233 4773 2247 4787
rect 2193 4593 2207 4607
rect 2173 4533 2187 4547
rect 2253 4493 2267 4507
rect 2193 4433 2207 4447
rect 2313 4713 2327 4727
rect 2293 4413 2307 4427
rect 2273 4373 2287 4387
rect 2233 4336 2247 4350
rect 2193 4073 2207 4087
rect 2293 4253 2307 4267
rect 2293 4153 2307 4167
rect 2173 4053 2187 4067
rect 2193 4010 2207 4024
rect 2253 4010 2267 4024
rect 2173 3893 2187 3907
rect 2153 3633 2167 3647
rect 2213 3833 2227 3847
rect 2213 3816 2227 3830
rect 2293 3893 2307 3907
rect 2313 3833 2327 3847
rect 2313 3793 2327 3807
rect 2233 3770 2247 3784
rect 2273 3753 2287 3767
rect 2193 3693 2207 3707
rect 2173 3533 2187 3547
rect 2153 3516 2167 3530
rect 2233 3533 2247 3547
rect 2133 3433 2147 3447
rect 2213 3433 2227 3447
rect 2153 3353 2167 3367
rect 2173 3353 2187 3367
rect 2113 3313 2127 3327
rect 2133 3250 2147 3264
rect 2213 3250 2227 3264
rect 2193 3193 2207 3207
rect 2173 3173 2187 3187
rect 2113 2996 2127 3010
rect 2173 2893 2187 2907
rect 2093 2833 2107 2847
rect 2153 2833 2167 2847
rect 2053 2776 2067 2790
rect 2173 2813 2187 2827
rect 2173 2773 2187 2787
rect 2213 3053 2227 3067
rect 2113 2713 2127 2727
rect 2193 2713 2207 2727
rect 2013 2553 2027 2567
rect 2213 2533 2227 2547
rect 2253 3516 2267 3530
rect 2253 3413 2267 3427
rect 2253 3353 2267 3367
rect 2293 3016 2307 3030
rect 2413 5213 2427 5227
rect 2373 5013 2387 5027
rect 2353 4893 2367 4907
rect 2353 4533 2367 4547
rect 2353 4493 2367 4507
rect 2533 6113 2547 6127
rect 2613 6636 2627 6650
rect 2613 6373 2627 6387
rect 2573 6313 2587 6327
rect 2733 7393 2747 7407
rect 2773 7393 2787 7407
rect 2713 7313 2727 7327
rect 2673 7193 2687 7207
rect 2653 7153 2667 7167
rect 2653 7093 2667 7107
rect 2673 7073 2687 7087
rect 2673 6973 2687 6987
rect 2773 7233 2787 7247
rect 2693 6873 2707 6887
rect 2733 6733 2747 6747
rect 2713 6713 2727 6727
rect 2753 6713 2767 6727
rect 2693 6636 2707 6650
rect 2933 8033 2947 8047
rect 2913 7793 2927 7807
rect 3013 8313 3027 8327
rect 2993 7813 3007 7827
rect 3113 8333 3127 8347
rect 3033 8153 3047 8167
rect 3053 8053 3067 8067
rect 3073 7930 3087 7944
rect 3013 7773 3027 7787
rect 2973 7753 2987 7767
rect 2933 7676 2947 7690
rect 3013 7673 3027 7687
rect 2873 7653 2887 7667
rect 2953 7630 2967 7644
rect 2873 7593 2887 7607
rect 2933 7593 2947 7607
rect 2813 7155 2827 7169
rect 2913 7109 2927 7123
rect 2973 7456 2987 7470
rect 3053 7629 3067 7643
rect 2993 7410 3007 7424
rect 2993 7373 3007 7387
rect 2973 7313 2987 7327
rect 2933 7073 2947 7087
rect 2873 7033 2887 7047
rect 2933 7033 2947 7047
rect 2913 7013 2927 7027
rect 2853 6973 2867 6987
rect 2793 6693 2807 6707
rect 2873 6953 2887 6967
rect 2853 6673 2867 6687
rect 2773 6613 2787 6627
rect 2673 6590 2687 6604
rect 2793 6593 2807 6607
rect 3033 7273 3047 7287
rect 2993 7213 3007 7227
rect 2973 7013 2987 7027
rect 3013 7133 3027 7147
rect 3033 7113 3047 7127
rect 3013 6993 3027 7007
rect 3173 8293 3187 8307
rect 3133 8253 3147 8267
rect 3113 7633 3127 7647
rect 3093 7456 3107 7470
rect 3093 7413 3107 7427
rect 3213 8196 3227 8210
rect 3233 8150 3247 8164
rect 3193 8053 3207 8067
rect 3173 8013 3187 8027
rect 3333 8013 3347 8027
rect 3153 7976 3167 7990
rect 3293 7976 3307 7990
rect 3173 7933 3187 7947
rect 3313 7893 3327 7907
rect 3313 7713 3327 7727
rect 3293 7675 3307 7689
rect 3193 7629 3207 7643
rect 3153 7553 3167 7567
rect 3253 7410 3267 7424
rect 3133 7313 3147 7327
rect 3073 7273 3087 7287
rect 3053 6953 3067 6967
rect 2953 6937 2967 6951
rect 2933 6893 2947 6907
rect 3053 6891 3067 6905
rect 2993 6753 3007 6767
rect 2953 6636 2967 6650
rect 3033 6636 3047 6650
rect 2793 6553 2807 6567
rect 2733 6453 2747 6467
rect 2693 6433 2707 6447
rect 2713 6370 2727 6384
rect 2753 6313 2767 6327
rect 2653 6253 2667 6267
rect 2673 6213 2687 6227
rect 2632 6153 2646 6167
rect 2653 6153 2667 6167
rect 2673 6133 2687 6147
rect 2813 6533 2827 6547
rect 2833 6416 2847 6430
rect 2793 6293 2807 6307
rect 2813 6213 2827 6227
rect 2813 6173 2827 6187
rect 2753 6093 2767 6107
rect 2593 6070 2607 6084
rect 2573 5896 2587 5910
rect 2553 5813 2567 5827
rect 2753 6033 2767 6047
rect 2713 5993 2727 6007
rect 2713 5913 2727 5927
rect 2693 5896 2707 5910
rect 2633 5850 2647 5864
rect 2713 5833 2727 5847
rect 2693 5813 2707 5827
rect 2673 5773 2687 5787
rect 2573 5713 2587 5727
rect 2673 5673 2687 5687
rect 2673 5596 2687 5610
rect 2613 5550 2627 5564
rect 2693 5553 2707 5567
rect 2653 5533 2667 5547
rect 2573 5453 2587 5467
rect 2533 5373 2547 5387
rect 2513 5356 2527 5370
rect 2673 5413 2687 5427
rect 2613 5373 2627 5387
rect 2653 5373 2667 5387
rect 2493 5313 2507 5327
rect 2473 5193 2487 5207
rect 2513 5173 2527 5187
rect 2433 5073 2447 5087
rect 2493 5073 2507 5087
rect 2573 5076 2587 5090
rect 2413 4633 2427 4647
rect 2393 4593 2407 4607
rect 2373 4473 2387 4487
rect 2373 4333 2387 4347
rect 2373 4290 2387 4304
rect 2353 4273 2367 4287
rect 2533 5030 2547 5044
rect 2593 5030 2607 5044
rect 2573 4993 2587 5007
rect 2493 4856 2507 4870
rect 2512 4813 2526 4827
rect 2533 4810 2547 4824
rect 2473 4753 2487 4767
rect 2473 4713 2487 4727
rect 2433 4573 2447 4587
rect 2493 4573 2507 4587
rect 2593 4813 2607 4827
rect 2573 4693 2587 4707
rect 2433 4533 2447 4547
rect 2433 4493 2447 4507
rect 2413 4473 2427 4487
rect 2393 4133 2407 4147
rect 2373 4113 2387 4127
rect 2353 4012 2367 4026
rect 2373 3933 2387 3947
rect 2373 3912 2387 3926
rect 2353 3793 2367 3807
rect 2393 3770 2407 3784
rect 2373 3713 2387 3727
rect 2433 4453 2447 4467
rect 2513 4510 2527 4524
rect 2593 4510 2607 4524
rect 2553 4453 2567 4467
rect 2473 4393 2487 4407
rect 2533 4336 2547 4350
rect 2513 4273 2527 4287
rect 2533 4193 2547 4207
rect 2473 4073 2487 4087
rect 2493 4036 2507 4050
rect 2433 3893 2447 3907
rect 2553 4173 2567 4187
rect 2553 4010 2567 4024
rect 2533 3853 2547 3867
rect 2533 3816 2547 3830
rect 2513 3753 2527 3767
rect 2453 3693 2467 3707
rect 2473 3673 2487 3687
rect 2413 3653 2427 3667
rect 2353 3613 2367 3627
rect 2593 4193 2607 4207
rect 2573 3593 2587 3607
rect 2473 3573 2487 3587
rect 2513 3553 2527 3567
rect 2413 3516 2427 3530
rect 2493 3513 2507 3527
rect 2393 3470 2407 3484
rect 2433 3413 2447 3427
rect 2413 3313 2427 3327
rect 2473 3293 2487 3307
rect 2393 3250 2407 3264
rect 2493 3250 2507 3264
rect 2633 5353 2647 5367
rect 2633 5113 2647 5127
rect 2633 4873 2647 4887
rect 2633 4393 2647 4407
rect 2673 5213 2687 5227
rect 2672 4993 2686 5007
rect 2693 4993 2707 5007
rect 2673 4893 2687 4907
rect 2653 4373 2667 4387
rect 2653 4293 2667 4307
rect 2633 4273 2647 4287
rect 2693 4653 2707 4667
rect 2693 4493 2707 4507
rect 2693 4293 2707 4307
rect 2673 4253 2687 4267
rect 2673 4113 2687 4127
rect 2633 4073 2647 4087
rect 2613 4036 2627 4050
rect 2613 3816 2627 3830
rect 2613 3713 2627 3727
rect 2733 5813 2747 5827
rect 2733 5153 2747 5167
rect 2733 5113 2747 5127
rect 2733 4913 2747 4927
rect 2773 5993 2787 6007
rect 2793 5893 2807 5907
rect 2793 5850 2807 5864
rect 2793 5813 2807 5827
rect 2833 6053 2847 6067
rect 2813 5673 2827 5687
rect 2793 5613 2807 5627
rect 2773 5596 2787 5610
rect 2793 5413 2807 5427
rect 2913 6493 2927 6507
rect 2913 6453 2927 6467
rect 2973 6533 2987 6547
rect 3033 6493 3047 6507
rect 2973 6416 2987 6430
rect 3013 6416 3027 6430
rect 2993 6370 3007 6384
rect 3033 6370 3047 6384
rect 3013 6333 3027 6347
rect 2993 6313 3007 6327
rect 2973 6213 2987 6227
rect 2873 6173 2887 6187
rect 2913 6133 2927 6147
rect 2873 5913 2887 5927
rect 2853 5753 2867 5767
rect 2853 5633 2867 5647
rect 3053 6273 3067 6287
rect 3033 6173 3047 6187
rect 2933 5933 2947 5947
rect 2973 5896 2987 5910
rect 3133 7173 3147 7187
rect 3173 7156 3187 7170
rect 3213 7156 3227 7170
rect 3153 7110 3167 7124
rect 3333 7675 3347 7689
rect 3333 7633 3347 7647
rect 3353 7456 3367 7470
rect 3333 7410 3347 7424
rect 3353 7373 3367 7387
rect 3353 7253 3367 7267
rect 3173 7093 3187 7107
rect 3213 7093 3227 7107
rect 3133 7073 3147 7087
rect 3133 6913 3147 6927
rect 3113 6673 3127 6687
rect 3113 6613 3127 6627
rect 3093 6413 3107 6427
rect 3073 6173 3087 6187
rect 3053 5993 3067 6007
rect 2953 5850 2967 5864
rect 2893 5773 2907 5787
rect 2953 5633 2967 5647
rect 2913 5596 2927 5610
rect 2973 5533 2987 5547
rect 2933 5512 2947 5526
rect 2893 5473 2907 5487
rect 2933 5473 2947 5487
rect 2832 5413 2846 5427
rect 2853 5413 2867 5427
rect 2893 5413 2907 5427
rect 2813 5330 2827 5344
rect 2853 5313 2867 5327
rect 2813 5233 2827 5247
rect 2813 5193 2827 5207
rect 2793 5173 2807 5187
rect 2793 5093 2807 5107
rect 2833 5076 2847 5090
rect 2873 5076 2887 5090
rect 2813 5030 2827 5044
rect 2853 5030 2867 5044
rect 2753 4873 2767 4887
rect 2773 4856 2787 4870
rect 2813 4856 2827 4870
rect 2853 4856 2867 4870
rect 2753 4753 2767 4767
rect 2733 4733 2747 4747
rect 2853 4813 2867 4827
rect 2753 4713 2767 4727
rect 2793 4713 2807 4727
rect 2733 4633 2747 4647
rect 2713 4153 2727 4167
rect 2713 4073 2727 4087
rect 2693 3913 2707 3927
rect 2693 3653 2707 3667
rect 2673 3553 2687 3567
rect 2753 4613 2767 4627
rect 2773 4567 2787 4570
rect 2773 4556 2787 4567
rect 2813 4556 2827 4570
rect 2873 4713 2887 4727
rect 2933 5373 2947 5387
rect 2973 5330 2987 5344
rect 2933 5312 2947 5326
rect 2913 5093 2927 5107
rect 2973 5253 2987 5267
rect 2953 5133 2967 5147
rect 2953 5053 2967 5067
rect 2933 5013 2947 5027
rect 2933 4913 2947 4927
rect 2933 4793 2947 4807
rect 2953 4753 2967 4767
rect 2933 4733 2947 4747
rect 2913 4613 2927 4627
rect 2893 4556 2907 4570
rect 2793 4513 2807 4527
rect 2773 4493 2787 4507
rect 2873 4510 2887 4524
rect 2913 4510 2927 4524
rect 2833 4473 2847 4487
rect 2753 4393 2767 4407
rect 2813 4393 2827 4407
rect 2813 4293 2827 4307
rect 2793 4253 2807 4267
rect 2773 3990 2787 4004
rect 2733 3816 2747 3830
rect 2773 3816 2787 3830
rect 2833 4193 2847 4207
rect 2913 4393 2927 4407
rect 2873 4373 2887 4387
rect 2853 4113 2867 4127
rect 2813 4073 2827 4087
rect 2733 3613 2747 3627
rect 2713 3573 2727 3587
rect 2773 3613 2787 3627
rect 2753 3533 2767 3547
rect 2733 3516 2747 3530
rect 2773 3513 2787 3527
rect 2753 3470 2767 3484
rect 2713 3433 2727 3447
rect 2713 3353 2727 3367
rect 2633 3313 2647 3327
rect 2673 3296 2687 3310
rect 2713 3296 2727 3310
rect 2773 3296 2787 3310
rect 2633 3250 2647 3264
rect 2693 3250 2707 3264
rect 2733 3213 2747 3227
rect 2593 3193 2607 3207
rect 2513 3173 2527 3187
rect 2593 3133 2607 3147
rect 2793 3253 2807 3267
rect 2473 3093 2487 3107
rect 2773 3093 2787 3107
rect 2433 3073 2447 3087
rect 2753 3073 2767 3087
rect 2433 3016 2447 3030
rect 2373 2996 2387 3010
rect 2413 2973 2427 2987
rect 2353 2893 2367 2907
rect 2433 2953 2447 2967
rect 2453 2893 2467 2907
rect 2433 2873 2447 2887
rect 2413 2853 2427 2867
rect 2393 2793 2407 2807
rect 2353 2776 2367 2790
rect 2453 2730 2467 2744
rect 2593 2976 2607 2990
rect 2793 3033 2807 3047
rect 2913 4253 2927 4267
rect 2893 4173 2907 4187
rect 2953 4693 2967 4707
rect 2933 4073 2947 4087
rect 2853 4036 2867 4050
rect 2893 4036 2907 4050
rect 2873 3990 2887 4004
rect 3033 5850 3047 5864
rect 3073 5933 3087 5947
rect 3053 5772 3067 5786
rect 3073 5713 3087 5727
rect 3153 6813 3167 6827
rect 3333 7013 3347 7027
rect 3253 6993 3267 7007
rect 3293 6973 3307 6987
rect 3273 6890 3287 6904
rect 3333 6793 3347 6807
rect 3393 8433 3407 8447
rect 3473 8213 3487 8227
rect 3432 8196 3446 8210
rect 3453 8196 3467 8210
rect 3473 8113 3487 8127
rect 3453 8073 3467 8087
rect 3393 7793 3407 7807
rect 3453 7593 3467 7607
rect 3593 8833 3607 8847
rect 3573 8716 3587 8730
rect 3553 8633 3567 8647
rect 3573 8413 3587 8427
rect 3613 8773 3627 8787
rect 3593 8293 3607 8307
rect 3553 8253 3567 8267
rect 3613 8153 3627 8167
rect 3773 9213 3787 9227
rect 3713 8973 3727 8987
rect 3833 9213 3847 9227
rect 3813 9133 3827 9147
rect 3873 9153 3887 9167
rect 3833 9073 3847 9087
rect 3973 9490 3987 9504
rect 4013 9490 4027 9504
rect 4193 9736 4207 9750
rect 4353 9653 4367 9667
rect 4273 9633 4287 9647
rect 4233 9536 4247 9550
rect 4453 9730 4467 9744
rect 4393 9713 4407 9727
rect 4393 9653 4407 9667
rect 4533 9833 4547 9847
rect 4513 9613 4527 9627
rect 4373 9593 4387 9607
rect 4353 9553 4367 9567
rect 4213 9393 4227 9407
rect 4253 9393 4267 9407
rect 3933 9353 3947 9367
rect 4333 9333 4347 9347
rect 4233 9313 4247 9327
rect 3933 9253 3947 9267
rect 3933 9213 3947 9227
rect 4073 9216 4087 9230
rect 4193 9210 4207 9224
rect 4293 9213 4307 9227
rect 3913 9113 3927 9127
rect 4013 9113 4027 9127
rect 3873 9033 3887 9047
rect 3973 9033 3987 9047
rect 3853 9016 3867 9030
rect 3913 8996 3927 9010
rect 3793 8972 3807 8986
rect 3773 8932 3787 8946
rect 3833 8970 3847 8984
rect 3893 8953 3907 8967
rect 3932 8953 3946 8967
rect 3953 8953 3967 8967
rect 3813 8933 3827 8947
rect 3873 8933 3887 8947
rect 3793 8873 3807 8887
rect 3833 8873 3847 8887
rect 3833 8852 3847 8866
rect 3793 8793 3807 8807
rect 3753 8670 3767 8684
rect 3713 8513 3727 8527
rect 3813 8493 3827 8507
rect 3713 8450 3727 8464
rect 3753 8413 3767 8427
rect 3693 8213 3707 8227
rect 3693 8196 3707 8210
rect 3633 8113 3647 8127
rect 3533 8073 3547 8087
rect 3593 8073 3607 8087
rect 3533 7976 3547 7990
rect 3693 8113 3707 8127
rect 3633 8033 3647 8047
rect 3673 8033 3687 8047
rect 3633 7976 3647 7990
rect 3513 7733 3527 7747
rect 3613 7913 3627 7927
rect 3633 7753 3647 7767
rect 3573 7733 3587 7747
rect 3613 7653 3627 7667
rect 3513 7630 3527 7644
rect 3553 7630 3567 7644
rect 3573 7593 3587 7607
rect 3473 7513 3487 7527
rect 3533 7513 3547 7527
rect 3473 7456 3487 7470
rect 3413 7173 3427 7187
rect 3373 6773 3387 6787
rect 3353 6753 3367 6767
rect 3273 6713 3287 6727
rect 3313 6713 3327 6727
rect 3273 6653 3287 6667
rect 3233 6636 3247 6650
rect 3353 6636 3367 6650
rect 3313 6613 3327 6627
rect 3173 6593 3187 6607
rect 3213 6590 3227 6604
rect 3253 6573 3267 6587
rect 3173 6493 3187 6507
rect 3153 6473 3167 6487
rect 3153 6413 3167 6427
rect 3153 6370 3167 6384
rect 3253 6473 3267 6487
rect 3213 6433 3227 6447
rect 3173 6333 3187 6347
rect 3153 6313 3167 6327
rect 3153 6233 3167 6247
rect 3133 6193 3147 6207
rect 3113 6173 3127 6187
rect 3293 6433 3307 6447
rect 3293 6353 3307 6367
rect 3273 6233 3287 6247
rect 3193 6116 3207 6130
rect 3253 6116 3267 6130
rect 3113 6073 3127 6087
rect 3093 5596 3107 5610
rect 3073 5573 3087 5587
rect 3053 5553 3067 5567
rect 3153 6033 3167 6047
rect 3133 5793 3147 5807
rect 3273 6033 3287 6047
rect 3253 5993 3267 6007
rect 3253 5933 3267 5947
rect 3213 5896 3227 5910
rect 3313 6133 3327 6147
rect 3353 6033 3367 6047
rect 3313 5933 3327 5947
rect 3273 5850 3287 5864
rect 3173 5813 3187 5827
rect 3213 5813 3227 5827
rect 3153 5713 3167 5727
rect 3193 5713 3207 5727
rect 3273 5693 3287 5707
rect 3253 5673 3267 5687
rect 3233 5596 3247 5610
rect 3353 5913 3367 5927
rect 3353 5733 3367 5747
rect 3313 5633 3327 5647
rect 3293 5613 3307 5627
rect 3273 5596 3287 5610
rect 3213 5550 3227 5564
rect 3113 5533 3127 5547
rect 3213 5529 3227 5543
rect 3073 5493 3087 5507
rect 3033 5433 3047 5447
rect 3013 5373 3027 5387
rect 3153 5376 3167 5390
rect 3193 5353 3207 5367
rect 3073 5293 3087 5307
rect 3173 5273 3187 5287
rect 3133 5233 3147 5247
rect 3093 5193 3107 5207
rect 3053 5093 3067 5107
rect 3093 5093 3107 5107
rect 3133 5076 3147 5090
rect 3073 5013 3087 5027
rect 3013 4953 3027 4967
rect 3153 4933 3167 4947
rect 3113 4913 3127 4927
rect 2993 4893 3007 4907
rect 2993 4856 3007 4870
rect 3053 4856 3067 4870
rect 2973 4653 2987 4667
rect 2973 4553 2987 4567
rect 2913 3933 2927 3947
rect 2833 3853 2847 3867
rect 2833 3813 2847 3827
rect 2873 3816 2887 3830
rect 3133 4853 3147 4867
rect 3013 4793 3027 4807
rect 3033 4773 3047 4787
rect 3193 5053 3207 5067
rect 3253 5373 3267 5387
rect 3233 5233 3247 5247
rect 3253 5113 3267 5127
rect 3233 4993 3247 5007
rect 3253 4933 3267 4947
rect 3193 4793 3207 4807
rect 3173 4753 3187 4767
rect 3013 4673 3027 4687
rect 3033 4633 3047 4647
rect 3053 4556 3067 4570
rect 3033 4513 3047 4527
rect 3213 4773 3227 4787
rect 3133 4556 3147 4570
rect 3213 4593 3227 4607
rect 3153 4510 3167 4524
rect 3013 4493 3027 4507
rect 3053 4493 3067 4507
rect 3013 4333 3027 4347
rect 3093 4336 3107 4350
rect 3033 4290 3047 4304
rect 3073 4253 3087 4267
rect 3013 4233 3027 4247
rect 3053 4233 3067 4247
rect 3013 4153 3027 4167
rect 3053 4153 3067 4167
rect 2973 3933 2987 3947
rect 2953 3873 2967 3887
rect 3033 4133 3047 4147
rect 3053 4036 3067 4050
rect 3033 4013 3047 4027
rect 3053 3993 3067 4007
rect 3053 3873 3067 3887
rect 3013 3833 3027 3847
rect 2973 3816 2987 3830
rect 3033 3753 3047 3767
rect 2993 3733 3007 3747
rect 2933 3673 2947 3687
rect 2913 3470 2927 3484
rect 2973 3653 2987 3667
rect 2973 3613 2987 3627
rect 3013 3516 3027 3530
rect 2873 3253 2887 3267
rect 2893 3153 2907 3167
rect 2813 3013 2827 3027
rect 2813 2973 2827 2987
rect 2913 3113 2927 3127
rect 2793 2933 2807 2947
rect 2753 2893 2767 2907
rect 2753 2853 2767 2867
rect 2753 2832 2767 2846
rect 2633 2776 2647 2790
rect 2613 2730 2627 2744
rect 2653 2730 2667 2744
rect 2373 2693 2387 2707
rect 2313 2613 2327 2627
rect 1857 2493 1871 2507
rect 2132 2493 2146 2507
rect 2153 2493 2167 2507
rect 2233 2493 2247 2507
rect 2273 2493 2287 2507
rect 2333 2593 2347 2607
rect 2333 2493 2347 2507
rect 2633 2493 2647 2507
rect 2713 2493 2727 2507
rect 2773 2793 2787 2807
rect 2793 2773 2807 2787
rect 2773 2730 2787 2744
rect 1773 2450 1787 2464
rect 1873 2450 1887 2464
rect 1993 2456 2007 2470
rect 2133 2413 2147 2427
rect 1713 2313 1727 2327
rect 2053 2313 2067 2327
rect 2613 2473 2627 2487
rect 2173 2456 2187 2470
rect 1673 2253 1687 2267
rect 2053 2253 2067 2267
rect 1733 2236 1747 2250
rect 1853 2230 1867 2244
rect 2013 2230 2027 2244
rect 2113 2236 2127 2250
rect 2153 2236 2167 2250
rect 1593 2210 1607 2224
rect 1653 2213 1667 2227
rect 1633 2173 1647 2187
rect 1513 2133 1527 2147
rect 1473 1993 1487 2007
rect 2033 2193 2047 2207
rect 1793 2113 1807 2127
rect 2013 2113 2027 2127
rect 1693 1976 1707 1990
rect 1513 1956 1527 1970
rect 1593 1956 1607 1970
rect 1493 1910 1507 1924
rect 1673 1893 1687 1907
rect 1653 1813 1667 1827
rect 1633 1737 1647 1751
rect 1673 1773 1687 1787
rect 1373 1493 1387 1507
rect 1373 1436 1387 1450
rect 1353 1373 1367 1387
rect 1413 1373 1427 1387
rect 1433 1353 1447 1367
rect 1533 1691 1547 1705
rect 1533 1633 1547 1647
rect 1553 1593 1567 1607
rect 1533 1433 1547 1447
rect 1493 1333 1507 1347
rect 1513 1313 1527 1327
rect 1553 1373 1567 1387
rect 1533 1193 1547 1207
rect 2033 2073 2047 2087
rect 2033 2033 2047 2047
rect 1973 1993 1987 2007
rect 1953 1956 1967 1970
rect 1753 1893 1767 1907
rect 1693 1633 1707 1647
rect 1713 1473 1727 1487
rect 1693 1390 1707 1404
rect 1952 1913 1966 1927
rect 2073 1956 2087 1970
rect 2213 2433 2227 2447
rect 2193 2413 2207 2427
rect 1973 1910 1987 1924
rect 2013 1910 2027 1924
rect 2053 1910 2067 1924
rect 2173 1913 2187 1927
rect 1773 1873 1787 1887
rect 2073 1833 2087 1847
rect 1873 1736 1887 1750
rect 2053 1733 2067 1747
rect 1853 1690 1867 1704
rect 1953 1693 1967 1707
rect 1893 1493 1907 1507
rect 1993 1493 2007 1507
rect 1933 1390 1947 1404
rect 1973 1390 1987 1404
rect 1653 1373 1667 1387
rect 1753 1373 1767 1387
rect 2053 1690 2067 1704
rect 2053 1433 2067 1447
rect 2053 1390 2067 1404
rect 2033 1333 2047 1347
rect 1913 1253 1927 1267
rect 2033 1253 2047 1267
rect 1713 1190 1727 1204
rect 2213 2253 2227 2267
rect 2273 2453 2287 2467
rect 2333 2453 2347 2467
rect 2253 2133 2267 2147
rect 2333 2313 2347 2327
rect 2373 2456 2387 2470
rect 2473 2456 2487 2470
rect 2373 2413 2387 2427
rect 2633 2450 2647 2464
rect 2673 2450 2687 2464
rect 2753 2453 2767 2467
rect 2733 2433 2747 2447
rect 2493 2333 2507 2347
rect 2473 2313 2487 2327
rect 2293 2273 2307 2287
rect 2353 2273 2367 2287
rect 2393 2253 2407 2267
rect 2293 2013 2307 2027
rect 2393 2173 2407 2187
rect 2333 1956 2347 1970
rect 2373 1956 2387 1970
rect 2473 1956 2487 1970
rect 2213 1853 2227 1867
rect 2193 1833 2207 1847
rect 2153 1813 2167 1827
rect 2132 1773 2146 1787
rect 2153 1773 2167 1787
rect 2173 1736 2187 1750
rect 2113 1690 2127 1704
rect 2233 1736 2247 1750
rect 2233 1693 2247 1707
rect 2153 1673 2167 1687
rect 2213 1673 2227 1687
rect 2373 1910 2387 1924
rect 2313 1893 2327 1907
rect 2293 1853 2307 1867
rect 2253 1453 2267 1467
rect 1973 1213 1987 1227
rect 2073 1216 2087 1230
rect 1473 1170 1487 1184
rect 1873 1173 1887 1187
rect 1553 1150 1567 1164
rect 1553 1073 1567 1087
rect 1353 993 1367 1007
rect 1453 993 1467 1007
rect 1633 993 1647 1007
rect 1333 916 1347 930
rect 693 853 707 867
rect 653 793 667 807
rect 633 693 647 707
rect 793 873 807 887
rect 753 833 767 847
rect 713 733 727 747
rect 633 650 647 664
rect 673 650 687 664
rect 513 593 527 607
rect 133 493 147 507
rect 353 493 367 507
rect 453 493 467 507
rect 513 493 527 507
rect 93 370 107 384
rect 133 370 147 384
rect 293 376 307 390
rect 392 376 406 390
rect 693 453 707 467
rect 413 370 427 384
rect 493 373 507 387
rect 973 870 987 884
rect 1053 870 1067 884
rect 1053 793 1067 807
rect 1293 793 1307 807
rect 1353 793 1367 807
rect 1013 753 1027 767
rect 993 733 1007 747
rect 1073 753 1087 767
rect 1013 633 1027 647
rect 1053 633 1067 647
rect 1293 713 1307 727
rect 1293 613 1307 627
rect 1073 493 1087 507
rect 1233 493 1247 507
rect 893 433 907 447
rect 953 433 967 447
rect 953 396 967 410
rect 893 350 907 364
rect 933 350 947 364
rect 973 350 987 364
rect 393 333 407 347
rect 753 333 767 347
rect 33 273 47 287
rect 193 273 207 287
rect 533 233 547 247
rect 713 233 727 247
rect 753 233 767 247
rect 473 176 487 190
rect 213 130 227 144
rect 673 173 687 187
rect 713 176 727 190
rect 813 176 827 190
rect 493 113 507 127
rect 533 113 547 127
rect 733 130 747 144
rect 1033 176 1047 190
rect 1173 453 1187 467
rect 1353 433 1367 447
rect 1213 413 1227 427
rect 1273 413 1287 427
rect 1193 350 1207 364
rect 1173 233 1187 247
rect 1113 193 1127 207
rect 913 130 927 144
rect 1053 130 1067 144
rect 673 93 687 107
rect 773 93 787 107
rect 813 93 827 107
rect 1013 93 1027 107
rect 1113 93 1127 107
rect 1213 173 1227 187
rect 1593 916 1607 930
rect 2233 1436 2247 1450
rect 2393 1690 2407 1704
rect 2373 1453 2387 1467
rect 2313 1433 2327 1447
rect 2213 1390 2227 1404
rect 2253 1390 2267 1404
rect 2293 1390 2307 1404
rect 2273 1333 2287 1347
rect 2193 1216 2207 1230
rect 2153 1133 2167 1147
rect 1993 993 2007 1007
rect 2113 993 2127 1007
rect 2193 993 2207 1007
rect 1833 973 1847 987
rect 1873 973 1887 987
rect 1613 870 1627 884
rect 1933 933 1947 947
rect 1893 916 1907 930
rect 2093 916 2107 930
rect 1873 870 1887 884
rect 1953 870 1967 884
rect 1993 870 2007 884
rect 2093 873 2107 887
rect 1833 833 1847 847
rect 1913 833 1927 847
rect 1573 793 1587 807
rect 1533 733 1547 747
rect 1853 733 1867 747
rect 1493 713 1507 727
rect 1573 693 1587 707
rect 1753 696 1767 710
rect 1793 696 1807 710
rect 1513 650 1527 664
rect 1513 433 1527 447
rect 1352 393 1366 407
rect 1373 393 1387 407
rect 1453 393 1467 407
rect 1273 313 1287 327
rect 1253 253 1267 267
rect 1333 213 1347 227
rect 1773 650 1787 664
rect 1773 553 1787 567
rect 1793 533 1807 547
rect 1753 453 1767 467
rect 1813 493 1827 507
rect 1533 350 1547 364
rect 1573 350 1587 364
rect 1493 293 1507 307
rect 1773 313 1787 327
rect 1753 293 1767 307
rect 1793 293 1807 307
rect 1733 253 1747 267
rect 1373 193 1387 207
rect 1253 152 1267 166
rect 1453 156 1467 170
rect 1573 150 1587 164
rect 2073 853 2087 867
rect 2033 793 2047 807
rect 2073 793 2087 807
rect 2153 953 2167 967
rect 2213 933 2227 947
rect 2213 870 2227 884
rect 2173 813 2187 827
rect 2153 773 2167 787
rect 2073 713 2087 727
rect 2113 713 2127 727
rect 2093 650 2107 664
rect 2053 613 2067 627
rect 2033 493 2047 507
rect 2173 650 2187 664
rect 2073 453 2087 467
rect 2153 453 2167 467
rect 2193 413 2207 427
rect 2053 350 2067 364
rect 2093 350 2107 364
rect 2113 273 2127 287
rect 2113 233 2127 247
rect 2013 213 2027 227
rect 2093 213 2107 227
rect 1993 176 2007 190
rect 1273 113 1287 127
rect 1353 130 1367 144
rect 1413 110 1427 124
rect 2053 176 2067 190
rect 2093 176 2107 190
rect 2193 153 2207 167
rect 2233 393 2247 407
rect 2333 915 2347 929
rect 2653 2393 2667 2407
rect 2753 2333 2767 2347
rect 2513 2293 2527 2307
rect 2632 2293 2646 2307
rect 2653 2293 2667 2307
rect 2713 2273 2727 2287
rect 2593 2256 2607 2270
rect 2613 2210 2627 2224
rect 2613 2153 2627 2167
rect 2513 2013 2527 2027
rect 2573 1956 2587 1970
rect 2553 1910 2567 1924
rect 2593 1910 2607 1924
rect 2673 1813 2687 1827
rect 2513 1613 2527 1627
rect 2493 1593 2507 1607
rect 2473 1513 2487 1527
rect 2393 1413 2407 1427
rect 2453 1390 2467 1404
rect 2513 1390 2527 1404
rect 2393 1353 2407 1367
rect 2453 1170 2467 1184
rect 2393 1073 2407 1087
rect 2373 733 2387 747
rect 2353 650 2367 664
rect 2353 613 2367 627
rect 2313 553 2327 567
rect 2333 453 2347 467
rect 2613 1733 2627 1747
rect 2793 2210 2807 2224
rect 2773 2113 2787 2127
rect 2733 1953 2747 1967
rect 2793 1955 2807 1969
rect 2853 2913 2867 2927
rect 2913 2913 2927 2927
rect 2853 2833 2867 2847
rect 2913 2833 2927 2847
rect 2873 2793 2887 2807
rect 2833 2773 2847 2787
rect 3033 3470 3047 3484
rect 3033 3053 3047 3067
rect 2993 2996 3007 3010
rect 3093 4113 3107 4127
rect 3233 4513 3247 4527
rect 3193 4336 3207 4350
rect 3193 4193 3207 4207
rect 3173 4113 3187 4127
rect 3113 4073 3127 4087
rect 3153 4036 3167 4050
rect 3193 4036 3207 4050
rect 3173 3990 3187 4004
rect 3313 5550 3327 5564
rect 3353 5493 3367 5507
rect 3313 5413 3327 5427
rect 3433 7110 3447 7124
rect 3553 7453 3567 7467
rect 3413 6573 3427 6587
rect 3393 6353 3407 6367
rect 3393 6193 3407 6207
rect 3473 6853 3487 6867
rect 3533 7110 3547 7124
rect 3613 7533 3627 7547
rect 3573 7093 3587 7107
rect 3553 7013 3567 7027
rect 3673 7513 3687 7527
rect 3713 7913 3727 7927
rect 3793 8149 3807 8163
rect 3753 7833 3767 7847
rect 3753 7812 3767 7826
rect 3713 7573 3727 7587
rect 3693 7453 3707 7467
rect 3793 7713 3807 7727
rect 3933 8753 3947 8767
rect 4033 9033 4047 9047
rect 4033 8993 4047 9007
rect 4173 8990 4187 9004
rect 4313 9190 4327 9204
rect 4333 9153 4347 9167
rect 4393 9513 4407 9527
rect 4373 9453 4387 9467
rect 4413 9413 4427 9427
rect 4473 9353 4487 9367
rect 4413 9313 4427 9327
rect 4653 10593 4667 10607
rect 4593 9973 4607 9987
rect 4633 9973 4647 9987
rect 4573 9513 4587 9527
rect 4553 9473 4567 9487
rect 4493 9333 4507 9347
rect 4533 9333 4547 9347
rect 4473 9293 4487 9307
rect 4393 9253 4407 9267
rect 4373 9193 4387 9207
rect 4493 9273 4507 9287
rect 4513 9236 4527 9250
rect 4573 9236 4587 9250
rect 4793 10770 4807 10784
rect 4833 10770 4847 10784
rect 4833 10673 4847 10687
rect 4813 10633 4827 10647
rect 4753 10613 4767 10627
rect 4773 10576 4787 10590
rect 4873 10793 4887 10807
rect 4793 10530 4807 10544
rect 4853 10530 4867 10544
rect 4693 10493 4707 10507
rect 4673 10213 4687 10227
rect 4673 10113 4687 10127
rect 4713 10413 4727 10427
rect 4753 10373 4767 10387
rect 4873 10373 4887 10387
rect 4813 10353 4827 10367
rect 4873 10313 4887 10327
rect 4793 10276 4807 10290
rect 4713 10233 4727 10247
rect 4693 10013 4707 10027
rect 4713 9993 4727 10007
rect 4773 10173 4787 10187
rect 4873 10153 4887 10167
rect 4773 10053 4787 10067
rect 4833 10056 4847 10070
rect 4753 10013 4767 10027
rect 4733 9933 4747 9947
rect 4673 9833 4687 9847
rect 4713 9793 4727 9807
rect 4633 9753 4647 9767
rect 4673 9756 4687 9770
rect 5033 11173 5047 11187
rect 5053 11050 5067 11064
rect 5013 11013 5027 11027
rect 5053 10993 5067 11007
rect 5093 11193 5107 11207
rect 5073 10953 5087 10967
rect 4933 10873 4947 10887
rect 5033 10873 5047 10887
rect 4913 10493 4927 10507
rect 4953 10813 4967 10827
rect 5113 11053 5127 11067
rect 5153 10933 5167 10947
rect 5093 10813 5107 10827
rect 5073 10750 5087 10764
rect 5133 10713 5147 10727
rect 4973 10633 4987 10647
rect 4953 10593 4967 10607
rect 5033 10593 5047 10607
rect 5073 10576 5087 10590
rect 5033 10513 5047 10527
rect 4933 10353 4947 10367
rect 4933 10276 4947 10290
rect 4933 10213 4947 10227
rect 4893 10033 4907 10047
rect 5093 10493 5107 10507
rect 5153 10593 5167 10607
rect 5153 10572 5167 10586
rect 5053 10473 5067 10487
rect 5133 10473 5147 10487
rect 5073 10276 5087 10290
rect 4973 10230 4987 10244
rect 5013 10230 5027 10244
rect 5053 10230 5067 10244
rect 5193 11393 5207 11407
rect 5313 11373 5327 11387
rect 5353 11353 5367 11367
rect 5433 11453 5447 11467
rect 5413 11433 5427 11447
rect 5233 11253 5247 11267
rect 5233 11096 5247 11110
rect 5193 11013 5207 11027
rect 5273 11050 5287 11064
rect 5253 10953 5267 10967
rect 5213 10793 5227 10807
rect 5353 11133 5367 11147
rect 5393 11050 5407 11064
rect 5393 10993 5407 11007
rect 5373 10973 5387 10987
rect 5353 10953 5367 10967
rect 5332 10913 5346 10927
rect 5353 10913 5367 10927
rect 5293 10833 5307 10847
rect 5333 10796 5347 10810
rect 5253 10750 5267 10764
rect 5313 10750 5327 10764
rect 5193 10693 5207 10707
rect 5173 10493 5187 10507
rect 5233 10533 5247 10547
rect 5213 10413 5227 10427
rect 5193 10373 5207 10387
rect 5233 10293 5247 10307
rect 5213 10153 5227 10167
rect 5153 10133 5167 10147
rect 5073 10030 5087 10044
rect 4813 10010 4827 10024
rect 4773 9893 4787 9907
rect 4753 9773 4767 9787
rect 4893 9993 4907 10007
rect 4853 9953 4867 9967
rect 4873 9756 4887 9770
rect 4693 9710 4707 9724
rect 4733 9710 4747 9724
rect 4813 9713 4827 9727
rect 4853 9713 4867 9727
rect 4833 9693 4847 9707
rect 4633 9673 4647 9687
rect 4633 9473 4647 9487
rect 4693 9433 4707 9447
rect 4633 9353 4647 9367
rect 4793 9633 4807 9647
rect 4793 9593 4807 9607
rect 4813 9513 4827 9527
rect 4793 9493 4807 9507
rect 4773 9413 4787 9427
rect 4793 9393 4807 9407
rect 4693 9273 4707 9287
rect 4353 9033 4367 9047
rect 4313 8993 4327 9007
rect 4453 9190 4467 9204
rect 4573 9193 4587 9207
rect 4493 9173 4507 9187
rect 4553 9153 4567 9167
rect 4713 9236 4727 9250
rect 4753 9236 4767 9250
rect 4793 9236 4807 9250
rect 4873 9673 4887 9687
rect 4853 9653 4867 9667
rect 5333 10673 5347 10687
rect 5273 10633 5287 10647
rect 5353 10653 5367 10667
rect 5473 11570 5487 11584
rect 5453 11353 5467 11367
rect 5453 11316 5467 11330
rect 5433 11193 5447 11207
rect 5473 11213 5487 11227
rect 5693 11773 5707 11787
rect 5673 11753 5687 11767
rect 5653 11653 5667 11667
rect 5573 11616 5587 11630
rect 5613 11616 5627 11630
rect 5593 11570 5607 11584
rect 5633 11570 5647 11584
rect 5513 11493 5527 11507
rect 5893 11816 5907 11830
rect 5873 11773 5887 11787
rect 5813 11713 5827 11727
rect 5753 11693 5767 11707
rect 5833 11613 5847 11627
rect 5933 11853 5947 11867
rect 6273 11833 6287 11847
rect 6073 11816 6087 11830
rect 5933 11793 5947 11807
rect 5933 11616 5947 11630
rect 6013 11616 6027 11630
rect 5813 11570 5827 11584
rect 5853 11473 5867 11487
rect 5673 11453 5687 11467
rect 5853 11433 5867 11447
rect 5653 11413 5667 11427
rect 5573 11316 5587 11330
rect 5613 11316 5627 11330
rect 5833 11353 5847 11367
rect 5693 11316 5707 11330
rect 5873 11316 5887 11330
rect 5933 11316 5947 11330
rect 5593 11270 5607 11284
rect 5653 11273 5667 11287
rect 5693 11273 5707 11287
rect 5853 11270 5867 11284
rect 5913 11273 5927 11287
rect 5513 11253 5527 11267
rect 5553 11253 5567 11267
rect 5853 11213 5867 11227
rect 5453 11173 5467 11187
rect 5493 11173 5507 11187
rect 5573 11173 5587 11187
rect 5433 11096 5447 11110
rect 5433 10873 5447 10887
rect 5433 10833 5447 10847
rect 5413 10633 5427 10647
rect 5333 10613 5347 10627
rect 5413 10612 5427 10626
rect 5273 10576 5287 10590
rect 5313 10576 5327 10590
rect 5353 10576 5367 10590
rect 5333 10530 5347 10544
rect 5373 10530 5387 10544
rect 5413 10530 5427 10544
rect 5413 10493 5427 10507
rect 5273 10473 5287 10487
rect 5333 10473 5347 10487
rect 5373 10373 5387 10387
rect 5253 10233 5267 10247
rect 5293 10230 5307 10244
rect 5273 10153 5287 10167
rect 5253 10093 5267 10107
rect 5253 10030 5267 10044
rect 5333 10173 5347 10187
rect 5333 10133 5347 10147
rect 5293 10033 5307 10047
rect 4993 9893 5007 9907
rect 5233 9893 5247 9907
rect 5213 9853 5227 9867
rect 5193 9793 5207 9807
rect 5033 9756 5047 9770
rect 5073 9753 5087 9767
rect 4913 9613 4927 9627
rect 4893 9553 4907 9567
rect 5013 9710 5027 9724
rect 5253 9833 5267 9847
rect 5333 9833 5347 9847
rect 5293 9793 5307 9807
rect 5333 9773 5347 9787
rect 5213 9710 5227 9724
rect 5273 9710 5287 9724
rect 5313 9710 5327 9724
rect 5193 9633 5207 9647
rect 5273 9633 5287 9647
rect 5073 9613 5087 9627
rect 4973 9593 4987 9607
rect 5293 9613 5307 9627
rect 5293 9573 5307 9587
rect 5313 9553 5327 9567
rect 5353 9553 5367 9567
rect 4993 9516 5007 9530
rect 5113 9510 5127 9524
rect 4873 9490 4887 9504
rect 5273 9516 5287 9530
rect 5313 9516 5327 9530
rect 5393 10353 5407 10367
rect 5393 9573 5407 9587
rect 5373 9533 5387 9547
rect 5253 9473 5267 9487
rect 5293 9473 5307 9487
rect 5353 9473 5367 9487
rect 5273 9433 5287 9447
rect 4953 9413 4967 9427
rect 5153 9393 5167 9407
rect 4873 9353 4887 9367
rect 4713 9133 4727 9147
rect 4553 9093 4567 9107
rect 4693 9093 4707 9107
rect 4553 8990 4567 9004
rect 4313 8953 4327 8967
rect 4173 8893 4187 8907
rect 4013 8853 4027 8867
rect 4033 8753 4047 8767
rect 3993 8716 4007 8730
rect 4013 8670 4027 8684
rect 3953 8633 3967 8647
rect 3893 8613 3907 8627
rect 3913 8593 3927 8607
rect 4013 8533 4027 8547
rect 3953 8513 3967 8527
rect 3973 8513 3987 8527
rect 4153 8813 4167 8827
rect 4173 8773 4187 8787
rect 4153 8716 4167 8730
rect 4333 8873 4347 8887
rect 4313 8813 4327 8827
rect 4253 8716 4267 8730
rect 4293 8716 4307 8730
rect 4333 8716 4347 8730
rect 4233 8653 4247 8667
rect 4333 8673 4347 8687
rect 4193 8633 4207 8647
rect 4273 8633 4287 8647
rect 4173 8613 4187 8627
rect 4153 8593 4167 8607
rect 4213 8470 4227 8484
rect 3913 8453 3927 8467
rect 3913 8293 3927 8307
rect 3893 8033 3907 8047
rect 4773 9190 4787 9204
rect 4813 9190 4827 9204
rect 4773 9153 4787 9167
rect 4773 9113 4787 9127
rect 4753 9093 4767 9107
rect 4733 8993 4747 9007
rect 4813 9013 4827 9027
rect 4733 8953 4747 8967
rect 4853 8953 4867 8967
rect 4413 8893 4427 8907
rect 4713 8893 4727 8907
rect 4613 8833 4627 8847
rect 4593 8813 4607 8827
rect 4513 8753 4527 8767
rect 4553 8716 4567 8730
rect 4533 8670 4547 8684
rect 4533 8613 4547 8627
rect 4473 8593 4487 8607
rect 4412 8573 4426 8587
rect 4433 8573 4447 8587
rect 4413 8493 4427 8507
rect 4433 8470 4447 8484
rect 4473 8413 4487 8427
rect 4053 8393 4067 8407
rect 4373 8393 4387 8407
rect 4353 8333 4367 8347
rect 4153 8273 4167 8287
rect 3993 8253 4007 8267
rect 4033 8253 4047 8267
rect 4073 8253 4087 8267
rect 3933 8195 3947 8209
rect 4033 8193 4047 8207
rect 4033 8149 4047 8163
rect 3953 8073 3967 8087
rect 3913 7976 3927 7990
rect 4033 8033 4047 8047
rect 3993 7993 4007 8007
rect 3973 7976 3987 7990
rect 3893 7930 3907 7944
rect 3953 7930 3967 7944
rect 3853 7893 3867 7907
rect 3913 7833 3927 7847
rect 3853 7733 3867 7747
rect 3813 7676 3827 7690
rect 3893 7676 3907 7690
rect 3833 7553 3847 7567
rect 3793 7513 3807 7527
rect 3853 7456 3867 7470
rect 3773 7410 3787 7424
rect 3633 7193 3647 7207
rect 3673 7193 3687 7207
rect 3693 7156 3707 7170
rect 3633 7093 3647 7107
rect 3673 7093 3687 7107
rect 3613 6993 3627 7007
rect 3593 6973 3607 6987
rect 3553 6936 3567 6950
rect 3693 7073 3707 7087
rect 3653 6973 3667 6987
rect 3633 6937 3647 6951
rect 3513 6893 3527 6907
rect 3493 6793 3507 6807
rect 3473 6753 3487 6767
rect 3573 6890 3587 6904
rect 3533 6853 3547 6867
rect 3572 6793 3586 6807
rect 3593 6793 3607 6807
rect 3533 6773 3547 6787
rect 3453 6653 3467 6667
rect 3513 6653 3527 6667
rect 3493 6636 3507 6650
rect 3593 6713 3607 6727
rect 3613 6693 3627 6707
rect 3593 6613 3607 6627
rect 3513 6553 3527 6567
rect 3573 6553 3587 6567
rect 3453 6353 3467 6367
rect 3433 6273 3447 6287
rect 3653 6890 3667 6904
rect 3653 6833 3667 6847
rect 3653 6713 3667 6727
rect 3633 6573 3647 6587
rect 3613 6553 3627 6567
rect 3593 6493 3607 6507
rect 3573 6416 3587 6430
rect 3593 6370 3607 6384
rect 3553 6333 3567 6347
rect 3633 6313 3647 6327
rect 3513 6233 3527 6247
rect 3593 6233 3607 6247
rect 3413 6133 3427 6147
rect 3473 6053 3487 6067
rect 3533 6053 3547 6067
rect 3433 6013 3447 6027
rect 3493 6013 3507 6027
rect 3493 5973 3507 5987
rect 3553 6013 3567 6027
rect 3393 5733 3407 5747
rect 3373 5453 3387 5467
rect 3513 5850 3527 5864
rect 3413 5673 3427 5687
rect 3553 5793 3567 5807
rect 3553 5753 3567 5767
rect 3473 5633 3487 5647
rect 3533 5633 3547 5647
rect 3513 5593 3527 5607
rect 3433 5553 3447 5567
rect 3413 5473 3427 5487
rect 3313 5333 3327 5347
rect 3373 5330 3387 5344
rect 3393 5213 3407 5227
rect 3393 5173 3407 5187
rect 3413 5153 3427 5167
rect 3493 5550 3507 5564
rect 3453 5513 3467 5527
rect 3473 5473 3487 5487
rect 3453 5433 3467 5447
rect 3473 5153 3487 5167
rect 3433 5113 3447 5127
rect 3292 5076 3306 5090
rect 3313 5076 3327 5090
rect 3373 5076 3387 5090
rect 3453 5092 3467 5106
rect 3393 5030 3407 5044
rect 3313 4893 3327 4907
rect 3333 4856 3347 4870
rect 3453 4953 3467 4967
rect 3413 4833 3427 4847
rect 3273 4513 3287 4527
rect 3313 4810 3327 4824
rect 3313 4753 3327 4767
rect 3293 4453 3307 4467
rect 3273 4332 3287 4346
rect 3273 4032 3287 4046
rect 3133 3953 3147 3967
rect 3093 3893 3107 3907
rect 3093 3713 3107 3727
rect 3093 3516 3107 3530
rect 3093 3353 3107 3367
rect 3133 3913 3147 3927
rect 3253 3973 3267 3987
rect 3273 3933 3287 3947
rect 3273 3893 3287 3907
rect 3253 3833 3267 3847
rect 3513 5193 3527 5207
rect 3473 4810 3487 4824
rect 3413 4773 3427 4787
rect 3453 4773 3467 4787
rect 3453 4733 3467 4747
rect 3353 4713 3367 4727
rect 3413 4713 3427 4727
rect 3373 4556 3387 4570
rect 3453 4556 3467 4570
rect 3333 4393 3347 4407
rect 3313 4333 3327 4347
rect 3493 4553 3507 4567
rect 3433 4510 3447 4524
rect 3413 4373 3427 4387
rect 3393 4290 3407 4304
rect 3373 4213 3387 4227
rect 3353 4173 3367 4187
rect 3313 4073 3327 4087
rect 3293 3833 3307 3847
rect 3313 3813 3327 3827
rect 3213 3673 3227 3687
rect 3293 3770 3307 3784
rect 3273 3753 3287 3767
rect 3153 3613 3167 3627
rect 3253 3613 3267 3627
rect 3313 3613 3327 3627
rect 3153 3553 3167 3567
rect 3153 3513 3167 3527
rect 3233 3516 3247 3530
rect 3253 3470 3267 3484
rect 3313 3473 3327 3487
rect 3233 3296 3247 3310
rect 3273 3293 3287 3307
rect 3193 3250 3207 3264
rect 3153 3193 3167 3207
rect 3133 3153 3147 3167
rect 3113 3113 3127 3127
rect 3113 2996 3127 3010
rect 3193 3093 3207 3107
rect 3033 2933 3047 2947
rect 3013 2873 3027 2887
rect 2973 2853 2987 2867
rect 2973 2793 2987 2807
rect 2953 2753 2967 2767
rect 3013 2753 3027 2767
rect 3193 2993 3207 3007
rect 3133 2933 3147 2947
rect 3193 2933 3207 2947
rect 3353 3813 3367 3827
rect 3353 3770 3367 3784
rect 3353 3573 3367 3587
rect 3453 4173 3467 4187
rect 3393 4113 3407 4127
rect 3393 4033 3407 4047
rect 3493 4513 3507 4527
rect 3613 6053 3627 6067
rect 3613 5893 3627 5907
rect 3613 5850 3627 5864
rect 3773 7353 3787 7367
rect 3753 7193 3767 7207
rect 3733 7073 3747 7087
rect 3713 6893 3727 6907
rect 3753 6891 3767 6905
rect 3713 6853 3727 6867
rect 3733 6833 3747 6847
rect 3733 6793 3747 6807
rect 3693 6673 3707 6687
rect 3833 7313 3847 7327
rect 3793 7293 3807 7307
rect 3673 6653 3687 6667
rect 3773 6653 3787 6667
rect 3693 6613 3707 6627
rect 3673 6590 3687 6604
rect 3673 6493 3687 6507
rect 3813 7213 3827 7227
rect 3813 7156 3827 7170
rect 3813 7113 3827 7127
rect 3873 7213 3887 7227
rect 3933 7773 3947 7787
rect 3913 7353 3927 7367
rect 3933 7333 3947 7347
rect 4173 8233 4187 8247
rect 4173 8153 4187 8167
rect 4153 8113 4167 8127
rect 4153 7993 4167 8007
rect 4253 8195 4267 8209
rect 4213 8073 4227 8087
rect 4193 7973 4207 7987
rect 4173 7930 4187 7944
rect 4173 7893 4187 7907
rect 4113 7873 4127 7887
rect 4113 7813 4127 7827
rect 4073 7753 4087 7767
rect 4113 7733 4127 7747
rect 4073 7676 4087 7690
rect 4093 7573 4107 7587
rect 4033 7456 4047 7470
rect 4193 7456 4207 7470
rect 4013 7410 4027 7424
rect 4173 7413 4187 7427
rect 3973 7293 3987 7307
rect 3933 7233 3947 7247
rect 3933 7192 3947 7206
rect 3973 7156 3987 7170
rect 3953 7110 3967 7124
rect 3873 7093 3887 7107
rect 3853 7053 3867 7067
rect 3873 7033 3887 7047
rect 3893 7013 3907 7027
rect 3993 6993 4007 7007
rect 3913 6937 3927 6951
rect 3953 6933 3967 6947
rect 3933 6913 3947 6927
rect 3813 6891 3827 6905
rect 3913 6873 3927 6887
rect 3913 6753 3927 6767
rect 3813 6673 3827 6687
rect 3733 6590 3747 6604
rect 3893 6653 3907 6667
rect 3853 6453 3867 6467
rect 3813 6416 3827 6430
rect 3693 6370 3707 6384
rect 3793 6370 3807 6384
rect 3793 6353 3807 6367
rect 3673 6333 3687 6347
rect 3713 6333 3727 6347
rect 3793 6253 3807 6267
rect 3713 6193 3727 6207
rect 3673 6173 3687 6187
rect 3753 6173 3767 6187
rect 3713 6116 3727 6130
rect 3693 6073 3707 6087
rect 3773 6070 3787 6084
rect 3993 6873 4007 6887
rect 4273 8150 4287 8164
rect 4273 8113 4287 8127
rect 4233 8033 4247 8047
rect 4233 7893 4247 7907
rect 4313 8093 4327 8107
rect 4333 7933 4347 7947
rect 4373 8195 4387 8209
rect 4473 8153 4487 8167
rect 4533 8333 4547 8347
rect 4653 8753 4667 8767
rect 4693 8713 4707 8727
rect 4693 8653 4707 8667
rect 4633 8533 4647 8547
rect 4573 8413 4587 8427
rect 4653 8493 4667 8507
rect 4793 8716 4807 8730
rect 5133 9373 5147 9387
rect 5113 9353 5127 9367
rect 4913 9333 4927 9347
rect 5133 9333 5147 9347
rect 4893 9190 4907 9204
rect 5033 9236 5047 9250
rect 5113 9236 5127 9250
rect 4993 9193 5007 9207
rect 5053 9190 5067 9204
rect 4933 9153 4947 9167
rect 4913 8813 4927 8827
rect 4873 8753 4887 8767
rect 4913 8733 4927 8747
rect 4853 8716 4867 8730
rect 4913 8693 4927 8707
rect 5113 9133 5127 9147
rect 5073 9033 5087 9047
rect 5113 9033 5127 9047
rect 5133 9013 5147 9027
rect 5013 8993 5027 9007
rect 5093 8970 5107 8984
rect 5133 8973 5147 8987
rect 5053 8933 5067 8947
rect 5053 8793 5067 8807
rect 5013 8773 5027 8787
rect 4733 8613 4747 8627
rect 4733 8573 4747 8587
rect 4793 8493 4807 8507
rect 4653 8433 4667 8447
rect 4633 8373 4647 8387
rect 4573 8293 4587 8307
rect 4553 8273 4567 8287
rect 4573 8253 4587 8267
rect 4553 8196 4567 8210
rect 4593 8196 4607 8210
rect 4533 8150 4547 8164
rect 4653 8196 4667 8210
rect 4493 8113 4507 8127
rect 4433 8093 4447 8107
rect 4393 7993 4407 8007
rect 4593 8133 4607 8147
rect 4573 8093 4587 8107
rect 4533 8073 4547 8087
rect 4573 8053 4587 8067
rect 4493 8033 4507 8047
rect 4493 7993 4507 8007
rect 4513 7956 4527 7970
rect 4593 7953 4607 7967
rect 4353 7913 4367 7927
rect 4453 7930 4467 7944
rect 4433 7913 4447 7927
rect 4413 7873 4427 7887
rect 4353 7676 4367 7690
rect 4413 7673 4427 7687
rect 4413 7630 4427 7644
rect 4373 7553 4387 7567
rect 4313 7456 4327 7470
rect 4192 7373 4206 7387
rect 4213 7373 4227 7387
rect 4293 7393 4307 7407
rect 4273 7373 4287 7387
rect 4073 7293 4087 7307
rect 4113 7293 4127 7307
rect 4253 7293 4267 7307
rect 4053 7193 4067 7207
rect 4053 7110 4067 7124
rect 4133 7156 4147 7170
rect 4193 7156 4207 7170
rect 4233 7156 4247 7170
rect 4173 7110 4187 7124
rect 4173 7073 4187 7087
rect 4133 7033 4147 7047
rect 4113 6973 4127 6987
rect 4253 7113 4267 7127
rect 4253 7073 4267 7087
rect 4213 7033 4227 7047
rect 4193 6973 4207 6987
rect 4233 6953 4247 6967
rect 4213 6933 4227 6947
rect 4233 6916 4247 6930
rect 4333 7293 4347 7307
rect 4293 7173 4307 7187
rect 4293 6993 4307 7007
rect 4273 6913 4287 6927
rect 4073 6873 4087 6887
rect 4013 6853 4027 6867
rect 4053 6833 4067 6847
rect 3953 6773 3967 6787
rect 4053 6773 4067 6787
rect 3973 6673 3987 6687
rect 4013 6636 4027 6650
rect 3933 6613 3947 6627
rect 4133 6853 4147 6867
rect 3893 6273 3907 6287
rect 3833 6193 3847 6207
rect 3733 6033 3747 6047
rect 3813 6033 3827 6047
rect 3793 6013 3807 6027
rect 3693 5973 3707 5987
rect 3733 5973 3747 5987
rect 3673 5850 3687 5864
rect 3653 5773 3667 5787
rect 3633 5593 3647 5607
rect 3793 5896 3807 5910
rect 3953 6590 3967 6604
rect 3993 6590 4007 6604
rect 3933 6233 3947 6247
rect 3853 6070 3867 6084
rect 3913 6116 3927 6130
rect 3893 6052 3907 6066
rect 3873 5993 3887 6007
rect 3893 5896 3907 5910
rect 3773 5850 3787 5864
rect 3813 5813 3827 5827
rect 3793 5753 3807 5767
rect 3773 5653 3787 5667
rect 3713 5550 3727 5564
rect 3633 5513 3647 5527
rect 3573 5472 3587 5486
rect 3533 5153 3547 5167
rect 3533 4913 3547 4927
rect 3533 4733 3547 4747
rect 3533 4553 3547 4567
rect 3513 4253 3527 4267
rect 3493 4213 3507 4227
rect 3513 4133 3527 4147
rect 3493 4113 3507 4127
rect 3473 4073 3487 4087
rect 3573 5413 3587 5427
rect 3573 5376 3587 5390
rect 3673 5376 3687 5390
rect 3733 5353 3747 5367
rect 3653 5330 3667 5344
rect 3713 5330 3727 5344
rect 3613 5273 3627 5287
rect 3633 5253 3647 5267
rect 3593 5153 3607 5167
rect 3593 5073 3607 5087
rect 3713 5273 3727 5287
rect 3653 5233 3667 5247
rect 3733 5233 3747 5247
rect 3693 5193 3707 5207
rect 3673 5093 3687 5107
rect 3873 5673 3887 5687
rect 3933 6070 3947 6084
rect 3933 5993 3947 6007
rect 3913 5753 3927 5767
rect 3893 5653 3907 5667
rect 3873 5633 3887 5647
rect 4033 6553 4047 6567
rect 4113 6593 4127 6607
rect 4173 6873 4187 6887
rect 4213 6873 4227 6887
rect 4093 6513 4107 6527
rect 4073 6473 4087 6487
rect 4053 6413 4067 6427
rect 4133 6416 4147 6430
rect 4193 6553 4207 6567
rect 4193 6513 4207 6527
rect 4173 6413 4187 6427
rect 4053 6273 4067 6287
rect 3973 6193 3987 6207
rect 4033 6173 4047 6187
rect 4033 6133 4047 6147
rect 3993 6116 4007 6130
rect 3973 6053 3987 6067
rect 4053 6070 4067 6084
rect 4013 6053 4027 6067
rect 4153 6370 4167 6384
rect 4133 6133 4147 6147
rect 4053 6033 4067 6047
rect 4113 6033 4127 6047
rect 4013 5896 4027 5910
rect 4113 5973 4127 5987
rect 4093 5953 4107 5967
rect 4033 5850 4047 5864
rect 3993 5773 4007 5787
rect 3953 5753 3967 5767
rect 3973 5596 3987 5610
rect 4013 5593 4027 5607
rect 3833 5550 3847 5564
rect 3993 5550 4007 5564
rect 3812 5473 3826 5487
rect 3833 5473 3847 5487
rect 3833 5452 3847 5466
rect 3813 5433 3827 5447
rect 3813 5376 3827 5390
rect 3793 5313 3807 5327
rect 3853 5413 3867 5427
rect 3893 5376 3907 5390
rect 3933 5376 3947 5390
rect 3833 5313 3847 5327
rect 3773 5273 3787 5287
rect 3753 5093 3767 5107
rect 3693 5073 3707 5087
rect 3653 5030 3667 5044
rect 3613 5013 3627 5027
rect 3653 5009 3667 5023
rect 3693 5013 3707 5027
rect 3573 4933 3587 4947
rect 3613 4893 3627 4907
rect 3593 4793 3607 4807
rect 3633 4753 3647 4767
rect 3573 4453 3587 4467
rect 3573 4413 3587 4427
rect 3573 4373 3587 4387
rect 3553 4153 3567 4167
rect 3553 4053 3567 4067
rect 3533 4033 3547 4047
rect 3413 3833 3427 3847
rect 3393 3572 3407 3586
rect 3373 3516 3387 3530
rect 3513 3990 3527 4004
rect 3473 3953 3487 3967
rect 3673 4673 3687 4687
rect 3713 4993 3727 5007
rect 3753 5053 3767 5067
rect 3773 4993 3787 5007
rect 3813 4953 3827 4967
rect 3793 4913 3807 4927
rect 3773 4833 3787 4847
rect 3753 4793 3767 4807
rect 3733 4753 3747 4767
rect 3753 4733 3767 4747
rect 3733 4673 3747 4687
rect 3713 4653 3727 4667
rect 3713 4613 3727 4627
rect 3653 4573 3667 4587
rect 3693 4573 3707 4587
rect 3733 4593 3747 4607
rect 3653 4533 3667 4547
rect 3633 4513 3647 4527
rect 3693 4510 3707 4524
rect 3653 4336 3667 4350
rect 3713 4333 3727 4347
rect 3653 4273 3667 4287
rect 3633 4233 3647 4247
rect 3653 4213 3667 4227
rect 3653 4113 3667 4127
rect 3633 4093 3647 4107
rect 3553 3973 3567 3987
rect 3513 3913 3527 3927
rect 3573 3853 3587 3867
rect 3673 4036 3687 4050
rect 3793 4290 3807 4304
rect 3773 4273 3787 4287
rect 4013 5373 4027 5387
rect 4053 5813 4067 5827
rect 4073 5793 4087 5807
rect 4073 5653 4087 5667
rect 4073 5550 4087 5564
rect 4093 5513 4107 5527
rect 4073 5493 4087 5507
rect 4053 5453 4067 5467
rect 4033 5333 4047 5347
rect 4013 5273 4027 5287
rect 4133 5873 4147 5887
rect 4193 6333 4207 6347
rect 4193 6253 4207 6267
rect 4173 6193 4187 6207
rect 4173 6133 4187 6147
rect 4173 6093 4187 6107
rect 4193 6070 4207 6084
rect 4173 5913 4187 5927
rect 4353 7233 4367 7247
rect 4493 7913 4507 7927
rect 4553 7913 4567 7927
rect 4493 7733 4507 7747
rect 4653 8133 4667 8147
rect 4753 8450 4767 8464
rect 4893 8453 4907 8467
rect 4813 8433 4827 8447
rect 4933 8653 4947 8667
rect 4713 8413 4727 8427
rect 4913 8413 4927 8427
rect 4793 8353 4807 8367
rect 4733 8233 4747 8247
rect 4773 8233 4787 8247
rect 4773 8153 4787 8167
rect 4873 8196 4887 8210
rect 4853 8150 4867 8164
rect 4793 8093 4807 8107
rect 4653 8053 4667 8067
rect 4773 7950 4787 7964
rect 5073 8716 5087 8730
rect 5253 9373 5267 9387
rect 5173 9353 5187 9367
rect 5153 8713 5167 8727
rect 4953 8633 4967 8647
rect 4953 8593 4967 8607
rect 4993 8496 5007 8510
rect 4933 8393 4947 8407
rect 4913 8133 4927 8147
rect 5093 8670 5107 8684
rect 5193 9253 5207 9267
rect 5253 9236 5267 9250
rect 5253 9193 5267 9207
rect 5193 8933 5207 8947
rect 5293 9413 5307 9427
rect 5353 9293 5367 9307
rect 5313 9236 5327 9250
rect 5373 9153 5387 9167
rect 5333 9113 5347 9127
rect 5493 11133 5507 11147
rect 5533 10973 5547 10987
rect 5493 10913 5507 10927
rect 5473 10873 5487 10887
rect 5473 10793 5487 10807
rect 5453 10613 5467 10627
rect 5433 10433 5447 10447
rect 5433 10193 5447 10207
rect 5413 9073 5427 9087
rect 5293 9033 5307 9047
rect 5353 9016 5367 9030
rect 5293 8953 5307 8967
rect 5333 8953 5347 8967
rect 5193 8773 5207 8787
rect 5213 8713 5227 8727
rect 5213 8633 5227 8647
rect 5513 10813 5527 10827
rect 5753 11153 5767 11167
rect 5753 11096 5767 11110
rect 5793 11096 5807 11110
rect 5773 11050 5787 11064
rect 5673 10953 5687 10967
rect 5613 10853 5627 10867
rect 5933 11253 5947 11267
rect 6033 11553 6047 11567
rect 5992 11093 6006 11107
rect 6013 11096 6027 11110
rect 5993 11050 6007 11064
rect 5913 10913 5927 10927
rect 5993 10873 6007 10887
rect 5973 10813 5987 10827
rect 5693 10773 5707 10787
rect 5533 10753 5547 10767
rect 5513 10693 5527 10707
rect 5513 10653 5527 10667
rect 5493 10530 5507 10544
rect 5473 10233 5487 10247
rect 5673 10733 5687 10747
rect 5593 10693 5607 10707
rect 5553 10653 5567 10667
rect 5673 10653 5687 10667
rect 5593 10613 5607 10627
rect 5553 10573 5567 10587
rect 5633 10593 5647 10607
rect 5693 10576 5707 10590
rect 5613 10530 5627 10544
rect 5553 10493 5567 10507
rect 5653 10493 5667 10507
rect 5593 10473 5607 10487
rect 5553 10453 5567 10467
rect 5533 10413 5547 10427
rect 5553 10393 5567 10407
rect 5573 10373 5587 10387
rect 5833 10776 5847 10790
rect 5973 10733 5987 10747
rect 5973 10673 5987 10687
rect 5753 10653 5767 10667
rect 5593 10293 5607 10307
rect 5613 10276 5627 10290
rect 5653 10276 5667 10290
rect 5513 10193 5527 10207
rect 5553 10193 5567 10207
rect 5693 10273 5707 10287
rect 5693 10233 5707 10247
rect 5693 10173 5707 10187
rect 5593 10153 5607 10167
rect 5593 10093 5607 10107
rect 5453 10056 5467 10070
rect 5553 10056 5567 10070
rect 5433 8933 5447 8947
rect 5433 8912 5447 8926
rect 5273 8892 5287 8906
rect 5373 8893 5387 8907
rect 5413 8893 5427 8907
rect 5253 8793 5267 8807
rect 5373 8853 5387 8867
rect 5353 8733 5367 8747
rect 5313 8716 5327 8730
rect 5493 10033 5507 10047
rect 5473 9933 5487 9947
rect 5713 10093 5727 10107
rect 5613 10010 5627 10024
rect 5653 10010 5667 10024
rect 5693 10010 5707 10024
rect 5573 9953 5587 9967
rect 5513 9813 5527 9827
rect 5493 9753 5507 9767
rect 5673 9893 5687 9907
rect 5713 9853 5727 9867
rect 5673 9833 5687 9847
rect 5513 9713 5527 9727
rect 5493 9653 5507 9667
rect 5653 9713 5667 9727
rect 5633 9653 5647 9667
rect 5673 9653 5687 9667
rect 5593 9613 5607 9627
rect 5573 9573 5587 9587
rect 5473 9553 5487 9567
rect 5513 9553 5527 9567
rect 5553 9553 5567 9567
rect 5493 9493 5507 9507
rect 5473 9013 5487 9027
rect 5473 8973 5487 8987
rect 5473 8952 5487 8966
rect 5453 8853 5467 8867
rect 5433 8833 5447 8847
rect 5473 8793 5487 8807
rect 5413 8773 5427 8787
rect 5533 9433 5547 9447
rect 5513 9153 5527 9167
rect 5513 9053 5527 9067
rect 5513 8993 5527 9007
rect 5773 10633 5787 10647
rect 5813 10613 5827 10627
rect 5913 10613 5927 10627
rect 5793 10573 5807 10587
rect 5773 10272 5787 10286
rect 5753 10193 5767 10207
rect 5873 10576 5887 10590
rect 5953 10533 5967 10547
rect 5893 10473 5907 10487
rect 5813 10433 5827 10447
rect 5853 10276 5867 10290
rect 5893 10276 5907 10290
rect 5933 10276 5947 10290
rect 5793 10230 5807 10244
rect 5833 10230 5847 10244
rect 5793 10193 5807 10207
rect 5833 10193 5847 10207
rect 5873 10193 5887 10207
rect 5733 9490 5747 9504
rect 5733 9373 5747 9387
rect 5653 9353 5667 9367
rect 5613 9333 5627 9347
rect 5573 9253 5587 9267
rect 5593 9133 5607 9147
rect 5773 10056 5787 10070
rect 5733 9113 5747 9127
rect 5573 9033 5587 9047
rect 5613 9016 5627 9030
rect 5633 8970 5647 8984
rect 5733 8970 5747 8984
rect 5593 8953 5607 8967
rect 5933 10173 5947 10187
rect 6153 11533 6167 11547
rect 6213 11793 6227 11807
rect 6273 11713 6287 11727
rect 6213 11553 6227 11567
rect 6293 11553 6307 11567
rect 6413 11973 6427 11987
rect 6373 11873 6387 11887
rect 6793 12153 6807 12167
rect 6933 12153 6947 12167
rect 8353 12153 8367 12167
rect 8453 12153 8467 12167
rect 6713 12113 6727 12127
rect 6912 12116 6926 12130
rect 7753 12136 7767 12150
rect 7953 12136 7967 12150
rect 6933 12110 6947 12124
rect 7033 12110 7047 12124
rect 7193 12116 7207 12130
rect 7233 12116 7247 12130
rect 7293 12116 7307 12130
rect 7333 12116 7347 12130
rect 6693 12013 6707 12027
rect 6673 11973 6687 11987
rect 6533 11933 6547 11947
rect 6493 11913 6507 11927
rect 6453 11836 6467 11850
rect 6533 11836 6547 11850
rect 6633 11836 6647 11850
rect 6373 11793 6387 11807
rect 6413 11793 6427 11807
rect 6513 11790 6527 11804
rect 6533 11773 6547 11787
rect 6373 11633 6387 11647
rect 6473 11633 6487 11647
rect 6333 11533 6347 11547
rect 6493 11533 6507 11547
rect 6173 11413 6187 11427
rect 6373 11413 6387 11427
rect 6113 11316 6127 11330
rect 6073 11153 6087 11167
rect 6093 11133 6107 11147
rect 6133 11096 6147 11110
rect 6073 11050 6087 11064
rect 6113 11013 6127 11027
rect 6153 10953 6167 10967
rect 6113 10933 6127 10947
rect 6033 10853 6047 10867
rect 6253 11373 6267 11387
rect 6193 11353 6207 11367
rect 6173 10933 6187 10947
rect 6153 10893 6167 10907
rect 6013 10813 6027 10827
rect 6113 10813 6127 10827
rect 6293 11313 6307 11327
rect 6333 11316 6347 11330
rect 6353 11270 6367 11284
rect 6313 11093 6327 11107
rect 6453 11213 6467 11227
rect 6393 11096 6407 11110
rect 6553 11570 6567 11584
rect 6633 11433 6647 11447
rect 6553 11373 6567 11387
rect 6593 11333 6607 11347
rect 7193 12073 7207 12087
rect 6873 12053 6887 12067
rect 6813 12033 6827 12047
rect 6853 12033 6867 12047
rect 6793 11913 6807 11927
rect 6773 11893 6787 11907
rect 6713 11836 6727 11850
rect 6753 11836 6767 11850
rect 6873 11993 6887 12007
rect 6933 11993 6947 12007
rect 6773 11790 6787 11804
rect 6713 11773 6727 11787
rect 6853 11793 6867 11807
rect 6813 11753 6827 11767
rect 6713 11733 6727 11747
rect 6693 11353 6707 11367
rect 6673 11333 6687 11347
rect 6613 11270 6627 11284
rect 6693 11273 6707 11287
rect 6813 11713 6827 11727
rect 6773 11673 6787 11687
rect 6793 11570 6807 11584
rect 6713 11233 6727 11247
rect 6513 11213 6527 11227
rect 6493 11153 6507 11167
rect 6473 11133 6487 11147
rect 6893 11473 6907 11487
rect 6953 11973 6967 11987
rect 7513 11993 7527 12007
rect 7293 11953 7307 11967
rect 7333 11953 7347 11967
rect 6953 11836 6967 11850
rect 7053 11836 7067 11850
rect 7093 11836 7107 11850
rect 7293 11836 7307 11850
rect 7333 11836 7347 11850
rect 6933 11313 6947 11327
rect 6873 11253 6887 11267
rect 6793 11173 6807 11187
rect 6493 11073 6507 11087
rect 6573 11070 6587 11084
rect 6713 11070 6727 11084
rect 6833 11076 6847 11090
rect 6913 11073 6927 11087
rect 6333 11050 6347 11064
rect 6413 11050 6427 11064
rect 6473 11033 6487 11047
rect 6313 11013 6327 11027
rect 6193 10833 6207 10847
rect 6013 10773 6027 10787
rect 5993 10593 6007 10607
rect 5973 10273 5987 10287
rect 5833 10010 5847 10024
rect 5953 10013 5967 10027
rect 5873 9953 5887 9967
rect 5833 9813 5847 9827
rect 5913 9933 5927 9947
rect 5853 9710 5867 9724
rect 5973 9893 5987 9907
rect 5913 9573 5927 9587
rect 5913 9536 5927 9550
rect 6033 10733 6047 10747
rect 6033 10693 6047 10707
rect 6033 10513 6047 10527
rect 6013 10233 6027 10247
rect 6113 10773 6127 10787
rect 6173 10773 6187 10787
rect 6093 10493 6107 10507
rect 6073 10453 6087 10467
rect 6173 10693 6187 10707
rect 6313 10776 6327 10790
rect 6452 10776 6466 10790
rect 6873 11030 6887 11044
rect 6473 10770 6487 10784
rect 6513 10770 6527 10784
rect 6573 10770 6587 10784
rect 6513 10733 6527 10747
rect 6473 10713 6487 10727
rect 6193 10673 6207 10687
rect 6313 10653 6327 10667
rect 6513 10653 6527 10667
rect 6133 10613 6147 10627
rect 6173 10593 6187 10607
rect 6253 10556 6267 10570
rect 6353 10550 6367 10564
rect 6513 10550 6527 10564
rect 7253 11813 7267 11827
rect 7073 11790 7087 11804
rect 7313 11773 7327 11787
rect 7053 11753 7067 11767
rect 7253 11753 7267 11767
rect 7333 11753 7347 11767
rect 7013 11673 7027 11687
rect 7153 11733 7167 11747
rect 7093 11693 7107 11707
rect 7293 11653 7307 11667
rect 7293 11613 7307 11627
rect 7373 11616 7387 11630
rect 7473 11593 7487 11607
rect 7113 11570 7127 11584
rect 7153 11570 7167 11584
rect 7013 11533 7027 11547
rect 7073 11533 7087 11547
rect 6973 11513 6987 11527
rect 7353 11493 7367 11507
rect 7473 11533 7487 11547
rect 7393 11473 7407 11487
rect 7013 11433 7027 11447
rect 7073 11433 7087 11447
rect 6973 11270 6987 11284
rect 6953 11253 6967 11267
rect 6993 11173 7007 11187
rect 6973 11093 6987 11107
rect 6953 11053 6967 11067
rect 6933 11030 6947 11044
rect 6733 10893 6747 10907
rect 6873 10893 6887 10907
rect 6933 10893 6947 10907
rect 6653 10833 6667 10847
rect 6653 10770 6667 10784
rect 6713 10653 6727 10667
rect 6193 10513 6207 10527
rect 6153 10493 6167 10507
rect 6193 10492 6207 10506
rect 6073 10313 6087 10327
rect 6153 10333 6167 10347
rect 6153 10276 6167 10290
rect 6293 10433 6307 10447
rect 6353 10413 6367 10427
rect 6293 10393 6307 10407
rect 6673 10413 6687 10427
rect 6773 10793 6787 10807
rect 6833 10796 6847 10810
rect 6733 10413 6747 10427
rect 6813 10673 6827 10687
rect 6813 10633 6827 10647
rect 6853 10633 6867 10647
rect 6793 10533 6807 10547
rect 6933 10613 6947 10627
rect 6913 10576 6927 10590
rect 6973 10833 6987 10847
rect 6813 10493 6827 10507
rect 6793 10333 6807 10347
rect 6773 10313 6787 10327
rect 6693 10273 6707 10287
rect 6773 10276 6787 10290
rect 6153 10173 6167 10187
rect 6093 10093 6107 10107
rect 6293 10250 6307 10264
rect 6333 10256 6347 10270
rect 6493 10256 6507 10270
rect 6253 10233 6267 10247
rect 6233 10173 6247 10187
rect 6233 10093 6247 10107
rect 6173 10073 6187 10087
rect 6213 10073 6227 10087
rect 6093 10010 6107 10024
rect 6033 9893 6047 9907
rect 5893 9490 5907 9504
rect 5953 9493 5967 9507
rect 5993 9493 6007 9507
rect 5933 9433 5947 9447
rect 5793 9373 5807 9387
rect 5873 9273 5887 9287
rect 5833 9236 5847 9250
rect 5913 9236 5927 9250
rect 5853 9190 5867 9204
rect 5913 9093 5927 9107
rect 5873 8970 5887 8984
rect 5813 8933 5827 8947
rect 5773 8913 5787 8927
rect 5813 8813 5827 8827
rect 5513 8753 5527 8767
rect 5493 8733 5507 8747
rect 5373 8713 5387 8727
rect 5393 8693 5407 8707
rect 5333 8670 5347 8684
rect 5273 8633 5287 8647
rect 5233 8533 5247 8547
rect 5213 8513 5227 8527
rect 5193 8496 5207 8510
rect 5253 8496 5267 8510
rect 5153 8353 5167 8367
rect 5133 8333 5147 8347
rect 5053 8293 5067 8307
rect 5093 8273 5107 8287
rect 5053 8253 5067 8267
rect 4993 8196 5007 8210
rect 5033 8196 5047 8210
rect 5033 8153 5047 8167
rect 4993 8033 5007 8047
rect 4953 7953 4967 7967
rect 4993 7956 5007 7970
rect 5093 8233 5107 8247
rect 5093 8196 5107 8210
rect 5092 8133 5106 8147
rect 5113 8133 5127 8147
rect 4933 7910 4947 7924
rect 4973 7913 4987 7927
rect 4753 7853 4767 7867
rect 4613 7813 4627 7827
rect 4713 7813 4727 7827
rect 4613 7792 4627 7806
rect 4633 7630 4647 7644
rect 4593 7593 4607 7607
rect 4633 7593 4647 7607
rect 4553 7573 4567 7587
rect 4533 7495 4547 7509
rect 4513 7410 4527 7424
rect 4453 7393 4467 7407
rect 4553 7393 4567 7407
rect 4613 7233 4627 7247
rect 4393 7213 4407 7227
rect 4433 7213 4447 7227
rect 4353 7109 4367 7123
rect 4553 7109 4567 7123
rect 4513 7071 4527 7085
rect 4493 6910 4507 6924
rect 4653 7573 4667 7587
rect 4693 7573 4707 7587
rect 4633 7113 4647 7127
rect 4633 7053 4647 7067
rect 4693 7453 4707 7467
rect 4673 7393 4687 7407
rect 4653 6933 4667 6947
rect 4693 6953 4707 6967
rect 4633 6910 4647 6924
rect 4673 6913 4687 6927
rect 4693 6893 4707 6907
rect 4673 6873 4687 6887
rect 4653 6853 4667 6867
rect 4473 6813 4487 6827
rect 4333 6713 4347 6727
rect 4453 6713 4467 6727
rect 4393 6673 4407 6687
rect 4233 6636 4247 6650
rect 4293 6590 4307 6604
rect 4253 6473 4267 6487
rect 4253 6333 4267 6347
rect 4233 6213 4247 6227
rect 4333 6553 4347 6567
rect 4353 6453 4367 6467
rect 4313 6413 4327 6427
rect 4393 6416 4407 6430
rect 4293 6373 4307 6387
rect 4273 6173 4287 6187
rect 4373 6370 4387 6384
rect 4373 6333 4387 6347
rect 4333 6133 4347 6147
rect 4313 6093 4327 6107
rect 4253 6070 4267 6084
rect 4333 6073 4347 6087
rect 4413 6273 4427 6287
rect 4253 5973 4267 5987
rect 4352 5973 4366 5987
rect 4373 5973 4387 5987
rect 4453 6253 4467 6267
rect 4433 6173 4447 6187
rect 4273 5893 4287 5907
rect 4313 5913 4327 5927
rect 4393 5913 4407 5927
rect 4353 5896 4367 5910
rect 4253 5813 4267 5827
rect 4213 5753 4227 5767
rect 4173 5693 4187 5707
rect 4133 5493 4147 5507
rect 4113 5413 4127 5427
rect 4253 5693 4267 5707
rect 4213 5673 4227 5687
rect 4253 5633 4267 5647
rect 4253 5593 4267 5607
rect 4313 5813 4327 5827
rect 4293 5653 4307 5667
rect 4293 5613 4307 5627
rect 4273 5553 4287 5567
rect 4253 5513 4267 5527
rect 4233 5493 4247 5507
rect 4233 5413 4247 5427
rect 4173 5393 4187 5407
rect 4073 5376 4087 5390
rect 4153 5376 4167 5390
rect 4193 5376 4207 5390
rect 4173 5330 4187 5344
rect 4233 5333 4247 5347
rect 4093 5233 4107 5247
rect 4053 5213 4067 5227
rect 3913 5193 3927 5207
rect 4093 5193 4107 5207
rect 4153 5213 4167 5227
rect 4133 5113 4147 5127
rect 3853 5093 3867 5107
rect 4213 5113 4227 5127
rect 3993 5056 4007 5070
rect 4173 5053 4187 5067
rect 3853 5013 3867 5027
rect 4033 4953 4047 4967
rect 3933 4933 3947 4947
rect 3933 4873 3947 4887
rect 3993 4873 4007 4887
rect 3893 4856 3907 4870
rect 3973 4853 3987 4867
rect 3873 4773 3887 4787
rect 3973 4773 3987 4787
rect 3853 4753 3867 4767
rect 3913 4753 3927 4767
rect 3853 4732 3867 4746
rect 3833 4273 3847 4287
rect 3773 4233 3787 4247
rect 3793 4153 3807 4167
rect 3752 4113 3766 4127
rect 3773 4113 3787 4127
rect 3753 4036 3767 4050
rect 3653 3990 3667 4004
rect 3793 4033 3807 4047
rect 3733 3990 3747 4004
rect 3672 3953 3686 3967
rect 3693 3953 3707 3967
rect 3633 3733 3647 3747
rect 3653 3713 3667 3727
rect 3553 3693 3567 3707
rect 3593 3693 3607 3707
rect 3553 3653 3567 3667
rect 3433 3633 3447 3647
rect 3393 3296 3407 3310
rect 3533 3516 3547 3530
rect 3493 3433 3507 3447
rect 3533 3413 3547 3427
rect 3513 3393 3527 3407
rect 3533 3353 3547 3367
rect 3353 3113 3367 3127
rect 3373 3053 3387 3067
rect 3353 2953 3367 2967
rect 3333 2913 3347 2927
rect 3273 2873 3287 2887
rect 3073 2813 3087 2827
rect 3053 2773 3067 2787
rect 3433 3153 3447 3167
rect 3513 3113 3527 3127
rect 3453 3053 3467 3067
rect 3473 3033 3487 3047
rect 3433 2933 3447 2947
rect 3413 2873 3427 2887
rect 3433 2853 3447 2867
rect 3433 2773 3447 2787
rect 3233 2750 3247 2764
rect 3353 2756 3367 2770
rect 3433 2752 3447 2766
rect 3073 2733 3087 2747
rect 2913 2713 2927 2727
rect 2893 2693 2907 2707
rect 2853 2553 2867 2567
rect 2873 2533 2887 2547
rect 2893 2473 2907 2487
rect 2893 2333 2907 2347
rect 2893 2293 2907 2307
rect 2873 2273 2887 2287
rect 2993 2653 3007 2667
rect 2972 2476 2986 2490
rect 3033 2613 3047 2627
rect 3453 2673 3467 2687
rect 3593 3133 3607 3147
rect 3553 2993 3567 3007
rect 3493 2933 3507 2947
rect 3473 2653 3487 2667
rect 3433 2613 3447 2627
rect 3073 2533 3087 2547
rect 3353 2513 3367 2527
rect 2993 2473 3007 2487
rect 2953 2430 2967 2444
rect 2953 2393 2967 2407
rect 2993 2353 3007 2367
rect 2933 2333 2947 2347
rect 2913 2273 2927 2287
rect 2973 2273 2987 2287
rect 2913 2210 2927 2224
rect 2973 2213 2987 2227
rect 2873 2073 2887 2087
rect 2833 1976 2847 1990
rect 2913 2073 2927 2087
rect 2713 1733 2727 1747
rect 2593 1493 2607 1507
rect 2653 1653 2667 1667
rect 2733 1633 2747 1647
rect 2693 1613 2707 1627
rect 2733 1473 2747 1487
rect 2633 1433 2647 1447
rect 2613 1390 2627 1404
rect 2613 1253 2627 1267
rect 2613 1173 2627 1187
rect 2533 1113 2547 1127
rect 2513 1033 2527 1047
rect 2573 993 2587 1007
rect 2433 915 2447 929
rect 2493 831 2507 845
rect 2573 833 2587 847
rect 2553 813 2567 827
rect 2693 1390 2707 1404
rect 2693 1253 2707 1267
rect 2733 1216 2747 1230
rect 2713 1133 2727 1147
rect 2833 1955 2847 1969
rect 2953 2013 2967 2027
rect 2932 1973 2946 1987
rect 2953 1973 2967 1987
rect 2793 1913 2807 1927
rect 2773 993 2787 1007
rect 2853 1910 2867 1924
rect 2913 1913 2927 1927
rect 3193 2456 3207 2470
rect 3453 2450 3467 2464
rect 3353 2433 3367 2447
rect 3393 2433 3407 2447
rect 3453 2413 3467 2427
rect 3333 2273 3347 2287
rect 3193 2256 3207 2270
rect 3233 2256 3247 2270
rect 3153 2210 3167 2224
rect 3293 2133 3307 2147
rect 3233 2053 3247 2067
rect 3193 2013 3207 2027
rect 3173 1993 3187 2007
rect 3133 1956 3147 1970
rect 3193 1956 3207 1970
rect 2993 1853 3007 1867
rect 2853 1833 2867 1847
rect 2933 1833 2947 1847
rect 2833 1473 2847 1487
rect 2833 1170 2847 1184
rect 2953 1813 2967 1827
rect 2913 1736 2927 1750
rect 2873 1573 2887 1587
rect 2893 1553 2907 1567
rect 2873 1513 2887 1527
rect 2973 1690 2987 1704
rect 3013 1693 3027 1707
rect 3153 1910 3167 1924
rect 3173 1893 3187 1907
rect 3233 1893 3247 1907
rect 2973 1593 2987 1607
rect 2933 1493 2947 1507
rect 2973 1436 2987 1450
rect 3113 1690 3127 1704
rect 3153 1633 3167 1647
rect 3033 1513 3047 1527
rect 3153 1493 3167 1507
rect 3033 1433 3047 1447
rect 3073 1410 3087 1424
rect 2873 1390 2887 1404
rect 2953 1390 2967 1404
rect 2993 1313 3007 1327
rect 3153 1416 3167 1430
rect 3133 1333 3147 1347
rect 3153 1313 3167 1327
rect 3073 1273 3087 1287
rect 2933 1213 2947 1227
rect 2993 1216 3007 1230
rect 3053 1213 3067 1227
rect 2973 1170 2987 1184
rect 3013 1170 3027 1184
rect 2933 1133 2947 1147
rect 2853 1013 2867 1027
rect 2793 973 2807 987
rect 2853 973 2867 987
rect 2713 933 2727 947
rect 2773 933 2787 947
rect 2813 916 2827 930
rect 2713 853 2727 867
rect 2753 793 2767 807
rect 2633 773 2647 787
rect 2773 733 2787 747
rect 2533 696 2547 710
rect 2593 696 2607 710
rect 2633 696 2647 710
rect 2693 696 2707 710
rect 2533 613 2547 627
rect 2613 650 2627 664
rect 2573 553 2587 567
rect 2773 650 2787 664
rect 2653 533 2667 547
rect 2573 493 2587 507
rect 2393 416 2407 430
rect 3113 1216 3127 1230
rect 3073 1170 3087 1184
rect 2993 1013 3007 1027
rect 3033 1013 3047 1027
rect 2873 916 2887 930
rect 2973 916 2987 930
rect 2873 873 2887 887
rect 2973 793 2987 807
rect 2893 753 2907 767
rect 2933 696 2947 710
rect 2973 693 2987 707
rect 2853 653 2867 667
rect 2693 413 2707 427
rect 2793 413 2807 427
rect 2333 396 2347 410
rect 2233 350 2247 364
rect 2273 353 2287 367
rect 2353 333 2367 347
rect 2273 293 2287 307
rect 2553 376 2567 390
rect 2693 376 2707 390
rect 2753 353 2767 367
rect 2813 353 2827 367
rect 2753 313 2767 327
rect 2433 273 2447 287
rect 2493 273 2507 287
rect 2353 253 2367 267
rect 2333 150 2347 164
rect 2013 130 2027 144
rect 2073 130 2087 144
rect 2173 110 2187 124
rect 1733 93 1747 107
rect 2113 93 2127 107
rect 1173 33 1187 47
rect 2593 253 2607 267
rect 2533 156 2547 170
rect 2773 233 2787 247
rect 2753 156 2767 170
rect 2873 650 2887 664
rect 2913 650 2927 664
rect 2953 653 2967 667
rect 2973 613 2987 627
rect 3073 916 3087 930
rect 3133 993 3147 1007
rect 3113 913 3127 927
rect 3053 870 3067 884
rect 3113 773 3127 787
rect 3113 733 3127 747
rect 3113 650 3127 664
rect 3233 1736 3247 1750
rect 3313 2113 3327 2127
rect 3313 1813 3327 1827
rect 3213 1653 3227 1667
rect 3513 2913 3527 2927
rect 3493 2333 3507 2347
rect 3533 2873 3547 2887
rect 3513 2273 3527 2287
rect 3493 2256 3507 2270
rect 3473 2210 3487 2224
rect 3433 2173 3447 2187
rect 3493 2113 3507 2127
rect 3473 2013 3487 2027
rect 3453 1956 3467 1970
rect 3513 2053 3527 2067
rect 3573 2913 3587 2927
rect 3553 2673 3567 2687
rect 3553 2513 3567 2527
rect 3553 2450 3567 2464
rect 3553 2256 3567 2270
rect 3553 2213 3567 2227
rect 3553 2173 3567 2187
rect 3533 1993 3547 2007
rect 3533 1972 3547 1986
rect 3433 1910 3447 1924
rect 3493 1910 3507 1924
rect 3493 1773 3507 1787
rect 3633 3516 3647 3530
rect 3633 3473 3647 3487
rect 3633 3193 3647 3207
rect 3653 3173 3667 3187
rect 3633 3113 3647 3127
rect 3673 3133 3687 3147
rect 3673 2953 3687 2967
rect 3773 3933 3787 3947
rect 4013 4853 4027 4867
rect 3993 4633 4007 4647
rect 3873 4613 3887 4627
rect 3953 4613 3967 4627
rect 3893 4553 3907 4567
rect 4073 4933 4087 4947
rect 4033 4553 4047 4567
rect 3893 4510 3907 4524
rect 3933 4510 3947 4524
rect 3913 4453 3927 4467
rect 3873 4373 3887 4387
rect 3973 4433 3987 4447
rect 3992 4373 4006 4387
rect 4013 4373 4027 4387
rect 3873 4272 3887 4286
rect 3893 4233 3907 4247
rect 3893 4133 3907 4147
rect 3913 4053 3927 4067
rect 3873 3953 3887 3967
rect 3893 3913 3907 3927
rect 3893 3873 3907 3887
rect 3853 3853 3867 3867
rect 3753 3770 3767 3784
rect 3813 3770 3827 3784
rect 3853 3770 3867 3784
rect 3733 3493 3747 3507
rect 3713 3333 3727 3347
rect 3893 3613 3907 3627
rect 3893 3573 3907 3587
rect 3793 3553 3807 3567
rect 3833 3516 3847 3530
rect 3893 3516 3907 3530
rect 3813 3470 3827 3484
rect 3853 3470 3867 3484
rect 3953 4093 3967 4107
rect 4013 4213 4027 4227
rect 3993 4053 4007 4067
rect 3973 3993 3987 4007
rect 3953 3973 3967 3987
rect 3933 3633 3947 3647
rect 3913 3470 3927 3484
rect 3893 3413 3907 3427
rect 3833 3373 3847 3387
rect 3753 3296 3767 3310
rect 3773 3250 3787 3264
rect 3953 3553 3967 3567
rect 3953 3513 3967 3527
rect 3893 3353 3907 3367
rect 3933 3353 3947 3367
rect 3873 3293 3887 3307
rect 3733 3193 3747 3207
rect 3833 3193 3847 3207
rect 3733 3053 3747 3067
rect 3773 2996 3787 3010
rect 3753 2950 3767 2964
rect 3853 3093 3867 3107
rect 3693 2873 3707 2887
rect 3733 2873 3747 2887
rect 3653 2813 3667 2827
rect 3653 2776 3667 2790
rect 3773 2813 3787 2827
rect 3633 2730 3647 2744
rect 3733 2733 3747 2747
rect 3633 2673 3647 2687
rect 3773 2633 3787 2647
rect 3633 2553 3647 2567
rect 3713 2476 3727 2490
rect 3813 2553 3827 2567
rect 3793 2476 3807 2490
rect 3633 2313 3647 2327
rect 3733 2413 3747 2427
rect 3773 2413 3787 2427
rect 3613 2253 3627 2267
rect 3693 2253 3707 2267
rect 3593 2053 3607 2067
rect 3593 1993 3607 2007
rect 3573 1956 3587 1970
rect 3533 1753 3547 1767
rect 3393 1690 3407 1704
rect 3473 1690 3487 1704
rect 3513 1593 3527 1607
rect 3393 1553 3407 1567
rect 3513 1533 3527 1547
rect 3333 1513 3347 1527
rect 3193 1456 3207 1470
rect 3493 1456 3507 1470
rect 3333 1416 3347 1430
rect 3453 1410 3467 1424
rect 3533 1413 3547 1427
rect 3193 1373 3207 1387
rect 3453 1373 3467 1387
rect 3573 1373 3587 1387
rect 3253 1313 3267 1327
rect 3333 1253 3347 1267
rect 3293 1216 3307 1230
rect 3273 1170 3287 1184
rect 3333 1170 3347 1184
rect 3313 1113 3327 1127
rect 3253 953 3267 967
rect 3353 953 3367 967
rect 3253 870 3267 884
rect 3213 753 3227 767
rect 3173 696 3187 710
rect 3193 650 3207 664
rect 3293 870 3307 884
rect 3333 833 3347 847
rect 3553 1255 3567 1269
rect 3593 1217 3607 1231
rect 3473 1133 3487 1147
rect 3713 2210 3727 2224
rect 3793 2253 3807 2267
rect 3833 2193 3847 2207
rect 3793 2153 3807 2167
rect 3773 2113 3787 2127
rect 3833 2093 3847 2107
rect 3773 2053 3787 2067
rect 3653 2033 3667 2047
rect 3713 1893 3727 1907
rect 3753 1893 3767 1907
rect 3653 1753 3667 1767
rect 3793 1853 3807 1867
rect 3833 1813 3847 1827
rect 3773 1773 3787 1787
rect 3693 1736 3707 1750
rect 3733 1736 3747 1750
rect 3653 1693 3667 1707
rect 3793 1690 3807 1704
rect 3833 1613 3847 1627
rect 3693 1573 3707 1587
rect 3753 1573 3767 1587
rect 3673 1493 3687 1507
rect 3753 1493 3767 1507
rect 3793 1436 3807 1450
rect 3693 1390 3707 1404
rect 3733 1390 3747 1404
rect 3673 1313 3687 1327
rect 3633 1153 3647 1167
rect 3613 953 3627 967
rect 3593 916 3607 930
rect 4033 3933 4047 3947
rect 4093 4893 4107 4907
rect 4073 3913 4087 3927
rect 4193 4993 4207 5007
rect 4213 4953 4227 4967
rect 4173 4933 4187 4947
rect 4233 4893 4247 4907
rect 4133 4853 4147 4867
rect 4173 4856 4187 4870
rect 4133 4813 4147 4827
rect 4293 5513 4307 5527
rect 4273 5373 4287 5387
rect 4333 5473 4347 5487
rect 4313 5293 4327 5307
rect 4313 5092 4327 5106
rect 4293 5073 4307 5087
rect 4273 5053 4287 5067
rect 4293 5033 4307 5047
rect 4273 4953 4287 4967
rect 4153 4793 4167 4807
rect 4193 4793 4207 4807
rect 4153 4556 4167 4570
rect 4133 4493 4147 4507
rect 4133 4472 4147 4486
rect 4153 4433 4167 4447
rect 4133 4336 4147 4350
rect 4153 4273 4167 4287
rect 4153 4173 4167 4187
rect 4173 4033 4187 4047
rect 4113 3993 4127 4007
rect 4013 3833 4027 3847
rect 4093 3833 4107 3847
rect 4053 3816 4067 3830
rect 4113 3816 4127 3830
rect 4013 3770 4027 3784
rect 4133 3773 4147 3787
rect 4173 3773 4187 3787
rect 4153 3753 4167 3767
rect 4093 3733 4107 3747
rect 4013 3653 4027 3667
rect 4053 3653 4067 3667
rect 4013 3573 4027 3587
rect 4073 3516 4087 3530
rect 4033 3493 4047 3507
rect 3993 3373 4007 3387
rect 3933 3313 3947 3327
rect 3973 3313 3987 3327
rect 3913 3293 3927 3307
rect 3913 3213 3927 3227
rect 3893 3033 3907 3047
rect 3913 3013 3927 3027
rect 3873 2950 3887 2964
rect 4113 3433 4127 3447
rect 4033 3296 4047 3310
rect 4093 3293 4107 3307
rect 3973 3250 3987 3264
rect 3953 3153 3967 3167
rect 4053 3250 4067 3264
rect 4053 3193 4067 3207
rect 4093 3093 4107 3107
rect 4133 3413 4147 3427
rect 4113 3073 4127 3087
rect 4013 3053 4027 3067
rect 4013 3013 4027 3027
rect 4053 2996 4067 3010
rect 3973 2933 3987 2947
rect 3953 2913 3967 2927
rect 3973 2833 3987 2847
rect 3893 2776 3907 2790
rect 3933 2776 3947 2790
rect 3873 2733 3887 2747
rect 3813 1153 3827 1167
rect 3973 2653 3987 2667
rect 4073 2950 4087 2964
rect 4073 2933 4087 2947
rect 4133 2933 4147 2947
rect 4073 2873 4087 2887
rect 4033 2833 4047 2847
rect 4013 2776 4027 2790
rect 4253 4793 4267 4807
rect 4233 4773 4247 4787
rect 4233 4673 4247 4687
rect 4313 4993 4327 5007
rect 4293 4753 4307 4767
rect 4313 4733 4327 4747
rect 4273 4653 4287 4667
rect 4273 4556 4287 4570
rect 4233 4473 4247 4487
rect 4293 4493 4307 4507
rect 4253 4293 4267 4307
rect 4273 4273 4287 4287
rect 4213 4073 4227 4087
rect 4193 3753 4207 3767
rect 4193 3693 4207 3707
rect 4313 4193 4327 4207
rect 4313 4153 4327 4167
rect 4213 3613 4227 3627
rect 4233 3573 4247 3587
rect 4193 3333 4207 3347
rect 4113 2833 4127 2847
rect 4113 2773 4127 2787
rect 4113 2713 4127 2727
rect 4093 2693 4107 2707
rect 4033 2593 4047 2607
rect 4013 2533 4027 2547
rect 3933 2513 3947 2527
rect 3993 2513 4007 2527
rect 3913 2476 3927 2490
rect 3913 2333 3927 2347
rect 3893 2153 3907 2167
rect 3993 2476 4007 2490
rect 4073 2553 4087 2567
rect 4013 2430 4027 2444
rect 3973 2353 3987 2367
rect 4053 2333 4067 2347
rect 3953 2256 3967 2270
rect 3993 2256 4007 2270
rect 4033 2256 4047 2270
rect 4013 2210 4027 2224
rect 4053 2210 4067 2224
rect 4093 2253 4107 2267
rect 4073 2193 4087 2207
rect 3973 1973 3987 1987
rect 4073 1913 4087 1927
rect 4013 1893 4027 1907
rect 4053 1893 4067 1907
rect 3953 1773 3967 1787
rect 3993 1773 4007 1787
rect 3893 1690 3907 1704
rect 3933 1413 3947 1427
rect 3893 1393 3907 1407
rect 3813 1132 3827 1146
rect 3873 1133 3887 1147
rect 3793 1053 3807 1067
rect 3773 973 3787 987
rect 3673 916 3687 930
rect 3573 870 3587 884
rect 3133 613 3147 627
rect 3233 613 3247 627
rect 3053 396 3067 410
rect 2993 350 3007 364
rect 3033 350 3047 364
rect 3373 653 3387 667
rect 3333 613 3347 627
rect 3253 353 3267 367
rect 3293 350 3307 364
rect 3133 333 3147 347
rect 2973 176 2987 190
rect 3053 176 3067 190
rect 3433 650 3447 664
rect 3473 613 3487 627
rect 3413 393 3427 407
rect 3413 350 3427 364
rect 3633 696 3647 710
rect 3713 913 3727 927
rect 3713 773 3727 787
rect 3733 733 3747 747
rect 3613 650 3627 664
rect 3613 593 3627 607
rect 3693 696 3707 710
rect 3853 1013 3867 1027
rect 3893 916 3907 930
rect 3913 870 3927 884
rect 4113 2233 4127 2247
rect 4093 1773 4107 1787
rect 4093 1736 4107 1750
rect 3993 1690 4007 1704
rect 4033 1690 4047 1704
rect 4093 1573 4107 1587
rect 4033 1436 4047 1450
rect 4013 1353 4027 1367
rect 4033 1273 4047 1287
rect 4053 1170 4067 1184
rect 4113 1533 4127 1547
rect 4173 2893 4187 2907
rect 4173 2813 4187 2827
rect 4233 3473 4247 3487
rect 4273 3913 4287 3927
rect 4293 3873 4307 3887
rect 4393 5612 4407 5626
rect 4373 5413 4387 5427
rect 4393 5353 4407 5367
rect 4393 5273 4407 5287
rect 4352 5193 4366 5207
rect 4373 5193 4387 5207
rect 4433 5872 4447 5886
rect 4593 6793 4607 6807
rect 4493 6636 4507 6650
rect 4653 6713 4667 6727
rect 4633 6636 4647 6650
rect 4573 6573 4587 6587
rect 4653 6573 4667 6587
rect 4613 6553 4627 6567
rect 4533 6473 4547 6487
rect 4513 6453 4527 6467
rect 4513 6333 4527 6347
rect 4493 6313 4507 6327
rect 4493 6173 4507 6187
rect 4473 6133 4487 6147
rect 4593 6413 4607 6427
rect 4673 6453 4687 6467
rect 4793 7833 4807 7847
rect 4773 7793 4787 7807
rect 4753 7752 4767 7766
rect 4733 7453 4747 7467
rect 4733 7410 4747 7424
rect 4773 7653 4787 7667
rect 4833 7773 4847 7787
rect 4853 7773 4867 7787
rect 4813 7733 4827 7747
rect 4913 7753 4927 7767
rect 5233 8433 5247 8447
rect 5273 8413 5287 8427
rect 5353 8353 5367 8367
rect 5313 8293 5327 8307
rect 5293 8253 5307 8267
rect 5233 8093 5247 8107
rect 5193 8073 5207 8087
rect 5413 8633 5427 8647
rect 5433 8613 5447 8627
rect 5413 8293 5427 8307
rect 5393 8193 5407 8207
rect 5833 8753 5847 8767
rect 5533 8733 5547 8747
rect 5813 8733 5827 8747
rect 5673 8696 5687 8710
rect 5533 8673 5547 8687
rect 5513 8653 5527 8667
rect 5813 8693 5827 8707
rect 5673 8593 5687 8607
rect 5793 8593 5807 8607
rect 5473 8533 5487 8547
rect 5553 8496 5567 8510
rect 5493 8453 5507 8467
rect 5473 8373 5487 8387
rect 5433 8233 5447 8247
rect 5533 8433 5547 8447
rect 5573 8413 5587 8427
rect 5613 8373 5627 8387
rect 5593 8353 5607 8367
rect 5573 8313 5587 8327
rect 5493 8293 5507 8307
rect 5553 8293 5567 8307
rect 5453 8213 5467 8227
rect 5493 8213 5507 8227
rect 5573 8253 5587 8267
rect 5573 8213 5587 8227
rect 5473 8153 5487 8167
rect 5433 8133 5447 8147
rect 5373 8113 5387 8127
rect 5373 8092 5387 8106
rect 5153 8053 5167 8067
rect 5313 8053 5327 8067
rect 5253 7950 5267 7964
rect 5433 8013 5447 8027
rect 5373 7893 5387 7907
rect 5413 7893 5427 7907
rect 5453 7913 5467 7927
rect 5093 7873 5107 7887
rect 5033 7793 5047 7807
rect 5053 7753 5067 7767
rect 4973 7733 4987 7747
rect 5033 7733 5047 7747
rect 4933 7693 4947 7707
rect 4813 7633 4827 7647
rect 4873 7630 4887 7644
rect 4793 7456 4807 7470
rect 4853 7433 4867 7447
rect 4753 7373 4767 7387
rect 4773 7233 4787 7247
rect 4933 7613 4947 7627
rect 4893 7410 4907 7424
rect 4873 7353 4887 7367
rect 4853 7273 4867 7287
rect 4893 7253 4907 7267
rect 4873 7133 4887 7147
rect 4733 7113 4747 7127
rect 4793 7053 4807 7067
rect 4753 6993 4767 7007
rect 4793 6973 4807 6987
rect 4773 6933 4787 6947
rect 4753 6833 4767 6847
rect 4753 6773 4767 6787
rect 4733 6713 4747 6727
rect 4853 7013 4867 7027
rect 4853 6933 4867 6947
rect 4973 7653 4987 7667
rect 5453 7872 5467 7886
rect 5433 7853 5447 7867
rect 5393 7733 5407 7747
rect 5073 7696 5087 7710
rect 5372 7696 5386 7710
rect 4953 7553 4967 7567
rect 4953 7353 4967 7367
rect 4913 7073 4927 7087
rect 5013 7650 5027 7664
rect 5053 7650 5067 7664
rect 5393 7693 5407 7707
rect 5213 7656 5227 7670
rect 5333 7650 5347 7664
rect 5413 7653 5427 7667
rect 5073 7613 5087 7627
rect 5053 7573 5067 7587
rect 5353 7573 5367 7587
rect 5013 7533 5027 7547
rect 4973 7093 4987 7107
rect 4972 7033 4986 7047
rect 4993 7033 5007 7047
rect 4973 6993 4987 7007
rect 4953 6913 4967 6927
rect 5053 7513 5067 7527
rect 5073 7473 5087 7487
rect 5313 7456 5327 7470
rect 5413 7473 5427 7487
rect 5393 7453 5407 7467
rect 5173 7313 5187 7327
rect 5073 7213 5087 7227
rect 5133 7213 5147 7227
rect 5053 7193 5067 7207
rect 5133 7173 5147 7187
rect 5033 7092 5047 7106
rect 5073 7093 5087 7107
rect 5013 6973 5027 6987
rect 4873 6890 4887 6904
rect 4833 6853 4847 6867
rect 4793 6793 4807 6807
rect 4833 6753 4847 6767
rect 4933 6893 4947 6907
rect 4913 6833 4927 6847
rect 4913 6733 4927 6747
rect 4873 6673 4887 6687
rect 4873 6636 4887 6650
rect 4593 6370 4607 6384
rect 4633 6370 4647 6384
rect 4673 6370 4687 6384
rect 4673 6333 4687 6347
rect 4713 6372 4727 6386
rect 4753 6373 4767 6387
rect 4693 6293 4707 6307
rect 4673 6116 4687 6130
rect 4453 5753 4467 5767
rect 4513 6070 4527 6084
rect 4573 6073 4587 6087
rect 4653 6033 4667 6047
rect 4573 5953 4587 5967
rect 4613 5913 4627 5927
rect 4473 5596 4487 5610
rect 4573 5833 4587 5847
rect 4513 5550 4527 5564
rect 4493 5453 4507 5467
rect 4473 5433 4487 5447
rect 4433 5393 4447 5407
rect 4473 5392 4487 5406
rect 4533 5413 4547 5427
rect 4493 5373 4507 5387
rect 4513 5353 4527 5367
rect 4453 5330 4467 5344
rect 4513 5293 4527 5307
rect 4553 5113 4567 5127
rect 4593 5793 4607 5807
rect 4593 5753 4607 5767
rect 4413 5093 4427 5107
rect 4533 5093 4547 5107
rect 4573 5093 4587 5107
rect 4433 5076 4447 5090
rect 4473 5053 4487 5067
rect 4353 4813 4367 4827
rect 4413 5030 4427 5044
rect 4453 5033 4467 5047
rect 4393 4873 4407 4887
rect 4533 5053 4547 5067
rect 4513 5013 4527 5027
rect 4493 4993 4507 5007
rect 4473 4953 4487 4967
rect 4493 4933 4507 4947
rect 4413 4813 4427 4827
rect 4433 4793 4447 4807
rect 4453 4773 4467 4787
rect 4373 4693 4387 4707
rect 4353 4673 4367 4687
rect 4353 4652 4367 4666
rect 4393 4653 4407 4667
rect 4433 4613 4447 4627
rect 4433 4556 4447 4570
rect 4413 4493 4427 4507
rect 4393 4473 4407 4487
rect 4373 4432 4387 4446
rect 4353 4373 4367 4387
rect 4433 4373 4447 4387
rect 4413 4336 4427 4350
rect 4353 4293 4367 4307
rect 4393 4290 4407 4304
rect 4453 3953 4467 3967
rect 4373 3913 4387 3927
rect 4413 3893 4427 3907
rect 4373 3816 4387 3830
rect 4333 3773 4347 3787
rect 4393 3770 4407 3784
rect 4433 3770 4447 3784
rect 4313 3693 4327 3707
rect 4373 3653 4387 3667
rect 4333 3516 4347 3530
rect 4573 4933 4587 4947
rect 4553 4913 4567 4927
rect 4553 4793 4567 4807
rect 4533 4773 4547 4787
rect 4513 4556 4527 4570
rect 4573 4513 4587 4527
rect 4553 4473 4567 4487
rect 4533 4433 4547 4447
rect 4533 4373 4547 4387
rect 4633 5633 4647 5647
rect 4613 5433 4627 5447
rect 4693 5953 4707 5967
rect 4693 5853 4707 5867
rect 4673 5713 4687 5727
rect 4733 6293 4747 6307
rect 4733 6173 4747 6187
rect 4733 6133 4747 6147
rect 4713 5833 4727 5847
rect 4693 5693 4707 5707
rect 4793 6116 4807 6130
rect 4953 6833 4967 6847
rect 5253 7253 5267 7267
rect 5173 7093 5187 7107
rect 5333 7353 5347 7367
rect 5293 7233 5307 7247
rect 5353 7193 5367 7207
rect 5393 7156 5407 7170
rect 5293 7093 5307 7107
rect 5113 7073 5127 7087
rect 5253 7073 5267 7087
rect 5373 7110 5387 7124
rect 5413 7113 5427 7127
rect 5353 7093 5367 7107
rect 5333 7053 5347 7067
rect 5093 6933 5107 6947
rect 5233 6910 5247 6924
rect 5433 7073 5447 7087
rect 5372 6993 5386 7007
rect 5393 6993 5407 7007
rect 5413 6973 5427 6987
rect 5393 6933 5407 6947
rect 5093 6873 5107 6887
rect 5393 6853 5407 6867
rect 5353 6813 5367 6827
rect 5073 6793 5087 6807
rect 5253 6793 5267 6807
rect 4953 6753 4967 6767
rect 5093 6733 5107 6747
rect 4953 6636 4967 6650
rect 5053 6636 5067 6650
rect 5093 6636 5107 6650
rect 5133 6636 5147 6650
rect 4953 6553 4967 6567
rect 4933 6513 4947 6527
rect 4993 6513 5007 6527
rect 4953 6473 4967 6487
rect 4933 6433 4947 6447
rect 4752 6073 4766 6087
rect 4773 6070 4787 6084
rect 4773 5993 4787 6007
rect 4853 6070 4867 6084
rect 4893 6093 4907 6107
rect 4893 6033 4907 6047
rect 4773 5833 4787 5847
rect 4753 5793 4767 5807
rect 4733 5633 4747 5647
rect 4853 5973 4867 5987
rect 4813 5953 4827 5967
rect 4853 5896 4867 5910
rect 4933 6133 4947 6147
rect 4973 6373 4987 6387
rect 4953 6073 4967 6087
rect 4913 5993 4927 6007
rect 4933 5973 4947 5987
rect 4853 5833 4867 5847
rect 4893 5833 4907 5847
rect 4773 5613 4787 5627
rect 4693 5596 4707 5610
rect 4733 5596 4747 5610
rect 4653 5553 4667 5567
rect 4873 5793 4887 5807
rect 5013 6433 5027 6447
rect 5053 6253 5067 6267
rect 5033 6233 5047 6247
rect 5273 6753 5287 6767
rect 5253 6473 5267 6487
rect 5193 6416 5207 6430
rect 5033 6193 5047 6207
rect 5133 6153 5147 6167
rect 5013 6133 5027 6147
rect 5013 6112 5027 6126
rect 5073 6116 5087 6130
rect 5033 6073 5047 6087
rect 5013 6013 5027 6027
rect 4753 5550 4767 5564
rect 4793 5550 4807 5564
rect 4832 5553 4846 5567
rect 4853 5553 4867 5567
rect 4693 5493 4707 5507
rect 4653 5453 4667 5467
rect 4653 5333 4667 5347
rect 4633 5293 4647 5307
rect 4693 5293 4707 5307
rect 4793 5253 4807 5267
rect 4873 5313 4887 5327
rect 4833 5233 4847 5247
rect 4913 5573 4927 5587
rect 4933 5513 4947 5527
rect 4913 5213 4927 5227
rect 4913 5113 4927 5127
rect 4613 5093 4627 5107
rect 4893 5093 4907 5107
rect 4613 5056 4627 5070
rect 4753 5056 4767 5070
rect 5013 5673 5027 5687
rect 5133 6073 5147 6087
rect 5213 6253 5227 6267
rect 5213 6232 5227 6246
rect 5213 6193 5227 6207
rect 5153 6013 5167 6027
rect 5092 5933 5106 5947
rect 5113 5933 5127 5947
rect 5073 5896 5087 5910
rect 5213 5993 5227 6007
rect 5073 5853 5087 5867
rect 5133 5833 5147 5847
rect 5173 5773 5187 5787
rect 5093 5753 5107 5767
rect 5093 5732 5107 5746
rect 5073 5693 5087 5707
rect 5033 5653 5047 5667
rect 4993 5596 5007 5610
rect 5013 5550 5027 5564
rect 4993 5493 5007 5507
rect 4973 5173 4987 5187
rect 4853 5053 4867 5067
rect 4613 5013 4627 5027
rect 4853 4953 4867 4967
rect 4693 4913 4707 4927
rect 4733 4873 4747 4887
rect 4833 4873 4847 4887
rect 4613 4653 4627 4667
rect 4613 4613 4627 4627
rect 4593 4473 4607 4487
rect 4653 4573 4667 4587
rect 4613 4413 4627 4427
rect 4773 4793 4787 4807
rect 4733 4753 4747 4767
rect 4713 4693 4727 4707
rect 4693 4513 4707 4527
rect 4613 4293 4627 4307
rect 4673 4290 4687 4304
rect 4593 4253 4607 4267
rect 4573 4233 4587 4247
rect 4573 4193 4587 4207
rect 4573 4153 4587 4167
rect 4553 4093 4567 4107
rect 4513 3990 4527 4004
rect 4573 3990 4587 4004
rect 4493 3853 4507 3867
rect 4493 3793 4507 3807
rect 4493 3693 4507 3707
rect 4473 3593 4487 3607
rect 4413 3553 4427 3567
rect 4473 3493 4487 3507
rect 4293 3373 4307 3387
rect 4393 3470 4407 3484
rect 4433 3473 4447 3487
rect 4393 3433 4407 3447
rect 4353 3413 4367 3427
rect 4413 3413 4427 3427
rect 4353 3373 4367 3387
rect 4313 3353 4327 3367
rect 4313 3296 4327 3310
rect 4413 3333 4427 3347
rect 4253 3253 4267 3267
rect 4233 2873 4247 2887
rect 4193 2793 4207 2807
rect 4213 2776 4227 2790
rect 4253 2776 4267 2790
rect 4193 2730 4207 2744
rect 4153 2713 4167 2727
rect 4253 2730 4267 2744
rect 4232 2693 4246 2707
rect 4253 2693 4267 2707
rect 4193 2673 4207 2687
rect 4173 2553 4187 2567
rect 4153 2413 4167 2427
rect 4153 2153 4167 2167
rect 4133 1393 4147 1407
rect 4113 1273 4127 1287
rect 4233 2633 4247 2647
rect 4333 3250 4347 3264
rect 4393 3250 4407 3264
rect 4293 3213 4307 3227
rect 4373 3213 4387 3227
rect 4313 3053 4327 3067
rect 4393 3053 4407 3067
rect 4353 2950 4367 2964
rect 4313 2893 4327 2907
rect 4293 2813 4307 2827
rect 4293 2553 4307 2567
rect 4273 2533 4287 2547
rect 4273 2476 4287 2490
rect 4353 2873 4367 2887
rect 4373 2813 4387 2827
rect 4333 2793 4347 2807
rect 4353 2772 4367 2786
rect 4333 2730 4347 2744
rect 4333 2673 4347 2687
rect 4253 2413 4267 2427
rect 4293 2393 4307 2407
rect 4293 2313 4307 2327
rect 4233 2256 4247 2270
rect 4253 2193 4267 2207
rect 4293 2193 4307 2207
rect 4213 2153 4227 2167
rect 4353 2133 4367 2147
rect 4213 2013 4227 2027
rect 4253 2013 4267 2027
rect 4293 2013 4307 2027
rect 4173 1956 4187 1970
rect 4253 1956 4267 1970
rect 4273 1910 4287 1924
rect 4253 1833 4267 1847
rect 4313 1773 4327 1787
rect 4293 1736 4307 1750
rect 4353 1736 4367 1750
rect 4313 1690 4327 1704
rect 4253 1533 4267 1547
rect 4213 1493 4227 1507
rect 4293 1493 4307 1507
rect 4153 1233 4167 1247
rect 4113 1217 4127 1231
rect 4113 1173 4127 1187
rect 4093 1053 4107 1067
rect 4253 1473 4267 1487
rect 4273 1390 4287 1404
rect 4273 1253 4287 1267
rect 4273 1216 4287 1230
rect 4313 1216 4327 1230
rect 4333 1170 4347 1184
rect 4293 1113 4307 1127
rect 4053 993 4067 1007
rect 4213 993 4227 1007
rect 3953 853 3967 867
rect 3873 833 3887 847
rect 3873 753 3887 767
rect 3813 693 3827 707
rect 3993 696 4007 710
rect 3793 673 3807 687
rect 3713 650 3727 664
rect 3753 650 3767 664
rect 3813 650 3827 664
rect 4253 973 4267 987
rect 4093 933 4107 947
rect 4173 933 4187 947
rect 4213 933 4227 947
rect 4193 870 4207 884
rect 4153 793 4167 807
rect 4273 933 4287 947
rect 4293 916 4307 930
rect 4273 873 4287 887
rect 4293 813 4307 827
rect 4313 733 4327 747
rect 4413 2793 4427 2807
rect 4473 3433 4487 3447
rect 4493 3213 4507 3227
rect 4453 3173 4467 3187
rect 4493 3153 4507 3167
rect 4533 3913 4547 3927
rect 4633 4233 4647 4247
rect 4713 4213 4727 4227
rect 4673 4193 4687 4207
rect 4633 4053 4647 4067
rect 4693 4133 4707 4147
rect 4673 3893 4687 3907
rect 4713 4093 4727 4107
rect 4773 4713 4787 4727
rect 4813 4493 4827 4507
rect 4793 4433 4807 4447
rect 4773 4393 4787 4407
rect 4773 4353 4787 4367
rect 4813 4313 4827 4327
rect 4793 4273 4807 4287
rect 4733 4033 4747 4047
rect 4773 4036 4787 4050
rect 4713 3993 4727 4007
rect 4793 3973 4807 3987
rect 4733 3953 4747 3967
rect 4813 3953 4827 3967
rect 4733 3893 4747 3907
rect 4773 3893 4787 3907
rect 4713 3853 4727 3867
rect 4753 3833 4767 3847
rect 4593 3770 4607 3784
rect 4653 3770 4667 3784
rect 4753 3770 4767 3784
rect 4793 3853 4807 3867
rect 4793 3733 4807 3747
rect 4553 3713 4567 3727
rect 4713 3713 4727 3727
rect 4533 3533 4547 3547
rect 4673 3673 4687 3687
rect 4593 3513 4607 3527
rect 4633 3516 4647 3530
rect 4773 3633 4787 3647
rect 4773 3593 4787 3607
rect 4713 3553 4727 3567
rect 4753 3533 4767 3547
rect 4553 3453 4567 3467
rect 4693 3453 4707 3467
rect 4733 3453 4747 3467
rect 4653 3413 4667 3427
rect 4593 3333 4607 3347
rect 4633 3333 4647 3347
rect 4533 3293 4547 3307
rect 4593 3296 4607 3310
rect 4713 3293 4727 3307
rect 4513 3093 4527 3107
rect 4453 2813 4467 2827
rect 4473 2793 4487 2807
rect 4433 2773 4447 2787
rect 4513 2776 4527 2790
rect 4613 3250 4627 3264
rect 4693 3253 4707 3267
rect 4673 3193 4687 3207
rect 4573 3153 4587 3167
rect 4633 3093 4647 3107
rect 4593 2996 4607 3010
rect 4613 2950 4627 2964
rect 4553 2933 4567 2947
rect 4653 2913 4667 2927
rect 4573 2753 4587 2767
rect 4453 2730 4467 2744
rect 4493 2713 4507 2727
rect 4513 2633 4527 2647
rect 4413 2593 4427 2607
rect 4553 2533 4567 2547
rect 4613 2593 4627 2607
rect 4573 2513 4587 2527
rect 4653 2512 4667 2526
rect 4613 2476 4627 2490
rect 4713 3153 4727 3167
rect 4753 3250 4767 3264
rect 4693 2773 4707 2787
rect 4793 3133 4807 3147
rect 4833 3693 4847 3707
rect 4833 3513 4847 3527
rect 4913 4813 4927 4827
rect 4913 4773 4927 4787
rect 4913 4713 4927 4727
rect 4893 4693 4907 4707
rect 4873 4433 4887 4447
rect 4913 4653 4927 4667
rect 5073 5550 5087 5564
rect 5053 5473 5067 5487
rect 5013 5453 5027 5467
rect 4993 4953 5007 4967
rect 5053 5433 5067 5447
rect 5073 5393 5087 5407
rect 5153 5613 5167 5627
rect 5133 5413 5147 5427
rect 5053 5313 5067 5327
rect 5033 5253 5047 5267
rect 5073 5073 5087 5087
rect 5173 5593 5187 5607
rect 5153 5213 5167 5227
rect 5193 5473 5207 5487
rect 5253 6293 5267 6307
rect 5253 6193 5267 6207
rect 5253 6113 5267 6127
rect 5253 6033 5267 6047
rect 5433 6733 5447 6747
rect 5352 6693 5366 6707
rect 5373 6693 5387 6707
rect 5293 6636 5307 6650
rect 5413 6636 5427 6650
rect 5313 6613 5327 6627
rect 5293 6313 5307 6327
rect 5293 6273 5307 6287
rect 5353 6593 5367 6607
rect 5333 6553 5347 6567
rect 5593 8093 5607 8107
rect 5533 8073 5547 8087
rect 5493 7913 5507 7927
rect 5473 7533 5487 7547
rect 5473 7453 5487 7467
rect 5473 7373 5487 7387
rect 5473 7352 5487 7366
rect 5573 8053 5587 8067
rect 5553 8033 5567 8047
rect 6093 9773 6107 9787
rect 6173 9933 6187 9947
rect 6253 10013 6267 10027
rect 6233 9793 6247 9807
rect 6213 9773 6227 9787
rect 6053 9613 6067 9627
rect 5973 9193 5987 9207
rect 6033 9193 6047 9207
rect 5973 9013 5987 9027
rect 5973 8913 5987 8927
rect 5953 8653 5967 8667
rect 5873 8613 5887 8627
rect 5953 8613 5967 8627
rect 5873 8592 5887 8606
rect 5913 8593 5927 8607
rect 5693 8573 5707 8587
rect 5813 8573 5827 8587
rect 5673 8353 5687 8367
rect 5793 8533 5807 8547
rect 5733 8513 5747 8527
rect 5693 8313 5707 8327
rect 5713 8293 5727 8307
rect 5673 8150 5687 8164
rect 5713 8150 5727 8164
rect 5593 8033 5607 8047
rect 5673 8033 5687 8047
rect 5593 7993 5607 8007
rect 5633 7976 5647 7990
rect 5573 7930 5587 7944
rect 5653 7930 5667 7944
rect 5693 7930 5707 7944
rect 5833 8496 5847 8510
rect 5753 8450 5767 8464
rect 5813 8450 5827 8464
rect 5773 8433 5787 8447
rect 5853 8433 5867 8447
rect 5933 8513 5947 8527
rect 5913 8433 5927 8447
rect 5953 8393 5967 8407
rect 5773 8313 5787 8327
rect 5773 8253 5787 8267
rect 5753 8053 5767 8067
rect 5753 7973 5767 7987
rect 5753 7930 5767 7944
rect 5733 7913 5747 7927
rect 5553 7893 5567 7907
rect 5553 7872 5567 7886
rect 5533 7853 5547 7867
rect 5593 7853 5607 7867
rect 5553 7813 5567 7827
rect 5753 7813 5767 7827
rect 5533 7733 5547 7747
rect 5713 7733 5727 7747
rect 5553 7693 5567 7707
rect 5613 7676 5627 7690
rect 5553 7630 5567 7644
rect 5593 7630 5607 7644
rect 5533 7613 5547 7627
rect 5613 7613 5627 7627
rect 5673 7630 5687 7644
rect 5593 7593 5607 7607
rect 5593 7553 5607 7567
rect 5633 7573 5647 7587
rect 5673 7573 5687 7587
rect 5653 7553 5667 7567
rect 5733 7676 5747 7690
rect 5573 7533 5587 7547
rect 5613 7533 5627 7547
rect 5713 7553 5727 7567
rect 5693 7533 5707 7547
rect 5673 7513 5687 7527
rect 5653 7453 5667 7467
rect 5713 7473 5727 7487
rect 5733 7433 5747 7447
rect 5513 7333 5527 7347
rect 5513 7173 5527 7187
rect 5513 7152 5527 7166
rect 5493 7072 5507 7086
rect 5473 7052 5487 7066
rect 5473 6813 5487 6827
rect 5493 6773 5507 6787
rect 5473 6753 5487 6767
rect 5393 6553 5407 6567
rect 5453 6553 5467 6567
rect 5373 6493 5387 6507
rect 5373 6373 5387 6387
rect 5353 6333 5367 6347
rect 5353 6153 5367 6167
rect 5333 6070 5347 6084
rect 5553 7410 5567 7424
rect 5593 7393 5607 7407
rect 5673 7393 5687 7407
rect 5733 7393 5747 7407
rect 5633 7353 5647 7367
rect 5553 7253 5567 7267
rect 5533 7113 5547 7127
rect 5533 6773 5547 6787
rect 5533 6613 5547 6627
rect 5513 6593 5527 6607
rect 5533 6553 5547 6567
rect 5493 6513 5507 6527
rect 5453 6493 5467 6507
rect 5453 6433 5467 6447
rect 5493 6416 5507 6430
rect 5613 7213 5627 7227
rect 5713 7373 5727 7387
rect 5733 7353 5747 7367
rect 5733 7332 5747 7346
rect 5733 7293 5747 7307
rect 5793 8233 5807 8247
rect 5773 7773 5787 7787
rect 5773 7733 5787 7747
rect 5833 8150 5847 8164
rect 5853 7993 5867 8007
rect 5853 7693 5867 7707
rect 5833 7673 5847 7687
rect 5933 8213 5947 8227
rect 6073 9573 6087 9587
rect 6333 10153 6347 10167
rect 6673 10253 6687 10267
rect 6393 10056 6407 10070
rect 6533 10053 6547 10067
rect 6413 10010 6427 10024
rect 6513 10010 6527 10024
rect 6473 9993 6487 10007
rect 6333 9813 6347 9827
rect 6153 9613 6167 9627
rect 6293 9613 6307 9627
rect 6213 9573 6227 9587
rect 6113 9533 6127 9547
rect 6173 9536 6187 9550
rect 6253 9536 6267 9550
rect 6313 9536 6327 9550
rect 6193 9433 6207 9447
rect 6233 9433 6247 9447
rect 6113 9253 6127 9267
rect 6153 9236 6167 9250
rect 6213 9236 6227 9250
rect 6133 9190 6147 9204
rect 6173 9190 6187 9204
rect 6073 9153 6087 9167
rect 6133 9153 6147 9167
rect 6053 8813 6067 8827
rect 6033 8753 6047 8767
rect 6113 8753 6127 8767
rect 6013 8733 6027 8747
rect 5993 8713 6007 8727
rect 6073 8716 6087 8730
rect 5993 8673 6007 8687
rect 6013 8653 6027 8667
rect 5993 8353 6007 8367
rect 5953 8150 5967 8164
rect 5993 8013 6007 8027
rect 5913 7993 5927 8007
rect 5933 7976 5947 7990
rect 5953 7930 5967 7944
rect 5993 7930 6007 7944
rect 5913 7853 5927 7867
rect 6033 8593 6047 8607
rect 6013 7813 6027 7827
rect 5913 7693 5927 7707
rect 5953 7676 5967 7690
rect 6013 7673 6027 7687
rect 5793 7553 5807 7567
rect 5773 7533 5787 7547
rect 5933 7533 5947 7547
rect 6013 7473 6027 7487
rect 5773 7433 5787 7447
rect 6053 8493 6067 8507
rect 6173 9073 6187 9087
rect 6153 8933 6167 8947
rect 6133 8593 6147 8607
rect 6313 9273 6327 9287
rect 6253 9253 6267 9267
rect 6233 9053 6247 9067
rect 6313 9236 6327 9250
rect 6313 9193 6327 9207
rect 6313 9113 6327 9127
rect 6273 8953 6287 8967
rect 6193 8893 6207 8907
rect 6233 8893 6247 8907
rect 6193 8733 6207 8747
rect 6173 8652 6187 8666
rect 6153 8533 6167 8547
rect 6153 8496 6167 8510
rect 6053 8453 6067 8467
rect 6093 8450 6107 8464
rect 6133 8450 6147 8464
rect 6053 8432 6067 8446
rect 6053 8393 6067 8407
rect 6133 8313 6147 8327
rect 6173 8313 6187 8327
rect 6133 8273 6147 8287
rect 6113 8093 6127 8107
rect 6093 8053 6107 8067
rect 6033 7453 6047 7467
rect 5913 7430 5927 7444
rect 6013 7430 6027 7444
rect 6113 7930 6127 7944
rect 6113 7813 6127 7827
rect 6093 7493 6107 7507
rect 5773 7393 5787 7407
rect 6073 7390 6087 7404
rect 6073 7333 6087 7347
rect 6013 7313 6027 7327
rect 5993 7253 6007 7267
rect 5753 7233 5767 7247
rect 5773 7193 5787 7207
rect 5813 7193 5827 7207
rect 5753 7173 5767 7187
rect 5573 6913 5587 6927
rect 5633 6890 5647 6904
rect 5713 7110 5727 7124
rect 5733 7093 5747 7107
rect 5713 6973 5727 6987
rect 5613 6853 5627 6867
rect 5673 6853 5687 6867
rect 5713 6853 5727 6867
rect 5573 6833 5587 6847
rect 5573 6793 5587 6807
rect 5593 6693 5607 6707
rect 5573 6513 5587 6527
rect 5673 6693 5687 6707
rect 5613 6633 5627 6647
rect 5813 7156 5827 7170
rect 5873 7156 5887 7170
rect 5913 7156 5927 7170
rect 5953 7156 5967 7170
rect 5793 7053 5807 7067
rect 5853 7110 5867 7124
rect 5813 7033 5827 7047
rect 5932 7053 5946 7067
rect 5953 7053 5967 7067
rect 5973 7033 5987 7047
rect 5893 7013 5907 7027
rect 5933 7013 5947 7027
rect 5893 6992 5907 7006
rect 5933 6973 5947 6987
rect 5833 6913 5847 6927
rect 5793 6893 5807 6907
rect 5773 6753 5787 6767
rect 5753 6693 5767 6707
rect 5733 6673 5747 6687
rect 5633 6573 5647 6587
rect 5613 6493 5627 6507
rect 5593 6433 5607 6447
rect 5613 6413 5627 6427
rect 5553 6393 5567 6407
rect 5593 6396 5607 6410
rect 5413 6373 5427 6387
rect 5333 6033 5347 6047
rect 5393 6033 5407 6047
rect 5313 5993 5327 6007
rect 5273 5853 5287 5867
rect 5293 5633 5307 5647
rect 5413 5993 5427 6007
rect 5473 6370 5487 6384
rect 5493 6353 5507 6367
rect 5552 6353 5566 6367
rect 5573 6353 5587 6367
rect 5613 6353 5627 6367
rect 5473 6333 5487 6347
rect 5453 6113 5467 6127
rect 5453 6053 5467 6067
rect 5433 5973 5447 5987
rect 5393 5896 5407 5910
rect 5353 5853 5367 5867
rect 5333 5733 5347 5747
rect 5313 5596 5327 5610
rect 5393 5813 5407 5827
rect 5373 5773 5387 5787
rect 5373 5693 5387 5707
rect 5373 5613 5387 5627
rect 5353 5593 5367 5607
rect 5273 5473 5287 5487
rect 5233 5453 5247 5467
rect 5213 5413 5227 5427
rect 5213 5353 5227 5367
rect 5193 5133 5207 5147
rect 5113 5093 5127 5107
rect 5173 5093 5187 5107
rect 5053 5033 5067 5047
rect 5033 4973 5047 4987
rect 5073 4913 5087 4927
rect 5013 4873 5027 4887
rect 5193 5076 5207 5090
rect 5113 4873 5127 4887
rect 4973 4852 4987 4866
rect 5033 4856 5047 4870
rect 5073 4856 5087 4870
rect 5113 4852 5127 4866
rect 5013 4810 5027 4824
rect 5093 4773 5107 4787
rect 5053 4713 5067 4727
rect 4973 4556 4987 4570
rect 5013 4556 5027 4570
rect 5073 4556 5087 4570
rect 4933 4452 4947 4466
rect 4933 4373 4947 4387
rect 4913 4290 4927 4304
rect 4893 4273 4907 4287
rect 4873 4056 4887 4070
rect 4953 4193 4967 4207
rect 4933 4073 4947 4087
rect 4893 3913 4907 3927
rect 5033 4493 5047 4507
rect 5153 5030 5167 5044
rect 5173 4973 5187 4987
rect 5153 4873 5167 4887
rect 5153 4833 5167 4847
rect 5173 4753 5187 4767
rect 5153 4673 5167 4687
rect 5313 5433 5327 5447
rect 5253 5373 5267 5387
rect 5473 5813 5487 5827
rect 5413 5773 5427 5787
rect 5433 5653 5447 5667
rect 5333 5330 5347 5344
rect 5433 5333 5447 5347
rect 5273 5233 5287 5247
rect 5233 5013 5247 5027
rect 5313 5153 5327 5167
rect 5293 5133 5307 5147
rect 5233 4893 5247 4907
rect 5273 4893 5287 4907
rect 5213 4493 5227 4507
rect 5133 4473 5147 4487
rect 5113 4373 5127 4387
rect 5153 4336 5167 4350
rect 5313 5076 5327 5090
rect 5513 6293 5527 6307
rect 5513 6073 5527 6087
rect 5493 5773 5507 5787
rect 5473 5753 5487 5767
rect 5553 6313 5567 6327
rect 5613 6313 5627 6327
rect 5593 6273 5607 6287
rect 5573 6113 5587 6127
rect 5693 6590 5707 6604
rect 5733 6590 5747 6604
rect 5873 6890 5887 6904
rect 5913 6890 5927 6904
rect 5973 6890 5987 6904
rect 5933 6873 5947 6887
rect 5873 6833 5887 6847
rect 5833 6573 5847 6587
rect 6013 7093 6027 7107
rect 6033 6913 6047 6927
rect 6073 6893 6087 6907
rect 6073 6853 6087 6867
rect 6053 6833 6067 6847
rect 5993 6793 6007 6807
rect 6073 6753 6087 6767
rect 6013 6733 6027 6747
rect 5913 6636 5927 6650
rect 5993 6573 6007 6587
rect 5933 6553 5947 6567
rect 5873 6533 5887 6547
rect 5653 6493 5667 6507
rect 5973 6473 5987 6487
rect 5653 6433 5667 6447
rect 5973 6433 5987 6447
rect 5793 6390 5807 6404
rect 5913 6396 5927 6410
rect 5993 6392 6007 6406
rect 5653 6353 5667 6367
rect 5953 6350 5967 6364
rect 5953 6313 5967 6327
rect 6033 6653 6047 6667
rect 6053 6633 6067 6647
rect 6053 6593 6067 6607
rect 6033 6473 6047 6487
rect 6013 6313 6027 6327
rect 5953 6253 5967 6267
rect 5792 6233 5806 6247
rect 5813 6233 5827 6247
rect 5633 6173 5647 6187
rect 5693 6173 5707 6187
rect 5753 6173 5767 6187
rect 5633 6116 5647 6130
rect 5653 6070 5667 6084
rect 5733 6153 5747 6167
rect 5653 6033 5667 6047
rect 5693 6033 5707 6047
rect 5633 5993 5647 6007
rect 5613 5813 5627 5827
rect 5553 5753 5567 5767
rect 5553 5673 5567 5687
rect 5593 5673 5607 5687
rect 5473 5633 5487 5647
rect 5533 5633 5547 5647
rect 5453 5293 5467 5307
rect 5533 5596 5547 5610
rect 5593 5613 5607 5627
rect 5473 5233 5487 5247
rect 5413 5213 5427 5227
rect 5373 5193 5387 5207
rect 5453 5076 5467 5090
rect 5493 5076 5507 5090
rect 5353 4973 5367 4987
rect 5313 4933 5327 4947
rect 5333 4856 5347 4870
rect 5433 5013 5447 5027
rect 5453 4933 5467 4947
rect 5493 4933 5507 4947
rect 5393 4853 5407 4867
rect 5373 4813 5387 4827
rect 5313 4793 5327 4807
rect 5313 4573 5327 4587
rect 5353 4556 5367 4570
rect 5293 4473 5307 4487
rect 5253 4336 5267 4350
rect 5053 4293 5067 4307
rect 5173 4290 5187 4304
rect 5213 4290 5227 4304
rect 5033 4233 5047 4247
rect 5133 4233 5147 4247
rect 5253 4153 5267 4167
rect 5073 4133 5087 4147
rect 5053 4073 5067 4087
rect 4973 4033 4987 4047
rect 5013 4036 5027 4050
rect 5313 4453 5327 4467
rect 5313 4373 5327 4387
rect 5293 4193 5307 4207
rect 5373 4290 5387 4304
rect 5433 4853 5447 4867
rect 5433 4793 5447 4807
rect 5413 4533 5427 4547
rect 5413 4493 5427 4507
rect 5493 4873 5507 4887
rect 5453 4413 5467 4427
rect 5493 4773 5507 4787
rect 5493 4673 5507 4687
rect 5533 5533 5547 5547
rect 5533 5473 5547 5487
rect 5553 5373 5567 5387
rect 5593 5573 5607 5587
rect 5613 5473 5627 5487
rect 5673 5973 5687 5987
rect 5713 5953 5727 5967
rect 5693 5933 5707 5947
rect 5793 6153 5807 6167
rect 5753 6116 5767 6130
rect 5793 6033 5807 6047
rect 5753 5973 5767 5987
rect 5713 5913 5727 5927
rect 5713 5850 5727 5864
rect 5713 5793 5727 5807
rect 5693 5613 5707 5627
rect 5693 5373 5707 5387
rect 5593 5330 5607 5344
rect 5673 5330 5687 5344
rect 5633 5293 5647 5307
rect 5673 5233 5687 5247
rect 5653 5213 5667 5227
rect 5633 5013 5647 5027
rect 5613 4953 5627 4967
rect 5573 4893 5587 4907
rect 5553 4873 5567 4887
rect 5573 4856 5587 4870
rect 5553 4810 5567 4824
rect 5593 4773 5607 4787
rect 5593 4752 5607 4766
rect 5553 4673 5567 4687
rect 5613 4653 5627 4667
rect 5533 4613 5547 4627
rect 5513 4593 5527 4607
rect 5513 4453 5527 4467
rect 5493 4393 5507 4407
rect 5493 4372 5507 4386
rect 5453 4353 5467 4367
rect 5513 4333 5527 4347
rect 5653 4810 5667 4824
rect 5653 4733 5667 4747
rect 5573 4510 5587 4524
rect 5653 4513 5667 4527
rect 5653 4492 5667 4506
rect 5573 4393 5587 4407
rect 5553 4373 5567 4387
rect 5433 4290 5447 4304
rect 5533 4293 5547 4307
rect 5513 4253 5527 4267
rect 5393 4173 5407 4187
rect 5313 4133 5327 4147
rect 5433 4133 5447 4147
rect 5273 4113 5287 4127
rect 5113 4056 5127 4070
rect 5073 4033 5087 4047
rect 5133 4013 5147 4027
rect 4973 3993 4987 4007
rect 4953 3953 4967 3967
rect 4993 3953 5007 3967
rect 4952 3893 4966 3907
rect 4973 3893 4987 3907
rect 4933 3873 4947 3887
rect 4873 3733 4887 3747
rect 4973 3753 4987 3767
rect 4933 3633 4947 3647
rect 4893 3553 4907 3567
rect 4953 3516 4967 3530
rect 4933 3470 4947 3484
rect 5113 3953 5127 3967
rect 5053 3933 5067 3947
rect 5033 3913 5047 3927
rect 5093 3893 5107 3907
rect 5073 3613 5087 3627
rect 5033 3553 5047 3567
rect 5013 3433 5027 3447
rect 4853 3393 4867 3407
rect 4933 3353 4947 3367
rect 4833 3333 4847 3347
rect 4973 3333 4987 3347
rect 4953 3313 4967 3327
rect 4873 3296 4887 3310
rect 4913 3296 4927 3310
rect 4893 3233 4907 3247
rect 4853 3213 4867 3227
rect 4953 3193 4967 3207
rect 4953 3153 4967 3167
rect 4893 3133 4907 3147
rect 4893 3093 4907 3107
rect 4893 2996 4907 3010
rect 4813 2932 4827 2946
rect 4753 2793 4767 2807
rect 4733 2730 4747 2744
rect 4773 2730 4787 2744
rect 4693 2713 4707 2727
rect 4673 2476 4687 2490
rect 4513 2430 4527 2444
rect 4473 2393 4487 2407
rect 4473 2293 4487 2307
rect 4513 2256 4527 2270
rect 4593 2430 4607 2444
rect 4653 2433 4667 2447
rect 4653 2333 4667 2347
rect 4633 2273 4647 2287
rect 4393 2133 4407 2147
rect 4393 2093 4407 2107
rect 4393 1933 4407 1947
rect 4533 2210 4547 2224
rect 4573 2210 4587 2224
rect 4613 2193 4627 2207
rect 4553 2133 4567 2147
rect 4533 2093 4547 2107
rect 4493 2073 4507 2087
rect 4453 2053 4467 2067
rect 4553 2033 4567 2047
rect 4533 2013 4547 2027
rect 4453 1973 4467 1987
rect 4633 2093 4647 2107
rect 4613 1993 4627 2007
rect 4513 1893 4527 1907
rect 4493 1873 4507 1887
rect 4493 1833 4507 1847
rect 4553 1833 4567 1847
rect 4413 1813 4427 1827
rect 4473 1813 4487 1827
rect 4413 1773 4427 1787
rect 4633 1893 4647 1907
rect 4553 1773 4567 1787
rect 4613 1773 4627 1787
rect 4413 1513 4427 1527
rect 4393 1170 4407 1184
rect 4433 1413 4447 1427
rect 4413 1153 4427 1167
rect 4593 1736 4607 1750
rect 4513 1693 4527 1707
rect 4473 1473 4487 1487
rect 4573 1633 4587 1647
rect 4533 1573 4547 1587
rect 4513 1453 4527 1467
rect 4573 1436 4587 1450
rect 4613 1436 4627 1450
rect 4513 1390 4527 1404
rect 4753 2673 4767 2687
rect 4713 2473 4727 2487
rect 4693 2193 4707 2207
rect 4673 2153 4687 2167
rect 4693 2133 4707 2147
rect 4673 2073 4687 2087
rect 4653 1732 4667 1746
rect 4653 1613 4667 1627
rect 4673 1573 4687 1587
rect 4633 1393 4647 1407
rect 4553 1353 4567 1367
rect 4733 2333 4747 2347
rect 4773 2573 4787 2587
rect 4753 2293 4767 2307
rect 4913 2933 4927 2947
rect 4873 2873 4887 2887
rect 4933 2873 4947 2887
rect 4853 2853 4867 2867
rect 4913 2833 4927 2847
rect 4853 2730 4867 2744
rect 4873 2693 4887 2707
rect 4833 2673 4847 2687
rect 4813 2473 4827 2487
rect 4913 2653 4927 2667
rect 4933 2633 4947 2647
rect 4933 2593 4947 2607
rect 4893 2473 4907 2487
rect 4793 2453 4807 2467
rect 4773 2273 4787 2287
rect 4753 2053 4767 2067
rect 4733 1973 4747 1987
rect 4633 1333 4647 1347
rect 4693 1333 4707 1347
rect 4693 1293 4707 1307
rect 4553 1216 4567 1230
rect 4633 1216 4647 1230
rect 4693 1196 4707 1210
rect 4893 2433 4907 2447
rect 4873 2393 4887 2407
rect 4793 2133 4807 2147
rect 4853 2133 4867 2147
rect 4773 1973 4787 1987
rect 4913 2313 4927 2327
rect 4893 2013 4907 2027
rect 4833 1956 4847 1970
rect 4753 1933 4767 1947
rect 4813 1873 4827 1887
rect 4833 1753 4847 1767
rect 4893 1873 4907 1887
rect 4753 1736 4767 1750
rect 4793 1736 4807 1750
rect 4873 1733 4887 1747
rect 4853 1690 4867 1704
rect 4813 1653 4827 1667
rect 4813 1573 4827 1587
rect 4753 1553 4767 1567
rect 4753 1513 4767 1527
rect 4793 1473 4807 1487
rect 4893 1473 4907 1487
rect 4753 1453 4767 1467
rect 4833 1436 4847 1450
rect 4813 1390 4827 1404
rect 4753 1333 4767 1347
rect 4893 1390 4907 1404
rect 4873 1313 4887 1327
rect 4933 1956 4947 1970
rect 4933 1613 4947 1627
rect 4933 1353 4947 1367
rect 4973 2996 4987 3010
rect 5093 3473 5107 3487
rect 5133 3633 5147 3647
rect 5273 4016 5287 4030
rect 5453 4113 5467 4127
rect 5513 4113 5527 4127
rect 5453 4053 5467 4067
rect 5633 4253 5647 4267
rect 5613 4173 5627 4187
rect 5453 4013 5467 4027
rect 5433 3993 5447 4007
rect 5253 3913 5267 3927
rect 5353 3913 5367 3927
rect 5353 3873 5367 3887
rect 5393 3873 5407 3887
rect 5273 3853 5287 3867
rect 5373 3852 5387 3866
rect 5333 3753 5347 3767
rect 5293 3653 5307 3667
rect 5233 3633 5247 3647
rect 5193 3593 5207 3607
rect 5233 3533 5247 3547
rect 5193 3516 5207 3530
rect 5313 3593 5327 3607
rect 5213 3470 5227 3484
rect 5293 3470 5307 3484
rect 5253 3433 5267 3447
rect 5113 3373 5127 3387
rect 5173 3296 5187 3310
rect 5093 3233 5107 3247
rect 4993 2873 5007 2887
rect 4973 2792 4987 2806
rect 5033 3073 5047 3087
rect 5073 3213 5087 3227
rect 5073 3192 5087 3206
rect 5073 3133 5087 3147
rect 5073 3073 5087 3087
rect 5053 2913 5067 2927
rect 5033 2813 5047 2827
rect 5033 2776 5047 2790
rect 5193 3233 5207 3247
rect 5133 3213 5147 3227
rect 5213 3133 5227 3147
rect 5153 3113 5167 3127
rect 5193 3093 5207 3107
rect 5153 3033 5167 3047
rect 5133 2996 5147 3010
rect 5013 2730 5027 2744
rect 5053 2730 5067 2744
rect 5113 2730 5127 2744
rect 4993 2613 5007 2627
rect 5173 2773 5187 2787
rect 5153 2573 5167 2587
rect 5073 2553 5087 2567
rect 5033 2476 5047 2490
rect 5213 3053 5227 3067
rect 5213 2973 5227 2987
rect 5213 2913 5227 2927
rect 5213 2793 5227 2807
rect 5213 2613 5227 2627
rect 5213 2573 5227 2587
rect 5193 2553 5207 2567
rect 5293 3373 5307 3387
rect 5273 3296 5287 3310
rect 5273 3073 5287 3087
rect 5373 3733 5387 3747
rect 5353 3633 5367 3647
rect 5533 3993 5547 4007
rect 5453 3953 5467 3967
rect 5513 3893 5527 3907
rect 5593 3953 5607 3967
rect 5573 3833 5587 3847
rect 5453 3770 5467 3784
rect 5433 3753 5447 3767
rect 5532 3770 5546 3784
rect 5553 3770 5567 3784
rect 5493 3733 5507 3747
rect 5433 3673 5447 3687
rect 5413 3653 5427 3667
rect 5453 3573 5467 3587
rect 5433 3533 5447 3547
rect 5553 3613 5567 3627
rect 5553 3573 5567 3587
rect 5453 3470 5467 3484
rect 5413 3333 5427 3347
rect 5553 3453 5567 3467
rect 5473 3393 5487 3407
rect 5393 3313 5407 3327
rect 5373 3292 5387 3306
rect 5433 3296 5447 3310
rect 5353 3253 5367 3267
rect 5413 3250 5427 3264
rect 5493 3296 5507 3310
rect 5473 3213 5487 3227
rect 5453 3193 5467 3207
rect 5493 3133 5507 3147
rect 5333 3033 5347 3047
rect 5373 2996 5387 3010
rect 5333 2950 5347 2964
rect 5413 2950 5427 2964
rect 5313 2933 5327 2947
rect 5433 2933 5447 2947
rect 5293 2793 5307 2807
rect 5313 2776 5327 2790
rect 5433 2773 5447 2787
rect 5473 2776 5487 2790
rect 5333 2730 5347 2744
rect 5453 2730 5467 2744
rect 5293 2713 5307 2727
rect 5493 2733 5507 2747
rect 5533 2933 5547 2947
rect 5653 3993 5667 4007
rect 5633 3933 5647 3947
rect 5653 3813 5667 3827
rect 5693 5193 5707 5207
rect 5733 5733 5747 5747
rect 5773 5693 5787 5707
rect 5893 6173 5907 6187
rect 5833 6133 5847 6147
rect 5993 6093 6007 6107
rect 5853 6070 5867 6084
rect 5873 6053 5887 6067
rect 5873 5973 5887 5987
rect 5913 5973 5927 5987
rect 5853 5933 5867 5947
rect 5873 5913 5887 5927
rect 5893 5896 5907 5910
rect 5893 5813 5907 5827
rect 5833 5793 5847 5807
rect 5813 5733 5827 5747
rect 5893 5653 5907 5667
rect 5793 5613 5807 5627
rect 5813 5596 5827 5610
rect 5873 5596 5887 5610
rect 5733 5533 5747 5547
rect 5833 5550 5847 5564
rect 5793 5393 5807 5407
rect 6033 6033 6047 6047
rect 6253 8673 6267 8687
rect 6233 8653 6247 8667
rect 6233 8573 6247 8587
rect 6253 8450 6267 8464
rect 6233 8433 6247 8447
rect 6213 8393 6227 8407
rect 6193 8213 6207 8227
rect 6213 8196 6227 8210
rect 6193 8150 6207 8164
rect 6153 8133 6167 8147
rect 6233 8133 6247 8147
rect 6213 7976 6227 7990
rect 6193 7930 6207 7944
rect 6233 7913 6247 7927
rect 6233 7833 6247 7847
rect 6193 7773 6207 7787
rect 6193 7676 6207 7690
rect 6213 7633 6227 7647
rect 6173 7593 6187 7607
rect 6153 7573 6167 7587
rect 6153 7533 6167 7547
rect 6173 7493 6187 7507
rect 6153 7373 6167 7387
rect 6313 8933 6327 8947
rect 6313 8873 6327 8887
rect 6313 8773 6327 8787
rect 6413 9756 6427 9770
rect 6393 9673 6407 9687
rect 6513 9673 6527 9687
rect 6473 9613 6487 9627
rect 6373 9490 6387 9504
rect 6433 9490 6447 9504
rect 6353 9413 6367 9427
rect 6393 9273 6407 9287
rect 6433 9236 6447 9250
rect 6473 9490 6487 9504
rect 6613 10053 6627 10067
rect 6753 10113 6767 10127
rect 6653 10010 6667 10024
rect 6693 9973 6707 9987
rect 6573 9853 6587 9867
rect 6533 9573 6547 9587
rect 6513 9473 6527 9487
rect 6533 9453 6547 9467
rect 6513 9433 6527 9447
rect 6533 9236 6547 9250
rect 6633 9756 6647 9770
rect 6713 9753 6727 9767
rect 6713 9653 6727 9667
rect 6773 10013 6787 10027
rect 6833 10313 6847 10327
rect 6893 10230 6907 10244
rect 6913 10113 6927 10127
rect 6953 10433 6967 10447
rect 6953 10373 6967 10387
rect 6933 10093 6947 10107
rect 6953 10056 6967 10070
rect 7693 12093 7707 12107
rect 7533 11873 7547 11887
rect 7733 11873 7747 11887
rect 7633 11836 7647 11850
rect 7673 11836 7687 11850
rect 7613 11733 7627 11747
rect 7713 11773 7727 11787
rect 7613 11693 7627 11707
rect 7673 11693 7687 11707
rect 7573 11653 7587 11667
rect 7573 11616 7587 11630
rect 7653 11616 7667 11630
rect 7633 11553 7647 11567
rect 7993 12133 8007 12147
rect 8053 12116 8067 12130
rect 8253 12110 8267 12124
rect 8352 12110 8366 12124
rect 8373 12116 8387 12130
rect 8453 12113 8467 12127
rect 7773 12093 7787 12107
rect 7573 11473 7587 11487
rect 7673 11473 7687 11487
rect 7753 11473 7767 11487
rect 7133 11413 7147 11427
rect 7513 11413 7527 11427
rect 7633 11413 7647 11427
rect 7073 11373 7087 11387
rect 7633 11336 7647 11350
rect 7133 11316 7147 11330
rect 7173 11270 7187 11284
rect 7173 11193 7187 11207
rect 7213 11173 7227 11187
rect 7473 11296 7487 11310
rect 7572 11296 7586 11310
rect 7593 11290 7607 11304
rect 7573 11253 7587 11267
rect 7613 11253 7627 11267
rect 7333 11173 7347 11187
rect 7273 11133 7287 11147
rect 7093 11096 7107 11110
rect 7533 11096 7547 11110
rect 7573 11096 7587 11110
rect 7353 11050 7367 11064
rect 7533 11053 7547 11067
rect 7653 11053 7667 11067
rect 7653 11013 7667 11027
rect 7113 10913 7127 10927
rect 7033 10853 7047 10867
rect 7013 10533 7027 10547
rect 7013 10230 7027 10244
rect 7113 10813 7127 10827
rect 7593 10933 7607 10947
rect 7493 10833 7507 10847
rect 7173 10816 7187 10830
rect 7093 10796 7107 10810
rect 7133 10796 7147 10810
rect 7113 10750 7127 10764
rect 7153 10753 7167 10767
rect 7073 10733 7087 10747
rect 7053 10713 7067 10727
rect 7053 10576 7067 10590
rect 7053 10533 7067 10547
rect 7133 10693 7147 10707
rect 7093 10573 7107 10587
rect 7073 10433 7087 10447
rect 7333 10776 7347 10790
rect 7493 10753 7507 10767
rect 7213 10693 7227 10707
rect 7253 10653 7267 10667
rect 7153 10573 7167 10587
rect 7193 10576 7207 10590
rect 7533 10733 7547 10747
rect 7593 10693 7607 10707
rect 7553 10673 7567 10687
rect 7513 10653 7527 10667
rect 7493 10633 7507 10647
rect 7273 10573 7287 10587
rect 7393 10576 7407 10590
rect 7433 10576 7447 10590
rect 7473 10576 7487 10590
rect 7213 10530 7227 10544
rect 7193 10453 7207 10467
rect 7073 10273 7087 10287
rect 7133 10276 7147 10290
rect 7053 10193 7067 10207
rect 7033 10093 7047 10107
rect 7013 10053 7027 10067
rect 6933 10010 6947 10024
rect 7033 10012 7047 10026
rect 7012 9973 7026 9987
rect 7033 9973 7047 9987
rect 6833 9813 6847 9827
rect 6973 9793 6987 9807
rect 6913 9756 6927 9770
rect 6893 9653 6907 9667
rect 6813 9633 6827 9647
rect 6873 9633 6887 9647
rect 6613 9613 6627 9627
rect 6753 9613 6767 9627
rect 6593 9536 6607 9550
rect 6593 9413 6607 9427
rect 6593 9373 6607 9387
rect 6653 9536 6667 9550
rect 6693 9536 6707 9550
rect 6673 9473 6687 9487
rect 6693 9453 6707 9467
rect 6613 9333 6627 9347
rect 6593 9236 6607 9250
rect 6413 9190 6427 9204
rect 6573 9193 6587 9207
rect 6653 9190 6667 9204
rect 6533 9173 6547 9187
rect 6593 9173 6607 9187
rect 6453 9133 6467 9147
rect 6373 9093 6387 9107
rect 6413 9093 6427 9107
rect 6353 8953 6367 8967
rect 6413 9053 6427 9067
rect 6453 9033 6467 9047
rect 6453 9012 6467 9026
rect 6493 9016 6507 9030
rect 6633 9113 6647 9127
rect 6613 9053 6627 9067
rect 6413 8970 6427 8984
rect 6373 8833 6387 8847
rect 6413 8773 6427 8787
rect 6333 8733 6347 8747
rect 6353 8716 6367 8730
rect 6513 8970 6527 8984
rect 6553 8970 6567 8984
rect 6613 8970 6627 8984
rect 6533 8933 6547 8947
rect 6513 8853 6527 8867
rect 6473 8833 6487 8847
rect 6473 8716 6487 8730
rect 6432 8673 6446 8687
rect 6453 8673 6467 8687
rect 6373 8633 6387 8647
rect 6333 8613 6347 8627
rect 6373 8533 6387 8547
rect 6333 8493 6347 8507
rect 6393 8496 6407 8510
rect 6313 8333 6327 8347
rect 6293 8273 6307 8287
rect 6373 8450 6387 8464
rect 6453 8453 6467 8467
rect 6353 8433 6367 8447
rect 6473 8433 6487 8447
rect 6333 8293 6347 8307
rect 6313 8153 6327 8167
rect 6293 8133 6307 8147
rect 6373 8353 6387 8367
rect 6353 8053 6367 8067
rect 6293 7893 6307 7907
rect 6273 7633 6287 7647
rect 6353 7513 6367 7527
rect 6253 7453 6267 7467
rect 6293 7456 6307 7470
rect 6233 7353 6247 7367
rect 6133 7333 6147 7347
rect 6173 7333 6187 7347
rect 6193 7233 6207 7247
rect 6153 7213 6167 7227
rect 6193 7156 6207 7170
rect 6173 7110 6187 7124
rect 6113 7073 6127 7087
rect 6213 7073 6227 7087
rect 6153 6953 6167 6967
rect 6133 6890 6147 6904
rect 6153 6853 6167 6867
rect 6113 6833 6127 6847
rect 6093 6350 6107 6364
rect 6093 6293 6107 6307
rect 6133 6636 6147 6650
rect 6333 7413 6347 7427
rect 6313 7373 6327 7387
rect 6313 7333 6327 7347
rect 6273 7156 6287 7170
rect 6253 6993 6267 7007
rect 6233 6973 6247 6987
rect 6213 6833 6227 6847
rect 6233 6793 6247 6807
rect 6193 6636 6207 6650
rect 6173 6590 6187 6604
rect 6213 6533 6227 6547
rect 6253 6453 6267 6467
rect 6213 6416 6227 6430
rect 6133 6373 6147 6387
rect 6193 6370 6207 6384
rect 6113 6233 6127 6247
rect 6093 6193 6107 6207
rect 6193 6193 6207 6207
rect 6073 6133 6087 6147
rect 6093 6116 6107 6130
rect 6153 6116 6167 6130
rect 5933 5953 5947 5967
rect 6032 5953 6046 5967
rect 6053 5953 6067 5967
rect 5913 5553 5927 5567
rect 5893 5453 5907 5467
rect 5973 5896 5987 5910
rect 6173 6070 6187 6084
rect 6193 6053 6207 6067
rect 6153 5893 6167 5907
rect 6093 5876 6107 5890
rect 6013 5853 6027 5867
rect 5993 5753 6007 5767
rect 5973 5593 5987 5607
rect 5973 5376 5987 5390
rect 5733 5330 5747 5344
rect 5873 5333 5887 5347
rect 5713 5153 5727 5167
rect 5953 5330 5967 5344
rect 5913 5253 5927 5267
rect 6053 5833 6067 5847
rect 6113 5833 6127 5847
rect 6053 5793 6067 5807
rect 6153 5813 6167 5827
rect 6133 5753 6147 5767
rect 6113 5693 6127 5707
rect 6053 5596 6067 5610
rect 6073 5550 6087 5564
rect 6133 5413 6147 5427
rect 6113 5333 6127 5347
rect 6013 5293 6027 5307
rect 6133 5233 6147 5247
rect 5973 5153 5987 5167
rect 5813 5113 5827 5127
rect 6113 5093 6127 5107
rect 5733 5073 5747 5087
rect 5773 5073 5787 5087
rect 5853 5050 5867 5064
rect 5973 5056 5987 5070
rect 5753 5030 5767 5044
rect 5713 5013 5727 5027
rect 5693 4893 5707 4907
rect 5733 4993 5747 5007
rect 6173 5713 6187 5727
rect 6173 5533 6187 5547
rect 6593 8753 6607 8767
rect 6553 8673 6567 8687
rect 6533 8413 6547 8427
rect 6513 8253 6527 8267
rect 6473 8196 6487 8210
rect 6513 8196 6527 8210
rect 6473 8013 6487 8027
rect 6413 7973 6427 7987
rect 6513 8073 6527 8087
rect 6493 7993 6507 8007
rect 6433 7913 6447 7927
rect 6413 7893 6427 7907
rect 6393 7793 6407 7807
rect 6373 7413 6387 7427
rect 6493 7930 6507 7944
rect 6453 7793 6467 7807
rect 6493 7676 6507 7690
rect 6433 7613 6447 7627
rect 6393 7373 6407 7387
rect 6353 7313 6367 7327
rect 6353 7292 6367 7306
rect 6293 6553 6307 6567
rect 6293 6416 6307 6430
rect 6293 6373 6307 6387
rect 6273 6053 6287 6067
rect 6333 6993 6347 7007
rect 6333 6733 6347 6747
rect 6653 8773 6667 8787
rect 6633 8553 6647 8567
rect 6593 8450 6607 8464
rect 6633 8353 6647 8367
rect 6653 8253 6667 8267
rect 6773 9490 6787 9504
rect 6833 9490 6847 9504
rect 6833 9413 6847 9427
rect 6873 9413 6887 9427
rect 6713 9393 6727 9407
rect 6713 9273 6727 9287
rect 6713 9190 6727 9204
rect 6713 9133 6727 9147
rect 6713 9013 6727 9027
rect 6753 9013 6767 9027
rect 6793 9016 6807 9030
rect 6853 9333 6867 9347
rect 7053 9873 7067 9887
rect 7033 9693 7047 9707
rect 6973 9573 6987 9587
rect 7013 9553 7027 9567
rect 6953 9536 6967 9550
rect 6993 9536 7007 9550
rect 6993 9493 7007 9507
rect 6973 9453 6987 9467
rect 6973 9373 6987 9387
rect 6893 9272 6907 9286
rect 6953 9273 6967 9287
rect 6933 9236 6947 9250
rect 6853 9190 6867 9204
rect 6953 9190 6967 9204
rect 6913 9073 6927 9087
rect 6893 9053 6907 9067
rect 6733 8973 6747 8987
rect 6773 8973 6787 8987
rect 6753 8893 6767 8907
rect 6733 8716 6747 8730
rect 6713 8593 6727 8607
rect 6713 8450 6727 8464
rect 6753 8670 6767 8684
rect 6733 8353 6747 8367
rect 6853 8970 6867 8984
rect 6893 8970 6907 8984
rect 6813 8853 6827 8867
rect 6813 8753 6827 8767
rect 6853 8753 6867 8767
rect 6853 8716 6867 8730
rect 6893 8713 6907 8727
rect 6833 8670 6847 8684
rect 6873 8670 6887 8684
rect 6873 8593 6887 8607
rect 6933 9016 6947 9030
rect 6933 8933 6947 8947
rect 6973 8716 6987 8730
rect 6953 8653 6967 8667
rect 6973 8513 6987 8527
rect 6953 8493 6967 8507
rect 6793 8353 6807 8367
rect 6773 8253 6787 8267
rect 6733 8196 6747 8210
rect 6893 8313 6907 8327
rect 6973 8273 6987 8287
rect 7053 9613 7067 9627
rect 7053 9393 7067 9407
rect 7053 9236 7067 9250
rect 7173 10233 7187 10247
rect 7113 10213 7127 10227
rect 7093 10093 7107 10107
rect 7133 10113 7147 10127
rect 7133 10033 7147 10047
rect 7153 9933 7167 9947
rect 7533 10573 7547 10587
rect 7453 10530 7467 10544
rect 7393 10513 7407 10527
rect 7433 10513 7447 10527
rect 7473 10513 7487 10527
rect 7272 10473 7286 10487
rect 7293 10473 7307 10487
rect 7253 10373 7267 10387
rect 7213 10313 7227 10327
rect 7213 10233 7227 10247
rect 7253 10233 7267 10247
rect 7193 10213 7207 10227
rect 7233 10056 7247 10070
rect 7173 9873 7187 9887
rect 7233 9833 7247 9847
rect 7273 9793 7287 9807
rect 7273 9772 7287 9786
rect 7193 9756 7207 9770
rect 7233 9756 7247 9770
rect 7113 9693 7127 9707
rect 7233 9673 7247 9687
rect 7213 9613 7227 9627
rect 7173 9553 7187 9567
rect 7113 9393 7127 9407
rect 7233 9490 7247 9504
rect 7253 9473 7267 9487
rect 7193 9393 7207 9407
rect 7133 9333 7147 9347
rect 7213 9313 7227 9327
rect 7133 9273 7147 9287
rect 7133 9193 7147 9207
rect 7073 9113 7087 9127
rect 7073 9016 7087 9030
rect 7033 8793 7047 8807
rect 7033 8373 7047 8387
rect 7113 8933 7127 8947
rect 7193 9190 7207 9204
rect 7153 8833 7167 8847
rect 7113 8716 7127 8730
rect 7173 8653 7187 8667
rect 7133 8573 7147 8587
rect 7093 8553 7107 8567
rect 7073 8533 7087 8547
rect 7053 8333 7067 8347
rect 7013 8253 7027 8267
rect 7173 8496 7187 8510
rect 7093 8413 7107 8427
rect 6993 8213 7007 8227
rect 7073 8213 7087 8227
rect 6893 8193 6907 8207
rect 6653 7976 6667 7990
rect 6653 7913 6667 7927
rect 6793 8150 6807 8164
rect 6753 8113 6767 8127
rect 6693 8033 6707 8047
rect 6673 7833 6687 7847
rect 6733 7976 6747 7990
rect 6753 7873 6767 7887
rect 6693 7813 6707 7827
rect 6693 7753 6707 7767
rect 6633 7733 6647 7747
rect 6553 7613 6567 7627
rect 6673 7713 6687 7727
rect 6713 7676 6727 7690
rect 6693 7630 6707 7644
rect 6633 7593 6647 7607
rect 7013 8150 7027 8164
rect 6853 8073 6867 8087
rect 6893 8073 6907 8087
rect 6873 8013 6887 8027
rect 6853 7853 6867 7867
rect 7073 8033 7087 8047
rect 6973 7973 6987 7987
rect 7033 7976 7047 7990
rect 7173 8433 7187 8447
rect 7153 8393 7167 8407
rect 7153 8372 7167 8386
rect 7113 8253 7127 8267
rect 6953 7833 6967 7847
rect 6813 7773 6827 7787
rect 6893 7676 6907 7690
rect 6933 7676 6947 7690
rect 7053 7930 7067 7944
rect 7013 7893 7027 7907
rect 7053 7893 7067 7907
rect 7033 7713 7047 7727
rect 7033 7673 7047 7687
rect 6893 7633 6907 7647
rect 6993 7630 7007 7644
rect 7033 7630 7047 7644
rect 7033 7593 7047 7607
rect 6713 7553 6727 7567
rect 6753 7553 6767 7567
rect 6953 7553 6967 7567
rect 7013 7553 7027 7567
rect 6573 7513 6587 7527
rect 6613 7513 6627 7527
rect 6993 7493 7007 7507
rect 6833 7430 6847 7444
rect 7013 7453 7027 7467
rect 7093 7753 7107 7767
rect 7153 8153 7167 8167
rect 7153 8013 7167 8027
rect 7133 7973 7147 7987
rect 7133 7630 7147 7644
rect 7113 7493 7127 7507
rect 7053 7433 7067 7447
rect 7093 7436 7107 7450
rect 6493 7390 6507 7404
rect 6493 7313 6507 7327
rect 6433 7293 6447 7307
rect 6513 7293 6527 7307
rect 6513 7253 6527 7267
rect 6413 7213 6427 7227
rect 6513 7173 6527 7187
rect 6373 7156 6387 7170
rect 6433 7156 6447 7170
rect 6473 7156 6487 7170
rect 6373 7113 6387 7127
rect 6413 7110 6427 7124
rect 6373 7073 6387 7087
rect 6413 7073 6427 7087
rect 6353 6693 6367 6707
rect 6353 6233 6367 6247
rect 6333 6153 6347 6167
rect 6313 6033 6327 6047
rect 6493 7093 6507 7107
rect 6453 7033 6467 7047
rect 6413 6936 6427 6950
rect 6433 6673 6447 6687
rect 6593 7410 6607 7424
rect 6993 7410 7007 7424
rect 6553 7373 6567 7387
rect 6633 7373 6647 7387
rect 6613 7333 6627 7347
rect 6553 7156 6567 7170
rect 6533 7093 6547 7107
rect 6553 7073 6567 7087
rect 6513 7053 6527 7067
rect 6533 7033 6547 7047
rect 6573 6773 6587 6787
rect 6533 6673 6547 6687
rect 6493 6636 6507 6650
rect 6473 6590 6487 6604
rect 6613 7213 6627 7227
rect 6613 7156 6627 7170
rect 6613 7113 6627 7127
rect 6613 6936 6627 6950
rect 6673 7333 6687 7347
rect 6853 7333 6867 7347
rect 6773 7293 6787 7307
rect 6653 7233 6667 7247
rect 6713 7156 6727 7170
rect 6753 7156 6767 7170
rect 6793 7156 6807 7170
rect 6693 7093 6707 7107
rect 6733 7073 6747 7087
rect 6773 7053 6787 7067
rect 6653 6993 6667 7007
rect 6693 6936 6707 6950
rect 6593 6693 6607 6707
rect 6493 6553 6507 6567
rect 6433 6473 6447 6487
rect 6453 6370 6467 6384
rect 6493 6373 6507 6387
rect 6513 6333 6527 6347
rect 6413 6193 6427 6207
rect 6453 6116 6467 6130
rect 6493 6116 6507 6130
rect 6413 6070 6427 6084
rect 6253 5973 6267 5987
rect 6373 5973 6387 5987
rect 6213 5893 6227 5907
rect 6513 6070 6527 6084
rect 6353 5870 6367 5884
rect 6452 5870 6466 5884
rect 6473 5876 6487 5890
rect 6213 5833 6227 5847
rect 6513 5830 6527 5844
rect 6593 6293 6607 6307
rect 6573 6116 6587 6130
rect 6593 5873 6607 5887
rect 6553 5793 6567 5807
rect 6273 5713 6287 5727
rect 6793 7013 6807 7027
rect 6873 7313 6887 7327
rect 6933 7213 6947 7227
rect 7113 7393 7127 7407
rect 7093 7253 7107 7267
rect 7073 7213 7087 7227
rect 7093 7193 7107 7207
rect 7033 7173 7047 7187
rect 7033 7156 7047 7170
rect 7093 7156 7107 7170
rect 7153 7333 7167 7347
rect 7153 7213 7167 7227
rect 6933 7113 6947 7127
rect 6873 6993 6887 7007
rect 6993 6993 7007 7007
rect 6893 6953 6907 6967
rect 6853 6936 6867 6950
rect 6933 6936 6947 6950
rect 7053 7110 7067 7124
rect 7113 7133 7127 7147
rect 7093 7073 7107 7087
rect 7013 6973 7027 6987
rect 7053 6953 7067 6967
rect 6773 6913 6787 6927
rect 6733 6890 6747 6904
rect 6813 6873 6827 6887
rect 6693 6753 6707 6767
rect 6673 6636 6687 6650
rect 6633 6473 6647 6487
rect 7093 6913 7107 6927
rect 7053 6873 7067 6887
rect 6913 6853 6927 6867
rect 7133 7053 7147 7067
rect 7133 6973 7147 6987
rect 7113 6833 7127 6847
rect 7133 6793 7147 6807
rect 7193 8393 7207 8407
rect 7253 9153 7267 9167
rect 7493 10453 7507 10467
rect 7473 10433 7487 10447
rect 7313 10373 7327 10387
rect 7513 10413 7527 10427
rect 7473 10333 7487 10347
rect 7453 10313 7467 10327
rect 7333 10276 7347 10290
rect 7413 10276 7427 10290
rect 7433 10230 7447 10244
rect 7593 10576 7607 10590
rect 7553 10533 7567 10547
rect 7553 10273 7567 10287
rect 7533 10193 7547 10207
rect 7433 10153 7447 10167
rect 7352 10053 7366 10067
rect 7373 10053 7387 10067
rect 7493 10093 7507 10107
rect 7453 10056 7467 10070
rect 7613 10493 7627 10507
rect 7693 11293 7707 11307
rect 8073 12073 8087 12087
rect 7933 12033 7947 12047
rect 7793 11833 7807 11847
rect 7853 11836 7867 11850
rect 7913 11833 7927 11847
rect 7873 11790 7887 11804
rect 7913 11790 7927 11804
rect 7833 11773 7847 11787
rect 7873 11713 7887 11727
rect 7993 11713 8007 11727
rect 7833 11616 7847 11630
rect 7913 11616 7927 11630
rect 8413 11993 8427 12007
rect 8193 11873 8207 11887
rect 8233 11853 8247 11867
rect 8133 11836 8147 11850
rect 8193 11836 8207 11850
rect 8113 11753 8127 11767
rect 8233 11733 8247 11747
rect 8173 11713 8187 11727
rect 8073 11613 8087 11627
rect 8253 11590 8267 11604
rect 8413 11853 8427 11867
rect 8473 11836 8487 11850
rect 8533 11836 8547 11850
rect 8453 11713 8467 11727
rect 8393 11693 8407 11707
rect 8393 11590 8407 11604
rect 7893 11553 7907 11567
rect 7833 11533 7847 11547
rect 7793 11373 7807 11387
rect 7813 11316 7827 11330
rect 8413 11533 8427 11547
rect 7953 11493 7967 11507
rect 7913 11473 7927 11487
rect 7873 11316 7887 11330
rect 8313 11473 8327 11487
rect 8033 11453 8047 11467
rect 7953 11393 7967 11407
rect 7833 11273 7847 11287
rect 7893 11270 7907 11284
rect 7893 11096 7907 11110
rect 7873 11050 7887 11064
rect 8013 11313 8027 11327
rect 7993 11096 8007 11110
rect 7953 11013 7967 11027
rect 7993 11013 8007 11027
rect 7813 10893 7827 10907
rect 7813 10796 7827 10810
rect 7873 10796 7887 10810
rect 7773 10733 7787 10747
rect 7813 10733 7827 10747
rect 7753 10576 7767 10590
rect 7733 10530 7747 10544
rect 7713 10493 7727 10507
rect 7673 10473 7687 10487
rect 7653 10373 7667 10387
rect 7953 10693 7967 10707
rect 7873 10633 7887 10647
rect 7853 10473 7867 10487
rect 7973 10530 7987 10544
rect 7973 10513 7987 10527
rect 7873 10453 7887 10467
rect 8013 10433 8027 10447
rect 8093 11316 8107 11330
rect 8173 11316 8187 11330
rect 8133 11233 8147 11247
rect 8093 11193 8107 11207
rect 8453 11393 8467 11407
rect 8493 11333 8507 11347
rect 8373 11293 8387 11307
rect 8313 11213 8327 11227
rect 8153 11153 8167 11167
rect 8073 11133 8087 11147
rect 8133 11133 8147 11147
rect 8053 10793 8067 10807
rect 8053 10673 8067 10687
rect 7873 10393 7887 10407
rect 8033 10393 8047 10407
rect 7853 10333 7867 10347
rect 7813 10293 7827 10307
rect 7713 10276 7727 10290
rect 7833 10250 7847 10264
rect 8213 11093 8227 11107
rect 8113 11050 8127 11064
rect 8253 11013 8267 11027
rect 8213 10913 8227 10927
rect 8253 10913 8267 10927
rect 8113 10833 8127 10847
rect 8173 10796 8187 10810
rect 8153 10750 8167 10764
rect 8113 10653 8127 10667
rect 8233 10796 8247 10810
rect 8273 10793 8287 10807
rect 8273 10750 8287 10764
rect 8253 10653 8267 10667
rect 8233 10633 8247 10647
rect 8213 10576 8227 10590
rect 8433 11253 8447 11267
rect 8653 12136 8667 12150
rect 8733 12136 8747 12150
rect 8673 12090 8687 12104
rect 8633 12033 8647 12047
rect 9093 12153 9107 12167
rect 9793 12153 9807 12167
rect 9353 12133 9367 12147
rect 9253 12110 9267 12124
rect 9373 12116 9387 12130
rect 9513 12116 9527 12130
rect 9633 12110 9647 12124
rect 8573 11993 8587 12007
rect 8733 11993 8747 12007
rect 8553 11810 8567 11824
rect 8553 11613 8567 11627
rect 8533 11253 8547 11267
rect 9093 12090 9107 12104
rect 9389 12073 9403 12087
rect 9497 12073 9511 12087
rect 9433 12053 9447 12067
rect 9473 12053 9487 12067
rect 8933 11953 8947 11967
rect 8813 11893 8827 11907
rect 8693 11873 8707 11887
rect 8733 11836 8747 11850
rect 8613 11713 8627 11727
rect 10413 12193 10427 12207
rect 9893 12133 9907 12147
rect 10113 12136 10127 12150
rect 10373 12136 10387 12150
rect 10453 12173 10467 12187
rect 11393 12173 11407 12187
rect 11473 12173 11487 12187
rect 9933 12110 9947 12124
rect 9793 12033 9807 12047
rect 10593 12136 10607 12150
rect 10653 12136 10667 12150
rect 10693 12136 10707 12150
rect 10753 12136 10767 12150
rect 10913 12136 10927 12150
rect 10953 12136 10967 12150
rect 11053 12136 11067 12150
rect 11193 12136 11207 12150
rect 11373 12136 11387 12150
rect 10133 12073 10147 12087
rect 9933 12013 9947 12027
rect 10013 11993 10027 12007
rect 9493 11893 9507 11907
rect 8973 11873 8987 11887
rect 9433 11873 9447 11887
rect 8933 11833 8947 11847
rect 9013 11833 9027 11847
rect 9153 11836 9167 11850
rect 9193 11836 9207 11850
rect 9233 11836 9247 11850
rect 9293 11836 9307 11850
rect 8753 11773 8767 11787
rect 8813 11773 8827 11787
rect 8953 11773 8967 11787
rect 8713 11673 8727 11687
rect 8713 11616 8727 11630
rect 8893 11616 8907 11630
rect 8613 11570 8627 11584
rect 8653 11570 8667 11584
rect 8593 11553 8607 11567
rect 8693 11553 8707 11567
rect 8753 11553 8767 11567
rect 8733 11533 8747 11547
rect 8693 11513 8707 11527
rect 8593 11333 8607 11347
rect 8733 11336 8747 11350
rect 8573 11293 8587 11307
rect 8553 11233 8567 11247
rect 8473 11213 8487 11227
rect 8493 11153 8507 11167
rect 8373 11096 8387 11110
rect 8413 11096 8427 11110
rect 8353 11050 8367 11064
rect 8393 11013 8407 11027
rect 8453 11053 8467 11067
rect 8453 10973 8467 10987
rect 8433 10913 8447 10927
rect 8653 11313 8667 11327
rect 8653 11270 8667 11284
rect 8693 11270 8707 11284
rect 8793 11273 8807 11287
rect 8873 11273 8887 11287
rect 8853 11233 8867 11247
rect 8973 11513 8987 11527
rect 8933 11473 8947 11487
rect 9253 11790 9267 11804
rect 9293 11773 9307 11787
rect 9233 11693 9247 11707
rect 9273 11693 9287 11707
rect 9413 11693 9427 11707
rect 9253 11570 9267 11584
rect 9213 11553 9227 11567
rect 9153 11453 9167 11467
rect 9213 11373 9227 11387
rect 9213 11336 9227 11350
rect 9053 11296 9067 11310
rect 9273 11373 9287 11387
rect 9173 11290 9187 11304
rect 9253 11293 9267 11307
rect 9173 11253 9187 11267
rect 8893 11193 8907 11207
rect 9013 11193 9027 11207
rect 8873 11153 8887 11167
rect 9053 11153 9067 11167
rect 9013 11096 9027 11110
rect 8613 11070 8627 11084
rect 8753 11070 8767 11084
rect 8873 11076 8887 11090
rect 8953 11073 8967 11087
rect 8613 11033 8627 11047
rect 8873 10993 8887 11007
rect 8913 10993 8927 11007
rect 8733 10973 8747 10987
rect 8633 10933 8647 10947
rect 8593 10833 8607 10847
rect 8393 10796 8407 10810
rect 8453 10793 8467 10807
rect 8753 10933 8767 10947
rect 8733 10913 8747 10927
rect 8733 10873 8747 10887
rect 8693 10816 8707 10830
rect 8673 10796 8687 10810
rect 8413 10733 8427 10747
rect 8313 10613 8327 10627
rect 8433 10553 8447 10567
rect 8193 10530 8207 10544
rect 8413 10533 8427 10547
rect 8273 10513 8287 10527
rect 8233 10453 8247 10467
rect 8193 10433 8207 10447
rect 8073 10373 8087 10387
rect 8173 10373 8187 10387
rect 8613 10733 8627 10747
rect 8553 10673 8567 10687
rect 8513 10576 8527 10590
rect 8533 10530 8547 10544
rect 8573 10530 8587 10544
rect 8472 10473 8486 10487
rect 8493 10473 8507 10487
rect 8513 10433 8527 10447
rect 8493 10413 8507 10427
rect 8473 10393 8487 10407
rect 8453 10373 8467 10387
rect 8573 10373 8587 10387
rect 8613 10373 8627 10387
rect 8413 10353 8427 10367
rect 8193 10313 8207 10327
rect 8253 10313 8267 10327
rect 8173 10293 8187 10307
rect 8033 10256 8047 10270
rect 7673 10230 7687 10244
rect 7773 10233 7787 10247
rect 7593 10193 7607 10207
rect 7693 10193 7707 10207
rect 7673 10153 7687 10167
rect 7553 10056 7567 10070
rect 7353 10010 7367 10024
rect 7393 9953 7407 9967
rect 7373 9873 7387 9887
rect 7333 9773 7347 9787
rect 7313 9493 7327 9507
rect 7293 9313 7307 9327
rect 7293 9190 7307 9204
rect 7353 9213 7367 9227
rect 7333 9153 7347 9167
rect 7393 9813 7407 9827
rect 7433 9933 7447 9947
rect 7513 10010 7527 10024
rect 7573 9993 7587 10007
rect 7553 9973 7567 9987
rect 7613 9913 7627 9927
rect 7433 9793 7447 9807
rect 7553 9793 7567 9807
rect 7593 9793 7607 9807
rect 7493 9756 7507 9770
rect 7413 9732 7427 9746
rect 7513 9710 7527 9724
rect 7553 9710 7567 9724
rect 7473 9613 7487 9627
rect 7413 9593 7427 9607
rect 7553 9593 7567 9607
rect 7493 9536 7507 9550
rect 7533 9493 7547 9507
rect 7513 9373 7527 9387
rect 7513 9313 7527 9327
rect 7473 9273 7487 9287
rect 7433 9236 7447 9250
rect 7413 9190 7427 9204
rect 7353 9113 7367 9127
rect 7333 9016 7347 9030
rect 7293 8953 7307 8967
rect 7333 8953 7347 8967
rect 7273 8893 7287 8907
rect 7293 8713 7307 8727
rect 7293 8593 7307 8607
rect 7313 8493 7327 8507
rect 7313 8450 7327 8464
rect 7233 8433 7247 8447
rect 7213 8373 7227 8387
rect 7253 8253 7267 8267
rect 7293 8196 7307 8210
rect 7233 8150 7247 8164
rect 7213 8033 7227 8047
rect 7273 7973 7287 7987
rect 7213 7930 7227 7944
rect 7253 7930 7267 7944
rect 7293 7930 7307 7944
rect 7193 7893 7207 7907
rect 7213 7676 7227 7690
rect 7273 7676 7287 7690
rect 7313 7676 7327 7690
rect 7233 7630 7247 7644
rect 7253 7613 7267 7627
rect 7193 7553 7207 7567
rect 7213 7493 7227 7507
rect 7233 7456 7247 7470
rect 7213 7436 7227 7450
rect 7213 7313 7227 7327
rect 7233 7193 7247 7207
rect 7193 7133 7207 7147
rect 7273 7593 7287 7607
rect 7353 8893 7367 8907
rect 7333 7613 7347 7627
rect 7453 8873 7467 8887
rect 7413 8753 7427 8767
rect 7373 8716 7387 8730
rect 7453 8716 7467 8730
rect 7433 8670 7447 8684
rect 7493 8670 7507 8684
rect 7433 8573 7447 8587
rect 7393 8553 7407 8567
rect 7433 8513 7447 8527
rect 7373 8493 7387 8507
rect 7453 8496 7467 8510
rect 7493 8496 7507 8510
rect 7433 8450 7447 8464
rect 7513 8453 7527 8467
rect 7493 8433 7507 8447
rect 7473 8413 7487 8427
rect 7453 8393 7467 8407
rect 7393 8333 7407 8347
rect 7453 8333 7467 8347
rect 7373 8033 7387 8047
rect 7453 8053 7467 8067
rect 7433 7930 7447 7944
rect 7433 7893 7447 7907
rect 7413 7733 7427 7747
rect 7353 7593 7367 7607
rect 7413 7553 7427 7567
rect 7413 7513 7427 7527
rect 7353 7493 7367 7507
rect 7373 7456 7387 7470
rect 7413 7453 7427 7467
rect 7293 7410 7307 7424
rect 7353 7410 7367 7424
rect 7393 7410 7407 7424
rect 7273 7393 7287 7407
rect 7333 7393 7347 7407
rect 7313 7213 7327 7227
rect 7253 7153 7267 7167
rect 7433 7213 7447 7227
rect 7413 7193 7427 7207
rect 7533 8433 7547 8447
rect 7573 9373 7587 9387
rect 7833 10092 7847 10106
rect 7753 10056 7767 10070
rect 7793 10056 7807 10070
rect 7693 9913 7707 9927
rect 7633 9853 7647 9867
rect 7672 9853 7686 9867
rect 7693 9853 7707 9867
rect 7633 9756 7647 9770
rect 7813 9793 7827 9807
rect 7733 9756 7747 9770
rect 7773 9756 7787 9770
rect 7833 9756 7847 9770
rect 7673 9713 7687 9727
rect 7753 9710 7767 9724
rect 7653 9633 7667 9647
rect 7713 9633 7727 9647
rect 8173 10253 8187 10267
rect 8153 10113 8167 10127
rect 7913 10073 7927 10087
rect 7913 9813 7927 9827
rect 7873 9753 7887 9767
rect 8013 10093 8027 10107
rect 7973 10056 7987 10070
rect 8273 10233 8287 10247
rect 8213 10173 8227 10187
rect 8173 10056 8187 10070
rect 7993 9993 8007 10007
rect 8233 10113 8247 10127
rect 8213 9953 8227 9967
rect 8413 10256 8427 10270
rect 8293 10113 8307 10127
rect 8373 10113 8387 10127
rect 8333 10056 8347 10070
rect 8273 9993 8287 10007
rect 8393 10056 8407 10070
rect 8493 10056 8507 10070
rect 8533 10056 8547 10070
rect 8693 10750 8707 10764
rect 8713 10613 8727 10627
rect 8733 10530 8747 10544
rect 8653 10293 8667 10307
rect 8713 10273 8727 10287
rect 8393 10013 8407 10027
rect 8313 9993 8327 10007
rect 8373 9993 8387 10007
rect 8553 10010 8567 10024
rect 8493 9933 8507 9947
rect 8033 9913 8047 9927
rect 7993 9853 8007 9867
rect 8113 9873 8127 9887
rect 8033 9793 8047 9807
rect 8113 9773 8127 9787
rect 8213 9773 8227 9787
rect 8513 9776 8527 9790
rect 8033 9756 8047 9770
rect 8093 9730 8107 9744
rect 8133 9733 8147 9747
rect 7933 9693 7947 9707
rect 7873 9673 7887 9687
rect 8053 9710 8067 9724
rect 8093 9710 8107 9724
rect 8013 9653 8027 9667
rect 7853 9593 7867 9607
rect 8033 9553 8047 9567
rect 7673 9533 7687 9547
rect 7753 9536 7767 9550
rect 7973 9533 7987 9547
rect 7673 9490 7687 9504
rect 7653 9473 7667 9487
rect 7773 9490 7787 9504
rect 7973 9490 7987 9504
rect 8013 9490 8027 9504
rect 8053 9473 8067 9487
rect 7733 9453 7747 9467
rect 8113 9433 8127 9447
rect 7653 9393 7667 9407
rect 7713 9373 7727 9387
rect 7793 9256 7807 9270
rect 7673 9213 7687 9227
rect 7833 9210 7847 9224
rect 7953 9216 7967 9230
rect 8093 9216 8107 9230
rect 8093 9173 8107 9187
rect 7753 9133 7767 9147
rect 7793 9133 7807 9147
rect 7633 9093 7647 9107
rect 7613 9033 7627 9047
rect 7753 9033 7767 9047
rect 7673 8793 7687 8807
rect 7613 8712 7627 8726
rect 7713 8773 7727 8787
rect 7613 8670 7627 8684
rect 7653 8670 7667 8684
rect 7693 8670 7707 8684
rect 7753 8673 7767 8687
rect 7753 8613 7767 8627
rect 7573 8553 7587 8567
rect 7553 8413 7567 8427
rect 7513 8373 7527 8387
rect 7653 8533 7667 8547
rect 7613 8513 7627 8527
rect 7593 8473 7607 8487
rect 7593 8353 7607 8367
rect 7613 8333 7627 8347
rect 7573 8253 7587 8267
rect 8213 9733 8227 9747
rect 8353 9736 8367 9750
rect 8153 9693 8167 9707
rect 8293 9633 8307 9647
rect 8193 9613 8207 9627
rect 8213 9553 8227 9567
rect 8193 9490 8207 9504
rect 8253 9536 8267 9550
rect 8413 9573 8427 9587
rect 8273 9490 8287 9504
rect 8313 9473 8327 9487
rect 8333 9413 8347 9427
rect 8213 9333 8227 9347
rect 8153 9273 8167 9287
rect 8253 9273 8267 9287
rect 8133 9256 8147 9270
rect 8153 9210 8167 9224
rect 8253 9210 8267 9224
rect 8113 9093 8127 9107
rect 8213 9093 8227 9107
rect 7873 9016 7887 9030
rect 7913 9013 7927 9027
rect 7973 8996 7987 9010
rect 8173 8990 8187 9004
rect 8353 9333 8367 9347
rect 8333 9133 8347 9147
rect 8313 9053 8327 9067
rect 8313 8990 8327 9004
rect 8393 9253 8407 9267
rect 7833 8973 7847 8987
rect 7793 8533 7807 8547
rect 8333 8950 8347 8964
rect 8313 8893 8327 8907
rect 8393 8950 8407 8964
rect 7853 8753 7867 8767
rect 8013 8716 8027 8730
rect 8053 8713 8067 8727
rect 7873 8670 7887 8684
rect 7993 8670 8007 8684
rect 7893 8593 7907 8607
rect 7953 8593 7967 8607
rect 7873 8573 7887 8587
rect 7853 8513 7867 8527
rect 7793 8476 7807 8490
rect 7913 8476 7927 8490
rect 8053 8470 8067 8484
rect 8213 8753 8227 8767
rect 8253 8716 8267 8730
rect 8193 8573 8207 8587
rect 8273 8673 8287 8687
rect 8233 8533 8247 8547
rect 8193 8470 8207 8484
rect 7913 8433 7927 8447
rect 7893 8393 7907 8407
rect 8173 8393 8187 8407
rect 8033 8293 8047 8307
rect 7713 8253 7727 8267
rect 7653 8213 7667 8227
rect 7553 8196 7567 8210
rect 7533 8133 7547 8147
rect 7553 8053 7567 8067
rect 7533 8013 7547 8027
rect 7493 7893 7507 7907
rect 7493 7833 7507 7847
rect 7553 7833 7567 7847
rect 7493 7773 7507 7787
rect 7593 8153 7607 8167
rect 7673 8153 7687 8167
rect 8253 8433 8267 8447
rect 8213 8373 8227 8387
rect 8273 8373 8287 8387
rect 8193 8313 8207 8327
rect 7873 8176 7887 8190
rect 7973 8176 7987 8190
rect 8013 8173 8027 8187
rect 8073 8173 8087 8187
rect 8113 8173 8127 8187
rect 7993 8153 8007 8167
rect 7713 8133 7727 8147
rect 7613 8093 7627 8107
rect 7633 8013 7647 8027
rect 7593 7933 7607 7947
rect 7573 7813 7587 7827
rect 7553 7733 7567 7747
rect 7593 7713 7607 7727
rect 7693 7976 7707 7990
rect 7733 7973 7747 7987
rect 7793 7956 7807 7970
rect 7833 7956 7847 7970
rect 7633 7693 7647 7707
rect 7613 7650 7627 7664
rect 7513 7593 7527 7607
rect 7553 7593 7567 7607
rect 7473 7493 7487 7507
rect 7333 7173 7347 7187
rect 7453 7173 7467 7187
rect 7233 7093 7247 7107
rect 7353 7113 7367 7127
rect 7333 7093 7347 7107
rect 7293 7073 7307 7087
rect 7213 7033 7227 7047
rect 7233 7013 7247 7027
rect 7313 7013 7327 7027
rect 7213 6973 7227 6987
rect 7253 6973 7267 6987
rect 7093 6753 7107 6767
rect 7153 6753 7167 6767
rect 6873 6693 6887 6707
rect 7173 6653 7187 6667
rect 6713 6636 6727 6650
rect 6773 6636 6787 6650
rect 6813 6636 6827 6650
rect 6893 6613 6907 6627
rect 6713 6593 6727 6607
rect 6753 6493 6767 6507
rect 6713 6473 6727 6487
rect 6693 6453 6707 6467
rect 6653 6433 6667 6447
rect 6693 6353 6707 6367
rect 6773 6353 6787 6367
rect 6673 6293 6687 6307
rect 6633 6116 6647 6130
rect 6633 5973 6647 5987
rect 6273 5653 6287 5667
rect 6293 5633 6307 5647
rect 6353 5573 6367 5587
rect 6313 5513 6327 5527
rect 6193 5473 6207 5487
rect 6273 5473 6287 5487
rect 6213 5433 6227 5447
rect 6193 5330 6207 5344
rect 6193 5113 6207 5127
rect 6153 5093 6167 5107
rect 6133 5056 6147 5070
rect 6133 5013 6147 5027
rect 5853 4973 5867 4987
rect 6133 4973 6147 4987
rect 6173 4973 6187 4987
rect 5773 4953 5787 4967
rect 5813 4893 5827 4907
rect 6133 4952 6147 4966
rect 5913 4933 5927 4947
rect 5973 4913 5987 4927
rect 5953 4893 5967 4907
rect 5933 4873 5947 4887
rect 5833 4810 5847 4824
rect 5873 4810 5887 4824
rect 5773 4753 5787 4767
rect 5753 4673 5767 4687
rect 5893 4673 5907 4687
rect 5793 4653 5807 4667
rect 5873 4653 5887 4667
rect 5913 4653 5927 4667
rect 5773 4633 5787 4647
rect 5853 4613 5867 4627
rect 5713 4493 5727 4507
rect 5753 4493 5767 4507
rect 5853 4573 5867 4587
rect 5873 4556 5887 4570
rect 5853 4510 5867 4524
rect 5893 4513 5907 4527
rect 5813 4493 5827 4507
rect 5853 4473 5867 4487
rect 5893 4472 5907 4486
rect 5773 4453 5787 4467
rect 5853 4452 5867 4466
rect 5913 4453 5927 4467
rect 5793 4433 5807 4447
rect 5733 4373 5747 4387
rect 5753 4290 5767 4304
rect 5813 4290 5827 4304
rect 5793 4273 5807 4287
rect 5753 4233 5767 4247
rect 5713 4213 5727 4227
rect 5713 4173 5727 4187
rect 5773 4213 5787 4227
rect 5753 4073 5767 4087
rect 5913 4373 5927 4387
rect 6033 4810 6047 4824
rect 5993 4733 6007 4747
rect 6013 4613 6027 4627
rect 6013 4533 6027 4547
rect 6033 4493 6047 4507
rect 5973 4453 5987 4467
rect 6013 4453 6027 4467
rect 5953 4433 5967 4447
rect 5953 4353 5967 4367
rect 5853 4193 5867 4207
rect 5793 4173 5807 4187
rect 5813 4053 5827 4067
rect 5713 4033 5727 4047
rect 5773 4036 5787 4050
rect 5873 4033 5887 4047
rect 5693 3692 5707 3706
rect 5673 3473 5687 3487
rect 5753 3973 5767 3987
rect 5753 3913 5767 3927
rect 5873 3973 5887 3987
rect 5873 3933 5887 3947
rect 5793 3893 5807 3907
rect 5853 3893 5867 3907
rect 5753 3816 5767 3830
rect 5793 3816 5807 3830
rect 5813 3770 5827 3784
rect 5873 3733 5887 3747
rect 5793 3713 5807 3727
rect 5733 3593 5747 3607
rect 5713 3513 5727 3527
rect 5773 3553 5787 3567
rect 5873 3693 5887 3707
rect 5913 4233 5927 4247
rect 5913 4173 5927 4187
rect 5933 4073 5947 4087
rect 5913 4053 5927 4067
rect 5933 3816 5947 3830
rect 5913 3733 5927 3747
rect 5933 3553 5947 3567
rect 5872 3473 5886 3487
rect 5853 3453 5867 3467
rect 5753 3433 5767 3447
rect 5693 3393 5707 3407
rect 5713 3373 5727 3387
rect 5673 3353 5687 3367
rect 5653 3293 5667 3307
rect 5833 3353 5847 3367
rect 5813 3333 5827 3347
rect 5773 3313 5787 3327
rect 5693 3250 5707 3264
rect 5733 3250 5747 3264
rect 5793 3293 5807 3307
rect 5773 3173 5787 3187
rect 5813 3250 5827 3264
rect 5813 3213 5827 3227
rect 5813 3173 5827 3187
rect 5613 3153 5627 3167
rect 5653 3153 5667 3167
rect 5793 3153 5807 3167
rect 5753 3073 5767 3087
rect 5653 3033 5667 3047
rect 5593 2996 5607 3010
rect 5573 2853 5587 2867
rect 5553 2776 5567 2790
rect 5753 3013 5767 3027
rect 5693 2996 5707 3010
rect 5633 2953 5647 2967
rect 5613 2773 5627 2787
rect 5573 2730 5587 2744
rect 5473 2693 5487 2707
rect 5253 2673 5267 2687
rect 5513 2693 5527 2707
rect 5493 2613 5507 2627
rect 5193 2513 5207 2527
rect 5233 2513 5247 2527
rect 5173 2493 5187 2507
rect 5493 2493 5507 2507
rect 5113 2476 5127 2490
rect 5033 2413 5047 2427
rect 4993 2313 5007 2327
rect 4993 2292 5007 2306
rect 5033 2292 5047 2306
rect 5013 2256 5027 2270
rect 5073 2256 5087 2270
rect 5033 2210 5047 2224
rect 5013 2153 5027 2167
rect 4993 2093 5007 2107
rect 4993 1793 5007 1807
rect 5093 2113 5107 2127
rect 5073 2093 5087 2107
rect 5193 2433 5207 2447
rect 5133 2053 5147 2067
rect 5033 1956 5047 1970
rect 5113 1956 5127 1970
rect 5153 1956 5167 1970
rect 5013 1573 5027 1587
rect 4973 1436 4987 1450
rect 4993 1413 5007 1427
rect 4913 1293 4927 1307
rect 4953 1293 4967 1307
rect 4733 1213 4747 1227
rect 4573 1153 4587 1167
rect 4673 1153 4687 1167
rect 4473 993 4487 1007
rect 4533 973 4547 987
rect 4433 916 4447 930
rect 4453 870 4467 884
rect 4493 870 4507 884
rect 4533 870 4547 884
rect 4593 993 4607 1007
rect 4513 733 4527 747
rect 4373 696 4387 710
rect 4113 673 4127 687
rect 4093 653 4107 667
rect 4093 573 4107 587
rect 3773 493 3787 507
rect 3973 493 3987 507
rect 3633 393 3647 407
rect 4113 533 4127 547
rect 4173 393 4187 407
rect 3673 370 3687 384
rect 3553 350 3567 364
rect 3473 213 3487 227
rect 3773 370 3787 384
rect 3933 376 3947 390
rect 3733 293 3747 307
rect 3913 213 3927 227
rect 3593 193 3607 207
rect 3633 193 3647 207
rect 3673 193 3687 207
rect 2773 133 2787 147
rect 3853 176 3867 190
rect 4033 173 4047 187
rect 2833 130 2847 144
rect 2833 93 2847 107
rect 3673 130 3687 144
rect 3833 130 3847 144
rect 3913 130 3927 144
rect 4133 376 4147 390
rect 4073 213 4087 227
rect 4433 696 4447 710
rect 4273 651 4287 665
rect 4333 651 4347 665
rect 4412 651 4426 665
rect 4433 653 4447 667
rect 4293 533 4307 547
rect 4293 493 4307 507
rect 4493 453 4507 467
rect 4353 396 4367 410
rect 4293 350 4307 364
rect 4333 350 4347 364
rect 4233 176 4247 190
rect 4153 130 4167 144
rect 4653 913 4667 927
rect 4653 870 4667 884
rect 4553 693 4567 707
rect 4593 696 4607 710
rect 4533 633 4547 647
rect 4533 453 4547 467
rect 4513 393 4527 407
rect 4633 653 4647 667
rect 4613 633 4627 647
rect 4573 433 4587 447
rect 4613 433 4627 447
rect 4893 1190 4907 1204
rect 5213 2153 5227 2167
rect 5133 1910 5147 1924
rect 5193 1910 5207 1924
rect 5093 1773 5107 1787
rect 5113 1736 5127 1750
rect 5353 2456 5367 2470
rect 5493 2450 5507 2464
rect 5533 2573 5547 2587
rect 5653 2933 5667 2947
rect 5533 2493 5547 2507
rect 5633 2493 5647 2507
rect 5553 2450 5567 2464
rect 5573 2433 5587 2447
rect 5473 2353 5487 2367
rect 5513 2353 5527 2367
rect 5453 2313 5467 2327
rect 5293 2256 5307 2270
rect 5433 2253 5447 2267
rect 5273 2210 5287 2224
rect 5293 2193 5307 2207
rect 5253 2013 5267 2027
rect 5233 1753 5247 1767
rect 5153 1653 5167 1667
rect 5073 1633 5087 1647
rect 5093 1633 5107 1647
rect 5133 1473 5147 1487
rect 5033 1393 5047 1407
rect 5093 1390 5107 1404
rect 5033 1273 5047 1287
rect 5073 1273 5087 1287
rect 5113 1213 5127 1227
rect 5073 1190 5087 1204
rect 5013 1113 5027 1127
rect 4993 1073 5007 1087
rect 4733 1033 4747 1047
rect 4773 1033 4787 1047
rect 4773 916 4787 930
rect 4833 913 4847 927
rect 5013 1033 5027 1047
rect 4753 870 4767 884
rect 4813 873 4827 887
rect 5013 870 5027 884
rect 5033 833 5047 847
rect 4973 733 4987 747
rect 4913 697 4927 711
rect 5013 713 5027 727
rect 4933 651 4947 665
rect 5012 651 5026 665
rect 5033 653 5047 667
rect 4833 633 4847 647
rect 4853 613 4867 627
rect 4713 593 4727 607
rect 5113 1013 5127 1027
rect 5173 1573 5187 1587
rect 5233 1390 5247 1404
rect 5433 2210 5447 2224
rect 5333 2193 5347 2207
rect 5313 2173 5327 2187
rect 5373 2073 5387 2087
rect 5373 1993 5387 2007
rect 5493 2256 5507 2270
rect 5533 2256 5547 2270
rect 5613 2313 5627 2327
rect 5613 2273 5627 2287
rect 5473 2153 5487 2167
rect 5413 1956 5427 1970
rect 5453 1956 5467 1970
rect 5293 1793 5307 1807
rect 5273 1773 5287 1787
rect 5273 1690 5287 1704
rect 5273 1553 5287 1567
rect 5213 1353 5227 1367
rect 5173 1133 5187 1147
rect 5153 1073 5167 1087
rect 5133 973 5147 987
rect 5173 916 5187 930
rect 5113 733 5127 747
rect 5073 573 5087 587
rect 5113 573 5127 587
rect 4853 553 4867 567
rect 4793 453 4807 467
rect 4673 413 4687 427
rect 4573 393 4587 407
rect 4633 396 4647 410
rect 5333 1910 5347 1924
rect 5393 1910 5407 1924
rect 5433 1910 5447 1924
rect 5553 2210 5567 2224
rect 5713 2933 5727 2947
rect 5673 2913 5687 2927
rect 5693 2893 5707 2907
rect 5753 2873 5767 2887
rect 5713 2853 5727 2867
rect 5693 2813 5707 2827
rect 5693 2773 5707 2787
rect 5673 2693 5687 2707
rect 5673 2633 5687 2647
rect 5733 2793 5747 2807
rect 5713 2513 5727 2527
rect 5713 2492 5727 2506
rect 5693 2393 5707 2407
rect 5673 2313 5687 2327
rect 5653 2193 5667 2207
rect 5593 2153 5607 2167
rect 5513 2093 5527 2107
rect 5573 2093 5587 2107
rect 5493 1753 5507 1767
rect 5353 1736 5367 1750
rect 5393 1736 5407 1750
rect 5573 1910 5587 1924
rect 5593 1773 5607 1787
rect 5513 1713 5527 1727
rect 5673 2093 5687 2107
rect 5673 2013 5687 2027
rect 5713 1956 5727 1970
rect 5853 3250 5867 3264
rect 5893 3453 5907 3467
rect 5893 3353 5907 3367
rect 5873 3153 5887 3167
rect 5853 3033 5867 3047
rect 5833 2793 5847 2807
rect 5773 2773 5787 2787
rect 5753 2633 5767 2647
rect 5853 2776 5867 2790
rect 5893 2713 5907 2727
rect 5853 2692 5867 2706
rect 5793 2653 5807 2667
rect 5853 2553 5867 2567
rect 5773 2476 5787 2490
rect 5933 3433 5947 3447
rect 5953 3373 5967 3387
rect 6013 4373 6027 4387
rect 6133 4873 6147 4887
rect 6073 4773 6087 4787
rect 6113 4773 6127 4787
rect 6173 4773 6187 4787
rect 6173 4752 6187 4766
rect 6173 4693 6187 4707
rect 6253 4973 6267 4987
rect 6233 4893 6247 4907
rect 6233 4810 6247 4824
rect 6213 4713 6227 4727
rect 6213 4613 6227 4627
rect 6113 4593 6127 4607
rect 6193 4593 6207 4607
rect 6073 4553 6087 4567
rect 6253 4753 6267 4767
rect 6253 4673 6267 4687
rect 6293 5373 6307 5387
rect 6273 4653 6287 4667
rect 6233 4573 6247 4587
rect 6173 4533 6187 4547
rect 6093 4493 6107 4507
rect 6073 4473 6087 4487
rect 6053 4433 6067 4447
rect 6013 4290 6027 4304
rect 6073 4290 6087 4304
rect 6053 4233 6067 4247
rect 6073 4213 6087 4227
rect 6013 4073 6027 4087
rect 6113 4373 6127 4387
rect 6113 4333 6127 4347
rect 6093 4173 6107 4187
rect 6213 4533 6227 4547
rect 6193 4473 6207 4487
rect 6173 4453 6187 4467
rect 6193 4433 6207 4447
rect 6133 4313 6147 4327
rect 6073 4053 6087 4067
rect 6053 4036 6067 4050
rect 6073 3953 6087 3967
rect 6013 3933 6027 3947
rect 6013 3893 6027 3907
rect 6113 3893 6127 3907
rect 5993 3813 6007 3827
rect 6153 3993 6167 4007
rect 6053 3853 6067 3867
rect 6093 3816 6107 3830
rect 5993 3770 6007 3784
rect 6033 3770 6047 3784
rect 6073 3753 6087 3767
rect 6113 3733 6127 3747
rect 5993 3713 6007 3727
rect 6073 3713 6087 3727
rect 6053 3613 6067 3627
rect 5993 3593 6007 3607
rect 6013 3533 6027 3547
rect 5993 3513 6007 3527
rect 6073 3593 6087 3607
rect 5973 3353 5987 3367
rect 6093 3473 6107 3487
rect 6073 3393 6087 3407
rect 6093 3373 6107 3387
rect 6053 3333 6067 3347
rect 6033 3313 6047 3327
rect 5993 3296 6007 3310
rect 5973 3250 5987 3264
rect 6053 3233 6067 3247
rect 6013 3213 6027 3227
rect 5973 3153 5987 3167
rect 6013 3133 6027 3147
rect 5973 3093 5987 3107
rect 6093 3033 6107 3047
rect 5953 2913 5967 2927
rect 5933 2813 5947 2827
rect 5913 2573 5927 2587
rect 5793 2453 5807 2467
rect 5933 2513 5947 2527
rect 5873 2430 5887 2444
rect 5913 2430 5927 2444
rect 5833 2373 5847 2387
rect 5873 2373 5887 2387
rect 5793 2293 5807 2307
rect 5753 2273 5767 2287
rect 5773 2253 5787 2267
rect 5833 2256 5847 2270
rect 5753 2173 5767 2187
rect 5853 1993 5867 2007
rect 5693 1773 5707 1787
rect 5693 1736 5707 1750
rect 5413 1690 5427 1704
rect 5593 1690 5607 1704
rect 5633 1690 5647 1704
rect 5673 1690 5687 1704
rect 5713 1690 5727 1704
rect 5373 1593 5387 1607
rect 5453 1513 5467 1527
rect 5313 1493 5327 1507
rect 5333 1473 5347 1487
rect 5313 1390 5327 1404
rect 5313 1273 5327 1287
rect 5613 1473 5627 1487
rect 5573 1436 5587 1450
rect 5733 1433 5747 1447
rect 5553 1333 5567 1347
rect 5533 1253 5547 1267
rect 5513 1233 5527 1247
rect 5453 1213 5467 1227
rect 5333 1170 5347 1184
rect 5373 1170 5387 1184
rect 5333 1133 5347 1147
rect 5293 1093 5307 1107
rect 5233 993 5247 1007
rect 5253 916 5267 930
rect 5393 973 5407 987
rect 5313 870 5327 884
rect 5273 773 5287 787
rect 5393 773 5407 787
rect 5293 733 5307 747
rect 5273 673 5287 687
rect 5213 650 5227 664
rect 5273 553 5287 567
rect 5173 533 5187 547
rect 4553 313 4567 327
rect 4653 350 4667 364
rect 4713 373 4727 387
rect 4693 313 4707 327
rect 4533 293 4547 307
rect 4613 293 4627 307
rect 4753 370 4767 384
rect 4793 376 4807 390
rect 4953 376 4967 390
rect 5193 453 5207 467
rect 5073 370 5087 384
rect 5153 373 5167 387
rect 4713 273 4727 287
rect 4633 176 4647 190
rect 4493 153 4507 167
rect 4393 130 4407 144
rect 4073 93 4087 107
rect 4233 93 4247 107
rect 4433 93 4447 107
rect 5213 433 5227 447
rect 4953 176 4967 190
rect 5193 176 5207 190
rect 5693 1293 5707 1307
rect 5593 1233 5607 1247
rect 5533 1216 5547 1230
rect 5453 713 5467 727
rect 5513 1170 5527 1184
rect 5553 1170 5567 1184
rect 5593 1113 5607 1127
rect 5613 1073 5627 1087
rect 5593 1033 5607 1047
rect 5613 993 5627 1007
rect 5533 916 5547 930
rect 5573 916 5587 930
rect 5653 953 5667 967
rect 5533 813 5547 827
rect 5573 733 5587 747
rect 5413 513 5427 527
rect 5373 396 5387 410
rect 5293 350 5307 364
rect 5333 350 5347 364
rect 5553 393 5567 407
rect 5553 293 5567 307
rect 5413 176 5427 190
rect 5473 173 5487 187
rect 4753 53 4767 67
rect 5433 130 5447 144
rect 5513 173 5527 187
rect 5513 93 5527 107
rect 5633 870 5647 884
rect 5633 697 5647 711
rect 5733 1153 5747 1167
rect 5773 1953 5787 1967
rect 5793 1773 5807 1787
rect 5773 1653 5787 1667
rect 5773 1433 5787 1447
rect 5833 1736 5847 1750
rect 5833 1553 5847 1567
rect 5973 2776 5987 2790
rect 6033 2950 6047 2964
rect 6093 2950 6107 2964
rect 6113 2913 6127 2927
rect 6173 3473 6187 3487
rect 6253 4530 6267 4544
rect 6273 4453 6287 4467
rect 6233 4413 6247 4427
rect 6213 4213 6227 4227
rect 6213 4036 6227 4050
rect 6213 3873 6227 3887
rect 6213 3793 6227 3807
rect 6213 3653 6227 3667
rect 6253 4393 6267 4407
rect 6273 4373 6287 4387
rect 6253 4352 6267 4366
rect 6313 5273 6327 5287
rect 6333 5153 6347 5167
rect 6333 4953 6347 4967
rect 6573 5553 6587 5567
rect 6553 5533 6567 5547
rect 6433 5473 6447 5487
rect 6453 5330 6467 5344
rect 6513 5076 6527 5090
rect 6373 4893 6387 4907
rect 6313 4813 6327 4827
rect 6393 4810 6407 4824
rect 6433 4753 6447 4767
rect 6473 4753 6487 4767
rect 6333 4713 6347 4727
rect 6833 6453 6847 6467
rect 7033 6616 7047 6630
rect 7173 6613 7187 6627
rect 6973 6416 6987 6430
rect 7173 6413 7187 6427
rect 7213 6833 7227 6847
rect 7273 6753 7287 6767
rect 7333 6893 7347 6907
rect 7213 6653 7227 6667
rect 7213 6613 7227 6627
rect 7293 6610 7307 6624
rect 7233 6513 7247 6527
rect 7293 6453 7307 6467
rect 7253 6416 7267 6430
rect 6913 6253 6927 6267
rect 6873 6233 6887 6247
rect 6793 6193 6807 6207
rect 6713 6116 6727 6130
rect 6753 6116 6767 6130
rect 6813 6116 6827 6130
rect 6733 6070 6747 6084
rect 6813 6073 6827 6087
rect 6693 6033 6707 6047
rect 6673 5833 6687 5847
rect 6773 5913 6787 5927
rect 6813 5896 6827 5910
rect 6713 5850 6727 5864
rect 6753 5850 6767 5864
rect 6753 5829 6767 5843
rect 6733 5773 6747 5787
rect 6713 5753 6727 5767
rect 6793 5773 6807 5787
rect 6753 5753 6767 5767
rect 6733 5733 6747 5747
rect 6693 5693 6707 5707
rect 6673 5596 6687 5610
rect 6573 5433 6587 5447
rect 6633 5433 6647 5447
rect 6613 5376 6627 5390
rect 6653 5376 6667 5390
rect 6833 5596 6847 5610
rect 6753 5553 6767 5567
rect 6813 5533 6827 5547
rect 6793 5513 6807 5527
rect 6773 5473 6787 5487
rect 7033 6373 7047 6387
rect 6933 6193 6947 6207
rect 6913 6153 6927 6167
rect 7013 6333 7027 6347
rect 7173 6370 7187 6384
rect 7233 6370 7247 6384
rect 7273 6370 7287 6384
rect 7113 6253 7127 6267
rect 7033 6233 7047 6247
rect 7013 6153 7027 6167
rect 7053 6116 7067 6130
rect 7033 6070 7047 6084
rect 7413 7133 7427 7147
rect 7393 6973 7407 6987
rect 7373 6853 7387 6867
rect 7393 6833 7407 6847
rect 7353 6753 7367 6767
rect 7333 6573 7347 6587
rect 7373 6713 7387 6727
rect 7393 6673 7407 6687
rect 7373 6610 7387 6624
rect 7353 6553 7367 6567
rect 7333 6473 7347 6487
rect 7173 6173 7187 6187
rect 7313 6173 7327 6187
rect 6973 6033 6987 6047
rect 7073 6033 7087 6047
rect 6933 5993 6947 6007
rect 7013 5896 7027 5910
rect 7153 6013 7167 6027
rect 7093 5850 7107 5864
rect 7133 5850 7147 5864
rect 7013 5713 7027 5727
rect 7053 5713 7067 5727
rect 7113 5693 7127 5707
rect 6893 5633 6907 5647
rect 6893 5533 6907 5547
rect 6913 5377 6927 5391
rect 6953 5377 6967 5391
rect 7013 5377 7027 5391
rect 6713 5330 6727 5344
rect 6753 5330 6767 5344
rect 6793 5333 6807 5347
rect 6673 5273 6687 5287
rect 6653 5133 6667 5147
rect 6733 5113 6747 5127
rect 6613 5073 6627 5087
rect 6653 5073 6667 5087
rect 6613 4856 6627 4870
rect 6693 4893 6707 4907
rect 6573 4813 6587 4827
rect 6633 4810 6647 4824
rect 6553 4673 6567 4687
rect 6433 4633 6447 4647
rect 6653 4613 6667 4627
rect 6313 4573 6327 4587
rect 6613 4576 6627 4590
rect 6453 4536 6467 4550
rect 6573 4530 6587 4544
rect 6313 4493 6327 4507
rect 6633 4493 6647 4507
rect 6533 4433 6547 4447
rect 6433 4393 6447 4407
rect 6293 4353 6307 4367
rect 6313 4273 6327 4287
rect 6373 4273 6387 4287
rect 6353 4213 6367 4227
rect 6333 4193 6347 4207
rect 6273 4036 6287 4050
rect 6293 3990 6307 4004
rect 6293 3953 6307 3967
rect 6233 3513 6247 3527
rect 6193 3293 6207 3307
rect 6293 3816 6307 3830
rect 6273 3713 6287 3727
rect 6273 3633 6287 3647
rect 6453 4373 6467 4387
rect 6393 4253 6407 4267
rect 6433 4253 6447 4267
rect 6373 3973 6387 3987
rect 6353 3953 6367 3967
rect 6473 4336 6487 4350
rect 6513 4336 6527 4350
rect 6493 4233 6507 4247
rect 6473 4213 6487 4227
rect 6473 4173 6487 4187
rect 6393 3933 6407 3947
rect 6373 3816 6387 3830
rect 6453 3816 6467 3830
rect 6353 3770 6367 3784
rect 6333 3693 6347 3707
rect 6373 3693 6387 3707
rect 6293 3573 6307 3587
rect 6393 3633 6407 3647
rect 6293 3533 6307 3547
rect 6353 3513 6367 3527
rect 6233 3233 6247 3247
rect 6193 3153 6207 3167
rect 6233 3153 6247 3167
rect 6153 2953 6167 2967
rect 6153 2833 6167 2847
rect 6053 2776 6067 2790
rect 6093 2776 6107 2790
rect 6073 2730 6087 2744
rect 6173 2730 6187 2744
rect 5993 2693 6007 2707
rect 6113 2693 6127 2707
rect 5973 2673 5987 2687
rect 5973 2293 5987 2307
rect 5953 2213 5967 2227
rect 5933 2033 5947 2047
rect 6013 2593 6027 2607
rect 6173 2593 6187 2607
rect 6013 2553 6027 2567
rect 6133 2553 6147 2567
rect 6093 2476 6107 2490
rect 6273 3113 6287 3127
rect 6212 2773 6226 2787
rect 6233 2773 6247 2787
rect 6193 2493 6207 2507
rect 5993 1993 6007 2007
rect 5933 1956 5947 1970
rect 5913 1893 5927 1907
rect 5953 1773 5967 1787
rect 5893 1733 5907 1747
rect 5953 1736 5967 1750
rect 5933 1690 5947 1704
rect 5933 1653 5947 1667
rect 5893 1593 5907 1607
rect 6133 2373 6147 2387
rect 6113 2313 6127 2327
rect 6053 2256 6067 2270
rect 6053 2033 6067 2047
rect 6033 2013 6047 2027
rect 6033 1853 6047 1867
rect 5973 1553 5987 1567
rect 5873 1513 5887 1527
rect 5853 1456 5867 1470
rect 5933 1453 5947 1467
rect 5813 1433 5827 1447
rect 5853 1435 5867 1449
rect 5913 1433 5927 1447
rect 5793 1390 5807 1404
rect 5833 1390 5847 1404
rect 5813 1216 5827 1230
rect 5853 1216 5867 1230
rect 5793 1153 5807 1167
rect 5833 1153 5847 1167
rect 5873 1153 5887 1167
rect 5913 1153 5927 1167
rect 5773 870 5787 884
rect 5753 753 5767 767
rect 5773 693 5787 707
rect 5593 653 5607 667
rect 5613 453 5627 467
rect 5713 393 5727 407
rect 5653 350 5667 364
rect 5713 350 5727 364
rect 5633 313 5647 327
rect 5673 213 5687 227
rect 5753 313 5767 327
rect 5733 193 5747 207
rect 5713 176 5727 190
rect 5633 133 5647 147
rect 5893 1113 5907 1127
rect 5813 1013 5827 1027
rect 5893 993 5907 1007
rect 5813 870 5827 884
rect 5853 870 5867 884
rect 5913 773 5927 787
rect 5893 753 5907 767
rect 5833 493 5847 507
rect 5813 373 5827 387
rect 5813 293 5827 307
rect 5913 613 5927 627
rect 6113 2213 6127 2227
rect 6093 1910 6107 1924
rect 6133 1633 6147 1647
rect 6233 2653 6247 2667
rect 6233 2430 6247 2444
rect 6213 2252 6227 2266
rect 6273 2813 6287 2827
rect 6293 2653 6307 2667
rect 6273 2253 6287 2267
rect 6273 2073 6287 2087
rect 6253 1956 6267 1970
rect 6193 1910 6207 1924
rect 6233 1853 6247 1867
rect 6193 1736 6207 1750
rect 6273 1733 6287 1747
rect 6173 1693 6187 1707
rect 6153 1593 6167 1607
rect 6113 1573 6127 1587
rect 6093 1453 6107 1467
rect 6133 1453 6147 1467
rect 5993 1253 6007 1267
rect 6013 1213 6027 1227
rect 5993 953 6007 967
rect 6013 916 6027 930
rect 6073 1390 6087 1404
rect 6153 1393 6167 1407
rect 6213 1690 6227 1704
rect 6233 1633 6247 1647
rect 6213 1353 6227 1367
rect 6173 1333 6187 1347
rect 6093 1273 6107 1287
rect 6133 1273 6147 1287
rect 6133 1216 6147 1230
rect 6213 1073 6227 1087
rect 6153 1033 6167 1047
rect 6193 1033 6207 1047
rect 6113 993 6127 1007
rect 6153 993 6167 1007
rect 6113 916 6127 930
rect 6133 870 6147 884
rect 6193 873 6207 887
rect 6033 833 6047 847
rect 6353 3213 6367 3227
rect 6433 3733 6447 3747
rect 6353 2933 6367 2947
rect 6373 2913 6387 2927
rect 6333 2893 6347 2907
rect 6333 2813 6347 2827
rect 6413 3473 6427 3487
rect 6453 3653 6467 3667
rect 6573 4290 6587 4304
rect 6573 4253 6587 4267
rect 6533 4193 6547 4207
rect 6513 4093 6527 4107
rect 6493 4073 6507 4087
rect 6633 4192 6647 4206
rect 6613 4073 6627 4087
rect 6533 3990 6547 4004
rect 6513 3973 6527 3987
rect 6493 3953 6507 3967
rect 6433 2913 6447 2927
rect 6353 2730 6367 2744
rect 6393 2673 6407 2687
rect 6613 3993 6627 4007
rect 6633 3816 6647 3830
rect 6673 4533 6687 4547
rect 6673 4290 6687 4304
rect 6573 3793 6587 3807
rect 6553 3593 6567 3607
rect 6613 3770 6627 3784
rect 6713 4856 6727 4870
rect 6793 5076 6807 5090
rect 6753 5013 6767 5027
rect 6733 4653 6747 4667
rect 6713 4576 6727 4590
rect 6693 4032 6707 4046
rect 6813 4993 6827 5007
rect 6773 4953 6787 4967
rect 7073 5373 7087 5387
rect 7093 5377 7107 5391
rect 6773 4913 6787 4927
rect 6913 4913 6927 4927
rect 6813 4856 6827 4870
rect 6853 4856 6867 4870
rect 6893 4856 6907 4870
rect 6813 4813 6827 4827
rect 6773 4453 6787 4467
rect 6812 4673 6826 4687
rect 6833 4673 6847 4687
rect 6993 5331 7007 5345
rect 7053 5313 7067 5327
rect 7093 5293 7107 5307
rect 7033 5076 7047 5090
rect 7073 5076 7087 5090
rect 7013 4993 7027 5007
rect 6973 4856 6987 4870
rect 6933 4633 6947 4647
rect 6873 4613 6887 4627
rect 7033 4933 7047 4947
rect 7013 4810 7027 4824
rect 6833 4555 6847 4569
rect 6933 4509 6947 4523
rect 6813 4493 6827 4507
rect 6933 4453 6947 4467
rect 6833 4336 6847 4350
rect 6873 4336 6887 4350
rect 6913 4336 6927 4350
rect 6753 4213 6767 4227
rect 6773 4193 6787 4207
rect 6913 4293 6927 4307
rect 6853 4253 6867 4267
rect 6813 4233 6827 4247
rect 6873 4233 6887 4247
rect 6853 4193 6867 4207
rect 6793 4133 6807 4147
rect 6793 4073 6807 4087
rect 6753 4036 6767 4050
rect 6713 3953 6727 3967
rect 6693 3816 6707 3830
rect 6693 3733 6707 3747
rect 6673 3713 6687 3727
rect 6713 3713 6727 3727
rect 6653 3693 6667 3707
rect 6813 3990 6827 4004
rect 6773 3933 6787 3947
rect 6913 4213 6927 4227
rect 6893 4173 6907 4187
rect 6913 3893 6927 3907
rect 6793 3833 6807 3847
rect 6853 3833 6867 3847
rect 6753 3813 6767 3827
rect 6733 3673 6747 3687
rect 6573 3553 6587 3567
rect 6713 3533 6727 3547
rect 6593 3516 6607 3530
rect 6673 3513 6687 3527
rect 6613 3470 6627 3484
rect 6573 3433 6587 3447
rect 6513 3296 6527 3310
rect 6553 3296 6567 3310
rect 6613 3296 6627 3310
rect 6653 3293 6667 3307
rect 6473 3233 6487 3247
rect 6533 3250 6547 3264
rect 6493 3213 6507 3227
rect 6553 3213 6567 3227
rect 6513 3193 6527 3207
rect 6493 3173 6507 3187
rect 6453 2773 6467 2787
rect 6433 2633 6447 2647
rect 6413 2613 6427 2627
rect 6353 2553 6367 2567
rect 6413 2533 6427 2547
rect 6413 2493 6427 2507
rect 6393 2430 6407 2444
rect 6313 2373 6327 2387
rect 6353 2373 6367 2387
rect 6373 2333 6387 2347
rect 6333 2256 6347 2270
rect 6353 2193 6367 2207
rect 6333 2153 6347 2167
rect 6393 2153 6407 2167
rect 6353 2073 6367 2087
rect 6453 2033 6467 2047
rect 6413 1953 6427 1967
rect 6533 2933 6547 2947
rect 6513 2653 6527 2667
rect 6513 2513 6527 2527
rect 6513 2453 6527 2467
rect 6593 2950 6607 2964
rect 6673 3250 6687 3264
rect 6713 3213 6727 3227
rect 6873 3816 6887 3830
rect 6813 3770 6827 3784
rect 6853 3770 6867 3784
rect 6833 3693 6847 3707
rect 6893 3673 6907 3687
rect 6833 3653 6847 3667
rect 6793 3516 6807 3530
rect 6913 3473 6927 3487
rect 6853 3432 6867 3446
rect 6753 3293 6767 3307
rect 6813 3296 6827 3310
rect 6793 3253 6807 3267
rect 6773 3173 6787 3187
rect 6733 3073 6747 3087
rect 6733 2996 6747 3010
rect 6833 3193 6847 3207
rect 6833 3033 6847 3047
rect 6713 2950 6727 2964
rect 6653 2853 6667 2867
rect 6633 2776 6647 2790
rect 6553 2693 6567 2707
rect 6653 2730 6667 2744
rect 6653 2713 6667 2727
rect 6553 2672 6567 2686
rect 6613 2673 6627 2687
rect 6533 2393 6547 2407
rect 6633 2476 6647 2490
rect 6733 2473 6747 2487
rect 6693 2413 6707 2427
rect 6653 2373 6667 2387
rect 6613 2333 6627 2347
rect 6713 2333 6727 2347
rect 6653 2256 6667 2270
rect 6693 2253 6707 2267
rect 6513 2153 6527 2167
rect 6373 1853 6387 1867
rect 6373 1793 6387 1807
rect 6313 1693 6327 1707
rect 6313 1653 6327 1667
rect 6353 1573 6367 1587
rect 6293 1293 6307 1307
rect 6313 1213 6327 1227
rect 6473 1910 6487 1924
rect 6433 1813 6447 1827
rect 6413 1233 6427 1247
rect 6373 1216 6387 1230
rect 6553 1910 6567 1924
rect 6453 1773 6467 1787
rect 6513 1773 6527 1787
rect 6333 1173 6347 1187
rect 6393 1170 6407 1184
rect 6313 1013 6327 1027
rect 6273 973 6287 987
rect 6313 913 6327 927
rect 6393 916 6407 930
rect 6253 893 6267 907
rect 6253 853 6267 867
rect 6293 773 6307 787
rect 6233 733 6247 747
rect 6293 733 6307 747
rect 6273 696 6287 710
rect 5893 396 5907 410
rect 5933 395 5947 409
rect 5873 313 5887 327
rect 5913 313 5927 327
rect 6253 650 6267 664
rect 6193 633 6207 647
rect 6273 573 6287 587
rect 6513 1736 6527 1750
rect 6593 2193 6607 2207
rect 6673 2153 6687 2167
rect 6613 2113 6627 2127
rect 6593 2033 6607 2047
rect 6593 1956 6607 1970
rect 6473 1053 6487 1067
rect 6453 873 6467 887
rect 6373 833 6387 847
rect 6613 1913 6627 1927
rect 6593 1633 6607 1647
rect 6553 1533 6567 1547
rect 6593 1513 6607 1527
rect 6593 1473 6607 1487
rect 6673 1613 6687 1627
rect 6633 1436 6647 1450
rect 6613 1390 6627 1404
rect 6653 1333 6667 1347
rect 6713 2173 6727 2187
rect 6833 2913 6847 2927
rect 6793 2853 6807 2867
rect 6773 2813 6787 2827
rect 6773 2430 6787 2444
rect 6753 2073 6767 2087
rect 6833 2653 6847 2667
rect 6813 2393 6827 2407
rect 6813 2313 6827 2327
rect 6873 3296 6887 3310
rect 6893 2993 6907 3007
rect 6893 2950 6907 2964
rect 6953 4293 6967 4307
rect 7053 4893 7067 4907
rect 7133 5013 7147 5027
rect 7193 6133 7207 6147
rect 7273 6053 7287 6067
rect 7213 5993 7227 6007
rect 7193 5773 7207 5787
rect 7193 5713 7207 5727
rect 7173 4933 7187 4947
rect 7273 5953 7287 5967
rect 7393 6052 7407 6066
rect 7313 5896 7327 5910
rect 7233 5813 7247 5827
rect 7213 5473 7227 5487
rect 7213 5173 7227 5187
rect 7213 5076 7227 5090
rect 7213 5033 7227 5047
rect 7213 4973 7227 4987
rect 7213 4873 7227 4887
rect 7033 4555 7047 4569
rect 7033 4413 7047 4427
rect 7093 4853 7107 4867
rect 7153 4856 7167 4870
rect 7073 4773 7087 4787
rect 7133 4810 7147 4824
rect 7173 4810 7187 4824
rect 7213 4810 7227 4824
rect 7093 4753 7107 4767
rect 7093 4732 7107 4746
rect 7093 4593 7107 4607
rect 7133 4593 7147 4607
rect 7353 5850 7367 5864
rect 7373 5793 7387 5807
rect 7353 5753 7367 5767
rect 7433 7113 7447 7127
rect 7453 7053 7467 7067
rect 7453 6993 7467 7007
rect 7533 7553 7547 7567
rect 7573 7553 7587 7567
rect 7553 7533 7567 7547
rect 7533 7513 7547 7527
rect 7513 7410 7527 7424
rect 7632 7456 7646 7470
rect 7673 7893 7687 7907
rect 7993 7950 8007 7964
rect 8133 8033 8147 8047
rect 8173 8213 8187 8227
rect 8173 8073 8187 8087
rect 8133 7950 8147 7964
rect 8173 7953 8187 7967
rect 7833 7833 7847 7847
rect 7953 7833 7967 7847
rect 7973 7713 7987 7727
rect 7673 7693 7687 7707
rect 7953 7693 7967 7707
rect 7813 7656 7827 7670
rect 8153 7910 8167 7924
rect 8193 7913 8207 7927
rect 8153 7813 8167 7827
rect 8133 7713 8147 7727
rect 8073 7673 8087 7687
rect 7933 7650 7947 7664
rect 8053 7653 8067 7667
rect 7673 7613 7687 7627
rect 7733 7513 7747 7527
rect 7653 7453 7667 7467
rect 7673 7436 7687 7450
rect 7773 7453 7787 7467
rect 7553 7333 7567 7347
rect 7613 7313 7627 7327
rect 7573 7293 7587 7307
rect 7933 7430 7947 7444
rect 8073 7553 8087 7567
rect 8113 7513 8127 7527
rect 8113 7430 8127 7444
rect 8273 8333 8287 8347
rect 8353 8793 8367 8807
rect 8333 8393 8347 8407
rect 8373 8450 8387 8464
rect 8453 9533 8467 9547
rect 8493 9653 8507 9667
rect 8693 10233 8707 10247
rect 8633 10193 8647 10207
rect 8613 9693 8627 9707
rect 8593 9573 8607 9587
rect 8533 9553 8547 9567
rect 8573 9536 8587 9550
rect 8773 10893 8787 10907
rect 8773 10833 8787 10847
rect 8973 10953 8987 10967
rect 8793 10793 8807 10807
rect 8793 10750 8807 10764
rect 8833 10576 8847 10590
rect 8813 10513 8827 10527
rect 8913 10796 8927 10810
rect 8933 10673 8947 10687
rect 8913 10473 8927 10487
rect 8873 10273 8887 10287
rect 8893 10230 8907 10244
rect 8773 10193 8787 10207
rect 9133 11096 9147 11110
rect 9253 11093 9267 11107
rect 9053 11033 9067 11047
rect 9173 11033 9187 11047
rect 9153 10893 9167 10907
rect 9113 10813 9127 10827
rect 9293 11316 9307 11330
rect 9973 11873 9987 11887
rect 9493 11853 9507 11867
rect 10013 11833 10027 11847
rect 9613 11810 9627 11824
rect 9813 11816 9827 11830
rect 9473 11790 9487 11804
rect 9553 11793 9567 11807
rect 9513 11633 9527 11647
rect 9753 11616 9767 11630
rect 9493 11570 9507 11584
rect 9653 11553 9667 11567
rect 9493 11413 9507 11427
rect 9433 11373 9447 11387
rect 9453 11316 9467 11330
rect 9733 11533 9747 11547
rect 9813 11533 9827 11547
rect 9773 11493 9787 11507
rect 9773 11333 9787 11347
rect 9413 11270 9427 11284
rect 9513 11270 9527 11284
rect 9653 11270 9667 11284
rect 9733 11270 9747 11284
rect 9293 11253 9307 11267
rect 9473 11253 9487 11267
rect 9553 11133 9567 11147
rect 9453 11096 9467 11110
rect 9493 11096 9507 11110
rect 9433 11050 9447 11064
rect 9473 11033 9487 11047
rect 9273 10993 9287 11007
rect 9473 10953 9487 10967
rect 9253 10913 9267 10927
rect 9213 10833 9227 10847
rect 9413 10833 9427 10847
rect 9453 10833 9467 10847
rect 9433 10813 9447 10827
rect 9473 10813 9487 10827
rect 9553 11096 9567 11110
rect 9233 10750 9247 10764
rect 9453 10750 9467 10764
rect 9533 10753 9547 10767
rect 9173 10733 9187 10747
rect 9213 10733 9227 10747
rect 9073 10576 9087 10590
rect 9113 10576 9127 10590
rect 9093 10530 9107 10544
rect 9053 10473 9067 10487
rect 9153 10473 9167 10487
rect 9093 10373 9107 10387
rect 9033 10293 9047 10307
rect 8753 10113 8767 10127
rect 8893 10113 8907 10127
rect 8733 10056 8747 10070
rect 8773 10056 8787 10070
rect 8813 10056 8827 10070
rect 8713 9776 8727 9790
rect 8873 10053 8887 10067
rect 8773 9993 8787 10007
rect 8793 9913 8807 9927
rect 8833 9753 8847 9767
rect 8553 9490 8567 9504
rect 8493 9473 8507 9487
rect 8493 9236 8507 9250
rect 8473 9173 8487 9187
rect 8433 9033 8447 9047
rect 8453 9016 8467 9030
rect 8573 9236 8587 9250
rect 8633 9493 8647 9507
rect 8593 9093 8607 9107
rect 8593 9053 8607 9067
rect 8553 9016 8567 9030
rect 8773 9633 8787 9647
rect 8913 10093 8927 10107
rect 8893 9913 8907 9927
rect 8873 9736 8887 9750
rect 8833 9653 8847 9667
rect 8853 9593 8867 9607
rect 8813 9573 8827 9587
rect 8793 9533 8807 9547
rect 8893 9573 8907 9587
rect 8773 9513 8787 9527
rect 8753 9393 8767 9407
rect 8653 9273 8667 9287
rect 8733 9273 8747 9287
rect 8613 9033 8627 9047
rect 8893 9453 8907 9467
rect 9093 10230 9107 10244
rect 9133 10230 9147 10244
rect 9173 10230 9187 10244
rect 9093 10093 9107 10107
rect 9093 10056 9107 10070
rect 9133 10056 9147 10070
rect 9033 10010 9047 10024
rect 9073 10010 9087 10024
rect 9113 9913 9127 9927
rect 9053 9813 9067 9827
rect 9013 9756 9027 9770
rect 9153 9756 9167 9770
rect 8993 9713 9007 9727
rect 8953 9553 8967 9567
rect 8693 9236 8707 9250
rect 8733 9236 8747 9250
rect 8673 9093 8687 9107
rect 8653 9013 8667 9027
rect 8613 8970 8627 8984
rect 8633 8873 8647 8887
rect 8693 8933 8707 8947
rect 8633 8813 8647 8827
rect 8533 8793 8547 8807
rect 8453 8753 8467 8767
rect 8513 8753 8527 8767
rect 8593 8753 8607 8767
rect 8433 8673 8447 8687
rect 8553 8670 8567 8684
rect 8593 8673 8607 8687
rect 8513 8573 8527 8587
rect 8513 8533 8527 8547
rect 8733 9093 8747 9107
rect 8733 8970 8747 8984
rect 8653 8633 8667 8647
rect 8613 8613 8627 8627
rect 8613 8553 8627 8567
rect 8553 8513 8567 8527
rect 8833 9233 8847 9247
rect 8773 9053 8787 9067
rect 8813 9053 8827 9067
rect 8793 8996 8807 9010
rect 8773 8873 8787 8887
rect 8813 8893 8827 8907
rect 8793 8853 8807 8867
rect 8753 8773 8767 8787
rect 8873 9073 8887 9087
rect 8973 9533 8987 9547
rect 8973 9313 8987 9327
rect 9033 9710 9047 9724
rect 9033 9613 9047 9627
rect 9093 9536 9107 9550
rect 9033 9490 9047 9504
rect 9113 9490 9127 9504
rect 9193 10013 9207 10027
rect 9173 9573 9187 9587
rect 9173 9493 9187 9507
rect 9193 9413 9207 9427
rect 9073 9393 9087 9407
rect 9153 9393 9167 9407
rect 9013 9353 9027 9367
rect 9053 9273 9067 9287
rect 9093 9273 9107 9287
rect 9033 9190 9047 9204
rect 8953 9133 8967 9147
rect 9053 9133 9067 9147
rect 9013 9013 9027 9027
rect 8953 8996 8967 9010
rect 9033 8933 9047 8947
rect 8893 8913 8907 8927
rect 8853 8833 8867 8847
rect 8773 8716 8787 8730
rect 8693 8670 8707 8684
rect 8753 8670 8767 8684
rect 8493 8450 8507 8464
rect 8673 8453 8687 8467
rect 8793 8633 8807 8647
rect 8773 8553 8787 8567
rect 8813 8513 8827 8527
rect 8413 8353 8427 8367
rect 8653 8353 8667 8367
rect 8673 8333 8687 8347
rect 8393 8313 8407 8327
rect 8653 8313 8667 8327
rect 8373 8253 8387 8267
rect 8353 8233 8367 8247
rect 8417 8213 8431 8227
rect 8693 8213 8707 8227
rect 8313 8196 8327 8210
rect 8373 8173 8387 8187
rect 8293 8150 8307 8164
rect 8333 8150 8347 8164
rect 8253 8093 8267 8107
rect 8233 8013 8247 8027
rect 8433 8170 8447 8184
rect 8553 8176 8567 8190
rect 8733 8450 8747 8464
rect 8813 8413 8827 8427
rect 8793 8213 8807 8227
rect 8713 8173 8727 8187
rect 8433 8113 8447 8127
rect 8713 8113 8727 8127
rect 8413 8033 8427 8047
rect 8273 7953 8287 7967
rect 8233 7833 8247 7847
rect 8233 7773 8247 7787
rect 8213 7733 8227 7747
rect 8193 7676 8207 7690
rect 8153 7613 8167 7627
rect 8093 7353 8107 7367
rect 8133 7353 8147 7367
rect 8113 7313 8127 7327
rect 7953 7293 7967 7307
rect 7773 7273 7787 7287
rect 7833 7273 7847 7287
rect 7493 7173 7507 7187
rect 7793 7176 7807 7190
rect 7633 7136 7647 7150
rect 7732 7136 7746 7150
rect 7493 7113 7507 7127
rect 7753 7130 7767 7144
rect 7733 7093 7747 7107
rect 7653 7033 7667 7047
rect 7533 6936 7547 6950
rect 7593 6916 7607 6930
rect 7893 7213 7907 7227
rect 7893 7176 7907 7190
rect 7853 7133 7867 7147
rect 7853 7093 7867 7107
rect 8133 7293 8147 7307
rect 8073 7253 8087 7267
rect 8113 7253 8127 7267
rect 8033 7156 8047 7170
rect 8073 7156 8087 7170
rect 7993 7113 8007 7127
rect 8053 7110 8067 7124
rect 7973 7093 7987 7107
rect 7913 7053 7927 7067
rect 7953 7053 7967 7067
rect 7893 7033 7907 7047
rect 7693 7013 7707 7027
rect 7833 7013 7847 7027
rect 7473 6893 7487 6907
rect 8073 7073 8087 7087
rect 8053 7053 8067 7067
rect 8033 7033 8047 7047
rect 7993 6953 8007 6967
rect 7973 6933 7987 6947
rect 7853 6910 7867 6924
rect 8033 6913 8047 6927
rect 7553 6873 7567 6887
rect 7693 6873 7707 6887
rect 7453 6773 7467 6787
rect 8013 6870 8027 6884
rect 7493 6733 7507 6747
rect 7473 6573 7487 6587
rect 7633 6813 7647 6827
rect 7613 6793 7627 6807
rect 7573 6753 7587 6767
rect 7573 6636 7587 6650
rect 7513 6593 7527 6607
rect 7613 6573 7627 6587
rect 7553 6493 7567 6507
rect 7493 6473 7507 6487
rect 7453 6433 7467 6447
rect 7433 6333 7447 6347
rect 7433 6273 7447 6287
rect 7433 5853 7447 5867
rect 7412 5813 7426 5827
rect 7433 5813 7447 5827
rect 7413 5753 7427 5767
rect 7372 5713 7386 5727
rect 7393 5713 7407 5727
rect 7413 5673 7427 5687
rect 7253 5653 7267 5667
rect 7353 5653 7367 5667
rect 7313 5596 7327 5610
rect 7353 5533 7367 5547
rect 7353 5433 7367 5447
rect 7313 5376 7327 5390
rect 7313 5293 7327 5307
rect 7373 5273 7387 5287
rect 7353 5233 7367 5247
rect 7273 5193 7287 5207
rect 7293 5133 7307 5147
rect 7353 5113 7367 5127
rect 7313 5030 7327 5044
rect 7273 4993 7287 5007
rect 7253 4933 7267 4947
rect 7093 4513 7107 4527
rect 7193 4510 7207 4524
rect 7233 4513 7247 4527
rect 7273 4713 7287 4727
rect 7073 4393 7087 4407
rect 7133 4393 7147 4407
rect 7093 4290 7107 4304
rect 7133 4273 7147 4287
rect 7113 4253 7127 4267
rect 7013 4173 7027 4187
rect 7073 4133 7087 4147
rect 7113 4133 7127 4147
rect 6993 4093 7007 4107
rect 7073 4053 7087 4067
rect 7053 4036 7067 4050
rect 7093 4036 7107 4050
rect 6972 3993 6986 4007
rect 6993 3993 7007 4007
rect 6993 3953 7007 3967
rect 6953 3473 6967 3487
rect 6932 3433 6946 3447
rect 6953 3433 6967 3447
rect 6973 3373 6987 3387
rect 7073 3990 7087 4004
rect 7033 3893 7047 3907
rect 7013 3693 7027 3707
rect 7013 3633 7027 3647
rect 7113 3873 7127 3887
rect 7053 3833 7067 3847
rect 7153 4073 7167 4087
rect 7193 4393 7207 4407
rect 7313 4810 7327 4824
rect 7293 4273 7307 4287
rect 7393 5233 7407 5247
rect 7393 4933 7407 4947
rect 7473 6416 7487 6430
rect 7553 6416 7567 6430
rect 7453 5313 7467 5327
rect 7453 5133 7467 5147
rect 7453 5030 7467 5044
rect 7513 6370 7527 6384
rect 7533 6133 7547 6147
rect 7533 6116 7547 6130
rect 7553 6053 7567 6067
rect 7513 6013 7527 6027
rect 7653 6793 7667 6807
rect 7673 6773 7687 6787
rect 7653 6713 7667 6727
rect 7753 6733 7767 6747
rect 7673 6673 7687 6687
rect 7653 6633 7667 6647
rect 7693 6636 7707 6650
rect 7633 6553 7647 6567
rect 7633 6513 7647 6527
rect 7633 6453 7647 6467
rect 7633 6416 7647 6430
rect 7633 6253 7647 6267
rect 7713 6573 7727 6587
rect 7693 6493 7707 6507
rect 7673 6373 7687 6387
rect 7653 6112 7667 6126
rect 7613 5973 7627 5987
rect 7513 5896 7527 5910
rect 7593 5896 7607 5910
rect 7613 5850 7627 5864
rect 7613 5653 7627 5667
rect 7553 5613 7567 5627
rect 7693 5773 7707 5787
rect 7673 5733 7687 5747
rect 7673 5593 7687 5607
rect 7653 5493 7667 5507
rect 7573 5413 7587 5427
rect 7693 5433 7707 5447
rect 7673 5393 7687 5407
rect 7613 5376 7627 5390
rect 7513 5313 7527 5327
rect 7573 5293 7587 5307
rect 7633 5293 7647 5307
rect 7693 5273 7707 5287
rect 7633 5253 7647 5267
rect 7593 5173 7607 5187
rect 7433 4953 7447 4967
rect 7493 4953 7507 4967
rect 7453 4913 7467 4927
rect 7413 4873 7427 4887
rect 7493 4873 7507 4887
rect 7433 4810 7447 4824
rect 7473 4753 7487 4767
rect 7493 4693 7507 4707
rect 7493 4613 7507 4627
rect 7433 4573 7447 4587
rect 7473 4573 7487 4587
rect 7373 4473 7387 4487
rect 7433 4433 7447 4447
rect 7413 4413 7427 4427
rect 7393 4353 7407 4367
rect 7353 4336 7367 4350
rect 7313 4253 7327 4267
rect 7233 4233 7247 4247
rect 7273 4233 7287 4247
rect 7253 4173 7267 4187
rect 7193 4113 7207 4127
rect 7233 4053 7247 4067
rect 7193 4013 7207 4027
rect 7173 3953 7187 3967
rect 7153 3933 7167 3947
rect 7153 3912 7167 3926
rect 7193 3893 7207 3907
rect 7153 3853 7167 3867
rect 7133 3833 7147 3847
rect 7153 3816 7167 3830
rect 7133 3770 7147 3784
rect 7193 3773 7207 3787
rect 7113 3713 7127 3727
rect 7073 3573 7087 3587
rect 7053 3533 7067 3547
rect 7213 3713 7227 3727
rect 7193 3613 7207 3627
rect 7113 3533 7127 3547
rect 7173 3533 7187 3547
rect 7133 3470 7147 3484
rect 7093 3433 7107 3447
rect 7013 3373 7027 3387
rect 7153 3353 7167 3367
rect 7033 3333 7047 3347
rect 7073 3296 7087 3310
rect 7113 3296 7127 3310
rect 6993 3253 7007 3267
rect 7093 3253 7107 3267
rect 7053 3213 7067 3227
rect 6973 3173 6987 3187
rect 7033 3113 7047 3127
rect 7013 3033 7027 3047
rect 6973 2996 6987 3010
rect 6953 2950 6967 2964
rect 6993 2933 7007 2947
rect 6913 2775 6927 2789
rect 6893 2713 6907 2727
rect 7033 2693 7047 2707
rect 7013 2593 7027 2607
rect 6993 2573 7007 2587
rect 7033 2573 7047 2587
rect 6993 2533 7007 2547
rect 6953 2476 6967 2490
rect 6913 2430 6927 2444
rect 6933 2393 6947 2407
rect 6913 2256 6927 2270
rect 6853 2213 6867 2227
rect 6833 2113 6847 2127
rect 6813 2093 6827 2107
rect 6793 2053 6807 2067
rect 6873 2053 6887 2067
rect 6753 2033 6767 2047
rect 6853 2013 6867 2027
rect 6793 1993 6807 2007
rect 6793 1956 6807 1970
rect 6773 1910 6787 1924
rect 6833 1913 6847 1927
rect 6813 1893 6827 1907
rect 6833 1853 6847 1867
rect 6853 1813 6867 1827
rect 6753 1736 6767 1750
rect 6793 1736 6807 1750
rect 6693 1273 6707 1287
rect 6593 1233 6607 1247
rect 6573 1216 6587 1230
rect 6513 793 6527 807
rect 6693 1216 6707 1230
rect 6693 1153 6707 1167
rect 6633 1133 6647 1147
rect 6673 1133 6687 1147
rect 6593 916 6607 930
rect 6633 916 6647 930
rect 6713 1093 6727 1107
rect 6553 833 6567 847
rect 6533 773 6547 787
rect 6473 650 6487 664
rect 6533 650 6547 664
rect 6573 633 6587 647
rect 6673 793 6687 807
rect 6653 673 6667 687
rect 6633 613 6647 627
rect 6453 513 6467 527
rect 6853 1693 6867 1707
rect 6773 1653 6787 1667
rect 6753 1613 6767 1627
rect 6913 2213 6927 2227
rect 6953 2113 6967 2127
rect 6913 1853 6927 1867
rect 6933 1833 6947 1847
rect 6893 1736 6907 1750
rect 6853 1473 6867 1487
rect 6813 1113 6827 1127
rect 6753 1093 6767 1107
rect 6733 1053 6747 1067
rect 6773 973 6787 987
rect 6813 913 6827 927
rect 6733 853 6747 867
rect 6773 853 6787 867
rect 6753 773 6767 787
rect 6813 733 6827 747
rect 6933 1690 6947 1704
rect 6953 1633 6967 1647
rect 6913 1553 6927 1567
rect 7013 2513 7027 2527
rect 7033 2333 7047 2347
rect 6993 1953 7007 1967
rect 7093 3133 7107 3147
rect 7133 3133 7147 3147
rect 7113 3093 7127 3107
rect 7073 2973 7087 2987
rect 7153 2933 7167 2947
rect 7073 2893 7087 2907
rect 7193 3213 7207 3227
rect 7233 3633 7247 3647
rect 7233 3213 7247 3227
rect 7233 3113 7247 3127
rect 7373 4253 7387 4267
rect 7413 4253 7427 4267
rect 7353 4073 7367 4087
rect 7333 4036 7347 4050
rect 7313 3990 7327 4004
rect 7333 3953 7347 3967
rect 7273 3893 7287 3907
rect 7413 4133 7427 4147
rect 7393 4033 7407 4047
rect 7393 3990 7407 4004
rect 7513 4473 7527 4487
rect 7493 4353 7507 4367
rect 7473 4336 7487 4350
rect 7493 4213 7507 4227
rect 7453 3993 7467 4007
rect 7433 3816 7447 3830
rect 7373 3773 7387 3787
rect 7453 3753 7467 3767
rect 7293 3713 7307 3727
rect 7413 3713 7427 3727
rect 7273 3633 7287 3647
rect 7273 3533 7287 3547
rect 7353 3533 7367 3547
rect 7413 3516 7427 3530
rect 7393 3433 7407 3447
rect 7393 3393 7407 3407
rect 7273 3333 7287 3347
rect 7333 3313 7347 3327
rect 7293 3296 7307 3310
rect 7313 3250 7327 3264
rect 7393 3250 7407 3264
rect 7253 3013 7267 3027
rect 7313 3013 7327 3027
rect 7173 2873 7187 2887
rect 7253 2933 7267 2947
rect 7273 2913 7287 2927
rect 7193 2833 7207 2847
rect 7233 2833 7247 2847
rect 7072 2773 7086 2787
rect 7093 2773 7107 2787
rect 7153 2776 7167 2790
rect 7193 2776 7207 2790
rect 7073 2733 7087 2747
rect 7133 2730 7147 2744
rect 7213 2730 7227 2744
rect 7173 2673 7187 2687
rect 7093 2653 7107 2667
rect 7073 2633 7087 2647
rect 7093 2553 7107 2567
rect 7133 2513 7147 2527
rect 7253 2776 7267 2790
rect 7233 2513 7247 2527
rect 7213 2476 7227 2490
rect 7133 2430 7147 2444
rect 7173 2430 7187 2444
rect 7253 2373 7267 2387
rect 7153 2313 7167 2327
rect 7113 2293 7127 2307
rect 7173 2256 7187 2270
rect 7153 2173 7167 2187
rect 7113 2113 7127 2127
rect 7093 2013 7107 2027
rect 7053 1833 7067 1847
rect 7013 1813 7027 1827
rect 7033 1690 7047 1704
rect 7133 2093 7147 2107
rect 7153 2033 7167 2047
rect 7133 1793 7147 1807
rect 7153 1773 7167 1787
rect 7093 1653 7107 1667
rect 7173 1653 7187 1667
rect 7053 1633 7067 1647
rect 7013 1553 7027 1567
rect 6893 1353 6907 1367
rect 6913 1293 6927 1307
rect 6873 1273 6887 1287
rect 6853 1233 6867 1247
rect 6853 873 6867 887
rect 6773 713 6787 727
rect 6833 713 6847 727
rect 6753 633 6767 647
rect 6733 493 6747 507
rect 6313 433 6327 447
rect 6593 433 6607 447
rect 5913 233 5927 247
rect 5973 233 5987 247
rect 5793 193 5807 207
rect 5733 130 5747 144
rect 5773 130 5787 144
rect 5693 93 5707 107
rect 5573 33 5587 47
rect 5833 213 5847 227
rect 5813 93 5827 107
rect 5453 13 5467 27
rect 5493 13 5507 27
rect 5713 13 5727 27
rect 5793 13 5807 27
rect 5953 176 5967 190
rect 6093 396 6107 410
rect 6173 396 6187 410
rect 6213 396 6227 410
rect 6053 373 6067 387
rect 6133 373 6147 387
rect 6293 376 6307 390
rect 6093 313 6107 327
rect 6113 173 6127 187
rect 6233 350 6247 364
rect 6193 313 6207 327
rect 6293 313 6307 327
rect 6233 176 6247 190
rect 6133 153 6147 167
rect 6113 130 6127 144
rect 6213 130 6227 144
rect 6253 130 6267 144
rect 6433 376 6447 390
rect 6593 350 6607 364
rect 6693 333 6707 347
rect 6733 333 6747 347
rect 6673 313 6687 327
rect 6633 293 6647 307
rect 6513 253 6527 267
rect 6453 173 6467 187
rect 6553 213 6567 227
rect 6453 130 6467 144
rect 6493 130 6507 144
rect 6533 130 6547 144
rect 6693 273 6707 287
rect 6753 273 6767 287
rect 6673 253 6687 267
rect 6893 1253 6907 1267
rect 6973 1393 6987 1407
rect 7033 1390 7047 1404
rect 7013 1333 7027 1347
rect 6933 1253 6947 1267
rect 6913 1216 6927 1230
rect 6973 1216 6987 1230
rect 7013 1213 7027 1227
rect 6893 1170 6907 1184
rect 6953 1170 6967 1184
rect 6993 1093 7007 1107
rect 7073 1293 7087 1307
rect 7073 1212 7087 1226
rect 7213 1933 7227 1947
rect 7233 1913 7247 1927
rect 7293 2873 7307 2887
rect 7293 2673 7307 2687
rect 7293 2473 7307 2487
rect 7353 3073 7367 3087
rect 7393 3073 7407 3087
rect 7353 2933 7367 2947
rect 7353 2776 7367 2790
rect 7393 2776 7407 2790
rect 7553 5030 7567 5044
rect 7573 4873 7587 4887
rect 7553 4393 7567 4407
rect 7733 6533 7747 6547
rect 7813 6636 7827 6650
rect 7853 6636 7867 6650
rect 7833 6590 7847 6604
rect 7793 6573 7807 6587
rect 7853 6553 7867 6567
rect 7753 6493 7767 6507
rect 7773 6416 7787 6430
rect 7813 6370 7827 6384
rect 7813 6333 7827 6347
rect 7753 6173 7767 6187
rect 7973 6573 7987 6587
rect 7913 6533 7927 6547
rect 7993 6553 8007 6567
rect 7993 6473 8007 6487
rect 7973 6453 7987 6467
rect 8113 6953 8127 6967
rect 8093 6933 8107 6947
rect 8073 6833 8087 6847
rect 8213 7630 8227 7644
rect 8213 7456 8227 7470
rect 8173 7293 8187 7307
rect 8173 7133 8187 7147
rect 8333 7975 8347 7989
rect 8373 7975 8387 7989
rect 8493 8073 8507 8087
rect 8653 8073 8667 8087
rect 8393 7913 8407 7927
rect 8333 7893 8347 7907
rect 8792 8173 8806 8187
rect 8753 8133 8767 8147
rect 8753 8093 8767 8107
rect 8633 8033 8647 8047
rect 8733 8033 8747 8047
rect 8593 7976 8607 7990
rect 8493 7873 8507 7887
rect 8393 7833 8407 7847
rect 8433 7833 8447 7847
rect 8353 7493 8367 7507
rect 8593 7793 8607 7807
rect 8473 7773 8487 7787
rect 8433 7733 8447 7747
rect 8573 7733 8587 7747
rect 8553 7673 8567 7687
rect 8293 7393 8307 7407
rect 8413 7413 8427 7427
rect 8373 7393 8387 7407
rect 8333 7313 8347 7327
rect 8393 7313 8407 7327
rect 8273 7156 8287 7170
rect 8173 6893 8187 6907
rect 8153 6873 8167 6887
rect 8252 7073 8266 7087
rect 8273 7073 8287 7087
rect 8213 7013 8227 7027
rect 8313 6936 8327 6950
rect 8393 7073 8407 7087
rect 8433 7213 8447 7227
rect 8413 6953 8427 6967
rect 8393 6933 8407 6947
rect 8213 6813 8227 6827
rect 8293 6873 8307 6887
rect 8253 6793 8267 6807
rect 8193 6773 8207 6787
rect 8133 6733 8147 6747
rect 8173 6733 8187 6747
rect 8333 6733 8347 6747
rect 8333 6656 8347 6670
rect 8033 6633 8047 6647
rect 8173 6616 8187 6630
rect 8033 6593 8047 6607
rect 8093 6493 8107 6507
rect 8013 6433 8027 6447
rect 7993 6413 8007 6427
rect 8253 6473 8267 6487
rect 7913 6373 7927 6387
rect 7873 6233 7887 6247
rect 7853 6133 7867 6147
rect 7833 6053 7847 6067
rect 7793 5993 7807 6007
rect 7813 5896 7827 5910
rect 8073 6370 8087 6384
rect 7993 6353 8007 6367
rect 8273 6416 8287 6430
rect 8333 6573 8347 6587
rect 8333 6493 8347 6507
rect 8373 6473 8387 6487
rect 8313 6453 8327 6467
rect 8313 6416 8327 6430
rect 8353 6416 8367 6430
rect 8393 6416 8407 6430
rect 8273 6373 8287 6387
rect 8253 6353 8267 6367
rect 7993 6233 8007 6247
rect 7973 6193 7987 6207
rect 7913 5953 7927 5967
rect 7953 5933 7967 5947
rect 7913 5896 7927 5910
rect 7813 5853 7827 5867
rect 7893 5850 7907 5864
rect 7953 5850 7967 5864
rect 7773 5713 7787 5727
rect 7733 5673 7747 5687
rect 7753 5473 7767 5487
rect 7733 5413 7747 5427
rect 7733 5392 7747 5406
rect 7733 5113 7747 5127
rect 7713 4933 7727 4947
rect 7633 4856 7647 4870
rect 7693 4856 7707 4870
rect 7613 4753 7627 4767
rect 7593 4713 7607 4727
rect 7613 4673 7627 4687
rect 7873 5633 7887 5647
rect 7833 5613 7847 5627
rect 7913 5596 7927 5610
rect 7853 5550 7867 5564
rect 7893 5473 7907 5487
rect 7853 5413 7867 5427
rect 7933 5376 7947 5390
rect 7793 5330 7807 5344
rect 7873 5330 7887 5344
rect 7913 5330 7927 5344
rect 7853 5293 7867 5307
rect 7773 4993 7787 5007
rect 7713 4810 7727 4824
rect 7753 4813 7767 4827
rect 7673 4633 7687 4647
rect 7633 4556 7647 4570
rect 7733 4556 7747 4570
rect 7613 4433 7627 4447
rect 7573 4353 7587 4367
rect 7613 4336 7627 4350
rect 7713 4510 7727 4524
rect 7893 5233 7907 5247
rect 7833 5030 7847 5044
rect 8013 6213 8027 6227
rect 8233 6153 8247 6167
rect 8073 6133 8087 6147
rect 7993 6013 8007 6027
rect 7993 5953 8007 5967
rect 7973 5773 7987 5787
rect 7993 5550 8007 5564
rect 7993 5493 8007 5507
rect 7993 4993 8007 5007
rect 7973 4933 7987 4947
rect 7873 4893 7887 4907
rect 7793 4793 7807 4807
rect 7973 4793 7987 4807
rect 7953 4773 7967 4787
rect 8013 4573 8027 4587
rect 7733 4393 7747 4407
rect 7713 4333 7727 4347
rect 7673 4290 7687 4304
rect 7713 4290 7727 4304
rect 7633 4273 7647 4287
rect 7593 4036 7607 4050
rect 7573 3990 7587 4004
rect 7573 3933 7587 3947
rect 7553 3816 7567 3830
rect 7553 3713 7567 3727
rect 7553 3516 7567 3530
rect 7553 3433 7567 3447
rect 7613 3893 7627 3907
rect 7673 3953 7687 3967
rect 7633 3873 7647 3887
rect 7653 3816 7667 3830
rect 7613 3793 7627 3807
rect 7673 3770 7687 3784
rect 7713 3713 7727 3727
rect 7613 3653 7627 3667
rect 7593 3573 7607 3587
rect 7573 3393 7587 3407
rect 7633 3633 7647 3647
rect 7613 3553 7627 3567
rect 7693 3553 7707 3567
rect 7633 3516 7647 3530
rect 7613 3473 7627 3487
rect 7593 3333 7607 3347
rect 7653 3470 7667 3484
rect 7693 3470 7707 3484
rect 7613 3313 7627 3327
rect 7573 3296 7587 3310
rect 7613 3250 7627 3264
rect 7553 3213 7567 3227
rect 7533 3193 7547 3207
rect 7453 3033 7467 3047
rect 7513 3033 7527 3047
rect 7573 3193 7587 3207
rect 7553 3013 7567 3027
rect 7513 2996 7527 3010
rect 7493 2933 7507 2947
rect 7453 2913 7467 2927
rect 7353 2733 7367 2747
rect 7333 2473 7347 2487
rect 7313 2333 7327 2347
rect 7293 2210 7307 2224
rect 7273 1993 7287 2007
rect 7333 1993 7347 2007
rect 7373 2693 7387 2707
rect 7413 2693 7427 2707
rect 7453 2653 7467 2667
rect 7433 2593 7447 2607
rect 7593 3113 7607 3127
rect 7573 2913 7587 2927
rect 7613 2893 7627 2907
rect 7593 2873 7607 2887
rect 7593 2833 7607 2847
rect 7513 2493 7527 2507
rect 7553 2493 7567 2507
rect 7473 2476 7487 2490
rect 7433 2393 7447 2407
rect 7493 2393 7507 2407
rect 7453 2373 7467 2387
rect 7473 2353 7487 2367
rect 7433 2313 7447 2327
rect 7473 2256 7487 2270
rect 7413 2210 7427 2224
rect 7373 2093 7387 2107
rect 7353 1973 7367 1987
rect 7293 1953 7307 1967
rect 7333 1956 7347 1970
rect 7253 1893 7267 1907
rect 7213 1673 7227 1687
rect 7193 1613 7207 1627
rect 7253 1613 7267 1627
rect 7193 1513 7207 1527
rect 7153 1493 7167 1507
rect 7113 1433 7127 1447
rect 7173 1313 7187 1327
rect 7133 1233 7147 1247
rect 7113 1170 7127 1184
rect 7053 1133 7067 1147
rect 7093 1133 7107 1147
rect 7033 1073 7047 1087
rect 7073 1053 7087 1067
rect 7013 1013 7027 1027
rect 7053 1013 7067 1027
rect 7013 973 7027 987
rect 6953 953 6967 967
rect 6933 915 6947 929
rect 6993 915 7007 929
rect 7033 833 7047 847
rect 6873 793 6887 807
rect 6972 793 6986 807
rect 6993 793 7007 807
rect 6933 733 6947 747
rect 7253 1313 7267 1327
rect 7253 1233 7267 1247
rect 7333 1893 7347 1907
rect 7353 1873 7367 1887
rect 7393 1813 7407 1827
rect 7293 1633 7307 1647
rect 7293 1573 7307 1587
rect 7333 1673 7347 1687
rect 7313 1493 7327 1507
rect 7353 1593 7367 1607
rect 7353 1553 7367 1567
rect 7333 1353 7347 1367
rect 7193 1170 7207 1184
rect 7153 1093 7167 1107
rect 7233 1033 7247 1047
rect 7593 2173 7607 2187
rect 7673 3250 7687 3264
rect 7953 4473 7967 4487
rect 7853 4433 7867 4447
rect 7993 4433 8007 4447
rect 7773 4113 7787 4127
rect 8013 4413 8027 4427
rect 7993 4393 8007 4407
rect 7873 4353 7887 4367
rect 7933 4353 7947 4367
rect 7853 4036 7867 4050
rect 7773 3990 7787 4004
rect 7813 3990 7827 4004
rect 7873 3993 7887 4007
rect 7753 3793 7767 3807
rect 7753 3733 7767 3747
rect 7733 3633 7747 3647
rect 7773 3693 7787 3707
rect 7753 3513 7767 3527
rect 7693 3053 7707 3067
rect 7673 2993 7687 3007
rect 7673 2950 7687 2964
rect 7813 3793 7827 3807
rect 7793 3633 7807 3647
rect 7773 3453 7787 3467
rect 7753 3033 7767 3047
rect 7753 2996 7767 3010
rect 7733 2950 7747 2964
rect 7733 2776 7747 2790
rect 7753 2713 7767 2727
rect 7793 2653 7807 2667
rect 7713 2613 7727 2627
rect 7633 2553 7647 2567
rect 7753 2513 7767 2527
rect 7773 2430 7787 2444
rect 7653 2293 7667 2307
rect 7733 2293 7747 2307
rect 7793 2293 7807 2307
rect 7693 2256 7707 2270
rect 7733 2256 7747 2270
rect 7613 2133 7627 2147
rect 7453 2073 7467 2087
rect 7453 1956 7467 1970
rect 7573 1956 7587 1970
rect 7613 1956 7627 1970
rect 7713 2210 7727 2224
rect 7773 2133 7787 2147
rect 7753 2073 7767 2087
rect 7713 1993 7727 2007
rect 7633 1910 7647 1924
rect 7673 1913 7687 1927
rect 7453 1873 7467 1887
rect 7593 1873 7607 1887
rect 7673 1873 7687 1887
rect 7553 1813 7567 1827
rect 7593 1773 7607 1787
rect 7633 1736 7647 1750
rect 7453 1593 7467 1607
rect 7573 1593 7587 1607
rect 7393 1533 7407 1547
rect 7373 1390 7387 1404
rect 7493 1493 7507 1507
rect 7493 1436 7507 1450
rect 7633 1633 7647 1647
rect 7613 1573 7627 1587
rect 7613 1436 7627 1450
rect 7433 1390 7447 1404
rect 7393 1293 7407 1307
rect 7573 1390 7587 1404
rect 7473 1273 7487 1287
rect 7573 1273 7587 1287
rect 7513 1253 7527 1267
rect 7473 1216 7487 1230
rect 7453 1173 7467 1187
rect 7593 1216 7607 1230
rect 7353 1053 7367 1067
rect 7232 973 7246 987
rect 7253 973 7267 987
rect 7293 973 7307 987
rect 7132 915 7146 929
rect 7153 913 7167 927
rect 7293 915 7307 929
rect 7533 1170 7547 1184
rect 7573 1170 7587 1184
rect 7553 1133 7567 1147
rect 7473 1093 7487 1107
rect 7493 1093 7507 1107
rect 7453 916 7467 930
rect 7253 869 7267 883
rect 7333 869 7347 883
rect 7393 853 7407 867
rect 7153 813 7167 827
rect 7213 733 7227 747
rect 7253 733 7267 747
rect 7133 696 7147 710
rect 7173 696 7187 710
rect 7073 673 7087 687
rect 6793 613 6807 627
rect 6773 253 6787 267
rect 6893 651 6907 665
rect 6993 651 7007 665
rect 6993 573 7007 587
rect 6833 553 6847 567
rect 6813 433 6827 447
rect 7193 650 7207 664
rect 7233 633 7247 647
rect 7233 533 7247 547
rect 7133 513 7147 527
rect 6933 433 6947 447
rect 6993 433 7007 447
rect 6873 373 6887 387
rect 7033 370 7047 384
rect 7153 376 7167 390
rect 6913 333 6927 347
rect 7493 650 7507 664
rect 7533 396 7547 410
rect 7413 353 7427 367
rect 7453 353 7467 367
rect 7353 293 7367 307
rect 6993 253 7007 267
rect 6793 213 6807 227
rect 6713 173 6727 187
rect 6753 176 6767 190
rect 7293 176 7307 190
rect 7353 173 7367 187
rect 7753 1956 7767 1970
rect 7713 1736 7727 1750
rect 7713 1453 7727 1467
rect 7793 1953 7807 1967
rect 7793 1673 7807 1687
rect 7773 1473 7787 1487
rect 7853 3973 7867 3987
rect 7913 4273 7927 4287
rect 7893 3973 7907 3987
rect 7993 4033 8007 4047
rect 7993 3990 8007 4004
rect 8093 6070 8107 6084
rect 8193 6053 8207 6067
rect 8153 5933 8167 5947
rect 8113 5896 8127 5910
rect 8133 5850 8147 5864
rect 8193 5853 8207 5867
rect 8173 5713 8187 5727
rect 8173 5673 8187 5687
rect 8073 5596 8087 5610
rect 8133 5596 8147 5610
rect 8213 5633 8227 5647
rect 8113 5493 8127 5507
rect 8153 5493 8167 5507
rect 8213 5433 8227 5447
rect 8093 5393 8107 5407
rect 8073 5153 8087 5167
rect 8073 5113 8087 5127
rect 8133 5376 8147 5390
rect 8173 5376 8187 5390
rect 8213 5376 8227 5390
rect 8153 5293 8167 5307
rect 8213 5293 8227 5307
rect 8153 5272 8167 5286
rect 8153 5133 8167 5147
rect 8153 5076 8167 5090
rect 8333 6333 8347 6347
rect 8473 7613 8487 7627
rect 8513 7413 8527 7427
rect 8553 7193 8567 7207
rect 8713 8013 8727 8027
rect 8673 7976 8687 7990
rect 8753 7993 8767 8007
rect 8733 7930 8747 7944
rect 8693 7913 8707 7927
rect 8813 8170 8827 8184
rect 8833 8153 8847 8167
rect 8813 8133 8827 8147
rect 8772 7873 8786 7887
rect 8793 7873 8807 7887
rect 8693 7733 8707 7747
rect 8673 7676 8687 7690
rect 8733 7676 8747 7690
rect 8633 7653 8647 7667
rect 8673 7633 8687 7647
rect 8613 7613 8627 7627
rect 8713 7613 8727 7627
rect 8633 7513 8647 7527
rect 8673 7513 8687 7527
rect 8653 7456 8667 7470
rect 8613 7353 8627 7367
rect 8613 7156 8627 7170
rect 8653 7156 8667 7170
rect 8533 6993 8547 7007
rect 8593 7093 8607 7107
rect 8653 7053 8667 7067
rect 8593 7033 8607 7047
rect 8553 6973 8567 6987
rect 8453 6753 8467 6767
rect 8473 6733 8487 6747
rect 8453 6713 8467 6727
rect 8453 6656 8467 6670
rect 8453 6293 8467 6307
rect 8433 6253 8447 6267
rect 8353 6173 8367 6187
rect 8393 6116 8407 6130
rect 8333 6070 8347 6084
rect 8373 6053 8387 6067
rect 8393 5973 8407 5987
rect 8333 5850 8347 5864
rect 8313 5653 8327 5667
rect 8253 5596 8267 5610
rect 8253 5533 8267 5547
rect 8273 5393 8287 5407
rect 8273 5076 8287 5090
rect 8253 5053 8267 5067
rect 8072 5033 8086 5047
rect 8093 5033 8107 5047
rect 8053 4993 8067 5007
rect 8053 4573 8067 4587
rect 8073 4510 8087 4524
rect 8073 4473 8087 4487
rect 8053 4413 8067 4427
rect 8053 4333 8067 4347
rect 8133 5030 8147 5044
rect 8153 4953 8167 4967
rect 8153 4793 8167 4807
rect 8113 4733 8127 4747
rect 8093 4293 8107 4307
rect 8053 4273 8067 4287
rect 8093 4093 8107 4107
rect 8273 5033 8287 5047
rect 8233 4993 8247 5007
rect 8273 4856 8287 4870
rect 8173 4693 8187 4707
rect 8213 4773 8227 4787
rect 8253 4733 8267 4747
rect 8193 4673 8207 4687
rect 8413 5850 8427 5864
rect 8553 6853 8567 6867
rect 8533 6813 8547 6827
rect 8513 6673 8527 6687
rect 8493 6533 8507 6547
rect 8693 6936 8707 6950
rect 8693 6853 8707 6867
rect 8553 6693 8567 6707
rect 8593 6693 8607 6707
rect 8813 7456 8827 7470
rect 8753 7433 8767 7447
rect 8873 8773 8887 8787
rect 8933 8893 8947 8907
rect 8913 8873 8927 8887
rect 8893 8753 8907 8767
rect 8873 7930 8887 7944
rect 8853 7833 8867 7847
rect 8893 7613 8907 7627
rect 8932 8793 8946 8807
rect 8953 8793 8967 8807
rect 9733 11173 9747 11187
rect 9713 11033 9727 11047
rect 9713 10953 9727 10967
rect 9653 10933 9667 10947
rect 9573 10813 9587 10827
rect 9753 10833 9767 10847
rect 10013 11633 10027 11647
rect 10053 11633 10067 11647
rect 10033 11570 10047 11584
rect 9993 11533 10007 11547
rect 9993 11433 10007 11447
rect 9853 11353 9867 11367
rect 9573 10753 9587 10767
rect 9693 10750 9707 10764
rect 9733 10750 9747 10764
rect 9233 10713 9247 10727
rect 9253 10673 9267 10687
rect 9233 10576 9247 10590
rect 9233 9853 9247 9867
rect 9433 10633 9447 10647
rect 9353 10576 9367 10590
rect 9333 10530 9347 10544
rect 9493 10576 9507 10590
rect 9413 10230 9427 10244
rect 9573 10613 9587 10627
rect 9613 10576 9627 10590
rect 9653 10576 9667 10590
rect 9533 10533 9547 10547
rect 9593 10530 9607 10544
rect 9673 10493 9687 10507
rect 9653 10433 9667 10447
rect 9693 10333 9707 10347
rect 9453 10193 9467 10207
rect 9493 10193 9507 10207
rect 9273 10053 9287 10067
rect 9333 10056 9347 10070
rect 9533 10056 9547 10070
rect 9573 10056 9587 10070
rect 9613 10056 9627 10070
rect 9353 10010 9367 10024
rect 9293 9973 9307 9987
rect 9273 9873 9287 9887
rect 9253 9753 9267 9767
rect 9333 9953 9347 9967
rect 9333 9913 9347 9927
rect 9453 9913 9467 9927
rect 9233 9713 9247 9727
rect 9273 9710 9287 9724
rect 9253 9553 9267 9567
rect 9233 9533 9247 9547
rect 9253 9513 9267 9527
rect 9233 9413 9247 9427
rect 9393 9653 9407 9667
rect 9353 9536 9367 9550
rect 9413 9536 9427 9550
rect 9313 9513 9327 9527
rect 9373 9490 9387 9504
rect 9433 9453 9447 9467
rect 9273 9353 9287 9367
rect 9273 9293 9287 9307
rect 9213 9233 9227 9247
rect 9313 9236 9327 9250
rect 9253 9190 9267 9204
rect 9093 9093 9107 9107
rect 9293 9093 9307 9107
rect 9333 9093 9347 9107
rect 9393 9236 9407 9250
rect 9213 8990 9227 9004
rect 9313 8990 9327 9004
rect 9393 8993 9407 9007
rect 9373 8950 9387 8964
rect 9213 8873 9227 8887
rect 9193 8853 9207 8867
rect 9053 8713 9067 8727
rect 9113 8713 9127 8727
rect 9173 8670 9187 8684
rect 9113 8653 9127 8667
rect 8933 8613 8947 8627
rect 9073 8613 9087 8627
rect 9053 8593 9067 8607
rect 8933 8573 8947 8587
rect 8933 8496 8947 8510
rect 8973 8496 8987 8510
rect 9013 8496 9027 8510
rect 8993 8450 9007 8464
rect 8993 8353 9007 8367
rect 8973 8196 8987 8210
rect 8953 8133 8967 8147
rect 8933 7933 8947 7947
rect 8913 7533 8927 7547
rect 9053 8413 9067 8427
rect 9053 8333 9067 8347
rect 9033 8313 9047 8327
rect 9093 8253 9107 8267
rect 9053 8196 9067 8210
rect 9173 8613 9187 8627
rect 9173 8493 9187 8507
rect 9153 8173 9167 8187
rect 9113 8133 9127 8147
rect 9073 8113 9087 8127
rect 9133 8093 9147 8107
rect 9253 8753 9267 8767
rect 9233 8653 9247 8667
rect 9213 8633 9227 8647
rect 9233 8533 9247 8547
rect 9213 8196 9227 8210
rect 9333 8716 9347 8730
rect 9353 8653 9367 8667
rect 9313 8633 9327 8647
rect 9313 8496 9327 8510
rect 9253 8450 9267 8464
rect 9293 8450 9307 8464
rect 9333 8450 9347 8464
rect 9433 8973 9447 8987
rect 9433 8873 9447 8887
rect 9633 9993 9647 10007
rect 9593 9893 9607 9907
rect 9553 9813 9567 9827
rect 9693 10073 9707 10087
rect 9673 9933 9687 9947
rect 9593 9772 9607 9786
rect 9633 9773 9647 9787
rect 9633 9710 9647 9724
rect 9573 9693 9587 9707
rect 9673 9653 9687 9667
rect 9513 9613 9527 9627
rect 9553 9613 9567 9627
rect 9693 9613 9707 9627
rect 9493 9553 9507 9567
rect 9473 9513 9487 9527
rect 9473 8753 9487 8767
rect 9653 9536 9667 9550
rect 9633 9490 9647 9504
rect 9733 10173 9747 10187
rect 9593 9393 9607 9407
rect 9553 9293 9567 9307
rect 9513 9236 9527 9250
rect 9553 9236 9567 9250
rect 9593 9236 9607 9250
rect 9633 9236 9647 9250
rect 9573 9093 9587 9107
rect 9553 9033 9567 9047
rect 9633 9033 9647 9047
rect 9533 9013 9547 9027
rect 9533 8893 9547 8907
rect 9553 8873 9567 8887
rect 9713 9333 9727 9347
rect 9713 9193 9727 9207
rect 9713 9073 9727 9087
rect 9653 8933 9667 8947
rect 9693 8933 9707 8947
rect 9653 8873 9667 8887
rect 9513 8813 9527 8827
rect 9593 8813 9607 8827
rect 9633 8813 9647 8827
rect 9593 8716 9607 8730
rect 9553 8670 9567 8684
rect 9573 8593 9587 8607
rect 9513 8553 9527 8567
rect 9493 8493 9507 8507
rect 9473 8450 9487 8464
rect 9493 8293 9507 8307
rect 9373 8273 9387 8287
rect 9453 8273 9467 8287
rect 9333 8196 9347 8210
rect 9233 8133 9247 8147
rect 9213 8113 9227 8127
rect 9393 8150 9407 8164
rect 9253 8093 9267 8107
rect 9353 8093 9367 8107
rect 9193 8073 9207 8087
rect 9113 8033 9127 8047
rect 8993 7993 9007 8007
rect 9013 7976 9027 7990
rect 9053 7973 9067 7987
rect 9053 7956 9067 7970
rect 9153 7973 9167 7987
rect 8953 7773 8967 7787
rect 8993 7930 9007 7944
rect 9033 7913 9047 7927
rect 8993 7793 9007 7807
rect 9113 7873 9127 7887
rect 9093 7833 9107 7847
rect 9033 7676 9047 7690
rect 8953 7633 8967 7647
rect 9013 7630 9027 7644
rect 8993 7533 9007 7547
rect 9033 7533 9047 7547
rect 8953 7513 8967 7527
rect 8933 7473 8947 7487
rect 8893 7456 8907 7470
rect 8973 7473 8987 7487
rect 8913 7410 8927 7424
rect 8873 7253 8887 7267
rect 8833 7213 8847 7227
rect 8993 7410 9007 7424
rect 8753 7193 8767 7207
rect 8853 7193 8867 7207
rect 8973 7193 8987 7207
rect 8753 7110 8767 7124
rect 8833 7110 8847 7124
rect 8813 7033 8827 7047
rect 8773 6936 8787 6950
rect 8793 6890 8807 6904
rect 8833 6890 8847 6904
rect 9013 7110 9027 7124
rect 8933 7093 8947 7107
rect 8893 6993 8907 7007
rect 8893 6890 8907 6904
rect 8733 6753 8747 6767
rect 8873 6753 8887 6767
rect 8713 6673 8727 6687
rect 8553 6653 8567 6667
rect 8573 6636 8587 6650
rect 8553 6593 8567 6607
rect 8553 6553 8567 6567
rect 8533 6533 8547 6547
rect 8513 6433 8527 6447
rect 8513 6253 8527 6267
rect 8473 5793 8487 5807
rect 8393 5733 8407 5747
rect 8373 5713 8387 5727
rect 8393 5693 8407 5707
rect 8333 5633 8347 5647
rect 8453 5596 8467 5610
rect 8433 5550 8447 5564
rect 8373 5453 8387 5467
rect 8373 5353 8387 5367
rect 8413 5293 8427 5307
rect 8493 5333 8507 5347
rect 8473 5173 8487 5187
rect 8393 5076 8407 5090
rect 8433 5076 8447 5090
rect 8353 4852 8367 4866
rect 8333 4573 8347 4587
rect 8133 4556 8147 4570
rect 8193 4556 8207 4570
rect 8233 4556 8247 4570
rect 8313 4556 8327 4570
rect 8213 4510 8227 4524
rect 8273 4510 8287 4524
rect 8253 4473 8267 4487
rect 8193 4373 8207 4387
rect 8233 4336 8247 4350
rect 8173 4293 8187 4307
rect 8133 4193 8147 4207
rect 8133 4036 8147 4050
rect 8033 3973 8047 3987
rect 7973 3933 7987 3947
rect 8013 3913 8027 3927
rect 7933 3853 7947 3867
rect 7973 3816 7987 3830
rect 7953 3770 7967 3784
rect 8013 3773 8027 3787
rect 7913 3733 7927 3747
rect 7993 3733 8007 3747
rect 7873 3713 7887 3727
rect 7933 3533 7947 3547
rect 7973 3533 7987 3547
rect 7873 3516 7887 3530
rect 7913 3470 7927 3484
rect 7893 3453 7907 3467
rect 7973 3413 7987 3427
rect 7833 3250 7847 3264
rect 7873 3250 7887 3264
rect 7913 3250 7927 3264
rect 7893 3213 7907 3227
rect 7832 3073 7846 3087
rect 7853 3073 7867 3087
rect 7833 2833 7847 2847
rect 7853 2776 7867 2790
rect 7833 2713 7847 2727
rect 7853 2573 7867 2587
rect 7833 2153 7847 2167
rect 7873 2553 7887 2567
rect 7913 3133 7927 3147
rect 7973 3296 7987 3310
rect 7973 3233 7987 3247
rect 8013 3633 8027 3647
rect 8073 3990 8087 4004
rect 8113 3990 8127 4004
rect 8073 3969 8087 3983
rect 8053 3816 8067 3830
rect 8053 3713 8067 3727
rect 8053 3533 8067 3547
rect 8033 3353 8047 3367
rect 8033 3293 8047 3307
rect 8013 3193 8027 3207
rect 7993 3133 8007 3147
rect 7913 3053 7927 3067
rect 7953 3033 7967 3047
rect 7993 2996 8007 3010
rect 8053 3113 8067 3127
rect 8113 3853 8127 3867
rect 8093 3753 8107 3767
rect 8213 4273 8227 4287
rect 8233 4193 8247 4207
rect 8213 4036 8227 4050
rect 8193 3933 8207 3947
rect 8173 3853 8187 3867
rect 8253 4093 8267 4107
rect 8253 4036 8267 4050
rect 8253 3913 8267 3927
rect 8153 3753 8167 3767
rect 8213 3753 8227 3767
rect 8133 3573 8147 3587
rect 8193 3573 8207 3587
rect 8173 3533 8187 3547
rect 8133 3513 8147 3527
rect 8233 3693 8247 3707
rect 8232 3653 8246 3667
rect 8253 3653 8267 3667
rect 8213 3516 8227 3530
rect 8253 3516 8267 3530
rect 8153 3470 8167 3484
rect 8193 3413 8207 3427
rect 8193 3373 8207 3387
rect 8213 3353 8227 3367
rect 8153 3333 8167 3347
rect 8193 3333 8207 3347
rect 8093 3250 8107 3264
rect 8073 2993 8087 3007
rect 8053 2950 8067 2964
rect 8013 2793 8027 2807
rect 8053 2873 8067 2887
rect 7913 2533 7927 2547
rect 8033 2773 8047 2787
rect 7993 2730 8007 2744
rect 7953 2473 7967 2487
rect 8013 2476 8027 2490
rect 8073 2733 8087 2747
rect 8073 2673 8087 2687
rect 8073 2633 8087 2647
rect 8053 2473 8067 2487
rect 7933 2430 7947 2444
rect 7913 2393 7927 2407
rect 7893 2256 7907 2270
rect 7993 2430 8007 2444
rect 8033 2333 8047 2347
rect 7853 2013 7867 2027
rect 7953 2253 7967 2267
rect 7993 2256 8007 2270
rect 7973 2210 7987 2224
rect 8033 2210 8047 2224
rect 7973 2073 7987 2087
rect 7833 1893 7847 1907
rect 7873 1893 7887 1907
rect 7853 1853 7867 1867
rect 7913 1873 7927 1887
rect 7973 1873 7987 1887
rect 7853 1690 7867 1704
rect 7873 1633 7887 1647
rect 7853 1593 7867 1607
rect 7853 1473 7867 1487
rect 7733 1390 7747 1404
rect 7713 1293 7727 1307
rect 7673 1273 7687 1287
rect 7733 1253 7747 1267
rect 7773 1233 7787 1247
rect 7733 1213 7747 1227
rect 7813 1216 7827 1230
rect 7793 1170 7807 1184
rect 7833 1173 7847 1187
rect 7813 1153 7827 1167
rect 7593 993 7607 1007
rect 7573 953 7587 967
rect 7713 933 7727 947
rect 7613 916 7627 930
rect 7793 1113 7807 1127
rect 7773 890 7787 904
rect 7633 870 7647 884
rect 7713 870 7727 884
rect 7673 813 7687 827
rect 7813 993 7827 1007
rect 7793 753 7807 767
rect 7653 733 7667 747
rect 7573 650 7587 664
rect 7733 713 7747 727
rect 7833 833 7847 847
rect 7773 650 7787 664
rect 7813 653 7827 667
rect 7653 613 7667 627
rect 7633 350 7647 364
rect 7553 273 7567 287
rect 7913 1613 7927 1627
rect 7893 1513 7907 1527
rect 8013 1873 8027 1887
rect 8053 1690 8067 1704
rect 7993 1533 8007 1547
rect 7913 1233 7927 1247
rect 7893 1213 7907 1227
rect 7873 1153 7887 1167
rect 7873 1033 7887 1047
rect 7873 953 7887 967
rect 8113 3173 8127 3187
rect 8093 1953 8107 1967
rect 8193 3253 8207 3267
rect 8173 3233 8187 3247
rect 8152 3193 8166 3207
rect 8173 3193 8187 3207
rect 8173 3113 8187 3127
rect 8153 2573 8167 2587
rect 8133 2113 8147 2127
rect 8173 2476 8187 2490
rect 8253 3253 8267 3267
rect 8293 4433 8307 4447
rect 8273 3173 8287 3187
rect 8233 3113 8247 3127
rect 8233 3053 8247 3067
rect 8453 5030 8467 5044
rect 8493 5030 8507 5044
rect 8413 4993 8427 5007
rect 8373 4793 8387 4807
rect 8393 4510 8407 4524
rect 8353 4393 8367 4407
rect 8313 4336 8327 4350
rect 8693 6593 8707 6607
rect 8633 6553 8647 6567
rect 8653 6553 8667 6567
rect 8593 6533 8607 6547
rect 8573 6433 8587 6447
rect 8553 6413 8567 6427
rect 8613 6416 8627 6430
rect 8693 6493 8707 6507
rect 8593 6370 8607 6384
rect 8633 6353 8647 6367
rect 8533 5853 8547 5867
rect 8533 5553 8547 5567
rect 8533 5393 8547 5407
rect 8533 5330 8547 5344
rect 8613 6116 8627 6130
rect 8573 6070 8587 6084
rect 8573 6013 8587 6027
rect 8573 5913 8587 5927
rect 8573 5593 8587 5607
rect 8553 5193 8567 5207
rect 8553 5153 8567 5167
rect 8533 5133 8547 5147
rect 8533 5013 8547 5027
rect 8513 4993 8527 5007
rect 8433 4973 8447 4987
rect 8513 4933 8527 4947
rect 8633 5993 8647 6007
rect 8693 5913 8707 5927
rect 8613 5896 8627 5910
rect 8653 5896 8667 5910
rect 8673 5850 8687 5864
rect 8713 5833 8727 5847
rect 8693 5813 8707 5827
rect 8713 5773 8727 5787
rect 8633 5753 8647 5767
rect 8613 5513 8627 5527
rect 8653 5733 8667 5747
rect 9053 7156 9067 7170
rect 9093 7573 9107 7587
rect 9133 7673 9147 7687
rect 9113 7553 9127 7567
rect 9093 7333 9107 7347
rect 9313 7950 9327 7964
rect 9493 8150 9507 8164
rect 9553 8433 9567 8447
rect 9633 8433 9647 8447
rect 9553 8353 9567 8367
rect 9613 8273 9627 8287
rect 9553 8233 9567 8247
rect 9533 8193 9547 8207
rect 9513 7930 9527 7944
rect 9173 7793 9187 7807
rect 9293 7733 9307 7747
rect 9473 7713 9487 7727
rect 9293 7676 9307 7690
rect 9533 7853 9547 7867
rect 9673 8493 9687 8507
rect 9673 8273 9687 8287
rect 9653 8233 9667 8247
rect 9653 8196 9667 8210
rect 9593 8133 9607 8147
rect 9573 8013 9587 8027
rect 9553 7833 9567 7847
rect 9633 8113 9647 8127
rect 9753 9833 9767 9847
rect 9753 9693 9767 9707
rect 9753 9573 9767 9587
rect 9753 9490 9767 9504
rect 9913 11093 9927 11107
rect 9953 11096 9967 11110
rect 10033 11316 10047 11330
rect 10092 11313 10106 11327
rect 10113 11313 10127 11327
rect 10053 11270 10067 11284
rect 10053 11113 10067 11127
rect 9873 10913 9887 10927
rect 9873 10713 9887 10727
rect 10073 11096 10087 11110
rect 10052 11050 10066 11064
rect 10073 11053 10087 11067
rect 10013 10873 10027 10887
rect 9913 10673 9927 10687
rect 9833 10513 9847 10527
rect 9993 10750 10007 10764
rect 10033 10750 10047 10764
rect 10013 10613 10027 10627
rect 10113 11270 10127 11284
rect 10393 12090 10407 12104
rect 10453 12090 10467 12104
rect 10513 12053 10527 12067
rect 10353 11953 10367 11967
rect 10233 11853 10247 11867
rect 10213 11836 10227 11850
rect 10573 11893 10587 11907
rect 10533 11853 10547 11867
rect 10173 11816 10187 11830
rect 10373 11790 10387 11804
rect 10213 11773 10227 11787
rect 10253 11773 10267 11787
rect 10153 11493 10167 11507
rect 10353 11753 10367 11767
rect 10293 11713 10307 11727
rect 10253 11633 10267 11647
rect 10353 11613 10367 11627
rect 10273 11570 10287 11584
rect 10313 11570 10327 11584
rect 10353 11570 10367 11584
rect 10333 11413 10347 11427
rect 10213 11333 10227 11347
rect 10173 11313 10187 11327
rect 10273 11316 10287 11330
rect 10153 11253 10167 11267
rect 10133 10853 10147 10867
rect 10053 10593 10067 10607
rect 10093 10593 10107 10607
rect 10013 10493 10027 10507
rect 9953 10373 9967 10387
rect 9873 10253 9887 10267
rect 10033 10253 10047 10267
rect 9933 10230 9947 10244
rect 9933 10173 9947 10187
rect 9933 10093 9947 10107
rect 9893 10073 9907 10087
rect 9833 10053 9847 10067
rect 10013 10230 10027 10244
rect 9993 10073 10007 10087
rect 9973 10056 9987 10070
rect 9833 10010 9847 10024
rect 9873 10010 9887 10024
rect 9913 10010 9927 10024
rect 9813 9913 9827 9927
rect 9953 9853 9967 9867
rect 9873 9756 9887 9770
rect 9853 9710 9867 9724
rect 9953 9693 9967 9707
rect 9853 9613 9867 9627
rect 9853 9533 9867 9547
rect 9913 9536 9927 9550
rect 9853 9490 9867 9504
rect 9893 9490 9907 9504
rect 9933 9490 9947 9504
rect 9833 9373 9847 9387
rect 9753 9313 9767 9327
rect 9793 9313 9807 9327
rect 9753 8873 9767 8887
rect 9953 9373 9967 9387
rect 9933 9093 9947 9107
rect 9913 9073 9927 9087
rect 9913 9033 9927 9047
rect 9893 9016 9907 9030
rect 9833 8933 9847 8947
rect 9813 8853 9827 8867
rect 9773 8713 9787 8727
rect 9913 8970 9927 8984
rect 9953 8970 9967 8984
rect 9873 8893 9887 8907
rect 9933 8793 9947 8807
rect 9753 8670 9767 8684
rect 9813 8670 9827 8684
rect 9933 8673 9947 8687
rect 9953 8633 9967 8647
rect 9853 8613 9867 8627
rect 10033 9692 10047 9706
rect 10013 9673 10027 9687
rect 9993 9233 10007 9247
rect 9973 8553 9987 8567
rect 9773 8493 9787 8507
rect 9813 8450 9827 8464
rect 9873 8353 9887 8367
rect 9833 8293 9847 8307
rect 9733 8273 9747 8287
rect 9713 8013 9727 8027
rect 9593 7976 9607 7990
rect 9693 7976 9707 7990
rect 9793 8193 9807 8207
rect 9773 8113 9787 8127
rect 10013 9193 10027 9207
rect 10013 8970 10027 8984
rect 10013 8727 10027 8730
rect 10013 8716 10027 8727
rect 10113 10576 10127 10590
rect 10293 11270 10307 11284
rect 10333 11270 10347 11284
rect 10253 11253 10267 11267
rect 10253 11096 10267 11110
rect 10233 11050 10247 11064
rect 10293 10873 10307 10887
rect 10253 10796 10267 10810
rect 10273 10750 10287 10764
rect 10313 10750 10327 10764
rect 10273 10713 10287 10727
rect 10253 10573 10267 10587
rect 10093 10530 10107 10544
rect 10173 10530 10187 10544
rect 10253 10530 10267 10544
rect 10213 10393 10227 10407
rect 10093 10293 10107 10307
rect 10073 10010 10087 10024
rect 10153 10230 10167 10244
rect 10193 10230 10207 10244
rect 10213 10193 10227 10207
rect 10313 10576 10327 10590
rect 10533 11790 10547 11804
rect 10493 11713 10507 11727
rect 10393 11633 10407 11647
rect 10513 11616 10527 11630
rect 10633 12073 10647 12087
rect 10753 12093 10767 12107
rect 10713 12053 10727 12067
rect 10673 12013 10687 12027
rect 10733 11873 10747 11887
rect 10853 11873 10867 11887
rect 10693 11836 10707 11850
rect 10813 11836 10827 11850
rect 10593 11693 10607 11707
rect 10613 11616 10627 11630
rect 10393 11573 10407 11587
rect 10413 11316 10427 11330
rect 10593 11570 10607 11584
rect 10553 11553 10567 11567
rect 10793 11790 10807 11804
rect 10853 11790 10867 11804
rect 10753 11693 10767 11707
rect 10853 11616 10867 11630
rect 10693 11533 10707 11547
rect 10593 11393 10607 11407
rect 10633 11393 10647 11407
rect 10553 11353 10567 11367
rect 10393 11096 10407 11110
rect 10513 11313 10527 11327
rect 10593 11316 10607 11330
rect 10633 11293 10647 11307
rect 10673 11293 10687 11307
rect 10473 11270 10487 11284
rect 10533 11270 10547 11284
rect 10573 11233 10587 11247
rect 10493 11050 10507 11064
rect 10453 11013 10467 11027
rect 10413 10873 10427 10887
rect 10633 10873 10647 10887
rect 10533 10833 10547 10847
rect 10433 10796 10447 10810
rect 10593 10796 10607 10810
rect 10393 10713 10407 10727
rect 10453 10753 10467 10767
rect 10433 10613 10447 10627
rect 10413 10576 10427 10590
rect 10233 10173 10247 10187
rect 10273 10173 10287 10187
rect 10133 9993 10147 10007
rect 10213 10013 10227 10027
rect 10193 9953 10207 9967
rect 10172 9913 10186 9927
rect 10193 9913 10207 9927
rect 10233 9873 10247 9887
rect 10093 9853 10107 9867
rect 10073 9793 10087 9807
rect 10073 9753 10087 9767
rect 10133 9756 10147 9770
rect 10233 9753 10247 9767
rect 10293 9756 10307 9770
rect 10073 9710 10087 9724
rect 10073 9573 10087 9587
rect 10073 9490 10087 9504
rect 10073 9273 10087 9287
rect 10053 9233 10067 9247
rect 10113 9710 10127 9724
rect 10173 9713 10187 9727
rect 10153 9693 10167 9707
rect 10113 9633 10127 9647
rect 10293 9673 10307 9687
rect 10273 9613 10287 9627
rect 10173 9535 10187 9549
rect 10193 9490 10207 9504
rect 10113 9453 10127 9467
rect 10253 9433 10267 9447
rect 10213 9413 10227 9427
rect 10213 9333 10227 9347
rect 10193 9313 10207 9327
rect 10133 9273 10147 9287
rect 10093 9233 10107 9247
rect 10253 9236 10267 9250
rect 10093 9193 10107 9207
rect 10113 9133 10127 9147
rect 10153 9133 10167 9147
rect 10093 9033 10107 9047
rect 10153 9016 10167 9030
rect 10133 8970 10147 8984
rect 10093 8933 10107 8947
rect 10173 8933 10187 8947
rect 10153 8773 10167 8787
rect 10113 8716 10127 8730
rect 10133 8670 10147 8684
rect 10293 9533 10307 9547
rect 10293 9190 10307 9204
rect 10573 10693 10587 10707
rect 10833 11433 10847 11447
rect 10893 11353 10907 11367
rect 10753 11316 10767 11330
rect 10853 11316 10867 11330
rect 10713 11153 10727 11167
rect 10873 11233 10887 11247
rect 10813 11213 10827 11227
rect 10833 11173 10847 11187
rect 10773 11050 10787 11064
rect 10813 11050 10827 11064
rect 10773 10953 10787 10967
rect 10833 10853 10847 10867
rect 10733 10833 10747 10847
rect 10813 10833 10827 10847
rect 10713 10796 10727 10810
rect 10853 10796 10867 10810
rect 10893 10796 10907 10810
rect 10673 10750 10687 10764
rect 10353 10530 10367 10544
rect 10393 10530 10407 10544
rect 10453 10530 10467 10544
rect 10533 10533 10547 10547
rect 10473 10453 10487 10467
rect 10353 10333 10367 10347
rect 10353 10230 10367 10244
rect 10453 10230 10467 10244
rect 10493 10173 10507 10187
rect 10433 10093 10447 10107
rect 10453 10010 10467 10024
rect 10393 9973 10407 9987
rect 10513 9973 10527 9987
rect 10453 9833 10467 9847
rect 10353 9793 10367 9807
rect 10393 9793 10407 9807
rect 10353 9756 10367 9770
rect 10373 9535 10387 9549
rect 10493 9793 10507 9807
rect 10373 9253 10387 9267
rect 10513 9493 10527 9507
rect 10573 10393 10587 10407
rect 10553 10153 10567 10167
rect 10553 10073 10567 10087
rect 10553 9753 10567 9767
rect 10533 9473 10547 9487
rect 10493 9373 10507 9387
rect 10513 9253 10527 9267
rect 10353 9190 10367 9204
rect 10393 9190 10407 9204
rect 10433 9190 10447 9204
rect 10393 9016 10407 9030
rect 10513 9053 10527 9067
rect 10333 8713 10347 8727
rect 10373 8716 10387 8730
rect 10593 10276 10607 10290
rect 10653 10530 10667 10544
rect 10653 10393 10667 10407
rect 10793 10750 10807 10764
rect 10833 10733 10847 10747
rect 11013 12093 11027 12107
rect 11033 12073 11047 12087
rect 10973 12033 10987 12047
rect 11093 12093 11107 12107
rect 11373 12073 11387 12087
rect 11213 11853 11227 11867
rect 11353 11853 11367 11867
rect 11433 12136 11447 12150
rect 11993 12153 12007 12167
rect 11653 12136 11667 12150
rect 11693 12136 11707 12150
rect 11733 12136 11747 12150
rect 11773 12136 11787 12150
rect 12033 12136 12047 12150
rect 12073 12136 12087 12150
rect 12233 12136 12247 12150
rect 12333 12136 12347 12150
rect 11393 12053 11407 12067
rect 11453 12053 11467 12067
rect 11713 12090 11727 12104
rect 11653 11893 11667 11907
rect 11113 11836 11127 11850
rect 10953 11733 10967 11747
rect 10953 11616 10967 11630
rect 10953 11316 10967 11330
rect 11073 11753 11087 11767
rect 11053 11616 11067 11630
rect 11193 11773 11207 11787
rect 11033 11533 11047 11547
rect 11013 11273 11027 11287
rect 11073 11513 11087 11527
rect 11113 11353 11127 11367
rect 11093 11316 11107 11330
rect 11133 11316 11147 11330
rect 11113 11270 11127 11284
rect 11053 11253 11067 11267
rect 10953 11133 10967 11147
rect 10953 11096 10967 11110
rect 11013 11096 11027 11110
rect 11113 11173 11127 11187
rect 10953 11013 10967 11027
rect 10933 10733 10947 10747
rect 10833 10673 10847 10687
rect 10713 10353 10727 10367
rect 10793 10353 10807 10367
rect 10693 10333 10707 10347
rect 10693 10276 10707 10290
rect 10733 10276 10747 10290
rect 10773 10276 10787 10290
rect 10773 10153 10787 10167
rect 10713 10113 10727 10127
rect 10673 10056 10687 10070
rect 10893 10613 10907 10627
rect 10873 10530 10887 10544
rect 10913 10530 10927 10544
rect 10853 10413 10867 10427
rect 10833 10113 10847 10127
rect 10913 10493 10927 10507
rect 10873 10373 10887 10387
rect 11033 10973 11047 10987
rect 11013 10796 11027 10810
rect 10993 10673 11007 10687
rect 10973 10573 10987 10587
rect 10973 10530 10987 10544
rect 10953 10293 10967 10307
rect 10973 10213 10987 10227
rect 10953 10133 10967 10147
rect 10873 10113 10887 10127
rect 10853 10093 10867 10107
rect 10793 10053 10807 10067
rect 10713 9913 10727 9927
rect 10753 9913 10767 9927
rect 10613 9833 10627 9847
rect 10653 9756 10667 9770
rect 10713 9756 10727 9770
rect 10773 9756 10787 9770
rect 10773 9713 10787 9727
rect 10693 9693 10707 9707
rect 10753 9693 10767 9707
rect 10753 9653 10767 9667
rect 10693 9633 10707 9647
rect 10653 9613 10667 9627
rect 10693 9536 10707 9550
rect 10673 9490 10687 9504
rect 10853 9553 10867 9567
rect 10833 9533 10847 9547
rect 10613 9353 10627 9367
rect 10593 9233 10607 9247
rect 10713 9473 10727 9487
rect 10693 9313 10707 9327
rect 10673 9273 10687 9287
rect 10653 9236 10667 9250
rect 10633 9133 10647 9147
rect 10573 8893 10587 8907
rect 10673 8813 10687 8827
rect 10553 8753 10567 8767
rect 10653 8753 10667 8767
rect 10493 8716 10507 8730
rect 10613 8716 10627 8730
rect 10153 8633 10167 8647
rect 10273 8633 10287 8647
rect 10033 8513 10047 8527
rect 10073 8496 10087 8510
rect 10133 8493 10147 8507
rect 10013 8453 10027 8467
rect 10093 8433 10107 8447
rect 10053 8393 10067 8407
rect 10313 8513 10327 8527
rect 10393 8633 10407 8647
rect 10153 8433 10167 8447
rect 10093 8373 10107 8387
rect 10133 8373 10147 8387
rect 9933 8233 9947 8247
rect 9993 8233 10007 8247
rect 9853 8170 9867 8184
rect 9833 7993 9847 8007
rect 9893 8133 9907 8147
rect 9873 8053 9887 8067
rect 9833 7953 9847 7967
rect 9873 7950 9887 7964
rect 9713 7930 9727 7944
rect 9773 7913 9787 7927
rect 9573 7793 9587 7807
rect 9713 7793 9727 7807
rect 9593 7753 9607 7767
rect 9553 7676 9567 7690
rect 9373 7613 9387 7627
rect 9533 7613 9547 7627
rect 9353 7593 9367 7607
rect 9273 7553 9287 7567
rect 9173 7533 9187 7547
rect 9153 7493 9167 7507
rect 9193 7456 9207 7470
rect 9333 7493 9347 7507
rect 9353 7430 9367 7444
rect 9173 7410 9187 7424
rect 9113 7233 9127 7247
rect 9133 7156 9147 7170
rect 9173 7156 9187 7170
rect 9113 7110 9127 7124
rect 9153 7093 9167 7107
rect 9073 7073 9087 7087
rect 9133 7073 9147 7087
rect 9173 7073 9187 7087
rect 9053 6973 9067 6987
rect 9033 6933 9047 6947
rect 9073 6893 9087 6907
rect 9153 6936 9167 6950
rect 9013 6733 9027 6747
rect 9053 6713 9067 6727
rect 9093 6853 9107 6867
rect 8893 6616 8907 6630
rect 8973 6473 8987 6487
rect 8913 6453 8927 6467
rect 8833 6413 8847 6427
rect 8873 6416 8887 6430
rect 8753 6353 8767 6367
rect 8853 6373 8867 6387
rect 8933 6370 8947 6384
rect 9093 6593 9107 6607
rect 9053 6533 9067 6547
rect 9033 6416 9047 6430
rect 9033 6333 9047 6347
rect 8973 6233 8987 6247
rect 8853 6153 8867 6167
rect 8913 6153 8927 6167
rect 8833 6133 8847 6147
rect 8793 6116 8807 6130
rect 8873 6116 8887 6130
rect 8853 6070 8867 6084
rect 8793 5973 8807 5987
rect 8773 5793 8787 5807
rect 8753 5733 8767 5747
rect 8733 5653 8747 5667
rect 8693 5633 8707 5647
rect 8733 5596 8747 5610
rect 8713 5550 8727 5564
rect 8733 5533 8747 5547
rect 8713 5513 8727 5527
rect 8653 5473 8667 5487
rect 8633 5413 8647 5427
rect 8653 5376 8667 5390
rect 8633 5330 8647 5344
rect 8673 5253 8687 5267
rect 8753 5473 8767 5487
rect 8732 5233 8746 5247
rect 8753 5233 8767 5247
rect 8753 5193 8767 5207
rect 8753 5172 8767 5186
rect 8713 5153 8727 5167
rect 8593 5073 8607 5087
rect 8613 5076 8627 5090
rect 8693 5076 8707 5090
rect 8593 4933 8607 4947
rect 8573 4893 8587 4907
rect 8553 4856 8567 4870
rect 8453 4773 8467 4787
rect 8513 4773 8527 4787
rect 8493 4733 8507 4747
rect 8433 4613 8447 4627
rect 8493 4613 8507 4627
rect 8553 4793 8567 4807
rect 8533 4753 8547 4767
rect 8493 4573 8507 4587
rect 8473 4510 8487 4524
rect 8513 4493 8527 4507
rect 8433 4473 8447 4487
rect 8513 4393 8527 4407
rect 8473 4373 8487 4387
rect 8433 4273 8447 4287
rect 8413 4253 8427 4267
rect 8413 4193 8427 4207
rect 8393 4053 8407 4067
rect 8373 4036 8387 4050
rect 8493 4290 8507 4304
rect 8573 4553 8587 4567
rect 8473 4253 8487 4267
rect 8453 4133 8467 4147
rect 8313 3993 8327 4007
rect 8353 3973 8367 3987
rect 8333 3873 8347 3887
rect 8313 3853 8327 3867
rect 8333 3773 8347 3787
rect 8313 3673 8327 3687
rect 8333 3493 8347 3507
rect 8313 3293 8327 3307
rect 8313 3253 8327 3267
rect 8453 3933 8467 3947
rect 8453 3853 8467 3867
rect 8413 3816 8427 3830
rect 8513 4053 8527 4067
rect 8473 3833 8487 3847
rect 8533 3973 8547 3987
rect 8573 4133 8587 4147
rect 8713 5030 8727 5044
rect 8753 5033 8767 5047
rect 8893 6033 8907 6047
rect 8933 5913 8947 5927
rect 8853 5896 8867 5910
rect 8813 5753 8827 5767
rect 8793 5596 8807 5610
rect 8793 5493 8807 5507
rect 8873 5813 8887 5827
rect 8853 5553 8867 5567
rect 8893 5673 8907 5687
rect 8893 5633 8907 5647
rect 8893 5533 8907 5547
rect 8813 5473 8827 5487
rect 8833 5413 8847 5427
rect 8813 5373 8827 5387
rect 8813 5313 8827 5327
rect 8813 5253 8827 5267
rect 8793 5193 8807 5207
rect 8813 5013 8827 5027
rect 8953 5850 8967 5864
rect 9133 6733 9147 6747
rect 9233 7413 9247 7427
rect 9353 7393 9367 7407
rect 9273 7293 9287 7307
rect 9233 7156 9247 7170
rect 9253 7133 9267 7147
rect 9253 6893 9267 6907
rect 9213 6813 9227 6827
rect 9233 6773 9247 6787
rect 9193 6733 9207 6747
rect 9173 6573 9187 6587
rect 9153 6533 9167 6547
rect 9113 6473 9127 6487
rect 9073 6453 9087 6467
rect 9153 6416 9167 6430
rect 9253 6713 9267 6727
rect 9253 6673 9267 6687
rect 9233 6616 9247 6630
rect 9173 6353 9187 6367
rect 9133 6293 9147 6307
rect 9153 6173 9167 6187
rect 9093 6133 9107 6147
rect 9213 6116 9227 6130
rect 9133 6053 9147 6067
rect 9173 6053 9187 6067
rect 9073 5953 9087 5967
rect 9113 5913 9127 5927
rect 9113 5850 9127 5864
rect 9213 6033 9227 6047
rect 9573 7533 9587 7547
rect 9393 7473 9407 7487
rect 9533 7430 9547 7444
rect 9753 7713 9767 7727
rect 9673 7673 9687 7687
rect 9733 7533 9747 7547
rect 9673 7433 9687 7447
rect 9393 7393 9407 7407
rect 9693 7353 9707 7367
rect 9373 7273 9387 7287
rect 9413 7273 9427 7287
rect 9873 7833 9887 7847
rect 9833 7676 9847 7690
rect 9833 7613 9847 7627
rect 9813 7493 9827 7507
rect 9773 7473 9787 7487
rect 9793 7433 9807 7447
rect 9813 7373 9827 7387
rect 9753 7353 9767 7367
rect 9853 7513 9867 7527
rect 9853 7453 9867 7467
rect 9833 7293 9847 7307
rect 9573 7233 9587 7247
rect 9733 7233 9747 7247
rect 10053 8170 10067 8184
rect 9993 8133 10007 8147
rect 10473 8593 10487 8607
rect 10473 8533 10487 8547
rect 10453 8513 10467 8527
rect 10813 9453 10827 9467
rect 10773 9393 10787 9407
rect 10753 9233 10767 9247
rect 10753 8813 10767 8827
rect 10513 8670 10527 8684
rect 10593 8670 10607 8684
rect 10493 8393 10507 8407
rect 10473 8353 10487 8367
rect 10453 8313 10467 8327
rect 10433 8233 10447 8247
rect 10413 8216 10427 8230
rect 10253 8176 10267 8190
rect 9953 8093 9967 8107
rect 10093 8093 10107 8107
rect 10293 8073 10307 8087
rect 9913 8053 9927 8067
rect 10093 8053 10107 8067
rect 10053 7950 10067 7964
rect 10173 7956 10187 7970
rect 10253 7953 10267 7967
rect 10213 7893 10227 7907
rect 10213 7713 10227 7727
rect 10073 7676 10087 7690
rect 10113 7676 10127 7690
rect 10153 7673 10167 7687
rect 9893 7613 9907 7627
rect 9953 7593 9967 7607
rect 10053 7593 10067 7607
rect 9913 7573 9927 7587
rect 10053 7493 10067 7507
rect 9993 7456 10007 7470
rect 10113 7513 10127 7527
rect 10093 7430 10107 7444
rect 10313 8033 10327 8047
rect 10393 8173 10407 8187
rect 10473 8073 10487 8087
rect 10433 7993 10447 8007
rect 10673 8670 10687 8684
rect 10733 8670 10747 8684
rect 10653 8593 10667 8607
rect 10533 8553 10547 8567
rect 10633 8553 10647 8567
rect 10613 8496 10627 8510
rect 10713 8553 10727 8567
rect 10633 8433 10647 8447
rect 10553 8233 10567 8247
rect 10533 8153 10547 8167
rect 10533 8013 10547 8027
rect 10513 7953 10527 7967
rect 10393 7893 10407 7907
rect 10453 7833 10467 7847
rect 10333 7733 10347 7747
rect 10313 7673 10327 7687
rect 10373 7693 10387 7707
rect 10293 7633 10307 7647
rect 10353 7630 10367 7644
rect 10313 7430 10327 7444
rect 10533 7753 10547 7767
rect 10513 7733 10527 7747
rect 10493 7673 10507 7687
rect 10513 7593 10527 7607
rect 9973 7410 9987 7424
rect 10153 7410 10167 7424
rect 9873 7213 9887 7227
rect 9893 7176 9907 7190
rect 9353 7130 9367 7144
rect 9533 7130 9547 7144
rect 9573 7136 9587 7150
rect 9733 7136 9747 7150
rect 9953 7176 9967 7190
rect 9853 7130 9867 7144
rect 9933 7133 9947 7147
rect 9493 7093 9507 7107
rect 9433 7073 9447 7087
rect 9473 7073 9487 7087
rect 9493 7053 9507 7067
rect 9533 7053 9547 7067
rect 10013 7373 10027 7387
rect 9993 7213 10007 7227
rect 9973 7053 9987 7067
rect 9813 7033 9827 7047
rect 9953 7033 9967 7047
rect 9473 7013 9487 7027
rect 9513 7013 9527 7027
rect 9613 7013 9627 7027
rect 9673 7013 9687 7027
rect 9433 6993 9447 7007
rect 9373 6973 9387 6987
rect 9313 6936 9327 6950
rect 9333 6890 9347 6904
rect 9413 6853 9427 6867
rect 9373 6753 9387 6767
rect 9313 6673 9327 6687
rect 9273 6633 9287 6647
rect 9373 6613 9387 6627
rect 9333 6590 9347 6604
rect 9293 6533 9307 6547
rect 9413 6533 9427 6547
rect 9473 6713 9487 6727
rect 9493 6636 9507 6650
rect 9493 6513 9507 6527
rect 9793 6936 9807 6950
rect 9793 6893 9807 6907
rect 9913 6953 9927 6967
rect 9873 6936 9887 6950
rect 9853 6853 9867 6867
rect 9933 6890 9947 6904
rect 9893 6793 9907 6807
rect 9653 6713 9667 6727
rect 9813 6713 9827 6727
rect 9553 6673 9567 6687
rect 9953 6653 9967 6667
rect 9613 6636 9627 6650
rect 9693 6610 9707 6624
rect 9813 6616 9827 6630
rect 9553 6573 9567 6587
rect 9433 6453 9447 6467
rect 9473 6453 9487 6467
rect 10033 7273 10047 7287
rect 10013 7013 10027 7027
rect 9993 6890 10007 6904
rect 10513 7393 10527 7407
rect 10473 7353 10487 7367
rect 10153 7233 10167 7247
rect 10493 7233 10507 7247
rect 10133 7156 10147 7170
rect 10373 7156 10387 7170
rect 10413 7156 10427 7170
rect 10333 7133 10347 7147
rect 10213 7033 10227 7047
rect 10213 6953 10227 6967
rect 10273 6953 10287 6967
rect 10113 6936 10127 6950
rect 10173 6936 10187 6950
rect 10093 6753 10107 6767
rect 10093 6693 10107 6707
rect 10033 6653 10047 6667
rect 9973 6610 9987 6624
rect 10013 6610 10027 6624
rect 9953 6573 9967 6587
rect 9993 6533 10007 6547
rect 9833 6513 9847 6527
rect 9953 6513 9967 6527
rect 9653 6453 9667 6467
rect 9493 6433 9507 6447
rect 9553 6433 9567 6447
rect 9593 6433 9607 6447
rect 9453 6416 9467 6430
rect 9433 6370 9447 6384
rect 9273 6353 9287 6367
rect 9433 6353 9447 6367
rect 9253 6013 9267 6027
rect 9233 5933 9247 5947
rect 9193 5896 9207 5910
rect 9053 5813 9067 5827
rect 8933 5613 8947 5627
rect 8973 5613 8987 5627
rect 9013 5596 9027 5610
rect 9173 5850 9187 5864
rect 9573 6353 9587 6367
rect 9473 6193 9487 6207
rect 9493 6153 9507 6167
rect 9393 6116 9407 6130
rect 9453 6116 9467 6130
rect 9413 5933 9427 5947
rect 9533 6033 9547 6047
rect 9573 5896 9587 5910
rect 9633 6293 9647 6307
rect 9513 5850 9527 5864
rect 9273 5813 9287 5827
rect 9533 5813 9547 5827
rect 9213 5793 9227 5807
rect 9513 5713 9527 5727
rect 9513 5593 9527 5607
rect 8993 5533 9007 5547
rect 9053 5533 9067 5547
rect 8953 5493 8967 5507
rect 8933 5413 8947 5427
rect 8913 5393 8927 5407
rect 8893 5376 8907 5390
rect 9093 5376 9107 5390
rect 8993 5353 9007 5367
rect 8853 5330 8867 5344
rect 8673 4973 8687 4987
rect 8773 4973 8787 4987
rect 8833 4973 8847 4987
rect 8693 4856 8707 4870
rect 8613 4773 8627 4787
rect 8673 4673 8687 4687
rect 8633 4473 8647 4487
rect 8633 4413 8647 4427
rect 8613 4393 8627 4407
rect 8633 4373 8647 4387
rect 8613 4333 8627 4347
rect 8633 4273 8647 4287
rect 8653 4253 8667 4267
rect 8653 4173 8667 4187
rect 8613 4153 8627 4167
rect 8513 3773 8527 3787
rect 8373 3753 8387 3767
rect 8433 3753 8447 3767
rect 8413 3633 8427 3647
rect 8553 3816 8567 3830
rect 8553 3713 8567 3727
rect 8413 3573 8427 3587
rect 8453 3573 8467 3587
rect 8533 3573 8547 3587
rect 8553 3513 8567 3527
rect 8513 3470 8527 3484
rect 8553 3470 8567 3484
rect 8413 3373 8427 3387
rect 8473 3373 8487 3387
rect 8453 3296 8467 3310
rect 8493 3296 8507 3310
rect 8433 3250 8447 3264
rect 8633 4133 8647 4147
rect 8613 4033 8627 4047
rect 8713 4613 8727 4627
rect 8693 4373 8707 4387
rect 8813 4953 8827 4967
rect 8853 4933 8867 4947
rect 8813 4893 8827 4907
rect 8793 4873 8807 4887
rect 8833 4856 8847 4870
rect 8773 4810 8787 4824
rect 8853 4810 8867 4824
rect 8913 5330 8927 5344
rect 8953 5313 8967 5327
rect 9013 5253 9027 5267
rect 8993 5153 9007 5167
rect 9013 5133 9027 5147
rect 8953 5076 8967 5090
rect 8993 5076 9007 5090
rect 9033 5076 9047 5090
rect 8893 5053 8907 5067
rect 8753 4773 8767 4787
rect 8793 4773 8807 4787
rect 8833 4773 8847 4787
rect 8873 4773 8887 4787
rect 8733 4553 8747 4567
rect 8813 4733 8827 4747
rect 8773 4510 8787 4524
rect 8813 4373 8827 4387
rect 8693 4290 8707 4304
rect 8673 4153 8687 4167
rect 8753 4273 8767 4287
rect 8793 4273 8807 4287
rect 8733 4253 8747 4267
rect 8713 4133 8727 4147
rect 8713 4093 8727 4107
rect 8693 4073 8707 4087
rect 8593 3953 8607 3967
rect 8593 3873 8607 3887
rect 8673 3990 8687 4004
rect 8713 3953 8727 3967
rect 8653 3833 8667 3847
rect 8633 3773 8647 3787
rect 8593 3373 8607 3387
rect 8733 3873 8747 3887
rect 8793 4233 8807 4247
rect 8913 5033 8927 5047
rect 8913 4933 8927 4947
rect 8973 5030 8987 5044
rect 9093 5033 9107 5047
rect 9313 5576 9327 5590
rect 9433 5570 9447 5584
rect 9313 5473 9327 5487
rect 9373 5473 9387 5487
rect 9173 5413 9187 5427
rect 9213 5376 9227 5390
rect 9113 5013 9127 5027
rect 9033 4993 9047 5007
rect 9093 4973 9107 4987
rect 9093 4893 9107 4907
rect 9113 4873 9127 4887
rect 8933 4856 8947 4870
rect 8973 4853 8987 4867
rect 9073 4856 9087 4870
rect 8933 4813 8947 4827
rect 9053 4810 9067 4824
rect 8913 4793 8927 4807
rect 9053 4773 9067 4787
rect 8933 4753 8947 4767
rect 9033 4753 9047 4767
rect 8893 4733 8907 4747
rect 8873 4713 8887 4727
rect 8853 4653 8867 4667
rect 8873 4633 8887 4647
rect 8853 4510 8867 4524
rect 8833 4173 8847 4187
rect 8793 4153 8807 4167
rect 8813 4093 8827 4107
rect 8793 3953 8807 3967
rect 8713 3816 8727 3830
rect 8793 3816 8807 3830
rect 8733 3733 8747 3747
rect 8753 3516 8767 3530
rect 8713 3470 8727 3484
rect 8773 3470 8787 3484
rect 8593 3293 8607 3307
rect 8653 3293 8667 3307
rect 8713 3296 8727 3310
rect 8513 3233 8527 3247
rect 8573 3233 8587 3247
rect 8353 3213 8367 3227
rect 8293 3033 8307 3047
rect 8373 3033 8387 3047
rect 8413 3033 8427 3047
rect 8213 3013 8227 3027
rect 8253 2996 8267 3010
rect 8293 2996 8307 3010
rect 8333 2996 8347 3010
rect 8313 2913 8327 2927
rect 8353 2893 8367 2907
rect 8253 2853 8267 2867
rect 8253 2793 8267 2807
rect 8293 2776 8307 2790
rect 8273 2730 8287 2744
rect 8233 2693 8247 2707
rect 8253 2476 8267 2490
rect 8273 2353 8287 2367
rect 8353 2353 8367 2367
rect 8273 2293 8287 2307
rect 8213 2256 8227 2270
rect 8393 2776 8407 2790
rect 8473 2996 8487 3010
rect 8432 2853 8446 2867
rect 8453 2853 8467 2867
rect 8433 2773 8447 2787
rect 8413 2730 8427 2744
rect 8433 2693 8447 2707
rect 8413 2573 8427 2587
rect 8393 2393 8407 2407
rect 8213 2193 8227 2207
rect 8253 2193 8267 2207
rect 8433 2493 8447 2507
rect 8433 2373 8447 2387
rect 8433 2352 8447 2366
rect 8433 2233 8447 2247
rect 8193 2173 8207 2187
rect 8293 2173 8307 2187
rect 8413 2173 8427 2187
rect 8173 2153 8187 2167
rect 8273 2153 8287 2167
rect 8193 2113 8207 2127
rect 8153 2033 8167 2047
rect 8153 1956 8167 1970
rect 8253 2033 8267 2047
rect 8113 1913 8127 1927
rect 8173 1910 8187 1924
rect 8213 1910 8227 1924
rect 8093 1873 8107 1887
rect 8153 1873 8167 1887
rect 8193 1813 8207 1827
rect 8193 1773 8207 1787
rect 8233 1773 8247 1787
rect 8072 1633 8086 1647
rect 8093 1633 8107 1647
rect 8233 1693 8247 1707
rect 8173 1593 8187 1607
rect 8213 1553 8227 1567
rect 8133 1473 8147 1487
rect 8013 1390 8027 1404
rect 8153 1353 8167 1367
rect 7973 1293 7987 1307
rect 8733 3250 8747 3264
rect 8613 3193 8627 3207
rect 8713 3173 8727 3187
rect 8553 2996 8567 3010
rect 8633 2996 8647 3010
rect 8513 2953 8527 2967
rect 8573 2950 8587 2964
rect 8573 2833 8587 2847
rect 8653 2833 8667 2847
rect 8533 2776 8547 2790
rect 8553 2730 8567 2744
rect 8613 2730 8627 2744
rect 8513 2673 8527 2687
rect 8533 2533 8547 2547
rect 8573 2476 8587 2490
rect 8453 2093 8467 2107
rect 8453 2033 8467 2047
rect 8313 1956 8327 1970
rect 8413 1956 8427 1970
rect 8453 1956 8467 1970
rect 8293 1773 8307 1787
rect 8273 1673 8287 1687
rect 8513 2393 8527 2407
rect 8573 2413 8587 2427
rect 8553 2333 8567 2347
rect 8533 2256 8547 2270
rect 8593 2353 8607 2367
rect 8593 2256 8607 2270
rect 8553 2173 8567 2187
rect 8613 2113 8627 2127
rect 8593 1956 8607 1970
rect 8493 1913 8507 1927
rect 8573 1873 8587 1887
rect 8433 1833 8447 1847
rect 8433 1773 8447 1787
rect 8373 1736 8387 1750
rect 8473 1736 8487 1750
rect 8513 1736 8527 1750
rect 8313 1593 8327 1607
rect 8253 1513 8267 1527
rect 8353 1573 8367 1587
rect 8273 1390 8287 1404
rect 8353 1390 8367 1404
rect 8213 1333 8227 1347
rect 7953 1213 7967 1227
rect 8073 1216 8087 1230
rect 8153 1216 8167 1230
rect 8293 1216 8307 1230
rect 7933 1173 7947 1187
rect 8053 1170 8067 1184
rect 8093 1170 8107 1184
rect 7973 1113 7987 1127
rect 7953 1073 7967 1087
rect 7973 1053 7987 1067
rect 8213 1073 8227 1087
rect 8413 1690 8427 1704
rect 8393 1673 8407 1687
rect 8453 1593 8467 1607
rect 8413 1553 8427 1567
rect 8473 1513 8487 1527
rect 8393 1393 8407 1407
rect 8453 1170 8467 1184
rect 8373 1073 8387 1087
rect 8053 1033 8067 1047
rect 8213 1033 8227 1047
rect 8333 1033 8347 1047
rect 8413 1033 8427 1047
rect 7913 1013 7927 1027
rect 7893 933 7907 947
rect 8093 953 8107 967
rect 8413 953 8427 967
rect 8093 913 8107 927
rect 7993 890 8007 904
rect 7873 733 7887 747
rect 7873 693 7887 707
rect 7853 633 7867 647
rect 7953 853 7967 867
rect 7933 793 7947 807
rect 7893 613 7907 627
rect 8253 896 8267 910
rect 8373 890 8387 904
rect 8413 873 8427 887
rect 8453 873 8467 887
rect 8053 833 8067 847
rect 7953 773 7967 787
rect 7993 753 8007 767
rect 7953 693 7967 707
rect 8293 733 8307 747
rect 8033 696 8047 710
rect 8333 696 8347 710
rect 7933 533 7947 547
rect 7913 396 7927 410
rect 8053 633 8067 647
rect 8013 553 8027 567
rect 8433 813 8447 827
rect 8353 613 8367 627
rect 8413 613 8427 627
rect 8453 773 8467 787
rect 8453 653 8467 667
rect 8433 573 8447 587
rect 8313 493 8327 507
rect 8512 1473 8526 1487
rect 8533 1473 8547 1487
rect 8533 1433 8547 1447
rect 8673 2313 8687 2327
rect 8653 2213 8667 2227
rect 8793 3433 8807 3447
rect 8793 3293 8807 3307
rect 8793 3250 8807 3264
rect 8833 3893 8847 3907
rect 8833 3693 8847 3707
rect 9013 4713 9027 4727
rect 8953 4693 8967 4707
rect 8953 4553 8967 4567
rect 8993 4556 9007 4570
rect 9113 4793 9127 4807
rect 9093 4633 9107 4647
rect 9073 4556 9087 4570
rect 8973 4510 8987 4524
rect 9013 4510 9027 4524
rect 9093 4513 9107 4527
rect 9073 4473 9087 4487
rect 8873 4413 8887 4427
rect 8933 4413 8947 4427
rect 9073 4353 9087 4367
rect 9033 4336 9047 4350
rect 9053 4293 9067 4307
rect 8993 4253 9007 4267
rect 8953 4233 8967 4247
rect 9013 4213 9027 4227
rect 9033 4193 9047 4207
rect 9013 4153 9027 4167
rect 8953 4133 8967 4147
rect 8953 4093 8967 4107
rect 8973 4073 8987 4087
rect 8933 4036 8947 4050
rect 9053 4113 9067 4127
rect 9033 4033 9047 4047
rect 9013 4013 9027 4027
rect 9093 4313 9107 4327
rect 9093 4173 9107 4187
rect 9093 4093 9107 4107
rect 8953 3973 8967 3987
rect 8913 3816 8927 3830
rect 8873 3733 8887 3747
rect 8893 3673 8907 3687
rect 8873 3333 8887 3347
rect 8893 3173 8907 3187
rect 8873 3153 8887 3167
rect 8853 3053 8867 3067
rect 8813 3033 8827 3047
rect 8833 2996 8847 3010
rect 8973 3816 8987 3830
rect 9013 3816 9027 3830
rect 8953 3773 8967 3787
rect 8953 3733 8967 3747
rect 8993 3733 9007 3747
rect 8993 3593 9007 3607
rect 8993 3553 9007 3567
rect 8933 3513 8947 3527
rect 8933 3470 8947 3484
rect 8973 3470 8987 3484
rect 8933 3353 8947 3367
rect 8993 3313 9007 3327
rect 8933 3293 8947 3307
rect 9033 3273 9047 3287
rect 8933 3253 8947 3267
rect 8773 2893 8787 2907
rect 8853 2913 8867 2927
rect 8913 2773 8927 2787
rect 8733 2673 8747 2687
rect 8773 2653 8787 2667
rect 8713 2633 8727 2647
rect 8753 2553 8767 2567
rect 8733 2533 8747 2547
rect 8693 2133 8707 2147
rect 8673 2053 8687 2067
rect 8873 2493 8887 2507
rect 8813 2413 8827 2427
rect 8853 2373 8867 2387
rect 8833 2256 8847 2270
rect 8793 2053 8807 2067
rect 8693 2033 8707 2047
rect 8753 2033 8767 2047
rect 8693 1956 8707 1970
rect 8713 1910 8727 1924
rect 8713 1853 8727 1867
rect 8653 1793 8667 1807
rect 8633 1673 8647 1687
rect 8753 1736 8767 1750
rect 8693 1673 8707 1687
rect 8733 1673 8747 1687
rect 8673 1613 8687 1627
rect 8613 1533 8627 1547
rect 8593 1493 8607 1507
rect 8613 1436 8627 1450
rect 8653 1436 8667 1450
rect 8553 1353 8567 1367
rect 8593 1216 8607 1230
rect 8513 1173 8527 1187
rect 8553 1173 8567 1187
rect 8513 953 8527 967
rect 8493 893 8507 907
rect 8513 813 8527 827
rect 8493 793 8507 807
rect 8533 773 8547 787
rect 8493 696 8507 710
rect 8473 553 8487 567
rect 8493 533 8507 547
rect 8473 433 8487 447
rect 8113 413 8127 427
rect 8433 416 8447 430
rect 7853 350 7867 364
rect 7893 350 7907 364
rect 8013 353 8027 367
rect 7933 313 7947 327
rect 8093 353 8107 367
rect 8093 313 8107 327
rect 7653 253 7667 267
rect 7833 253 7847 267
rect 8073 253 8087 267
rect 7653 173 7667 187
rect 6693 133 6707 147
rect 6633 53 6647 67
rect 7593 156 7607 170
rect 7693 150 7707 164
rect 7853 150 7867 164
rect 7973 156 7987 170
rect 8053 153 8067 167
rect 6773 130 6787 144
rect 6713 13 6727 27
rect 6773 13 6787 27
rect 7273 130 7287 144
rect 7513 130 7527 144
rect 8013 110 8027 124
rect 8273 376 8287 390
rect 8273 273 8287 287
rect 8173 253 8187 267
rect 8113 110 8127 124
rect 8253 130 8267 144
rect 8293 130 8307 144
rect 8573 1073 8587 1087
rect 8653 1073 8667 1087
rect 8573 993 8587 1007
rect 8633 953 8647 967
rect 8593 753 8607 767
rect 8553 693 8567 707
rect 8813 1956 8827 1970
rect 8853 2193 8867 2207
rect 8833 1853 8847 1867
rect 8953 3173 8967 3187
rect 8952 3053 8966 3067
rect 8973 3053 8987 3067
rect 8993 2933 9007 2947
rect 9013 2853 9027 2867
rect 9093 3993 9107 4007
rect 9093 3952 9107 3966
rect 9093 3453 9107 3467
rect 9073 3313 9087 3327
rect 9173 5293 9187 5307
rect 9193 5273 9207 5287
rect 9253 5113 9267 5127
rect 9213 5076 9227 5090
rect 9173 4873 9187 4887
rect 9273 5030 9287 5044
rect 9353 5413 9367 5427
rect 9193 4793 9207 4807
rect 9193 4753 9207 4767
rect 9173 4693 9187 4707
rect 9173 4672 9187 4686
rect 9193 4510 9207 4524
rect 9193 4433 9207 4447
rect 9193 4293 9207 4307
rect 9253 5013 9267 5027
rect 9233 4853 9247 4867
rect 9273 4953 9287 4967
rect 9233 4773 9247 4787
rect 9613 5850 9627 5864
rect 9613 5813 9627 5827
rect 9573 5793 9587 5807
rect 9553 5673 9567 5687
rect 9553 5493 9567 5507
rect 9533 5413 9547 5427
rect 9393 5376 9407 5390
rect 9433 5376 9447 5390
rect 9473 5330 9487 5344
rect 9393 5233 9407 5247
rect 9433 5233 9447 5247
rect 9413 5076 9427 5090
rect 9373 5033 9387 5047
rect 9393 4953 9407 4967
rect 9393 4913 9407 4927
rect 9413 4893 9427 4907
rect 9393 4856 9407 4870
rect 9313 4810 9327 4824
rect 9293 4773 9307 4787
rect 9373 4810 9387 4824
rect 9373 4773 9387 4787
rect 9353 4733 9367 4747
rect 9313 4673 9327 4687
rect 9333 4653 9347 4667
rect 9273 4593 9287 4607
rect 9273 4556 9287 4570
rect 9333 4556 9347 4570
rect 9253 4510 9267 4524
rect 9293 4510 9307 4524
rect 9353 4513 9367 4527
rect 9253 4433 9267 4447
rect 9333 4393 9347 4407
rect 9293 4336 9307 4350
rect 9273 4290 9287 4304
rect 9273 4233 9287 4247
rect 9213 4193 9227 4207
rect 9253 4133 9267 4147
rect 9213 4036 9227 4050
rect 9153 3953 9167 3967
rect 9193 3990 9207 4004
rect 9253 3953 9267 3967
rect 9193 3913 9207 3927
rect 9173 3873 9187 3887
rect 9133 3673 9147 3687
rect 9213 3873 9227 3887
rect 9193 3773 9207 3787
rect 9193 3752 9207 3766
rect 9193 3673 9207 3687
rect 9133 3613 9147 3627
rect 9173 3613 9187 3627
rect 9153 3513 9167 3527
rect 9133 3253 9147 3267
rect 9453 5213 9467 5227
rect 9433 4733 9447 4747
rect 9593 5376 9607 5390
rect 9593 5333 9607 5347
rect 9573 5293 9587 5307
rect 9473 5153 9487 5167
rect 9553 5153 9567 5167
rect 9593 5093 9607 5107
rect 9513 5076 9527 5090
rect 9553 5076 9567 5090
rect 9533 5030 9547 5044
rect 9593 4993 9607 5007
rect 9533 4973 9547 4987
rect 9713 6433 9727 6447
rect 9753 6416 9767 6430
rect 9733 6333 9747 6347
rect 9953 6416 9967 6430
rect 9913 6393 9927 6407
rect 9833 6313 9847 6327
rect 9773 6293 9787 6307
rect 9673 6253 9687 6267
rect 9653 5570 9667 5584
rect 9733 6116 9747 6130
rect 9773 6116 9787 6130
rect 9893 6116 9907 6130
rect 9893 6070 9907 6084
rect 9753 6013 9767 6027
rect 9713 5973 9727 5987
rect 9873 5953 9887 5967
rect 9793 5933 9807 5947
rect 9713 5896 9727 5910
rect 9833 5896 9847 5910
rect 9873 5896 9887 5910
rect 9773 5853 9787 5867
rect 9713 5613 9727 5627
rect 9773 5596 9787 5610
rect 9753 5550 9767 5564
rect 9793 5550 9807 5564
rect 9673 5473 9687 5487
rect 9733 5473 9747 5487
rect 9653 5453 9667 5467
rect 9693 5376 9707 5390
rect 9653 5330 9667 5344
rect 9753 5330 9767 5344
rect 9733 5293 9747 5307
rect 9793 5293 9807 5307
rect 9713 5233 9727 5247
rect 9633 5213 9647 5227
rect 9673 5113 9687 5127
rect 9633 5053 9647 5067
rect 9473 4793 9487 4807
rect 9473 4753 9487 4767
rect 9453 4633 9467 4647
rect 9393 4553 9407 4567
rect 9393 4433 9407 4447
rect 9433 4433 9447 4447
rect 9413 4413 9427 4427
rect 9373 4293 9387 4307
rect 9333 4213 9347 4227
rect 9353 4193 9367 4207
rect 9293 4113 9307 4127
rect 9333 4073 9347 4087
rect 9293 3990 9307 4004
rect 9333 3993 9347 4007
rect 9273 3873 9287 3887
rect 9293 3770 9307 3784
rect 9253 3693 9267 3707
rect 9253 3633 9267 3647
rect 9293 3516 9307 3530
rect 9433 4313 9447 4327
rect 9473 4336 9487 4350
rect 9513 4856 9527 4870
rect 9553 4933 9567 4947
rect 9573 4856 9587 4870
rect 9693 5076 9707 5090
rect 9673 5033 9687 5047
rect 9673 4856 9687 4870
rect 9553 4810 9567 4824
rect 9553 4713 9567 4727
rect 9533 4673 9547 4687
rect 9513 4573 9527 4587
rect 9613 4810 9627 4824
rect 9573 4693 9587 4707
rect 9553 4553 9567 4567
rect 9673 4593 9687 4607
rect 9593 4513 9607 4527
rect 9653 4513 9667 4527
rect 9533 4493 9547 4507
rect 9513 4353 9527 4367
rect 9553 4336 9567 4350
rect 9453 4233 9467 4247
rect 9433 4173 9447 4187
rect 9533 4290 9547 4304
rect 9473 4113 9487 4127
rect 9453 3990 9467 4004
rect 9413 3953 9427 3967
rect 9413 3913 9427 3927
rect 9413 3873 9427 3887
rect 9393 3816 9407 3830
rect 9373 3770 9387 3784
rect 9213 3413 9227 3427
rect 9253 3413 9267 3427
rect 9193 3296 9207 3310
rect 9333 3473 9347 3487
rect 9273 3353 9287 3367
rect 9313 3353 9327 3367
rect 9273 3313 9287 3327
rect 9173 3253 9187 3267
rect 9213 3250 9227 3264
rect 9253 3253 9267 3267
rect 9173 3213 9187 3227
rect 9233 3213 9247 3227
rect 9153 3053 9167 3067
rect 9113 3033 9127 3047
rect 9213 3033 9227 3047
rect 9153 2996 9167 3010
rect 9093 2950 9107 2964
rect 9053 2873 9067 2887
rect 9113 2853 9127 2867
rect 9033 2833 9047 2847
rect 9013 2793 9027 2807
rect 8993 2730 9007 2744
rect 8973 2653 8987 2667
rect 8993 2513 9007 2527
rect 8953 2253 8967 2267
rect 8933 2153 8947 2167
rect 8873 2133 8887 2147
rect 8853 1733 8867 1747
rect 8813 1613 8827 1627
rect 8793 1593 8807 1607
rect 9073 2776 9087 2790
rect 9153 2933 9167 2947
rect 9193 2873 9207 2887
rect 9153 2853 9167 2867
rect 9133 2793 9147 2807
rect 9053 2730 9067 2744
rect 9073 2713 9087 2727
rect 9073 2673 9087 2687
rect 9093 2653 9107 2667
rect 9153 2553 9167 2567
rect 9053 2533 9067 2547
rect 9093 2493 9107 2507
rect 9053 2476 9067 2490
rect 9053 2430 9067 2444
rect 9113 2430 9127 2444
rect 9093 2256 9107 2270
rect 9073 2173 9087 2187
rect 9092 2153 9106 2167
rect 9113 2153 9127 2167
rect 9013 2053 9027 2067
rect 9073 2013 9087 2027
rect 8973 1956 8987 1970
rect 8913 1793 8927 1807
rect 8893 1753 8907 1767
rect 9073 1913 9087 1927
rect 9053 1853 9067 1867
rect 8993 1753 9007 1767
rect 8913 1673 8927 1687
rect 8973 1673 8987 1687
rect 8893 1653 8907 1667
rect 8933 1653 8947 1667
rect 9033 1673 9047 1687
rect 9073 1753 9087 1767
rect 9073 1653 9087 1667
rect 8972 1633 8986 1647
rect 8993 1633 9007 1647
rect 9053 1633 9067 1647
rect 8953 1613 8967 1627
rect 8852 1553 8866 1567
rect 8873 1553 8887 1567
rect 8833 1533 8847 1547
rect 8833 1433 8847 1447
rect 8753 1393 8767 1407
rect 8693 1273 8707 1287
rect 8713 1253 8727 1267
rect 8813 1390 8827 1404
rect 8853 1353 8867 1367
rect 8813 1273 8827 1287
rect 8773 1213 8787 1227
rect 8813 1216 8827 1230
rect 8913 1293 8927 1307
rect 8773 1170 8787 1184
rect 8873 1170 8887 1184
rect 8833 1133 8847 1147
rect 8733 1113 8747 1127
rect 8713 1053 8727 1067
rect 8733 1033 8747 1047
rect 8733 915 8747 929
rect 8813 893 8827 907
rect 8713 853 8727 867
rect 8773 773 8787 787
rect 8693 697 8707 711
rect 8933 1216 8947 1230
rect 9173 2133 9187 2147
rect 9173 2093 9187 2107
rect 9173 2033 9187 2047
rect 9253 3153 9267 3167
rect 9253 3053 9267 3067
rect 9253 2996 9267 3010
rect 9313 3173 9327 3187
rect 9353 3373 9367 3387
rect 9533 3853 9547 3867
rect 9473 3816 9487 3830
rect 9533 3816 9547 3830
rect 9513 3753 9527 3767
rect 9473 3733 9487 3747
rect 9513 3713 9527 3727
rect 9553 3673 9567 3687
rect 9533 3633 9547 3647
rect 9473 3533 9487 3547
rect 9453 3473 9467 3487
rect 9533 3513 9547 3527
rect 9473 3453 9487 3467
rect 9513 3453 9527 3467
rect 9413 3413 9427 3427
rect 9493 3393 9507 3407
rect 9533 3433 9547 3447
rect 9613 4473 9627 4487
rect 9613 4393 9627 4407
rect 9593 3413 9607 3427
rect 9493 3353 9507 3367
rect 9533 3353 9547 3367
rect 9453 3296 9467 3310
rect 9493 3296 9507 3310
rect 9533 3296 9547 3310
rect 9373 3193 9387 3207
rect 9373 3153 9387 3167
rect 9533 3213 9547 3227
rect 9493 3193 9507 3207
rect 9493 3133 9507 3147
rect 9533 3133 9547 3147
rect 9473 3113 9487 3127
rect 9273 2913 9287 2927
rect 9253 2573 9267 2587
rect 9233 2433 9247 2447
rect 9413 2893 9427 2907
rect 9333 2853 9347 2867
rect 9313 2713 9327 2727
rect 9473 2713 9487 2727
rect 9273 2413 9287 2427
rect 9353 2573 9367 2587
rect 9473 2573 9487 2587
rect 9433 2493 9447 2507
rect 9373 2430 9387 2444
rect 9353 2413 9367 2427
rect 9413 2273 9427 2287
rect 9253 2073 9267 2087
rect 9213 2013 9227 2027
rect 9193 1956 9207 1970
rect 9173 1872 9187 1886
rect 9193 1853 9207 1867
rect 9393 2213 9407 2227
rect 9413 2193 9427 2207
rect 9373 2153 9387 2167
rect 9373 2093 9387 2107
rect 9313 1993 9327 2007
rect 9253 1956 9267 1970
rect 9293 1956 9307 1970
rect 9353 1956 9367 1970
rect 9213 1833 9227 1847
rect 9273 1910 9287 1924
rect 9313 1910 9327 1924
rect 9213 1690 9227 1704
rect 9173 1653 9187 1667
rect 9213 1633 9227 1647
rect 9453 2333 9467 2347
rect 9533 3093 9547 3107
rect 9653 4373 9667 4387
rect 9633 4336 9647 4350
rect 9653 4273 9667 4287
rect 9633 4253 9647 4267
rect 9713 4413 9727 4427
rect 9693 4273 9707 4287
rect 9693 4173 9707 4187
rect 9873 5853 9887 5867
rect 9873 5433 9887 5447
rect 9813 5193 9827 5207
rect 9853 5193 9867 5207
rect 9853 5133 9867 5147
rect 9833 5076 9847 5090
rect 9773 5030 9787 5044
rect 9813 5030 9827 5044
rect 9873 5030 9887 5044
rect 10013 6370 10027 6384
rect 9973 6333 9987 6347
rect 10053 6313 10067 6327
rect 9933 6233 9947 6247
rect 9993 6193 10007 6207
rect 10093 6173 10107 6187
rect 10073 6153 10087 6167
rect 9973 6070 9987 6084
rect 10013 6013 10027 6027
rect 9933 5933 9947 5947
rect 9913 5873 9927 5887
rect 9953 5793 9967 5807
rect 10093 6093 10107 6107
rect 10093 6033 10107 6047
rect 10153 6853 10167 6867
rect 10133 6793 10147 6807
rect 10233 6890 10247 6904
rect 10273 6890 10287 6904
rect 10233 6733 10247 6747
rect 10173 6673 10187 6687
rect 10153 6553 10167 6567
rect 10133 6333 10147 6347
rect 10133 6153 10147 6167
rect 10113 6013 10127 6027
rect 10053 5850 10067 5864
rect 10013 5753 10027 5767
rect 10033 5733 10047 5747
rect 10033 5613 10047 5627
rect 9993 5596 10007 5610
rect 10133 5813 10147 5827
rect 10093 5733 10107 5747
rect 10093 5693 10107 5707
rect 10053 5593 10067 5607
rect 10013 5550 10027 5564
rect 9973 5533 9987 5547
rect 9953 5513 9967 5527
rect 9933 5373 9947 5387
rect 9953 5053 9967 5067
rect 9773 4993 9787 5007
rect 9893 4993 9907 5007
rect 9953 4973 9967 4987
rect 9893 4953 9907 4967
rect 9893 4913 9907 4927
rect 9833 4893 9847 4907
rect 9873 4856 9887 4870
rect 9913 4856 9927 4870
rect 9933 4793 9947 4807
rect 10113 5593 10127 5607
rect 10113 5550 10127 5564
rect 10093 5513 10107 5527
rect 10033 5376 10047 5390
rect 10093 5376 10107 5390
rect 10013 5313 10027 5327
rect 9993 5233 10007 5247
rect 9993 5113 10007 5127
rect 9993 5053 10007 5067
rect 9913 4773 9927 4787
rect 9973 4773 9987 4787
rect 9893 4613 9907 4627
rect 9893 4553 9907 4567
rect 9773 4453 9787 4467
rect 9793 4433 9807 4447
rect 9733 4373 9747 4387
rect 9793 4336 9807 4350
rect 9773 4233 9787 4247
rect 9713 4153 9727 4167
rect 9673 4093 9687 4107
rect 9813 4093 9827 4107
rect 9693 4053 9707 4067
rect 9653 4033 9667 4047
rect 9733 4036 9747 4050
rect 9693 3853 9707 3867
rect 9653 3770 9667 3784
rect 9633 3753 9647 3767
rect 9613 3313 9627 3327
rect 9593 3233 9607 3247
rect 9673 3653 9687 3667
rect 9653 3553 9667 3567
rect 9653 3453 9667 3467
rect 9633 3093 9647 3107
rect 9753 3990 9767 4004
rect 9853 4452 9867 4466
rect 9873 4336 9887 4350
rect 9873 4153 9887 4167
rect 9833 3993 9847 4007
rect 9813 3816 9827 3830
rect 9853 3816 9867 3830
rect 9753 3770 9767 3784
rect 9793 3753 9807 3767
rect 9713 3633 9727 3647
rect 9893 3770 9907 3784
rect 9873 3713 9887 3727
rect 9853 3573 9867 3587
rect 9793 3533 9807 3547
rect 9833 3473 9847 3487
rect 9773 3393 9787 3407
rect 9813 3393 9827 3407
rect 9753 3313 9767 3327
rect 9713 3296 9727 3310
rect 9673 3253 9687 3267
rect 9773 3250 9787 3264
rect 9653 3013 9667 3027
rect 9713 3013 9727 3027
rect 9633 2996 9647 3010
rect 9733 2993 9747 3007
rect 9673 2950 9687 2964
rect 9713 2950 9727 2964
rect 9573 2913 9587 2927
rect 9613 2893 9627 2907
rect 9693 2813 9707 2827
rect 9633 2713 9647 2727
rect 9553 2613 9567 2627
rect 9493 2373 9507 2387
rect 9513 2210 9527 2224
rect 9633 2553 9647 2567
rect 9593 2473 9607 2487
rect 9713 2473 9727 2487
rect 9653 2430 9667 2444
rect 9693 2433 9707 2447
rect 9613 2413 9627 2427
rect 9613 2293 9627 2307
rect 9593 2210 9607 2224
rect 9513 2173 9527 2187
rect 9473 2093 9487 2107
rect 9433 2033 9447 2047
rect 9373 1713 9387 1727
rect 9253 1613 9267 1627
rect 9353 1613 9367 1627
rect 9193 1593 9207 1607
rect 9153 1433 9167 1447
rect 9053 1393 9067 1407
rect 9153 1333 9167 1347
rect 9153 1253 9167 1267
rect 8953 1173 8967 1187
rect 9093 1173 9107 1187
rect 9213 1213 9227 1227
rect 8933 1133 8947 1147
rect 9093 1133 9107 1147
rect 9193 1133 9207 1147
rect 9033 993 9047 1007
rect 8913 933 8927 947
rect 8833 853 8847 867
rect 8733 693 8747 707
rect 8813 693 8827 707
rect 8593 651 8607 665
rect 8673 433 8687 447
rect 8973 813 8987 827
rect 8933 753 8947 767
rect 9053 773 9067 787
rect 9033 697 9047 711
rect 8993 650 9007 664
rect 9033 633 9047 647
rect 8993 613 9007 627
rect 8753 553 8767 567
rect 8913 553 8927 567
rect 8953 553 8967 567
rect 9013 553 9027 567
rect 8693 350 8707 364
rect 8733 350 8747 364
rect 8913 433 8927 447
rect 8953 433 8967 447
rect 8933 350 8947 364
rect 9073 433 9087 447
rect 8473 153 8487 167
rect 9213 1073 9227 1087
rect 9193 1053 9207 1067
rect 9193 1013 9207 1027
rect 9433 1953 9447 1967
rect 9413 1693 9427 1707
rect 9613 2193 9627 2207
rect 9553 2173 9567 2187
rect 9533 1953 9547 1967
rect 9453 1910 9467 1924
rect 9513 1893 9527 1907
rect 9573 1893 9587 1907
rect 9513 1813 9527 1827
rect 9473 1753 9487 1767
rect 9473 1736 9487 1750
rect 9493 1690 9507 1704
rect 9533 1673 9547 1687
rect 9593 1833 9607 1847
rect 9593 1673 9607 1687
rect 9573 1573 9587 1587
rect 9493 1553 9507 1567
rect 9473 1493 9487 1507
rect 9433 1390 9447 1404
rect 9333 1253 9347 1267
rect 9373 1216 9387 1230
rect 9393 1133 9407 1147
rect 9353 1093 9367 1107
rect 9433 1093 9447 1107
rect 9293 1033 9307 1047
rect 9133 973 9147 987
rect 9233 973 9247 987
rect 9213 933 9227 947
rect 9353 915 9367 929
rect 9333 853 9347 867
rect 9393 773 9407 787
rect 9273 693 9287 707
rect 9193 613 9207 627
rect 9193 433 9207 447
rect 9173 396 9187 410
rect 9133 353 9147 367
rect 9093 313 9107 327
rect 9193 313 9207 327
rect 9213 193 9227 207
rect 9473 1053 9487 1067
rect 9473 733 9487 747
rect 9653 2133 9667 2147
rect 9633 2073 9647 2087
rect 9653 1913 9667 1927
rect 9673 1793 9687 1807
rect 9633 1736 9647 1750
rect 9673 1690 9687 1704
rect 9793 3153 9807 3167
rect 9833 3153 9847 3167
rect 9893 3633 9907 3647
rect 9873 3473 9887 3487
rect 9953 4493 9967 4507
rect 9933 4473 9947 4487
rect 9933 4290 9947 4304
rect 10093 5253 10107 5267
rect 10033 5233 10047 5247
rect 10032 5173 10046 5187
rect 10053 5173 10067 5187
rect 10033 5073 10047 5087
rect 10113 5153 10127 5167
rect 10233 6590 10247 6604
rect 10213 6453 10227 6467
rect 10393 7110 10407 7124
rect 10493 7110 10507 7124
rect 10333 6673 10347 6687
rect 10353 6636 10367 6650
rect 10333 6590 10347 6604
rect 10353 6573 10367 6587
rect 10333 6533 10347 6547
rect 10353 6513 10367 6527
rect 10333 6493 10347 6507
rect 10253 6433 10267 6447
rect 10293 6433 10307 6447
rect 10213 6370 10227 6384
rect 10273 6370 10287 6384
rect 10233 6333 10247 6347
rect 10193 6253 10207 6267
rect 10173 6233 10187 6247
rect 10173 5913 10187 5927
rect 10273 6193 10287 6207
rect 10293 6013 10307 6027
rect 10253 5913 10267 5927
rect 10193 5833 10207 5847
rect 10173 5313 10187 5327
rect 10373 6370 10387 6384
rect 10673 8393 10687 8407
rect 10593 7976 10607 7990
rect 10573 7953 10587 7967
rect 10613 7873 10627 7887
rect 10753 8493 10767 8507
rect 10753 8450 10767 8464
rect 10713 8013 10727 8027
rect 10733 7976 10747 7990
rect 10633 7793 10647 7807
rect 10693 7793 10707 7807
rect 10613 7676 10627 7690
rect 10653 7630 10667 7644
rect 10693 7630 10707 7644
rect 10593 7573 10607 7587
rect 10753 7613 10767 7627
rect 10673 7493 10687 7507
rect 10713 7493 10727 7507
rect 10593 7456 10607 7470
rect 10653 7456 10667 7470
rect 10573 7413 10587 7427
rect 10693 7456 10707 7470
rect 10653 7293 10667 7307
rect 10573 7273 10587 7287
rect 10573 7193 10587 7207
rect 10553 7156 10567 7170
rect 10513 7033 10527 7047
rect 10473 6993 10487 7007
rect 10633 7156 10647 7170
rect 10713 7410 10727 7424
rect 10693 7110 10707 7124
rect 10653 7033 10667 7047
rect 10693 6993 10707 7007
rect 10453 6853 10467 6867
rect 10473 6713 10487 6727
rect 10453 6653 10467 6667
rect 10433 6633 10447 6647
rect 10433 6533 10447 6547
rect 10413 6333 10427 6347
rect 10353 6033 10367 6047
rect 10373 5913 10387 5927
rect 10333 5896 10347 5910
rect 10313 5850 10327 5864
rect 10253 5733 10267 5747
rect 10213 5593 10227 5607
rect 10253 5596 10267 5610
rect 10193 5153 10207 5167
rect 10193 5093 10207 5107
rect 10073 4933 10087 4947
rect 10073 4653 10087 4667
rect 10053 4433 10067 4447
rect 9993 4336 10007 4350
rect 10093 4336 10107 4350
rect 9973 4193 9987 4207
rect 9953 4093 9967 4107
rect 9933 3993 9947 4007
rect 10033 4290 10047 4304
rect 10073 4253 10087 4267
rect 10052 4233 10066 4247
rect 9973 4036 9987 4050
rect 9993 4053 10007 4067
rect 10033 4036 10047 4050
rect 10113 4193 10127 4207
rect 10013 3990 10027 4004
rect 10053 3990 10067 4004
rect 10093 3990 10107 4004
rect 9993 3953 10007 3967
rect 10033 3953 10047 3967
rect 10113 3953 10127 3967
rect 9993 3853 10007 3867
rect 9953 3833 9967 3847
rect 10073 3816 10087 3830
rect 9913 3193 9927 3207
rect 9833 3053 9847 3067
rect 10053 3770 10067 3784
rect 10273 5513 10287 5527
rect 10273 5413 10287 5427
rect 10293 5330 10307 5344
rect 10253 5273 10267 5287
rect 10273 5253 10287 5267
rect 10213 4873 10227 4887
rect 10253 4873 10267 4887
rect 10153 4793 10167 4807
rect 10193 4773 10207 4787
rect 10173 4573 10187 4587
rect 10153 4510 10167 4524
rect 10153 4373 10167 4387
rect 10173 4333 10187 4347
rect 10153 4193 10167 4207
rect 10173 3833 10187 3847
rect 10153 3770 10167 3784
rect 10053 3733 10067 3747
rect 10013 3673 10027 3687
rect 10113 3693 10127 3707
rect 10093 3516 10107 3530
rect 10013 3473 10027 3487
rect 10073 3470 10087 3484
rect 10093 3453 10107 3467
rect 10033 3296 10047 3310
rect 9993 3233 10007 3247
rect 9953 3133 9967 3147
rect 9893 3033 9907 3047
rect 9933 3033 9947 3047
rect 9793 2950 9807 2964
rect 9853 2913 9867 2927
rect 9773 2893 9787 2907
rect 9953 2950 9967 2964
rect 10053 3233 10067 3247
rect 10013 2973 10027 2987
rect 9993 2873 10007 2887
rect 9913 2813 9927 2827
rect 9893 2776 9907 2790
rect 9773 2730 9787 2744
rect 9873 2730 9887 2744
rect 9733 2233 9747 2247
rect 9713 1953 9727 1967
rect 9633 1593 9647 1607
rect 9693 1593 9707 1607
rect 9713 1453 9727 1467
rect 9593 1390 9607 1404
rect 9633 1353 9647 1367
rect 9613 1293 9627 1307
rect 9613 1253 9627 1267
rect 9653 1093 9667 1107
rect 9673 1013 9687 1027
rect 9633 973 9647 987
rect 9653 870 9667 884
rect 9613 853 9627 867
rect 9573 813 9587 827
rect 9513 713 9527 727
rect 9693 713 9707 727
rect 9573 673 9587 687
rect 9433 650 9447 664
rect 9493 650 9507 664
rect 9853 2693 9867 2707
rect 9913 2593 9927 2607
rect 9893 2533 9907 2547
rect 9973 2430 9987 2444
rect 9873 2373 9887 2387
rect 9853 2293 9867 2307
rect 9793 2256 9807 2270
rect 9833 2256 9847 2270
rect 9953 2353 9967 2367
rect 9933 2273 9947 2287
rect 9773 2193 9787 2207
rect 9773 2172 9787 2186
rect 9853 2173 9867 2187
rect 9793 2073 9807 2087
rect 9893 2013 9907 2027
rect 9813 1956 9827 1970
rect 9873 1956 9887 1970
rect 9793 1910 9807 1924
rect 9813 1813 9827 1827
rect 9773 1736 9787 1750
rect 9793 1690 9807 1704
rect 9893 1833 9907 1847
rect 9893 1733 9907 1747
rect 9833 1633 9847 1647
rect 9813 1553 9827 1567
rect 9853 1553 9867 1567
rect 9753 1313 9767 1327
rect 9733 853 9747 867
rect 9713 693 9727 707
rect 9873 1533 9887 1547
rect 10033 2873 10047 2887
rect 10013 2413 10027 2427
rect 9973 2333 9987 2347
rect 9953 2213 9967 2227
rect 9933 2173 9947 2187
rect 9933 1873 9947 1887
rect 9953 1736 9967 1750
rect 9933 1713 9947 1727
rect 9953 1633 9967 1647
rect 9953 1612 9967 1626
rect 9913 1453 9927 1467
rect 9853 1373 9867 1387
rect 9893 1353 9907 1367
rect 9913 1273 9927 1287
rect 9833 1216 9847 1230
rect 9873 1216 9887 1230
rect 9813 1153 9827 1167
rect 9913 1153 9927 1167
rect 9893 1133 9907 1147
rect 10073 3193 10087 3207
rect 10053 2353 10067 2367
rect 9993 2193 10007 2207
rect 10033 2073 10047 2087
rect 10113 3233 10127 3247
rect 10413 5793 10427 5807
rect 10393 5330 10407 5344
rect 10353 5253 10367 5267
rect 10293 5193 10307 5207
rect 10533 6890 10547 6904
rect 10573 6890 10587 6904
rect 10673 6773 10687 6787
rect 10593 6653 10607 6667
rect 10533 6636 10547 6650
rect 10573 6636 10587 6650
rect 10633 6636 10647 6650
rect 10533 6593 10547 6607
rect 10593 6593 10607 6607
rect 10493 6573 10507 6587
rect 10533 6513 10547 6527
rect 10473 6370 10487 6384
rect 10553 6370 10567 6384
rect 10553 6070 10567 6084
rect 10513 6053 10527 6067
rect 10493 5893 10507 5907
rect 10493 5673 10507 5687
rect 10453 5633 10467 5647
rect 10673 6593 10687 6607
rect 10613 6453 10627 6467
rect 10993 10093 11007 10107
rect 11073 10893 11087 10907
rect 11073 10796 11087 10810
rect 11313 11836 11327 11850
rect 11413 11833 11427 11847
rect 11633 11836 11647 11850
rect 11333 11790 11347 11804
rect 11393 11793 11407 11807
rect 11693 11790 11707 11804
rect 11593 11773 11607 11787
rect 11413 11693 11427 11707
rect 11473 11693 11487 11707
rect 11233 11616 11247 11630
rect 11293 11616 11307 11630
rect 11333 11616 11347 11630
rect 11213 11213 11227 11227
rect 11213 11133 11227 11147
rect 11193 10813 11207 10827
rect 11033 10453 11047 10467
rect 11033 10393 11047 10407
rect 11013 10073 11027 10087
rect 10933 9973 10947 9987
rect 10993 9933 11007 9947
rect 10973 9913 10987 9927
rect 10973 9773 10987 9787
rect 10933 9756 10947 9770
rect 10913 9710 10927 9724
rect 10913 9573 10927 9587
rect 10873 9536 10887 9550
rect 10853 9453 10867 9467
rect 10833 9393 10847 9407
rect 10873 9313 10887 9327
rect 10953 9536 10967 9550
rect 11013 9733 11027 9747
rect 11013 9573 11027 9587
rect 10973 9413 10987 9427
rect 10933 9373 10947 9387
rect 10913 9272 10927 9286
rect 10893 9190 10907 9204
rect 10853 9173 10867 9187
rect 10813 8793 10827 8807
rect 10813 7693 10827 7707
rect 10853 9016 10867 9030
rect 10993 9253 11007 9267
rect 10993 9190 11007 9204
rect 10953 9133 10967 9147
rect 10953 9093 10967 9107
rect 10913 9016 10927 9030
rect 10953 9016 10967 9030
rect 10853 8873 10867 8887
rect 10873 8753 10887 8767
rect 10933 8753 10947 8767
rect 10913 8716 10927 8730
rect 10953 8716 10967 8730
rect 11013 8716 11027 8730
rect 10973 8653 10987 8667
rect 10933 8553 10947 8567
rect 10993 8553 11007 8567
rect 10873 8496 10887 8510
rect 10893 8433 10907 8447
rect 10993 8433 11007 8447
rect 10993 8333 11007 8347
rect 10873 8313 10887 8327
rect 10913 8233 10927 8247
rect 10953 8196 10967 8210
rect 10933 8113 10947 8127
rect 10893 8093 10907 8107
rect 10893 7993 10907 8007
rect 10913 7973 10927 7987
rect 11013 7973 11027 7987
rect 10873 7930 10887 7944
rect 10953 7930 10967 7944
rect 10993 7853 11007 7867
rect 10913 7693 10927 7707
rect 10973 7693 10987 7707
rect 10893 7676 10907 7690
rect 11013 7673 11027 7687
rect 10913 7630 10927 7644
rect 10973 7630 10987 7644
rect 10873 7613 10887 7627
rect 10833 7573 10847 7587
rect 10893 7553 10907 7567
rect 10873 7456 10887 7470
rect 10853 7253 10867 7267
rect 10793 7193 10807 7207
rect 10833 7173 10847 7187
rect 10793 7033 10807 7047
rect 10773 6953 10787 6967
rect 10713 6935 10727 6949
rect 10753 6935 10767 6949
rect 10693 6253 10707 6267
rect 10693 6193 10707 6207
rect 10613 6173 10627 6187
rect 10673 6053 10687 6067
rect 10533 5973 10547 5987
rect 10592 5973 10606 5987
rect 10613 5973 10627 5987
rect 10593 5913 10607 5927
rect 10533 5833 10547 5847
rect 10633 5850 10647 5864
rect 10613 5833 10627 5847
rect 10573 5793 10587 5807
rect 10453 5333 10467 5347
rect 10453 5233 10467 5247
rect 10333 5076 10347 5090
rect 10393 5076 10407 5090
rect 10433 5072 10447 5086
rect 10293 4773 10307 4787
rect 10533 5550 10547 5564
rect 10513 5473 10527 5487
rect 10553 5376 10567 5390
rect 10593 5376 10607 5390
rect 10533 5330 10547 5344
rect 10533 5293 10547 5307
rect 10593 5293 10607 5307
rect 10473 5213 10487 5227
rect 10513 5153 10527 5167
rect 10493 5113 10507 5127
rect 10493 5053 10507 5067
rect 10433 5013 10447 5027
rect 10473 5013 10487 5027
rect 10393 4893 10407 4907
rect 10393 4853 10407 4867
rect 10513 4853 10527 4867
rect 10453 4810 10467 4824
rect 10493 4810 10507 4824
rect 10373 4793 10387 4807
rect 10513 4753 10527 4767
rect 10433 4733 10447 4747
rect 10313 4693 10327 4707
rect 10353 4693 10367 4707
rect 10273 4613 10287 4627
rect 10353 4556 10367 4570
rect 10393 4556 10407 4570
rect 10293 4510 10307 4524
rect 10333 4453 10347 4467
rect 10333 4393 10347 4407
rect 10413 4493 10427 4507
rect 10393 4373 10407 4387
rect 10373 4336 10387 4350
rect 10413 4336 10427 4350
rect 10273 4290 10287 4304
rect 10353 4253 10367 4267
rect 10353 4193 10367 4207
rect 10313 4053 10327 4067
rect 10213 3893 10227 3907
rect 10213 3693 10227 3707
rect 10173 3553 10187 3567
rect 10173 3516 10187 3530
rect 10173 3473 10187 3487
rect 10153 3453 10167 3467
rect 10213 3413 10227 3427
rect 10153 3296 10167 3310
rect 10133 3053 10147 3067
rect 10133 3032 10147 3046
rect 10273 3990 10287 4004
rect 10353 3990 10367 4004
rect 10353 3853 10367 3867
rect 10313 3833 10327 3847
rect 10253 3816 10267 3830
rect 10293 3770 10307 3784
rect 10293 3713 10307 3727
rect 10253 3516 10267 3530
rect 10413 4233 10427 4247
rect 10333 3573 10347 3587
rect 10373 3573 10387 3587
rect 10413 3873 10427 3887
rect 10413 3816 10427 3830
rect 10413 3593 10427 3607
rect 10413 3572 10427 3586
rect 10313 3516 10327 3530
rect 10253 3293 10267 3307
rect 10333 3470 10347 3484
rect 10393 3433 10407 3447
rect 10333 3296 10347 3310
rect 10373 3296 10387 3310
rect 10273 3250 10287 3264
rect 10233 2993 10247 3007
rect 10173 2913 10187 2927
rect 10213 2913 10227 2927
rect 10093 2733 10107 2747
rect 10173 2733 10187 2747
rect 10133 2476 10147 2490
rect 10113 2430 10127 2444
rect 10173 2433 10187 2447
rect 10173 2393 10187 2407
rect 10293 3173 10307 3187
rect 10273 3133 10287 3147
rect 10253 2553 10267 2567
rect 10213 2473 10227 2487
rect 10233 2430 10247 2444
rect 10213 2373 10227 2387
rect 10153 2353 10167 2367
rect 10193 2353 10207 2367
rect 10213 2333 10227 2347
rect 10193 2256 10207 2270
rect 10073 1956 10087 1970
rect 10113 1956 10127 1970
rect 9993 1913 10007 1927
rect 10093 1910 10107 1924
rect 10053 1853 10067 1867
rect 10033 1736 10047 1750
rect 9993 1713 10007 1727
rect 10253 2393 10267 2407
rect 10393 3213 10407 3227
rect 10513 4633 10527 4647
rect 10473 4613 10487 4627
rect 10473 4213 10487 4227
rect 10633 5513 10647 5527
rect 10633 5273 10647 5287
rect 10633 5030 10647 5044
rect 10593 4893 10607 4907
rect 10553 4856 10567 4870
rect 10553 4593 10567 4607
rect 10593 4810 10607 4824
rect 10633 4653 10647 4667
rect 10593 4573 10607 4587
rect 10753 6853 10767 6867
rect 10733 6433 10747 6447
rect 10773 6553 10787 6567
rect 11013 7473 11027 7487
rect 10953 7456 10967 7470
rect 10993 7456 11007 7470
rect 11353 11570 11367 11584
rect 11293 11413 11307 11427
rect 11353 11353 11367 11367
rect 11453 11353 11467 11367
rect 11393 11316 11407 11330
rect 11433 11316 11447 11330
rect 11433 11173 11447 11187
rect 11373 11133 11387 11147
rect 11273 11050 11287 11064
rect 11233 11013 11247 11027
rect 11233 10913 11247 10927
rect 11213 10692 11227 10706
rect 11253 10853 11267 10867
rect 11233 10673 11247 10687
rect 11293 11013 11307 11027
rect 11273 10750 11287 10764
rect 11253 10653 11267 10667
rect 11173 10576 11187 10590
rect 11213 10576 11227 10590
rect 11273 10576 11287 10590
rect 11153 10530 11167 10544
rect 11253 10530 11267 10544
rect 11073 10473 11087 10487
rect 11053 9273 11067 9287
rect 11093 10413 11107 10427
rect 11093 10273 11107 10287
rect 11093 9710 11107 9724
rect 11073 9233 11087 9247
rect 11053 9173 11067 9187
rect 11133 10053 11147 10067
rect 11173 10353 11187 10367
rect 11213 10433 11227 10447
rect 11193 10273 11207 10287
rect 11193 10230 11207 10244
rect 11233 10230 11247 10244
rect 11173 10133 11187 10147
rect 11133 9773 11147 9787
rect 11313 10973 11327 10987
rect 11373 10833 11387 10847
rect 11453 11096 11467 11110
rect 11453 11053 11467 11067
rect 11433 10773 11447 10787
rect 11353 10750 11367 10764
rect 11313 10733 11327 10747
rect 11313 10633 11327 10647
rect 11293 10513 11307 10527
rect 11313 10313 11327 10327
rect 11273 10213 11287 10227
rect 11273 10073 11287 10087
rect 11313 10073 11327 10087
rect 11253 10056 11267 10070
rect 11273 9973 11287 9987
rect 11193 9933 11207 9947
rect 11233 9873 11247 9887
rect 11193 9833 11207 9847
rect 11273 9753 11287 9767
rect 11153 9653 11167 9667
rect 11233 9536 11247 9550
rect 11133 9293 11147 9307
rect 11173 9293 11187 9307
rect 11113 9233 11127 9247
rect 11213 9253 11227 9267
rect 11153 9190 11167 9204
rect 11213 9113 11227 9127
rect 11213 9013 11227 9027
rect 11193 8970 11207 8984
rect 11093 8953 11107 8967
rect 11153 8953 11167 8967
rect 11253 9193 11267 9207
rect 11293 9413 11307 9427
rect 11273 9173 11287 9187
rect 11253 9053 11267 9067
rect 11253 9016 11267 9030
rect 11353 10576 11367 10590
rect 11413 10576 11427 10590
rect 11373 10533 11387 10547
rect 11353 10473 11367 10487
rect 11433 10530 11447 10544
rect 11413 10493 11427 10507
rect 11373 10413 11387 10427
rect 11593 11616 11607 11630
rect 11613 11570 11627 11584
rect 11493 11333 11507 11347
rect 11573 11333 11587 11347
rect 11713 11733 11727 11747
rect 11693 11573 11707 11587
rect 11593 11270 11607 11284
rect 11633 11270 11647 11284
rect 11673 11270 11687 11284
rect 11573 11233 11587 11247
rect 11633 11233 11647 11247
rect 11533 11096 11547 11110
rect 11533 10813 11547 10827
rect 11493 10573 11507 10587
rect 11473 10393 11487 10407
rect 11393 10373 11407 10387
rect 11453 10276 11467 10290
rect 11513 10273 11527 10287
rect 11393 10230 11407 10244
rect 11433 10230 11447 10244
rect 11513 10133 11527 10147
rect 11393 10093 11407 10107
rect 11533 10093 11547 10107
rect 11353 10013 11367 10027
rect 11353 9793 11367 9807
rect 11413 10053 11427 10067
rect 11593 11050 11607 11064
rect 11673 11173 11687 11187
rect 11572 10893 11586 10907
rect 11593 10893 11607 10907
rect 11633 10893 11647 10907
rect 11553 10053 11567 10067
rect 11533 9973 11547 9987
rect 11493 9913 11507 9927
rect 11413 9873 11427 9887
rect 11393 9693 11407 9707
rect 11333 9536 11347 9550
rect 11453 9756 11467 9770
rect 11493 9693 11507 9707
rect 11533 9573 11547 9587
rect 11493 9536 11507 9550
rect 11333 9490 11347 9504
rect 11413 9490 11427 9504
rect 11513 9490 11527 9504
rect 11473 9433 11487 9447
rect 11453 9393 11467 9407
rect 11373 9353 11387 9367
rect 11413 9353 11427 9367
rect 11333 9253 11347 9267
rect 11293 8970 11307 8984
rect 11253 8853 11267 8867
rect 11233 8793 11247 8807
rect 11153 8716 11167 8730
rect 11233 8716 11247 8730
rect 11133 8553 11147 8567
rect 11073 8493 11087 8507
rect 11213 8653 11227 8667
rect 11253 8633 11267 8647
rect 11313 8713 11327 8727
rect 11353 8716 11367 8730
rect 11293 8593 11307 8607
rect 11153 8533 11167 8547
rect 11173 8496 11187 8510
rect 11273 8493 11287 8507
rect 11053 8213 11067 8227
rect 11053 7613 11067 7627
rect 11093 8253 11107 8267
rect 11153 8450 11167 8464
rect 11153 8433 11167 8447
rect 11273 8413 11287 8427
rect 11333 8693 11347 8707
rect 11313 8450 11327 8464
rect 11153 8213 11167 8227
rect 11153 8196 11167 8210
rect 11193 8213 11207 8227
rect 11273 8213 11287 8227
rect 11293 8213 11307 8227
rect 11273 8173 11287 8187
rect 11113 8153 11127 8167
rect 11173 8150 11187 8164
rect 11093 8113 11107 8127
rect 11273 8053 11287 8067
rect 11193 7973 11207 7987
rect 11233 7976 11247 7990
rect 11513 9236 11527 9250
rect 11473 9153 11487 9167
rect 11513 9153 11527 9167
rect 11473 9033 11487 9047
rect 11433 9016 11447 9030
rect 11413 8970 11427 8984
rect 11553 8853 11567 8867
rect 11493 8716 11507 8730
rect 11533 8716 11547 8730
rect 11633 10833 11647 10847
rect 11653 10733 11667 10747
rect 11593 10693 11607 10707
rect 11613 10573 11627 10587
rect 11673 10576 11687 10590
rect 11733 11593 11747 11607
rect 11733 11513 11747 11527
rect 11893 11893 11907 11907
rect 11773 11836 11787 11850
rect 11853 11836 11867 11850
rect 11873 11790 11887 11804
rect 11913 11790 11927 11804
rect 11973 11793 11987 11807
rect 11893 11753 11907 11767
rect 11773 11733 11787 11747
rect 11813 11633 11827 11647
rect 11853 11633 11867 11647
rect 11913 11570 11927 11584
rect 11973 11570 11987 11584
rect 12013 11573 12027 11587
rect 11873 11533 11887 11547
rect 11813 11433 11827 11447
rect 11953 11433 11967 11447
rect 11773 11313 11787 11327
rect 11913 11316 11927 11330
rect 11753 11273 11767 11287
rect 11893 11233 11907 11247
rect 11773 11092 11787 11106
rect 11813 11096 11827 11110
rect 11773 11053 11787 11067
rect 11833 11050 11847 11064
rect 11833 11013 11847 11027
rect 11893 11013 11907 11027
rect 11953 11013 11967 11027
rect 11793 10796 11807 10810
rect 11773 10773 11787 10787
rect 11733 10733 11747 10747
rect 11693 10530 11707 10544
rect 11733 10530 11747 10544
rect 11613 10493 11627 10507
rect 11613 10093 11627 10107
rect 11593 9973 11607 9987
rect 11613 9913 11627 9927
rect 11593 9573 11607 9587
rect 11593 8773 11607 8787
rect 11573 8733 11587 8747
rect 11373 8670 11387 8684
rect 11373 8633 11387 8647
rect 11453 8513 11467 8527
rect 11353 8496 11367 8510
rect 11413 8496 11427 8510
rect 11513 8670 11527 8684
rect 11333 8393 11347 8407
rect 11473 8493 11487 8507
rect 11393 8450 11407 8464
rect 11433 8450 11447 8464
rect 11353 8253 11367 8267
rect 11413 8253 11427 8267
rect 11373 8233 11387 8247
rect 11253 7930 11267 7944
rect 11293 7930 11307 7944
rect 11333 7930 11347 7944
rect 11193 7873 11207 7887
rect 11173 7773 11187 7787
rect 11193 7753 11207 7767
rect 11133 7676 11147 7690
rect 11153 7630 11167 7644
rect 11193 7630 11207 7644
rect 11113 7573 11127 7587
rect 11073 7553 11087 7567
rect 11073 7473 11087 7487
rect 10953 7253 10967 7267
rect 10893 7153 10907 7167
rect 11013 7410 11027 7424
rect 10973 7173 10987 7187
rect 10893 7113 10907 7127
rect 10873 6993 10887 7007
rect 10853 6853 10867 6867
rect 10953 6993 10967 7007
rect 10913 6693 10927 6707
rect 10933 6673 10947 6687
rect 10893 6635 10907 6649
rect 11313 7853 11327 7867
rect 11233 7673 11247 7687
rect 11293 7593 11307 7607
rect 11233 7472 11247 7486
rect 11133 7453 11147 7467
rect 11213 7453 11227 7467
rect 11093 7410 11107 7424
rect 11073 6993 11087 7007
rect 10973 6936 10987 6950
rect 11013 6936 11027 6950
rect 11053 6936 11067 6950
rect 10953 6633 10967 6647
rect 10873 6590 10887 6604
rect 10913 6553 10927 6567
rect 10833 6453 10847 6467
rect 10813 6433 10827 6447
rect 10753 6370 10767 6384
rect 10793 6370 10807 6384
rect 10793 6333 10807 6347
rect 10793 6293 10807 6307
rect 10733 6153 10747 6167
rect 10733 6113 10747 6127
rect 10873 6370 10887 6384
rect 10853 6133 10867 6147
rect 10833 6113 10847 6127
rect 10793 6033 10807 6047
rect 10773 5633 10787 5647
rect 10733 5593 10747 5607
rect 10953 6070 10967 6084
rect 10933 5993 10947 6007
rect 10813 5896 10827 5910
rect 10873 5896 10887 5910
rect 10913 5896 10927 5910
rect 10813 5853 10827 5867
rect 10813 5596 10827 5610
rect 10753 5550 10767 5564
rect 10793 5550 10807 5564
rect 10713 5513 10727 5527
rect 10893 5813 10907 5827
rect 10873 5573 10887 5587
rect 10853 5433 10867 5447
rect 10833 5413 10847 5427
rect 10773 5376 10787 5390
rect 10812 5373 10826 5387
rect 10833 5376 10847 5390
rect 10933 5433 10947 5447
rect 10753 5293 10767 5307
rect 10813 5293 10827 5307
rect 10933 5293 10947 5307
rect 10713 5073 10727 5087
rect 10713 5030 10727 5044
rect 10753 4933 10767 4947
rect 10733 4913 10747 4927
rect 10733 4873 10747 4887
rect 10713 4856 10727 4870
rect 10753 4856 10767 4870
rect 10673 4773 10687 4787
rect 10713 4733 10727 4747
rect 10693 4573 10707 4587
rect 10653 4510 10667 4524
rect 10613 4493 10627 4507
rect 10693 4492 10707 4506
rect 10613 4373 10627 4387
rect 10653 4336 10667 4350
rect 10593 4290 10607 4304
rect 10633 4290 10647 4304
rect 10673 4290 10687 4304
rect 10653 4253 10667 4267
rect 10653 4093 10667 4107
rect 10513 4073 10527 4087
rect 10493 4036 10507 4050
rect 10473 3953 10487 3967
rect 10493 3913 10507 3927
rect 10553 4036 10567 4050
rect 10593 4036 10607 4050
rect 10573 3990 10587 4004
rect 10593 3953 10607 3967
rect 10533 3833 10547 3847
rect 10473 3733 10487 3747
rect 10513 3733 10527 3747
rect 10453 3470 10467 3484
rect 10333 3113 10347 3127
rect 10373 3113 10387 3127
rect 10633 3853 10647 3867
rect 10613 3753 10627 3767
rect 10653 3753 10667 3767
rect 10533 3673 10547 3687
rect 10573 3673 10587 3687
rect 10553 3653 10567 3667
rect 10613 3633 10627 3647
rect 10613 3593 10627 3607
rect 10452 3053 10466 3067
rect 10473 3053 10487 3067
rect 10453 3013 10467 3027
rect 10393 2953 10407 2967
rect 10433 2950 10447 2964
rect 10333 2893 10347 2907
rect 10613 3516 10627 3530
rect 10573 3470 10587 3484
rect 10573 3353 10587 3367
rect 10533 3313 10547 3327
rect 10633 3313 10647 3327
rect 10513 3250 10527 3264
rect 10493 2853 10507 2867
rect 10433 2793 10447 2807
rect 10493 2793 10507 2807
rect 10393 2776 10407 2790
rect 10453 2733 10467 2747
rect 10413 2633 10427 2647
rect 10373 2553 10387 2567
rect 10413 2513 10427 2527
rect 10373 2476 10387 2490
rect 10413 2476 10427 2490
rect 10353 2430 10367 2444
rect 10473 2476 10487 2490
rect 10473 2433 10487 2447
rect 10273 2373 10287 2387
rect 10253 2256 10267 2270
rect 10373 2256 10387 2270
rect 10433 2256 10447 2270
rect 10172 2153 10186 2167
rect 10193 2153 10207 2167
rect 10193 2113 10207 2127
rect 10133 1793 10147 1807
rect 10113 1773 10127 1787
rect 10053 1690 10067 1704
rect 10093 1693 10107 1707
rect 10113 1613 10127 1627
rect 10093 1533 10107 1547
rect 10133 1513 10147 1527
rect 10093 1390 10107 1404
rect 10133 1390 10147 1404
rect 10313 2113 10327 2127
rect 10413 2210 10427 2224
rect 10373 1956 10387 1970
rect 10293 1910 10307 1924
rect 10333 1893 10347 1907
rect 10293 1793 10307 1807
rect 10333 1736 10347 1750
rect 10593 3250 10607 3264
rect 10593 3233 10607 3247
rect 10693 4036 10707 4050
rect 10733 4653 10747 4667
rect 10733 4593 10747 4607
rect 10733 4433 10747 4447
rect 10773 4773 10787 4787
rect 10753 4393 10767 4407
rect 10753 4213 10767 4227
rect 10733 4033 10747 4047
rect 10713 3993 10727 4007
rect 10713 3613 10727 3627
rect 10693 3513 10707 3527
rect 10673 3373 10687 3387
rect 10593 3212 10607 3226
rect 10633 3213 10647 3227
rect 10553 3173 10567 3187
rect 10553 3093 10567 3107
rect 10533 3053 10547 3067
rect 10533 2733 10547 2747
rect 10513 2513 10527 2527
rect 10513 2373 10527 2387
rect 10493 2153 10507 2167
rect 10493 2013 10507 2027
rect 10253 1593 10267 1607
rect 10253 1553 10267 1567
rect 10233 1453 10247 1467
rect 10153 1373 10167 1387
rect 10213 1373 10227 1387
rect 10153 1233 10167 1247
rect 10133 1216 10147 1230
rect 10173 1216 10187 1230
rect 10253 1333 10267 1347
rect 10253 1216 10267 1230
rect 9973 1173 9987 1187
rect 10153 1170 10167 1184
rect 10233 1173 10247 1187
rect 10313 1690 10327 1704
rect 10373 1693 10387 1707
rect 10353 1613 10367 1627
rect 10333 1216 10347 1230
rect 10253 1133 10267 1147
rect 9953 1093 9967 1107
rect 10173 1053 10187 1067
rect 10253 1053 10267 1067
rect 10293 1053 10307 1067
rect 9973 953 9987 967
rect 9933 813 9947 827
rect 10033 813 10047 827
rect 10153 813 10167 827
rect 9833 773 9847 787
rect 9893 773 9907 787
rect 9973 773 9987 787
rect 9533 613 9547 627
rect 9473 533 9487 547
rect 9413 433 9427 447
rect 9293 396 9307 410
rect 9773 650 9787 664
rect 9773 473 9787 487
rect 9713 433 9727 447
rect 9573 393 9587 407
rect 9813 453 9827 467
rect 9773 396 9787 410
rect 9453 333 9467 347
rect 9533 333 9547 347
rect 9293 273 9307 287
rect 9293 193 9307 207
rect 9533 176 9547 190
rect 10213 773 10227 787
rect 10233 733 10247 747
rect 9933 633 9947 647
rect 9993 513 10007 527
rect 10193 613 10207 627
rect 10033 473 10047 487
rect 10013 453 10027 467
rect 9953 396 9967 410
rect 9993 396 10007 410
rect 9933 353 9947 367
rect 9733 313 9747 327
rect 9813 313 9827 327
rect 9893 313 9907 327
rect 9613 176 9627 190
rect 10093 393 10107 407
rect 10013 350 10027 364
rect 10073 313 10087 327
rect 10093 273 10107 287
rect 10113 213 10127 227
rect 10112 173 10126 187
rect 10133 173 10147 187
rect 8513 130 8527 144
rect 8733 130 8747 144
rect 8993 130 9007 144
rect 9073 130 9087 144
rect 9213 130 9227 144
rect 9253 130 9267 144
rect 9293 130 9307 144
rect 9553 130 9567 144
rect 9613 133 9627 147
rect 9793 130 9807 144
rect 9953 133 9967 147
rect 10053 130 10067 144
rect 10413 1436 10427 1450
rect 10393 1390 10407 1404
rect 10433 1373 10447 1387
rect 10473 1313 10487 1327
rect 10433 1273 10447 1287
rect 10393 1253 10407 1267
rect 10433 1252 10447 1266
rect 10393 1216 10407 1230
rect 10573 2853 10587 2867
rect 10553 2256 10567 2270
rect 10713 3470 10727 3484
rect 10693 3250 10707 3264
rect 10613 3173 10627 3187
rect 10673 3173 10687 3187
rect 10753 3933 10767 3947
rect 10833 5273 10847 5287
rect 11033 6890 11047 6904
rect 10993 6733 11007 6747
rect 11013 6633 11027 6647
rect 11033 6413 11047 6427
rect 11013 6370 11027 6384
rect 11013 6153 11027 6167
rect 10993 6133 11007 6147
rect 11013 6013 11027 6027
rect 11013 5933 11027 5947
rect 10993 5813 11007 5827
rect 10953 5113 10967 5127
rect 10873 5076 10887 5090
rect 10933 5076 10947 5090
rect 10913 4973 10927 4987
rect 10913 4853 10927 4867
rect 10913 4810 10927 4824
rect 10913 4753 10927 4767
rect 10813 4733 10827 4747
rect 10953 4873 10967 4887
rect 10953 4753 10967 4767
rect 10933 4733 10947 4747
rect 10913 4613 10927 4627
rect 10813 4556 10827 4570
rect 10873 4556 10887 4570
rect 10833 4473 10847 4487
rect 10953 4510 10967 4524
rect 10893 4473 10907 4487
rect 10853 4393 10867 4407
rect 10953 4373 10967 4387
rect 10853 4333 10867 4347
rect 10913 4336 10927 4350
rect 10953 4336 10967 4350
rect 10873 4290 10887 4304
rect 10953 4253 10967 4267
rect 10813 4153 10827 4167
rect 10953 4153 10967 4167
rect 10813 4113 10827 4127
rect 10833 4073 10847 4087
rect 10793 4033 10807 4047
rect 10873 4036 10887 4050
rect 10913 4033 10927 4047
rect 10773 3833 10787 3847
rect 10773 3673 10787 3687
rect 10753 3413 10767 3427
rect 10853 3913 10867 3927
rect 10853 3873 10867 3887
rect 10913 3853 10927 3867
rect 10893 3816 10907 3830
rect 10933 3813 10947 3827
rect 10873 3733 10887 3747
rect 10913 3733 10927 3747
rect 10873 3712 10887 3726
rect 10813 3513 10827 3527
rect 10913 3553 10927 3567
rect 10933 3516 10947 3530
rect 11053 6173 11067 6187
rect 11153 7156 11167 7170
rect 11193 7156 11207 7170
rect 11213 7110 11227 7124
rect 11333 7673 11347 7687
rect 11533 8493 11547 8507
rect 11433 8150 11447 8164
rect 11513 8053 11527 8067
rect 11533 8013 11547 8027
rect 11453 7973 11467 7987
rect 11493 7973 11507 7987
rect 11593 8196 11607 8210
rect 11393 7676 11407 7690
rect 11593 8013 11607 8027
rect 11573 7953 11587 7967
rect 11513 7930 11527 7944
rect 11513 7753 11527 7767
rect 11573 7713 11587 7727
rect 11313 7413 11327 7427
rect 11153 7073 11167 7087
rect 11253 7073 11267 7087
rect 11233 6953 11247 6967
rect 11133 6733 11147 6747
rect 11213 6733 11227 6747
rect 11153 6673 11167 6687
rect 11173 6590 11187 6604
rect 11113 6513 11127 6527
rect 11093 6413 11107 6427
rect 11153 6416 11167 6430
rect 11153 6333 11167 6347
rect 11133 6233 11147 6247
rect 11113 6116 11127 6130
rect 11153 6116 11167 6130
rect 11193 6092 11207 6106
rect 11133 6070 11147 6084
rect 11093 6033 11107 6047
rect 11013 5596 11027 5610
rect 11073 5596 11087 5610
rect 11113 5973 11127 5987
rect 11093 5550 11107 5564
rect 11053 5513 11067 5527
rect 11033 5393 11047 5407
rect 11033 5376 11047 5390
rect 11093 5373 11107 5387
rect 10993 5133 11007 5147
rect 10993 5076 11007 5090
rect 11053 5330 11067 5344
rect 11193 5933 11207 5947
rect 11193 5896 11207 5910
rect 11233 6412 11247 6426
rect 11193 5833 11207 5847
rect 11173 5793 11187 5807
rect 11153 5596 11167 5610
rect 11033 5273 11047 5287
rect 11073 5093 11087 5107
rect 11053 5013 11067 5027
rect 11033 4953 11047 4967
rect 11033 4893 11047 4907
rect 11073 4853 11087 4867
rect 11013 4810 11027 4824
rect 11153 5493 11167 5507
rect 11213 5733 11227 5747
rect 11193 5333 11207 5347
rect 11153 5273 11167 5287
rect 11133 5093 11147 5107
rect 11173 5076 11187 5090
rect 11213 5076 11227 5090
rect 11313 6993 11327 7007
rect 11333 6953 11347 6967
rect 11433 7630 11447 7644
rect 11473 7613 11487 7627
rect 11553 7673 11567 7687
rect 11493 7593 11507 7607
rect 11513 7513 11527 7527
rect 11413 7413 11427 7427
rect 11393 7153 11407 7167
rect 11293 6890 11307 6904
rect 11333 6853 11347 6867
rect 11293 6753 11307 6767
rect 11273 6673 11287 6687
rect 11293 6590 11307 6604
rect 11353 6590 11367 6604
rect 11393 6713 11407 6727
rect 11493 7410 11507 7424
rect 11473 7156 11487 7170
rect 11453 7110 11467 7124
rect 11493 7033 11507 7047
rect 11513 7013 11527 7027
rect 11473 6953 11487 6967
rect 11453 6933 11467 6947
rect 11453 6753 11467 6767
rect 11413 6673 11427 6687
rect 11413 6636 11427 6650
rect 11433 6590 11447 6604
rect 11433 6513 11447 6527
rect 11293 6113 11307 6127
rect 11273 6033 11287 6047
rect 11253 5833 11267 5847
rect 11293 5693 11307 5707
rect 11273 5673 11287 5687
rect 11373 6416 11387 6430
rect 11473 6453 11487 6467
rect 11413 6371 11427 6385
rect 11473 6353 11487 6367
rect 11573 7013 11587 7027
rect 11653 10513 11667 10527
rect 11693 10353 11707 10367
rect 11693 10276 11707 10290
rect 11653 10173 11667 10187
rect 11633 9793 11647 9807
rect 11713 10230 11727 10244
rect 11693 10213 11707 10227
rect 11673 10153 11687 10167
rect 11813 10733 11827 10747
rect 11793 10633 11807 10647
rect 11793 10576 11807 10590
rect 11773 10433 11787 10447
rect 11873 10796 11887 10810
rect 11913 10796 11927 10810
rect 11893 10733 11907 10747
rect 11933 10733 11947 10747
rect 11933 10576 11947 10590
rect 12033 11353 12047 11367
rect 12013 11313 12027 11327
rect 11993 11253 12007 11267
rect 11993 10693 12007 10707
rect 11953 10530 11967 10544
rect 12013 10530 12027 10544
rect 11953 10473 11967 10487
rect 11913 10433 11927 10447
rect 11953 10276 11967 10290
rect 12013 10273 12027 10287
rect 11833 10233 11847 10247
rect 11873 10230 11887 10244
rect 11813 10173 11827 10187
rect 11793 10073 11807 10087
rect 11853 10053 11867 10067
rect 11693 10010 11707 10024
rect 11733 10010 11747 10024
rect 11673 9933 11687 9947
rect 11813 9993 11827 10007
rect 11773 9893 11787 9907
rect 11733 9756 11747 9770
rect 11793 9756 11807 9770
rect 11713 9710 11727 9724
rect 11753 9653 11767 9667
rect 11753 9573 11767 9587
rect 11793 9373 11807 9387
rect 11653 9353 11667 9367
rect 11733 9353 11747 9367
rect 11673 9273 11687 9287
rect 11813 9273 11827 9287
rect 11733 9236 11747 9250
rect 11673 9190 11687 9204
rect 11633 9113 11647 9127
rect 11753 9190 11767 9204
rect 11673 9093 11687 9107
rect 11713 9093 11727 9107
rect 11653 9033 11667 9047
rect 11653 8970 11667 8984
rect 11633 8593 11647 8607
rect 11713 9053 11727 9067
rect 11833 9213 11847 9227
rect 11753 9016 11767 9030
rect 11813 9016 11827 9030
rect 11733 8970 11747 8984
rect 11773 8970 11787 8984
rect 11753 8813 11767 8827
rect 11793 8733 11807 8747
rect 11673 8553 11687 8567
rect 11653 8513 11667 8527
rect 11713 8496 11727 8510
rect 11693 8433 11707 8447
rect 11813 8670 11827 8684
rect 11813 8553 11827 8567
rect 11793 8493 11807 8507
rect 11733 8433 11747 8447
rect 11773 8433 11787 8447
rect 11653 8353 11667 8367
rect 11653 8193 11667 8207
rect 11713 8196 11727 8210
rect 11673 8153 11687 8167
rect 11673 8093 11687 8107
rect 11793 8013 11807 8027
rect 11673 7976 11687 7990
rect 11733 7976 11747 7990
rect 11773 7976 11787 7990
rect 11833 8496 11847 8510
rect 11833 8113 11847 8127
rect 11673 7933 11687 7947
rect 11653 7893 11667 7907
rect 11753 7893 11767 7907
rect 11693 7693 11707 7707
rect 11673 7676 11687 7690
rect 11793 7773 11807 7787
rect 11793 7693 11807 7707
rect 11653 7630 11667 7644
rect 11693 7630 11707 7644
rect 11773 7630 11787 7644
rect 11613 7613 11627 7627
rect 11653 7613 11667 7627
rect 11753 7593 11767 7607
rect 11833 7673 11847 7687
rect 11813 7573 11827 7587
rect 11793 7513 11807 7527
rect 11753 7393 11767 7407
rect 11633 7373 11647 7387
rect 11613 7153 11627 7167
rect 11553 6953 11567 6967
rect 11593 6953 11607 6967
rect 11573 6936 11587 6950
rect 11673 7333 11687 7347
rect 11633 7110 11647 7124
rect 11633 6953 11647 6967
rect 11613 6933 11627 6947
rect 11553 6890 11567 6904
rect 11533 6853 11547 6867
rect 11593 6793 11607 6807
rect 11713 7253 11727 7267
rect 11753 7156 11767 7170
rect 11773 7110 11787 7124
rect 11753 6973 11767 6987
rect 11733 6873 11747 6887
rect 11673 6853 11687 6867
rect 11593 6633 11607 6647
rect 11533 6370 11547 6384
rect 11353 6173 11367 6187
rect 11473 6153 11487 6167
rect 11353 6116 11367 6130
rect 11453 6073 11467 6087
rect 11393 6033 11407 6047
rect 11413 5933 11427 5947
rect 11473 6033 11487 6047
rect 11333 5733 11347 5747
rect 11313 5633 11327 5647
rect 11313 5596 11327 5610
rect 11293 5550 11307 5564
rect 11333 5550 11347 5564
rect 11313 5533 11327 5547
rect 11293 5393 11307 5407
rect 11313 5373 11327 5387
rect 11253 5333 11267 5347
rect 11133 5013 11147 5027
rect 11113 4853 11127 4867
rect 11033 4733 11047 4747
rect 11013 4453 11027 4467
rect 10993 3753 11007 3767
rect 10973 3633 10987 3647
rect 10793 3393 10807 3407
rect 10773 3353 10787 3367
rect 10753 3213 10767 3227
rect 10913 3470 10927 3484
rect 10993 3553 11007 3567
rect 10853 3433 10867 3447
rect 10973 3433 10987 3447
rect 10833 3250 10847 3264
rect 10773 3193 10787 3207
rect 10793 3113 10807 3127
rect 10753 3013 10767 3027
rect 10673 2996 10687 3010
rect 10733 2992 10747 3006
rect 10613 2950 10627 2964
rect 10653 2950 10667 2964
rect 10693 2913 10707 2927
rect 10693 2873 10707 2887
rect 10733 2853 10747 2867
rect 10713 2813 10727 2827
rect 10673 2776 10687 2790
rect 10593 2733 10607 2747
rect 10653 2593 10667 2607
rect 10653 2513 10667 2527
rect 10733 2776 10747 2790
rect 10733 2733 10747 2747
rect 10693 2493 10707 2507
rect 10693 2476 10707 2490
rect 10673 2430 10687 2444
rect 10633 2393 10647 2407
rect 10613 2353 10627 2367
rect 10593 2293 10607 2307
rect 10573 2233 10587 2247
rect 10533 2193 10547 2207
rect 10533 2033 10547 2047
rect 10533 1973 10547 1987
rect 10553 1956 10567 1970
rect 10633 2313 10647 2327
rect 10733 2273 10747 2287
rect 10673 2256 10687 2270
rect 10613 2193 10627 2207
rect 10633 2113 10647 2127
rect 10713 2210 10727 2224
rect 10673 2193 10687 2207
rect 10653 1953 10667 1967
rect 10573 1910 10587 1924
rect 10613 1910 10627 1924
rect 10593 1893 10607 1907
rect 10513 1833 10527 1847
rect 10573 1833 10587 1847
rect 10613 1773 10627 1787
rect 10593 1690 10607 1704
rect 10553 1653 10567 1667
rect 10553 1533 10567 1547
rect 10593 1533 10607 1547
rect 10353 1113 10367 1127
rect 10413 1170 10427 1184
rect 10493 1173 10507 1187
rect 10373 973 10387 987
rect 10473 973 10487 987
rect 10353 953 10367 967
rect 10353 873 10367 887
rect 10333 813 10347 827
rect 10253 650 10267 664
rect 10233 553 10247 567
rect 10213 473 10227 487
rect 10313 650 10327 664
rect 10273 513 10287 527
rect 10393 916 10407 930
rect 10433 916 10447 930
rect 10453 870 10467 884
rect 10493 853 10507 867
rect 10393 653 10407 667
rect 10693 1993 10707 2007
rect 10693 1693 10707 1707
rect 10653 1390 10667 1404
rect 10573 1373 10587 1387
rect 10653 1353 10667 1367
rect 10573 1253 10587 1267
rect 10693 1253 10707 1267
rect 10653 1216 10667 1230
rect 10673 1170 10687 1184
rect 10693 1113 10707 1127
rect 10753 1736 10767 1750
rect 10733 1073 10747 1087
rect 10573 873 10587 887
rect 10673 870 10687 884
rect 10713 833 10727 847
rect 10613 793 10627 807
rect 10613 673 10627 687
rect 10793 2996 10807 3010
rect 10873 3193 10887 3207
rect 10833 3173 10847 3187
rect 10813 2813 10827 2827
rect 10813 2593 10827 2607
rect 10813 2513 10827 2527
rect 10793 2476 10807 2490
rect 10993 3113 11007 3127
rect 10993 3053 11007 3067
rect 10953 2996 10967 3010
rect 11053 4413 11067 4427
rect 11053 3990 11067 4004
rect 11033 3773 11047 3787
rect 10933 2893 10947 2907
rect 10893 2776 10907 2790
rect 10973 2813 10987 2827
rect 10993 2776 11007 2790
rect 10873 2693 10887 2707
rect 10973 2730 10987 2744
rect 10913 2653 10927 2667
rect 10853 2613 10867 2627
rect 10833 2393 10847 2407
rect 10833 2293 10847 2307
rect 10833 2210 10847 2224
rect 10813 2133 10827 2147
rect 10953 2573 10967 2587
rect 10993 2533 11007 2547
rect 10993 2476 11007 2490
rect 10893 2430 10907 2444
rect 10933 2430 10947 2444
rect 10913 2333 10927 2347
rect 10873 2273 10887 2287
rect 10853 2093 10867 2107
rect 10793 2073 10807 2087
rect 10813 2013 10827 2027
rect 10973 2393 10987 2407
rect 10953 2293 10967 2307
rect 10933 2210 10947 2224
rect 10873 1993 10887 2007
rect 10813 1955 10827 1969
rect 10933 1973 10947 1987
rect 10893 1955 10907 1969
rect 10833 1910 10847 1924
rect 10853 1892 10867 1906
rect 10913 1893 10927 1907
rect 10793 1853 10807 1867
rect 10793 1773 10807 1787
rect 10933 1753 10947 1767
rect 10893 1736 10907 1750
rect 10793 1693 10807 1707
rect 10833 1690 10847 1704
rect 10873 1673 10887 1687
rect 10933 1573 10947 1587
rect 10793 1513 10807 1527
rect 10993 2373 11007 2387
rect 10993 2073 11007 2087
rect 10993 1873 11007 1887
rect 10993 1673 11007 1687
rect 10973 1513 10987 1527
rect 10793 1373 10807 1387
rect 10853 1353 10867 1367
rect 10793 953 10807 967
rect 10953 1373 10967 1387
rect 10913 1353 10927 1367
rect 10873 1253 10887 1267
rect 10953 1253 10967 1267
rect 10913 1216 10927 1230
rect 10933 1170 10947 1184
rect 10993 1153 11007 1167
rect 10873 1133 10887 1147
rect 10953 1073 10967 1087
rect 10913 953 10927 967
rect 10853 873 10867 887
rect 10813 753 10827 767
rect 10773 693 10787 707
rect 10973 870 10987 884
rect 10933 713 10947 727
rect 10893 693 10907 707
rect 10493 650 10507 664
rect 10373 453 10387 467
rect 10573 650 10587 664
rect 10753 653 10767 667
rect 10533 613 10547 627
rect 10753 396 10767 410
rect 10793 393 10807 407
rect 10213 350 10227 364
rect 10273 350 10287 364
rect 10373 350 10387 364
rect 10513 350 10527 364
rect 10293 313 10307 327
rect 10333 233 10347 247
rect 10293 176 10307 190
rect 10773 350 10787 364
rect 10813 350 10827 364
rect 10873 573 10887 587
rect 10733 313 10747 327
rect 10833 313 10847 327
rect 10453 156 10467 170
rect 10493 156 10507 170
rect 10193 133 10207 147
rect 10313 130 10327 144
rect 9033 113 9047 127
rect 9293 113 9307 127
rect 8773 93 8787 107
rect 10653 150 10667 164
rect 10773 156 10787 170
rect 10853 153 10867 167
rect 10813 110 10827 124
rect 10993 676 11007 690
rect 10933 633 10947 647
rect 11033 2256 11047 2270
rect 11033 2213 11047 2227
rect 11033 1953 11047 1967
rect 10893 193 10907 207
rect 11013 552 11027 566
rect 11013 396 11027 410
rect 11093 4653 11107 4667
rect 11093 4493 11107 4507
rect 11193 5030 11207 5044
rect 11233 5033 11247 5047
rect 11313 5333 11327 5347
rect 11273 5293 11287 5307
rect 11333 5313 11347 5327
rect 11313 5273 11327 5287
rect 11293 5213 11307 5227
rect 11273 5053 11287 5067
rect 11153 4993 11167 5007
rect 11153 4953 11167 4967
rect 11213 4933 11227 4947
rect 11173 4693 11187 4707
rect 11133 4673 11147 4687
rect 11213 4556 11227 4570
rect 11253 4993 11267 5007
rect 11132 4513 11146 4527
rect 11153 4510 11167 4524
rect 11113 4433 11127 4447
rect 11193 4493 11207 4507
rect 11193 4373 11207 4387
rect 11133 4290 11147 4304
rect 11153 4273 11167 4287
rect 11233 4273 11247 4287
rect 11213 4233 11227 4247
rect 11173 4213 11187 4227
rect 11213 4036 11227 4050
rect 11193 3990 11207 4004
rect 11133 3933 11147 3947
rect 11213 3933 11227 3947
rect 11212 3873 11226 3887
rect 11233 3873 11247 3887
rect 11133 3853 11147 3867
rect 11093 3773 11107 3787
rect 11193 3673 11207 3687
rect 11113 3553 11127 3567
rect 11153 3553 11167 3567
rect 11113 3513 11127 3527
rect 11153 3516 11167 3530
rect 11213 3513 11227 3527
rect 11133 3470 11147 3484
rect 11133 3433 11147 3447
rect 11093 3373 11107 3387
rect 11173 3373 11187 3387
rect 11173 3296 11187 3310
rect 11193 3233 11207 3247
rect 11153 3213 11167 3227
rect 11093 3133 11107 3147
rect 11133 3093 11147 3107
rect 11113 3033 11127 3047
rect 11073 2293 11087 2307
rect 11053 1673 11067 1687
rect 11153 2996 11167 3010
rect 11133 2913 11147 2927
rect 11193 3212 11207 3226
rect 11193 3173 11207 3187
rect 11353 5073 11367 5087
rect 11333 5053 11347 5067
rect 11313 4853 11327 4867
rect 11433 5850 11447 5864
rect 11473 5793 11487 5807
rect 11493 5673 11507 5687
rect 11413 5633 11427 5647
rect 11393 5493 11407 5507
rect 11453 5173 11467 5187
rect 11413 5073 11427 5087
rect 11593 6590 11607 6604
rect 11653 6590 11667 6604
rect 11593 6493 11607 6507
rect 11693 6493 11707 6507
rect 11973 10230 11987 10244
rect 11933 10153 11947 10167
rect 11973 9893 11987 9907
rect 11893 9833 11907 9847
rect 12093 11893 12107 11907
rect 12153 11853 12167 11867
rect 12093 11790 12107 11804
rect 12133 11790 12147 11804
rect 12173 11753 12187 11767
rect 12253 11693 12267 11707
rect 12173 11616 12187 11630
rect 12313 11616 12327 11630
rect 12213 11570 12227 11584
rect 12253 11570 12267 11584
rect 12153 11353 12167 11367
rect 12153 11316 12167 11330
rect 12133 11253 12147 11267
rect 12073 11233 12087 11247
rect 12093 11096 12107 11110
rect 12073 11050 12087 11064
rect 12053 10796 12067 10810
rect 12053 10733 12067 10747
rect 12113 11013 12127 11027
rect 12093 10973 12107 10987
rect 12173 10973 12187 10987
rect 12173 10796 12187 10810
rect 12213 10796 12227 10810
rect 12093 10733 12107 10747
rect 12153 10733 12167 10747
rect 12073 10653 12087 10667
rect 12073 10313 12087 10327
rect 12213 10713 12227 10727
rect 12193 10673 12207 10687
rect 12153 10633 12167 10647
rect 12133 10276 12147 10290
rect 12133 10233 12147 10247
rect 12133 10173 12147 10187
rect 12093 10133 12107 10147
rect 12053 10093 12067 10107
rect 12033 10053 12047 10067
rect 12073 9993 12087 10007
rect 12073 9893 12087 9907
rect 11873 9713 11887 9727
rect 11873 9013 11887 9027
rect 11873 7713 11887 7727
rect 11913 9793 11927 9807
rect 11993 9793 12007 9807
rect 11953 9756 11967 9770
rect 11973 9710 11987 9724
rect 12053 9753 12067 9767
rect 11953 9533 11967 9547
rect 12013 9536 12027 9550
rect 12073 9713 12087 9727
rect 12113 9533 12127 9547
rect 11953 9490 11967 9504
rect 11993 9490 12007 9504
rect 12073 9490 12087 9504
rect 12033 9273 12047 9287
rect 11993 9236 12007 9250
rect 12033 9236 12047 9250
rect 12093 9236 12107 9250
rect 12013 9190 12027 9204
rect 11973 9053 11987 9067
rect 12033 9053 12047 9067
rect 11933 8970 11947 8984
rect 11993 8970 12007 8984
rect 12033 8973 12047 8987
rect 11913 8693 11927 8707
rect 12013 8853 12027 8867
rect 12053 8716 12067 8730
rect 11933 8673 11947 8687
rect 12033 8670 12047 8684
rect 11933 8593 11947 8607
rect 11993 8496 12007 8510
rect 12073 8495 12087 8509
rect 11953 8450 11967 8464
rect 12013 8450 12027 8464
rect 12053 8450 12067 8464
rect 11953 8196 11967 8210
rect 12073 8413 12087 8427
rect 12073 8193 12087 8207
rect 12073 8150 12087 8164
rect 11933 8113 11947 8127
rect 12013 8013 12027 8027
rect 12053 7976 12067 7990
rect 11913 7713 11927 7727
rect 11973 7676 11987 7690
rect 11853 6973 11867 6987
rect 11933 7613 11947 7627
rect 12073 7753 12087 7767
rect 11953 7533 11967 7547
rect 12033 7533 12047 7547
rect 11933 7473 11947 7487
rect 11933 7093 11947 7107
rect 11613 6453 11627 6467
rect 11753 6453 11767 6467
rect 11593 6393 11607 6407
rect 11553 6070 11567 6084
rect 11533 5850 11547 5864
rect 11653 6413 11667 6427
rect 11733 6416 11747 6430
rect 11793 6935 11807 6949
rect 11833 6935 11847 6949
rect 11873 6935 11887 6949
rect 11633 6153 11647 6167
rect 11713 6370 11727 6384
rect 11773 6373 11787 6387
rect 11753 6353 11767 6367
rect 11753 6233 11767 6247
rect 11673 6116 11687 6130
rect 11653 6070 11667 6084
rect 11613 6033 11627 6047
rect 11653 5993 11667 6007
rect 11693 5993 11707 6007
rect 11633 5933 11647 5947
rect 11693 5953 11707 5967
rect 11653 5893 11667 5907
rect 11773 6033 11787 6047
rect 11773 5953 11787 5967
rect 11753 5913 11767 5927
rect 11733 5896 11747 5910
rect 11633 5793 11647 5807
rect 11613 5773 11627 5787
rect 11753 5853 11767 5867
rect 11693 5833 11707 5847
rect 11673 5693 11687 5707
rect 11593 5673 11607 5687
rect 11513 5633 11527 5647
rect 11633 5633 11647 5647
rect 11673 5633 11687 5647
rect 11513 5593 11527 5607
rect 11573 5596 11587 5610
rect 11493 5075 11507 5089
rect 11613 5550 11627 5564
rect 11613 5513 11627 5527
rect 11533 5377 11547 5391
rect 11573 5377 11587 5391
rect 11713 5773 11727 5787
rect 11673 5473 11687 5487
rect 11733 5693 11747 5707
rect 11673 5331 11687 5345
rect 11713 5333 11727 5347
rect 11613 5313 11627 5327
rect 11393 5013 11407 5027
rect 11433 5013 11447 5027
rect 11393 4893 11407 4907
rect 11373 4853 11387 4867
rect 11293 4811 11307 4825
rect 11513 5033 11527 5047
rect 11473 4973 11487 4987
rect 11353 4793 11367 4807
rect 11433 4793 11447 4807
rect 11333 4753 11347 4767
rect 11333 4573 11347 4587
rect 11273 4513 11287 4527
rect 11313 4433 11327 4447
rect 11293 4373 11307 4387
rect 11273 4333 11287 4347
rect 11273 4290 11287 4304
rect 11293 4233 11307 4247
rect 11293 4212 11307 4226
rect 11273 4113 11287 4127
rect 11273 4036 11287 4050
rect 11253 3433 11267 3447
rect 11313 3873 11327 3887
rect 11373 4673 11387 4687
rect 11433 4613 11447 4627
rect 11513 4813 11527 4827
rect 11513 4792 11527 4806
rect 11493 4773 11507 4787
rect 11453 4573 11467 4587
rect 11473 4556 11487 4570
rect 11493 4513 11507 4527
rect 11453 4493 11467 4507
rect 11513 4453 11527 4467
rect 11473 4393 11487 4407
rect 11413 4373 11427 4387
rect 11433 4336 11447 4350
rect 11413 4233 11427 4247
rect 11433 4233 11447 4247
rect 11393 4133 11407 4147
rect 11493 4293 11507 4307
rect 11453 4073 11467 4087
rect 11493 4193 11507 4207
rect 11513 4133 11527 4147
rect 11473 4036 11487 4050
rect 11393 3993 11407 4007
rect 11453 3990 11467 4004
rect 11393 3953 11407 3967
rect 11373 3933 11387 3947
rect 11473 3933 11487 3947
rect 11433 3816 11447 3830
rect 11333 3713 11347 3727
rect 11333 3493 11347 3507
rect 11413 3753 11427 3767
rect 11413 3553 11427 3567
rect 11453 3516 11467 3530
rect 11373 3473 11387 3487
rect 11433 3470 11447 3484
rect 11313 3273 11327 3287
rect 11293 3250 11307 3264
rect 11253 3233 11267 3247
rect 11233 3033 11247 3047
rect 11273 3133 11287 3147
rect 11213 2996 11227 3010
rect 11253 2996 11267 3010
rect 11173 2953 11187 2967
rect 11273 2953 11287 2967
rect 11233 2913 11247 2927
rect 11153 2853 11167 2867
rect 11233 2853 11247 2867
rect 11133 2773 11147 2787
rect 11193 2776 11207 2790
rect 11173 2730 11187 2744
rect 11213 2693 11227 2707
rect 11133 2573 11147 2587
rect 11213 2573 11227 2587
rect 11133 2533 11147 2547
rect 11173 2473 11187 2487
rect 11293 2793 11307 2807
rect 11313 2593 11327 2607
rect 11273 2553 11287 2567
rect 11313 2553 11327 2567
rect 11273 2476 11287 2490
rect 11133 2373 11147 2387
rect 11233 2413 11247 2427
rect 11153 2256 11167 2270
rect 11253 2353 11267 2367
rect 11233 2193 11247 2207
rect 11213 2153 11227 2167
rect 11173 2133 11187 2147
rect 11153 2013 11167 2027
rect 11113 1953 11127 1967
rect 11093 1793 11107 1807
rect 11133 1753 11147 1767
rect 11173 1733 11187 1747
rect 11113 1690 11127 1704
rect 11233 1953 11247 1967
rect 11213 1673 11227 1687
rect 11173 1653 11187 1667
rect 11133 1413 11147 1427
rect 11073 1353 11087 1367
rect 11073 1216 11087 1230
rect 11213 1313 11227 1327
rect 11173 1293 11187 1307
rect 11173 1233 11187 1247
rect 11173 1216 11187 1230
rect 11133 1173 11147 1187
rect 11193 1170 11207 1184
rect 11213 1133 11227 1147
rect 11213 1093 11227 1107
rect 11153 913 11167 927
rect 11273 2253 11287 2267
rect 11373 3253 11387 3267
rect 11353 3113 11367 3127
rect 11393 3193 11407 3207
rect 11513 3753 11527 3767
rect 11513 3593 11527 3607
rect 11493 3433 11507 3447
rect 11493 3393 11507 3407
rect 11513 3253 11527 3267
rect 11473 3213 11487 3227
rect 11393 3053 11407 3067
rect 11433 3053 11447 3067
rect 11373 2913 11387 2927
rect 11353 2613 11367 2627
rect 11353 2533 11367 2547
rect 11333 2253 11347 2267
rect 11333 2232 11347 2246
rect 11313 2113 11327 2127
rect 11293 2093 11307 2107
rect 11293 1910 11307 1924
rect 11273 1793 11287 1807
rect 11253 913 11267 927
rect 11073 753 11087 767
rect 11113 713 11127 727
rect 11093 650 11107 664
rect 10993 350 11007 364
rect 11033 313 11047 327
rect 10993 233 11007 247
rect 11133 393 11147 407
rect 11093 293 11107 307
rect 11173 813 11187 827
rect 11233 833 11247 847
rect 11253 773 11267 787
rect 11193 713 11207 727
rect 11233 713 11247 727
rect 11253 650 11267 664
rect 11233 433 11247 447
rect 11193 413 11207 427
rect 11173 313 11187 327
rect 11153 176 11167 190
rect 11273 473 11287 487
rect 11373 2273 11387 2287
rect 11373 2210 11387 2224
rect 11413 2996 11427 3010
rect 11513 2996 11527 3010
rect 11693 5153 11707 5167
rect 11633 5133 11647 5147
rect 11593 5076 11607 5090
rect 11553 5033 11567 5047
rect 11573 4973 11587 4987
rect 11553 4853 11567 4867
rect 11553 4432 11567 4446
rect 11593 4933 11607 4947
rect 11633 4933 11647 4947
rect 11773 5713 11787 5727
rect 11773 5593 11787 5607
rect 11753 5393 11767 5407
rect 11733 5113 11747 5127
rect 11693 5076 11707 5090
rect 11733 5076 11747 5090
rect 11653 4855 11667 4869
rect 11633 4810 11647 4824
rect 11653 4673 11667 4687
rect 11633 4510 11647 4524
rect 11573 4273 11587 4287
rect 11553 4153 11567 4167
rect 11553 4073 11567 4087
rect 11613 4413 11627 4427
rect 11753 5030 11767 5044
rect 11753 4953 11767 4967
rect 11733 4556 11747 4570
rect 11713 4510 11727 4524
rect 11673 4453 11687 4467
rect 11653 4413 11667 4427
rect 11773 4453 11787 4467
rect 11753 4393 11767 4407
rect 11673 4336 11687 4350
rect 11693 4293 11707 4307
rect 11653 4193 11667 4207
rect 11613 3933 11627 3947
rect 11733 4273 11747 4287
rect 11713 4233 11727 4247
rect 11693 4033 11707 4047
rect 11753 4193 11767 4207
rect 11773 4073 11787 4087
rect 11673 4013 11687 4027
rect 11553 3013 11567 3027
rect 11453 2950 11467 2964
rect 11473 2913 11487 2927
rect 11493 2893 11507 2907
rect 11533 2793 11547 2807
rect 11493 2693 11507 2707
rect 11493 2513 11507 2527
rect 11453 2476 11467 2490
rect 11453 2413 11467 2427
rect 11493 2333 11507 2347
rect 11493 2293 11507 2307
rect 11453 2256 11467 2270
rect 11653 3873 11667 3887
rect 11593 3853 11607 3867
rect 11633 3816 11647 3830
rect 11773 3990 11787 4004
rect 11713 3953 11727 3967
rect 11733 3913 11747 3927
rect 11593 3773 11607 3787
rect 11633 3733 11647 3747
rect 11613 3713 11627 3727
rect 11593 3516 11607 3530
rect 11693 3770 11707 3784
rect 11753 3873 11767 3887
rect 11733 3733 11747 3747
rect 11652 3713 11666 3727
rect 11673 3713 11687 3727
rect 11753 3713 11767 3727
rect 11633 3473 11647 3487
rect 11613 3452 11627 3466
rect 11713 3633 11727 3647
rect 11833 6873 11847 6887
rect 11813 6793 11827 6807
rect 11793 3633 11807 3647
rect 11853 6653 11867 6667
rect 11873 6633 11887 6647
rect 12033 7473 12047 7487
rect 11993 7393 12007 7407
rect 12033 7373 12047 7387
rect 11993 7313 12007 7327
rect 11973 7153 11987 7167
rect 12053 7333 12067 7347
rect 12113 8716 12127 8730
rect 12113 8670 12127 8684
rect 12293 11093 12307 11107
rect 12273 10796 12287 10810
rect 12273 10713 12287 10727
rect 12253 10633 12267 10647
rect 12233 10530 12247 10544
rect 12193 10473 12207 10487
rect 12213 10313 12227 10327
rect 12253 10276 12267 10290
rect 12193 10213 12207 10227
rect 12233 9833 12247 9847
rect 12233 9756 12247 9770
rect 12153 9233 12167 9247
rect 12173 9013 12187 9027
rect 12153 8973 12167 8987
rect 12133 8613 12147 8627
rect 12133 7633 12147 7647
rect 12113 7553 12127 7567
rect 12113 7373 12127 7387
rect 12093 7313 12107 7327
rect 12113 7253 12127 7267
rect 12073 7156 12087 7170
rect 12033 7093 12047 7107
rect 11993 6936 12007 6950
rect 11973 6793 11987 6807
rect 11953 6733 11967 6747
rect 11913 6653 11927 6667
rect 11933 6573 11947 6587
rect 11873 6553 11887 6567
rect 11913 6553 11927 6567
rect 11913 6453 11927 6467
rect 11873 6373 11887 6387
rect 11873 6313 11887 6327
rect 11893 6273 11907 6287
rect 11973 6593 11987 6607
rect 11953 6453 11967 6467
rect 12053 7072 12067 7086
rect 12093 7073 12107 7087
rect 11993 6573 12007 6587
rect 12033 6573 12047 6587
rect 12113 6936 12127 6950
rect 12093 6873 12107 6887
rect 12073 6812 12087 6826
rect 12053 6433 12067 6447
rect 12033 6416 12047 6430
rect 11973 6353 11987 6367
rect 11933 6253 11947 6267
rect 11973 6193 11987 6207
rect 11913 6173 11927 6187
rect 11913 6133 11927 6147
rect 11893 6053 11907 6067
rect 11873 5853 11887 5867
rect 12033 6173 12047 6187
rect 12013 6053 12027 6067
rect 11933 6033 11947 6047
rect 11973 6033 11987 6047
rect 11933 5993 11947 6007
rect 11913 5873 11927 5887
rect 11873 5653 11887 5667
rect 11853 5593 11867 5607
rect 11913 5793 11927 5807
rect 11893 5633 11907 5647
rect 12053 6033 12067 6047
rect 12033 5993 12047 6007
rect 12013 5913 12027 5927
rect 12033 5833 12047 5847
rect 11993 5753 12007 5767
rect 12033 5653 12047 5667
rect 11913 5593 11927 5607
rect 11953 5593 11967 5607
rect 12013 5573 12027 5587
rect 11833 4993 11847 5007
rect 11913 5549 11927 5563
rect 11973 5513 11987 5527
rect 11933 5473 11947 5487
rect 11973 5473 11987 5487
rect 11873 5433 11887 5447
rect 11933 5413 11947 5427
rect 12013 5473 12027 5487
rect 12013 5413 12027 5427
rect 11993 5393 12007 5407
rect 11873 5330 11887 5344
rect 11913 5330 11927 5344
rect 11953 5330 11967 5344
rect 11913 5153 11927 5167
rect 11873 5076 11887 5090
rect 12053 5330 12067 5344
rect 12253 9710 12267 9724
rect 12213 9653 12227 9667
rect 12313 10173 12327 10187
rect 12293 9490 12307 9504
rect 12253 9236 12267 9250
rect 12233 9190 12247 9204
rect 12273 9053 12287 9067
rect 12233 9016 12247 9030
rect 12293 8970 12307 8984
rect 12213 8713 12227 8727
rect 12293 8716 12307 8730
rect 12273 8670 12287 8684
rect 12333 8613 12347 8627
rect 12233 8513 12247 8527
rect 12213 8495 12227 8509
rect 12233 8450 12247 8464
rect 12313 8353 12327 8367
rect 12213 8233 12227 8247
rect 12173 8193 12187 8207
rect 12293 8193 12307 8207
rect 12233 8150 12247 8164
rect 12193 8093 12207 8107
rect 12233 7753 12247 7767
rect 12213 7713 12227 7727
rect 12253 7676 12267 7690
rect 12173 7633 12187 7647
rect 12193 7573 12207 7587
rect 12193 7552 12207 7566
rect 12193 6873 12207 6887
rect 12173 6813 12187 6827
rect 12273 7633 12287 7647
rect 12233 6713 12247 6727
rect 12233 6673 12247 6687
rect 12093 6473 12107 6487
rect 12093 6433 12107 6447
rect 12093 6313 12107 6327
rect 12093 6273 12107 6287
rect 12073 5193 12087 5207
rect 11932 5113 11946 5127
rect 11953 5113 11967 5127
rect 12033 5113 12047 5127
rect 11913 5030 11927 5044
rect 11873 4953 11887 4967
rect 11893 4856 11907 4870
rect 11933 4856 11947 4870
rect 11873 4793 11887 4807
rect 11833 4553 11847 4567
rect 11933 4753 11947 4767
rect 11913 4593 11927 4607
rect 11893 4573 11907 4587
rect 11873 4336 11887 4350
rect 11873 4253 11887 4267
rect 11873 4033 11887 4047
rect 11873 3893 11887 3907
rect 12053 5076 12067 5090
rect 12033 5030 12047 5044
rect 12053 4993 12067 5007
rect 12033 4953 12047 4967
rect 11993 4933 12007 4947
rect 12013 4853 12027 4867
rect 11973 4673 11987 4687
rect 11953 4573 11967 4587
rect 11933 4553 11947 4567
rect 12113 6133 12127 6147
rect 12113 6073 12127 6087
rect 12113 5313 12127 5327
rect 12113 5073 12127 5087
rect 12053 4813 12067 4827
rect 12033 4773 12047 4787
rect 12033 4653 12047 4667
rect 12053 4613 12067 4627
rect 12033 4553 12047 4567
rect 11993 4510 12007 4524
rect 11993 4433 12007 4447
rect 11953 4393 11967 4407
rect 11953 4336 11967 4350
rect 11973 4290 11987 4304
rect 12053 4290 12067 4304
rect 11933 4253 11947 4267
rect 11913 4013 11927 4027
rect 11953 4213 11967 4227
rect 12053 4213 12067 4227
rect 11993 4036 12007 4050
rect 11913 3973 11927 3987
rect 11893 3853 11907 3867
rect 11873 3816 11887 3830
rect 11913 3816 11927 3830
rect 12013 3990 12027 4004
rect 11973 3973 11987 3987
rect 12013 3853 12027 3867
rect 11833 3633 11847 3647
rect 11813 3593 11827 3607
rect 11753 3553 11767 3567
rect 11793 3553 11807 3567
rect 11693 3473 11707 3487
rect 11673 3333 11687 3347
rect 11733 3353 11747 3367
rect 11773 3353 11787 3367
rect 11713 3313 11727 3327
rect 11773 3332 11787 3346
rect 11593 3093 11607 3107
rect 11673 3250 11687 3264
rect 11713 3153 11727 3167
rect 11673 3113 11687 3127
rect 11633 3013 11647 3027
rect 11633 2992 11647 3006
rect 11573 2912 11587 2926
rect 11573 2853 11587 2867
rect 11473 2210 11487 2224
rect 11513 2213 11527 2227
rect 11413 2173 11427 2187
rect 11353 2153 11367 2167
rect 11393 2153 11407 2167
rect 11353 1993 11367 2007
rect 11333 1793 11347 1807
rect 11473 2153 11487 2167
rect 11393 1910 11407 1924
rect 11413 1853 11427 1867
rect 11353 1736 11367 1750
rect 11373 1673 11387 1687
rect 11333 1593 11347 1607
rect 11313 1513 11327 1527
rect 11333 1436 11347 1450
rect 11453 1793 11467 1807
rect 11453 1633 11467 1647
rect 11473 1593 11487 1607
rect 11373 1413 11387 1427
rect 11373 1293 11387 1307
rect 11333 1213 11347 1227
rect 11373 1170 11387 1184
rect 11433 1436 11447 1450
rect 11513 1493 11527 1507
rect 11493 1433 11507 1447
rect 11473 1373 11487 1387
rect 11433 1353 11447 1367
rect 11433 1273 11447 1287
rect 11473 1233 11487 1247
rect 11473 1216 11487 1230
rect 11453 1170 11467 1184
rect 11393 1113 11407 1127
rect 11313 1013 11327 1027
rect 11393 916 11407 930
rect 11453 916 11467 930
rect 11333 793 11347 807
rect 11333 753 11347 767
rect 11313 733 11327 747
rect 11473 870 11487 884
rect 11473 813 11487 827
rect 11393 713 11407 727
rect 11413 676 11427 690
rect 11613 2353 11627 2367
rect 11713 3073 11727 3087
rect 11753 3213 11767 3227
rect 11733 2950 11747 2964
rect 11693 2853 11707 2867
rect 11693 2793 11707 2807
rect 11773 2853 11787 2867
rect 11673 2733 11687 2747
rect 11713 2653 11727 2667
rect 11673 2633 11687 2647
rect 11653 2513 11667 2527
rect 11613 2253 11627 2267
rect 11593 2213 11607 2227
rect 11633 2232 11647 2246
rect 11813 2893 11827 2907
rect 11793 2776 11807 2790
rect 11793 2593 11807 2607
rect 11713 2553 11727 2567
rect 11773 2553 11787 2567
rect 11673 2393 11687 2407
rect 11753 2476 11767 2490
rect 11793 2476 11807 2490
rect 11773 2430 11787 2444
rect 11773 2393 11787 2407
rect 11733 2293 11747 2307
rect 11713 2273 11727 2287
rect 11693 2256 11707 2270
rect 11813 2273 11827 2287
rect 11613 2173 11627 2187
rect 11733 2113 11747 2127
rect 11673 1956 11687 1970
rect 11573 1913 11587 1927
rect 11553 993 11567 1007
rect 11653 1910 11667 1924
rect 11633 1793 11647 1807
rect 11673 1736 11687 1750
rect 11713 1910 11727 1924
rect 11693 1733 11707 1747
rect 11753 2073 11767 2087
rect 11753 1993 11767 2007
rect 11753 1893 11767 1907
rect 11733 1853 11747 1867
rect 11753 1793 11767 1807
rect 11733 1736 11747 1750
rect 11653 1673 11667 1687
rect 11713 1673 11727 1687
rect 11633 1593 11647 1607
rect 11593 1553 11607 1567
rect 11593 1473 11607 1487
rect 11613 1436 11627 1450
rect 11593 1353 11607 1367
rect 11633 1390 11647 1404
rect 11753 1690 11767 1704
rect 11733 1473 11747 1487
rect 11693 1436 11707 1450
rect 11733 1436 11747 1450
rect 11793 1433 11807 1447
rect 11713 1390 11727 1404
rect 11713 1353 11727 1367
rect 11653 1273 11667 1287
rect 11753 1213 11767 1227
rect 11653 1170 11667 1184
rect 11693 1170 11707 1184
rect 11613 1133 11627 1147
rect 11793 1133 11807 1147
rect 11633 1113 11647 1127
rect 11573 973 11587 987
rect 11813 1033 11827 1047
rect 11813 973 11827 987
rect 11673 916 11687 930
rect 11713 916 11727 930
rect 11673 853 11687 867
rect 11813 853 11827 867
rect 11793 833 11807 847
rect 11633 813 11647 827
rect 11733 813 11747 827
rect 11553 773 11567 787
rect 11793 753 11807 767
rect 11913 3753 11927 3767
rect 11893 3593 11907 3607
rect 11873 3553 11887 3567
rect 11873 3473 11887 3487
rect 11853 3172 11867 3186
rect 11853 713 11867 727
rect 11953 3713 11967 3727
rect 11933 3673 11947 3687
rect 11933 3573 11947 3587
rect 11973 3633 11987 3647
rect 12053 3753 12067 3767
rect 12053 3633 12067 3647
rect 12013 3573 12027 3587
rect 11973 3553 11987 3567
rect 12013 3516 12027 3530
rect 12053 3513 12067 3527
rect 11953 3473 11967 3487
rect 11933 3432 11947 3446
rect 11913 3413 11927 3427
rect 11913 3293 11927 3307
rect 11893 3173 11907 3187
rect 11893 3152 11907 3166
rect 11893 2433 11907 2447
rect 11993 3470 12007 3484
rect 12053 3473 12067 3487
rect 12033 3433 12047 3447
rect 11973 3413 11987 3427
rect 11953 3293 11967 3307
rect 12013 3296 12027 3310
rect 12053 3253 12067 3267
rect 12033 3193 12047 3207
rect 11993 2996 12007 3010
rect 11933 2950 11947 2964
rect 11973 2950 11987 2964
rect 12013 2913 12027 2927
rect 11973 2833 11987 2847
rect 12013 2776 12027 2790
rect 11973 2633 11987 2647
rect 11953 2493 11967 2507
rect 11933 2473 11947 2487
rect 11913 2252 11927 2266
rect 11913 2173 11927 2187
rect 12053 2533 12067 2547
rect 12013 2513 12027 2527
rect 11993 2493 12007 2507
rect 12033 2476 12047 2490
rect 12153 6632 12167 6646
rect 12193 6636 12207 6650
rect 12333 7713 12347 7727
rect 12313 6713 12327 6727
rect 12293 6673 12307 6687
rect 12273 6633 12287 6647
rect 12153 6293 12167 6307
rect 12193 6573 12207 6587
rect 12213 6533 12227 6547
rect 12213 6473 12227 6487
rect 12273 6453 12287 6467
rect 12333 6413 12347 6427
rect 12233 6353 12247 6367
rect 12333 6373 12347 6387
rect 12313 6253 12327 6267
rect 12213 6070 12227 6084
rect 12173 6032 12187 6046
rect 12253 5953 12267 5967
rect 12193 5896 12207 5910
rect 12233 5896 12247 5910
rect 12253 5833 12267 5847
rect 12193 5793 12207 5807
rect 12253 5753 12267 5767
rect 12193 5596 12207 5610
rect 12212 5553 12226 5567
rect 12233 5550 12247 5564
rect 12273 5550 12287 5564
rect 12213 5513 12227 5527
rect 12233 5376 12247 5390
rect 12293 5513 12307 5527
rect 12273 5373 12287 5387
rect 12153 5313 12167 5327
rect 12213 5333 12227 5347
rect 12173 5233 12187 5247
rect 12193 5076 12207 5090
rect 12153 4953 12167 4967
rect 12153 4856 12167 4870
rect 12273 5333 12287 5347
rect 12273 5273 12287 5287
rect 12273 5233 12287 5247
rect 12213 5033 12227 5047
rect 12113 4812 12127 4826
rect 12113 4313 12127 4327
rect 12093 4253 12107 4267
rect 12173 4810 12187 4824
rect 12173 4773 12187 4787
rect 12153 4673 12167 4687
rect 12133 4253 12147 4267
rect 12093 3713 12107 3727
rect 12093 3673 12107 3687
rect 12093 2833 12107 2847
rect 12093 2730 12107 2744
rect 11953 2430 11967 2444
rect 12013 2430 12027 2444
rect 11973 2293 11987 2307
rect 12033 2413 12047 2427
rect 12012 2255 12026 2269
rect 12053 2373 12067 2387
rect 12033 2253 12047 2267
rect 11993 2210 12007 2224
rect 11933 2153 11947 2167
rect 12033 1973 12047 1987
rect 11913 1956 11927 1970
rect 12013 1953 12027 1967
rect 11933 1893 11947 1907
rect 11913 1773 11927 1787
rect 11953 1753 11967 1767
rect 12013 1736 12027 1750
rect 11973 1690 11987 1704
rect 11913 1633 11927 1647
rect 11893 1453 11907 1467
rect 11933 1533 11947 1547
rect 12013 1533 12027 1547
rect 12053 1913 12067 1927
rect 12093 1833 12107 1847
rect 12073 1753 12087 1767
rect 12073 1690 12087 1704
rect 12033 1453 12047 1467
rect 11913 1273 11927 1287
rect 11933 1233 11947 1247
rect 12033 1390 12047 1404
rect 12033 1213 12047 1227
rect 11993 1170 12007 1184
rect 12093 1393 12107 1407
rect 11953 1133 11967 1147
rect 11933 993 11947 1007
rect 11893 712 11907 726
rect 11513 670 11527 684
rect 11673 670 11687 684
rect 11793 676 11807 690
rect 11373 650 11387 664
rect 11833 573 11847 587
rect 11333 553 11347 567
rect 11733 553 11747 567
rect 11413 433 11427 447
rect 11293 413 11307 427
rect 11313 333 11327 347
rect 11813 473 11827 487
rect 11573 376 11587 390
rect 11793 393 11807 407
rect 11693 370 11707 384
rect 11773 373 11787 387
rect 11413 333 11427 347
rect 11793 333 11807 347
rect 11293 313 11307 327
rect 11373 313 11387 327
rect 11033 130 11047 144
rect 11133 130 11147 144
rect 11193 130 11207 144
rect 10873 110 10887 124
rect 11613 273 11627 287
rect 11333 253 11347 267
rect 11373 176 11387 190
rect 11673 173 11687 187
rect 11913 353 11927 367
rect 11873 176 11887 190
rect 11973 1013 11987 1027
rect 12033 1170 12047 1184
rect 12073 953 12087 967
rect 12133 4033 12147 4047
rect 12133 1973 12147 1987
rect 12233 4813 12247 4827
rect 12213 4753 12227 4767
rect 12213 4713 12227 4727
rect 12193 4573 12207 4587
rect 12293 5193 12307 5207
rect 12273 4813 12287 4827
rect 12313 4713 12327 4727
rect 12293 4673 12307 4687
rect 12253 4573 12267 4587
rect 12313 4573 12327 4587
rect 12333 4553 12347 4567
rect 12233 4513 12247 4527
rect 12213 4493 12227 4507
rect 12273 4393 12287 4407
rect 12333 4513 12347 4527
rect 12313 4493 12327 4507
rect 12293 4333 12307 4347
rect 12193 4233 12207 4247
rect 12253 4290 12267 4304
rect 12293 4293 12307 4307
rect 12253 4233 12267 4247
rect 12293 4033 12307 4047
rect 12293 3993 12307 4007
rect 12273 3933 12287 3947
rect 12233 3913 12247 3927
rect 12253 3873 12267 3887
rect 12193 3813 12207 3827
rect 12253 3816 12267 3830
rect 12193 3733 12207 3747
rect 12233 3773 12247 3787
rect 12253 3753 12267 3767
rect 12233 3573 12247 3587
rect 12213 3553 12227 3567
rect 12213 3516 12227 3530
rect 12313 3753 12327 3767
rect 12333 3733 12347 3747
rect 12293 3653 12307 3667
rect 12273 3533 12287 3547
rect 12193 3393 12207 3407
rect 12253 3516 12267 3530
rect 12333 3553 12347 3567
rect 12333 3513 12347 3527
rect 12273 3470 12287 3484
rect 12313 3470 12327 3484
rect 12233 3433 12247 3447
rect 12213 3373 12227 3387
rect 12193 3333 12207 3347
rect 12293 3433 12307 3447
rect 12273 3373 12287 3387
rect 12253 3313 12267 3327
rect 12293 3333 12307 3347
rect 12333 3393 12347 3407
rect 12313 3293 12327 3307
rect 12213 3253 12227 3267
rect 12213 3213 12227 3227
rect 12193 3193 12207 3207
rect 12293 3250 12307 3264
rect 12313 3213 12327 3227
rect 12293 3193 12307 3207
rect 12253 3113 12267 3127
rect 12193 3033 12207 3047
rect 12253 3013 12267 3027
rect 12253 2730 12267 2744
rect 12173 2373 12187 2387
rect 12173 1993 12187 2007
rect 12233 2153 12247 2167
rect 12233 1956 12247 1970
rect 12033 870 12047 884
rect 12073 870 12087 884
rect 11993 853 12007 867
rect 12073 833 12087 847
rect 11993 693 12007 707
rect 11973 673 11987 687
rect 11953 633 11967 647
rect 11993 433 12007 447
rect 11973 396 11987 410
rect 12093 773 12107 787
rect 12073 713 12087 727
rect 12053 696 12067 710
rect 12073 650 12087 664
rect 12053 633 12067 647
rect 11993 350 12007 364
rect 11353 130 11367 144
rect 11393 113 11407 127
rect 11633 130 11647 144
rect 11673 130 11687 144
rect 11813 130 11827 144
rect 11853 130 11867 144
rect 11593 93 11607 107
rect 11813 93 11827 107
rect 11953 113 11967 127
rect 12153 1913 12167 1927
rect 12253 1913 12267 1927
rect 12213 1873 12227 1887
rect 12213 1736 12227 1750
rect 12293 1993 12307 2007
rect 12273 1833 12287 1847
rect 12193 1690 12207 1704
rect 12233 1493 12247 1507
rect 12253 1390 12267 1404
rect 12173 1373 12187 1387
rect 12233 1373 12247 1387
rect 12173 1273 12187 1287
rect 12213 1170 12227 1184
rect 12193 1033 12207 1047
rect 12173 433 12187 447
rect 12233 870 12247 884
rect 12253 433 12267 447
rect 12193 413 12207 427
rect 12173 353 12187 367
rect 12233 350 12247 364
rect 12153 293 12167 307
rect 12133 176 12147 190
rect 12173 176 12187 190
rect 12053 133 12067 147
rect 12153 130 12167 144
rect 12033 93 12047 107
rect 12213 93 12227 107
rect 12313 273 12327 287
rect 12333 253 12347 267
rect 8173 53 8187 67
rect 10493 53 10507 67
rect 11293 53 11307 67
rect 11893 53 11907 67
rect 12293 53 12307 67
rect 7513 13 7527 27
rect 7553 13 7567 27
rect 7693 13 7707 27
<< metal3 >>
rect 4107 12236 4173 12244
rect 2247 12216 2453 12224
rect 9067 12216 9833 12224
rect 2847 12196 3613 12204
rect 4587 12196 4673 12204
rect 9387 12196 10413 12204
rect 407 12176 493 12184
rect 2327 12176 2433 12184
rect 3156 12176 3833 12184
rect 247 12139 313 12147
rect 427 12136 453 12144
rect 716 12136 753 12144
rect 716 12107 724 12136
rect 847 12136 993 12144
rect 1067 12136 1253 12144
rect 1547 12139 1573 12147
rect 1707 12139 1753 12147
rect 1807 12136 2033 12144
rect 2087 12136 2113 12144
rect 2167 12136 2353 12144
rect 2787 12136 2953 12144
rect 2967 12136 2993 12144
rect 2447 12113 2573 12121
rect 2596 12116 2833 12124
rect 3156 12124 3164 12176
rect 4547 12176 4713 12184
rect 6047 12176 6213 12184
rect 8567 12176 9053 12184
rect 10467 12176 11393 12184
rect 11487 12176 11724 12184
rect 3767 12156 3873 12164
rect 3887 12156 6673 12164
rect 6687 12156 6753 12164
rect 6807 12156 6933 12164
rect 8367 12156 8453 12164
rect 9107 12156 9793 12164
rect 11716 12164 11724 12176
rect 11716 12156 11993 12164
rect 3567 12136 3633 12144
rect 3687 12136 4093 12144
rect 4387 12136 4553 12144
rect 4647 12136 4984 12144
rect 5787 12136 5892 12144
rect 227 12096 393 12104
rect 2596 12104 2604 12116
rect 787 12093 833 12101
rect 1247 12093 1353 12101
rect 2107 12093 2153 12101
rect 2387 12096 2604 12104
rect 2896 12087 2904 12116
rect 3287 12116 3353 12124
rect 4976 12124 4984 12136
rect 5927 12139 6073 12147
rect 6247 12136 6384 12144
rect 7767 12139 7953 12147
rect 7967 12136 7993 12144
rect 5107 12116 5173 12124
rect 6187 12119 6213 12127
rect 6376 12124 6384 12136
rect 8667 12139 8733 12147
rect 9256 12136 9353 12144
rect 3867 12093 3913 12101
rect 4407 12096 4532 12104
rect 4567 12093 4613 12101
rect 5907 12093 6013 12101
rect 6116 12087 6124 12116
rect 6507 12116 6713 12124
rect 6727 12116 6912 12124
rect 6947 12113 7033 12121
rect 7207 12119 7233 12127
rect 7307 12119 7333 12127
rect 7707 12096 7773 12104
rect 8056 12104 8064 12116
rect 8267 12113 8352 12121
rect 8387 12116 8453 12124
rect 9256 12124 9264 12136
rect 9907 12136 10113 12144
rect 10387 12136 10593 12144
rect 10607 12139 10653 12147
rect 10707 12139 10753 12147
rect 10927 12139 10953 12147
rect 11067 12139 11193 12147
rect 11387 12139 11433 12147
rect 11667 12139 11693 12147
rect 11747 12139 11773 12147
rect 12047 12139 12073 12147
rect 12247 12139 12333 12147
rect 9387 12116 9404 12124
rect 7787 12100 8084 12104
rect 7787 12096 8087 12100
rect 8073 12087 8087 12096
rect 8687 12093 9093 12101
rect 9396 12087 9404 12116
rect 747 12076 1053 12084
rect 1747 12076 1793 12084
rect 2896 12076 2913 12087
rect 2900 12073 2913 12076
rect 5767 12076 6053 12084
rect 6116 12076 6133 12087
rect 6120 12073 6133 12076
rect 6227 12076 7193 12084
rect 9403 12076 9404 12087
rect 9496 12116 9513 12124
rect 9496 12087 9504 12116
rect 9647 12113 9933 12121
rect 10407 12093 10453 12101
rect 10767 12096 11013 12104
rect 11107 12096 11713 12104
rect 9496 12076 9497 12087
rect 10147 12076 10633 12084
rect 11047 12076 11373 12084
rect 3927 12056 4573 12064
rect 6547 12056 6873 12064
rect 9447 12056 9473 12064
rect 10527 12056 10713 12064
rect 11407 12056 11453 12064
rect 1707 12036 1733 12044
rect 2427 12036 3673 12044
rect 5447 12036 5513 12044
rect 5527 12036 5833 12044
rect 6827 12036 6853 12044
rect 7947 12036 8633 12044
rect 9807 12036 10973 12044
rect 4367 12016 4653 12024
rect 4667 12016 4973 12024
rect 6067 12016 6693 12024
rect 9947 12016 10673 12024
rect 2927 11996 3193 12004
rect 3207 11996 3533 12004
rect 6227 11996 6333 12004
rect 6887 11996 6933 12004
rect 7527 11996 8413 12004
rect 8587 11996 8733 12004
rect 8747 11996 10013 12004
rect 5147 11976 5333 11984
rect 5807 11976 6133 11984
rect 6147 11976 6413 11984
rect 6687 11976 6953 11984
rect 4147 11956 4173 11964
rect 4187 11956 4773 11964
rect 7307 11956 7333 11964
rect 8947 11956 10353 11964
rect 687 11936 2193 11944
rect 2427 11936 2553 11944
rect 6247 11936 6533 11944
rect 527 11916 913 11924
rect 4987 11916 5273 11924
rect 5287 11916 5753 11924
rect 5927 11916 6484 11924
rect 3327 11896 4233 11904
rect 4247 11896 4713 11904
rect 6476 11904 6484 11916
rect 6507 11916 6793 11924
rect 6476 11896 6773 11904
rect 8827 11896 9493 11904
rect 10587 11896 11653 11904
rect 11667 11896 11893 11904
rect 11907 11896 12093 11904
rect 427 11876 793 11884
rect 1647 11876 1793 11884
rect 5387 11876 5653 11884
rect 6387 11876 7533 11884
rect 7747 11876 8193 11884
rect 8707 11876 8973 11884
rect 9447 11876 9973 11884
rect 10076 11876 10733 11884
rect 1207 11856 1413 11864
rect 4727 11859 4753 11867
rect 4767 11856 5133 11864
rect 5847 11856 5933 11864
rect 8247 11856 8413 11864
rect 8536 11856 8724 11864
rect 8536 11850 8544 11856
rect 467 11839 493 11847
rect 587 11839 753 11847
rect 927 11839 1053 11847
rect 1107 11839 1173 11847
rect 1687 11839 1753 11847
rect 1927 11839 2133 11847
rect 536 11824 544 11836
rect 2347 11836 2373 11844
rect 2387 11839 2473 11847
rect 3247 11836 3433 11844
rect 3447 11839 3473 11847
rect 3527 11836 3713 11844
rect 3727 11836 3824 11844
rect 5027 11839 5053 11847
rect 5187 11839 5233 11847
rect 5287 11840 5364 11844
rect 5287 11836 5367 11840
rect 536 11816 593 11824
rect 2516 11824 2524 11836
rect 2516 11816 2573 11824
rect 2627 11819 2713 11827
rect 3816 11824 3824 11836
rect 596 11804 604 11813
rect 2907 11813 2973 11821
rect 3867 11816 3913 11824
rect 4567 11819 4653 11827
rect 5353 11827 5367 11836
rect 6287 11836 6453 11844
rect 6547 11839 6633 11847
rect 6727 11839 6753 11847
rect 6967 11839 7053 11847
rect 7107 11836 7293 11844
rect 7647 11839 7673 11847
rect 347 11796 604 11804
rect 727 11793 773 11801
rect 1027 11796 1073 11804
rect 1527 11793 1693 11801
rect 1707 11796 1893 11804
rect 1947 11796 2053 11804
rect 2187 11793 2373 11801
rect 2447 11796 2493 11804
rect 196 11764 204 11789
rect 527 11776 573 11784
rect 1287 11776 1653 11784
rect 2536 11776 2613 11784
rect 196 11756 253 11764
rect 267 11756 313 11764
rect 327 11756 453 11764
rect 1127 11756 1193 11764
rect 1347 11756 1393 11764
rect 2536 11764 2544 11776
rect 2227 11756 2544 11764
rect 3447 11756 3893 11764
rect 407 11736 793 11744
rect 2927 11736 3013 11744
rect 3027 11736 3113 11744
rect 2427 11716 2533 11724
rect 2587 11716 2893 11724
rect 3587 11716 3793 11724
rect 3807 11716 4033 11724
rect 1327 11696 1573 11704
rect 2007 11696 2293 11704
rect 4076 11704 4084 11816
rect 4907 11793 4953 11801
rect 5496 11804 5504 11816
rect 5667 11813 5693 11821
rect 5907 11819 6073 11827
rect 7336 11824 7344 11836
rect 7807 11836 7853 11844
rect 7927 11836 8133 11844
rect 8207 11836 8473 11844
rect 8487 11839 8533 11847
rect 8716 11844 8724 11856
rect 10076 11864 10084 11876
rect 10867 11876 11884 11884
rect 9507 11856 10084 11864
rect 10247 11856 10533 11864
rect 11227 11856 11353 11864
rect 11876 11864 11884 11876
rect 11876 11856 12153 11864
rect 8716 11836 8733 11844
rect 8947 11836 9013 11844
rect 9167 11839 9193 11847
rect 9247 11839 9293 11847
rect 10027 11836 10213 11844
rect 10707 11839 10813 11847
rect 11127 11839 11313 11847
rect 11427 11836 11633 11844
rect 11787 11839 11853 11847
rect 7267 11816 7344 11824
rect 8567 11813 9613 11821
rect 9827 11819 10173 11827
rect 5167 11796 5504 11804
rect 5947 11796 6213 11804
rect 6227 11796 6373 11804
rect 6427 11796 6513 11804
rect 6787 11796 6844 11804
rect 4667 11776 4933 11784
rect 5207 11776 5373 11784
rect 5707 11776 5873 11784
rect 6547 11776 6713 11784
rect 6836 11784 6844 11796
rect 6867 11796 7073 11804
rect 7887 11793 7913 11801
rect 7936 11796 9253 11804
rect 6836 11776 7313 11784
rect 7727 11776 7833 11784
rect 7936 11784 7944 11796
rect 9487 11796 9553 11804
rect 10387 11793 10533 11801
rect 10807 11793 10853 11801
rect 11347 11796 11393 11804
rect 11707 11793 11873 11801
rect 11927 11796 11973 11804
rect 12107 11793 12133 11801
rect 7847 11776 7944 11784
rect 8767 11776 8813 11784
rect 8967 11776 9293 11784
rect 10227 11776 10253 11784
rect 10267 11776 11193 11784
rect 11207 11776 11593 11784
rect 4287 11756 5173 11764
rect 5687 11756 6813 11764
rect 7067 11756 7253 11764
rect 7347 11756 8113 11764
rect 10367 11756 11073 11764
rect 11907 11756 12173 11764
rect 4867 11736 5153 11744
rect 5176 11736 6713 11744
rect 5176 11724 5184 11736
rect 7167 11736 7613 11744
rect 7627 11736 8233 11744
rect 10967 11736 11713 11744
rect 11727 11736 11773 11744
rect 4787 11716 5184 11724
rect 5827 11716 6273 11724
rect 6827 11716 7873 11724
rect 8007 11716 8173 11724
rect 8187 11716 8453 11724
rect 8467 11716 8613 11724
rect 10307 11716 10493 11724
rect 4007 11696 4084 11704
rect 4327 11696 4373 11704
rect 4507 11696 5753 11704
rect 7107 11696 7613 11704
rect 7627 11696 7673 11704
rect 8407 11696 9233 11704
rect 9287 11696 9413 11704
rect 9427 11696 10593 11704
rect 10607 11696 10753 11704
rect 10767 11696 11413 11704
rect 11487 11696 12253 11704
rect 247 11676 673 11684
rect 787 11676 873 11684
rect 887 11676 2333 11684
rect 5367 11676 5493 11684
rect 6787 11676 7013 11684
rect 7027 11676 8713 11684
rect 2427 11656 2793 11664
rect 3087 11656 3113 11664
rect 3127 11656 3833 11664
rect 3847 11656 3873 11664
rect 3887 11656 4353 11664
rect 4367 11656 4713 11664
rect 4727 11656 4793 11664
rect 4807 11656 5293 11664
rect 5307 11656 5653 11664
rect 7307 11656 7573 11664
rect 287 11636 333 11644
rect 827 11636 853 11644
rect 1127 11636 1153 11644
rect 1867 11636 2044 11644
rect 2036 11630 2044 11636
rect 2387 11636 2493 11644
rect 2567 11636 2824 11644
rect 296 11616 493 11624
rect 707 11619 753 11627
rect 296 11604 304 11616
rect 907 11616 1073 11624
rect 1207 11619 1353 11627
rect 1907 11619 1933 11627
rect 2047 11619 2093 11627
rect 2627 11616 2693 11624
rect 2816 11624 2824 11636
rect 3747 11636 3773 11644
rect 6387 11636 6473 11644
rect 6487 11636 6924 11644
rect 2816 11616 3413 11624
rect 3467 11619 3492 11627
rect 3527 11616 3713 11624
rect 4427 11619 4533 11627
rect 4587 11616 4733 11624
rect 4807 11619 4893 11627
rect 5407 11619 5573 11627
rect 5627 11616 5833 11624
rect 5947 11619 6013 11627
rect 6916 11624 6924 11636
rect 9527 11636 10013 11644
rect 10067 11636 10253 11644
rect 10267 11636 10393 11644
rect 11827 11636 11853 11644
rect 6916 11616 7293 11624
rect 7587 11619 7653 11627
rect 7847 11619 7913 11627
rect 236 11596 304 11604
rect 236 11584 244 11596
rect 2487 11596 2593 11604
rect 2607 11596 2792 11604
rect 2827 11593 2913 11601
rect 3187 11599 3233 11607
rect 4356 11596 4404 11604
rect 227 11576 244 11584
rect 347 11573 513 11581
rect 607 11576 813 11584
rect 927 11573 1053 11581
rect 1167 11576 1333 11584
rect 4356 11584 4364 11596
rect 1767 11576 1873 11584
rect 2347 11573 2393 11581
rect 3787 11573 3973 11581
rect 4027 11573 4113 11581
rect 4347 11576 4364 11584
rect 4396 11584 4404 11596
rect 4787 11596 4973 11604
rect 7376 11604 7384 11616
rect 8087 11616 8553 11624
rect 8727 11619 8893 11627
rect 9767 11616 10353 11624
rect 10527 11619 10613 11627
rect 10867 11619 10953 11627
rect 11067 11619 11233 11627
rect 11307 11619 11333 11627
rect 11607 11616 11644 11624
rect 12187 11619 12313 11627
rect 5107 11593 5253 11601
rect 7376 11596 7473 11604
rect 11636 11604 11644 11616
rect 8267 11593 8393 11601
rect 11636 11596 11733 11604
rect 4396 11576 4493 11584
rect 4507 11576 4593 11584
rect 5487 11573 5593 11581
rect 5647 11573 5813 11581
rect 6567 11576 6793 11584
rect 7127 11573 7153 11581
rect 8627 11573 8653 11581
rect 9267 11576 9493 11584
rect 10047 11576 10273 11584
rect 10327 11573 10353 11581
rect 10407 11576 10593 11584
rect 11367 11576 11613 11584
rect 11627 11576 11693 11584
rect 11927 11573 11973 11581
rect 11987 11576 12013 11584
rect 12227 11573 12253 11581
rect 2547 11553 2753 11561
rect 3527 11556 4293 11564
rect 6047 11556 6213 11564
rect 6227 11556 6293 11564
rect 7647 11556 7893 11564
rect 8607 11556 8693 11564
rect 8767 11556 9213 11564
rect 9667 11556 10553 11564
rect 1807 11536 2093 11544
rect 2107 11536 2153 11544
rect 3707 11536 4033 11544
rect 4267 11536 4573 11544
rect 6167 11536 6333 11544
rect 6347 11536 6493 11544
rect 7027 11536 7073 11544
rect 7487 11536 7833 11544
rect 8427 11536 8733 11544
rect 9747 11536 9813 11544
rect 10007 11536 10693 11544
rect 11047 11536 11873 11544
rect 227 11516 253 11524
rect 2527 11516 2713 11524
rect 4127 11516 4793 11524
rect 6536 11516 6973 11524
rect 987 11496 1093 11504
rect 1107 11496 1873 11504
rect 1947 11496 2113 11504
rect 2127 11496 2173 11504
rect 4287 11496 4553 11504
rect 6536 11504 6544 11516
rect 8707 11516 8973 11524
rect 11087 11516 11733 11524
rect 5527 11496 6544 11504
rect 7367 11496 7953 11504
rect 9787 11496 10153 11504
rect 4447 11476 4693 11484
rect 5867 11476 6893 11484
rect 7407 11476 7573 11484
rect 7587 11476 7673 11484
rect 7767 11476 7913 11484
rect 8327 11476 8933 11484
rect 2727 11456 3233 11464
rect 4387 11456 4753 11464
rect 4767 11456 4933 11464
rect 4947 11456 5053 11464
rect 5447 11456 5673 11464
rect 8047 11456 9153 11464
rect 3627 11436 3884 11444
rect 467 11416 473 11424
rect 487 11416 693 11424
rect 707 11416 933 11424
rect 3876 11424 3884 11436
rect 3967 11436 4353 11444
rect 4396 11436 4724 11444
rect 4396 11424 4404 11436
rect 3876 11416 4404 11424
rect 4416 11416 4673 11424
rect 2907 11396 3213 11404
rect 4416 11404 4424 11416
rect 4716 11424 4724 11436
rect 5327 11436 5413 11444
rect 5427 11436 5853 11444
rect 6647 11436 7013 11444
rect 7027 11436 7073 11444
rect 10007 11436 10833 11444
rect 10847 11436 11813 11444
rect 11827 11436 11953 11444
rect 4716 11416 5173 11424
rect 5267 11416 5653 11424
rect 6187 11416 6373 11424
rect 7147 11416 7513 11424
rect 7527 11416 7633 11424
rect 9507 11416 10333 11424
rect 10347 11416 11293 11424
rect 3907 11396 4424 11404
rect 4707 11396 4873 11404
rect 4887 11396 5193 11404
rect 7967 11396 8453 11404
rect 10607 11396 10633 11404
rect 687 11376 793 11384
rect 1327 11376 1413 11384
rect 1427 11376 1593 11384
rect 4687 11376 5313 11384
rect 6267 11376 6553 11384
rect 7087 11376 7793 11384
rect 9227 11376 9273 11384
rect 9287 11376 9433 11384
rect 3227 11356 3693 11364
rect 3767 11356 4233 11364
rect 4247 11356 4304 11364
rect 567 11336 773 11344
rect 1047 11336 1193 11344
rect 1376 11336 1593 11344
rect 1376 11330 1384 11336
rect 3187 11336 3253 11344
rect 3307 11336 3613 11344
rect 4296 11344 4304 11356
rect 4347 11356 4533 11364
rect 5367 11356 5453 11364
rect 5467 11356 5833 11364
rect 6207 11356 6693 11364
rect 9867 11356 10553 11364
rect 10907 11356 11113 11364
rect 11127 11356 11353 11364
rect 11367 11356 11453 11364
rect 12047 11356 12153 11364
rect 4296 11336 4493 11344
rect 5067 11339 5113 11347
rect 6536 11336 6593 11344
rect 507 11319 613 11327
rect 1007 11319 1073 11327
rect 1287 11319 1373 11327
rect 1527 11319 1553 11327
rect 1667 11319 1733 11327
rect 1747 11319 1833 11327
rect 1927 11316 2033 11324
rect 2047 11319 2133 11327
rect 2187 11319 2233 11327
rect 2307 11319 2453 11327
rect 4147 11319 4273 11327
rect 5467 11319 5573 11327
rect 5627 11319 5693 11327
rect 5887 11319 5933 11327
rect 6127 11316 6293 11324
rect 247 11276 473 11284
rect 767 11273 873 11281
rect 927 11276 1013 11284
rect 1307 11276 1393 11284
rect 1587 11276 1893 11284
rect 2996 11284 3004 11316
rect 3467 11299 3593 11307
rect 3727 11293 3753 11301
rect 3996 11284 4004 11316
rect 4576 11304 4584 11316
rect 6307 11316 6333 11324
rect 6536 11324 6544 11336
rect 6607 11336 6673 11344
rect 7647 11336 7944 11344
rect 6347 11316 6544 11324
rect 6947 11316 7133 11324
rect 7827 11319 7873 11327
rect 7936 11324 7944 11336
rect 8507 11336 8593 11344
rect 8747 11339 9213 11347
rect 9787 11336 10213 11344
rect 11507 11336 11573 11344
rect 7936 11316 8013 11324
rect 8107 11319 8173 11327
rect 8187 11316 8653 11324
rect 9307 11319 9453 11327
rect 10047 11316 10092 11324
rect 10127 11316 10173 11324
rect 10187 11316 10273 11324
rect 10427 11319 10513 11327
rect 10527 11319 10593 11327
rect 10767 11319 10853 11327
rect 10967 11319 11093 11327
rect 11147 11316 11393 11324
rect 11407 11319 11433 11327
rect 11787 11316 11913 11324
rect 12027 11316 12153 11324
rect 4576 11296 4613 11304
rect 4707 11293 4733 11301
rect 2107 11276 2153 11284
rect 2427 11273 2493 11281
rect 2507 11276 2653 11284
rect 2907 11273 2973 11281
rect 2996 11276 3233 11284
rect 3736 11276 3973 11284
rect 3736 11264 3744 11276
rect 3996 11276 4253 11284
rect 4407 11276 4513 11284
rect 3607 11256 3744 11264
rect 4896 11264 4904 11296
rect 5027 11296 5093 11304
rect 7487 11299 7572 11307
rect 7607 11296 7693 11304
rect 8387 11296 8573 11304
rect 5607 11276 5653 11284
rect 5707 11276 5853 11284
rect 5927 11276 6353 11284
rect 6627 11276 6693 11284
rect 6987 11273 7173 11281
rect 7847 11276 7893 11284
rect 8667 11273 8693 11281
rect 8807 11276 8873 11284
rect 4896 11256 5013 11264
rect 5247 11256 5513 11264
rect 5567 11256 5933 11264
rect 5947 11256 6873 11264
rect 6887 11256 6953 11264
rect 7587 11256 7613 11264
rect 8447 11256 8533 11264
rect 1087 11236 1173 11244
rect 1187 11236 1333 11244
rect 1787 11236 1853 11244
rect 1867 11236 2013 11244
rect 3147 11236 3333 11244
rect 3667 11236 3833 11244
rect 4047 11236 4253 11244
rect 4307 11236 4413 11244
rect 4467 11236 4553 11244
rect 6727 11236 8133 11244
rect 8567 11236 8853 11244
rect 9056 11244 9064 11296
rect 9187 11296 9253 11304
rect 10647 11296 10673 11304
rect 10687 11296 11044 11304
rect 9427 11273 9513 11281
rect 9667 11273 9733 11281
rect 10067 11273 10113 11281
rect 10307 11273 10333 11281
rect 10487 11273 10533 11281
rect 10547 11276 11013 11284
rect 11036 11284 11044 11296
rect 11036 11276 11113 11284
rect 11607 11273 11633 11281
rect 11687 11276 11753 11284
rect 9187 11256 9293 11264
rect 9316 11256 9473 11264
rect 9316 11244 9324 11256
rect 10167 11256 10253 11264
rect 10267 11256 11053 11264
rect 12007 11256 12133 11264
rect 9056 11236 9324 11244
rect 10587 11236 10873 11244
rect 11587 11236 11633 11244
rect 11907 11236 12073 11244
rect 987 11216 1433 11224
rect 1447 11216 2193 11224
rect 3047 11216 4333 11224
rect 5087 11216 5473 11224
rect 5867 11216 6453 11224
rect 6467 11216 6513 11224
rect 8327 11216 8473 11224
rect 10827 11216 11213 11224
rect 4547 11196 4613 11204
rect 4627 11196 4913 11204
rect 5107 11196 5433 11204
rect 7187 11196 8093 11204
rect 8907 11196 9013 11204
rect 2147 11176 2233 11184
rect 2947 11176 3053 11184
rect 3607 11176 3893 11184
rect 5047 11176 5453 11184
rect 5507 11176 5573 11184
rect 6807 11176 6993 11184
rect 7227 11176 7333 11184
rect 9747 11176 10833 11184
rect 11127 11176 11433 11184
rect 11447 11176 11673 11184
rect 1047 11156 1153 11164
rect 3187 11156 4073 11164
rect 5767 11156 6073 11164
rect 6507 11156 7204 11164
rect 487 11136 573 11144
rect 767 11136 1253 11144
rect 1267 11136 1613 11144
rect 1627 11136 1713 11144
rect 1847 11136 1993 11144
rect 4727 11136 4873 11144
rect 5367 11136 5493 11144
rect 6107 11136 6473 11144
rect 7196 11144 7204 11156
rect 8167 11156 8493 11164
rect 8887 11156 9053 11164
rect 10727 11156 10984 11164
rect 7196 11136 7273 11144
rect 8087 11136 8133 11144
rect 9567 11136 10953 11144
rect 10976 11144 10984 11156
rect 10976 11136 11213 11144
rect 11227 11136 11373 11144
rect 2487 11116 2673 11124
rect 3627 11116 3693 11124
rect 10067 11116 10224 11124
rect 187 11099 233 11107
rect 627 11096 693 11104
rect 707 11099 753 11107
rect 807 11096 1073 11104
rect 1087 11099 1113 11107
rect 1307 11099 1393 11107
rect 1607 11096 1833 11104
rect 1887 11099 1913 11107
rect 1967 11096 2093 11104
rect 2107 11099 2233 11107
rect 2327 11099 2353 11107
rect 2407 11096 2453 11104
rect 3187 11096 3213 11104
rect 3287 11096 3313 11104
rect 3476 11096 3573 11104
rect 2627 11073 2893 11081
rect 3136 11076 3153 11084
rect 3476 11084 3484 11096
rect 3867 11099 3933 11107
rect 3947 11099 3953 11107
rect 4007 11096 4173 11104
rect 4227 11099 4293 11107
rect 4347 11096 4453 11104
rect 4767 11099 4793 11107
rect 4907 11099 5233 11107
rect 5447 11099 5753 11107
rect 5807 11096 5992 11104
rect 6027 11099 6133 11107
rect 6327 11096 6393 11104
rect 6987 11096 7093 11104
rect 7547 11099 7573 11107
rect 7907 11099 7993 11107
rect 8227 11096 8373 11104
rect 9027 11099 9133 11107
rect 227 11056 413 11064
rect 787 11056 973 11064
rect 1167 11053 1313 11061
rect 1727 11053 1813 11061
rect 1867 11053 1953 11061
rect 2007 11053 2113 11061
rect 3136 11064 3144 11076
rect 3607 11076 3673 11084
rect 6480 11084 6493 11087
rect 6476 11073 6493 11084
rect 2467 11053 2693 11061
rect 2707 11056 3144 11064
rect 3947 11056 3993 11064
rect 4087 11053 4153 11061
rect 4507 11056 4733 11064
rect 4747 11053 5053 11061
rect 5127 11056 5273 11064
rect 5407 11053 5773 11061
rect 6007 11053 6073 11061
rect 6347 11053 6413 11061
rect 6476 11047 6484 11073
rect 6587 11073 6713 11081
rect 6847 11076 6913 11084
rect 6967 11056 7353 11064
rect 7367 11056 7533 11064
rect 8416 11064 8424 11096
rect 9267 11096 9453 11104
rect 9507 11099 9553 11107
rect 9927 11096 9953 11104
rect 9967 11099 10073 11107
rect 10216 11104 10224 11116
rect 10216 11096 10253 11104
rect 10267 11099 10393 11107
rect 10967 11099 11013 11107
rect 11467 11099 11533 11107
rect 11776 11106 11813 11107
rect 11787 11099 11813 11106
rect 12107 11096 12293 11104
rect 8627 11073 8753 11081
rect 8887 11076 8953 11084
rect 7667 11056 7873 11064
rect 8127 11056 8353 11064
rect 8416 11056 8453 11064
rect 9447 11053 10052 11061
rect 10087 11056 10233 11064
rect 10247 11056 10493 11064
rect 10787 11053 10813 11061
rect 11287 11056 11453 11064
rect 11607 11056 11773 11064
rect 11847 11056 12073 11064
rect 2427 11036 2473 11044
rect 2547 11033 2733 11041
rect 3247 11036 3633 11044
rect 3647 11033 3693 11041
rect 4267 11036 4433 11044
rect 6887 11033 6933 11041
rect 9067 11036 9173 11044
rect 9487 11036 9713 11044
rect 3807 11016 4533 11024
rect 5027 11016 5193 11024
rect 5207 11016 6113 11024
rect 6127 11016 6313 11024
rect 7667 11016 7953 11024
rect 8007 11016 8253 11024
rect 8613 11024 8627 11033
rect 8407 11020 8627 11024
rect 8407 11016 8624 11020
rect 10467 11016 10953 11024
rect 11247 11016 11293 11024
rect 11847 11016 11893 11024
rect 11967 11016 12113 11024
rect 1067 10996 1393 11004
rect 2047 10996 2153 11004
rect 2727 10996 3313 11004
rect 3927 10996 4193 11004
rect 4207 10996 4493 11004
rect 5067 10996 5393 11004
rect 8887 10996 8913 11004
rect 8927 10996 9273 11004
rect 847 10976 1073 10984
rect 1127 10976 1273 10984
rect 1287 10976 1373 10984
rect 1387 10976 1453 10984
rect 1467 10976 1913 10984
rect 1927 10976 2073 10984
rect 2087 10976 2273 10984
rect 4307 10976 4793 10984
rect 4807 10976 5373 10984
rect 5387 10976 5533 10984
rect 8467 10976 8733 10984
rect 11047 10976 11313 10984
rect 12107 10976 12173 10984
rect 3987 10956 4853 10964
rect 4867 10956 5073 10964
rect 5267 10956 5353 10964
rect 5687 10956 6153 10964
rect 8156 10956 8244 10964
rect 587 10936 2373 10944
rect 3327 10936 3853 10944
rect 4027 10936 4513 10944
rect 4527 10936 5153 10944
rect 5167 10936 6113 10944
rect 6127 10936 6173 10944
rect 8156 10944 8164 10956
rect 7607 10936 8164 10944
rect 8236 10944 8244 10956
rect 8987 10956 9473 10964
rect 9727 10956 10773 10964
rect 8236 10936 8633 10944
rect 8647 10936 8753 10944
rect 8767 10936 9653 10944
rect 4707 10916 5332 10924
rect 5367 10916 5493 10924
rect 5507 10916 5913 10924
rect 7127 10916 8213 10924
rect 8267 10916 8433 10924
rect 8747 10916 9253 10924
rect 9887 10916 11233 10924
rect 2327 10896 2353 10904
rect 2367 10896 2653 10904
rect 3647 10896 3773 10904
rect 3967 10896 4193 10904
rect 6167 10896 6733 10904
rect 6747 10896 6873 10904
rect 6947 10896 7813 10904
rect 8787 10896 9153 10904
rect 11087 10896 11572 10904
rect 11607 10896 11633 10904
rect 2927 10876 3053 10884
rect 4433 10884 4447 10893
rect 4433 10880 4933 10884
rect 4436 10876 4933 10880
rect 5047 10876 5433 10884
rect 5447 10876 5473 10884
rect 5896 10876 5993 10884
rect 5896 10864 5904 10876
rect 8747 10876 10013 10884
rect 10307 10876 10413 10884
rect 10427 10876 10633 10884
rect 5627 10856 5904 10864
rect 5996 10856 6033 10864
rect 327 10836 553 10844
rect 3487 10836 3593 10844
rect 3687 10836 3753 10844
rect 5307 10836 5433 10844
rect 5996 10844 6004 10856
rect 7047 10856 10133 10864
rect 10847 10856 11253 10864
rect 6180 10844 6193 10847
rect 5976 10840 6004 10844
rect 5973 10836 6004 10840
rect 827 10816 853 10824
rect 1087 10816 1213 10824
rect 1707 10819 2533 10827
rect 5973 10827 5987 10836
rect 6176 10833 6193 10844
rect 6667 10836 6973 10844
rect 7507 10836 8113 10844
rect 8607 10836 8773 10844
rect 9227 10836 9413 10844
rect 9467 10836 9753 10844
rect 10547 10836 10733 10844
rect 10747 10836 10813 10844
rect 11387 10836 11633 10844
rect 2547 10816 2573 10824
rect 2767 10816 3293 10824
rect 4967 10816 5093 10824
rect 5527 10816 5844 10824
rect 507 10799 533 10807
rect 1547 10799 1573 10807
rect 1316 10784 1324 10796
rect 2327 10796 2613 10804
rect 2627 10796 2713 10804
rect 3076 10796 3333 10804
rect 1316 10776 1413 10784
rect 687 10756 833 10764
rect 1347 10756 1513 10764
rect 1656 10764 1664 10793
rect 3076 10790 3084 10796
rect 3387 10796 3713 10804
rect 3756 10796 4013 10804
rect 196 10744 204 10749
rect 196 10736 633 10744
rect 1516 10744 1524 10753
rect 1647 10756 1664 10764
rect 1856 10764 1864 10776
rect 2127 10773 2173 10781
rect 3207 10776 3273 10784
rect 3756 10784 3764 10796
rect 3736 10776 3764 10784
rect 4296 10784 4304 10796
rect 4887 10796 5213 10804
rect 5227 10796 5333 10804
rect 5487 10800 5704 10804
rect 5487 10796 5707 10800
rect 4296 10776 4393 10784
rect 1856 10756 2033 10764
rect 2407 10756 2493 10764
rect 2727 10756 2873 10764
rect 3736 10764 3744 10776
rect 4547 10779 4753 10787
rect 5693 10787 5707 10796
rect 5836 10790 5844 10816
rect 4807 10773 4833 10781
rect 6016 10787 6024 10813
rect 6116 10787 6124 10813
rect 6176 10787 6184 10833
rect 7187 10819 8693 10827
rect 9127 10816 9433 10824
rect 9487 10816 9573 10824
rect 11207 10816 11533 10824
rect 6787 10796 6833 10804
rect 6327 10779 6452 10787
rect 6487 10773 6513 10781
rect 6587 10773 6653 10781
rect 3987 10756 4033 10764
rect 4327 10753 4693 10761
rect 5087 10753 5253 10761
rect 5327 10756 5533 10764
rect 7096 10764 7104 10796
rect 7116 10764 7124 10813
rect 7147 10796 7164 10804
rect 7887 10796 8053 10804
rect 7156 10767 7164 10796
rect 7816 10784 7824 10796
rect 8076 10796 8173 10804
rect 8187 10799 8233 10807
rect 8076 10784 8084 10796
rect 8287 10796 8393 10804
rect 8407 10796 8453 10804
rect 7816 10776 8084 10784
rect 8676 10784 8684 10796
rect 8807 10796 8913 10804
rect 10267 10799 10433 10807
rect 10607 10799 10713 10807
rect 10867 10799 10893 10807
rect 11027 10799 11073 10807
rect 11807 10799 11873 10807
rect 12067 10799 12173 10807
rect 12227 10799 12273 10807
rect 8676 10776 9244 10784
rect 7076 10760 7104 10764
rect 7073 10756 7104 10760
rect 7073 10747 7087 10756
rect 7336 10764 7344 10776
rect 7336 10756 7493 10764
rect 9236 10764 9244 10776
rect 11447 10776 11773 10784
rect 11916 10784 11924 10796
rect 11787 10776 11924 10784
rect 8167 10753 8273 10761
rect 8707 10753 8793 10761
rect 9467 10756 9533 10764
rect 9587 10756 9693 10764
rect 9747 10756 9993 10764
rect 10047 10756 10273 10764
rect 10327 10756 10453 10764
rect 10467 10756 10673 10764
rect 10687 10753 10793 10761
rect 11287 10753 11353 10761
rect 1516 10736 1593 10744
rect 2067 10736 2313 10744
rect 5687 10736 5973 10744
rect 6047 10736 6513 10744
rect 7547 10736 7773 10744
rect 7787 10736 7813 10744
rect 8427 10736 8613 10744
rect 9187 10736 9213 10744
rect 10847 10736 10933 10744
rect 11327 10736 11653 10744
rect 11747 10736 11813 10744
rect 11827 10736 11893 10744
rect 11947 10736 12053 10744
rect 12107 10736 12153 10744
rect 2087 10716 2153 10724
rect 2687 10716 3193 10724
rect 3567 10716 3773 10724
rect 4127 10716 4293 10724
rect 4407 10716 5133 10724
rect 6487 10716 7053 10724
rect 9247 10716 9873 10724
rect 10287 10716 10393 10724
rect 12227 10716 12273 10724
rect 567 10696 593 10704
rect 907 10696 1093 10704
rect 1507 10696 2373 10704
rect 2667 10696 3144 10704
rect 3136 10687 3144 10696
rect 3347 10696 3404 10704
rect 1307 10676 1373 10684
rect 2047 10676 2673 10684
rect 2927 10676 2973 10684
rect 3136 10676 3153 10687
rect 3140 10673 3153 10676
rect 3167 10676 3313 10684
rect 3396 10684 3404 10696
rect 3887 10696 5193 10704
rect 5527 10696 5593 10704
rect 6047 10696 6173 10704
rect 7147 10696 7213 10704
rect 7607 10696 7953 10704
rect 10587 10696 11213 10704
rect 11607 10696 11993 10704
rect 3396 10676 4493 10684
rect 4847 10676 5333 10684
rect 5987 10676 6193 10684
rect 6827 10676 7553 10684
rect 8067 10676 8553 10684
rect 8947 10676 9253 10684
rect 9267 10676 9913 10684
rect 10847 10676 10993 10684
rect 11247 10676 12193 10684
rect 507 10656 553 10664
rect 627 10656 693 10664
rect 707 10656 1013 10664
rect 2827 10656 3373 10664
rect 3387 10656 4173 10664
rect 5367 10656 5513 10664
rect 5527 10656 5553 10664
rect 5687 10656 5753 10664
rect 6327 10656 6513 10664
rect 6527 10656 6713 10664
rect 7267 10656 7513 10664
rect 8127 10656 8253 10664
rect 11267 10656 12073 10664
rect 2887 10636 3073 10644
rect 3747 10636 3893 10644
rect 4207 10636 4633 10644
rect 4827 10636 4973 10644
rect 4987 10636 5273 10644
rect 5427 10636 5773 10644
rect 6827 10636 6853 10644
rect 7507 10636 7873 10644
rect 8247 10636 9433 10644
rect 11327 10636 11793 10644
rect 12167 10636 12253 10644
rect 247 10616 773 10624
rect 947 10616 1313 10624
rect 1847 10616 2233 10624
rect 2507 10616 2793 10624
rect 3787 10616 3813 10624
rect 4767 10616 5184 10624
rect 4267 10596 4613 10604
rect 4667 10596 4953 10604
rect 5047 10596 5153 10604
rect 5176 10604 5184 10616
rect 5347 10616 5413 10624
rect 5467 10616 5593 10624
rect 5827 10616 5913 10624
rect 6147 10616 6933 10624
rect 8327 10616 8713 10624
rect 9587 10616 10013 10624
rect 10447 10616 10893 10624
rect 5176 10596 5633 10604
rect 6007 10596 6173 10604
rect 10067 10596 10093 10604
rect 247 10576 473 10584
rect 527 10579 613 10587
rect 667 10576 733 10584
rect 867 10579 993 10587
rect 1367 10577 1493 10584
rect 1356 10576 1493 10577
rect 1507 10576 1573 10584
rect 2127 10579 2193 10587
rect 2447 10576 2633 10584
rect 2767 10579 2873 10587
rect 2947 10579 3033 10587
rect 3267 10576 3453 10584
rect 2007 10556 2293 10564
rect 707 10533 793 10541
rect 1427 10536 1813 10544
rect 2367 10533 2433 10541
rect 2627 10533 2893 10541
rect 2967 10533 3173 10541
rect 3327 10533 3473 10541
rect 3527 10533 3713 10541
rect 3776 10527 3784 10576
rect 4416 10586 4453 10587
rect 3907 10576 3964 10584
rect 3956 10564 3964 10576
rect 4427 10579 4453 10586
rect 4567 10576 4773 10584
rect 5087 10576 5153 10584
rect 5287 10579 5313 10587
rect 5367 10576 5553 10584
rect 5707 10579 5793 10587
rect 5807 10579 5873 10587
rect 6927 10579 7053 10587
rect 7107 10576 7153 10584
rect 7207 10576 7273 10584
rect 7407 10579 7433 10587
rect 7487 10576 7533 10584
rect 7607 10579 7753 10587
rect 7767 10576 7904 10584
rect 8227 10576 8513 10584
rect 8847 10576 9073 10584
rect 9127 10579 9233 10587
rect 9367 10579 9493 10587
rect 9627 10579 9653 10587
rect 10127 10576 10253 10584
rect 3956 10556 4073 10564
rect 3836 10527 3844 10553
rect 4207 10556 4353 10564
rect 6176 10556 6253 10564
rect 7896 10564 7904 10576
rect 10327 10579 10413 10587
rect 10987 10576 11173 10584
rect 11227 10579 11273 10587
rect 11367 10579 11413 10587
rect 11427 10576 11493 10584
rect 11627 10576 11673 10584
rect 11807 10579 11933 10587
rect 4527 10533 4553 10541
rect 4807 10533 4853 10541
rect 4867 10536 5233 10544
rect 5033 10527 5047 10536
rect 5247 10536 5333 10544
rect 5387 10533 5413 10541
rect 5507 10533 5613 10541
rect 6176 10544 6184 10556
rect 6367 10553 6513 10561
rect 7896 10556 8433 10564
rect 5967 10536 6184 10544
rect 6807 10536 7013 10544
rect 7067 10536 7213 10544
rect 7227 10536 7453 10544
rect 7567 10536 7733 10544
rect 7987 10536 8193 10544
rect 8427 10536 8533 10544
rect 8587 10533 8733 10541
rect 9107 10536 9333 10544
rect 9547 10536 9593 10544
rect 10107 10533 10173 10541
rect 10267 10533 10353 10541
rect 10407 10533 10453 10541
rect 10467 10536 10533 10544
rect 10667 10536 10873 10544
rect 10927 10533 10973 10541
rect 11167 10533 11253 10541
rect 11387 10536 11433 10544
rect 11707 10533 11733 10541
rect 11967 10533 12013 10541
rect 12027 10536 12233 10544
rect 567 10516 1013 10524
rect 1467 10516 1593 10524
rect 3776 10516 3793 10527
rect 3780 10513 3793 10516
rect 6047 10516 6193 10524
rect 7407 10516 7433 10524
rect 7487 10516 7973 10524
rect 8287 10516 8813 10524
rect 9847 10516 11293 10524
rect 11307 10516 11653 10524
rect 1927 10496 2753 10504
rect 2927 10496 3433 10504
rect 4707 10496 4913 10504
rect 4927 10496 5093 10504
rect 5187 10496 5413 10504
rect 5567 10496 5653 10504
rect 6107 10496 6153 10504
rect 6167 10496 6193 10504
rect 6827 10496 7613 10504
rect 7727 10496 9673 10504
rect 10027 10496 10913 10504
rect 11427 10496 11613 10504
rect 1247 10476 1333 10484
rect 2367 10476 2473 10484
rect 3607 10476 3753 10484
rect 3767 10476 3813 10484
rect 3887 10476 4273 10484
rect 5067 10476 5133 10484
rect 5287 10476 5333 10484
rect 5607 10476 5893 10484
rect 6836 10476 7272 10484
rect 507 10456 973 10464
rect 987 10456 1453 10464
rect 1827 10456 1913 10464
rect 2287 10456 5553 10464
rect 6836 10464 6844 10476
rect 7307 10476 7673 10484
rect 7867 10476 8472 10484
rect 8507 10476 8913 10484
rect 9067 10476 9153 10484
rect 9676 10484 9684 10493
rect 9676 10476 11073 10484
rect 11087 10476 11353 10484
rect 11967 10476 12193 10484
rect 6087 10456 6844 10464
rect 7207 10456 7493 10464
rect 7887 10456 8233 10464
rect 10487 10456 11033 10464
rect 2187 10436 2913 10444
rect 3307 10436 4593 10444
rect 5447 10436 5813 10444
rect 6307 10436 6953 10444
rect 7087 10436 7473 10444
rect 8027 10436 8193 10444
rect 8527 10436 9653 10444
rect 11227 10436 11773 10444
rect 11787 10436 11913 10444
rect 467 10416 553 10424
rect 1827 10416 2093 10424
rect 3327 10416 3773 10424
rect 3947 10416 4073 10424
rect 4087 10416 4233 10424
rect 4727 10416 5213 10424
rect 5547 10416 6353 10424
rect 6687 10416 6733 10424
rect 7527 10416 8493 10424
rect 8516 10416 10853 10424
rect 767 10396 853 10404
rect 1107 10396 1673 10404
rect 3987 10396 4413 10404
rect 5567 10396 6293 10404
rect 7887 10396 8033 10404
rect 8516 10404 8524 10416
rect 11107 10416 11373 10424
rect 8487 10396 8524 10404
rect 10227 10396 10573 10404
rect 10587 10396 10653 10404
rect 11047 10396 11473 10404
rect 2387 10376 2713 10384
rect 3967 10376 4084 10384
rect 1547 10356 2053 10364
rect 2407 10356 2453 10364
rect 4076 10364 4084 10376
rect 4487 10376 4553 10384
rect 4567 10376 4753 10384
rect 4767 10376 4873 10384
rect 5207 10376 5373 10384
rect 5387 10376 5573 10384
rect 6967 10376 7253 10384
rect 7327 10376 7653 10384
rect 8087 10376 8173 10384
rect 8467 10376 8573 10384
rect 8627 10376 9093 10384
rect 9107 10376 9953 10384
rect 10887 10376 11393 10384
rect 4076 10356 4813 10364
rect 4947 10356 5393 10364
rect 10727 10356 10793 10364
rect 11187 10356 11693 10364
rect 3167 10336 3253 10344
rect 3927 10336 4013 10344
rect 6167 10336 6793 10344
rect 7487 10336 7853 10344
rect 227 10316 273 10324
rect 327 10316 773 10324
rect 2287 10316 2753 10324
rect 2767 10316 3053 10324
rect 3687 10316 3893 10324
rect 4096 10316 4097 10324
rect 4111 10324 4120 10327
rect 4111 10313 4124 10324
rect 4887 10316 6073 10324
rect 6787 10316 6833 10324
rect 7227 10316 7453 10324
rect 8207 10316 8253 10324
rect 2547 10296 2993 10304
rect 3627 10296 3653 10304
rect 247 10279 353 10287
rect 407 10279 513 10287
rect 567 10279 933 10287
rect 1027 10279 1053 10287
rect 1107 10279 1153 10287
rect 1587 10279 1653 10287
rect 1887 10279 1973 10287
rect 2127 10279 2153 10287
rect 2247 10279 2373 10287
rect 307 10233 393 10241
rect 807 10236 853 10244
rect 1367 10233 1653 10241
rect 1987 10236 2453 10244
rect 2476 10227 2484 10276
rect 2947 10276 2973 10284
rect 3047 10276 3133 10284
rect 3147 10279 3213 10287
rect 2516 10244 2524 10273
rect 3487 10259 3633 10267
rect 4076 10267 4084 10296
rect 3747 10253 3833 10261
rect 4076 10256 4092 10267
rect 4080 10253 4092 10256
rect 4116 10264 4124 10313
rect 5247 10296 5593 10304
rect 7827 10304 7840 10307
rect 7827 10293 7844 10304
rect 4947 10279 5073 10287
rect 5627 10279 5653 10287
rect 4247 10259 4413 10267
rect 4796 10264 4804 10276
rect 5776 10286 5853 10287
rect 5707 10276 5773 10284
rect 5787 10279 5853 10286
rect 5907 10279 5933 10287
rect 5987 10276 6153 10284
rect 6296 10276 6693 10284
rect 6296 10264 6304 10276
rect 4796 10256 5044 10264
rect 2507 10236 2524 10244
rect 2667 10236 2733 10244
rect 3067 10236 3233 10244
rect 3947 10233 4033 10241
rect 4607 10236 4713 10244
rect 5036 10244 5044 10256
rect 6347 10259 6493 10267
rect 6776 10264 6784 10276
rect 7087 10276 7133 10284
rect 7347 10279 7413 10287
rect 7567 10276 7713 10284
rect 7836 10264 7844 10293
rect 6687 10256 6784 10264
rect 8176 10267 8184 10293
rect 8416 10270 8424 10353
rect 9707 10336 10353 10344
rect 10707 10336 11164 10344
rect 11156 10324 11164 10336
rect 11156 10316 11313 10324
rect 12087 10316 12213 10324
rect 8667 10296 9033 10304
rect 10107 10296 10953 10304
rect 8727 10276 8873 10284
rect 10607 10279 10693 10287
rect 10747 10279 10773 10287
rect 11107 10276 11193 10284
rect 11467 10276 11513 10284
rect 11967 10276 12013 10284
rect 4987 10233 5013 10241
rect 5036 10236 5053 10244
rect 5267 10236 5293 10244
rect 5487 10236 5693 10244
rect 5807 10233 5833 10241
rect 6027 10236 6253 10244
rect 6907 10233 7013 10241
rect 7187 10236 7213 10244
rect 7267 10236 7433 10244
rect 7687 10236 7773 10244
rect 8036 10244 8044 10256
rect 9887 10256 10033 10264
rect 10047 10256 10164 10264
rect 8036 10236 8273 10244
rect 10156 10244 10164 10256
rect 8707 10236 8893 10244
rect 9107 10233 9133 10241
rect 9187 10236 9413 10244
rect 9947 10233 10013 10241
rect 10167 10233 10193 10241
rect 10367 10233 10453 10241
rect 11207 10233 11233 10241
rect 11407 10233 11433 10241
rect 11696 10227 11704 10276
rect 12147 10279 12253 10287
rect 11727 10233 11833 10241
rect 11847 10233 11873 10241
rect 11987 10236 12133 10244
rect 2227 10216 2273 10224
rect 2767 10216 2953 10224
rect 3187 10216 3353 10224
rect 3627 10216 3693 10224
rect 4447 10216 4533 10224
rect 4687 10216 4933 10224
rect 7127 10216 7193 10224
rect 10987 10216 11273 10224
rect 11876 10224 11884 10230
rect 11876 10216 12193 10224
rect 367 10196 533 10204
rect 647 10196 753 10204
rect 767 10196 1073 10204
rect 1327 10196 1733 10204
rect 1927 10196 2053 10204
rect 2187 10196 2313 10204
rect 3647 10196 3813 10204
rect 3987 10196 4393 10204
rect 5447 10196 5513 10204
rect 5527 10196 5553 10204
rect 5767 10196 5793 10204
rect 5847 10196 5873 10204
rect 7067 10196 7533 10204
rect 7607 10196 7693 10204
rect 8647 10196 8773 10204
rect 9467 10196 9493 10204
rect 9507 10196 10213 10204
rect 2467 10176 2533 10184
rect 4427 10176 4773 10184
rect 5347 10176 5693 10184
rect 5947 10176 6153 10184
rect 6167 10176 6233 10184
rect 8227 10176 9733 10184
rect 9747 10176 9933 10184
rect 10247 10176 10273 10184
rect 10287 10176 10493 10184
rect 11667 10176 11813 10184
rect 12147 10176 12313 10184
rect 3047 10156 3133 10164
rect 3147 10156 4873 10164
rect 5227 10156 5273 10164
rect 5607 10156 6333 10164
rect 7447 10156 7673 10164
rect 10567 10156 10773 10164
rect 11687 10156 11933 10164
rect 2567 10136 2633 10144
rect 3967 10136 4093 10144
rect 5167 10136 5333 10144
rect 10967 10136 11173 10144
rect 11527 10136 12093 10144
rect 2507 10116 2793 10124
rect 4507 10116 4673 10124
rect 6767 10116 6913 10124
rect 6927 10116 7133 10124
rect 8167 10116 8233 10124
rect 8247 10116 8293 10124
rect 8387 10116 8753 10124
rect 8767 10116 8893 10124
rect 10727 10116 10833 10124
rect 10847 10116 10873 10124
rect 267 10096 533 10104
rect 547 10096 753 10104
rect 1787 10096 1893 10104
rect 3207 10096 3673 10104
rect 5267 10096 5593 10104
rect 5727 10096 6093 10104
rect 6247 10096 6933 10104
rect 7047 10096 7093 10104
rect 7507 10096 7824 10104
rect 1447 10076 1533 10084
rect 1547 10076 1753 10084
rect 2587 10076 2733 10084
rect 4107 10076 4264 10084
rect 247 10056 453 10064
rect 1307 10059 1413 10067
rect 496 10007 504 10056
rect 1787 10064 1800 10067
rect 1787 10053 1804 10064
rect 1887 10056 1953 10064
rect 1967 10056 2053 10064
rect 2147 10056 2213 10064
rect 2227 10056 2553 10064
rect 2707 10056 3073 10064
rect 3867 10059 3973 10067
rect 4027 10059 4053 10067
rect 907 10013 1013 10021
rect 1027 10016 1113 10024
rect 1167 10016 1313 10024
rect 1796 10024 1804 10053
rect 3147 10039 3233 10047
rect 3527 10036 3613 10044
rect 4136 10040 4213 10044
rect 4133 10036 4213 10040
rect 4256 10044 4264 10076
rect 4507 10076 4553 10084
rect 6187 10076 6213 10084
rect 7816 10084 7824 10096
rect 7847 10096 8013 10104
rect 8927 10096 9093 10104
rect 9947 10096 10433 10104
rect 10447 10096 10824 10104
rect 7816 10076 7913 10084
rect 9707 10076 9893 10084
rect 10007 10076 10553 10084
rect 10816 10084 10824 10096
rect 10867 10096 10993 10104
rect 11407 10096 11533 10104
rect 11627 10096 12053 10104
rect 10816 10076 11013 10084
rect 11287 10076 11313 10084
rect 11327 10076 11793 10084
rect 4787 10056 4833 10064
rect 5467 10059 5553 10067
rect 5787 10059 6393 10067
rect 6547 10056 6613 10064
rect 6967 10056 7013 10064
rect 7247 10056 7352 10064
rect 7387 10056 7453 10064
rect 7467 10059 7553 10067
rect 7767 10059 7793 10067
rect 7816 10056 7973 10064
rect 7987 10059 8173 10067
rect 8347 10059 8393 10067
rect 8507 10059 8533 10067
rect 8747 10059 8773 10067
rect 8796 10056 8813 10064
rect 4256 10036 4333 10044
rect 1427 10016 1553 10024
rect 2587 10013 2693 10021
rect 3047 10013 3093 10021
rect 1847 9996 1873 10004
rect 2087 9996 2473 10004
rect 3396 10004 3404 10030
rect 4133 10027 4147 10036
rect 4607 10036 4784 10044
rect 4536 10007 4544 10036
rect 4707 10016 4753 10024
rect 4776 10024 4784 10036
rect 4776 10016 4813 10024
rect 4896 10007 4904 10033
rect 5087 10033 5253 10041
rect 5307 10036 5493 10044
rect 7816 10044 7824 10056
rect 7147 10036 7824 10044
rect 5627 10013 5653 10021
rect 5707 10013 5833 10021
rect 5967 10016 6093 10024
rect 6267 10016 6413 10024
rect 6527 10013 6653 10021
rect 6787 10016 6933 10024
rect 6947 10013 7033 10021
rect 7367 10013 7513 10021
rect 8796 10024 8804 10056
rect 8887 10056 9093 10064
rect 9136 10024 9144 10056
rect 9287 10056 9333 10064
rect 9547 10059 9573 10067
rect 9627 10056 9833 10064
rect 9987 10059 10673 10067
rect 10807 10056 11133 10064
rect 11147 10056 11253 10064
rect 11427 10056 11553 10064
rect 11867 10056 12033 10064
rect 8407 10016 8553 10024
rect 8776 10020 8804 10024
rect 8773 10016 8804 10020
rect 8773 10007 8787 10016
rect 9047 10013 9073 10021
rect 9136 10016 9193 10024
rect 9207 10016 9353 10024
rect 9847 10013 9873 10021
rect 9927 10013 10073 10021
rect 10227 10016 10453 10024
rect 11367 10016 11693 10024
rect 11707 10013 11733 10021
rect 3396 9996 3533 10004
rect 3807 9996 3993 10004
rect 4527 9996 4544 10007
rect 4527 9993 4540 9996
rect 4567 9996 4713 10004
rect 6487 9996 7573 10004
rect 8007 9996 8273 10004
rect 8327 9996 8373 10004
rect 9647 9996 10133 10004
rect 11827 9996 12073 10004
rect 227 9976 453 9984
rect 467 9976 513 9984
rect 2027 9976 2113 9984
rect 2307 9976 2333 9984
rect 2347 9976 2373 9984
rect 2607 9976 2913 9984
rect 3027 9976 3193 9984
rect 4607 9976 4633 9984
rect 6707 9976 7012 9984
rect 7047 9976 7553 9984
rect 9307 9976 10393 9984
rect 10527 9976 10933 9984
rect 11287 9976 11533 9984
rect 11547 9976 11593 9984
rect 3567 9956 3953 9964
rect 3967 9956 4033 9964
rect 4087 9956 4853 9964
rect 4867 9956 5573 9964
rect 5587 9956 5873 9964
rect 7407 9956 8213 9964
rect 9347 9956 10193 9964
rect 4036 9944 4044 9953
rect 4036 9936 4173 9944
rect 4747 9936 5473 9944
rect 5927 9936 6173 9944
rect 6187 9936 7153 9944
rect 7447 9936 8493 9944
rect 9687 9936 10993 9944
rect 11007 9936 11193 9944
rect 11207 9936 11673 9944
rect 3947 9916 4073 9924
rect 7627 9916 7693 9924
rect 8047 9916 8793 9924
rect 8907 9916 9113 9924
rect 9127 9916 9333 9924
rect 9467 9916 9624 9924
rect 267 9896 293 9904
rect 627 9896 993 9904
rect 1007 9896 1093 9904
rect 1107 9896 1613 9904
rect 1627 9896 1793 9904
rect 2207 9896 2573 9904
rect 3067 9896 3613 9904
rect 3627 9896 3673 9904
rect 3847 9896 3893 9904
rect 4127 9896 4773 9904
rect 5007 9896 5233 9904
rect 5687 9896 5973 9904
rect 6047 9896 9593 9904
rect 9616 9904 9624 9916
rect 9827 9916 10172 9924
rect 10207 9916 10713 9924
rect 10767 9916 10973 9924
rect 10987 9916 11493 9924
rect 11507 9916 11613 9924
rect 9616 9896 11773 9904
rect 11987 9896 12073 9904
rect 1947 9876 2173 9884
rect 2187 9876 2533 9884
rect 2547 9876 2873 9884
rect 2887 9876 7053 9884
rect 7187 9876 7373 9884
rect 8127 9876 9273 9884
rect 10247 9876 11233 9884
rect 11247 9876 11413 9884
rect 1227 9856 1853 9864
rect 2327 9856 2653 9864
rect 2667 9856 2833 9864
rect 2947 9856 3073 9864
rect 3887 9856 3953 9864
rect 4007 9856 4493 9864
rect 5227 9856 5713 9864
rect 6587 9856 7044 9864
rect 707 9836 1633 9844
rect 2727 9836 2773 9844
rect 3427 9836 3693 9844
rect 3707 9836 3753 9844
rect 3987 9836 4533 9844
rect 4687 9836 5253 9844
rect 5347 9836 5673 9844
rect 7036 9844 7044 9856
rect 7647 9856 7672 9864
rect 7707 9856 7993 9864
rect 9247 9856 9953 9864
rect 9967 9856 10093 9864
rect 7036 9836 7233 9844
rect 9767 9836 10453 9844
rect 10467 9836 10613 9844
rect 10627 9836 11193 9844
rect 11907 9836 12233 9844
rect 1667 9816 5324 9824
rect 1387 9796 1453 9804
rect 1467 9796 1593 9804
rect 2487 9796 2713 9804
rect 2787 9796 2904 9804
rect 2587 9776 2732 9784
rect 267 9759 433 9767
rect 487 9759 573 9767
rect 787 9756 873 9764
rect 196 9727 204 9753
rect 507 9716 693 9724
rect 736 9707 744 9756
rect 987 9759 1033 9767
rect 1047 9756 1113 9764
rect 1507 9759 1553 9767
rect 1647 9759 1893 9767
rect 1907 9756 2373 9764
rect 1276 9744 1284 9756
rect 1236 9736 1284 9744
rect 2416 9744 2424 9756
rect 2416 9736 2684 9744
rect 1236 9727 1244 9736
rect 1027 9716 1233 9724
rect 2676 9724 2684 9736
rect 2696 9724 2704 9756
rect 2756 9747 2764 9773
rect 2896 9750 2904 9796
rect 3796 9796 4013 9804
rect 3796 9787 3804 9796
rect 4367 9796 4713 9804
rect 5207 9796 5293 9804
rect 5316 9804 5324 9816
rect 5527 9816 5833 9824
rect 6347 9816 6833 9824
rect 6847 9816 7393 9824
rect 7927 9816 9053 9824
rect 9067 9816 9553 9824
rect 5316 9796 6233 9804
rect 6987 9796 7273 9804
rect 7447 9796 7553 9804
rect 7607 9796 7813 9804
rect 7827 9796 8033 9804
rect 10087 9796 10353 9804
rect 10367 9796 10393 9804
rect 10507 9796 11353 9804
rect 11647 9796 11913 9804
rect 11927 9796 11993 9804
rect 3047 9776 3073 9784
rect 3527 9776 3693 9784
rect 3707 9776 3793 9784
rect 4767 9776 5333 9784
rect 6107 9776 6213 9784
rect 7287 9776 7333 9784
rect 8100 9784 8113 9787
rect 8096 9773 8113 9784
rect 8227 9776 8513 9784
rect 8527 9779 8713 9787
rect 9156 9776 9593 9784
rect 3247 9756 3293 9764
rect 3307 9759 3373 9767
rect 3607 9759 3653 9767
rect 3947 9759 3993 9767
rect 4456 9756 4633 9764
rect 3067 9733 3093 9741
rect 4067 9739 4193 9747
rect 4456 9744 4464 9756
rect 4647 9756 4673 9764
rect 4887 9759 5033 9767
rect 5087 9756 5493 9764
rect 6427 9756 6633 9764
rect 6727 9756 6913 9764
rect 7207 9759 7233 9767
rect 7647 9759 7733 9767
rect 7787 9759 7833 9767
rect 4696 9736 5224 9744
rect 1447 9716 1573 9724
rect 1627 9713 1653 9721
rect 2067 9713 2093 9721
rect 2327 9713 2353 9721
rect 2696 9716 3073 9724
rect 3087 9716 3153 9724
rect 3407 9716 3593 9724
rect 3887 9716 4393 9724
rect 4696 9724 4704 9736
rect 4747 9716 4813 9724
rect 5216 9724 5224 9736
rect 7496 9744 7504 9756
rect 7887 9756 8033 9764
rect 8096 9744 8104 9773
rect 9156 9770 9164 9776
rect 9607 9776 9633 9784
rect 10987 9776 11133 9784
rect 8847 9756 9013 9764
rect 9027 9759 9153 9767
rect 9267 9764 9280 9767
rect 9267 9753 9284 9764
rect 9887 9756 10073 9764
rect 10147 9756 10184 9764
rect 7427 9736 7504 9744
rect 8147 9736 8213 9744
rect 8367 9739 8873 9747
rect 4867 9716 5013 9724
rect 5227 9713 5273 9721
rect 5327 9716 5513 9724
rect 5667 9716 5853 9724
rect 7527 9713 7553 9721
rect 7687 9716 7753 9724
rect 8067 9713 8093 9721
rect 9007 9716 9033 9724
rect 9047 9716 9233 9724
rect 9276 9724 9284 9753
rect 10176 9727 10184 9756
rect 10247 9756 10293 9764
rect 10307 9759 10353 9767
rect 10567 9756 10653 9764
rect 10727 9759 10773 9767
rect 10947 9756 10964 9764
rect 10956 9744 10964 9756
rect 11287 9756 11453 9764
rect 11747 9759 11793 9767
rect 11807 9756 11953 9764
rect 12067 9756 12233 9764
rect 10956 9736 11013 9744
rect 9647 9713 9853 9721
rect 10087 9713 10113 9721
rect 10787 9716 10913 9724
rect 10927 9713 11093 9721
rect 11727 9716 11873 9724
rect 11987 9716 12073 9724
rect 12087 9716 12253 9724
rect 1267 9696 1373 9704
rect 1847 9696 2013 9704
rect 3547 9696 3673 9704
rect 3727 9696 3753 9704
rect 3767 9696 4833 9704
rect 7047 9696 7113 9704
rect 7947 9696 8153 9704
rect 8167 9696 8613 9704
rect 9587 9696 9753 9704
rect 9967 9696 10033 9704
rect 10047 9696 10153 9704
rect 10707 9696 10753 9704
rect 11407 9696 11493 9704
rect 247 9676 724 9684
rect 716 9664 724 9676
rect 1207 9676 1293 9684
rect 2407 9676 2473 9684
rect 2687 9676 2753 9684
rect 3807 9676 3913 9684
rect 3967 9676 4053 9684
rect 4647 9676 4873 9684
rect 6407 9676 6513 9684
rect 7247 9676 7873 9684
rect 10027 9676 10293 9684
rect 716 9656 1173 9664
rect 2607 9656 2784 9664
rect 2996 9660 4353 9664
rect 587 9636 753 9644
rect 1876 9636 2553 9644
rect 1876 9627 1884 9636
rect 2776 9644 2784 9656
rect 2993 9656 4353 9660
rect 2993 9647 3007 9656
rect 4407 9656 4853 9664
rect 5507 9656 5633 9664
rect 5687 9656 6713 9664
rect 6907 9656 8013 9664
rect 8507 9656 8833 9664
rect 9407 9656 9673 9664
rect 10767 9656 11153 9664
rect 11767 9656 12213 9664
rect 2776 9636 2813 9644
rect 3567 9636 3753 9644
rect 4287 9636 4793 9644
rect 5207 9636 5273 9644
rect 6827 9636 6873 9644
rect 7667 9636 7713 9644
rect 8307 9636 8773 9644
rect 10127 9636 10693 9644
rect 1187 9616 1873 9624
rect 3127 9616 3513 9624
rect 4376 9616 4513 9624
rect 4376 9607 4384 9616
rect 4927 9616 5073 9624
rect 5307 9616 5593 9624
rect 6067 9616 6153 9624
rect 6307 9616 6473 9624
rect 6627 9616 6753 9624
rect 7067 9616 7213 9624
rect 7487 9616 8193 9624
rect 8207 9616 9033 9624
rect 9047 9616 9513 9624
rect 9567 9616 9693 9624
rect 9867 9616 10273 9624
rect 10287 9616 10653 9624
rect 2367 9596 2893 9604
rect 2907 9596 3093 9604
rect 3167 9596 3293 9604
rect 3627 9596 4373 9604
rect 4807 9596 4973 9604
rect 6216 9596 7413 9604
rect 6216 9587 6224 9596
rect 7567 9596 7853 9604
rect 8867 9596 8944 9604
rect 367 9576 653 9584
rect 947 9576 993 9584
rect 1007 9576 1313 9584
rect 1387 9576 1593 9584
rect 2627 9576 2853 9584
rect 5116 9576 5293 9584
rect 1487 9556 1553 9564
rect 1567 9556 1613 9564
rect 1807 9556 1973 9564
rect 1987 9556 2093 9564
rect 3027 9556 3164 9564
rect 667 9539 693 9547
rect 747 9536 833 9544
rect 887 9539 1033 9547
rect 1167 9539 1273 9547
rect 1867 9536 1933 9544
rect 2047 9536 2173 9544
rect 2347 9536 2393 9544
rect 2487 9539 2633 9547
rect 2947 9536 3133 9544
rect 3156 9544 3164 9556
rect 4367 9556 4893 9564
rect 3156 9536 3213 9544
rect 3807 9536 3953 9544
rect 4027 9536 4233 9544
rect 196 9504 204 9533
rect 3707 9519 3733 9527
rect 4407 9516 4573 9524
rect 4827 9516 4993 9524
rect 5116 9524 5124 9576
rect 5407 9576 5573 9584
rect 5587 9576 5913 9584
rect 6087 9576 6213 9584
rect 6547 9576 6973 9584
rect 8427 9576 8593 9584
rect 8827 9576 8893 9584
rect 8936 9584 8944 9596
rect 8936 9576 9173 9584
rect 9767 9576 10073 9584
rect 10927 9576 11013 9584
rect 11547 9576 11593 9584
rect 11607 9576 11753 9584
rect 5327 9556 5353 9564
rect 5487 9556 5513 9564
rect 5527 9556 5553 9564
rect 7027 9556 7173 9564
rect 8047 9556 8213 9564
rect 8547 9556 8953 9564
rect 9267 9556 9493 9564
rect 9507 9556 9644 9564
rect 5360 9544 5373 9547
rect 5356 9533 5373 9544
rect 5927 9536 6113 9544
rect 6187 9536 6244 9544
rect 6267 9539 6313 9547
rect 6607 9539 6653 9547
rect 6707 9536 6844 9544
rect 6967 9539 6993 9547
rect 7507 9536 7673 9544
rect 5287 9519 5313 9527
rect 196 9496 213 9504
rect 287 9496 433 9504
rect 447 9496 653 9504
rect 1036 9496 1053 9504
rect 1036 9484 1044 9496
rect 1247 9493 1293 9501
rect 2167 9493 2253 9501
rect 2367 9493 2413 9501
rect 2967 9493 3013 9501
rect 3107 9493 3193 9501
rect 847 9476 1044 9484
rect 1347 9476 1373 9484
rect 1507 9476 1593 9484
rect 1607 9476 1613 9484
rect 2587 9473 3273 9481
rect 567 9456 673 9464
rect 687 9456 753 9464
rect 1847 9456 2053 9464
rect 2067 9456 2273 9464
rect 2567 9456 2913 9464
rect 3167 9456 3233 9464
rect 3436 9464 3444 9510
rect 3987 9493 4013 9501
rect 4807 9496 4873 9504
rect 5356 9487 5364 9533
rect 6236 9524 6244 9536
rect 6236 9516 6284 9524
rect 5507 9496 5733 9504
rect 5747 9493 5893 9501
rect 5967 9496 5993 9504
rect 6276 9504 6284 9516
rect 6836 9504 6844 9536
rect 7767 9536 7973 9544
rect 7987 9536 8253 9544
rect 8467 9536 8573 9544
rect 8807 9536 8973 9544
rect 9107 9536 9233 9544
rect 9367 9539 9413 9547
rect 9636 9544 9644 9556
rect 10156 9556 10853 9564
rect 9636 9536 9653 9544
rect 9667 9536 9853 9544
rect 10156 9544 10164 9556
rect 9927 9536 10164 9544
rect 10187 9538 10293 9546
rect 10307 9538 10373 9546
rect 10707 9536 10833 9544
rect 10887 9539 10953 9547
rect 11247 9539 11333 9547
rect 11507 9536 11953 9544
rect 12027 9536 12113 9544
rect 8787 9516 9253 9524
rect 9327 9516 9473 9524
rect 6276 9496 6373 9504
rect 6447 9493 6473 9501
rect 6487 9496 6773 9504
rect 7007 9496 7233 9504
rect 7327 9496 7533 9504
rect 7687 9493 7773 9501
rect 7987 9493 8013 9501
rect 8207 9493 8273 9501
rect 8567 9496 8633 9504
rect 9047 9493 9113 9501
rect 9187 9496 9373 9504
rect 9647 9493 9753 9501
rect 9867 9493 9893 9501
rect 9947 9493 10073 9501
rect 10207 9496 10513 9504
rect 10687 9493 11333 9501
rect 11427 9493 11513 9501
rect 11967 9493 11993 9501
rect 12087 9493 12293 9501
rect 4567 9476 4633 9484
rect 5267 9476 5293 9484
rect 6527 9476 6673 9484
rect 7267 9476 7653 9484
rect 8067 9476 8313 9484
rect 8327 9476 8493 9484
rect 10547 9476 10713 9484
rect 3327 9456 3444 9464
rect 3787 9456 4373 9464
rect 6547 9456 6693 9464
rect 6987 9456 7733 9464
rect 8907 9456 9433 9464
rect 9447 9456 10113 9464
rect 10827 9456 10853 9464
rect 10867 9456 10944 9464
rect 967 9436 1153 9444
rect 1167 9436 1573 9444
rect 1627 9436 2113 9444
rect 4707 9436 5273 9444
rect 5547 9436 5933 9444
rect 6207 9436 6233 9444
rect 6247 9436 6513 9444
rect 8127 9436 10253 9444
rect 10936 9444 10944 9456
rect 10936 9436 11473 9444
rect 2527 9416 3153 9424
rect 3207 9416 3313 9424
rect 3727 9416 3793 9424
rect 4427 9416 4773 9424
rect 4787 9416 4953 9424
rect 5156 9420 5293 9424
rect 5153 9416 5293 9420
rect 5153 9407 5167 9416
rect 6367 9416 6593 9424
rect 6847 9416 6873 9424
rect 8347 9416 9193 9424
rect 9247 9416 10213 9424
rect 10987 9416 11293 9424
rect 407 9396 973 9404
rect 2567 9396 2613 9404
rect 3427 9396 4213 9404
rect 4267 9396 4793 9404
rect 6727 9396 7053 9404
rect 7127 9396 7193 9404
rect 7667 9396 8753 9404
rect 9087 9396 9153 9404
rect 9167 9396 9593 9404
rect 10787 9396 10833 9404
rect 10847 9396 11453 9404
rect 3207 9376 5133 9384
rect 5267 9376 5733 9384
rect 5747 9376 5793 9384
rect 6607 9376 6973 9384
rect 7527 9376 7573 9384
rect 7587 9376 7713 9384
rect 9696 9376 9824 9384
rect 1947 9356 2213 9364
rect 3447 9356 3813 9364
rect 3887 9356 3933 9364
rect 3947 9356 4473 9364
rect 4647 9356 4873 9364
rect 4887 9356 5113 9364
rect 5187 9356 5653 9364
rect 9027 9356 9273 9364
rect 9696 9364 9704 9376
rect 9287 9356 9704 9364
rect 9816 9364 9824 9376
rect 9847 9376 9953 9384
rect 9967 9376 10493 9384
rect 10947 9376 11793 9384
rect 9816 9356 10613 9364
rect 10976 9356 11373 9364
rect 1027 9336 2613 9344
rect 2627 9336 2973 9344
rect 3087 9336 3173 9344
rect 3267 9336 3733 9344
rect 4347 9336 4493 9344
rect 4547 9336 4913 9344
rect 5147 9336 5613 9344
rect 6627 9336 6853 9344
rect 6867 9336 7133 9344
rect 8227 9336 8353 9344
rect 8367 9336 9713 9344
rect 10976 9344 10984 9356
rect 11387 9356 11413 9364
rect 11427 9356 11653 9364
rect 11667 9356 11733 9364
rect 10227 9336 10984 9344
rect 1887 9316 2053 9324
rect 3767 9316 4233 9324
rect 4247 9316 4413 9324
rect 7227 9316 7293 9324
rect 7307 9316 7513 9324
rect 8987 9316 9753 9324
rect 9807 9316 10193 9324
rect 10707 9316 10873 9324
rect 787 9296 993 9304
rect 1007 9296 1153 9304
rect 1827 9296 2193 9304
rect 4487 9296 5353 9304
rect 9287 9296 9553 9304
rect 11147 9296 11173 9304
rect 267 9276 493 9284
rect 1207 9276 1553 9284
rect 1767 9276 2413 9284
rect 2427 9276 2473 9284
rect 2867 9276 3053 9284
rect 3596 9276 3713 9284
rect 227 9256 673 9264
rect 1147 9256 2153 9264
rect 2927 9256 2993 9264
rect 3427 9256 3453 9264
rect 256 9236 293 9244
rect 256 9224 264 9236
rect 387 9239 733 9247
rect 1047 9239 1113 9247
rect 1187 9236 1273 9244
rect 1327 9239 1373 9247
rect 1647 9236 1853 9244
rect 1907 9239 2073 9247
rect 2336 9246 2453 9247
rect 2196 9224 2204 9236
rect 2347 9239 2453 9246
rect 2467 9236 2553 9244
rect 2647 9239 2653 9247
rect 2667 9239 2693 9247
rect 2747 9239 2773 9247
rect 2787 9236 3013 9244
rect 3287 9236 3364 9244
rect 196 9220 264 9224
rect 193 9216 264 9220
rect 2056 9216 2204 9224
rect 3356 9224 3364 9236
rect 3596 9230 3604 9276
rect 4507 9276 4693 9284
rect 5887 9276 6313 9284
rect 6327 9276 6393 9284
rect 6727 9276 6893 9284
rect 6907 9276 6953 9284
rect 7147 9276 7473 9284
rect 8167 9276 8253 9284
rect 8267 9276 8653 9284
rect 8747 9276 9053 9284
rect 9107 9276 10073 9284
rect 10147 9276 10673 9284
rect 10927 9276 11053 9284
rect 11067 9276 11673 9284
rect 11827 9276 12033 9284
rect 3947 9256 4393 9264
rect 5207 9256 5573 9264
rect 6127 9256 6253 9264
rect 7807 9259 8133 9267
rect 8147 9256 8393 9264
rect 10387 9256 10513 9264
rect 11007 9256 11213 9264
rect 11227 9256 11333 9264
rect 3356 9216 3413 9224
rect 193 9207 207 9216
rect 287 9193 373 9201
rect 687 9196 753 9204
rect 847 9196 1013 9204
rect 1067 9193 1093 9201
rect 1167 9196 1293 9204
rect 2056 9204 2064 9216
rect 3736 9207 3744 9253
rect 3833 9244 3847 9253
rect 3776 9240 3847 9244
rect 3773 9236 3844 9240
rect 4527 9239 4573 9247
rect 4727 9239 4753 9247
rect 4807 9236 5033 9244
rect 5047 9239 5113 9247
rect 5267 9239 5313 9247
rect 5847 9239 5913 9247
rect 6167 9239 6213 9247
rect 6327 9239 6433 9247
rect 6547 9239 6593 9247
rect 6947 9239 7053 9247
rect 8507 9239 8573 9247
rect 8707 9239 8733 9247
rect 3773 9227 3787 9236
rect 3847 9216 3933 9224
rect 1407 9196 1793 9204
rect 1807 9193 1833 9201
rect 1847 9196 2064 9204
rect 2087 9196 2133 9204
rect 2567 9193 2673 9201
rect 2727 9196 2833 9204
rect 2847 9196 2953 9204
rect 3727 9196 3744 9207
rect 3727 9193 3740 9196
rect 1487 9176 1533 9184
rect 3336 9176 3453 9184
rect 3336 9167 3344 9176
rect 4076 9184 4084 9216
rect 4207 9216 4293 9224
rect 7436 9224 7444 9236
rect 8847 9236 9213 9244
rect 9327 9239 9393 9247
rect 9527 9239 9553 9247
rect 9607 9239 9633 9247
rect 10007 9236 10053 9244
rect 10267 9239 10593 9247
rect 10607 9239 10653 9247
rect 10667 9236 10753 9244
rect 11087 9236 11113 9244
rect 11527 9239 11733 9247
rect 11747 9236 11993 9244
rect 12047 9239 12093 9247
rect 7367 9216 7444 9224
rect 7687 9216 7833 9224
rect 7967 9219 8093 9227
rect 8167 9213 8253 9221
rect 10096 9207 10104 9233
rect 12036 9224 12044 9236
rect 12167 9236 12253 9244
rect 11847 9216 12044 9224
rect 4327 9193 4373 9201
rect 4387 9193 4453 9201
rect 4587 9196 4773 9204
rect 4827 9193 4893 9201
rect 4907 9196 4993 9204
rect 5067 9196 5253 9204
rect 5867 9196 5973 9204
rect 6047 9196 6133 9204
rect 6187 9196 6313 9204
rect 6427 9196 6573 9204
rect 6667 9193 6713 9201
rect 6867 9193 6953 9201
rect 7147 9196 7193 9204
rect 7307 9193 7413 9201
rect 9047 9196 9253 9204
rect 9727 9196 10013 9204
rect 10307 9193 10353 9201
rect 10407 9193 10433 9201
rect 10907 9193 10993 9201
rect 11167 9196 11253 9204
rect 11687 9193 11753 9201
rect 12027 9196 12233 9204
rect 4076 9176 4493 9184
rect 6547 9176 6593 9184
rect 8107 9176 8473 9184
rect 10867 9176 11053 9184
rect 11067 9176 11273 9184
rect 207 9156 233 9164
rect 527 9156 833 9164
rect 1387 9156 1573 9164
rect 2067 9156 2173 9164
rect 2447 9156 2773 9164
rect 3067 9156 3252 9164
rect 3287 9156 3333 9164
rect 3887 9156 4333 9164
rect 4567 9156 4773 9164
rect 4947 9156 5373 9164
rect 5387 9156 5513 9164
rect 6087 9156 6133 9164
rect 6616 9156 7253 9164
rect 267 9136 433 9144
rect 2407 9136 2473 9144
rect 2487 9136 2633 9144
rect 3827 9136 4713 9144
rect 5127 9136 5593 9144
rect 6616 9144 6624 9156
rect 7347 9156 7544 9164
rect 6467 9136 6624 9144
rect 7536 9144 7544 9156
rect 11487 9156 11513 9164
rect 6727 9136 7244 9144
rect 7536 9136 7753 9144
rect 947 9116 1193 9124
rect 1207 9116 1253 9124
rect 1707 9116 1873 9124
rect 3927 9116 4013 9124
rect 4787 9116 5333 9124
rect 5747 9116 6313 9124
rect 6647 9116 7073 9124
rect 7236 9124 7244 9136
rect 7807 9136 8333 9144
rect 8967 9136 9053 9144
rect 10127 9136 10153 9144
rect 10647 9136 10953 9144
rect 7236 9116 7353 9124
rect 11227 9116 11633 9124
rect 1827 9096 1953 9104
rect 2247 9096 2673 9104
rect 4707 9096 4753 9104
rect 5927 9096 6373 9104
rect 6427 9096 7633 9104
rect 8227 9096 8593 9104
rect 8607 9096 8673 9104
rect 8747 9096 9093 9104
rect 9307 9096 9333 9104
rect 9587 9096 9933 9104
rect 9947 9096 10953 9104
rect 11687 9096 11713 9104
rect 807 9076 1053 9084
rect 1227 9076 1593 9084
rect 3107 9076 3473 9084
rect 3647 9076 3833 9084
rect 1247 9056 1313 9064
rect 1847 9056 2213 9064
rect 2227 9056 2293 9064
rect 2616 9056 2753 9064
rect 2616 9047 2624 9056
rect 2796 9056 2833 9064
rect 847 9036 1033 9044
rect 1367 9036 1473 9044
rect 2607 9036 2624 9047
rect 2607 9033 2620 9036
rect 2796 9031 2804 9056
rect 3887 9036 3973 9044
rect 4047 9036 4353 9044
rect 287 9019 313 9027
rect 527 9016 753 9024
rect 1007 9019 1253 9027
rect 1427 9019 1553 9027
rect 1687 9016 1893 9024
rect 1947 9019 2053 9027
rect 2187 9016 2352 9024
rect 2387 9019 2433 9027
rect 2847 9016 3013 9024
rect 3147 9016 3333 9024
rect 3527 9019 3553 9027
rect 3867 9016 3904 9024
rect 267 8973 353 8981
rect 367 8976 413 8984
rect 1027 8973 1173 8981
rect 1267 8973 1333 8981
rect 1627 8973 1673 8981
rect 2207 8976 2373 8984
rect 2627 8974 2693 8982
rect 3287 8976 3353 8984
rect 3607 8976 3713 8984
rect 3807 8973 3833 8981
rect 3896 8967 3904 9016
rect 4020 9004 4033 9007
rect 3916 8967 3924 8996
rect 4016 8993 4033 9004
rect 4016 8984 4024 8993
rect 4556 9004 4564 9093
rect 5427 9076 6173 9084
rect 8113 9084 8127 9093
rect 6927 9080 8127 9084
rect 6927 9076 8124 9080
rect 8887 9076 9713 9084
rect 9727 9076 9913 9084
rect 5527 9056 6224 9064
rect 5087 9036 5113 9044
rect 5307 9036 5573 9044
rect 6216 9044 6224 9056
rect 6247 9056 6413 9064
rect 6627 9056 6893 9064
rect 8327 9056 8593 9064
rect 8787 9056 8813 9064
rect 10527 9056 11253 9064
rect 11727 9056 11973 9064
rect 12047 9056 12273 9064
rect 6216 9036 6453 9044
rect 7627 9036 7753 9044
rect 8447 9036 8613 9044
rect 9567 9036 9633 9044
rect 9927 9036 10093 9044
rect 11487 9036 11653 9044
rect 4827 9016 5133 9024
rect 5367 9016 5473 9024
rect 5627 9016 5973 9024
rect 6456 9026 6493 9027
rect 6467 9019 6493 9026
rect 6507 9016 6713 9024
rect 6767 9016 6793 9024
rect 6807 9019 6933 9027
rect 7087 9016 7333 9024
rect 7887 9016 7913 9024
rect 8467 9019 8553 9027
rect 8667 9016 9013 9024
rect 9547 9016 9893 9024
rect 10167 9016 10393 9024
rect 10867 9019 10913 9027
rect 11200 9024 11213 9027
rect 10967 9016 11213 9024
rect 11196 9013 11213 9016
rect 11267 9019 11433 9027
rect 11767 9019 11813 9027
rect 11827 9016 11873 9024
rect 12187 9016 12233 9024
rect 3996 8976 4024 8984
rect 1307 8956 1493 8964
rect 1587 8956 1813 8964
rect 1827 8956 1873 8964
rect 1987 8956 2153 8964
rect 2927 8956 3033 8964
rect 3527 8956 3553 8964
rect 3916 8956 3932 8967
rect 3920 8953 3932 8956
rect 3996 8964 4004 8976
rect 3967 8956 4004 8964
rect 547 8936 673 8944
rect 687 8936 733 8944
rect 747 8936 833 8944
rect 1927 8936 2093 8944
rect 2307 8936 2413 8944
rect 3067 8936 3113 8944
rect 3427 8936 3773 8944
rect 3827 8936 3873 8944
rect 2027 8916 2084 8924
rect 2076 8904 2084 8916
rect 4176 8907 4184 8990
rect 4316 8967 4324 8993
rect 5027 8996 5513 9004
rect 4736 8967 4744 8993
rect 5107 8976 5133 8984
rect 5487 8973 5633 8981
rect 5747 8973 5873 8981
rect 6427 8973 6513 8981
rect 6567 8973 6613 8981
rect 6747 8976 6773 8984
rect 6867 8973 6893 8981
rect 7976 8984 7984 8996
rect 8187 8993 8313 9001
rect 8807 8999 8953 9007
rect 9227 8993 9313 9001
rect 9393 8984 9407 8993
rect 7847 8976 7984 8984
rect 8627 8973 8733 8981
rect 9393 8980 9433 8984
rect 9396 8976 9433 8980
rect 11196 8984 11204 9013
rect 9927 8973 9953 8981
rect 10027 8973 10133 8981
rect 11307 8973 11413 8981
rect 11667 8973 11733 8981
rect 11787 8973 11933 8981
rect 12007 8976 12033 8984
rect 12167 8973 12293 8981
rect 4867 8956 5293 8964
rect 5307 8956 5333 8964
rect 5487 8956 5593 8964
rect 6287 8956 6353 8964
rect 7307 8956 7333 8964
rect 5067 8936 5193 8944
rect 5476 8944 5484 8952
rect 8347 8953 8393 8961
rect 8407 8956 9373 8964
rect 11107 8956 11153 8964
rect 5447 8936 5484 8944
rect 5827 8936 6153 8944
rect 6327 8936 6533 8944
rect 6947 8936 7113 8944
rect 8707 8936 9033 8944
rect 9667 8936 9693 8944
rect 9707 8936 9833 8944
rect 10107 8936 10173 8944
rect 5447 8916 5773 8924
rect 5987 8916 8893 8924
rect 2076 8896 2473 8904
rect 4427 8896 4713 8904
rect 5287 8896 5373 8904
rect 5427 8896 5964 8904
rect 787 8876 1113 8884
rect 1127 8876 1833 8884
rect 2607 8876 2893 8884
rect 3327 8876 3793 8884
rect 3847 8876 4333 8884
rect 5956 8884 5964 8896
rect 6207 8896 6233 8904
rect 6247 8896 6753 8904
rect 7287 8896 7353 8904
rect 8327 8896 8813 8904
rect 8947 8896 9533 8904
rect 9887 8896 10573 8904
rect 5956 8876 6313 8884
rect 7467 8876 8633 8884
rect 8787 8876 8913 8884
rect 9227 8876 9433 8884
rect 9567 8876 9653 8884
rect 9767 8876 10853 8884
rect 2027 8856 2933 8864
rect 2947 8856 3193 8864
rect 3847 8856 4013 8864
rect 5387 8856 5453 8864
rect 6527 8856 6813 8864
rect 8807 8856 9193 8864
rect 9216 8856 9813 8864
rect 707 8836 773 8844
rect 2887 8836 3593 8844
rect 4627 8836 5433 8844
rect 6387 8836 6473 8844
rect 6487 8836 7153 8844
rect 9216 8844 9224 8856
rect 11267 8856 11553 8864
rect 11567 8856 12013 8864
rect 8867 8836 9224 8844
rect 3187 8816 3533 8824
rect 4167 8816 4313 8824
rect 4607 8816 4913 8824
rect 5827 8816 6053 8824
rect 8647 8816 9513 8824
rect 9527 8816 9593 8824
rect 9647 8816 10673 8824
rect 10767 8816 11753 8824
rect 267 8796 493 8804
rect 607 8796 813 8804
rect 827 8796 993 8804
rect 1947 8796 2333 8804
rect 3807 8796 5053 8804
rect 5267 8796 5473 8804
rect 7047 8796 7673 8804
rect 8367 8796 8533 8804
rect 8547 8796 8932 8804
rect 8967 8796 9933 8804
rect 10827 8796 11233 8804
rect 2367 8776 2633 8784
rect 2647 8776 2733 8784
rect 3167 8776 3613 8784
rect 4187 8776 5013 8784
rect 5207 8776 5413 8784
rect 6327 8776 6413 8784
rect 6667 8776 7713 8784
rect 8767 8776 8873 8784
rect 10167 8776 11593 8784
rect 227 8756 433 8764
rect 1307 8756 1533 8764
rect 1547 8756 1573 8764
rect 2307 8756 2833 8764
rect 3947 8756 4033 8764
rect 4047 8756 4513 8764
rect 4667 8756 4873 8764
rect 5527 8756 5833 8764
rect 6047 8756 6113 8764
rect 6607 8756 6813 8764
rect 6867 8756 7413 8764
rect 7867 8756 8213 8764
rect 8227 8756 8453 8764
rect 8527 8756 8593 8764
rect 8907 8756 9253 8764
rect 9267 8756 9473 8764
rect 10567 8756 10653 8764
rect 10887 8756 10933 8764
rect 367 8736 493 8744
rect 507 8736 733 8744
rect 4927 8736 5353 8744
rect 5367 8736 5493 8744
rect 5547 8736 5813 8744
rect 5856 8736 6013 8744
rect 1067 8716 1113 8724
rect 1347 8719 1373 8727
rect 1627 8716 1853 8724
rect 2987 8718 3133 8726
rect 3387 8718 3433 8726
rect 3487 8719 3573 8727
rect 4167 8719 4253 8727
rect 4307 8719 4333 8727
rect 4567 8716 4693 8724
rect 3996 8704 4004 8716
rect 4707 8716 4793 8724
rect 4807 8719 4853 8727
rect 5087 8719 5153 8727
rect 5227 8716 5313 8724
rect 5856 8724 5864 8736
rect 6207 8736 6333 8744
rect 11587 8736 11793 8744
rect 5816 8720 5864 8724
rect 5373 8707 5387 8713
rect 5813 8716 5864 8720
rect 3996 8696 4913 8704
rect 5373 8700 5393 8707
rect 5376 8696 5393 8700
rect 5380 8693 5393 8696
rect 5813 8707 5827 8716
rect 6013 8724 6027 8733
rect 6013 8720 6073 8724
rect 6016 8716 6073 8720
rect 6367 8719 6473 8727
rect 6747 8719 6853 8727
rect 6987 8719 7113 8727
rect 7307 8716 7373 8724
rect 7387 8719 7453 8727
rect 7467 8716 7613 8724
rect 447 8676 513 8684
rect 687 8673 753 8681
rect 1007 8673 1073 8681
rect 1387 8676 1593 8684
rect 1747 8676 1833 8684
rect 2547 8676 2913 8684
rect 3236 8683 3453 8684
rect 3247 8676 3453 8683
rect 3767 8676 4013 8684
rect 4347 8676 4533 8684
rect 5107 8676 5333 8684
rect 5547 8684 5560 8687
rect 5547 8673 5564 8684
rect 1647 8656 2033 8664
rect 2047 8656 2073 8664
rect 2407 8656 2513 8664
rect 2947 8656 3053 8664
rect 4247 8656 4693 8664
rect 4947 8656 5513 8664
rect 347 8636 753 8644
rect 2827 8636 2913 8644
rect 3567 8636 3953 8644
rect 4207 8636 4273 8644
rect 4967 8636 5213 8644
rect 5287 8636 5413 8644
rect 5556 8644 5564 8673
rect 5536 8636 5564 8644
rect 307 8616 793 8624
rect 927 8616 1033 8624
rect 1047 8616 1613 8624
rect 1667 8616 2193 8624
rect 2727 8616 3193 8624
rect 3907 8616 4173 8624
rect 4547 8616 4733 8624
rect 5536 8624 5544 8636
rect 5447 8616 5544 8624
rect 5676 8607 5684 8696
rect 5996 8687 6004 8713
rect 6267 8676 6432 8684
rect 6467 8676 6553 8684
rect 6896 8684 6904 8713
rect 8016 8704 8024 8716
rect 8067 8716 8253 8724
rect 8267 8716 8773 8724
rect 9067 8716 9113 8724
rect 9347 8716 9593 8724
rect 9607 8716 9773 8724
rect 10027 8719 10113 8727
rect 10347 8716 10373 8724
rect 10507 8719 10613 8727
rect 10627 8716 10913 8724
rect 10967 8719 11013 8727
rect 11167 8719 11233 8727
rect 11247 8716 11313 8724
rect 11367 8719 11493 8727
rect 12067 8719 12113 8727
rect 8016 8696 8704 8704
rect 6767 8673 6833 8681
rect 6887 8676 6904 8684
rect 7447 8673 7493 8681
rect 7627 8673 7653 8681
rect 7707 8676 7753 8684
rect 7887 8673 7993 8681
rect 8287 8676 8433 8684
rect 8567 8676 8593 8684
rect 8696 8684 8704 8696
rect 11536 8704 11544 8716
rect 12227 8716 12293 8724
rect 11347 8696 11544 8704
rect 11816 8696 11913 8704
rect 8707 8673 8753 8681
rect 9187 8673 9553 8681
rect 9767 8673 9813 8681
rect 11816 8684 11824 8696
rect 9947 8676 10133 8684
rect 10527 8673 10593 8681
rect 10687 8673 10733 8681
rect 11387 8673 11513 8681
rect 11947 8676 12033 8684
rect 12127 8673 12273 8681
rect 5967 8656 6013 8664
rect 6187 8656 6233 8664
rect 6967 8656 7173 8664
rect 9127 8656 9233 8664
rect 9247 8656 9353 8664
rect 10987 8656 11213 8664
rect 6956 8644 6964 8653
rect 6387 8636 6964 8644
rect 8667 8636 8793 8644
rect 9227 8636 9313 8644
rect 9967 8636 10153 8644
rect 10287 8636 10393 8644
rect 11267 8636 11373 8644
rect 5887 8624 5900 8627
rect 5887 8613 5904 8624
rect 5967 8616 6333 8624
rect 7767 8616 8613 8624
rect 8947 8616 9073 8624
rect 9087 8616 9173 8624
rect 9336 8616 9853 8624
rect 5896 8607 5904 8613
rect 867 8596 2273 8604
rect 2287 8596 2373 8604
rect 2387 8596 3373 8604
rect 3927 8596 4153 8604
rect 4487 8596 4953 8604
rect 5807 8596 5873 8604
rect 5896 8596 5913 8607
rect 5900 8593 5913 8596
rect 6047 8596 6133 8604
rect 6727 8596 6873 8604
rect 6887 8596 7293 8604
rect 7907 8596 7953 8604
rect 9336 8604 9344 8616
rect 12147 8616 12333 8624
rect 9067 8596 9344 8604
rect 9587 8596 10473 8604
rect 10667 8596 11293 8604
rect 11647 8596 11933 8604
rect 1087 8576 1153 8584
rect 1167 8576 1773 8584
rect 2396 8576 3033 8584
rect 287 8556 353 8564
rect 2396 8564 2404 8576
rect 3427 8576 3513 8584
rect 3527 8576 4412 8584
rect 4447 8576 4733 8584
rect 5707 8576 5813 8584
rect 6247 8576 7133 8584
rect 7447 8576 7873 8584
rect 8207 8576 8513 8584
rect 8676 8576 8933 8584
rect 1767 8556 2404 8564
rect 3387 8556 6633 8564
rect 7107 8556 7393 8564
rect 7587 8556 7844 8564
rect 807 8536 1313 8544
rect 1627 8536 1693 8544
rect 2287 8536 2533 8544
rect 2847 8536 3413 8544
rect 4027 8536 4633 8544
rect 5247 8536 5473 8544
rect 5807 8536 6153 8544
rect 6167 8536 6373 8544
rect 7087 8536 7653 8544
rect 7667 8536 7793 8544
rect 7836 8544 7844 8556
rect 8676 8564 8684 8576
rect 8627 8556 8684 8564
rect 8787 8556 9513 8564
rect 9527 8556 9973 8564
rect 10547 8556 10633 8564
rect 10727 8556 10933 8564
rect 11007 8556 11133 8564
rect 11687 8556 11813 8564
rect 7836 8536 8233 8544
rect 8527 8536 9233 8544
rect 10487 8536 11153 8544
rect 3047 8516 3353 8524
rect 3527 8516 3713 8524
rect 3967 8513 3973 8527
rect 5227 8516 5733 8524
rect 5947 8516 6144 8524
rect 247 8496 313 8504
rect 327 8496 433 8504
rect 487 8496 973 8504
rect 1127 8499 1293 8507
rect 1347 8496 1473 8504
rect 1527 8499 1653 8507
rect 1867 8499 1893 8507
rect 2107 8499 2173 8507
rect 2247 8496 2433 8504
rect 2733 8504 2747 8513
rect 2547 8496 2753 8504
rect 3027 8496 3473 8504
rect 3487 8496 3813 8504
rect 4427 8496 4653 8504
rect 4756 8496 4793 8504
rect 3196 8476 3213 8484
rect 227 8456 293 8464
rect 347 8453 453 8461
rect 707 8453 733 8461
rect 1107 8453 1173 8461
rect 1687 8453 1773 8461
rect 3196 8464 3204 8476
rect 4227 8473 4433 8481
rect 2127 8456 2193 8464
rect 2387 8453 2413 8461
rect 2667 8453 2693 8461
rect 2747 8456 3204 8464
rect 3727 8456 3913 8464
rect 4756 8464 4764 8496
rect 5007 8499 5193 8507
rect 5236 8496 5253 8504
rect 5496 8496 5553 8504
rect 5847 8496 6053 8504
rect 5236 8484 5244 8496
rect 5216 8476 5244 8484
rect 5216 8464 5224 8476
rect 5496 8467 5504 8496
rect 6136 8504 6144 8516
rect 6987 8516 7433 8524
rect 7627 8516 7853 8524
rect 8567 8516 8813 8524
rect 10047 8516 10313 8524
rect 10327 8516 10453 8524
rect 11467 8516 11653 8524
rect 6136 8496 6153 8504
rect 6347 8496 6393 8504
rect 6407 8496 6953 8504
rect 7187 8496 7313 8504
rect 7387 8496 7453 8504
rect 8947 8499 8973 8507
rect 9027 8496 9173 8504
rect 7496 8467 7504 8496
rect 9327 8496 9493 8504
rect 9687 8496 9773 8504
rect 10087 8496 10133 8504
rect 10627 8496 10753 8504
rect 10887 8496 11073 8504
rect 11187 8496 11273 8504
rect 11367 8499 11413 8507
rect 11487 8496 11533 8504
rect 11727 8496 11793 8504
rect 11847 8499 11993 8507
rect 12087 8498 12213 8506
rect 12233 8504 12247 8513
rect 12233 8500 12264 8504
rect 12236 8496 12264 8500
rect 7607 8476 7793 8484
rect 7807 8479 7913 8487
rect 8067 8473 8193 8481
rect 4907 8456 5224 8464
rect 5767 8453 5813 8461
rect 6067 8453 6093 8461
rect 6147 8453 6253 8461
rect 6387 8456 6453 8464
rect 6607 8453 6713 8461
rect 7327 8453 7433 8461
rect 7496 8456 7513 8467
rect 7500 8453 7513 8456
rect 8387 8453 8493 8461
rect 8687 8456 8733 8464
rect 8747 8456 8993 8464
rect 9267 8453 9293 8461
rect 9347 8453 9473 8461
rect 9827 8456 10013 8464
rect 12256 8464 12264 8496
rect 10767 8453 11153 8461
rect 11327 8453 11393 8461
rect 11447 8456 11953 8464
rect 12027 8453 12053 8461
rect 12247 8456 12264 8464
rect 507 8436 653 8444
rect 787 8436 1053 8444
rect 1647 8436 1913 8444
rect 2567 8433 3053 8441
rect 3367 8436 3393 8444
rect 4667 8436 4813 8444
rect 5247 8436 5533 8444
rect 5547 8436 5773 8444
rect 5867 8436 5913 8444
rect 5927 8436 6053 8444
rect 6156 8436 6233 8444
rect 807 8416 853 8424
rect 1007 8416 1253 8424
rect 1967 8416 2233 8424
rect 2576 8416 2893 8424
rect 987 8396 1313 8404
rect 2576 8404 2584 8416
rect 3587 8416 3753 8424
rect 4487 8416 4573 8424
rect 4727 8416 4913 8424
rect 5287 8416 5504 8424
rect 2467 8396 2584 8404
rect 2927 8396 3033 8404
rect 4067 8396 4373 8404
rect 4387 8396 4933 8404
rect 5496 8404 5504 8416
rect 6156 8424 6164 8436
rect 6367 8436 6473 8444
rect 7187 8436 7233 8444
rect 7507 8436 7533 8444
rect 7927 8436 8253 8444
rect 9567 8436 9633 8444
rect 10107 8436 10153 8444
rect 10167 8436 10633 8444
rect 10907 8436 10993 8444
rect 11167 8436 11693 8444
rect 11747 8436 11773 8444
rect 5587 8416 6164 8424
rect 6547 8416 7093 8424
rect 7487 8416 7553 8424
rect 8827 8416 9053 8424
rect 11287 8416 12073 8424
rect 5496 8396 5953 8404
rect 6067 8396 6213 8404
rect 7167 8396 7193 8404
rect 7467 8396 7893 8404
rect 8187 8396 8333 8404
rect 10067 8396 10493 8404
rect 10507 8396 10673 8404
rect 10687 8396 11333 8404
rect 1367 8376 1753 8384
rect 1907 8376 2444 8384
rect 2436 8367 2444 8376
rect 2947 8376 2993 8384
rect 4647 8376 5473 8384
rect 5627 8376 7033 8384
rect 7167 8376 7213 8384
rect 7227 8376 7513 8384
rect 8227 8376 8273 8384
rect 10107 8376 10133 8384
rect 767 8356 953 8364
rect 2447 8356 2533 8364
rect 4807 8356 5153 8364
rect 5367 8356 5593 8364
rect 5687 8356 5993 8364
rect 6387 8356 6633 8364
rect 6647 8356 6733 8364
rect 6807 8356 7593 8364
rect 8427 8356 8653 8364
rect 9007 8356 9553 8364
rect 9887 8356 10473 8364
rect 11667 8356 12313 8364
rect 1247 8336 1793 8344
rect 1807 8336 2093 8344
rect 2267 8336 2453 8344
rect 2887 8336 3113 8344
rect 4367 8336 4533 8344
rect 5147 8336 6313 8344
rect 7067 8336 7393 8344
rect 7467 8336 7613 8344
rect 8287 8336 8673 8344
rect 9067 8336 10993 8344
rect 607 8316 633 8324
rect 647 8316 1152 8324
rect 1187 8316 1833 8324
rect 2367 8316 2553 8324
rect 2907 8316 3013 8324
rect 5587 8316 5693 8324
rect 5787 8316 6133 8324
rect 6187 8316 6893 8324
rect 8207 8316 8393 8324
rect 8667 8316 9033 8324
rect 10467 8316 10873 8324
rect 2047 8296 2524 8304
rect 467 8276 1973 8284
rect 2407 8276 2493 8284
rect 2516 8284 2524 8296
rect 3187 8296 3593 8304
rect 3607 8296 3913 8304
rect 4587 8296 5053 8304
rect 5327 8296 5413 8304
rect 5507 8296 5553 8304
rect 5727 8296 6333 8304
rect 8196 8304 8204 8313
rect 8047 8296 8204 8304
rect 9507 8296 9833 8304
rect 2516 8276 2833 8284
rect 4167 8276 4553 8284
rect 5107 8276 6064 8284
rect 3147 8256 3553 8264
rect 4007 8256 4033 8264
rect 4087 8256 4573 8264
rect 5067 8256 5293 8264
rect 5587 8256 5773 8264
rect 6056 8264 6064 8276
rect 6147 8276 6293 8284
rect 6307 8276 6973 8284
rect 9387 8276 9453 8284
rect 9496 8276 9613 8284
rect 6056 8256 6513 8264
rect 6667 8256 6773 8264
rect 7027 8256 7113 8264
rect 7267 8256 7573 8264
rect 7727 8256 8373 8264
rect 9496 8264 9504 8276
rect 9627 8276 9673 8284
rect 9687 8276 9733 8284
rect 9107 8256 9504 8264
rect 11107 8256 11353 8264
rect 11367 8256 11413 8264
rect 247 8236 553 8244
rect 847 8236 1253 8244
rect 1987 8236 2193 8244
rect 2527 8236 2553 8244
rect 4187 8236 4733 8244
rect 4787 8236 5093 8244
rect 5447 8236 5793 8244
rect 8296 8236 8353 8244
rect 2867 8216 2973 8224
rect 3487 8216 3693 8224
rect 5467 8216 5493 8224
rect 5507 8216 5573 8224
rect 5947 8216 6193 8224
rect 7007 8216 7073 8224
rect 7667 8216 8173 8224
rect 287 8199 313 8207
rect 267 8156 393 8164
rect 516 8147 524 8196
rect 727 8196 793 8204
rect 967 8196 1093 8204
rect 1147 8198 1193 8206
rect 1267 8199 1333 8207
rect 1447 8196 1533 8204
rect 1547 8199 1613 8207
rect 1947 8199 2073 8207
rect 2127 8199 2153 8207
rect 2413 8204 2427 8213
rect 2413 8200 2473 8204
rect 2416 8196 2473 8200
rect 3227 8199 3432 8207
rect 3707 8196 3933 8204
rect 1656 8184 1664 8196
rect 1507 8176 1664 8184
rect 1736 8176 1853 8184
rect 547 8153 873 8161
rect 887 8153 913 8161
rect 1736 8164 1744 8176
rect 2387 8176 2552 8184
rect 2587 8179 2673 8187
rect 3456 8184 3464 8196
rect 4047 8196 4253 8204
rect 4267 8198 4373 8206
rect 4387 8196 4553 8204
rect 4607 8199 4653 8207
rect 4887 8199 4993 8207
rect 5047 8199 5093 8207
rect 6227 8196 6473 8204
rect 6527 8196 6733 8204
rect 6747 8196 6893 8204
rect 7307 8196 7553 8204
rect 3236 8176 3464 8184
rect 1027 8156 1073 8164
rect 1647 8156 1744 8164
rect 1767 8156 1913 8164
rect 2927 8156 3033 8164
rect 3236 8164 3244 8176
rect 3627 8163 3804 8164
rect 4036 8163 4173 8164
rect 3627 8156 3793 8163
rect 3807 8152 4033 8160
rect 4047 8156 4173 8163
rect 4287 8156 4473 8164
rect 4547 8156 4773 8164
rect 4867 8156 5033 8164
rect 5396 8164 5404 8193
rect 7887 8179 7973 8187
rect 8027 8176 8073 8184
rect 8087 8176 8113 8184
rect 8296 8184 8304 8236
rect 9567 8236 9653 8244
rect 9947 8236 9993 8244
rect 10447 8236 10553 8244
rect 10567 8236 10913 8244
rect 11387 8236 12213 8244
rect 8416 8213 8417 8224
rect 8707 8216 8793 8224
rect 8327 8200 8384 8204
rect 8327 8196 8387 8200
rect 8373 8187 8387 8196
rect 8296 8176 8344 8184
rect 5396 8156 5473 8164
rect 5687 8153 5713 8161
rect 5847 8153 5953 8161
rect 6207 8153 6313 8161
rect 6327 8153 6793 8161
rect 7027 8156 7153 8164
rect 7167 8156 7233 8164
rect 7607 8156 7673 8164
rect 8336 8164 8344 8176
rect 8416 8184 8424 8213
rect 8816 8196 8973 8204
rect 8987 8199 9053 8207
rect 9227 8199 9333 8207
rect 8416 8176 8433 8184
rect 8007 8156 8293 8164
rect 587 8136 773 8144
rect 1367 8136 1573 8144
rect 2847 8136 2873 8144
rect 4607 8136 4653 8144
rect 4927 8136 5092 8144
rect 5127 8136 5284 8144
rect 1267 8116 1673 8124
rect 2127 8116 2453 8124
rect 3487 8116 3633 8124
rect 3707 8116 4153 8124
rect 4287 8116 4493 8124
rect 5276 8124 5284 8136
rect 5447 8136 6153 8144
rect 6247 8136 6293 8144
rect 7547 8136 7713 8144
rect 8556 8144 8564 8176
rect 8727 8176 8792 8184
rect 8816 8184 8824 8196
rect 9547 8196 9653 8204
rect 9667 8196 9793 8204
rect 8836 8180 9153 8184
rect 8833 8176 9153 8180
rect 8833 8167 8847 8176
rect 9867 8173 10053 8181
rect 10416 8187 10424 8216
rect 11067 8216 11153 8224
rect 11207 8216 11273 8224
rect 11287 8216 11293 8224
rect 11167 8199 11593 8207
rect 10256 8164 10264 8176
rect 10407 8176 10424 8187
rect 10956 8184 10964 8196
rect 11667 8196 11713 8204
rect 11967 8196 12073 8204
rect 12187 8196 12293 8204
rect 10956 8176 11273 8184
rect 10407 8173 10420 8176
rect 8856 8156 9393 8164
rect 8556 8136 8753 8144
rect 8856 8144 8864 8156
rect 9407 8153 9493 8161
rect 10256 8156 10533 8164
rect 11127 8156 11173 8164
rect 11447 8156 11673 8164
rect 12087 8153 12233 8161
rect 8827 8136 8864 8144
rect 8967 8136 9113 8144
rect 9127 8136 9233 8144
rect 9247 8136 9593 8144
rect 9907 8136 9993 8144
rect 5276 8116 5373 8124
rect 6767 8116 6964 8124
rect 327 8096 813 8104
rect 2187 8096 2553 8104
rect 4327 8096 4433 8104
rect 4587 8096 4793 8104
rect 5247 8096 5373 8104
rect 5607 8096 6113 8104
rect 6956 8104 6964 8116
rect 8447 8116 8713 8124
rect 9087 8116 9213 8124
rect 9647 8116 9773 8124
rect 10947 8116 11093 8124
rect 11276 8116 11833 8124
rect 6956 8096 7613 8104
rect 8116 8096 8253 8104
rect 2027 8076 2153 8084
rect 2227 8076 2312 8084
rect 2347 8076 2453 8084
rect 3467 8076 3533 8084
rect 3607 8076 3953 8084
rect 4227 8076 4533 8084
rect 5207 8076 5533 8084
rect 6527 8076 6853 8084
rect 8116 8084 8124 8096
rect 8767 8096 9133 8104
rect 9267 8096 9353 8104
rect 9967 8096 10093 8104
rect 11276 8104 11284 8116
rect 11847 8116 11933 8124
rect 10907 8096 11284 8104
rect 11687 8096 12193 8104
rect 6907 8076 8124 8084
rect 8187 8076 8493 8084
rect 8667 8076 9193 8084
rect 10307 8076 10473 8084
rect 3067 8056 3193 8064
rect 4587 8056 4653 8064
rect 5327 8056 5573 8064
rect 5767 8056 6093 8064
rect 6107 8056 6353 8064
rect 7467 8056 7553 8064
rect 9887 8056 9913 8064
rect 11287 8056 11513 8064
rect 1987 8036 2293 8044
rect 2427 8036 2933 8044
rect 2947 8036 3633 8044
rect 3647 8036 3673 8044
rect 3907 8036 4033 8044
rect 4247 8036 4493 8044
rect 5153 8044 5167 8053
rect 5007 8036 5553 8044
rect 5607 8036 5673 8044
rect 6707 8036 7073 8044
rect 7227 8036 7373 8044
rect 8147 8036 8413 8044
rect 8647 8036 8733 8044
rect 8747 8036 9113 8044
rect 10093 8044 10107 8053
rect 10093 8040 10313 8044
rect 10096 8036 10313 8040
rect 287 8016 313 8024
rect 1487 8016 1673 8024
rect 2367 8016 2433 8024
rect 2787 8016 2833 8024
rect 3187 8016 3333 8024
rect 5256 8016 5433 8024
rect 1067 7996 1393 8004
rect 1407 7996 1453 8004
rect 2027 7996 2173 8004
rect 2347 7996 2473 8004
rect 4007 7996 4153 8004
rect 4167 7996 4393 8004
rect 5256 8004 5264 8016
rect 6007 8016 6473 8024
rect 6887 8016 7153 8024
rect 7167 8016 7533 8024
rect 7547 8016 7633 8024
rect 8247 8016 8713 8024
rect 9587 8016 9713 8024
rect 10547 8016 10713 8024
rect 11547 8016 11593 8024
rect 11807 8016 12013 8024
rect 4507 7996 5264 8004
rect 5276 7996 5593 8004
rect 787 7979 913 7987
rect 1127 7976 1213 7984
rect 1227 7979 1293 7987
rect 1527 7979 1573 7987
rect 2256 7986 2293 7987
rect 2267 7979 2293 7986
rect 3167 7979 3293 7987
rect 3547 7979 3633 7987
rect 3927 7979 3973 7987
rect 5276 7984 5284 7996
rect 5867 7996 5913 8004
rect 8767 7996 8993 8004
rect 9847 7996 10433 8004
rect 10447 7996 10893 8004
rect 5256 7976 5284 7984
rect 1687 7953 1813 7961
rect 2087 7959 2133 7967
rect 2207 7956 2393 7964
rect 267 7936 493 7944
rect 507 7936 753 7944
rect 1327 7936 1413 7944
rect 1507 7936 1553 7944
rect 2247 7933 2353 7941
rect 827 7916 953 7924
rect 967 7916 1013 7924
rect 1027 7916 1484 7924
rect 327 7896 533 7904
rect 1476 7904 1484 7916
rect 1667 7916 2033 7924
rect 2436 7924 2444 7953
rect 2487 7953 2573 7961
rect 2847 7959 2873 7967
rect 3087 7936 3173 7944
rect 4196 7944 4204 7973
rect 3907 7933 3953 7941
rect 4187 7936 4204 7944
rect 4347 7936 4453 7944
rect 4516 7927 4524 7956
rect 2047 7916 2413 7924
rect 2427 7916 2444 7924
rect 3627 7916 3713 7924
rect 4367 7916 4433 7924
rect 4507 7916 4524 7927
rect 4507 7913 4520 7916
rect 4596 7924 4604 7953
rect 5256 7964 5264 7976
rect 5636 7964 5644 7976
rect 5767 7976 5933 7984
rect 6227 7976 6413 7984
rect 4567 7916 4604 7924
rect 1476 7896 1613 7904
rect 3327 7896 3853 7904
rect 4187 7896 4233 7904
rect 227 7876 673 7884
rect 687 7876 1053 7884
rect 2227 7876 2793 7884
rect 4127 7876 4413 7884
rect 4776 7867 4784 7950
rect 4956 7924 4964 7953
rect 4996 7927 5004 7956
rect 5636 7956 6004 7964
rect 5996 7944 6004 7956
rect 6496 7944 6504 7993
rect 6667 7979 6733 7987
rect 6987 7976 7033 7984
rect 7147 7976 7273 7984
rect 7707 7976 7733 7984
rect 8347 7978 8373 7986
rect 8607 7979 8673 7987
rect 9027 7976 9053 7984
rect 9167 7976 9304 7984
rect 9607 7979 9693 7987
rect 10607 7979 10733 7987
rect 7807 7959 7833 7967
rect 8007 7953 8133 7961
rect 8187 7956 8273 7964
rect 9036 7956 9053 7964
rect 9296 7964 9304 7976
rect 10927 7976 11013 7984
rect 11207 7976 11233 7984
rect 11467 7976 11493 7984
rect 11687 7979 11733 7987
rect 11787 7976 12053 7984
rect 9296 7956 9313 7964
rect 5587 7933 5653 7941
rect 5707 7933 5753 7941
rect 5967 7933 5993 7941
rect 6127 7933 6193 7941
rect 7067 7933 7213 7941
rect 7267 7933 7293 7941
rect 7447 7936 7593 7944
rect 8747 7933 8873 7941
rect 8947 7936 8993 7944
rect 9036 7927 9044 7956
rect 9833 7944 9847 7953
rect 9887 7953 10053 7961
rect 10187 7956 10253 7964
rect 10527 7956 10573 7964
rect 11256 7956 11573 7964
rect 11256 7944 11264 7956
rect 9527 7933 9713 7941
rect 9796 7940 9847 7944
rect 9796 7936 9844 7940
rect 9796 7927 9804 7936
rect 10887 7933 10953 7941
rect 11307 7933 11333 7941
rect 11527 7936 11673 7944
rect 4947 7916 4964 7924
rect 4987 7924 5004 7927
rect 4987 7916 5453 7924
rect 4987 7913 5000 7916
rect 5507 7916 5733 7924
rect 5747 7916 6233 7924
rect 6447 7916 6653 7924
rect 8167 7916 8193 7924
rect 8407 7916 8693 7924
rect 9787 7916 9804 7927
rect 9787 7913 9800 7916
rect 5387 7896 5413 7904
rect 5567 7896 6293 7904
rect 6427 7896 7013 7904
rect 7067 7896 7193 7904
rect 7447 7896 7493 7904
rect 7687 7896 8333 7904
rect 10227 7896 10393 7904
rect 11667 7896 11753 7904
rect 5107 7876 5453 7884
rect 5567 7876 6753 7884
rect 8507 7876 8772 7884
rect 8807 7876 9113 7884
rect 10627 7876 11193 7884
rect 4767 7856 4784 7867
rect 4767 7853 4780 7856
rect 5447 7856 5533 7864
rect 5607 7856 5913 7864
rect 6867 7856 9533 7864
rect 11007 7856 11313 7864
rect 3767 7836 3913 7844
rect 4807 7836 5064 7844
rect 667 7816 1793 7824
rect 1807 7816 2153 7824
rect 2167 7816 2313 7824
rect 2667 7816 2993 7824
rect 3767 7816 4113 7824
rect 4627 7816 4713 7824
rect 5056 7824 5064 7836
rect 6247 7836 6673 7844
rect 6967 7836 7493 7844
rect 7567 7836 7833 7844
rect 7967 7836 8233 7844
rect 8407 7836 8433 7844
rect 8447 7836 8853 7844
rect 9107 7836 9553 7844
rect 9887 7836 10453 7844
rect 5056 7816 5553 7824
rect 5767 7816 6013 7824
rect 6127 7816 6693 7824
rect 7587 7816 8153 7824
rect 2447 7796 2913 7804
rect 3407 7796 4613 7804
rect 4787 7796 5033 7804
rect 6407 7796 6453 7804
rect 8236 7796 8593 7804
rect 8236 7787 8244 7796
rect 8607 7796 8993 7804
rect 9187 7796 9573 7804
rect 9727 7796 10633 7804
rect 10647 7796 10693 7804
rect 1067 7776 1433 7784
rect 3027 7776 3933 7784
rect 4847 7773 4853 7787
rect 5096 7776 5773 7784
rect 547 7756 1993 7764
rect 2567 7756 2973 7764
rect 3647 7756 4073 7764
rect 4767 7756 4913 7764
rect 5096 7764 5104 7776
rect 6207 7776 6813 7784
rect 7507 7776 8233 7784
rect 8487 7776 8953 7784
rect 11187 7776 11793 7784
rect 5067 7756 5104 7764
rect 6707 7756 7093 7764
rect 9607 7756 10533 7764
rect 11207 7756 11513 7764
rect 12087 7756 12233 7764
rect 587 7736 633 7744
rect 1907 7736 3513 7744
rect 3587 7736 3853 7744
rect 3867 7736 4113 7744
rect 4127 7736 4493 7744
rect 4827 7736 4973 7744
rect 5047 7736 5393 7744
rect 5547 7736 5713 7744
rect 5787 7736 6633 7744
rect 7427 7736 7553 7744
rect 8227 7736 8433 7744
rect 8587 7736 8693 7744
rect 8707 7736 9293 7744
rect 10347 7736 10513 7744
rect 267 7716 533 7724
rect 1107 7716 1353 7724
rect 1607 7716 1733 7724
rect 1747 7716 2613 7724
rect 3327 7716 3793 7724
rect 6687 7716 7033 7724
rect 7607 7716 7704 7724
rect 4947 7696 5073 7704
rect 5087 7699 5372 7707
rect 5407 7696 5553 7704
rect 5867 7696 5913 7704
rect 7647 7696 7673 7704
rect 187 7679 213 7687
rect 427 7679 493 7687
rect 587 7676 613 7684
rect 667 7676 713 7684
rect 727 7679 793 7687
rect 1047 7676 1153 7684
rect 1167 7676 1313 7684
rect 1327 7679 1653 7687
rect 1847 7676 2053 7684
rect 2707 7679 2773 7687
rect 2947 7676 3013 7684
rect 776 7656 933 7664
rect 776 7644 784 7656
rect 2316 7664 2324 7675
rect 3307 7678 3333 7686
rect 3827 7679 3893 7687
rect 4087 7676 4353 7684
rect 4367 7676 4413 7684
rect 5627 7679 5733 7687
rect 5747 7676 5833 7684
rect 5847 7676 5953 7684
rect 6027 7676 6193 7684
rect 6507 7679 6713 7687
rect 6907 7679 6933 7687
rect 7047 7676 7213 7684
rect 7287 7679 7313 7687
rect 7696 7684 7704 7716
rect 7987 7716 8133 7724
rect 9487 7716 9753 7724
rect 9767 7716 10213 7724
rect 11587 7716 11873 7724
rect 11887 7716 11913 7724
rect 12227 7716 12333 7724
rect 7856 7696 7953 7704
rect 7856 7684 7864 7696
rect 10387 7696 10813 7704
rect 10927 7696 10973 7704
rect 11707 7696 11793 7704
rect 7636 7676 7704 7684
rect 7836 7676 7864 7684
rect 2136 7656 2873 7664
rect 287 7633 333 7641
rect 567 7633 593 7641
rect 607 7636 784 7644
rect 2136 7644 2144 7656
rect 3556 7656 3613 7664
rect 1047 7636 1073 7644
rect 1127 7633 1153 7641
rect 1867 7633 1893 7641
rect 2127 7636 2144 7644
rect 2687 7636 2953 7644
rect 3067 7633 3113 7640
rect 3127 7633 3193 7640
rect 3067 7632 3193 7633
rect 3556 7644 3564 7656
rect 4636 7656 4773 7664
rect 4636 7644 4644 7656
rect 4987 7656 5013 7664
rect 5027 7653 5053 7661
rect 5227 7656 5284 7664
rect 3347 7636 3513 7644
rect 4427 7633 4633 7641
rect 5276 7644 5284 7656
rect 5347 7656 5413 7664
rect 7636 7664 7644 7676
rect 7627 7656 7804 7664
rect 7836 7664 7844 7676
rect 8087 7676 8193 7684
rect 8207 7676 8553 7684
rect 8687 7679 8733 7687
rect 9047 7676 9133 7684
rect 9307 7676 9553 7684
rect 9567 7676 9673 7684
rect 9847 7676 10073 7684
rect 7827 7656 7844 7664
rect 4827 7636 4873 7644
rect 5276 7636 5304 7644
rect 527 7616 793 7624
rect 1187 7616 1613 7624
rect 1627 7616 1833 7624
rect 4947 7616 5073 7624
rect 5296 7624 5304 7636
rect 5567 7633 5593 7641
rect 6227 7636 6273 7644
rect 6707 7636 6893 7644
rect 7796 7644 7804 7656
rect 7947 7656 8053 7664
rect 8196 7656 8633 7664
rect 8196 7644 8204 7656
rect 7007 7633 7033 7641
rect 7147 7633 7233 7641
rect 7796 7636 8204 7644
rect 8227 7636 8673 7644
rect 10116 7644 10124 7676
rect 10167 7676 10313 7684
rect 10507 7676 10613 7684
rect 10907 7676 11013 7684
rect 11147 7676 11233 7684
rect 11347 7676 11393 7684
rect 11567 7676 11673 7684
rect 11847 7676 11973 7684
rect 10976 7656 11444 7664
rect 8967 7636 9013 7644
rect 10116 7636 10293 7644
rect 10976 7644 10984 7656
rect 11436 7644 11444 7656
rect 12256 7647 12264 7676
rect 10307 7636 10353 7644
rect 10667 7633 10693 7641
rect 10927 7633 10973 7641
rect 11167 7633 11193 7641
rect 11447 7636 11653 7644
rect 11707 7633 11773 7641
rect 12147 7636 12173 7644
rect 12256 7636 12273 7647
rect 12260 7633 12273 7636
rect 5296 7616 5533 7624
rect 5676 7624 5684 7630
rect 5627 7616 5684 7624
rect 6447 7616 6553 7624
rect 7267 7616 7333 7624
rect 7687 7616 8153 7624
rect 8487 7616 8613 7624
rect 8727 7616 8893 7624
rect 9387 7616 9533 7624
rect 9847 7616 9893 7624
rect 10767 7616 10873 7624
rect 10887 7616 11053 7624
rect 11487 7616 11613 7624
rect 11667 7616 11933 7624
rect 247 7596 373 7604
rect 707 7596 813 7604
rect 907 7596 1073 7604
rect 2887 7596 2933 7604
rect 3467 7596 3573 7604
rect 4607 7596 4633 7604
rect 5607 7596 6173 7604
rect 6647 7596 7033 7604
rect 7287 7596 7353 7604
rect 7527 7596 7553 7604
rect 9367 7596 9953 7604
rect 10067 7596 10513 7604
rect 11307 7596 11493 7604
rect 11507 7596 11753 7604
rect 187 7576 233 7584
rect 3727 7576 4093 7584
rect 4567 7576 4653 7584
rect 4707 7576 5053 7584
rect 5367 7576 5633 7584
rect 5687 7576 6153 7584
rect 9107 7576 9913 7584
rect 10607 7576 10833 7584
rect 10847 7576 11113 7584
rect 11827 7576 12193 7584
rect 2647 7556 3153 7564
rect 3847 7556 4373 7564
rect 4387 7556 4953 7564
rect 5607 7556 5653 7564
rect 5727 7556 5793 7564
rect 6727 7556 6753 7564
rect 6967 7556 7013 7564
rect 7207 7556 7413 7564
rect 7427 7556 7533 7564
rect 7587 7556 8073 7564
rect 9127 7556 9273 7564
rect 10907 7556 11073 7564
rect 12127 7556 12193 7564
rect 3836 7544 3844 7553
rect 3627 7536 3844 7544
rect 5027 7536 5473 7544
rect 5587 7536 5613 7544
rect 5707 7536 5773 7544
rect 6167 7536 7553 7544
rect 8927 7536 8993 7544
rect 9047 7536 9173 7544
rect 9587 7536 9733 7544
rect 11967 7536 12033 7544
rect 3487 7516 3533 7524
rect 3687 7516 3793 7524
rect 5067 7516 5673 7524
rect 1947 7496 2193 7504
rect 2207 7496 2393 7504
rect 2467 7498 4533 7506
rect 5936 7504 5944 7533
rect 6367 7516 6573 7524
rect 6627 7516 7413 7524
rect 7547 7516 7733 7524
rect 8127 7516 8633 7524
rect 8687 7516 8953 7524
rect 9867 7516 10113 7524
rect 11527 7516 11793 7524
rect 5936 7500 6024 7504
rect 5936 7496 6027 7500
rect 6013 7487 6027 7496
rect 6107 7496 6173 7504
rect 7007 7496 7113 7504
rect 7227 7496 7353 7504
rect 7487 7496 8353 7504
rect 9167 7496 9333 7504
rect 9827 7496 10053 7504
rect 10687 7496 10713 7504
rect 807 7476 873 7484
rect 887 7476 1353 7484
rect 5087 7476 5413 7484
rect 5427 7476 5713 7484
rect 8947 7476 8973 7484
rect 9336 7484 9344 7493
rect 9336 7476 9393 7484
rect 9407 7476 9773 7484
rect 9787 7476 9804 7484
rect 547 7459 573 7467
rect 767 7459 933 7467
rect 947 7456 993 7464
rect 1327 7464 1340 7467
rect 1327 7453 1344 7464
rect 1407 7459 1453 7467
rect 1547 7459 1693 7467
rect 1707 7456 2133 7464
rect 2387 7460 2413 7468
rect 2647 7459 2713 7467
rect 2987 7459 3093 7467
rect 3367 7459 3473 7467
rect 593 7424 607 7433
rect 1336 7424 1344 7453
rect 2756 7424 2764 7456
rect 3567 7456 3693 7464
rect 3867 7459 4033 7467
rect 4207 7459 4313 7467
rect 4327 7456 4693 7464
rect 4747 7456 4793 7464
rect 5327 7456 5393 7464
rect 5487 7456 5653 7464
rect 5716 7456 6033 7464
rect 5716 7444 5724 7456
rect 6267 7456 6293 7464
rect 6836 7456 7013 7464
rect 4867 7436 5724 7444
rect 5747 7436 5773 7444
rect 6836 7444 6844 7456
rect 7247 7459 7373 7467
rect 7427 7456 7632 7464
rect 7646 7456 7647 7470
rect 5927 7433 6013 7441
rect 7107 7439 7213 7447
rect 7636 7444 7644 7456
rect 7667 7456 7773 7464
rect 8227 7459 8653 7467
rect 8827 7459 8893 7467
rect 9796 7464 9804 7476
rect 11027 7476 11073 7484
rect 11087 7476 11233 7484
rect 11947 7476 12033 7484
rect 9207 7456 9244 7464
rect 9796 7456 9853 7464
rect 7636 7436 7673 7444
rect 567 7420 607 7424
rect 567 7416 604 7420
rect 827 7413 893 7421
rect 1107 7413 1133 7421
rect 1687 7416 1913 7424
rect 2067 7413 2153 7421
rect 2207 7413 2253 7421
rect 2756 7416 2993 7424
rect 3107 7416 3253 7424
rect 3347 7413 3773 7421
rect 4027 7416 4173 7424
rect 4527 7413 4733 7421
rect 4907 7413 5553 7421
rect 6347 7416 6373 7424
rect 7053 7424 7067 7433
rect 7947 7433 8113 7441
rect 8767 7436 9184 7444
rect 6607 7413 6993 7421
rect 7053 7420 7084 7424
rect 7056 7416 7084 7420
rect 267 7396 653 7404
rect 747 7396 1413 7404
rect 2747 7396 2773 7404
rect 4307 7396 4453 7404
rect 4567 7396 4673 7404
rect 5607 7396 5673 7404
rect 5747 7396 5773 7404
rect 7076 7404 7084 7416
rect 7307 7413 7353 7421
rect 7407 7413 7513 7421
rect 8427 7416 8513 7424
rect 9176 7424 9184 7436
rect 9236 7427 9244 7456
rect 10007 7459 10593 7467
rect 10667 7459 10693 7467
rect 10887 7459 10953 7467
rect 9367 7433 9533 7441
rect 9687 7436 9793 7444
rect 10107 7433 10313 7441
rect 8927 7413 8993 7421
rect 9987 7413 10153 7421
rect 10587 7416 10713 7424
rect 6087 7393 6493 7401
rect 7076 7396 7113 7404
rect 7287 7396 7333 7404
rect 8307 7396 8373 7404
rect 9367 7396 9393 7404
rect 10996 7404 11004 7456
rect 11147 7456 11213 7464
rect 11027 7413 11093 7421
rect 11327 7416 11413 7424
rect 11427 7416 11493 7424
rect 10527 7396 11144 7404
rect 1067 7376 1373 7384
rect 1647 7376 1733 7384
rect 3007 7376 3353 7384
rect 3896 7376 4192 7384
rect 227 7356 313 7364
rect 1267 7356 1613 7364
rect 1827 7356 3773 7364
rect 3896 7364 3904 7376
rect 4227 7376 4273 7384
rect 4767 7376 5473 7384
rect 5487 7376 5713 7384
rect 6167 7376 6313 7384
rect 6407 7376 6553 7384
rect 6567 7376 6633 7384
rect 8616 7376 9244 7384
rect 8616 7367 8624 7376
rect 3787 7356 3904 7364
rect 3927 7356 4873 7364
rect 4967 7356 5333 7364
rect 5347 7356 5473 7364
rect 5647 7356 5733 7364
rect 5936 7356 6233 7364
rect 2247 7336 2433 7344
rect 3947 7336 5513 7344
rect 5936 7344 5944 7356
rect 8107 7356 8133 7364
rect 8147 7356 8613 7364
rect 9236 7364 9244 7376
rect 9827 7376 10013 7384
rect 11136 7384 11144 7396
rect 11767 7396 11993 7404
rect 11136 7376 11633 7384
rect 12047 7376 12113 7384
rect 9236 7356 9693 7364
rect 9707 7356 9753 7364
rect 9767 7356 10473 7364
rect 5747 7336 5944 7344
rect 6087 7336 6133 7344
rect 6187 7336 6313 7344
rect 6627 7336 6673 7344
rect 6867 7336 7153 7344
rect 7567 7336 9093 7344
rect 11687 7336 12053 7344
rect 1627 7316 2713 7324
rect 2987 7316 3133 7324
rect 3847 7316 5173 7324
rect 6027 7316 6353 7324
rect 6616 7324 6624 7333
rect 6507 7316 6624 7324
rect 6887 7316 7213 7324
rect 7627 7316 8113 7324
rect 8347 7316 8393 7324
rect 12007 7316 12093 7324
rect 1847 7296 3793 7304
rect 3987 7296 4073 7304
rect 4127 7296 4253 7304
rect 4347 7296 5733 7304
rect 6367 7296 6433 7304
rect 6527 7296 6773 7304
rect 7587 7296 7953 7304
rect 8147 7296 8173 7304
rect 8187 7296 9273 7304
rect 9287 7296 9833 7304
rect 9847 7296 10653 7304
rect 707 7276 1813 7284
rect 2007 7276 3033 7284
rect 3087 7276 4853 7284
rect 7787 7276 7833 7284
rect 9387 7276 9413 7284
rect 10047 7276 10573 7284
rect 1667 7256 1973 7264
rect 3367 7256 4893 7264
rect 5267 7256 5553 7264
rect 6007 7256 6513 7264
rect 7107 7256 8073 7264
rect 8127 7256 8873 7264
rect 10867 7256 10953 7264
rect 10967 7256 11713 7264
rect 11727 7256 12113 7264
rect 1267 7236 1573 7244
rect 2567 7236 2773 7244
rect 3947 7236 4353 7244
rect 4627 7236 4773 7244
rect 5307 7236 5753 7244
rect 5767 7236 6193 7244
rect 6667 7236 9113 7244
rect 9587 7236 9733 7244
rect 10167 7236 10493 7244
rect 1887 7216 2593 7224
rect 3007 7216 3813 7224
rect 3887 7216 4393 7224
rect 4447 7216 5073 7224
rect 5147 7216 5404 7224
rect 227 7196 673 7204
rect 1827 7196 1853 7204
rect 2687 7196 3633 7204
rect 3687 7196 3753 7204
rect 3947 7196 4053 7204
rect 5067 7196 5353 7204
rect 5396 7204 5404 7216
rect 5627 7216 6153 7224
rect 6427 7216 6613 7224
rect 6947 7216 7073 7224
rect 7167 7216 7313 7224
rect 7447 7216 7893 7224
rect 8447 7216 8833 7224
rect 9887 7216 9993 7224
rect 5396 7196 5773 7204
rect 5827 7196 7093 7204
rect 7247 7196 7413 7204
rect 8567 7196 8753 7204
rect 8867 7196 8973 7204
rect 10587 7196 10793 7204
rect 507 7176 653 7184
rect 667 7176 1293 7184
rect 3147 7176 3413 7184
rect 4307 7176 5133 7184
rect 5527 7176 5753 7184
rect 6527 7176 7033 7184
rect 7467 7176 7493 7184
rect 7807 7179 7893 7187
rect 9907 7179 9953 7187
rect 10847 7176 10973 7184
rect 267 7159 313 7167
rect 447 7159 532 7167
rect 567 7156 593 7164
rect 687 7159 773 7167
rect 827 7159 873 7167
rect 887 7156 1053 7164
rect 1076 7156 1093 7164
rect 1107 7156 1333 7164
rect 1347 7159 1473 7167
rect 1587 7156 1784 7164
rect 1076 7144 1084 7156
rect 836 7136 1084 7144
rect 1776 7144 1784 7156
rect 1827 7156 1944 7164
rect 1936 7147 1944 7156
rect 2487 7156 2553 7164
rect 2667 7156 2813 7164
rect 3187 7159 3213 7167
rect 3707 7159 3813 7167
rect 3987 7156 4133 7164
rect 4147 7159 4193 7167
rect 5407 7166 5524 7167
rect 5407 7159 5513 7166
rect 1776 7136 1793 7144
rect 247 7116 333 7124
rect 467 7116 513 7124
rect 836 7124 844 7136
rect 1807 7136 1904 7144
rect 1936 7136 1953 7147
rect 587 7116 793 7124
rect 907 7116 1073 7124
rect 1147 7116 1313 7124
rect 1607 7116 1773 7124
rect 1896 7124 1904 7136
rect 1940 7133 1953 7136
rect 2007 7139 2093 7147
rect 2916 7136 3013 7144
rect 2916 7123 2924 7136
rect 4236 7127 4244 7156
rect 5827 7159 5873 7167
rect 5927 7159 5953 7167
rect 6207 7159 6273 7167
rect 6387 7159 6433 7167
rect 6487 7159 6553 7167
rect 6627 7159 6713 7167
rect 6767 7159 6793 7167
rect 7047 7159 7093 7167
rect 4887 7136 5064 7144
rect 3047 7116 3153 7124
rect 3447 7113 3533 7121
rect 3827 7116 3953 7124
rect 4067 7113 4173 7121
rect 4236 7116 4253 7127
rect 4240 7113 4253 7116
rect 4367 7112 4553 7120
rect 4647 7116 4733 7124
rect 5056 7124 5064 7136
rect 7127 7136 7193 7144
rect 5056 7116 5373 7124
rect 5427 7116 5533 7124
rect 5727 7113 5853 7121
rect 6187 7116 6373 7124
rect 6427 7116 6613 7124
rect 6627 7116 6933 7124
rect 7256 7124 7264 7153
rect 7336 7144 7344 7173
rect 8087 7159 8273 7167
rect 8627 7159 8653 7167
rect 9067 7159 9133 7167
rect 9187 7159 9233 7167
rect 10147 7156 10373 7164
rect 10427 7159 10553 7167
rect 7336 7136 7413 7144
rect 7647 7139 7732 7147
rect 7767 7136 7853 7144
rect 8036 7144 8044 7156
rect 8036 7136 8173 7144
rect 9267 7136 9353 7144
rect 9367 7133 9533 7141
rect 9587 7139 9733 7147
rect 9867 7136 9933 7144
rect 10636 7144 10644 7156
rect 11167 7159 11193 7167
rect 11407 7156 11473 7164
rect 11627 7156 11753 7164
rect 11987 7156 12073 7164
rect 10347 7136 10644 7144
rect 10896 7127 10904 7153
rect 6947 7116 7053 7124
rect 7256 7116 7353 7124
rect 7447 7116 7493 7124
rect 8007 7116 8053 7124
rect 8767 7113 8833 7121
rect 9027 7113 9113 7121
rect 10096 7116 10393 7124
rect 236 7103 413 7104
rect 247 7096 413 7103
rect 2387 7096 2573 7104
rect 2587 7096 2653 7104
rect 3187 7096 3213 7104
rect 3587 7096 3633 7104
rect 3687 7096 3873 7104
rect 4987 7096 5033 7104
rect 1067 7076 1193 7084
rect 1993 7084 2007 7093
rect 5087 7096 5173 7104
rect 5307 7096 5353 7104
rect 5747 7096 6013 7104
rect 6507 7096 6533 7104
rect 6547 7096 6693 7104
rect 7247 7096 7333 7104
rect 7747 7096 7853 7104
rect 7987 7096 8593 7104
rect 8947 7096 9153 7104
rect 10096 7104 10104 7116
rect 10507 7113 10693 7121
rect 11227 7116 11453 7124
rect 11647 7113 11773 7121
rect 9507 7096 10104 7104
rect 11947 7096 12033 7104
rect 1867 7080 2007 7084
rect 1867 7076 2004 7080
rect 2367 7076 2673 7084
rect 2947 7076 3133 7084
rect 3707 7076 3733 7084
rect 4187 7076 4253 7084
rect 4527 7076 4913 7084
rect 5127 7076 5253 7084
rect 5447 7076 5493 7084
rect 6127 7076 6213 7084
rect 6387 7076 6413 7084
rect 6567 7076 6733 7084
rect 7107 7076 7293 7084
rect 8087 7076 8252 7084
rect 8287 7076 8393 7084
rect 9087 7076 9133 7084
rect 9187 7076 9433 7084
rect 9447 7076 9473 7084
rect 11167 7076 11253 7084
rect 12067 7076 12093 7084
rect 1227 7056 1353 7064
rect 2956 7056 3853 7064
rect 2956 7047 2964 7056
rect 4647 7056 4793 7064
rect 5347 7056 5473 7064
rect 5807 7056 5932 7064
rect 5967 7056 6513 7064
rect 6787 7056 7133 7064
rect 7467 7056 7913 7064
rect 7653 7047 7667 7056
rect 7967 7056 8053 7064
rect 8667 7056 9493 7064
rect 9547 7056 9973 7064
rect 1527 7036 2173 7044
rect 2547 7036 2873 7044
rect 2947 7036 2964 7047
rect 2947 7033 2960 7036
rect 3887 7036 4133 7044
rect 4227 7036 4972 7044
rect 5007 7036 5813 7044
rect 5987 7036 6453 7044
rect 6547 7036 7213 7044
rect 7907 7036 8033 7044
rect 8607 7036 8813 7044
rect 9827 7036 9953 7044
rect 10227 7036 10513 7044
rect 10667 7036 10793 7044
rect 10807 7036 11493 7044
rect 2447 7016 2593 7024
rect 2927 7016 2973 7024
rect 3347 7016 3553 7024
rect 3907 7016 4853 7024
rect 4876 7016 5893 7024
rect 1927 6996 2293 7004
rect 3027 6996 3253 7004
rect 3267 6996 3613 7004
rect 4007 6996 4293 7004
rect 4876 7004 4884 7016
rect 5947 7016 6793 7024
rect 7247 7016 7313 7024
rect 7707 7016 7833 7024
rect 8227 7016 9473 7024
rect 9527 7016 9613 7024
rect 9687 7016 10013 7024
rect 11527 7016 11573 7024
rect 4767 6996 4884 7004
rect 4987 6996 5372 7004
rect 5407 6996 5893 7004
rect 6267 6996 6333 7004
rect 6347 6996 6653 7004
rect 6887 6996 6993 7004
rect 7467 6996 8164 7004
rect 687 6976 1113 6984
rect 1127 6976 1173 6984
rect 1407 6976 1533 6984
rect 1547 6976 2033 6984
rect 2687 6976 2853 6984
rect 3307 6976 3593 6984
rect 3607 6976 3653 6984
rect 4127 6976 4193 6984
rect 4807 6976 5013 6984
rect 5427 6976 5713 6984
rect 5947 6976 6233 6984
rect 6247 6976 7013 6984
rect 7147 6976 7213 6984
rect 7267 6976 7393 6984
rect 8156 6984 8164 6996
rect 8547 6996 8893 7004
rect 9447 6996 10473 7004
rect 10707 6996 10873 7004
rect 10967 6996 11073 7004
rect 11327 6996 11884 7004
rect 8156 6976 8553 6984
rect 8756 6976 9053 6984
rect 2887 6956 3053 6964
rect 4247 6956 4693 6964
rect 5876 6956 6153 6964
rect 507 6939 573 6947
rect 787 6939 893 6947
rect 947 6939 1013 6947
rect 1667 6936 1752 6944
rect 1787 6939 1833 6947
rect 1856 6936 1873 6944
rect 2107 6939 2133 6947
rect 2227 6939 2573 6947
rect 1856 6924 1864 6936
rect 1467 6916 1864 6924
rect 2956 6924 2964 6937
rect 3516 6936 3553 6944
rect 3647 6940 3913 6948
rect 2956 6916 3133 6924
rect 3516 6907 3524 6936
rect 3967 6936 4213 6944
rect 4667 6936 4773 6944
rect 4867 6936 5093 6944
rect 5256 6936 5393 6944
rect 3947 6916 4233 6924
rect 547 6896 733 6904
rect 747 6893 833 6901
rect 1387 6896 1613 6904
rect 1907 6896 2193 6904
rect 2207 6893 2233 6901
rect 2307 6896 2933 6904
rect 3067 6896 3273 6904
rect 3587 6893 3653 6901
rect 3727 6896 3753 6904
rect 3767 6894 3813 6902
rect 1867 6876 2153 6884
rect 2467 6876 2693 6884
rect 3927 6876 3993 6884
rect 4087 6876 4173 6884
rect 4276 6884 4284 6913
rect 4507 6913 4633 6921
rect 5256 6924 5264 6936
rect 4676 6887 4684 6913
rect 4953 6907 4967 6913
rect 5247 6916 5264 6924
rect 5587 6916 5833 6924
rect 4707 6896 4873 6904
rect 4947 6900 4967 6907
rect 4947 6896 4964 6900
rect 4947 6893 4960 6896
rect 5647 6896 5793 6904
rect 5876 6904 5884 6956
rect 7067 6956 7124 6964
rect 6427 6939 6613 6947
rect 6707 6939 6853 6947
rect 6893 6944 6907 6953
rect 6893 6940 6933 6944
rect 6896 6936 6933 6940
rect 7116 6944 7124 6956
rect 8007 6956 8113 6964
rect 8756 6964 8764 6976
rect 9067 6976 9373 6984
rect 11767 6976 11853 6984
rect 8427 6956 8764 6964
rect 9927 6956 10213 6964
rect 10287 6956 10773 6964
rect 11247 6956 11333 6964
rect 11487 6956 11553 6964
rect 11607 6956 11633 6964
rect 7116 6936 7533 6944
rect 7856 6936 7973 6944
rect 6047 6916 6773 6924
rect 7107 6916 7524 6924
rect 7856 6924 7864 6936
rect 8107 6936 8313 6944
rect 8327 6936 8393 6944
rect 8407 6936 8693 6944
rect 8707 6939 8773 6947
rect 8796 6936 9033 6944
rect 5927 6893 5973 6901
rect 6087 6896 6133 6904
rect 6147 6893 6733 6901
rect 7347 6896 7473 6904
rect 7516 6904 7524 6916
rect 7596 6904 7604 6916
rect 8033 6904 8047 6913
rect 7516 6896 7604 6904
rect 8016 6896 8173 6904
rect 4227 6876 4284 6884
rect 5107 6876 5933 6884
rect 6827 6876 7053 6884
rect 7567 6876 7693 6884
rect 8016 6884 8024 6896
rect 8796 6904 8804 6936
rect 9167 6939 9313 6947
rect 9807 6939 9873 6947
rect 10127 6939 10173 6947
rect 10727 6938 10753 6946
rect 10987 6939 11013 6947
rect 10716 6924 10724 6935
rect 11056 6924 11064 6936
rect 11467 6936 11573 6944
rect 11876 6949 11884 6996
rect 11807 6938 11833 6946
rect 12007 6939 12113 6947
rect 11613 6924 11627 6933
rect 10716 6916 11064 6924
rect 11596 6920 11627 6924
rect 11596 6916 11624 6920
rect 8847 6893 8893 6901
rect 9087 6896 9253 6904
rect 9347 6896 9793 6904
rect 11596 6904 11604 6916
rect 9947 6893 9993 6901
rect 10247 6893 10273 6901
rect 10547 6893 10573 6901
rect 11047 6896 11293 6904
rect 11567 6896 11604 6904
rect 8167 6876 8293 6884
rect 11747 6876 11833 6884
rect 12107 6876 12193 6884
rect 227 6856 313 6864
rect 327 6856 473 6864
rect 807 6856 873 6864
rect 1287 6856 2313 6864
rect 2327 6856 3473 6864
rect 3547 6856 3713 6864
rect 4027 6856 4133 6864
rect 4667 6856 4833 6864
rect 4847 6856 5393 6864
rect 5627 6856 5673 6864
rect 5727 6856 6073 6864
rect 6167 6856 6913 6864
rect 6927 6856 7373 6864
rect 7387 6856 7804 6864
rect 1307 6836 3653 6844
rect 3747 6836 4053 6844
rect 4767 6836 4913 6844
rect 4967 6836 5573 6844
rect 5887 6836 6053 6844
rect 6127 6836 6213 6844
rect 7127 6836 7213 6844
rect 7796 6844 7804 6856
rect 8567 6856 8693 6864
rect 8707 6856 9093 6864
rect 9107 6856 9413 6864
rect 9427 6856 9853 6864
rect 9867 6856 10153 6864
rect 10467 6856 10753 6864
rect 10767 6856 10853 6864
rect 11347 6856 11533 6864
rect 11547 6856 11673 6864
rect 7407 6836 7784 6844
rect 7796 6836 8073 6844
rect 407 6816 933 6824
rect 1047 6816 1113 6824
rect 1127 6816 1853 6824
rect 2107 6816 3153 6824
rect 3336 6816 4473 6824
rect 3336 6807 3344 6816
rect 5367 6816 5473 6824
rect 5487 6816 7633 6824
rect 7776 6824 7784 6836
rect 7776 6816 8213 6824
rect 8547 6816 9213 6824
rect 12087 6816 12173 6824
rect 2547 6796 3333 6804
rect 3507 6796 3572 6804
rect 3607 6796 3733 6804
rect 4607 6796 4793 6804
rect 5087 6796 5253 6804
rect 5587 6796 5993 6804
rect 6247 6796 7133 6804
rect 7147 6796 7613 6804
rect 7667 6796 8253 6804
rect 9907 6796 10133 6804
rect 11607 6796 11813 6804
rect 11827 6796 11973 6804
rect 267 6776 293 6784
rect 307 6776 1993 6784
rect 2527 6776 3373 6784
rect 3547 6776 3953 6784
rect 4067 6776 4753 6784
rect 5507 6776 5533 6784
rect 6587 6776 7453 6784
rect 7687 6776 8193 6784
rect 9247 6776 10673 6784
rect 787 6756 873 6764
rect 887 6756 1073 6764
rect 1087 6756 1893 6764
rect 3007 6756 3353 6764
rect 3487 6756 3913 6764
rect 4847 6756 4953 6764
rect 5287 6756 5473 6764
rect 5787 6756 6073 6764
rect 6707 6756 7093 6764
rect 7287 6756 7353 6764
rect 7587 6756 8453 6764
rect 8747 6756 8873 6764
rect 9387 6756 10093 6764
rect 11307 6756 11453 6764
rect 1347 6736 2493 6744
rect 2747 6736 4913 6744
rect 5107 6736 5433 6744
rect 6027 6736 6333 6744
rect 7153 6744 7167 6753
rect 6356 6736 7493 6744
rect 307 6716 953 6724
rect 2167 6716 2713 6724
rect 2767 6716 3273 6724
rect 3327 6716 3593 6724
rect 3667 6716 4333 6724
rect 4467 6716 4653 6724
rect 6356 6724 6364 6736
rect 7767 6736 8133 6744
rect 8187 6736 8333 6744
rect 8487 6736 9013 6744
rect 9207 6736 10233 6744
rect 11007 6736 11133 6744
rect 11227 6736 11953 6744
rect 4747 6716 6364 6724
rect 7387 6716 7653 6724
rect 8467 6716 9053 6724
rect 9133 6724 9147 6733
rect 9067 6720 9147 6724
rect 9067 6716 9144 6720
rect 9267 6716 9473 6724
rect 9487 6716 9653 6724
rect 9667 6716 9813 6724
rect 10487 6716 11393 6724
rect 12247 6716 12313 6724
rect 2807 6696 3613 6704
rect 3636 6696 5352 6704
rect -24 6676 513 6684
rect 1887 6676 2153 6684
rect 2347 6676 2853 6684
rect 2867 6676 3113 6684
rect 3636 6684 3644 6696
rect 5387 6696 5464 6704
rect 3127 6676 3644 6684
rect 3707 6676 3813 6684
rect 3987 6676 4393 6684
rect 5456 6684 5464 6696
rect 5607 6696 5673 6704
rect 5767 6696 6353 6704
rect 6607 6696 6873 6704
rect 8567 6696 8593 6704
rect 10107 6696 10913 6704
rect 4887 6676 5444 6684
rect 5456 6676 5733 6684
rect 447 6656 473 6664
rect 2207 6656 2273 6664
rect 3287 6656 3453 6664
rect 3527 6656 3673 6664
rect 3787 6656 3893 6664
rect 5436 6664 5444 6676
rect 6447 6676 6533 6684
rect 7407 6676 7673 6684
rect 8527 6676 8713 6684
rect 9267 6676 9313 6684
rect 9567 6676 9744 6684
rect 5436 6656 6033 6664
rect 7187 6656 7213 6664
rect 8347 6659 8453 6667
rect 8540 6664 8553 6667
rect 8536 6653 8553 6664
rect -24 6636 193 6644
rect 827 6636 973 6644
rect 987 6636 1113 6644
rect 1407 6639 1453 6647
rect 1356 6624 1364 6636
rect 1507 6636 1633 6644
rect 1927 6639 1973 6647
rect 2167 6636 2433 6644
rect 2627 6639 2693 6647
rect 2967 6639 3033 6647
rect 3247 6639 3353 6647
rect 4027 6639 4233 6647
rect 4507 6639 4633 6647
rect 4887 6639 4953 6647
rect 5067 6639 5093 6647
rect 5147 6639 5293 6647
rect 1356 6616 1713 6624
rect 2787 6616 3113 6624
rect 3136 6616 3313 6624
rect 467 6596 493 6604
rect 547 6593 633 6601
rect 707 6596 753 6604
rect 967 6596 1373 6604
rect 1427 6593 1493 6601
rect 1947 6596 2093 6604
rect 2147 6593 2333 6601
rect 2507 6596 2673 6604
rect 3136 6604 3144 6616
rect 3496 6624 3504 6636
rect 3496 6616 3593 6624
rect 3707 6616 3933 6624
rect 5416 6624 5424 6636
rect 5927 6636 6053 6644
rect 6147 6639 6193 6647
rect 6507 6639 6673 6647
rect 6727 6639 6773 6647
rect 6827 6640 6904 6644
rect 6827 6636 6907 6640
rect 7587 6636 7653 6644
rect 5327 6616 5533 6624
rect 2807 6596 3144 6604
rect 3187 6596 3213 6604
rect 3687 6593 3733 6601
rect 3967 6593 3993 6601
rect 4127 6596 4293 6604
rect 5367 6596 5513 6604
rect 5616 6587 5624 6633
rect 6893 6627 6907 6636
rect 7707 6639 7813 6647
rect 7867 6636 8033 6644
rect 8536 6644 8544 6653
rect 8476 6636 8544 6644
rect 8556 6636 8573 6644
rect 5707 6593 5733 6601
rect 6067 6593 6173 6601
rect 6487 6596 6713 6604
rect 267 6576 293 6584
rect 807 6576 913 6584
rect 1107 6576 1233 6584
rect 1487 6576 1833 6584
rect 1887 6576 2033 6584
rect 2047 6576 2133 6584
rect 2467 6576 2513 6584
rect 3267 6576 3413 6584
rect 3427 6576 3633 6584
rect 4587 6576 4653 6584
rect 5616 6576 5633 6587
rect 5620 6573 5633 6576
rect 5847 6576 5993 6584
rect 7036 6584 7044 6616
rect 7187 6616 7213 6624
rect 7307 6613 7373 6621
rect 8476 6624 8484 6636
rect 8187 6616 8484 6624
rect 8556 6607 8564 6636
rect 9507 6639 9613 6647
rect 9736 6644 9744 6676
rect 10187 6676 10333 6684
rect 10947 6676 11153 6684
rect 11287 6676 11413 6684
rect 12247 6676 12293 6684
rect 9967 6656 10033 6664
rect 10467 6656 10593 6664
rect 11867 6656 11913 6664
rect 9736 6636 9824 6644
rect 10367 6636 10433 6644
rect 8907 6619 9233 6627
rect 9273 6624 9287 6633
rect 9816 6630 9824 6636
rect 10547 6639 10573 6647
rect 10647 6636 10893 6644
rect 10967 6636 11013 6644
rect 11427 6636 11593 6644
rect 11887 6644 11900 6647
rect 12156 6646 12193 6647
rect 11887 6633 11904 6644
rect 9273 6620 9344 6624
rect 9276 6616 9344 6620
rect 7527 6596 7833 6604
rect 8047 6596 8544 6604
rect 7036 6576 7333 6584
rect 7487 6576 7613 6584
rect 7727 6576 7793 6584
rect 7987 6576 8333 6584
rect 8536 6584 8544 6596
rect 8707 6596 9093 6604
rect 9336 6604 9344 6616
rect 9387 6616 9693 6624
rect 11896 6624 11904 6633
rect 12167 6639 12193 6646
rect 12207 6636 12273 6644
rect 9987 6613 10013 6621
rect 11896 6620 11984 6624
rect 11896 6616 11987 6620
rect 11973 6607 11987 6616
rect 10247 6593 10333 6601
rect 10547 6596 10593 6604
rect 10687 6596 10873 6604
rect 11187 6593 11293 6601
rect 11367 6593 11433 6601
rect 11607 6593 11653 6601
rect 8536 6576 9173 6584
rect 9567 6576 9953 6584
rect 10367 6576 10493 6584
rect 11947 6576 11993 6584
rect 12047 6576 12193 6584
rect 467 6556 673 6564
rect 1507 6556 1853 6564
rect 1956 6556 2793 6564
rect 1956 6544 1964 6556
rect 3527 6556 3573 6564
rect 3627 6556 4033 6564
rect 4207 6556 4333 6564
rect 4347 6556 4613 6564
rect 4967 6556 5333 6564
rect 5407 6556 5453 6564
rect 5547 6556 5933 6564
rect 6307 6556 6493 6564
rect 7236 6556 7353 6564
rect 1067 6536 1964 6544
rect 2007 6536 2173 6544
rect 2827 6536 2973 6544
rect 5576 6540 5873 6544
rect 5573 6536 5873 6540
rect 5573 6527 5587 6536
rect 7236 6544 7244 6556
rect 7647 6556 7853 6564
rect 8007 6556 8553 6564
rect 8647 6556 8653 6564
rect 8667 6556 10153 6564
rect 10787 6556 10913 6564
rect 11887 6556 11913 6564
rect 6227 6536 7244 6544
rect 7747 6536 7913 6544
rect 7927 6536 8493 6544
rect 8547 6536 8593 6544
rect 9067 6536 9153 6544
rect 9307 6536 9413 6544
rect 10007 6536 10333 6544
rect 10447 6536 12213 6544
rect 1107 6516 1173 6524
rect 1467 6516 1913 6524
rect 2267 6516 4093 6524
rect 4207 6516 4933 6524
rect 5007 6516 5493 6524
rect 7247 6516 7633 6524
rect 9507 6516 9833 6524
rect 9967 6516 10353 6524
rect 10547 6516 11113 6524
rect 11127 6516 11433 6524
rect 587 6496 1053 6504
rect 1227 6496 1273 6504
rect 2287 6496 2913 6504
rect 3047 6496 3173 6504
rect 3187 6496 3593 6504
rect 3607 6496 3673 6504
rect 3687 6496 4544 6504
rect 4536 6487 4544 6496
rect 5387 6496 5453 6504
rect 5627 6496 5653 6504
rect 6767 6496 6864 6504
rect 267 6476 1893 6484
rect 3167 6476 3253 6484
rect 4087 6476 4253 6484
rect 4547 6476 4953 6484
rect 5267 6476 5973 6484
rect 6047 6476 6433 6484
rect 6647 6476 6713 6484
rect 6856 6484 6864 6496
rect 7567 6496 7693 6504
rect 7767 6496 8093 6504
rect 8347 6496 8693 6504
rect 10347 6496 11593 6504
rect 11607 6496 11693 6504
rect 6856 6476 7333 6484
rect 7507 6476 7993 6484
rect 8267 6476 8373 6484
rect 8987 6476 9113 6484
rect 12107 6476 12213 6484
rect 527 6456 1153 6464
rect 2127 6456 2153 6464
rect 2167 6456 2352 6464
rect 2387 6456 2733 6464
rect 2927 6456 3853 6464
rect 4367 6456 4513 6464
rect 4687 6456 5224 6464
rect 1787 6436 2693 6444
rect 3227 6436 3293 6444
rect 4947 6436 5013 6444
rect 5216 6444 5224 6456
rect 6267 6456 6693 6464
rect 6847 6456 7293 6464
rect 7647 6456 7973 6464
rect 8327 6456 8913 6464
rect 9087 6456 9433 6464
rect 9487 6456 9653 6464
rect 10227 6456 10613 6464
rect 10627 6456 10833 6464
rect 11487 6456 11613 6464
rect 11767 6456 11913 6464
rect 11967 6456 12273 6464
rect 5216 6436 5453 6444
rect 5607 6436 5653 6444
rect 5987 6436 6653 6444
rect 7467 6436 8013 6444
rect 8527 6436 8573 6444
rect 9507 6436 9553 6444
rect 9607 6436 9713 6444
rect 10267 6436 10293 6444
rect 10747 6436 10813 6444
rect 12067 6436 12093 6444
rect -24 6416 573 6424
rect 647 6419 733 6427
rect 1096 6404 1104 6416
rect 1147 6416 1273 6424
rect 2847 6419 2973 6427
rect 3027 6416 3093 6424
rect 3167 6416 3573 6424
rect 3827 6416 4053 6424
rect 4147 6416 4173 6424
rect 4187 6416 4313 6424
rect 4407 6416 4593 6424
rect 5207 6416 5464 6424
rect 1096 6400 1124 6404
rect 1096 6396 1127 6400
rect 1113 6387 1127 6396
rect -24 6376 193 6384
rect 447 6376 473 6384
rect 587 6376 753 6384
rect 947 6376 973 6384
rect 987 6373 1033 6381
rect 1196 6396 1213 6404
rect 1196 6367 1204 6396
rect 1427 6393 1693 6401
rect 1707 6396 2173 6404
rect 1436 6376 1953 6384
rect 1436 6364 1444 6376
rect 2627 6376 2713 6384
rect 2727 6376 2993 6384
rect 3047 6373 3153 6381
rect 3607 6373 3693 6381
rect 3807 6376 4153 6384
rect 4307 6376 4373 6384
rect 4607 6373 4633 6381
rect 4687 6373 4713 6381
rect 4767 6376 4973 6384
rect 5387 6376 5413 6384
rect 5456 6384 5464 6416
rect 5456 6376 5473 6384
rect 5496 6367 5504 6416
rect 5627 6416 5804 6424
rect 6227 6419 6293 6427
rect 6987 6416 7173 6424
rect 5796 6404 5804 6416
rect 7267 6419 7473 6427
rect 7567 6419 7633 6427
rect 7787 6416 7993 6424
rect 8287 6419 8313 6427
rect 8367 6419 8393 6427
rect 8627 6416 8833 6424
rect 8856 6416 8873 6424
rect 9047 6419 9153 6427
rect 9467 6416 9744 6424
rect 9767 6419 9953 6427
rect 5556 6367 5564 6393
rect 5596 6367 5604 6396
rect 5927 6396 5993 6404
rect 8553 6404 8567 6413
rect 8553 6400 8604 6404
rect 8556 6396 8604 6400
rect 6147 6376 6193 6384
rect 6307 6376 6453 6384
rect 6507 6376 7033 6384
rect 7187 6373 7233 6381
rect 7287 6376 7513 6384
rect 7527 6376 7673 6384
rect 7827 6376 7913 6384
rect 8087 6376 8273 6384
rect 8596 6384 8604 6396
rect 8856 6387 8864 6416
rect 9736 6404 9744 6416
rect 11047 6416 11093 6424
rect 11167 6426 11244 6427
rect 11167 6419 11233 6426
rect 11247 6416 11373 6424
rect 11667 6416 11733 6424
rect 12047 6416 12144 6424
rect 9736 6396 9913 6404
rect 11416 6396 11593 6404
rect 11416 6385 11424 6396
rect 8947 6376 9433 6384
rect 10027 6373 10213 6381
rect 10287 6373 10373 6381
rect 10487 6373 10553 6381
rect 10767 6373 10793 6381
rect 10887 6373 11013 6381
rect 11547 6373 11713 6381
rect 11787 6376 11873 6384
rect 1287 6356 1444 6364
rect 2407 6356 3293 6364
rect 3307 6356 3393 6364
rect 3467 6356 3793 6364
rect 5587 6356 5604 6367
rect 5587 6353 5600 6356
rect 5627 6356 5653 6364
rect 5967 6353 6093 6361
rect 6707 6356 6773 6364
rect 8007 6356 8253 6364
rect 8647 6356 8753 6364
rect 9187 6356 9273 6364
rect 9447 6356 9573 6364
rect 11487 6356 11753 6364
rect 11767 6356 11973 6364
rect 12136 6364 12144 6416
rect 12336 6387 12344 6413
rect 12136 6356 12233 6364
rect 767 6336 793 6344
rect 1827 6336 1873 6344
rect 2487 6336 2533 6344
rect 3027 6336 3173 6344
rect 3567 6336 3673 6344
rect 3727 6336 4193 6344
rect 4267 6336 4373 6344
rect 4527 6336 4673 6344
rect 5367 6336 5473 6344
rect 6527 6336 7013 6344
rect 7447 6336 7813 6344
rect 8347 6336 9033 6344
rect 9747 6336 9973 6344
rect 9987 6336 10133 6344
rect 10247 6336 10413 6344
rect 10807 6336 11153 6344
rect 1047 6316 1253 6324
rect 1587 6316 1773 6324
rect 2587 6316 2753 6324
rect 3007 6316 3153 6324
rect 3647 6316 4493 6324
rect 5307 6324 5320 6327
rect 5307 6313 5324 6324
rect 5567 6316 5613 6324
rect 5967 6316 6013 6324
rect 9847 6316 10053 6324
rect 11887 6316 12093 6324
rect 2807 6296 4693 6304
rect 4747 6296 5253 6304
rect 5316 6304 5324 6313
rect 5316 6296 5513 6304
rect 6107 6296 6593 6304
rect 6607 6296 6673 6304
rect 8416 6296 8453 6304
rect 887 6276 1073 6284
rect 1087 6276 1213 6284
rect 1687 6276 1993 6284
rect 2287 6276 2333 6284
rect 2347 6276 2513 6284
rect 3067 6276 3433 6284
rect 3907 6276 4044 6284
rect 2667 6256 3793 6264
rect 4036 6264 4044 6276
rect 4067 6276 4413 6284
rect 5307 6276 5593 6284
rect 8416 6284 8424 6296
rect 9147 6296 9633 6304
rect 9787 6296 10793 6304
rect 11616 6296 12153 6304
rect 11616 6284 11624 6296
rect 7447 6276 8424 6284
rect 10176 6276 11624 6284
rect 4036 6256 4193 6264
rect 4467 6256 5053 6264
rect 5227 6256 5953 6264
rect 6927 6256 7113 6264
rect 7647 6256 8433 6264
rect 8447 6256 8513 6264
rect 10176 6264 10184 6276
rect 11907 6276 12093 6284
rect 9687 6256 10184 6264
rect 10207 6256 10693 6264
rect 11947 6256 12313 6264
rect 847 6236 1913 6244
rect 1987 6244 2000 6247
rect 1987 6233 2004 6244
rect 2247 6236 3064 6244
rect 867 6216 1653 6224
rect 1996 6224 2004 6233
rect 1996 6216 2673 6224
rect 2827 6216 2973 6224
rect 3056 6224 3064 6236
rect 3167 6236 3273 6244
rect 3527 6236 3593 6244
rect 3947 6236 5033 6244
rect 5227 6236 5792 6244
rect 5827 6236 6113 6244
rect 6367 6236 6873 6244
rect 7047 6236 7873 6244
rect 8007 6236 8973 6244
rect 9947 6236 10173 6244
rect 11147 6236 11753 6244
rect 3056 6216 4233 6224
rect 4247 6216 8013 6224
rect -24 6196 213 6204
rect 447 6196 1113 6204
rect 3147 6196 3393 6204
rect 3407 6196 3713 6204
rect 3727 6196 3833 6204
rect 3987 6196 4173 6204
rect 5047 6196 5213 6204
rect 5267 6196 6093 6204
rect 6207 6196 6413 6204
rect 6427 6196 6793 6204
rect 6947 6196 7973 6204
rect 9487 6196 9993 6204
rect 10007 6196 10273 6204
rect 10707 6196 11973 6204
rect 627 6176 913 6184
rect 1007 6176 1813 6184
rect 2067 6176 2364 6184
rect -24 6156 13 6164
rect 1776 6156 1833 6164
rect 1547 6139 1593 6147
rect 1607 6139 1693 6147
rect 1776 6147 1784 6156
rect 2356 6164 2364 6176
rect 2476 6176 2813 6184
rect 2476 6164 2484 6176
rect 2887 6176 3033 6184
rect 3087 6176 3113 6184
rect 3127 6176 3673 6184
rect 3767 6176 4033 6184
rect 4287 6176 4433 6184
rect 4507 6176 4733 6184
rect 5647 6176 5693 6184
rect 5767 6176 5893 6184
rect 7187 6176 7313 6184
rect 7327 6176 7753 6184
rect 8367 6176 9153 6184
rect 10107 6176 10613 6184
rect 11067 6176 11353 6184
rect 11927 6176 12033 6184
rect 2356 6156 2484 6164
rect 2507 6156 2632 6164
rect 2667 6156 5133 6164
rect 5367 6156 5733 6164
rect 5807 6156 6333 6164
rect 6347 6156 6913 6164
rect 7027 6156 8233 6164
rect 8867 6156 8913 6164
rect 9507 6156 10073 6164
rect 10147 6156 10733 6164
rect 11027 6156 11473 6164
rect 11487 6156 11633 6164
rect 1760 6146 1784 6147
rect -24 6116 473 6124
rect 547 6116 813 6124
rect 827 6116 1033 6124
rect 1196 6104 1204 6133
rect 1767 6136 1784 6146
rect 1767 6133 1780 6136
rect 2687 6136 2913 6144
rect 3327 6136 3413 6144
rect 4047 6136 4133 6144
rect 4187 6136 4333 6144
rect 4487 6136 4733 6144
rect 4947 6136 5013 6144
rect 5847 6136 6073 6144
rect 7207 6136 7533 6144
rect 7867 6136 8073 6144
rect 8847 6136 9093 6144
rect 10867 6136 10993 6144
rect 11927 6136 12113 6144
rect 1807 6119 1893 6127
rect 2007 6119 2053 6127
rect 2107 6119 2413 6127
rect 2427 6116 2533 6124
rect 3207 6119 3253 6127
rect 3927 6119 3993 6127
rect 4687 6119 4793 6127
rect 1187 6096 1204 6104
rect 1387 6099 1473 6107
rect 1527 6096 1633 6104
rect 2767 6096 2864 6104
rect 807 6076 1113 6084
rect 1667 6076 1773 6084
rect 2856 6084 2864 6096
rect 3716 6087 3724 6116
rect 5027 6116 5073 6124
rect 5267 6116 5453 6124
rect 5647 6119 5753 6127
rect 6107 6119 6153 6127
rect 6436 6116 6453 6124
rect 6507 6119 6573 6127
rect 6647 6119 6713 6127
rect 6767 6119 6813 6127
rect 6836 6116 7053 6124
rect 7547 6126 7664 6127
rect 7547 6119 7653 6126
rect 4187 6096 4313 6104
rect 4327 6096 4893 6104
rect 5573 6104 5587 6113
rect 5573 6100 5993 6104
rect 5576 6096 5993 6100
rect 6436 6104 6444 6116
rect 6836 6104 6844 6116
rect 8407 6116 8613 6124
rect 8807 6119 8873 6127
rect 9227 6119 9393 6127
rect 9467 6116 9733 6124
rect 9787 6119 9893 6127
rect 10747 6116 10833 6124
rect 11127 6116 11144 6124
rect 11167 6116 11293 6124
rect 6176 6096 6444 6104
rect 6736 6096 6844 6104
rect 1907 6076 2073 6084
rect 2287 6073 2593 6081
rect 2856 6076 3113 6084
rect 3707 6076 3724 6087
rect 3707 6073 3720 6076
rect 3787 6073 3853 6081
rect 3947 6073 4053 6081
rect 4207 6073 4253 6081
rect 4347 6076 4513 6084
rect 4587 6076 4752 6084
rect 4787 6073 4853 6081
rect 4967 6076 5033 6084
rect 5147 6076 5333 6084
rect 6176 6084 6184 6096
rect 6736 6084 6744 6096
rect 11136 6104 11144 6116
rect 11367 6116 11673 6124
rect 10107 6096 10564 6104
rect 11136 6096 11193 6104
rect 5527 6076 5653 6084
rect 5667 6073 5853 6081
rect 6427 6073 6513 6081
rect 10556 6084 10564 6096
rect 6827 6076 7033 6084
rect 8107 6076 8333 6084
rect 8587 6073 8853 6081
rect 9907 6073 9973 6081
rect 10967 6073 11133 6081
rect 11467 6076 11553 6084
rect 11567 6073 11653 6081
rect 12127 6073 12213 6081
rect 1487 6056 1533 6064
rect 1927 6056 2833 6064
rect 3487 6056 3533 6064
rect 3627 6056 3893 6064
rect 3987 6056 4013 6064
rect 5467 6056 5873 6064
rect 6207 6056 6273 6064
rect 7287 6056 7393 6064
rect 7567 6056 7833 6064
rect 8207 6056 8373 6064
rect 9147 6056 9173 6064
rect 10527 6056 10673 6064
rect 11907 6056 12013 6064
rect 527 6036 853 6044
rect 1827 6036 2333 6044
rect 2487 6036 2753 6044
rect 3167 6036 3273 6044
rect 3367 6036 3733 6044
rect 3827 6036 4053 6044
rect 4127 6036 4653 6044
rect 4907 6036 5253 6044
rect 5347 6036 5393 6044
rect 5667 6036 5693 6044
rect 5807 6036 6033 6044
rect 6327 6036 6693 6044
rect 6987 6036 7073 6044
rect 8907 6036 9213 6044
rect 9547 6036 10093 6044
rect 10367 6036 10793 6044
rect 11107 6036 11273 6044
rect 11407 6036 11473 6044
rect 11627 6036 11773 6044
rect 11947 6036 11973 6044
rect 12067 6036 12173 6044
rect 1987 6016 2153 6024
rect 3447 6016 3493 6024
rect 3567 6016 3793 6024
rect 3936 6020 4144 6024
rect 3933 6016 4144 6020
rect 3933 6007 3947 6016
rect 267 5996 793 6004
rect 1047 5996 2113 6004
rect 2187 5996 2713 6004
rect 2787 5996 3053 6004
rect 3267 5996 3873 6004
rect 4136 6004 4144 6016
rect 5027 6016 5153 6024
rect 7167 6016 7513 6024
rect 8007 6016 8573 6024
rect 9267 6016 9753 6024
rect 10027 6016 10113 6024
rect 10307 6016 11013 6024
rect 4136 5996 4773 6004
rect 4927 5996 5213 6004
rect 5327 5996 5413 6004
rect 5647 5996 6933 6004
rect 7227 5996 7793 6004
rect 7836 5996 8633 6004
rect 1627 5976 1793 5984
rect 1907 5976 3493 5984
rect 3707 5976 3733 5984
rect 4127 5984 4140 5987
rect 4127 5973 4144 5984
rect 4267 5976 4352 5984
rect 4387 5976 4853 5984
rect 4867 5976 4933 5984
rect 5447 5976 5673 5984
rect 5767 5976 5873 5984
rect 5927 5976 6253 5984
rect 6387 5976 6633 5984
rect 7836 5984 7844 5996
rect 10476 5996 10933 6004
rect 7627 5976 7844 5984
rect 8407 5976 8793 5984
rect 10476 5984 10484 5996
rect 11667 5996 11693 6004
rect 11947 5996 12033 6004
rect 9727 5976 10484 5984
rect 10547 5976 10592 5984
rect 10627 5976 11113 5984
rect 1887 5956 4093 5964
rect 4136 5964 4144 5973
rect 4136 5956 4573 5964
rect 4707 5956 4813 5964
rect 5727 5956 5933 5964
rect 5947 5956 6032 5964
rect 6067 5956 7273 5964
rect 7927 5956 7993 5964
rect 8156 5956 9073 5964
rect -24 5936 33 5944
rect 667 5936 993 5944
rect 1007 5936 1273 5944
rect 1467 5936 1573 5944
rect 1687 5936 2933 5944
rect 3087 5936 3253 5944
rect 3327 5936 5092 5944
rect 5127 5936 5693 5944
rect 6056 5944 6064 5953
rect 8156 5947 8164 5956
rect 9887 5956 11693 5964
rect 11787 5956 12253 5964
rect 5867 5936 6064 5944
rect 7967 5936 8153 5944
rect 9247 5936 9413 5944
rect 9807 5936 9933 5944
rect 11027 5936 11193 5944
rect 11427 5936 11633 5944
rect 2727 5916 2873 5924
rect 3367 5916 4173 5924
rect 4327 5916 4393 5924
rect 4407 5916 4613 5924
rect 5887 5916 6773 5924
rect 8587 5916 8693 5924
rect 8947 5916 9113 5924
rect 10187 5916 10253 5924
rect 10267 5916 10373 5924
rect 10387 5916 10593 5924
rect 11767 5916 12013 5924
rect -24 5896 73 5904
rect 227 5899 453 5907
rect 736 5867 744 5896
rect 907 5896 1313 5904
rect 2167 5896 2393 5904
rect 2447 5899 2573 5907
rect 2707 5896 2793 5904
rect 2987 5896 3213 5904
rect 3627 5896 3793 5904
rect 3907 5899 4013 5907
rect 4287 5896 4353 5904
rect 5087 5899 5393 5907
rect 4120 5884 4133 5887
rect 4116 5873 4133 5884
rect -24 5856 52 5864
rect 87 5856 493 5864
rect 727 5856 744 5867
rect 727 5853 740 5856
rect 787 5856 1053 5864
rect 4116 5864 4124 5873
rect 4856 5884 4864 5896
rect 4447 5876 4864 5884
rect 1227 5853 1293 5861
rect 1887 5853 2133 5861
rect 2427 5853 2633 5861
rect 2807 5853 2953 5861
rect 3047 5853 3273 5861
rect 3527 5853 3613 5861
rect 3687 5853 3773 5861
rect 4047 5856 4124 5864
rect 4707 5856 5073 5864
rect 5287 5856 5353 5864
rect 5716 5864 5724 5913
rect 5907 5899 5973 5907
rect 6167 5896 6213 5904
rect 7027 5899 7313 5907
rect 7527 5899 7593 5907
rect 7827 5899 7913 5907
rect 7927 5896 8113 5904
rect 8627 5899 8653 5907
rect 8867 5899 9193 5907
rect 9587 5899 9713 5907
rect 9847 5899 9873 5907
rect 10347 5896 10493 5904
rect 6096 5864 6104 5876
rect 6367 5873 6452 5881
rect 6487 5876 6593 5884
rect 6816 5884 6824 5896
rect 10827 5899 10873 5907
rect 10927 5896 11193 5904
rect 11667 5896 11704 5904
rect 11747 5900 11924 5904
rect 11747 5896 11927 5900
rect 12207 5899 12233 5907
rect 6816 5876 6984 5884
rect 6976 5864 6984 5876
rect 9927 5876 10264 5884
rect 6027 5856 6104 5864
rect 6727 5853 6753 5861
rect 6976 5856 7093 5864
rect 7107 5853 7133 5861
rect 7367 5856 7433 5864
rect 7627 5856 7813 5864
rect 7907 5853 7953 5861
rect 8147 5856 8193 5864
rect 8347 5853 8413 5861
rect 8547 5856 8673 5864
rect 8687 5856 8953 5864
rect 9127 5853 9173 5861
rect 9527 5853 9613 5861
rect 9627 5856 9773 5864
rect 10256 5864 10264 5876
rect 9887 5856 10053 5864
rect 10256 5856 10313 5864
rect 10647 5856 10813 5864
rect 11447 5853 11533 5861
rect 11696 5847 11704 5896
rect 11913 5887 11927 5896
rect 11767 5856 11873 5864
rect 1587 5836 1693 5844
rect 2307 5836 2713 5844
rect 2976 5836 3244 5844
rect 27 5816 253 5824
rect 1767 5816 2173 5824
rect 2567 5816 2693 5824
rect 2747 5816 2793 5824
rect 2976 5824 2984 5836
rect 2807 5816 2984 5824
rect 3187 5816 3213 5824
rect 3236 5824 3244 5836
rect 3296 5836 3824 5844
rect 3296 5824 3304 5836
rect 3816 5827 3824 5836
rect 4587 5836 4713 5844
rect 4787 5836 4853 5844
rect 4907 5836 5133 5844
rect 6067 5836 6113 5844
rect 3236 5816 3304 5824
rect 3827 5816 4053 5824
rect 4267 5816 4313 5824
rect 5407 5816 5473 5824
rect 5627 5816 5893 5824
rect 6213 5824 6227 5833
rect 6527 5833 6673 5841
rect 6687 5833 6753 5841
rect 8727 5836 10193 5844
rect 10547 5836 10613 5844
rect 11207 5836 11253 5844
rect 12047 5836 12253 5844
rect 6167 5820 6227 5824
rect 6167 5816 6224 5820
rect 7247 5816 7412 5824
rect 7447 5816 8693 5824
rect 8887 5816 9053 5824
rect 9287 5816 9533 5824
rect 9627 5816 10133 5824
rect 10907 5816 10993 5824
rect 67 5796 772 5804
rect 807 5796 1673 5804
rect 2207 5796 3133 5804
rect 3567 5796 4073 5804
rect 4607 5796 4744 5804
rect 47 5776 993 5784
rect 1067 5776 1853 5784
rect 1967 5776 2273 5784
rect 2327 5776 2673 5784
rect 2907 5776 3053 5784
rect 3667 5776 3993 5784
rect 4736 5784 4744 5796
rect 4767 5796 4873 5804
rect 5727 5796 5833 5804
rect 6067 5796 6553 5804
rect 7387 5796 8473 5804
rect 8787 5796 9213 5804
rect 9587 5796 9953 5804
rect 10427 5796 10573 5804
rect 11187 5796 11473 5804
rect 11647 5796 11913 5804
rect 11927 5796 12193 5804
rect 4736 5776 5173 5784
rect 5387 5776 5413 5784
rect 5507 5776 6733 5784
rect 6807 5776 7193 5784
rect 7707 5776 7844 5784
rect 1407 5756 1713 5764
rect 2867 5756 3553 5764
rect 3807 5756 3913 5764
rect 3967 5756 4213 5764
rect 4467 5756 4593 5764
rect 5107 5756 5473 5764
rect 5567 5756 5993 5764
rect 6147 5756 6713 5764
rect 6767 5756 7353 5764
rect 7836 5764 7844 5776
rect 7987 5776 8713 5784
rect 11627 5776 11713 5784
rect 7427 5756 7824 5764
rect 7836 5756 8633 5764
rect 1267 5736 1673 5744
rect 2467 5736 3353 5744
rect 3367 5736 3393 5744
rect 5107 5736 5333 5744
rect 5747 5736 5813 5744
rect 6747 5736 7673 5744
rect 7816 5744 7824 5756
rect 8827 5756 10013 5764
rect 12007 5756 12253 5764
rect 7816 5736 8393 5744
rect 8667 5736 8753 5744
rect 10047 5736 10093 5744
rect 10107 5736 10253 5744
rect 11227 5736 11333 5744
rect 947 5716 1333 5724
rect 1807 5716 2173 5724
rect 2587 5716 3073 5724
rect 3167 5716 3193 5724
rect 3207 5716 4673 5724
rect 4687 5716 6173 5724
rect 6287 5716 7013 5724
rect 7067 5716 7193 5724
rect 7207 5716 7372 5724
rect 7407 5716 7773 5724
rect 8187 5716 8373 5724
rect 9527 5716 11773 5724
rect 727 5696 1253 5704
rect 1687 5696 2453 5704
rect 3287 5696 4173 5704
rect 4267 5696 4693 5704
rect 5087 5696 5373 5704
rect 5787 5696 6113 5704
rect 6707 5696 7113 5704
rect 8407 5696 10093 5704
rect 11307 5696 11673 5704
rect 11687 5696 11733 5704
rect 1667 5676 2313 5684
rect 2367 5676 2673 5684
rect 2827 5676 3253 5684
rect 3427 5676 3873 5684
rect 4227 5676 5013 5684
rect 5027 5676 5553 5684
rect 5607 5676 7413 5684
rect 7747 5676 8173 5684
rect 8907 5676 9553 5684
rect 10507 5676 11273 5684
rect 11507 5676 11593 5684
rect 827 5656 3773 5664
rect 3907 5656 4073 5664
rect 4307 5656 5033 5664
rect 5047 5656 5433 5664
rect 5907 5656 6273 5664
rect 7267 5656 7353 5664
rect 7627 5656 8244 5664
rect -24 5624 -16 5644
rect 27 5636 753 5644
rect 847 5636 1913 5644
rect 2007 5636 2133 5644
rect 2187 5636 2853 5644
rect 2967 5636 3313 5644
rect 3487 5636 3533 5644
rect 3887 5636 4253 5644
rect 4647 5636 4733 5644
rect 5307 5636 5473 5644
rect 5487 5636 5533 5644
rect 6307 5636 6893 5644
rect 7887 5636 8213 5644
rect 8236 5644 8244 5656
rect 8327 5656 8733 5664
rect 11887 5656 12033 5664
rect 8236 5636 8333 5644
rect 8707 5636 8893 5644
rect 10467 5636 10773 5644
rect 11327 5636 11413 5644
rect 11527 5636 11633 5644
rect 11687 5636 11893 5644
rect -44 5616 -16 5624
rect -44 5584 -36 5616
rect 1087 5616 1673 5624
rect 1807 5616 2033 5624
rect 2047 5616 2393 5624
rect 2407 5616 2793 5624
rect 3307 5616 4293 5624
rect 4407 5616 4773 5624
rect 4787 5616 5153 5624
rect 5387 5616 5593 5624
rect 5707 5616 5793 5624
rect 7567 5616 7833 5624
rect 8947 5616 8973 5624
rect 9727 5616 10033 5624
rect -24 5596 13 5604
rect 36 5596 213 5604
rect 36 5584 44 5596
rect 687 5596 993 5604
rect 1307 5599 1353 5607
rect 1567 5599 1633 5607
rect 2107 5599 2173 5607
rect 2687 5599 2773 5607
rect 2927 5599 3093 5607
rect 3247 5599 3273 5607
rect 3296 5596 3513 5604
rect -44 5576 44 5584
rect 1687 5576 2213 5584
rect 3296 5584 3304 5596
rect 3647 5596 3973 5604
rect 4027 5596 4253 5604
rect 4487 5596 4684 5604
rect 4707 5599 4733 5607
rect 5007 5599 5173 5607
rect 3087 5576 3304 5584
rect 4676 5584 4684 5596
rect 5187 5599 5313 5607
rect 5367 5596 5533 5604
rect 5827 5599 5873 5607
rect 5987 5596 6053 5604
rect 6687 5599 6833 5607
rect 7327 5596 7673 5604
rect 7687 5596 7913 5604
rect 8087 5599 8133 5607
rect 8267 5599 8453 5607
rect 8467 5596 8573 5604
rect 8747 5599 8793 5607
rect 8807 5596 9013 5604
rect 9316 5596 9513 5604
rect 9316 5590 9324 5596
rect 9787 5599 9993 5607
rect 10067 5596 10113 5604
rect 10127 5596 10213 5604
rect 10227 5596 10253 5604
rect 10747 5596 10804 5604
rect 10827 5599 11013 5607
rect 11087 5599 11153 5607
rect 4676 5576 4913 5584
rect 5607 5576 6353 5584
rect 10796 5584 10804 5596
rect 9447 5573 9653 5581
rect 10796 5576 10873 5584
rect 667 5556 733 5564
rect 1047 5553 1073 5561
rect 1087 5556 1133 5564
rect 1207 5556 1273 5564
rect 1827 5556 1873 5564
rect 1927 5556 2073 5564
rect 2267 5556 2373 5564
rect 2467 5556 2613 5564
rect 2707 5560 2984 5564
rect 2707 5556 2987 5560
rect 2973 5547 2987 5556
rect 3067 5556 3213 5564
rect 3327 5553 3433 5561
rect 3447 5553 3493 5561
rect 3727 5553 3833 5561
rect 4007 5553 4073 5561
rect 4287 5556 4513 5564
rect 4667 5556 4753 5564
rect 4807 5556 4832 5564
rect 4867 5556 5013 5564
rect 5027 5553 5073 5561
rect 5847 5556 5913 5564
rect 5927 5556 6073 5564
rect 6587 5556 6753 5564
rect 7867 5553 7993 5561
rect 8447 5556 8533 5564
rect 8727 5556 8853 5564
rect 10796 5564 10804 5576
rect 9767 5553 9793 5561
rect 10027 5553 10113 5561
rect 10547 5556 10753 5564
rect 11107 5553 11293 5561
rect 11316 5547 11324 5596
rect 11527 5596 11573 5604
rect 11787 5596 11853 5604
rect 11347 5556 11613 5564
rect 11916 5563 11924 5593
rect 11953 5584 11967 5593
rect 11953 5580 12013 5584
rect 11956 5576 12013 5580
rect 12196 5567 12204 5596
rect 12196 5556 12212 5567
rect 12200 5553 12212 5556
rect 12247 5553 12273 5561
rect 1247 5543 1284 5544
rect 1247 5536 1273 5543
rect 1587 5536 2653 5544
rect 3127 5543 3224 5544
rect 3127 5536 3213 5543
rect 5547 5536 5733 5544
rect 6187 5536 6553 5544
rect 6827 5536 6893 5544
rect 7367 5536 7684 5544
rect 267 5516 833 5524
rect 1627 5516 2933 5524
rect 3467 5516 3633 5524
rect 4107 5516 4253 5524
rect 4307 5516 4933 5524
rect 6327 5516 6793 5524
rect 7676 5524 7684 5536
rect 7876 5536 8253 5544
rect 7876 5524 7884 5536
rect 8747 5536 8824 5544
rect 7676 5516 7884 5524
rect 8627 5516 8713 5524
rect 8816 5524 8824 5536
rect 8907 5536 8993 5544
rect 9067 5536 9973 5544
rect 8816 5516 9953 5524
rect 10107 5516 10273 5524
rect 10287 5516 10633 5524
rect 10727 5516 11053 5524
rect 11627 5516 11973 5524
rect 12227 5516 12293 5524
rect 427 5496 633 5504
rect 647 5496 773 5504
rect 1327 5496 1533 5504
rect 1647 5496 2073 5504
rect 2227 5496 3073 5504
rect 3367 5496 4073 5504
rect 4147 5496 4233 5504
rect 4707 5496 4993 5504
rect 7667 5496 7993 5504
rect 8007 5496 8113 5504
rect 8167 5496 8793 5504
rect 8967 5496 9553 5504
rect 11167 5496 11393 5504
rect 1316 5484 1324 5493
rect 507 5476 1324 5484
rect 1676 5476 2033 5484
rect 1676 5464 1684 5476
rect 2127 5476 2893 5484
rect 2947 5476 3064 5484
rect 1447 5456 1684 5464
rect 1727 5456 2573 5464
rect 3056 5464 3064 5476
rect 3427 5476 3473 5484
rect 3587 5476 3812 5484
rect 3847 5476 4333 5484
rect 5067 5476 5193 5484
rect 5287 5476 5533 5484
rect 5627 5476 6193 5484
rect 6207 5476 6273 5484
rect 6287 5476 6433 5484
rect 6787 5476 7213 5484
rect 7767 5476 7893 5484
rect 8667 5476 8753 5484
rect 8827 5476 9313 5484
rect 9387 5476 9673 5484
rect 9747 5476 10513 5484
rect 11687 5476 11933 5484
rect 11987 5476 12013 5484
rect 3056 5456 3344 5464
rect 507 5436 813 5444
rect 1747 5436 3033 5444
rect 3336 5444 3344 5456
rect 3387 5456 3833 5464
rect 4067 5456 4493 5464
rect 4667 5456 5013 5464
rect 5027 5456 5233 5464
rect 5756 5456 5893 5464
rect 3336 5436 3453 5444
rect 3827 5436 4473 5444
rect 4627 5436 5053 5444
rect 5756 5444 5764 5456
rect 8387 5456 9653 5464
rect 5327 5436 5764 5444
rect 6227 5436 6573 5444
rect 6587 5436 6633 5444
rect 7367 5436 7693 5444
rect 8227 5436 9873 5444
rect 9887 5436 10853 5444
rect 10947 5436 11873 5444
rect 767 5416 1713 5424
rect 1867 5416 2473 5424
rect 2687 5416 2793 5424
rect 2807 5416 2832 5424
rect 2867 5416 2893 5424
rect 2916 5416 3313 5424
rect 1307 5396 1453 5404
rect 2916 5404 2924 5416
rect 3327 5416 3573 5424
rect 3867 5416 4113 5424
rect 4247 5416 4373 5424
rect 4547 5416 5133 5424
rect 5227 5416 6133 5424
rect 7587 5416 7733 5424
rect 7747 5416 7853 5424
rect 8647 5416 8833 5424
rect 8947 5416 9173 5424
rect 9367 5416 9533 5424
rect 10287 5416 10833 5424
rect 11947 5416 12013 5424
rect 2467 5396 2924 5404
rect 4187 5396 4433 5404
rect 4447 5396 4473 5404
rect 5087 5396 5793 5404
rect 7687 5396 7733 5404
rect 7747 5396 8093 5404
rect 8107 5396 8273 5404
rect 8287 5396 8533 5404
rect 8547 5396 8913 5404
rect 11047 5396 11293 5404
rect 11767 5396 11993 5404
rect 1547 5376 1733 5384
rect 1747 5379 1833 5387
rect 2047 5376 2193 5384
rect 2547 5376 2613 5384
rect 2667 5376 2933 5384
rect 3027 5376 3153 5384
rect 3267 5376 3573 5384
rect 3587 5379 3673 5387
rect 3827 5379 3893 5387
rect 3947 5376 4013 5384
rect 4087 5379 4153 5387
rect 4207 5376 4273 5384
rect 4507 5376 5253 5384
rect 5567 5376 5693 5384
rect 5987 5376 6293 5384
rect 6627 5379 6653 5387
rect 6927 5380 6953 5388
rect 7027 5387 7093 5388
rect 7027 5380 7073 5387
rect 7087 5380 7093 5387
rect 7116 5376 7313 5384
rect 7627 5376 7924 5384
rect 7947 5379 8133 5387
rect 8187 5379 8213 5387
rect 8667 5376 8813 5384
rect -24 5336 193 5344
rect 696 5344 704 5373
rect 987 5353 1193 5361
rect 1247 5359 1333 5367
rect 2327 5353 2453 5361
rect 2527 5356 2633 5364
rect 3207 5356 3733 5364
rect 4176 5356 4393 5364
rect 307 5336 473 5344
rect 696 5336 713 5344
rect 1767 5333 1853 5341
rect 1967 5336 2013 5344
rect 2067 5336 2813 5344
rect 2827 5333 2973 5341
rect 3327 5336 3373 5344
rect 3667 5333 3713 5341
rect 4176 5344 4184 5356
rect 4527 5356 5213 5364
rect 7116 5364 7124 5376
rect 6996 5356 7124 5364
rect 7916 5364 7924 5376
rect 9107 5379 9213 5387
rect 9407 5379 9433 5387
rect 9607 5379 9693 5387
rect 7916 5356 8373 5364
rect 4047 5336 4173 5344
rect 4187 5336 4233 5344
rect 4467 5336 4653 5344
rect 5347 5333 5433 5341
rect 5447 5333 5593 5341
rect 5687 5333 5733 5341
rect 5887 5336 5953 5344
rect 6127 5336 6193 5344
rect 6467 5336 6713 5344
rect 6727 5333 6753 5341
rect 6996 5345 7004 5356
rect 6807 5336 6993 5344
rect 7916 5344 7924 5356
rect 8896 5364 8904 5376
rect 9947 5376 10033 5384
rect 10047 5379 10093 5387
rect 10567 5379 10593 5387
rect 10787 5376 10812 5384
rect 10847 5379 11033 5387
rect 11547 5380 11573 5388
rect 8896 5356 8993 5364
rect 7807 5333 7873 5341
rect 8507 5336 8533 5344
rect 8547 5333 8633 5341
rect 8867 5333 8913 5341
rect 9487 5336 9593 5344
rect 9667 5333 9753 5341
rect 10307 5333 10393 5341
rect 11096 5344 11104 5373
rect 11316 5347 11324 5373
rect 12236 5347 12244 5376
rect 12276 5347 12284 5373
rect 10467 5336 10533 5344
rect 11067 5336 11104 5344
rect 11207 5336 11253 5344
rect 11687 5336 11713 5344
rect 11887 5333 11913 5341
rect 11967 5333 12053 5341
rect 12227 5336 12244 5347
rect 12227 5333 12240 5336
rect 647 5316 673 5324
rect 687 5316 773 5324
rect 1387 5316 1453 5324
rect 2467 5316 2493 5324
rect 2867 5316 2933 5324
rect 3807 5316 3833 5324
rect 4887 5316 5053 5324
rect 7067 5316 7453 5324
rect 7527 5316 8444 5324
rect 1487 5296 2053 5304
rect 3087 5300 3724 5304
rect 3087 5296 3727 5300
rect 3713 5287 3727 5296
rect 4327 5296 4513 5304
rect 4647 5296 4693 5304
rect 5056 5304 5064 5313
rect 5056 5296 5453 5304
rect 5647 5296 6013 5304
rect 7107 5296 7313 5304
rect 7327 5304 7340 5307
rect 7327 5296 7344 5304
rect 7327 5293 7340 5296
rect 7587 5296 7633 5304
rect 7867 5296 8153 5304
rect 8227 5296 8413 5304
rect 8436 5304 8444 5316
rect 8827 5316 8953 5324
rect 10027 5316 10173 5324
rect 11347 5316 11613 5324
rect 12127 5316 12153 5324
rect 8436 5296 9173 5304
rect 9187 5296 9573 5304
rect 9747 5296 9793 5304
rect 10547 5296 10593 5304
rect 10767 5296 10813 5304
rect 10947 5296 11273 5304
rect 407 5276 1433 5284
rect 1527 5276 1753 5284
rect 3187 5276 3613 5284
rect 3787 5276 4013 5284
rect 4027 5276 4393 5284
rect 6036 5276 6313 5284
rect 1807 5256 2333 5264
rect 2987 5256 3633 5264
rect 4807 5256 5033 5264
rect 6036 5264 6044 5276
rect 6687 5276 7373 5284
rect 7707 5276 8153 5284
rect 9207 5276 10253 5284
rect 10647 5276 10833 5284
rect 11047 5276 11153 5284
rect 11327 5276 12273 5284
rect 5927 5256 6044 5264
rect 7647 5256 8673 5264
rect 8827 5256 9013 5264
rect 10107 5256 10273 5264
rect 10287 5256 10353 5264
rect 827 5236 953 5244
rect 1547 5236 1812 5244
rect 1847 5236 1944 5244
rect 1936 5224 1944 5236
rect 2007 5236 2153 5244
rect 2827 5236 3133 5244
rect 3147 5236 3233 5244
rect 3247 5236 3653 5244
rect 3747 5236 4093 5244
rect 4847 5236 5273 5244
rect 5487 5236 5673 5244
rect 5687 5236 6133 5244
rect 7367 5236 7393 5244
rect 7907 5236 8732 5244
rect 8767 5236 9393 5244
rect 9407 5236 9433 5244
rect 9727 5236 9993 5244
rect 10047 5236 10453 5244
rect 12187 5236 12273 5244
rect 1936 5216 2113 5224
rect 2427 5216 2673 5224
rect 3407 5216 4053 5224
rect 4167 5216 4913 5224
rect 5167 5216 5413 5224
rect 5427 5216 5653 5224
rect 5667 5216 8804 5224
rect 8796 5207 8804 5216
rect 9467 5216 9633 5224
rect 10487 5216 11293 5224
rect 1707 5196 2133 5204
rect 2287 5196 2473 5204
rect 2487 5196 2813 5204
rect 3107 5196 3513 5204
rect 3707 5196 3913 5204
rect 4107 5196 4352 5204
rect 4387 5196 4904 5204
rect 1387 5176 1613 5184
rect 2107 5176 2513 5184
rect 2807 5176 3393 5184
rect 4896 5184 4904 5196
rect 5387 5196 5693 5204
rect 5707 5196 7273 5204
rect 7287 5196 8553 5204
rect 8567 5196 8753 5204
rect 8807 5196 9813 5204
rect 9867 5196 10293 5204
rect 12087 5196 12293 5204
rect 4896 5176 4973 5184
rect 7227 5176 7593 5184
rect 8076 5176 8473 5184
rect 8076 5167 8084 5176
rect 8767 5176 10032 5184
rect 10067 5176 11453 5184
rect 1027 5156 1593 5164
rect 1947 5156 2093 5164
rect 2747 5164 2760 5167
rect 2747 5153 2764 5164
rect 3427 5156 3473 5164
rect 3547 5156 3593 5164
rect 5327 5156 5713 5164
rect 5987 5156 6333 5164
rect 7456 5156 8073 5164
rect 2756 5144 2764 5153
rect 7456 5147 7464 5156
rect 8567 5156 8713 5164
rect 9007 5156 9473 5164
rect 9567 5156 10113 5164
rect 10207 5156 10513 5164
rect 11707 5156 11913 5164
rect 2756 5136 2953 5144
rect 5207 5136 5293 5144
rect 6667 5136 7293 5144
rect 7307 5136 7453 5144
rect 8167 5136 8533 5144
rect 9027 5136 9853 5144
rect 11007 5136 11633 5144
rect 1207 5116 1313 5124
rect 1447 5116 1493 5124
rect 1627 5116 1744 5124
rect 627 5096 653 5104
rect 967 5096 993 5104
rect 1007 5096 1573 5104
rect -24 5076 193 5084
rect 307 5076 473 5084
rect 1247 5079 1313 5087
rect 807 5059 1013 5067
rect 467 5036 653 5044
rect 1227 5036 1373 5044
rect 1456 5044 1464 5073
rect 1736 5070 1744 5116
rect 2047 5116 2633 5124
rect 2647 5116 2733 5124
rect 3267 5116 3433 5124
rect 4147 5116 4213 5124
rect 4567 5120 4624 5124
rect 4567 5116 4627 5120
rect 4613 5107 4627 5116
rect 4927 5116 5813 5124
rect 6207 5116 6733 5124
rect 7367 5116 7733 5124
rect 8087 5116 9253 5124
rect 9687 5116 9993 5124
rect 10507 5116 10953 5124
rect 11747 5116 11932 5124
rect 11967 5116 12033 5124
rect 2807 5096 2913 5104
rect 2927 5096 3053 5104
rect 3107 5096 3453 5104
rect 3687 5096 3724 5104
rect 2207 5076 2233 5084
rect 2447 5076 2493 5084
rect 2847 5079 2873 5087
rect 3147 5079 3292 5087
rect 3327 5079 3373 5087
rect 2576 5064 2584 5076
rect 3607 5076 3644 5084
rect 1947 5053 2033 5061
rect 2576 5056 2624 5064
rect 1456 5036 1553 5044
rect 2616 5044 2624 5056
rect 2967 5056 3193 5064
rect 2167 5036 2253 5044
rect 2547 5033 2593 5041
rect 2616 5036 2813 5044
rect 2867 5036 3393 5044
rect 3636 5027 3644 5076
rect 3696 5044 3704 5073
rect 3716 5064 3724 5096
rect 3767 5096 3853 5104
rect 4327 5096 4413 5104
rect 4520 5104 4533 5107
rect 4516 5093 4533 5104
rect 5127 5096 5173 5104
rect 6127 5096 6153 5104
rect 9607 5096 10193 5104
rect 11087 5096 11133 5104
rect 3996 5076 4293 5084
rect 3996 5070 4004 5076
rect 4516 5084 4524 5093
rect 4496 5076 4524 5084
rect 3716 5056 3753 5064
rect 4187 5056 4273 5064
rect 4436 5047 4444 5076
rect 4496 5067 4504 5076
rect 4487 5056 4504 5067
rect 4487 5053 4500 5056
rect 4576 5064 4584 5093
rect 4547 5056 4584 5064
rect 4627 5059 4753 5067
rect 4896 5064 4904 5093
rect 5087 5076 5193 5084
rect 5207 5079 5313 5087
rect 5467 5079 5493 5087
rect 6527 5076 6613 5084
rect 6627 5076 6653 5084
rect 6807 5076 7033 5084
rect 7087 5079 7213 5087
rect 8287 5079 8393 5087
rect 8447 5079 8593 5087
rect 4867 5056 4904 5064
rect 3667 5036 3704 5044
rect 4307 5036 4413 5044
rect 4436 5036 4453 5047
rect 4440 5033 4453 5036
rect 5736 5044 5744 5073
rect 5773 5064 5787 5073
rect 5773 5060 5853 5064
rect 5776 5056 5853 5060
rect 5987 5059 6133 5067
rect 8156 5064 8164 5076
rect 8607 5079 8613 5087
rect 9007 5079 9033 5087
rect 9227 5076 9413 5084
rect 9427 5079 9513 5087
rect 9707 5079 9833 5087
rect 8116 5056 8253 5064
rect 8116 5047 8124 5056
rect 8696 5064 8704 5076
rect 8696 5056 8893 5064
rect 5067 5036 5153 5044
rect 5736 5036 5753 5044
rect 7227 5036 7313 5044
rect 7467 5033 7553 5041
rect 7847 5036 8072 5044
rect 8107 5036 8124 5047
rect 8107 5033 8120 5036
rect 8147 5036 8273 5044
rect 8467 5033 8493 5041
rect 8727 5036 8753 5044
rect 8956 5044 8964 5076
rect 9556 5064 9564 5076
rect 10047 5076 10333 5084
rect 10407 5086 10444 5087
rect 10407 5079 10433 5086
rect 10727 5076 10873 5084
rect 10947 5079 10993 5087
rect 11187 5079 11213 5087
rect 11367 5076 11413 5084
rect 11607 5079 11693 5087
rect 11747 5079 11873 5087
rect 12067 5079 12113 5087
rect 9556 5056 9633 5064
rect 9776 5056 9953 5064
rect 8927 5036 8964 5044
rect 8987 5036 9093 5044
rect 9287 5036 9373 5044
rect 9547 5036 9673 5044
rect 9776 5044 9784 5056
rect 10007 5056 10493 5064
rect 11287 5056 11333 5064
rect 11496 5047 11504 5075
rect 12127 5079 12193 5087
rect 9827 5033 9873 5041
rect 10647 5033 10713 5041
rect 11207 5036 11233 5044
rect 11496 5036 11513 5047
rect 11500 5033 11513 5036
rect 11567 5036 11753 5044
rect 11927 5033 12033 5041
rect 12047 5036 12213 5044
rect 2007 5016 2373 5024
rect 2947 5016 3073 5024
rect 3087 5024 3100 5027
rect 3087 5016 3104 5024
rect 3216 5016 3613 5024
rect 3087 5013 3100 5016
rect 247 4996 433 5004
rect 1447 4996 1933 5004
rect 2587 4996 2672 5004
rect 3216 5004 3224 5016
rect 3636 5024 3660 5027
rect 3636 5023 3664 5024
rect 3636 5016 3653 5023
rect 3640 5013 3653 5016
rect 3707 5016 3853 5024
rect 4527 5016 4613 5024
rect 5247 5016 5433 5024
rect 5647 5016 5713 5024
rect 5836 5016 6133 5024
rect 2707 4996 3224 5004
rect 3247 4996 3713 5004
rect 3787 4996 4193 5004
rect 4327 4996 4493 5004
rect 5836 5004 5844 5016
rect 6767 5016 7133 5024
rect 8547 5016 8813 5024
rect 9127 5016 9253 5024
rect 10447 5016 10473 5024
rect 11067 5016 11133 5024
rect 11407 5016 11433 5024
rect 5747 4996 5844 5004
rect 6827 4996 7013 5004
rect 7287 4996 7773 5004
rect 7787 4996 7993 5004
rect 8067 4996 8233 5004
rect 8427 4996 8513 5004
rect 9047 4996 9593 5004
rect 9787 4996 9893 5004
rect 11167 4996 11253 5004
rect 11847 4996 12053 5004
rect 627 4976 1133 4984
rect 1427 4976 1493 4984
rect 5047 4976 5173 4984
rect 5367 4976 5853 4984
rect 6147 4976 6173 4984
rect 6267 4976 7213 4984
rect 8447 4976 8673 4984
rect 8687 4976 8773 4984
rect 8847 4976 8944 4984
rect 507 4956 673 4964
rect 1327 4956 1653 4964
rect 2127 4956 2293 4964
rect 2307 4956 3013 4964
rect 3467 4956 3813 4964
rect 4047 4956 4213 4964
rect 4287 4956 4473 4964
rect 4867 4956 4993 4964
rect 5627 4956 5773 4964
rect 6147 4956 6333 4964
rect 6787 4956 7433 4964
rect 7447 4956 7493 4964
rect 8167 4956 8813 4964
rect 8936 4964 8944 4976
rect 9107 4976 9533 4984
rect 9967 4976 10913 4984
rect 11487 4976 11573 4984
rect 8936 4956 9273 4964
rect 9407 4956 9893 4964
rect 11047 4956 11153 4964
rect 11767 4956 11873 4964
rect 12047 4956 12153 4964
rect 867 4936 1173 4944
rect 1187 4936 1273 4944
rect 1407 4936 1573 4944
rect 1787 4936 2213 4944
rect 3167 4936 3253 4944
rect 3587 4936 3933 4944
rect 4087 4936 4173 4944
rect 4507 4936 4573 4944
rect 5327 4936 5453 4944
rect 5507 4936 5913 4944
rect 7047 4936 7173 4944
rect 7267 4936 7393 4944
rect 7727 4936 7973 4944
rect 7987 4936 8513 4944
rect 8607 4936 8853 4944
rect 8927 4936 9553 4944
rect 10087 4936 10753 4944
rect 11227 4936 11593 4944
rect 11647 4936 11993 4944
rect 1887 4916 1973 4924
rect 2747 4916 2933 4924
rect 3127 4916 3533 4924
rect 3807 4916 4553 4924
rect 4707 4916 5073 4924
rect 5987 4916 6773 4924
rect 6787 4916 6913 4924
rect 7467 4916 9393 4924
rect 9907 4916 10733 4924
rect 827 4896 1013 4904
rect 1067 4896 1473 4904
rect 1847 4896 2133 4904
rect 2187 4896 2353 4904
rect 2687 4896 2993 4904
rect 3327 4896 3613 4904
rect 4107 4896 4233 4904
rect 5247 4896 5273 4904
rect 5587 4896 5693 4904
rect 5707 4896 5813 4904
rect 5967 4896 6233 4904
rect 6387 4896 6693 4904
rect 7067 4896 7873 4904
rect 8587 4896 8724 4904
rect 1627 4876 1733 4884
rect 2207 4876 2293 4884
rect 2647 4876 2753 4884
rect 3947 4876 3993 4884
rect 4407 4876 4733 4884
rect 4847 4876 5013 4884
rect 5127 4876 5153 4884
rect 5507 4876 5553 4884
rect 5947 4876 6133 4884
rect 7227 4876 7413 4884
rect 7507 4876 7573 4884
rect 8716 4884 8724 4896
rect 8827 4896 9093 4904
rect 9427 4896 9833 4904
rect 10407 4896 10593 4904
rect 11047 4896 11393 4904
rect 8716 4876 8793 4884
rect 9127 4876 9173 4884
rect 10227 4876 10253 4884
rect 10747 4876 10953 4884
rect 207 4859 293 4867
rect 307 4856 413 4864
rect 907 4856 1093 4864
rect 1147 4856 1253 4864
rect 1267 4859 1333 4867
rect 1347 4856 1593 4864
rect 2536 4856 2773 4864
rect 2827 4859 2853 4867
rect 3007 4859 3053 4867
rect 2496 4827 2504 4856
rect -24 4816 213 4824
rect 267 4816 493 4824
rect 567 4813 633 4821
rect 687 4816 833 4824
rect 847 4813 1033 4821
rect 1967 4813 2073 4821
rect 2087 4816 2193 4824
rect 2496 4816 2512 4827
rect 2500 4813 2512 4816
rect 2536 4824 2544 4856
rect 3147 4856 3333 4864
rect 3907 4856 3973 4864
rect 4027 4856 4133 4864
rect 3427 4836 3773 4844
rect 2607 4816 2853 4824
rect 3327 4813 3473 4821
rect 4176 4824 4184 4856
rect 4987 4856 5033 4864
rect 5087 4866 5124 4867
rect 5087 4859 5113 4866
rect 5347 4856 5393 4864
rect 5447 4856 5573 4864
rect 6627 4859 6713 4867
rect 6827 4859 6853 4867
rect 6907 4859 6973 4867
rect 7107 4856 7153 4864
rect 7647 4859 7693 4867
rect 8287 4866 8364 4867
rect 8287 4859 8353 4866
rect 8567 4859 8693 4867
rect 8847 4859 8933 4867
rect 8987 4856 9073 4864
rect 9247 4856 9393 4864
rect 9407 4859 9513 4867
rect 9587 4859 9673 4867
rect 9687 4856 9873 4864
rect 9927 4856 10393 4864
rect 10456 4856 10513 4864
rect 5016 4836 5153 4844
rect 4147 4816 4184 4824
rect 4367 4816 4413 4824
rect 4436 4820 4913 4824
rect 4433 4816 4913 4820
rect 4433 4807 4447 4816
rect 5016 4824 5024 4836
rect 5387 4816 5553 4824
rect 5667 4813 5833 4821
rect 5887 4813 6033 4821
rect 6247 4813 6313 4821
rect 6327 4813 6393 4821
rect 6587 4816 6633 4824
rect 6647 4816 6813 4824
rect 7027 4813 7133 4821
rect 7187 4813 7213 4821
rect 7327 4813 7433 4821
rect 7727 4816 7753 4824
rect 8787 4813 8853 4821
rect 10456 4824 10464 4856
rect 10567 4859 10713 4867
rect 10767 4856 10913 4864
rect 11087 4856 11113 4864
rect 11387 4856 11553 4864
rect 11667 4856 11893 4864
rect 11947 4859 12013 4867
rect 12027 4859 12153 4867
rect 8947 4816 9053 4824
rect 9327 4813 9373 4821
rect 9567 4813 9613 4821
rect 10507 4813 10593 4821
rect 10927 4813 11013 4821
rect 11316 4824 11324 4853
rect 11307 4816 11324 4824
rect 11527 4816 11633 4824
rect 12067 4816 12113 4824
rect 12127 4813 12173 4821
rect 12247 4816 12273 4824
rect 1407 4796 1433 4804
rect 1447 4796 1653 4804
rect 2947 4796 3013 4804
rect 3207 4796 3593 4804
rect 3767 4796 4153 4804
rect 4207 4796 4253 4804
rect 4567 4796 4773 4804
rect 5327 4796 5433 4804
rect 7807 4796 7973 4804
rect 7987 4796 8153 4804
rect 8387 4796 8553 4804
rect 8567 4796 8913 4804
rect 9127 4796 9193 4804
rect 9487 4796 9933 4804
rect 9947 4796 10153 4804
rect 10167 4796 10373 4804
rect 11367 4796 11433 4804
rect 11527 4796 11873 4804
rect 467 4776 573 4784
rect 807 4776 893 4784
rect 1687 4776 2013 4784
rect 2247 4776 3033 4784
rect 3227 4776 3413 4784
rect 3467 4776 3873 4784
rect 3987 4776 4233 4784
rect 4467 4776 4533 4784
rect 4927 4776 5093 4784
rect 5507 4776 5593 4784
rect 6087 4776 6113 4784
rect 6127 4776 6173 4784
rect 6976 4776 7073 4784
rect 1127 4756 1353 4764
rect 1367 4756 1633 4764
rect 1927 4756 2473 4764
rect 2767 4756 2953 4764
rect 3187 4756 3313 4764
rect 3647 4756 3733 4764
rect 3867 4756 3913 4764
rect 4307 4756 4733 4764
rect 5187 4756 5593 4764
rect 5787 4756 6173 4764
rect 6267 4756 6433 4764
rect 6976 4764 6984 4776
rect 7967 4776 8213 4784
rect 8467 4776 8513 4784
rect 8627 4776 8753 4784
rect 8767 4776 8793 4784
rect 8847 4776 8873 4784
rect 9067 4776 9233 4784
rect 9307 4776 9373 4784
rect 9927 4776 9973 4784
rect 10207 4776 10293 4784
rect 10687 4776 10773 4784
rect 10787 4776 11493 4784
rect 12047 4776 12173 4784
rect 6487 4756 6984 4764
rect 7107 4756 7473 4764
rect 7627 4756 8533 4764
rect 8547 4756 8933 4764
rect 9047 4756 9193 4764
rect 9207 4756 9473 4764
rect 10527 4756 10913 4764
rect 10967 4756 11333 4764
rect 11947 4756 12213 4764
rect 587 4736 1513 4744
rect 1667 4736 2733 4744
rect 2947 4736 3453 4744
rect 3547 4736 3753 4744
rect 3867 4736 4313 4744
rect 5667 4736 5993 4744
rect 6007 4736 7093 4744
rect 8127 4736 8253 4744
rect 8507 4736 8813 4744
rect 8907 4736 9353 4744
rect 9447 4736 10433 4744
rect 10727 4736 10813 4744
rect 10947 4736 11033 4744
rect 1307 4716 1553 4724
rect 2107 4716 2313 4724
rect 2487 4716 2753 4724
rect 2807 4716 2873 4724
rect 2887 4716 3353 4724
rect 3367 4716 3413 4724
rect 3427 4716 4724 4724
rect 4716 4707 4724 4716
rect 4787 4716 4913 4724
rect 5067 4716 6213 4724
rect 6347 4716 7273 4724
rect 7607 4716 8873 4724
rect 9027 4716 9553 4724
rect 12227 4716 12313 4724
rect 1187 4696 1653 4704
rect 1776 4696 2573 4704
rect 1776 4684 1784 4696
rect 2967 4696 4373 4704
rect 4727 4696 4893 4704
rect 5056 4704 5064 4713
rect 4907 4696 5064 4704
rect 5616 4696 5944 4704
rect 1687 4676 1784 4684
rect 2067 4676 2153 4684
rect 3027 4676 3673 4684
rect 3747 4676 4233 4684
rect 4247 4676 4353 4684
rect 5167 4676 5493 4684
rect 5616 4684 5624 4696
rect 5567 4676 5624 4684
rect 5767 4676 5893 4684
rect 5936 4684 5944 4696
rect 6187 4696 7493 4704
rect 8187 4696 8953 4704
rect 8967 4696 9173 4704
rect 9187 4696 9573 4704
rect 10056 4696 10313 4704
rect 5936 4676 6253 4684
rect 6567 4676 6812 4684
rect 6847 4676 7613 4684
rect 8207 4676 8673 4684
rect 9187 4676 9313 4684
rect 10056 4684 10064 4696
rect 10367 4696 11173 4704
rect 9547 4676 10064 4684
rect 10316 4684 10324 4693
rect 10316 4676 10664 4684
rect 1027 4656 1113 4664
rect 1527 4656 2693 4664
rect 2987 4656 3713 4664
rect 4287 4656 4353 4664
rect 4407 4656 4613 4664
rect 4927 4656 5613 4664
rect 5807 4656 5873 4664
rect 5927 4656 6273 4664
rect 6747 4656 8853 4664
rect 9347 4656 10073 4664
rect 10087 4656 10633 4664
rect 10656 4664 10664 4676
rect 11147 4676 11373 4684
rect 11667 4676 11973 4684
rect 12167 4676 12293 4684
rect 10656 4656 10733 4664
rect 11107 4656 12033 4664
rect 1267 4636 1413 4644
rect 1587 4636 2413 4644
rect 2747 4636 3033 4644
rect 4007 4636 5773 4644
rect 6947 4636 7673 4644
rect 8887 4636 9093 4644
rect 9467 4636 10513 4644
rect 667 4616 993 4624
rect 1007 4616 1073 4624
rect 1507 4616 2424 4624
rect -24 4596 513 4604
rect 1127 4596 1204 4604
rect 787 4576 1013 4584
rect -24 4556 173 4564
rect 347 4556 473 4564
rect 487 4559 553 4567
rect 707 4559 733 4567
rect 1093 4564 1107 4573
rect 1093 4560 1144 4564
rect 1096 4556 1144 4560
rect 847 4536 1113 4544
rect 267 4513 433 4521
rect 507 4516 693 4524
rect 1136 4524 1144 4556
rect 1196 4544 1204 4596
rect 1627 4596 1873 4604
rect 2207 4596 2393 4604
rect 2416 4604 2424 4616
rect 2767 4616 2913 4624
rect 3727 4616 3873 4624
rect 3967 4616 4433 4624
rect 4627 4616 5533 4624
rect 5867 4616 6013 4624
rect 6433 4624 6447 4633
rect 6227 4616 6284 4624
rect 6433 4620 6653 4624
rect 6436 4616 6653 4620
rect 2416 4596 3213 4604
rect 3747 4596 4664 4604
rect 4656 4587 4664 4596
rect 5527 4596 6113 4604
rect 6276 4604 6284 4616
rect 6667 4616 6873 4624
rect 7507 4616 8433 4624
rect 8507 4616 8713 4624
rect 9096 4624 9104 4633
rect 9096 4616 9893 4624
rect 10287 4616 10473 4624
rect 10927 4616 11433 4624
rect 11916 4616 12053 4624
rect 11916 4607 11924 4616
rect 6207 4596 6264 4604
rect 6276 4600 6324 4604
rect 6276 4596 6327 4600
rect 1413 4564 1427 4573
rect 1776 4576 2024 4584
rect 1776 4564 1784 4576
rect 1413 4560 1784 4564
rect 1416 4556 1784 4560
rect 2016 4564 2024 4576
rect 2447 4576 2493 4584
rect 3667 4576 3693 4584
rect 4667 4576 5313 4584
rect 2016 4556 2384 4564
rect 2787 4559 2813 4567
rect 2907 4556 2973 4564
rect 1196 4536 1233 4544
rect 1527 4536 1633 4544
rect 1867 4539 1993 4547
rect 2187 4536 2353 4544
rect 2376 4544 2384 4556
rect 3067 4559 3133 4567
rect 3387 4559 3453 4567
rect 3507 4556 3533 4564
rect 3907 4556 4033 4564
rect 4167 4559 4273 4567
rect 4447 4559 4513 4567
rect 4987 4559 5013 4567
rect 5087 4556 5353 4564
rect 2376 4536 2433 4544
rect 3456 4536 3653 4544
rect 1136 4516 1493 4524
rect 1607 4516 1873 4524
rect 2527 4513 2593 4521
rect 2807 4516 2873 4524
rect 2887 4513 2913 4521
rect 3047 4516 3153 4524
rect 3247 4516 3273 4524
rect 3456 4524 3464 4536
rect 5196 4536 5413 4544
rect 3447 4516 3493 4524
rect 3647 4516 3693 4524
rect 3907 4513 3933 4521
rect 4587 4516 4693 4524
rect 5196 4524 5204 4536
rect 4707 4516 5204 4524
rect 5587 4513 5653 4521
rect 5856 4524 5864 4573
rect 5876 4527 5884 4556
rect 6233 4564 6247 4573
rect 6087 4556 6164 4564
rect 6216 4560 6247 4564
rect 6156 4547 6164 4556
rect 6213 4556 6244 4560
rect 6213 4547 6227 4556
rect 6027 4536 6144 4544
rect 6156 4536 6173 4547
rect 5876 4516 5893 4527
rect 5880 4513 5893 4516
rect 6136 4524 6144 4536
rect 6160 4533 6173 4536
rect 6256 4544 6264 4596
rect 6313 4587 6327 4596
rect 7107 4596 7133 4604
rect 9287 4596 9673 4604
rect 10176 4596 10553 4604
rect 6627 4579 6713 4587
rect 10176 4587 10184 4596
rect 10747 4596 11913 4604
rect 7447 4576 7473 4584
rect 8027 4576 8053 4584
rect 8347 4576 8493 4584
rect 9527 4576 10173 4584
rect 10607 4576 10693 4584
rect 11347 4576 11453 4584
rect 11907 4576 11953 4584
rect 12207 4576 12253 4584
rect 12267 4576 12313 4584
rect 6847 4558 7033 4566
rect 7647 4559 7733 4567
rect 8147 4559 8193 4567
rect 8247 4559 8313 4567
rect 8587 4556 8733 4564
rect 8967 4564 8980 4567
rect 8967 4553 8984 4564
rect 9007 4559 9073 4567
rect 9287 4559 9333 4567
rect 9347 4556 9393 4564
rect 9567 4556 9893 4564
rect 10367 4559 10393 4567
rect 10827 4559 10873 4567
rect 11747 4556 11833 4564
rect 6376 4536 6453 4544
rect 6376 4524 6384 4536
rect 6587 4536 6673 4544
rect 6136 4516 6244 4524
rect 567 4496 793 4504
rect 847 4496 1433 4504
rect 1856 4496 1893 4504
rect 1856 4487 1864 4496
rect 2267 4496 2353 4504
rect 2447 4496 2693 4504
rect 2787 4496 3013 4504
rect 3027 4496 3053 4504
rect 3067 4496 3324 4504
rect 1847 4476 1864 4487
rect 1847 4473 1860 4476
rect 2387 4476 2413 4484
rect 2427 4476 2833 4484
rect 3316 4484 3324 4496
rect 4147 4496 4293 4504
rect 4427 4496 4813 4504
rect 5047 4496 5213 4504
rect 5427 4496 5524 4504
rect 3316 4476 4133 4484
rect 4247 4476 4393 4484
rect 4567 4476 4593 4484
rect 5147 4476 5293 4484
rect 5516 4484 5524 4496
rect 5667 4496 5713 4504
rect 5767 4496 5813 4504
rect 6047 4496 6093 4504
rect 6236 4504 6244 4516
rect 6296 4516 6384 4524
rect 6936 4523 7093 4524
rect 6296 4504 6304 4516
rect 6947 4516 7093 4523
rect 7207 4516 7233 4524
rect 8976 4524 8984 4553
rect 11216 4544 11224 4556
rect 11136 4540 11224 4544
rect 11133 4536 11224 4540
rect 11133 4527 11147 4536
rect 11476 4527 11484 4556
rect 12047 4556 12184 4564
rect 7727 4513 8073 4521
rect 8227 4513 8273 4521
rect 8407 4513 8473 4521
rect 8787 4513 8853 4521
rect 9027 4516 9093 4524
rect 9207 4513 9253 4521
rect 9307 4516 9353 4524
rect 9607 4516 9653 4524
rect 10167 4513 10293 4521
rect 10667 4513 10953 4521
rect 11146 4520 11147 4527
rect 11167 4516 11273 4524
rect 11476 4516 11493 4527
rect 11480 4513 11493 4516
rect 11936 4524 11944 4553
rect 12176 4544 12184 4556
rect 12176 4540 12244 4544
rect 12176 4536 12247 4540
rect 12233 4527 12247 4536
rect 12336 4527 12344 4553
rect 11647 4513 11713 4521
rect 11936 4516 11993 4524
rect 6236 4496 6304 4504
rect 6647 4496 6813 4504
rect 8527 4496 8664 4504
rect 5516 4476 5853 4484
rect 5907 4476 6004 4484
rect 5996 4467 6004 4476
rect 6087 4476 6193 4484
rect 6313 4484 6327 4493
rect 6313 4480 6384 4484
rect 6316 4476 6384 4480
rect 1507 4456 2433 4464
rect 2447 4456 2553 4464
rect 3307 4456 3573 4464
rect 3587 4456 3913 4464
rect 3927 4456 4933 4464
rect 5327 4456 5513 4464
rect 5787 4456 5853 4464
rect 5927 4456 5973 4464
rect 5996 4456 6013 4467
rect 6000 4453 6013 4456
rect 6187 4456 6273 4464
rect 6376 4464 6384 4476
rect 7387 4476 7513 4484
rect 7527 4476 7953 4484
rect 8087 4476 8253 4484
rect 8447 4476 8633 4484
rect 8656 4484 8664 4496
rect 9547 4496 9953 4504
rect 10427 4496 10613 4504
rect 10707 4496 11093 4504
rect 11207 4496 11453 4504
rect 12227 4496 12313 4504
rect 8656 4476 9073 4484
rect 9627 4476 9933 4484
rect 10847 4476 10893 4484
rect 6376 4460 6544 4464
rect 6376 4456 6547 4460
rect 6533 4447 6547 4456
rect 6787 4456 6933 4464
rect 9787 4456 9853 4464
rect 10347 4456 11013 4464
rect 11027 4456 11513 4464
rect 11687 4456 11773 4464
rect 787 4436 1033 4444
rect 1447 4436 2193 4444
rect 3987 4436 4153 4444
rect 4387 4436 4533 4444
rect 4807 4436 4873 4444
rect 5807 4436 5953 4444
rect 6067 4436 6193 4444
rect 7447 4436 7613 4444
rect 7867 4436 7993 4444
rect 8307 4436 9193 4444
rect 9267 4436 9393 4444
rect 9447 4436 9793 4444
rect 10067 4436 10733 4444
rect 10836 4436 11004 4444
rect 707 4416 1733 4424
rect 1867 4416 1973 4424
rect 2147 4416 2293 4424
rect 3587 4416 4613 4424
rect 5467 4416 6233 4424
rect 7047 4416 7413 4424
rect 8027 4416 8053 4424
rect 8647 4416 8873 4424
rect 8947 4416 9413 4424
rect 10836 4424 10844 4436
rect 9727 4416 10844 4424
rect 10996 4424 11004 4436
rect 11127 4436 11313 4444
rect 11567 4436 11993 4444
rect 10996 4416 11053 4424
rect 11627 4416 11653 4424
rect 1607 4396 1693 4404
rect 2487 4396 2633 4404
rect 2767 4396 2813 4404
rect 2927 4396 3333 4404
rect 3356 4396 4773 4404
rect 767 4376 873 4384
rect 887 4376 1493 4384
rect 1547 4376 1773 4384
rect 1787 4376 2273 4384
rect 2287 4376 2653 4384
rect 2667 4376 2873 4384
rect 3356 4384 3364 4396
rect 5507 4396 5573 4404
rect 6267 4396 6433 4404
rect 7087 4396 7133 4404
rect 7147 4396 7193 4404
rect 7567 4396 7733 4404
rect 8007 4396 8353 4404
rect 8367 4396 8513 4404
rect 8627 4396 9333 4404
rect 9376 4396 9613 4404
rect 2887 4376 3364 4384
rect 3427 4376 3573 4384
rect 3887 4376 3992 4384
rect 4027 4376 4353 4384
rect 4447 4376 4533 4384
rect 4947 4376 5113 4384
rect 5127 4376 5313 4384
rect 5507 4376 5553 4384
rect 5747 4376 5913 4384
rect 6027 4376 6113 4384
rect 6287 4376 6453 4384
rect 8207 4376 8473 4384
rect 8647 4376 8693 4384
rect 9376 4384 9384 4396
rect 10347 4396 10753 4404
rect 10867 4396 11473 4404
rect 11487 4396 11753 4404
rect 11767 4396 11953 4404
rect 11967 4396 12273 4404
rect 8827 4376 9384 4384
rect 9667 4376 9733 4384
rect 9747 4376 10153 4384
rect 10407 4376 10613 4384
rect 10967 4376 11193 4384
rect 11207 4376 11293 4384
rect 11307 4376 11413 4384
rect 1667 4356 1753 4364
rect 4787 4356 5453 4364
rect 5467 4356 5953 4364
rect 267 4339 413 4347
rect 507 4339 533 4347
rect 1387 4336 1413 4344
rect 1756 4344 1764 4353
rect 6267 4356 6293 4364
rect 7407 4356 7493 4364
rect 7587 4356 7873 4364
rect 7887 4356 7933 4364
rect 9087 4356 9513 4364
rect 1756 4336 1933 4344
rect 2047 4336 2233 4344
rect 2387 4336 2533 4344
rect 3027 4344 3040 4347
rect 3027 4333 3044 4344
rect 3107 4339 3193 4347
rect 607 4316 633 4324
rect 647 4316 833 4324
rect 887 4313 1033 4321
rect 1167 4316 1233 4324
rect -24 4296 213 4304
rect 427 4296 713 4304
rect 1447 4296 1613 4304
rect 1687 4296 1704 4304
rect 1696 4284 1704 4296
rect 2007 4293 2373 4301
rect 2667 4296 2693 4304
rect 2707 4296 2813 4304
rect 3036 4304 3044 4333
rect 3287 4336 3313 4344
rect 3667 4336 3713 4344
rect 4147 4336 4413 4344
rect 5167 4339 5253 4347
rect 5527 4336 6113 4344
rect 6487 4339 6513 4347
rect 6556 4336 6833 4344
rect 6887 4339 6913 4347
rect 7487 4339 7613 4347
rect 4827 4316 5224 4324
rect 3407 4293 3793 4301
rect 4267 4296 4353 4304
rect 4407 4296 4613 4304
rect 4687 4296 4913 4304
rect 5216 4304 5224 4316
rect 6556 4324 6564 4336
rect 6147 4316 6344 4324
rect 5067 4296 5173 4304
rect 5387 4293 5433 4301
rect 6336 4304 6344 4316
rect 6536 4316 6564 4324
rect 7356 4324 7364 4336
rect 7727 4336 8053 4344
rect 8247 4339 8313 4347
rect 8376 4336 8613 4344
rect 8376 4324 8384 4336
rect 9047 4336 9064 4344
rect 9307 4339 9473 4347
rect 9567 4339 9633 4347
rect 9807 4339 9873 4347
rect 10007 4339 10093 4347
rect 10107 4336 10173 4344
rect 7356 4316 8384 4324
rect 6536 4304 6544 4316
rect 9056 4307 9064 4336
rect 10387 4339 10413 4347
rect 10427 4336 10653 4344
rect 10927 4339 10953 4347
rect 11287 4336 11433 4344
rect 11687 4336 11704 4344
rect 11887 4339 11953 4347
rect 9107 4316 9433 4324
rect 5547 4296 5753 4304
rect 5827 4296 6013 4304
rect 6027 4293 6073 4301
rect 6336 4296 6544 4304
rect 6587 4293 6673 4301
rect 6927 4296 6953 4304
rect 6967 4296 7093 4304
rect 7687 4293 7713 4301
rect 8107 4296 8173 4304
rect 8507 4293 8693 4301
rect 9207 4296 9273 4304
rect 10856 4304 10864 4333
rect 11696 4307 11704 4336
rect 12127 4316 12244 4324
rect 9387 4296 9533 4304
rect 9947 4293 10033 4301
rect 10287 4293 10593 4301
rect 10647 4293 10673 4301
rect 10856 4296 10873 4304
rect 11147 4293 11273 4301
rect 11507 4296 11693 4304
rect 12236 4304 12244 4316
rect 12296 4307 12304 4333
rect 11987 4293 12053 4301
rect 12236 4296 12253 4304
rect 1696 4276 1733 4284
rect 2367 4276 2513 4284
rect 2527 4276 2633 4284
rect 3667 4276 3773 4284
rect 3847 4276 3873 4284
rect 4167 4276 4273 4284
rect 4807 4276 4893 4284
rect 5807 4276 6313 4284
rect 6327 4276 6373 4284
rect 7147 4276 7293 4284
rect 7647 4276 7913 4284
rect 8067 4276 8213 4284
rect 8236 4276 8433 4284
rect 1687 4256 1713 4264
rect 1967 4256 2033 4264
rect 2307 4256 2673 4264
rect 2807 4256 2913 4264
rect 3087 4256 3513 4264
rect 4607 4256 5513 4264
rect 5647 4256 6393 4264
rect 6447 4256 6573 4264
rect 6616 4256 6853 4264
rect 1707 4236 1753 4244
rect 3027 4236 3053 4244
rect 3647 4236 3773 4244
rect 3907 4236 4573 4244
rect 4647 4236 5033 4244
rect 5147 4236 5753 4244
rect 5927 4236 6053 4244
rect 6616 4244 6624 4256
rect 6867 4256 7113 4264
rect 7327 4256 7373 4264
rect 8236 4264 8244 4276
rect 8647 4276 8753 4284
rect 8807 4276 9653 4284
rect 9707 4276 10104 4284
rect 7427 4256 8244 4264
rect 8427 4256 8473 4264
rect 8667 4256 8733 4264
rect 9007 4256 9633 4264
rect 9647 4256 10073 4264
rect 10096 4264 10104 4276
rect 11167 4276 11233 4284
rect 11587 4276 11733 4284
rect 10096 4256 10353 4264
rect 10667 4256 10953 4264
rect 11887 4256 11933 4264
rect 12107 4256 12133 4264
rect 6507 4236 6624 4244
rect 6827 4236 6873 4244
rect 6887 4236 7233 4244
rect 7287 4236 8793 4244
rect 8967 4236 9273 4244
rect 9287 4236 9453 4244
rect 9787 4236 10052 4244
rect 10076 4244 10084 4253
rect 10076 4236 10413 4244
rect 11227 4236 11293 4244
rect 11307 4236 11413 4244
rect 11427 4236 11433 4244
rect 11447 4236 11713 4244
rect 12207 4236 12253 4244
rect 3387 4216 3493 4224
rect 3667 4216 4013 4224
rect 4727 4216 5713 4224
rect 5787 4216 6073 4224
rect 6227 4216 6353 4224
rect 6487 4216 6753 4224
rect 6767 4216 6913 4224
rect 7507 4216 9013 4224
rect 9776 4224 9784 4233
rect 9347 4216 9784 4224
rect 10487 4216 10753 4224
rect 11187 4216 11293 4224
rect 11967 4216 12053 4224
rect 1147 4196 1493 4204
rect 1507 4196 2533 4204
rect 2607 4196 2833 4204
rect 3207 4196 4313 4204
rect 4587 4196 4673 4204
rect 4967 4196 5293 4204
rect 5867 4196 6333 4204
rect 6547 4196 6633 4204
rect 6787 4196 6853 4204
rect 8147 4196 8233 4204
rect 8427 4196 9033 4204
rect 9227 4196 9353 4204
rect 9987 4196 10113 4204
rect 10167 4196 10353 4204
rect 10367 4196 11493 4204
rect 11667 4196 11753 4204
rect 547 4176 1953 4184
rect 2567 4176 2893 4184
rect 3367 4176 3453 4184
rect 3467 4176 4153 4184
rect 5407 4176 5613 4184
rect 5727 4176 5793 4184
rect 5927 4176 6093 4184
rect 6487 4176 6893 4184
rect 7027 4176 7253 4184
rect 8667 4176 8833 4184
rect 8847 4176 9093 4184
rect 9447 4176 9693 4184
rect 667 4156 813 4164
rect 827 4156 1193 4164
rect 1207 4156 1833 4164
rect 2147 4156 2293 4164
rect 2727 4156 3013 4164
rect 3067 4156 3184 4164
rect 307 4136 593 4144
rect 2407 4136 3033 4144
rect 3176 4144 3184 4156
rect 3567 4156 3793 4164
rect 4327 4156 4573 4164
rect 4587 4156 5253 4164
rect 5267 4156 8613 4164
rect 8687 4156 8793 4164
rect 9027 4156 9713 4164
rect 9887 4156 10813 4164
rect 10967 4156 11553 4164
rect 3176 4136 3513 4144
rect 3856 4136 3893 4144
rect 1827 4116 2373 4124
rect 2687 4116 2853 4124
rect 3107 4116 3173 4124
rect 3407 4116 3493 4124
rect 3667 4116 3752 4124
rect 3856 4124 3864 4136
rect 4707 4136 5073 4144
rect 5327 4136 5433 4144
rect 6807 4136 7073 4144
rect 7127 4136 7413 4144
rect 8467 4136 8573 4144
rect 8647 4136 8713 4144
rect 8967 4136 9253 4144
rect 11407 4136 11513 4144
rect 3787 4116 3864 4124
rect 5287 4116 5453 4124
rect 5527 4116 6044 4124
rect 767 4096 1393 4104
rect 1887 4096 3633 4104
rect 3967 4096 4553 4104
rect 4567 4096 4713 4104
rect 6036 4104 6044 4116
rect 7207 4116 7773 4124
rect 7787 4116 9053 4124
rect 9307 4116 9473 4124
rect 10827 4116 11273 4124
rect 6036 4096 6513 4104
rect 6527 4096 6993 4104
rect 8107 4096 8253 4104
rect 8727 4096 8813 4104
rect 8827 4096 8953 4104
rect 9687 4096 9813 4104
rect 9967 4096 10653 4104
rect 2487 4076 2633 4084
rect 2647 4076 2713 4084
rect 2827 4076 2933 4084
rect 3127 4084 3140 4087
rect 3127 4073 3144 4084
rect 3327 4076 3473 4084
rect 4227 4076 4464 4084
rect 567 4056 713 4064
rect 1387 4056 1453 4064
rect 1547 4056 1773 4064
rect 1787 4056 1813 4064
rect 2147 4056 2173 4064
rect -24 4036 213 4044
rect 307 4036 473 4044
rect 1647 4039 1733 4047
rect 2196 4044 2204 4073
rect 3136 4064 3144 4073
rect 3136 4056 3553 4064
rect 3927 4056 3993 4064
rect 4456 4064 4464 4076
rect 4947 4076 5053 4084
rect 5767 4076 5933 4084
rect 6027 4076 6493 4084
rect 6627 4076 6793 4084
rect 7167 4076 7353 4084
rect 8707 4076 8973 4084
rect 9093 4084 9107 4093
rect 9093 4080 9333 4084
rect 9096 4076 9333 4080
rect 10527 4076 10833 4084
rect 10847 4076 11453 4084
rect 11567 4076 11773 4084
rect 4456 4056 4633 4064
rect 4887 4059 5113 4067
rect 5827 4056 5913 4064
rect 6087 4064 6100 4067
rect 6087 4053 6104 4064
rect 7087 4056 7233 4064
rect 8407 4056 8513 4064
rect 9707 4056 9993 4064
rect 10007 4056 10313 4064
rect 2196 4036 2493 4044
rect 2627 4039 2853 4047
rect 2907 4039 3053 4047
rect 3207 4046 3284 4047
rect 3207 4039 3273 4046
rect 667 4016 852 4024
rect 887 4019 973 4027
rect 1247 4013 1373 4021
rect 1607 4019 1993 4027
rect 2196 4024 2204 4036
rect 2267 4013 2353 4021
rect 2367 4013 2553 4021
rect 3156 4024 3164 4036
rect 3407 4036 3533 4044
rect 3687 4039 3753 4047
rect 3807 4036 4173 4044
rect 4747 4036 4773 4044
rect 3047 4016 3164 4024
rect 4976 4007 4984 4033
rect 5016 4024 5024 4036
rect 5087 4036 5264 4044
rect 5016 4016 5133 4024
rect 5256 4024 5264 4036
rect 5256 4016 5273 4024
rect 5456 4027 5464 4053
rect 5727 4036 5773 4044
rect 5887 4036 6053 4044
rect 6096 4044 6104 4053
rect 6096 4036 6184 4044
rect 6227 4039 6273 4047
rect 6696 4046 6753 4047
rect 6176 4024 6184 4036
rect 6707 4039 6753 4046
rect 7107 4036 7333 4044
rect 7056 4024 7064 4036
rect 7407 4036 7593 4044
rect 7867 4036 7993 4044
rect 8147 4039 8213 4047
rect 8267 4039 8373 4047
rect 6176 4016 6204 4024
rect 7056 4016 7193 4024
rect 527 3996 573 4004
rect 1407 3996 1473 4004
rect 1707 3996 1793 4004
rect 1847 3996 2133 4004
rect 2787 3993 2873 4001
rect 3067 3996 3173 4004
rect 3496 3996 3513 4004
rect 507 3976 1533 3984
rect 3496 3984 3504 3996
rect 3667 3993 3733 4001
rect 3987 3996 4113 4004
rect 4527 3993 4573 4001
rect 4727 3996 4784 4004
rect 4776 3987 4784 3996
rect 5447 3996 5533 4004
rect 5667 3996 6153 4004
rect 6196 4004 6204 4016
rect 7596 4016 7844 4024
rect 6196 3996 6293 4004
rect 6547 3996 6613 4004
rect 6827 3996 6972 4004
rect 7007 3996 7073 4004
rect 7327 3993 7393 4001
rect 7596 4004 7604 4016
rect 7836 4004 7844 4016
rect 7467 3996 7573 4004
rect 7587 3996 7604 4004
rect 7787 3993 7813 4001
rect 7836 3996 7873 4004
rect 8007 3993 8073 4001
rect 8127 3996 8313 4004
rect 8616 4004 8624 4033
rect 8936 4024 8944 4036
rect 9047 4036 9213 4044
rect 9227 4036 9653 4044
rect 9667 4036 9733 4044
rect 9987 4039 10033 4047
rect 10507 4039 10553 4047
rect 10607 4039 10693 4047
rect 10747 4036 10793 4044
rect 10887 4036 10913 4044
rect 10927 4036 11213 4044
rect 11287 4039 11473 4047
rect 11707 4036 11873 4044
rect 12007 4036 12133 4044
rect 8936 4016 9013 4024
rect 11687 4016 11913 4024
rect 12296 4007 12304 4033
rect 8616 3996 8673 4004
rect 3267 3976 3504 3984
rect 3567 3976 3953 3984
rect 4776 3976 4793 3987
rect 4780 3973 4793 3976
rect 5767 3976 5873 3984
rect 6387 3976 6513 3984
rect 7867 3976 7893 3984
rect 8047 3983 8084 3984
rect 8047 3976 8073 3983
rect 8367 3976 8533 3984
rect 9093 3984 9107 3993
rect 9207 3993 9293 4001
rect 9347 3996 9453 4004
rect 9767 3996 9833 4004
rect 9947 3996 10013 4004
rect 10067 3993 10093 4001
rect 10287 3993 10353 4001
rect 10587 3996 10713 4004
rect 11067 3993 11193 4001
rect 11407 3996 11453 4004
rect 11787 3993 12013 4001
rect 8967 3980 9107 3984
rect 8967 3976 9104 3980
rect 11927 3976 11973 3984
rect 607 3956 693 3964
rect 747 3956 853 3964
rect 1567 3956 1873 3964
rect 1887 3956 3133 3964
rect 3487 3956 3672 3964
rect 3707 3956 3873 3964
rect 4467 3956 4733 3964
rect 4747 3956 4813 3964
rect 4967 3956 4993 3964
rect 5127 3956 5453 3964
rect 5607 3956 6073 3964
rect 6307 3956 6353 3964
rect 6507 3956 6713 3964
rect 7007 3956 7173 3964
rect 7347 3956 7673 3964
rect 8607 3956 8713 3964
rect 8807 3956 9093 3964
rect 9167 3956 9253 3964
rect 9427 3956 9993 3964
rect 10047 3956 10113 3964
rect 10487 3956 10593 3964
rect 11407 3956 11713 3964
rect 267 3936 553 3944
rect 1427 3936 1513 3944
rect 1687 3936 1733 3944
rect 2387 3936 2913 3944
rect 2987 3936 3124 3944
rect 3116 3927 3124 3936
rect 3287 3936 3773 3944
rect 4047 3936 5053 3944
rect 5256 3940 5633 3944
rect 5253 3936 5633 3940
rect 5253 3927 5267 3936
rect 5887 3936 6013 3944
rect 6407 3936 6773 3944
rect 6787 3936 7153 3944
rect 7587 3936 7973 3944
rect 8207 3936 8453 3944
rect 10767 3936 11133 3944
rect 11227 3936 11373 3944
rect 11487 3936 11613 3944
rect 11716 3944 11724 3953
rect 11716 3936 12273 3944
rect 636 3916 1173 3924
rect 636 3907 644 3916
rect 2027 3916 2344 3924
rect 367 3896 633 3904
rect 707 3896 1133 3904
rect 1176 3904 1184 3913
rect 1176 3896 1413 3904
rect 2187 3896 2293 3904
rect 2336 3904 2344 3916
rect 2387 3916 2693 3924
rect 3116 3916 3133 3927
rect 3120 3913 3133 3916
rect 3527 3916 3893 3924
rect 4087 3916 4273 3924
rect 4387 3916 4533 3924
rect 4907 3916 5033 3924
rect 5367 3916 5753 3924
rect 5776 3916 6244 3924
rect 2336 3896 2433 3904
rect 3107 3896 3273 3904
rect 3516 3896 4413 3904
rect 1407 3876 2953 3884
rect 3516 3884 3524 3896
rect 4687 3896 4733 3904
rect 4787 3896 4952 3904
rect 4987 3896 5093 3904
rect 5776 3904 5784 3916
rect 5527 3896 5784 3904
rect 5807 3896 5853 3904
rect 6027 3896 6113 3904
rect 6236 3904 6244 3916
rect 6796 3916 7153 3924
rect 6796 3904 6804 3916
rect 8027 3916 8253 3924
rect 9207 3916 9413 3924
rect 10507 3916 10853 3924
rect 11747 3916 12233 3924
rect 6236 3896 6804 3904
rect 6927 3896 7033 3904
rect 7207 3896 7273 3904
rect 7627 3896 8764 3904
rect 3067 3876 3524 3884
rect 3907 3876 4293 3884
rect 4947 3876 5353 3884
rect 5407 3876 6213 3884
rect 6227 3876 7113 3884
rect 7647 3876 8333 3884
rect 8607 3876 8733 3884
rect 8756 3884 8764 3896
rect 8847 3896 10213 3904
rect 11887 3896 12224 3904
rect 8756 3876 9173 3884
rect 9227 3876 9273 3884
rect 9427 3876 10413 3884
rect 10867 3876 11212 3884
rect 11247 3876 11313 3884
rect 11667 3876 11753 3884
rect 12216 3884 12224 3896
rect 12216 3876 12253 3884
rect 1447 3856 1753 3864
rect 2547 3856 2833 3864
rect 3587 3856 3853 3864
rect 4507 3856 4713 3864
rect 4807 3856 5273 3864
rect 5387 3856 6053 3864
rect 7167 3856 7933 3864
rect 8127 3856 8173 3864
rect 8327 3856 8453 3864
rect 9547 3856 9693 3864
rect 10007 3856 10353 3864
rect 10647 3856 10913 3864
rect 11147 3856 11593 3864
rect 11907 3856 12013 3864
rect 627 3836 673 3844
rect 2227 3836 2313 3844
rect 3027 3836 3253 3844
rect 3307 3836 3413 3844
rect 4027 3836 4093 3844
rect 4767 3836 5573 3844
rect 6807 3836 6853 3844
rect 7067 3836 7133 3844
rect 8487 3836 8653 3844
rect 9967 3836 10173 3844
rect 10187 3836 10313 3844
rect 10547 3836 10773 3844
rect 467 3816 513 3824
rect 1647 3819 1693 3827
rect 1967 3819 2213 3827
rect 2547 3819 2613 3827
rect 2747 3819 2773 3827
rect 2847 3816 2873 3824
rect 2887 3819 2973 3827
rect 3327 3816 3353 3824
rect 4067 3819 4113 3827
rect 4136 3816 4373 3824
rect -24 3776 13 3784
rect 576 3784 584 3796
rect 707 3793 833 3801
rect 196 3744 204 3771
rect 547 3776 584 3784
rect 667 3756 693 3764
rect 956 3747 964 3796
rect 1007 3756 1053 3764
rect 1096 3747 1104 3796
rect 1227 3793 1433 3801
rect 1507 3796 1573 3804
rect 1756 3796 2313 3804
rect 1756 3784 1764 3796
rect 2327 3796 2353 3804
rect 4136 3787 4144 3816
rect 5667 3816 5753 3824
rect 5807 3819 5933 3827
rect 6107 3819 6293 3827
rect 6387 3819 6453 3827
rect 6647 3819 6693 3827
rect 6767 3816 6873 3824
rect 7167 3816 7433 3824
rect 7567 3819 7653 3827
rect 7987 3819 8053 3827
rect 8427 3819 8553 3827
rect 8727 3819 8793 3827
rect 8927 3819 8973 3827
rect 9027 3819 9393 3827
rect 9487 3819 9533 3827
rect 9827 3819 9853 3827
rect 10087 3819 10253 3827
rect 10427 3819 10893 3827
rect 10907 3816 10933 3824
rect 11447 3816 11633 3824
rect 11647 3816 11873 3824
rect 11887 3819 11913 3827
rect 12267 3816 12384 3824
rect 4396 3796 4493 3804
rect 1667 3776 1713 3784
rect 1987 3776 2233 3784
rect 2247 3773 2393 3781
rect 3307 3773 3353 3781
rect 3767 3773 3813 3781
rect 3867 3773 4013 3781
rect 4187 3776 4333 3784
rect 4396 3784 4404 3796
rect 5996 3784 6004 3813
rect 6227 3796 6573 3804
rect 7156 3796 7613 3804
rect 7156 3784 7164 3796
rect 7767 3796 7813 3804
rect 4447 3773 4593 3781
rect 4667 3773 4753 3781
rect 5467 3773 5532 3781
rect 5567 3773 5813 3781
rect 6007 3773 6033 3781
rect 6367 3776 6613 3784
rect 6827 3773 6853 3781
rect 7147 3776 7164 3784
rect 7207 3776 7373 3784
rect 7687 3776 7953 3784
rect 7967 3776 8013 3784
rect 8347 3776 8513 3784
rect 8527 3776 8633 3784
rect 8647 3776 8764 3784
rect 2287 3756 2513 3764
rect 3047 3756 3273 3764
rect 4167 3756 4193 3764
rect 4987 3756 5333 3764
rect 5347 3756 5433 3764
rect 6087 3756 6144 3764
rect 196 3736 233 3744
rect 956 3736 969 3747
rect 960 3733 969 3736
rect 983 3736 984 3744
rect 1076 3736 1077 3744
rect 1091 3736 1104 3747
rect 1091 3733 1100 3736
rect 1767 3736 1873 3744
rect 1927 3736 2993 3744
rect 3647 3736 4093 3744
rect 4807 3736 4873 3744
rect 4887 3736 5373 3744
rect 5387 3736 5493 3744
rect 5507 3736 5873 3744
rect 5927 3736 6113 3744
rect 6136 3744 6144 3756
rect 7467 3756 8093 3764
rect 8167 3756 8213 3764
rect 8387 3756 8433 3764
rect 8756 3764 8764 3776
rect 8967 3776 9193 3784
rect 9307 3773 9373 3781
rect 9667 3773 9753 3781
rect 9907 3773 10053 3781
rect 10167 3773 10293 3781
rect 11047 3776 11093 3784
rect 12196 3784 12204 3813
rect 11607 3773 11693 3781
rect 12196 3776 12233 3784
rect 8756 3756 9193 3764
rect 9527 3756 9633 3764
rect 9647 3756 9793 3764
rect 10456 3756 10613 3764
rect 6136 3736 6433 3744
rect 6707 3736 7753 3744
rect 7927 3736 7993 3744
rect 8747 3736 8873 3744
rect 8887 3736 8953 3744
rect 9007 3736 9473 3744
rect 10456 3744 10464 3756
rect 10667 3756 10993 3764
rect 11427 3756 11513 3764
rect 11927 3756 12053 3764
rect 12267 3756 12313 3764
rect 10067 3736 10464 3744
rect 10487 3736 10513 3744
rect 10676 3736 10873 3744
rect 1936 3716 2373 3724
rect 1647 3696 1733 3704
rect 1936 3704 1944 3716
rect 2627 3716 3093 3724
rect 3667 3716 4553 3724
rect 4727 3716 5793 3724
rect 6007 3716 6073 3724
rect 6287 3716 6673 3724
rect 6727 3716 7113 3724
rect 7227 3716 7293 3724
rect 7427 3716 7553 3724
rect 7567 3716 7713 3724
rect 7887 3716 8053 3724
rect 8996 3724 9004 3733
rect 8567 3716 9004 3724
rect 9527 3716 9873 3724
rect 10676 3724 10684 3736
rect 10887 3736 10913 3744
rect 11647 3736 11733 3744
rect 12207 3736 12333 3744
rect 10307 3716 10684 3724
rect 10887 3716 11333 3724
rect 11627 3716 11652 3724
rect 11687 3716 11753 3724
rect 11967 3716 12093 3724
rect 1747 3696 1944 3704
rect 2207 3696 2453 3704
rect 2467 3696 3553 3704
rect 3607 3696 4193 3704
rect 4327 3696 4493 3704
rect 4847 3696 5693 3704
rect 5887 3696 6333 3704
rect 6387 3696 6653 3704
rect 6847 3696 7013 3704
rect 7027 3696 7773 3704
rect 8247 3696 8833 3704
rect 9267 3696 10113 3704
rect 10227 3696 11604 3704
rect 2487 3676 2933 3684
rect 3227 3676 4673 3684
rect 5447 3676 6733 3684
rect 6907 3676 8313 3684
rect 8907 3676 9133 3684
rect 9207 3676 9553 3684
rect 10027 3676 10533 3684
rect 10587 3676 10773 3684
rect 10787 3676 11193 3684
rect 11596 3684 11604 3696
rect 11596 3676 11933 3684
rect 11947 3676 12093 3684
rect 2087 3656 2413 3664
rect 2707 3656 2973 3664
rect 3567 3656 4013 3664
rect 4067 3656 4373 3664
rect 4556 3656 5293 3664
rect 1416 3636 1913 3644
rect 1416 3624 1424 3636
rect 2027 3636 2153 3644
rect 2356 3636 3433 3644
rect 2356 3627 2364 3636
rect 4556 3644 4564 3656
rect 5427 3656 6213 3664
rect 6467 3656 6833 3664
rect 7627 3656 8232 3664
rect 8267 3656 9673 3664
rect 10567 3656 12293 3664
rect 3947 3636 4564 3644
rect 4787 3636 4933 3644
rect 5147 3636 5233 3644
rect 5367 3636 6273 3644
rect 6407 3636 7013 3644
rect 7247 3636 7273 3644
rect 7647 3636 7733 3644
rect 7807 3636 8013 3644
rect 8427 3636 9244 3644
rect 27 3616 1424 3624
rect 1907 3616 2353 3624
rect 2747 3616 2773 3624
rect 2987 3616 3153 3624
rect 3267 3616 3313 3624
rect 3907 3616 4213 3624
rect 5087 3616 5553 3624
rect 6067 3616 7193 3624
rect 9147 3616 9173 3624
rect 9236 3624 9244 3636
rect 9267 3636 9533 3644
rect 9727 3636 9893 3644
rect 9907 3636 10613 3644
rect 10987 3636 11713 3644
rect 11807 3636 11833 3644
rect 11987 3636 12053 3644
rect 9236 3616 10713 3624
rect 1627 3596 1713 3604
rect 1727 3596 2573 3604
rect 2587 3596 4473 3604
rect 4487 3596 4773 3604
rect 5207 3596 5313 3604
rect 5747 3596 5993 3604
rect 6087 3596 6553 3604
rect 6567 3596 7124 3604
rect 547 3576 773 3584
rect 1347 3576 1373 3584
rect 1807 3576 2473 3584
rect 2727 3576 3353 3584
rect 3407 3576 3893 3584
rect 4027 3576 4233 3584
rect 5467 3576 5553 3584
rect 6307 3576 7073 3584
rect 7116 3584 7124 3596
rect 9007 3596 10413 3604
rect 10627 3596 11513 3604
rect 11827 3596 11893 3604
rect 7116 3576 7593 3584
rect 8147 3576 8193 3584
rect 8207 3576 8413 3584
rect 8467 3576 8533 3584
rect 9867 3576 10333 3584
rect 10387 3576 10413 3584
rect 11947 3576 12013 3584
rect 12247 3576 12364 3584
rect 227 3556 293 3564
rect 2527 3556 2673 3564
rect 3167 3556 3793 3564
rect 3807 3556 3953 3564
rect 4427 3556 4713 3564
rect 4907 3556 5033 3564
rect 5787 3556 5933 3564
rect 6587 3556 7613 3564
rect 7707 3556 8993 3564
rect 9667 3556 10173 3564
rect 10927 3556 10993 3564
rect 11127 3556 11153 3564
rect 11167 3556 11413 3564
rect 11427 3556 11753 3564
rect 11767 3556 11793 3564
rect 11807 3556 11873 3564
rect 11887 3556 11973 3564
rect 11987 3556 12213 3564
rect 12227 3556 12333 3564
rect 467 3536 553 3544
rect 567 3536 733 3544
rect 2187 3536 2233 3544
rect 4547 3536 4753 3544
rect 4767 3536 5224 3544
rect 267 3519 333 3527
rect 1027 3519 1053 3527
rect 1147 3519 1173 3527
rect 1387 3519 1433 3527
rect 247 3476 493 3484
rect 516 3467 524 3516
rect 816 3504 824 3516
rect 1436 3504 1444 3516
rect 1587 3516 1653 3524
rect 1667 3519 1693 3527
rect 2167 3519 2253 3527
rect 2427 3516 2493 3524
rect 2507 3516 2733 3524
rect 816 3496 1444 3504
rect 547 3476 653 3484
rect 807 3476 1013 3484
rect 1187 3476 1353 3484
rect 2756 3484 2764 3533
rect 2787 3516 3013 3524
rect 3027 3519 3093 3527
rect 3167 3516 3233 3524
rect 3247 3519 3373 3527
rect 3547 3519 3633 3527
rect 3847 3519 3893 3527
rect 3967 3516 4073 3524
rect 4347 3516 4444 3524
rect 3747 3496 4033 3504
rect 4436 3487 4444 3516
rect 4607 3516 4633 3524
rect 4847 3516 4953 3524
rect 4967 3516 5193 3524
rect 5216 3524 5224 3536
rect 5247 3536 5433 3544
rect 6027 3536 6293 3544
rect 6727 3536 7053 3544
rect 7127 3536 7173 3544
rect 7287 3536 7353 3544
rect 7947 3536 7973 3544
rect 8067 3536 8173 3544
rect 9487 3536 9793 3544
rect 5216 3516 5713 3524
rect 6007 3516 6233 3524
rect 6247 3516 6353 3524
rect 6607 3519 6673 3527
rect 6687 3519 6793 3527
rect 7427 3519 7553 3527
rect 7616 3516 7633 3524
rect 4487 3496 4924 3504
rect 1707 3476 1873 3484
rect 2007 3473 2393 3481
rect 2927 3473 3033 3481
rect 3267 3476 3313 3484
rect 3647 3476 3813 3484
rect 3867 3473 3913 3481
rect 4247 3473 4393 3481
rect 4916 3484 4924 3496
rect 7616 3487 7624 3516
rect 7767 3516 7873 3524
rect 8120 3524 8133 3527
rect 8116 3513 8133 3524
rect 8227 3519 8253 3527
rect 8567 3516 8753 3524
rect 8767 3516 8933 3524
rect 9167 3516 9293 3524
rect 8116 3504 8124 3513
rect 7916 3496 8124 3504
rect 8156 3496 8333 3504
rect 4916 3476 4933 3484
rect 5107 3476 5213 3484
rect 5307 3473 5453 3481
rect 5687 3476 5872 3484
rect 5896 3480 6093 3484
rect 5893 3476 6093 3480
rect 5893 3467 5907 3476
rect 6187 3476 6413 3484
rect 6627 3476 6913 3484
rect 6927 3476 6953 3484
rect 6967 3473 7133 3481
rect 7916 3484 7924 3496
rect 8156 3484 8164 3496
rect 9533 3504 9547 3513
rect 9916 3516 10093 3524
rect 10107 3519 10173 3527
rect 10267 3519 10313 3527
rect 10627 3516 10693 3524
rect 9916 3504 9924 3516
rect 10707 3516 10813 3524
rect 10827 3516 10933 3524
rect 11127 3524 11140 3527
rect 11127 3513 11144 3524
rect 9533 3500 9924 3504
rect 9536 3496 9924 3500
rect 7667 3473 7693 3481
rect 8527 3473 8553 3481
rect 8727 3473 8773 3481
rect 8947 3473 8973 3481
rect 9347 3476 9453 3484
rect 9847 3476 9873 3484
rect 10027 3476 10073 3484
rect 11136 3484 11144 3513
rect 11156 3504 11164 3516
rect 11227 3516 11453 3524
rect 11607 3519 12013 3527
rect 11156 3496 11333 3504
rect 10187 3476 10333 3484
rect 10467 3473 10573 3481
rect 10727 3473 10913 3481
rect 11387 3476 11433 3484
rect 1547 3456 1633 3464
rect 4567 3456 4693 3464
rect 4707 3456 4733 3464
rect 5567 3456 5853 3464
rect 7787 3456 7893 3464
rect 9107 3456 9473 3464
rect 9527 3456 9653 3464
rect 10107 3456 10153 3464
rect 11456 3464 11464 3516
rect 12227 3519 12253 3527
rect 12056 3487 12064 3513
rect 11647 3476 11693 3484
rect 11887 3476 11953 3484
rect 12007 3476 12053 3484
rect 12276 3484 12284 3533
rect 12333 3504 12347 3513
rect 12316 3500 12347 3504
rect 12316 3496 12344 3500
rect 12316 3484 12324 3496
rect 11456 3456 11613 3464
rect 347 3436 573 3444
rect 1127 3436 1293 3444
rect 1307 3436 2133 3444
rect 2227 3436 2713 3444
rect 3507 3436 4113 3444
rect 4407 3436 4473 3444
rect 5027 3436 5253 3444
rect 5276 3436 5753 3444
rect 1687 3416 1813 3424
rect 2267 3416 2433 3424
rect 3547 3416 3893 3424
rect 3907 3416 4133 3424
rect 4367 3416 4413 3424
rect 5276 3424 5284 3436
rect 5947 3436 6573 3444
rect 6867 3436 6932 3444
rect 6967 3436 7093 3444
rect 7107 3436 7393 3444
rect 7567 3436 7984 3444
rect 7976 3427 7984 3436
rect 8807 3436 9533 3444
rect 10407 3436 10853 3444
rect 10867 3436 10973 3444
rect 11147 3436 11253 3444
rect 11507 3436 11933 3444
rect 11947 3436 12033 3444
rect 12047 3436 12233 3444
rect 12356 3444 12364 3576
rect 12307 3436 12364 3444
rect 4667 3416 5284 3424
rect 7987 3416 8193 3424
rect 9227 3416 9253 3424
rect 9427 3416 9593 3424
rect 10227 3416 10753 3424
rect 11927 3416 11973 3424
rect 207 3396 273 3404
rect 847 3396 1073 3404
rect 1087 3396 3513 3404
rect 4867 3396 5473 3404
rect 5707 3396 6073 3404
rect 7407 3396 7573 3404
rect 9507 3396 9773 3404
rect 9827 3396 10793 3404
rect 10807 3396 11493 3404
rect 12207 3396 12333 3404
rect 327 3376 473 3384
rect 487 3376 1353 3384
rect 1607 3376 1733 3384
rect 3847 3376 3993 3384
rect 4307 3376 4353 3384
rect 5127 3376 5293 3384
rect 5727 3376 5953 3384
rect 6107 3376 6973 3384
rect 7027 3376 8193 3384
rect 8427 3376 8473 3384
rect 8607 3376 9353 3384
rect 9836 3376 10673 3384
rect 1007 3356 1153 3364
rect 2167 3356 2173 3364
rect 2187 3356 2253 3364
rect 2267 3356 2713 3364
rect 3107 3356 3533 3364
rect 3907 3356 3933 3364
rect 4327 3356 4933 3364
rect 5687 3356 5833 3364
rect 5907 3356 5973 3364
rect 7167 3356 8033 3364
rect 8596 3364 8604 3373
rect 8227 3356 8604 3364
rect 8947 3356 9273 3364
rect 9327 3356 9493 3364
rect 9836 3364 9844 3376
rect 11107 3376 11173 3384
rect 12227 3376 12273 3384
rect 9547 3356 9844 3364
rect 10587 3356 10773 3364
rect 11747 3356 11773 3364
rect 947 3336 1073 3344
rect 1407 3336 1513 3344
rect 1747 3336 1904 3344
rect 1896 3324 1904 3336
rect 3727 3336 4193 3344
rect 4427 3336 4593 3344
rect 4647 3336 4833 3344
rect 4987 3336 5413 3344
rect 5827 3336 6053 3344
rect 7047 3336 7273 3344
rect 7607 3336 8153 3344
rect 8207 3336 8873 3344
rect 11687 3336 11773 3344
rect 12207 3336 12293 3344
rect 1896 3316 2113 3324
rect 2427 3316 2633 3324
rect 3947 3316 3973 3324
rect 4967 3316 5393 3324
rect 5787 3316 6033 3324
rect 7347 3316 7613 3324
rect 9007 3316 9073 3324
rect 9287 3316 9613 3324
rect 9627 3316 9753 3324
rect 10547 3316 10633 3324
rect 11676 3316 11713 3324
rect 227 3299 293 3307
rect 567 3296 773 3304
rect 1047 3296 1233 3304
rect 1247 3296 1553 3304
rect 1567 3296 1613 3304
rect 1787 3296 1873 3304
rect 2487 3296 2673 3304
rect 2727 3299 2773 3307
rect 3247 3299 3273 3307
rect 3287 3299 3393 3307
rect 3767 3296 3873 3304
rect 3927 3296 4033 3304
rect 4107 3296 4313 3304
rect 4547 3296 4593 3304
rect 4727 3296 4873 3304
rect 4927 3296 5173 3304
rect 5187 3299 5273 3307
rect 5287 3296 5373 3304
rect 5447 3299 5493 3307
rect 5667 3296 5704 3304
rect 247 3256 453 3264
rect 507 3253 553 3261
rect 807 3253 833 3261
rect 1307 3253 1333 3261
rect 1447 3256 1653 3264
rect 1667 3253 1853 3261
rect 2147 3253 2213 3261
rect 2407 3253 2493 3261
rect 2647 3253 2693 3261
rect 2807 3256 2873 3264
rect 2887 3256 3193 3264
rect 3787 3256 3973 3264
rect 4067 3256 4253 3264
rect 4347 3253 4393 3261
rect 4627 3253 4693 3261
rect 4707 3253 4753 3261
rect 5696 3264 5704 3296
rect 5807 3296 5993 3304
rect 6007 3296 6193 3304
rect 6207 3296 6513 3304
rect 6567 3299 6613 3307
rect 6667 3296 6753 3304
rect 6827 3299 6873 3307
rect 7087 3299 7113 3307
rect 7156 3296 7293 3304
rect 7587 3299 7973 3307
rect 7156 3284 7164 3296
rect 8047 3296 8313 3304
rect 8467 3299 8493 3307
rect 8607 3296 8653 3304
rect 7136 3276 7164 3284
rect 8716 3284 8724 3296
rect 8807 3296 8933 3304
rect 9507 3299 9533 3307
rect 9556 3296 9713 3304
rect 10047 3299 10153 3307
rect 10167 3296 10253 3304
rect 8716 3276 9033 3284
rect 5367 3256 5413 3264
rect 5747 3253 5813 3261
rect 5867 3253 5973 3261
rect 6547 3253 6673 3261
rect 6807 3256 6993 3264
rect 7136 3264 7144 3276
rect 9196 3267 9204 3296
rect 9456 3284 9464 3296
rect 9556 3284 9564 3296
rect 10347 3299 10373 3307
rect 9456 3276 9564 3284
rect 11176 3284 11184 3296
rect 11176 3276 11313 3284
rect 7107 3256 7144 3264
rect 7327 3253 7393 3261
rect 7627 3253 7673 3261
rect 7847 3253 7873 3261
rect 7927 3253 8093 3261
rect 8207 3256 8253 3264
rect 8327 3256 8433 3264
rect 8747 3253 8793 3261
rect 8947 3256 9133 3264
rect 9187 3256 9204 3267
rect 9187 3253 9200 3256
rect 9227 3256 9253 3264
rect 9687 3256 9773 3264
rect 10287 3253 10513 3261
rect 10607 3253 10693 3261
rect 10707 3256 10824 3264
rect 4907 3236 5093 3244
rect 5107 3236 5193 3244
rect 6067 3236 6233 3244
rect 6247 3236 6473 3244
rect 7987 3236 8173 3244
rect 8527 3236 8573 3244
rect 9607 3236 9993 3244
rect 10067 3236 10113 3244
rect 10127 3236 10593 3244
rect 10816 3244 10824 3256
rect 10847 3253 11293 3261
rect 11387 3256 11513 3264
rect 11676 3264 11684 3316
rect 11927 3296 11953 3304
rect 12016 3264 12024 3296
rect 12016 3256 12053 3264
rect 12256 3264 12264 3313
rect 12300 3304 12313 3307
rect 12296 3293 12313 3304
rect 12296 3264 12304 3293
rect 12227 3256 12264 3264
rect 10816 3236 11193 3244
rect 11207 3236 11253 3244
rect 767 3216 1053 3224
rect 1067 3216 1373 3224
rect 1647 3216 1893 3224
rect 2747 3216 3913 3224
rect 4307 3216 4373 3224
rect 4507 3216 4853 3224
rect 5087 3216 5133 3224
rect 5487 3216 5813 3224
rect 6027 3216 6353 3224
rect 6507 3216 6553 3224
rect 6567 3216 6713 3224
rect 7067 3216 7193 3224
rect 7247 3216 7553 3224
rect 7907 3216 8353 3224
rect 9187 3216 9233 3224
rect 9547 3216 10393 3224
rect 10607 3216 10633 3224
rect 10767 3216 11153 3224
rect 11207 3216 11473 3224
rect 11487 3216 11753 3224
rect 12227 3216 12313 3224
rect 2207 3196 2593 3204
rect 3167 3196 3633 3204
rect 3747 3196 3833 3204
rect 4067 3196 4673 3204
rect 4687 3196 4953 3204
rect 5087 3196 5453 3204
rect 6527 3196 6833 3204
rect 7547 3196 7573 3204
rect 8027 3196 8152 3204
rect 8187 3196 8613 3204
rect 9387 3196 9493 3204
rect 9927 3196 10073 3204
rect 10787 3196 10873 3204
rect 11407 3196 12033 3204
rect 12207 3196 12293 3204
rect 2187 3176 2513 3184
rect 2527 3176 3653 3184
rect 4467 3176 5773 3184
rect 5827 3176 6493 3184
rect 6787 3176 6973 3184
rect 8127 3176 8273 3184
rect 8727 3176 8893 3184
rect 8967 3176 9313 3184
rect 9327 3176 10293 3184
rect 10307 3176 10553 3184
rect 10567 3176 10613 3184
rect 10687 3176 10833 3184
rect 10856 3176 11193 3184
rect 347 3156 1753 3164
rect 1907 3156 2893 3164
rect 3147 3156 3433 3164
rect 3967 3156 4493 3164
rect 4587 3156 4713 3164
rect 4967 3156 5613 3164
rect 5667 3156 5793 3164
rect 5887 3156 5973 3164
rect 6207 3156 6233 3164
rect 8887 3156 9253 3164
rect 9387 3156 9793 3164
rect 10856 3164 10864 3176
rect 11867 3176 11893 3184
rect 9847 3156 10864 3164
rect 11727 3156 11893 3164
rect 2607 3136 3593 3144
rect 3687 3136 4793 3144
rect 4907 3136 5073 3144
rect 5227 3136 5493 3144
rect 5507 3136 6013 3144
rect 6027 3136 7093 3144
rect 7147 3136 7913 3144
rect 8007 3136 9493 3144
rect 9547 3136 9664 3144
rect 1107 3116 1733 3124
rect 2927 3116 3113 3124
rect 3367 3116 3513 3124
rect 3647 3116 5153 3124
rect 6287 3116 7033 3124
rect 7247 3116 7593 3124
rect 8067 3116 8173 3124
rect 8247 3116 9473 3124
rect 9656 3124 9664 3136
rect 9967 3136 10273 3144
rect 11107 3136 11273 3144
rect 9656 3116 10333 3124
rect 10387 3116 10793 3124
rect 11007 3116 11353 3124
rect 11687 3116 12253 3124
rect 1907 3096 2473 3104
rect 2787 3096 3193 3104
rect 3867 3096 4093 3104
rect 4527 3096 4633 3104
rect 4647 3096 4893 3104
rect 5207 3096 5973 3104
rect 7127 3096 9533 3104
rect 9647 3096 10553 3104
rect 11147 3096 11593 3104
rect 187 3076 1284 3084
rect 1276 3067 1284 3076
rect 2447 3076 2753 3084
rect 2767 3076 3464 3084
rect 3456 3067 3464 3076
rect 4127 3076 5033 3084
rect 5087 3076 5273 3084
rect 5287 3076 5753 3084
rect 6747 3076 7353 3084
rect 7407 3076 7832 3084
rect 7867 3076 11713 3084
rect 1287 3056 1513 3064
rect 2227 3056 2504 3064
rect 887 3036 1273 3044
rect 2496 3044 2504 3056
rect 3047 3056 3373 3064
rect 3467 3056 3733 3064
rect 4027 3056 4313 3064
rect 4407 3056 4884 3064
rect 2496 3036 2793 3044
rect 3487 3036 3893 3044
rect 4876 3044 4884 3056
rect 5096 3056 5213 3064
rect 5096 3044 5104 3056
rect 6756 3056 7693 3064
rect 4876 3036 5104 3044
rect 5167 3036 5284 3044
rect 2307 3019 2433 3027
rect 3927 3016 4013 3024
rect 5276 3024 5284 3036
rect 5347 3036 5653 3044
rect 5736 3036 5853 3044
rect 5736 3024 5744 3036
rect 6756 3044 6764 3056
rect 7927 3056 8233 3064
rect 8867 3056 8952 3064
rect 8987 3056 9153 3064
rect 9267 3056 9833 3064
rect 10147 3056 10452 3064
rect 10487 3056 10533 3064
rect 11007 3056 11393 3064
rect 11447 3056 11684 3064
rect 6107 3036 6764 3044
rect 6847 3036 7013 3044
rect 7467 3036 7513 3044
rect 7767 3036 7953 3044
rect 8307 3036 8373 3044
rect 8427 3036 8813 3044
rect 9127 3036 9213 3044
rect 9227 3036 9893 3044
rect 9947 3036 10133 3044
rect 5276 3016 5744 3024
rect 6096 3024 6104 3033
rect 11127 3036 11233 3044
rect 11676 3044 11684 3056
rect 11676 3036 12193 3044
rect 5767 3016 6104 3024
rect 7267 3016 7313 3024
rect 7567 3016 8213 3024
rect 9667 3016 9713 3024
rect 10467 3016 10753 3024
rect 11567 3016 11624 3024
rect 187 3004 200 3007
rect 187 2993 204 3004
rect 227 2996 273 3004
rect 287 2996 393 3004
rect 587 2999 753 3007
rect 767 2996 893 3004
rect 196 2964 204 2993
rect 456 2984 464 2996
rect 1007 2996 1304 3004
rect 1567 2996 1813 3004
rect 456 2976 513 2984
rect 407 2953 433 2961
rect 747 2956 873 2964
rect 1296 2964 1304 2996
rect 947 2953 1013 2961
rect 1747 2953 1793 2961
rect 907 2936 1213 2944
rect 1856 2924 1864 2996
rect 2116 2984 2124 2996
rect 2376 2984 2384 2996
rect 2116 2976 2413 2984
rect 2816 2987 2824 3013
rect 3007 2999 3113 3007
rect 3207 2996 3553 3004
rect 3787 2996 4053 3004
rect 4336 2996 4593 3004
rect 4907 2999 4973 3007
rect 5387 2999 5593 3007
rect 5636 2996 5693 3004
rect 6747 2996 6893 3004
rect 2596 2964 2604 2976
rect 4336 2984 4344 2996
rect 4116 2976 4344 2984
rect 5136 2984 5144 2996
rect 5136 2976 5213 2984
rect 2447 2956 2604 2964
rect 3367 2956 3673 2964
rect 4116 2964 4124 2976
rect 5636 2967 5644 2996
rect 7527 2996 7673 3004
rect 6976 2984 6984 2996
rect 7767 2996 7993 3004
rect 8267 2999 8293 3007
rect 8347 2999 8473 3007
rect 8567 2999 8633 3007
rect 9167 2999 9253 3007
rect 9647 2996 9733 3004
rect 6976 2976 7073 2984
rect 3767 2953 3873 2961
rect 4087 2956 4124 2964
rect 4367 2956 4613 2964
rect 5347 2953 5413 2961
rect 6047 2953 6093 2961
rect 8076 2964 8084 2993
rect 6167 2956 6593 2964
rect 6607 2953 6713 2961
rect 6907 2953 6953 2961
rect 7687 2953 7733 2961
rect 8067 2956 8084 2964
rect 8836 2964 8844 2996
rect 10196 2996 10233 3004
rect 10196 2984 10204 2996
rect 10687 2996 10733 3004
rect 10807 2999 10953 3007
rect 11167 2999 11213 3007
rect 11267 2996 11344 3004
rect 11427 2999 11513 3007
rect 11616 3007 11624 3016
rect 11647 3016 12253 3024
rect 11616 3006 11640 3007
rect 11616 2996 11633 3006
rect 10027 2976 10204 2984
rect 8527 2956 8573 2964
rect 8836 2956 9093 2964
rect 9687 2953 9713 2961
rect 9807 2953 9953 2961
rect 10407 2956 10433 2964
rect 10627 2953 10653 2961
rect 11187 2956 11273 2964
rect 11336 2964 11344 2996
rect 11620 2993 11633 2996
rect 11736 2996 11993 3004
rect 11736 2964 11744 2996
rect 11336 2956 11453 2964
rect 11947 2953 11973 2961
rect 2807 2936 3033 2944
rect 3147 2936 3193 2944
rect 3447 2936 3493 2944
rect 3987 2936 4073 2944
rect 4147 2936 4553 2944
rect 4827 2936 4913 2944
rect 5327 2936 5433 2944
rect 5547 2936 5653 2944
rect 5667 2936 5713 2944
rect 6367 2936 6533 2944
rect 7007 2936 7153 2944
rect 7267 2936 7353 2944
rect 7367 2936 7493 2944
rect 9007 2936 9153 2944
rect 1807 2916 1864 2924
rect 2867 2916 2913 2924
rect 3347 2916 3513 2924
rect 3587 2916 3953 2924
rect 4667 2916 5053 2924
rect 5227 2916 5673 2924
rect 5967 2916 6113 2924
rect 6387 2916 6433 2924
rect 6447 2916 6833 2924
rect 7287 2916 7453 2924
rect 7587 2916 8313 2924
rect 8867 2916 9273 2924
rect 9587 2916 9853 2924
rect 10187 2916 10213 2924
rect 10707 2916 11133 2924
rect 11147 2916 11233 2924
rect 11387 2916 11473 2924
rect 467 2896 513 2904
rect 527 2896 933 2904
rect 947 2896 973 2904
rect 1207 2896 1533 2904
rect 1847 2896 2173 2904
rect 2367 2896 2453 2904
rect 2767 2896 4173 2904
rect 4187 2896 4313 2904
rect 5216 2904 5224 2913
rect 11587 2916 12013 2924
rect 4327 2896 5224 2904
rect 5707 2896 6333 2904
rect 7087 2896 7613 2904
rect 8367 2896 8773 2904
rect 8787 2896 9413 2904
rect 9627 2896 9773 2904
rect 10347 2896 10933 2904
rect 11507 2896 11813 2904
rect 1267 2876 2433 2884
rect 3027 2876 3273 2884
rect 3427 2876 3533 2884
rect 3707 2876 3733 2884
rect 4087 2876 4233 2884
rect 4367 2876 4873 2884
rect 4887 2876 4933 2884
rect 5007 2876 5753 2884
rect 7187 2876 7293 2884
rect 7607 2876 8053 2884
rect 9067 2876 9193 2884
rect 10007 2876 10033 2884
rect 10047 2876 10693 2884
rect 2427 2856 2753 2864
rect 2987 2856 3433 2864
rect 3536 2864 3544 2873
rect 3536 2856 4853 2864
rect 5587 2856 5713 2864
rect 6667 2856 6793 2864
rect 8267 2856 8432 2864
rect 8467 2856 9013 2864
rect 9027 2856 9113 2864
rect 9167 2856 9333 2864
rect 10507 2856 10573 2864
rect 10747 2856 11153 2864
rect 11247 2856 11573 2864
rect 11707 2856 11773 2864
rect 1367 2836 1833 2844
rect 2107 2836 2153 2844
rect 2767 2836 2853 2844
rect 2927 2836 3104 2844
rect 787 2816 993 2824
rect 1007 2816 1233 2824
rect 2187 2816 3073 2824
rect 3096 2824 3104 2836
rect 3456 2836 3973 2844
rect 3456 2824 3464 2836
rect 4047 2836 4113 2844
rect 4927 2836 6153 2844
rect 7207 2836 7233 2844
rect 7607 2836 7833 2844
rect 7847 2836 8573 2844
rect 8587 2836 8653 2844
rect 9047 2836 9704 2844
rect 9696 2827 9704 2836
rect 11987 2836 12093 2844
rect 3096 2816 3464 2824
rect 3667 2816 3773 2824
rect 4187 2816 4293 2824
rect 4387 2816 4453 2824
rect 5047 2816 5693 2824
rect 5947 2816 6273 2824
rect 6347 2816 6773 2824
rect 9707 2816 9913 2824
rect 9927 2816 10713 2824
rect 10827 2816 10973 2824
rect 1267 2796 1393 2804
rect 1407 2796 1553 2804
rect 1567 2796 1953 2804
rect 2407 2796 2773 2804
rect 2887 2796 2973 2804
rect 4207 2796 4333 2804
rect 4427 2796 4473 2804
rect 4767 2796 4973 2804
rect 5227 2796 5293 2804
rect 5747 2796 5833 2804
rect 8027 2796 8253 2804
rect 9027 2796 9133 2804
rect 10447 2796 10493 2804
rect 11307 2796 11533 2804
rect 11547 2796 11693 2804
rect 187 2776 233 2784
rect 287 2779 333 2787
rect 527 2776 673 2784
rect 687 2776 713 2784
rect 1047 2776 1073 2784
rect 2007 2776 2053 2784
rect 2187 2776 2353 2784
rect 2647 2776 2793 2784
rect 2847 2776 3053 2784
rect 3447 2779 3653 2787
rect 3947 2779 4013 2787
rect 3027 2764 3040 2767
rect 3027 2753 3044 2764
rect 467 2733 493 2741
rect 547 2736 913 2744
rect 927 2733 973 2741
rect 1327 2733 1353 2741
rect 1587 2736 1773 2744
rect 2467 2733 2613 2741
rect 2667 2733 2773 2741
rect 187 2716 253 2724
rect 267 2716 1133 2724
rect 1147 2716 1273 2724
rect 1287 2716 1373 2724
rect 2127 2716 2193 2724
rect 2956 2724 2964 2753
rect 3036 2744 3044 2753
rect 3367 2756 3433 2764
rect 3896 2764 3904 2776
rect 4127 2776 4213 2784
rect 4227 2779 4253 2787
rect 4367 2776 4433 2784
rect 4516 2764 4524 2776
rect 4707 2784 4720 2787
rect 4707 2773 4724 2784
rect 3896 2756 4204 2764
rect 4516 2756 4573 2764
rect 3036 2736 3073 2744
rect 3236 2744 3244 2750
rect 3236 2736 3633 2744
rect 3747 2736 3873 2744
rect 4196 2744 4204 2756
rect 4716 2744 4724 2773
rect 4776 2776 5033 2784
rect 4776 2744 4784 2776
rect 5187 2776 5313 2784
rect 5447 2776 5473 2784
rect 5487 2779 5553 2787
rect 5627 2776 5693 2784
rect 5787 2776 5853 2784
rect 5987 2779 6053 2787
rect 6107 2776 6212 2784
rect 6247 2776 6453 2784
rect 6467 2776 6633 2784
rect 6927 2776 7072 2784
rect 7107 2776 7153 2784
rect 7207 2779 7253 2787
rect 7367 2779 7393 2787
rect 7747 2779 7853 2787
rect 8307 2779 8393 2787
rect 8447 2776 8533 2784
rect 8927 2776 9073 2784
rect 9907 2776 10393 2784
rect 10687 2779 10733 2787
rect 10907 2779 10993 2787
rect 11147 2776 11193 2784
rect 11807 2779 12013 2787
rect 4207 2733 4253 2741
rect 4347 2733 4453 2741
rect 4716 2736 4733 2744
rect 4867 2733 5013 2741
rect 5067 2733 5113 2741
rect 5347 2733 5453 2741
rect 5507 2736 5573 2744
rect 6087 2733 6173 2741
rect 6367 2736 6653 2744
rect 7087 2736 7133 2744
rect 7147 2733 7213 2741
rect 7227 2736 7353 2744
rect 8036 2744 8044 2773
rect 8007 2736 8044 2744
rect 8087 2736 8273 2744
rect 8287 2733 8413 2741
rect 8567 2733 8613 2741
rect 9007 2733 9053 2741
rect 9787 2733 9873 2741
rect 10107 2736 10173 2744
rect 10467 2736 10533 2744
rect 10607 2736 10733 2744
rect 10987 2733 11173 2741
rect 11687 2736 12093 2744
rect 12107 2733 12253 2741
rect 2927 2716 2964 2724
rect 4127 2716 4153 2724
rect 4507 2716 4693 2724
rect 5307 2716 5893 2724
rect 6667 2716 6893 2724
rect 7767 2716 7833 2724
rect 9087 2716 9313 2724
rect 9487 2716 9633 2724
rect 227 2696 553 2704
rect 2387 2696 2893 2704
rect 4107 2696 4232 2704
rect 4267 2696 4873 2704
rect 5487 2696 5513 2704
rect 5687 2696 5853 2704
rect 6007 2696 6113 2704
rect 6567 2696 7033 2704
rect 7387 2696 7413 2704
rect 8247 2696 8433 2704
rect 9867 2696 10873 2704
rect 11227 2696 11493 2704
rect 1187 2676 1653 2684
rect 1707 2676 3453 2684
rect 3567 2676 3633 2684
rect 4207 2676 4333 2684
rect 4767 2676 4833 2684
rect 5267 2676 5973 2684
rect 6407 2676 6553 2684
rect 6567 2676 6613 2684
rect 7187 2676 7293 2684
rect 7307 2676 8073 2684
rect 8527 2676 8733 2684
rect 8747 2676 9073 2684
rect 567 2656 1893 2664
rect 3007 2656 3473 2664
rect 3987 2656 4913 2664
rect 5807 2656 6233 2664
rect 6247 2656 6293 2664
rect 6527 2656 6833 2664
rect 7107 2656 7453 2664
rect 7807 2656 8773 2664
rect 8987 2656 9093 2664
rect 10636 2656 10884 2664
rect 547 2636 1993 2644
rect 3787 2636 4233 2644
rect 4247 2636 4513 2644
rect 4947 2636 5673 2644
rect 5767 2636 6433 2644
rect 6447 2636 7073 2644
rect 8087 2636 8713 2644
rect 10636 2644 10644 2656
rect 10427 2636 10644 2644
rect 10876 2644 10884 2656
rect 10927 2656 11713 2664
rect 10876 2636 11673 2644
rect 11776 2636 11973 2644
rect 1167 2616 1353 2624
rect 1367 2616 1833 2624
rect 1847 2616 2313 2624
rect 2327 2616 3033 2624
rect 3047 2616 3433 2624
rect 5007 2616 5213 2624
rect 5507 2616 6413 2624
rect 7727 2616 9504 2624
rect 1667 2596 1813 2604
rect 1987 2596 2333 2604
rect 4047 2596 4413 2604
rect 4627 2596 4933 2604
rect 6027 2596 6173 2604
rect 7027 2596 7433 2604
rect 9496 2604 9504 2616
rect 9567 2616 10853 2624
rect 11776 2624 11784 2636
rect 11367 2616 11784 2624
rect 9496 2596 9913 2604
rect 9927 2596 10653 2604
rect 10827 2596 11313 2604
rect 11327 2596 11793 2604
rect 4787 2576 5153 2584
rect 5227 2576 5533 2584
rect 5927 2576 6993 2584
rect 7047 2576 7853 2584
rect 8167 2576 8413 2584
rect 9267 2576 9353 2584
rect 9367 2576 9473 2584
rect 10967 2576 11133 2584
rect 11147 2576 11213 2584
rect 2027 2556 2143 2564
rect 227 2536 433 2544
rect 447 2536 813 2544
rect 2135 2507 2143 2556
rect 2867 2556 3633 2564
rect 3827 2556 4073 2564
rect 4187 2556 4293 2564
rect 5087 2556 5193 2564
rect 5867 2556 6013 2564
rect 6147 2556 6353 2564
rect 7107 2556 7633 2564
rect 7887 2556 8753 2564
rect 9167 2556 9633 2564
rect 10267 2556 10373 2564
rect 11287 2556 11313 2564
rect 11727 2556 11773 2564
rect 2227 2536 2604 2544
rect 267 2496 293 2504
rect 307 2496 893 2504
rect 1667 2496 1693 2504
rect 1767 2504 1780 2507
rect 1767 2493 1784 2504
rect 507 2476 613 2484
rect 927 2479 993 2487
rect 1067 2479 1253 2487
rect 196 2447 204 2473
rect 1227 2456 1373 2464
rect 1776 2464 1784 2493
rect 1856 2493 1857 2504
rect 2167 2496 2233 2504
rect 1856 2464 1864 2493
rect 747 2436 913 2444
rect 1027 2436 1053 2444
rect 1516 2444 1524 2456
rect 1856 2456 1873 2464
rect 2007 2459 2173 2467
rect 2276 2467 2284 2493
rect 2336 2467 2344 2493
rect 2596 2487 2604 2536
rect 2887 2536 3073 2544
rect 4027 2536 4273 2544
rect 4287 2536 4553 2544
rect 6427 2536 6993 2544
rect 7927 2536 8533 2544
rect 8547 2536 8733 2544
rect 9067 2536 9893 2544
rect 11007 2536 11133 2544
rect 11367 2536 12053 2544
rect 2716 2516 3353 2524
rect 2716 2507 2724 2516
rect 3567 2516 3933 2524
rect 3947 2516 3993 2524
rect 4587 2516 4653 2524
rect 5207 2516 5233 2524
rect 5727 2516 5933 2524
rect 6527 2516 7013 2524
rect 7147 2516 7233 2524
rect 7767 2516 8324 2524
rect 2647 2496 2713 2504
rect 5187 2504 5200 2507
rect 5187 2493 5204 2504
rect 5507 2496 5533 2504
rect 5647 2496 5713 2504
rect 2596 2476 2613 2487
rect 2600 2473 2613 2476
rect 2907 2476 2972 2484
rect 3727 2479 3793 2487
rect 3927 2479 3993 2487
rect 4096 2476 4273 2484
rect 4627 2479 4673 2487
rect 2387 2459 2473 2467
rect 2647 2453 2673 2461
rect 2993 2464 3007 2473
rect 2767 2460 3007 2464
rect 2767 2456 3004 2460
rect 4096 2464 4104 2476
rect 4727 2476 4813 2484
rect 4880 2484 4893 2487
rect 4876 2473 4893 2484
rect 5047 2479 5113 2487
rect 1407 2436 1524 2444
rect 2636 2444 2644 2450
rect 2227 2436 2644 2444
rect 2747 2436 2953 2444
rect 987 2416 1073 2424
rect 1327 2416 1373 2424
rect 1387 2416 1653 2424
rect 2147 2416 2193 2424
rect 3196 2424 3204 2456
rect 3467 2453 3553 2461
rect 4016 2456 4104 2464
rect 3367 2436 3393 2444
rect 4016 2444 4024 2456
rect 4876 2464 4884 2473
rect 4807 2456 4884 2464
rect 5196 2447 5204 2493
rect 6207 2496 6413 2504
rect 7527 2496 7553 2504
rect 8316 2504 8324 2516
rect 9007 2516 10413 2524
rect 10527 2516 10653 2524
rect 10667 2516 10813 2524
rect 11507 2516 11653 2524
rect 11667 2516 12013 2524
rect 8316 2496 8433 2504
rect 8887 2496 9093 2504
rect 9447 2496 10693 2504
rect 11967 2496 11993 2504
rect 5787 2479 6093 2487
rect 6647 2476 6733 2484
rect 6747 2476 6953 2484
rect 7227 2476 7293 2484
rect 7347 2476 7473 2484
rect 7967 2476 8013 2484
rect 8067 2476 8173 2484
rect 8187 2479 8253 2487
rect 8587 2479 9053 2487
rect 9607 2476 9713 2484
rect 10147 2476 10213 2484
rect 10227 2476 10373 2484
rect 10427 2479 10473 2487
rect 10707 2479 10793 2487
rect 11007 2476 11173 2484
rect 11187 2476 11273 2484
rect 11467 2479 11753 2487
rect 11807 2476 11933 2484
rect 4527 2433 4593 2441
rect 4667 2436 4893 2444
rect 5356 2444 5364 2456
rect 5507 2453 5553 2461
rect 5807 2456 6513 2464
rect 5356 2436 5573 2444
rect 5887 2433 5913 2441
rect 6247 2433 6393 2441
rect 6787 2433 6913 2441
rect 7147 2433 7173 2441
rect 7787 2436 7933 2444
rect 7947 2433 7993 2441
rect 9067 2433 9113 2441
rect 9247 2436 9373 2444
rect 9667 2433 9693 2441
rect 9987 2433 10113 2441
rect 10187 2436 10233 2444
rect 10247 2433 10353 2441
rect 10487 2436 10673 2444
rect 10907 2433 10933 2441
rect 11787 2436 11893 2444
rect 11967 2433 12013 2441
rect 12036 2427 12044 2476
rect 3196 2416 3453 2424
rect 3747 2416 3773 2424
rect 4167 2416 4253 2424
rect 5047 2416 6693 2424
rect 8587 2416 8813 2424
rect 9287 2416 9353 2424
rect 9627 2416 10013 2424
rect 11247 2416 11453 2424
rect 2373 2404 2387 2413
rect 2373 2400 2653 2404
rect 2376 2396 2653 2400
rect 2967 2396 4293 2404
rect 4487 2396 4873 2404
rect 5707 2396 6533 2404
rect 6827 2396 6933 2404
rect 6947 2396 7433 2404
rect 7507 2396 7913 2404
rect 8407 2396 8513 2404
rect 8527 2396 10173 2404
rect 10267 2396 10633 2404
rect 10847 2396 10973 2404
rect 11687 2396 11773 2404
rect 1287 2376 1393 2384
rect 5847 2376 5873 2384
rect 6147 2376 6313 2384
rect 6367 2376 6653 2384
rect 7267 2376 7453 2384
rect 7467 2376 8384 2384
rect 3007 2356 3973 2364
rect 5487 2356 5513 2364
rect 7487 2356 8273 2364
rect 8287 2356 8353 2364
rect 8376 2364 8384 2376
rect 8447 2376 8853 2384
rect 9507 2376 9873 2384
rect 9887 2376 10213 2384
rect 10287 2376 10513 2384
rect 11007 2376 11133 2384
rect 12067 2376 12173 2384
rect 8376 2356 8433 2364
rect 8607 2356 9953 2364
rect 10067 2356 10153 2364
rect 10207 2356 10613 2364
rect 11267 2356 11613 2364
rect 2507 2336 2753 2344
rect 2907 2336 2933 2344
rect 3507 2336 3913 2344
rect 4067 2336 4653 2344
rect 4667 2336 4733 2344
rect 6387 2336 6613 2344
rect 6627 2336 6713 2344
rect 7047 2336 7313 2344
rect 8047 2336 8553 2344
rect 9467 2336 9973 2344
rect 10227 2336 10913 2344
rect 10936 2336 11493 2344
rect 267 2316 1153 2324
rect 1727 2316 2053 2324
rect 2347 2316 2473 2324
rect 2936 2324 2944 2333
rect 2936 2316 3624 2324
rect 687 2296 853 2304
rect 1527 2296 1613 2304
rect 2527 2296 2632 2304
rect 2667 2296 2893 2304
rect 3616 2304 3624 2316
rect 3647 2316 4293 2324
rect 4927 2316 4993 2324
rect 5467 2316 5613 2324
rect 5687 2316 6113 2324
rect 6127 2316 6813 2324
rect 7167 2316 7433 2324
rect 8687 2316 10184 2324
rect 3616 2296 4473 2304
rect 4767 2296 4993 2304
rect 5047 2296 5793 2304
rect 5987 2296 7113 2304
rect 7667 2296 7733 2304
rect 7807 2296 8273 2304
rect 9627 2296 9853 2304
rect 10176 2304 10184 2316
rect 10936 2324 10944 2336
rect 10647 2316 10944 2324
rect 10176 2296 10593 2304
rect 10847 2296 10953 2304
rect 11087 2296 11493 2304
rect 11747 2296 11973 2304
rect 1147 2276 1353 2284
rect 1367 2276 1433 2284
rect 2307 2276 2353 2284
rect 2727 2276 2873 2284
rect 2927 2276 2973 2284
rect 3347 2276 3513 2284
rect 4647 2276 4773 2284
rect 5627 2276 5753 2284
rect 9427 2276 9933 2284
rect 10747 2276 10873 2284
rect 10887 2276 11373 2284
rect 11727 2276 11813 2284
rect 407 2256 513 2264
rect 667 2256 813 2264
rect 836 2256 1093 2264
rect 1427 2259 1573 2267
rect 1587 2256 1673 2264
rect 196 2227 204 2253
rect 836 2244 844 2256
rect 2067 2256 2213 2264
rect 2407 2256 2593 2264
rect 3207 2259 3233 2267
rect 3507 2259 3553 2267
rect 3627 2256 3693 2264
rect 3807 2256 3953 2264
rect 4007 2259 4033 2267
rect 4107 2256 4233 2264
rect 4276 2256 4513 2264
rect 5027 2259 5073 2267
rect 5307 2256 5433 2264
rect 576 2236 844 2244
rect 1696 2236 1733 2244
rect 287 2213 333 2221
rect 576 2224 584 2236
rect 347 2213 453 2221
rect 807 2213 833 2221
rect 1447 2213 1593 2221
rect 1696 2224 1704 2236
rect 1867 2233 2013 2241
rect 2127 2239 2153 2247
rect 4276 2244 4284 2256
rect 5507 2259 5533 2267
rect 5787 2256 5833 2264
rect 6067 2266 6224 2267
rect 6067 2259 6213 2266
rect 6287 2256 6333 2264
rect 6667 2256 6693 2264
rect 6927 2259 7173 2267
rect 7487 2256 7693 2264
rect 7747 2259 7893 2267
rect 8007 2259 8213 2267
rect 8547 2259 8593 2267
rect 8847 2256 8953 2264
rect 8967 2256 9093 2264
rect 9807 2259 9833 2267
rect 10207 2259 10253 2267
rect 10387 2259 10433 2267
rect 10567 2259 10673 2267
rect 11047 2259 11153 2267
rect 11287 2256 11333 2264
rect 11467 2256 11613 2264
rect 4127 2236 4284 2244
rect 7953 2244 7967 2253
rect 7953 2240 8044 2244
rect 7956 2236 8044 2240
rect 1667 2216 1704 2224
rect 2627 2213 2793 2221
rect 2927 2216 2973 2224
rect 2987 2216 3153 2224
rect 3167 2216 3473 2224
rect 3567 2216 3713 2224
rect 4027 2213 4053 2221
rect 4547 2213 4573 2221
rect 5047 2216 5273 2224
rect 5447 2213 5553 2221
rect 5967 2216 6113 2224
rect 6867 2216 6913 2224
rect 8036 2224 8044 2236
rect 8447 2236 9733 2244
rect 10587 2236 11333 2244
rect 11696 2244 11704 2256
rect 11927 2258 12012 2266
rect 11647 2236 11704 2244
rect 7307 2213 7413 2221
rect 7727 2216 7973 2224
rect 8667 2216 9393 2224
rect 9527 2213 9593 2221
rect 9967 2216 10413 2224
rect 10727 2213 10833 2221
rect 10947 2216 11033 2224
rect 11387 2213 11473 2221
rect 11487 2216 11513 2224
rect 11527 2216 11593 2224
rect 12036 2224 12044 2253
rect 12007 2216 12044 2224
rect 627 2196 1073 2204
rect 1127 2196 1173 2204
rect 1187 2196 1373 2204
rect 2047 2196 3833 2204
rect 4087 2196 4253 2204
rect 4307 2196 4613 2204
rect 4707 2196 5293 2204
rect 5347 2196 5653 2204
rect 6367 2196 6593 2204
rect 8227 2196 8253 2204
rect 8867 2196 9413 2204
rect 9627 2196 9773 2204
rect 10007 2196 10533 2204
rect 10627 2196 10673 2204
rect 10687 2196 11233 2204
rect 547 2176 593 2184
rect 1076 2184 1084 2193
rect 1076 2176 1313 2184
rect 1647 2176 2393 2184
rect 3447 2176 3553 2184
rect 5327 2176 5753 2184
rect 6727 2176 7144 2184
rect 2627 2156 3793 2164
rect 3907 2156 4153 2164
rect 4227 2156 4664 2164
rect 547 2136 873 2144
rect 887 2136 1293 2144
rect 1307 2136 1513 2144
rect 2267 2136 3293 2144
rect 3307 2136 4353 2144
rect 4407 2136 4553 2144
rect 4656 2144 4664 2156
rect 4687 2156 5013 2164
rect 5227 2156 5473 2164
rect 5487 2156 5593 2164
rect 6347 2156 6393 2164
rect 6527 2156 6673 2164
rect 7136 2164 7144 2176
rect 7167 2176 7593 2184
rect 8207 2176 8293 2184
rect 8427 2176 8553 2184
rect 9087 2176 9513 2184
rect 9567 2176 9773 2184
rect 9787 2176 9853 2184
rect 9947 2176 11413 2184
rect 11627 2176 11913 2184
rect 7136 2156 7833 2164
rect 8187 2156 8273 2164
rect 8947 2156 9092 2164
rect 9127 2156 9373 2164
rect 9856 2164 9864 2173
rect 9856 2156 10172 2164
rect 10207 2156 10493 2164
rect 10507 2156 11213 2164
rect 11227 2156 11353 2164
rect 11407 2156 11473 2164
rect 11947 2156 12233 2164
rect 4656 2136 4693 2144
rect 4707 2136 4793 2144
rect 6336 2144 6344 2153
rect 4867 2136 6344 2144
rect 7627 2136 7773 2144
rect 8707 2136 8873 2144
rect 9187 2136 9653 2144
rect 10827 2136 11173 2144
rect 1807 2116 2013 2124
rect 2787 2116 3313 2124
rect 3507 2116 3773 2124
rect 3787 2116 5093 2124
rect 5107 2116 6613 2124
rect 6847 2116 6953 2124
rect 7127 2116 7384 2124
rect 7376 2107 7384 2116
rect 8147 2116 8193 2124
rect 8207 2116 8613 2124
rect 8627 2116 10193 2124
rect 10327 2116 10633 2124
rect 11327 2116 11733 2124
rect 507 2096 593 2104
rect 3847 2096 4393 2104
rect 4547 2096 4633 2104
rect 5007 2096 5073 2104
rect 5087 2096 5513 2104
rect 5587 2096 5673 2104
rect 6827 2096 7133 2104
rect 7387 2096 8453 2104
rect 8476 2096 9173 2104
rect 1387 2076 2033 2084
rect 2887 2076 2913 2084
rect 4507 2076 4673 2084
rect 5387 2076 6273 2084
rect 6367 2076 6753 2084
rect 7467 2076 7604 2084
rect 987 2056 1353 2064
rect 3247 2056 3513 2064
rect 3607 2056 3773 2064
rect 4236 2056 4453 2064
rect 2047 2036 2544 2044
rect 2307 2016 2513 2024
rect 2536 2024 2544 2036
rect 4236 2044 4244 2056
rect 4767 2056 5133 2064
rect 6807 2056 6873 2064
rect 7596 2064 7604 2076
rect 7767 2076 7973 2084
rect 8476 2084 8484 2096
rect 9387 2096 9473 2104
rect 10867 2096 11293 2104
rect 7987 2076 8484 2084
rect 9267 2076 9633 2084
rect 9647 2076 9793 2084
rect 9807 2076 10033 2084
rect 10807 2076 10993 2084
rect 11007 2076 11753 2084
rect 7596 2056 8673 2064
rect 8807 2056 9013 2064
rect 3667 2036 4244 2044
rect 4567 2036 5684 2044
rect 5676 2027 5684 2036
rect 5947 2036 6053 2044
rect 6467 2036 6593 2044
rect 6607 2036 6753 2044
rect 6767 2036 7153 2044
rect 8167 2036 8253 2044
rect 8467 2036 8693 2044
rect 8767 2036 9173 2044
rect 9187 2036 9433 2044
rect 9656 2036 10533 2044
rect 2536 2016 2953 2024
rect 3207 2016 3473 2024
rect 4227 2016 4253 2024
rect 4307 2016 4533 2024
rect 4907 2016 5253 2024
rect 5687 2016 6033 2024
rect 6867 2016 7093 2024
rect 7867 2016 9073 2024
rect 9656 2024 9664 2036
rect 9227 2016 9664 2024
rect 9907 2016 10493 2024
rect 10827 2016 11153 2024
rect 207 1996 293 2004
rect 507 1996 573 2004
rect 707 1996 773 2004
rect 1207 1996 1373 2004
rect 1487 1996 1973 2004
rect 3187 1996 3533 2004
rect 4627 1996 5373 2004
rect 5867 1996 5993 2004
rect 6807 1996 7273 2004
rect 7347 1996 7713 2004
rect 10707 1996 10873 2004
rect 11367 1996 11753 2004
rect 12187 1996 12293 2004
rect 847 1979 1693 1987
rect 2847 1976 2932 1984
rect 2967 1976 3533 1984
rect 187 1959 213 1967
rect 236 1924 244 1973
rect 3593 1984 3607 1993
rect 3593 1980 3973 1984
rect 3596 1976 3973 1980
rect 4467 1976 4733 1984
rect 4747 1976 4773 1984
rect 9313 1984 9327 1993
rect 8716 1980 9327 1984
rect 8716 1976 9324 1980
rect 267 1959 393 1967
rect 1527 1959 1593 1967
rect 1967 1959 2073 1967
rect 2347 1959 2373 1967
rect 2487 1959 2573 1967
rect 2587 1956 2733 1964
rect 2807 1958 2833 1966
rect 3147 1959 3193 1967
rect 3467 1959 3573 1967
rect 4187 1959 4253 1967
rect 4847 1959 4933 1967
rect 5047 1959 5113 1967
rect 5167 1956 5413 1964
rect 5467 1956 5713 1964
rect 5787 1956 5933 1964
rect 5947 1959 6253 1967
rect 6267 1956 6413 1964
rect 6607 1959 6793 1967
rect 7007 1956 7084 1964
rect 1007 1939 1153 1947
rect 1267 1933 1313 1941
rect 3156 1936 3204 1944
rect 236 1916 273 1924
rect 647 1913 733 1921
rect 1507 1916 1952 1924
rect 1987 1913 2013 1921
rect 2067 1916 2173 1924
rect 2387 1913 2553 1921
rect 2607 1916 2793 1924
rect 2867 1916 2913 1924
rect 3156 1924 3164 1936
rect 3196 1924 3204 1936
rect 4407 1936 4753 1944
rect 7076 1944 7084 1956
rect 7307 1956 7333 1964
rect 7076 1936 7213 1944
rect 3196 1916 3433 1924
rect 3447 1913 3493 1921
rect 4087 1916 4273 1924
rect 5147 1913 5193 1921
rect 5347 1913 5393 1921
rect 5447 1913 5573 1921
rect 6107 1913 6193 1921
rect 6487 1913 6553 1921
rect 6627 1916 6773 1924
rect 6847 1916 7233 1924
rect 1687 1896 1753 1904
rect 2076 1896 2313 1904
rect 607 1876 753 1884
rect 2076 1884 2084 1896
rect 3187 1896 3233 1904
rect 3727 1896 3753 1904
rect 4027 1896 4053 1904
rect 4527 1896 4633 1904
rect 6096 1904 6104 1910
rect 7356 1907 7364 1973
rect 7467 1959 7573 1967
rect 7627 1959 7753 1967
rect 7767 1956 7793 1964
rect 8107 1956 8153 1964
rect 8167 1956 8313 1964
rect 8327 1959 8413 1967
rect 8436 1956 8453 1964
rect 8467 1959 8593 1967
rect 8716 1964 8724 1976
rect 10547 1976 10933 1984
rect 12047 1976 12133 1984
rect 8707 1956 8724 1964
rect 8827 1959 8973 1967
rect 9207 1959 9253 1967
rect 9307 1959 9353 1967
rect 7647 1916 7673 1924
rect 8436 1924 8444 1956
rect 9447 1956 9533 1964
rect 9727 1956 9813 1964
rect 9827 1959 9873 1967
rect 10087 1959 10113 1967
rect 10387 1959 10553 1967
rect 10576 1956 10653 1964
rect 8127 1916 8173 1924
rect 8227 1916 8444 1924
rect 8507 1916 8713 1924
rect 9087 1916 9273 1924
rect 9327 1913 9453 1921
rect 9667 1916 9793 1924
rect 9807 1916 9993 1924
rect 10576 1924 10584 1956
rect 10827 1958 10893 1966
rect 11047 1956 11113 1964
rect 11247 1956 11673 1964
rect 11927 1956 12013 1964
rect 12236 1927 12244 1956
rect 10107 1913 10293 1921
rect 10627 1913 10833 1921
rect 11307 1913 11393 1921
rect 11407 1916 11573 1924
rect 11667 1913 11713 1921
rect 12067 1916 12153 1924
rect 12236 1916 12253 1927
rect 12240 1913 12253 1916
rect 5927 1896 6104 1904
rect 6827 1896 7253 1904
rect 7347 1896 7364 1907
rect 7347 1893 7360 1896
rect 7847 1896 7873 1904
rect 9527 1896 9573 1904
rect 10347 1896 10593 1904
rect 10867 1896 10913 1904
rect 11767 1896 11933 1904
rect 1787 1876 2084 1884
rect 4456 1876 4493 1884
rect 207 1856 373 1864
rect 387 1856 553 1864
rect 827 1856 1393 1864
rect 2227 1856 2293 1864
rect 2307 1856 2993 1864
rect 4456 1864 4464 1876
rect 4827 1876 4893 1884
rect 7367 1876 7453 1884
rect 7607 1876 7673 1884
rect 7927 1876 7973 1884
rect 8027 1876 8093 1884
rect 8107 1876 8153 1884
rect 8587 1876 9173 1884
rect 10856 1884 10864 1892
rect 9947 1876 10864 1884
rect 11007 1876 12213 1884
rect 3807 1856 4464 1864
rect 6047 1856 6233 1864
rect 6387 1856 6833 1864
rect 6927 1856 7853 1864
rect 8727 1856 8833 1864
rect 9067 1856 9193 1864
rect 10067 1856 10793 1864
rect 11427 1856 11733 1864
rect 1007 1836 1293 1844
rect 2087 1836 2193 1844
rect 2867 1836 2933 1844
rect 3816 1836 4253 1844
rect 1667 1816 2153 1824
rect 2687 1816 2953 1824
rect 3816 1824 3824 1836
rect 4507 1836 4553 1844
rect 6947 1836 7053 1844
rect 8447 1836 9213 1844
rect 9607 1836 9893 1844
rect 10527 1836 10573 1844
rect 12107 1836 12273 1844
rect 3327 1816 3824 1824
rect 3847 1816 4413 1824
rect 4487 1816 5304 1824
rect 5296 1807 5304 1816
rect 6447 1816 6853 1824
rect 6867 1816 7013 1824
rect 7407 1816 7553 1824
rect 7567 1816 8193 1824
rect 9527 1816 9813 1824
rect 347 1796 513 1804
rect 587 1796 673 1804
rect 687 1796 1033 1804
rect 1047 1796 4993 1804
rect 5307 1796 6373 1804
rect 7147 1796 8653 1804
rect 8927 1796 9504 1804
rect 1687 1776 2132 1784
rect 2167 1776 3493 1784
rect 3787 1776 3953 1784
rect 4007 1776 4093 1784
rect 4327 1776 4413 1784
rect 4567 1776 4613 1784
rect 5107 1776 5273 1784
rect 5607 1776 5693 1784
rect 5807 1776 5953 1784
rect 6467 1776 6513 1784
rect 7167 1776 7593 1784
rect 8207 1776 8233 1784
rect 8307 1776 8433 1784
rect 9496 1784 9504 1796
rect 9687 1796 10133 1804
rect 10307 1796 10824 1804
rect 9496 1776 10113 1784
rect 10627 1776 10793 1784
rect 10816 1784 10824 1796
rect 11107 1796 11273 1804
rect 11347 1796 11453 1804
rect 11647 1796 11753 1804
rect 10816 1776 11913 1784
rect 247 1756 313 1764
rect 507 1756 673 1764
rect 927 1756 1293 1764
rect 3547 1756 3653 1764
rect 4847 1756 5233 1764
rect 5356 1756 5493 1764
rect 256 1736 293 1744
rect 256 1704 264 1736
rect 1276 1737 1633 1744
rect 5356 1750 5364 1756
rect 8907 1756 8993 1764
rect 9087 1756 9473 1764
rect 10947 1756 11133 1764
rect 11967 1756 12073 1764
rect 1276 1736 1644 1737
rect 1887 1736 2053 1744
rect 167 1693 213 1701
rect 527 1696 553 1704
rect 1276 1704 1284 1736
rect 2187 1739 2233 1747
rect 2627 1736 2713 1744
rect 2927 1736 3233 1744
rect 3707 1739 3733 1747
rect 3776 1736 4093 1744
rect 4307 1739 4353 1747
rect 4607 1746 4664 1747
rect 4607 1739 4653 1746
rect 3776 1724 3784 1736
rect 3756 1716 3784 1724
rect 1327 1696 1533 1704
rect 1547 1696 1853 1704
rect 1867 1696 1953 1704
rect 2067 1693 2113 1701
rect 2247 1696 2393 1704
rect 2987 1693 3013 1701
rect 3027 1693 3113 1701
rect 3407 1693 3473 1701
rect 3756 1704 3764 1716
rect 4096 1704 4104 1736
rect 4767 1739 4793 1747
rect 4860 1744 4873 1747
rect 4856 1733 4873 1744
rect 5127 1736 5344 1744
rect 5376 1736 5393 1744
rect 5707 1739 5833 1747
rect 3667 1696 3764 1704
rect 3807 1693 3893 1701
rect 4007 1693 4033 1701
rect 4096 1696 4313 1704
rect 4327 1696 4513 1704
rect 4856 1704 4864 1733
rect 5336 1724 5344 1736
rect 5376 1724 5384 1736
rect 5907 1736 5953 1744
rect 6216 1736 6273 1744
rect 5336 1716 5384 1724
rect 6196 1724 6204 1736
rect 5527 1716 5664 1724
rect 6176 1720 6204 1724
rect 5656 1704 5664 1716
rect 6173 1716 6204 1720
rect 6173 1707 6187 1716
rect 5287 1693 5413 1701
rect 5607 1693 5633 1701
rect 5656 1696 5673 1704
rect 5727 1696 5933 1704
rect 6216 1704 6224 1736
rect 6527 1736 6753 1744
rect 6807 1739 6893 1747
rect 7647 1739 7713 1747
rect 8387 1739 8473 1747
rect 8527 1739 8753 1747
rect 8767 1736 8853 1744
rect 9487 1739 9633 1747
rect 9787 1736 9893 1744
rect 9967 1739 10033 1747
rect 10296 1736 10333 1744
rect 10767 1739 10893 1747
rect 9216 1716 9373 1724
rect 6327 1696 6853 1704
rect 6947 1693 7033 1701
rect 7867 1693 8053 1701
rect 9216 1704 9224 1716
rect 9796 1716 9933 1724
rect 8247 1696 8413 1704
rect 9796 1704 9804 1716
rect 10296 1724 10304 1736
rect 11187 1736 11353 1744
rect 11687 1739 11693 1747
rect 11707 1739 11733 1747
rect 12027 1739 12213 1747
rect 10007 1716 10304 1724
rect 9427 1696 9493 1704
rect 9507 1693 9673 1701
rect 10067 1696 10093 1704
rect 10327 1696 10373 1704
rect 10607 1696 10693 1704
rect 10807 1696 10833 1704
rect 10847 1696 11113 1704
rect 11767 1693 11973 1701
rect 12087 1693 12193 1701
rect 787 1676 813 1684
rect 2167 1676 2213 1684
rect 7227 1676 7333 1684
rect 7807 1676 8273 1684
rect 8287 1676 8393 1684
rect 8647 1676 8693 1684
rect 8747 1676 8913 1684
rect 8987 1676 9033 1684
rect 9547 1676 9593 1684
rect 10887 1676 10993 1684
rect 11007 1676 11053 1684
rect 11227 1676 11373 1684
rect 11667 1676 11713 1684
rect 367 1656 1193 1664
rect 2667 1656 3213 1664
rect 3227 1656 4584 1664
rect 4576 1647 4584 1656
rect 4827 1656 5153 1664
rect 5167 1656 5773 1664
rect 5947 1656 6313 1664
rect 6787 1656 7093 1664
rect 7187 1656 8893 1664
rect 8947 1656 9073 1664
rect 9187 1656 10553 1664
rect 10567 1656 11173 1664
rect 1547 1636 1693 1644
rect 2747 1636 3153 1644
rect 4587 1636 5073 1644
rect 5087 1636 5093 1644
rect 6147 1636 6233 1644
rect 6776 1644 6784 1653
rect 6607 1636 6784 1644
rect 6967 1636 7053 1644
rect 7307 1636 7633 1644
rect 7887 1636 8072 1644
rect 8107 1636 8972 1644
rect 9007 1636 9053 1644
rect 9227 1636 9833 1644
rect 9847 1636 9953 1644
rect 11467 1636 11913 1644
rect 2527 1616 2693 1624
rect 2707 1616 3833 1624
rect 4667 1616 4933 1624
rect 6687 1616 6753 1624
rect 7207 1616 7253 1624
rect 7267 1616 7913 1624
rect 7927 1616 8673 1624
rect 8687 1616 8813 1624
rect 8827 1616 8953 1624
rect 9267 1616 9353 1624
rect 9367 1616 9953 1624
rect 10127 1616 10353 1624
rect 1567 1596 2493 1604
rect 2987 1596 3513 1604
rect 5387 1596 5893 1604
rect 6167 1596 6724 1604
rect 2887 1576 3693 1584
rect 3767 1576 4093 1584
rect 4547 1576 4673 1584
rect 4687 1576 4813 1584
rect 5027 1576 5173 1584
rect 6127 1576 6353 1584
rect 6716 1584 6724 1596
rect 7367 1596 7453 1604
rect 7467 1596 7573 1604
rect 7587 1596 7853 1604
rect 8187 1596 8313 1604
rect 8467 1596 8793 1604
rect 8807 1596 9193 1604
rect 9647 1596 9693 1604
rect 9707 1596 10253 1604
rect 11347 1596 11473 1604
rect 11487 1596 11633 1604
rect 6716 1576 7293 1584
rect 7627 1576 8024 1584
rect 2907 1556 3393 1564
rect 4767 1556 5273 1564
rect 5847 1556 5973 1564
rect 5987 1556 6913 1564
rect 7027 1556 7353 1564
rect 8016 1564 8024 1576
rect 8367 1576 9573 1584
rect 9587 1576 10933 1584
rect 8016 1556 8213 1564
rect 8427 1556 8852 1564
rect 8887 1556 9493 1564
rect 9827 1556 9853 1564
rect 10267 1556 11593 1564
rect 3527 1536 4113 1544
rect 4267 1536 6553 1544
rect 6567 1536 7393 1544
rect 8007 1536 8613 1544
rect 8847 1536 9873 1544
rect 9887 1536 10093 1544
rect 10567 1536 10593 1544
rect 11947 1536 12013 1544
rect 2487 1516 2873 1524
rect 3047 1516 3333 1524
rect 4427 1516 4753 1524
rect 5467 1516 5873 1524
rect 5887 1516 6593 1524
rect 7207 1516 7893 1524
rect 8267 1516 8473 1524
rect 10147 1516 10793 1524
rect 10987 1516 11313 1524
rect 507 1496 613 1504
rect 627 1496 673 1504
rect 907 1496 1093 1504
rect 1147 1496 1213 1504
rect 1327 1496 1373 1504
rect 1907 1496 1993 1504
rect 2007 1496 2593 1504
rect 2607 1496 2933 1504
rect 3167 1496 3673 1504
rect 3687 1496 3753 1504
rect 4227 1496 4293 1504
rect 4307 1496 4904 1504
rect 4896 1487 4904 1496
rect 5327 1496 7153 1504
rect 7327 1496 7493 1504
rect 8607 1496 9473 1504
rect 11527 1496 12233 1504
rect 987 1476 1113 1484
rect 1287 1476 1713 1484
rect 2747 1476 2833 1484
rect 4267 1476 4473 1484
rect 4487 1476 4793 1484
rect 4907 1476 5133 1484
rect 5347 1476 5613 1484
rect 6607 1476 6853 1484
rect 7787 1476 7853 1484
rect 8147 1476 8512 1484
rect 8547 1476 10104 1484
rect 2267 1456 2373 1464
rect 3207 1459 3493 1467
rect 4527 1456 4753 1464
rect 5867 1456 5933 1464
rect 6107 1456 6133 1464
rect 7727 1456 7864 1464
rect 207 1438 333 1446
rect 767 1438 913 1446
rect 1087 1439 1173 1447
rect 1387 1436 1533 1444
rect 2067 1436 2233 1444
rect 2247 1436 2313 1444
rect 2647 1436 2973 1444
rect 3047 1436 3084 1444
rect 3807 1436 4033 1444
rect 4587 1439 4613 1447
rect 4847 1439 4973 1447
rect 5016 1436 5573 1444
rect 5587 1436 5733 1444
rect 2216 1416 2393 1424
rect 2216 1404 2224 1416
rect 3076 1424 3084 1436
rect 3167 1419 3333 1427
rect 5016 1427 5024 1436
rect 5787 1436 5813 1444
rect 5867 1436 5913 1444
rect 6647 1436 7113 1444
rect 7507 1439 7613 1447
rect 7856 1444 7864 1456
rect 9727 1456 9913 1464
rect 10096 1464 10104 1476
rect 11607 1476 11733 1484
rect 10096 1456 10233 1464
rect 11907 1456 12033 1464
rect 7856 1436 8533 1444
rect 8627 1439 8653 1447
rect 9167 1436 10413 1444
rect 11347 1439 11433 1447
rect 11447 1436 11493 1444
rect 11627 1439 11693 1447
rect 11747 1439 11793 1447
rect 3467 1416 3533 1424
rect 3947 1416 4433 1424
rect 5007 1416 5024 1427
rect 8833 1424 8847 1433
rect 8833 1420 9064 1424
rect 8836 1416 9067 1420
rect 5007 1413 5020 1416
rect 867 1392 893 1400
rect 1707 1396 1933 1404
rect 1987 1393 2053 1401
rect 2267 1393 2293 1401
rect 2467 1393 2513 1401
rect 2627 1393 2693 1401
rect 2887 1393 2953 1401
rect 3707 1393 3733 1401
rect 3907 1396 4133 1404
rect 4147 1396 4273 1404
rect 4527 1396 4633 1404
rect 4827 1393 4893 1401
rect 5047 1396 5093 1404
rect 5247 1393 5313 1401
rect 5807 1393 5833 1401
rect 6087 1396 6153 1404
rect 6627 1393 6973 1401
rect 6987 1393 7033 1401
rect 7387 1393 7433 1401
rect 7587 1393 7733 1401
rect 8027 1396 8273 1404
rect 8287 1393 8353 1401
rect 8407 1396 8753 1404
rect 8856 1404 8864 1416
rect 8827 1396 8864 1404
rect 9053 1407 9067 1416
rect 11147 1416 11373 1424
rect 9447 1393 9593 1401
rect 10107 1393 10133 1401
rect 10407 1396 10653 1404
rect 11647 1393 11713 1401
rect 12047 1396 12093 1404
rect 12107 1396 12253 1404
rect 1007 1376 1053 1384
rect 1067 1376 1273 1384
rect 1287 1376 1353 1384
rect 1427 1376 1553 1384
rect 1667 1376 1753 1384
rect 3076 1376 3193 1384
rect 787 1356 973 1364
rect 1087 1356 1133 1364
rect 1227 1356 1433 1364
rect 3076 1364 3084 1376
rect 3467 1376 3573 1384
rect 9867 1376 10153 1384
rect 10167 1376 10213 1384
rect 10447 1376 10573 1384
rect 10807 1376 10953 1384
rect 10967 1376 11473 1384
rect 12187 1376 12233 1384
rect 2407 1356 3084 1364
rect 4027 1356 4553 1364
rect 4947 1356 5213 1364
rect 5227 1356 5584 1364
rect 1187 1336 1493 1344
rect 2047 1336 2273 1344
rect 2287 1336 3133 1344
rect 4647 1336 4693 1344
rect 4767 1336 5553 1344
rect 5576 1344 5584 1356
rect 6227 1356 6704 1364
rect 5576 1336 6173 1344
rect 6187 1336 6653 1344
rect 6696 1344 6704 1356
rect 6907 1356 7044 1364
rect 6696 1336 7013 1344
rect 7036 1344 7044 1356
rect 7347 1356 8153 1364
rect 8176 1356 8553 1364
rect 8176 1344 8184 1356
rect 8867 1356 9633 1364
rect 9907 1356 10104 1364
rect 7036 1336 8184 1344
rect 8227 1336 9153 1344
rect 10096 1344 10104 1356
rect 10667 1356 10853 1364
rect 10927 1356 11073 1364
rect 11087 1356 11433 1364
rect 11607 1356 11713 1364
rect 10096 1336 10253 1344
rect 707 1316 993 1324
rect 1527 1316 2993 1324
rect 3167 1316 3253 1324
rect 3687 1316 4873 1324
rect 7187 1316 7253 1324
rect 9767 1316 10473 1324
rect 10487 1316 11213 1324
rect 996 1296 1093 1304
rect 447 1256 513 1264
rect 207 1219 333 1227
rect 447 1224 460 1227
rect 447 1213 464 1224
rect 527 1219 553 1227
rect 727 1216 813 1224
rect 456 1184 464 1213
rect 996 1204 1004 1296
rect 4707 1296 4913 1304
rect 4967 1296 5693 1304
rect 6307 1296 6913 1304
rect 6927 1296 7073 1304
rect 7407 1296 7713 1304
rect 7987 1296 8913 1304
rect 9627 1296 11173 1304
rect 11187 1296 11373 1304
rect 3087 1276 4033 1284
rect 4127 1276 5033 1284
rect 5087 1276 5313 1284
rect 6107 1276 6133 1284
rect 6707 1276 6873 1284
rect 7487 1276 7573 1284
rect 7587 1276 7673 1284
rect 8707 1276 8813 1284
rect 9927 1276 10433 1284
rect 11447 1276 11653 1284
rect 11927 1276 12173 1284
rect 1927 1256 2033 1264
rect 2627 1256 2693 1264
rect 3347 1256 3553 1264
rect 4287 1256 5533 1264
rect 6007 1256 6893 1264
rect 6947 1256 7513 1264
rect 7747 1256 8713 1264
rect 9167 1256 9333 1264
rect 9347 1256 9613 1264
rect 10407 1256 10433 1264
rect 10587 1256 10693 1264
rect 10887 1256 10953 1264
rect 4167 1236 5184 1244
rect 1987 1216 2073 1224
rect 2087 1219 2193 1227
rect 2747 1216 2933 1224
rect 3007 1216 3053 1224
rect 3127 1219 3293 1227
rect 3607 1220 4113 1228
rect 4296 1216 4313 1224
rect 4567 1219 4633 1227
rect 1256 1184 1264 1196
rect 1547 1204 1560 1207
rect 4276 1204 4284 1216
rect 1547 1193 1564 1204
rect 167 1176 213 1184
rect 1256 1176 1473 1184
rect 347 1156 753 1164
rect 1556 1164 1564 1193
rect 4096 1196 4284 1204
rect 1716 1184 1724 1190
rect 1716 1176 1873 1184
rect 2467 1176 2613 1184
rect 4096 1184 4104 1196
rect 2847 1173 2973 1181
rect 3027 1173 3073 1181
rect 3287 1173 3333 1181
rect 4067 1176 4104 1184
rect 4296 1184 4304 1216
rect 4747 1216 5113 1224
rect 5176 1224 5184 1236
rect 5527 1236 5593 1244
rect 6427 1236 6593 1244
rect 6867 1236 7104 1244
rect 5176 1216 5453 1224
rect 5547 1219 5813 1227
rect 5867 1216 6013 1224
rect 6147 1216 6313 1224
rect 6387 1219 6573 1227
rect 6927 1219 6973 1227
rect 4676 1196 4693 1204
rect 4127 1176 4304 1184
rect 4347 1173 4393 1181
rect 4676 1167 4684 1196
rect 4907 1193 5073 1201
rect 5347 1173 5373 1181
rect 5527 1173 5553 1181
rect 6347 1176 6393 1184
rect 6696 1167 6704 1216
rect 7027 1216 7073 1224
rect 7096 1224 7104 1236
rect 7147 1236 7253 1244
rect 7787 1236 7913 1244
rect 10167 1236 11173 1244
rect 11487 1236 11933 1244
rect 7096 1216 7473 1224
rect 7487 1219 7593 1227
rect 7607 1216 7733 1224
rect 7827 1216 7893 1224
rect 7967 1216 8073 1224
rect 8167 1219 8293 1227
rect 8607 1216 8773 1224
rect 8827 1219 8933 1227
rect 9227 1216 9373 1224
rect 9847 1219 9873 1227
rect 10187 1219 10253 1227
rect 10347 1219 10393 1227
rect 10667 1216 10913 1224
rect 10927 1219 11073 1227
rect 11187 1216 11333 1224
rect 9836 1204 9844 1216
rect 10136 1204 10144 1216
rect 11347 1216 11473 1224
rect 11767 1216 12033 1224
rect 7796 1200 7844 1204
rect 7796 1196 7847 1200
rect 9836 1196 10144 1204
rect 6907 1173 6953 1181
rect 7127 1173 7193 1181
rect 7207 1176 7453 1184
rect 7796 1184 7804 1196
rect 7833 1187 7847 1196
rect 7547 1173 7573 1181
rect 7947 1176 8053 1184
rect 8107 1173 8453 1181
rect 8527 1176 8553 1184
rect 8787 1173 8873 1181
rect 8967 1176 9093 1184
rect 9987 1176 10153 1184
rect 10247 1176 10413 1184
rect 10507 1176 10673 1184
rect 10947 1176 11133 1184
rect 11156 1176 11193 1184
rect 3647 1156 3813 1164
rect 4427 1156 4573 1164
rect 5747 1156 5793 1164
rect 5807 1156 5833 1164
rect 5887 1156 5913 1164
rect 7827 1156 7873 1164
rect 9827 1156 9913 1164
rect 11156 1164 11164 1176
rect 11387 1173 11453 1181
rect 11667 1173 11693 1181
rect 12007 1173 12033 1181
rect 12047 1176 12213 1184
rect 11007 1156 11164 1164
rect 427 1136 493 1144
rect 2167 1136 2713 1144
rect 2947 1136 3473 1144
rect 3827 1136 3873 1144
rect 5187 1136 5333 1144
rect 5347 1136 6633 1144
rect 6687 1136 7053 1144
rect 7107 1136 7553 1144
rect 7796 1136 8833 1144
rect 7796 1127 7804 1136
rect 8947 1136 9093 1144
rect 9207 1136 9393 1144
rect 9407 1136 9893 1144
rect 10267 1136 10873 1144
rect 11227 1136 11613 1144
rect 11807 1136 11953 1144
rect 707 1116 793 1124
rect 1267 1116 1293 1124
rect 2547 1116 3313 1124
rect 3327 1116 4293 1124
rect 4307 1116 5013 1124
rect 5607 1116 5893 1124
rect 6827 1116 7793 1124
rect 7987 1116 8733 1124
rect 10367 1116 10693 1124
rect 11407 1116 11633 1124
rect 5596 1104 5604 1113
rect 5307 1096 5604 1104
rect 6727 1096 6753 1104
rect 6767 1096 6993 1104
rect 7167 1096 7473 1104
rect 7487 1096 7493 1104
rect 9367 1096 9433 1104
rect 9447 1096 9653 1104
rect 9967 1096 11213 1104
rect 47 1076 513 1084
rect 527 1076 833 1084
rect 847 1076 1553 1084
rect 1567 1076 2393 1084
rect 5007 1076 5153 1084
rect 5627 1076 6213 1084
rect 7047 1076 7953 1084
rect 8227 1076 8373 1084
rect 8387 1076 8573 1084
rect 8667 1076 9213 1084
rect 10747 1076 10953 1084
rect 3807 1056 4093 1064
rect 4107 1056 6473 1064
rect 6487 1056 6733 1064
rect 6747 1056 7073 1064
rect 7367 1056 7973 1064
rect 8727 1056 9193 1064
rect 9487 1056 10173 1064
rect 10267 1056 10293 1064
rect 647 1036 2513 1044
rect 4747 1036 4773 1044
rect 5027 1036 5593 1044
rect 6167 1036 6193 1044
rect 7247 1036 7873 1044
rect 8067 1036 8213 1044
rect 8347 1036 8413 1044
rect 8747 1036 9293 1044
rect 11827 1036 12193 1044
rect 2867 1016 2993 1024
rect 3007 1016 3033 1024
rect 3047 1016 3853 1024
rect 5127 1016 5813 1024
rect 6327 1016 7013 1024
rect 7067 1016 7913 1024
rect 9207 1016 9673 1024
rect 11327 1016 11973 1024
rect 1367 996 1453 1004
rect 1467 996 1633 1004
rect 1647 996 1993 1004
rect 2127 996 2193 1004
rect 2207 996 2573 1004
rect 2787 996 3133 1004
rect 4067 996 4213 1004
rect 4487 996 4593 1004
rect 4736 996 5233 1004
rect 1847 976 1873 984
rect 2807 976 2853 984
rect 3787 976 4253 984
rect 4736 984 4744 996
rect 5247 996 5613 1004
rect 5907 996 6113 1004
rect 6127 996 6153 1004
rect 7607 996 7813 1004
rect 8587 996 9033 1004
rect 11567 996 11933 1004
rect 4547 976 4744 984
rect 5147 976 5393 984
rect 5407 976 6273 984
rect 6287 976 6773 984
rect 7027 976 7232 984
rect 7267 976 7293 984
rect 9147 976 9233 984
rect 9247 976 9633 984
rect 10387 976 10473 984
rect 11587 976 11813 984
rect 1007 956 2153 964
rect 2216 956 3253 964
rect 2216 947 2224 956
rect 3367 956 3613 964
rect 5667 956 5993 964
rect 6967 956 7573 964
rect 7887 956 8093 964
rect 8427 956 8513 964
rect 8647 956 9973 964
rect 10367 956 10793 964
rect 10927 956 12073 964
rect 56 933 57 944
rect 196 936 373 944
rect 56 904 64 933
rect 196 910 204 936
rect 1947 936 2213 944
rect 2727 936 2773 944
rect 4107 936 4173 944
rect 4227 936 4273 944
rect 7727 936 7893 944
rect 8927 936 9213 944
rect 56 896 73 904
rect 467 893 613 901
rect 367 876 393 884
rect 696 867 704 916
rect 1067 916 1333 924
rect 1347 919 1593 927
rect 1907 919 2093 927
rect 2347 918 2433 926
rect 2827 919 2873 927
rect 2987 919 3073 927
rect 3087 916 3113 924
rect 3607 919 3673 927
rect 3727 916 3893 924
rect 3907 919 4293 927
rect 4447 916 4653 924
rect 4787 916 4833 924
rect 5187 919 5253 927
rect 5547 919 5573 927
rect 6027 919 6113 927
rect 6327 916 6393 924
rect 6607 919 6633 927
rect 6827 916 6933 924
rect 7007 918 7132 926
rect 7167 916 7293 924
rect 7467 919 7613 927
rect 8107 916 8264 924
rect 8256 910 8264 916
rect 10407 919 10433 927
rect 5776 896 6253 904
rect 807 876 973 884
rect 987 873 1053 881
rect 1627 876 1873 884
rect 1967 873 1993 881
rect 2107 876 2213 884
rect 2887 876 3053 884
rect 3267 873 3293 881
rect 3307 876 3573 884
rect 3927 876 4193 884
rect 4287 876 4453 884
rect 4507 873 4533 881
rect 4667 873 4753 881
rect 5776 884 5784 896
rect 7787 893 7993 901
rect 8387 896 8493 904
rect 8736 904 8744 915
rect 8736 896 8813 904
rect 9356 904 9364 915
rect 11167 916 11253 924
rect 11407 919 11453 927
rect 11687 919 11713 927
rect 8827 896 9364 904
rect 4827 876 5013 884
rect 5296 876 5313 884
rect 996 856 2073 864
rect 567 836 753 844
rect 996 844 1004 856
rect 2536 856 2713 864
rect 767 836 1004 844
rect 1847 836 1913 844
rect 2536 844 2544 856
rect 5296 864 5304 876
rect 5647 873 5773 881
rect 5827 873 5853 881
rect 6147 876 6193 884
rect 6467 876 6853 884
rect 7267 872 7333 880
rect 7647 873 7713 881
rect 8427 876 8453 884
rect 9667 876 10353 884
rect 10467 876 10573 884
rect 10587 876 10673 884
rect 10867 876 10973 884
rect 10987 876 11473 884
rect 12047 873 12073 881
rect 12087 876 12233 884
rect 3967 856 5304 864
rect 6267 856 6733 864
rect 6787 856 7393 864
rect 7407 856 7953 864
rect 8727 856 8833 864
rect 9347 856 9613 864
rect 9627 856 9733 864
rect 10507 856 11673 864
rect 11827 856 11993 864
rect 2507 836 2544 844
rect 2587 836 3333 844
rect 3887 836 5033 844
rect 6047 836 6373 844
rect 6567 836 7033 844
rect 7847 836 8053 844
rect 10727 836 11233 844
rect 11807 836 12073 844
rect 2187 816 2553 824
rect 2567 816 3004 824
rect 667 796 1053 804
rect 1067 796 1293 804
rect 1367 796 1573 804
rect 1587 796 2033 804
rect 2087 796 2753 804
rect 2767 796 2973 804
rect 2996 804 3004 816
rect 4307 816 5533 824
rect 5547 816 7153 824
rect 7176 816 7673 824
rect 2996 796 4153 804
rect 6527 796 6673 804
rect 6887 796 6972 804
rect 7176 804 7184 816
rect 8447 816 8513 824
rect 8987 816 9573 824
rect 9947 816 10033 824
rect 10047 816 10153 824
rect 10167 816 10333 824
rect 11187 816 11473 824
rect 11647 816 11733 824
rect 7007 796 7184 804
rect 7947 796 8493 804
rect 10627 796 11333 804
rect 2167 776 2633 784
rect 3127 776 3713 784
rect 5287 776 5393 784
rect 5927 776 6293 784
rect 6547 776 6753 784
rect 7967 776 8453 784
rect 8547 776 8773 784
rect 8787 776 9053 784
rect 9067 776 9393 784
rect 9407 776 9833 784
rect 9847 776 9893 784
rect 9987 776 10213 784
rect 10227 776 10624 784
rect 1027 756 1073 764
rect 2907 756 3213 764
rect 3227 756 3873 764
rect 5767 756 5893 764
rect 7807 756 7993 764
rect 8607 756 8933 764
rect 10616 764 10624 776
rect 11267 776 11553 784
rect 11567 776 12093 784
rect 10616 756 10813 764
rect 10827 756 11073 764
rect 11347 756 11793 764
rect 387 736 713 744
rect 1007 736 1533 744
rect 1867 736 2373 744
rect 2387 736 2773 744
rect 2916 736 3113 744
rect 1307 716 1493 724
rect 2087 716 2113 724
rect 196 696 373 704
rect 56 676 73 684
rect 196 684 204 696
rect 467 696 633 704
rect 1587 696 1753 704
rect 1807 696 2533 704
rect 2547 699 2593 707
rect 2647 699 2693 707
rect 56 647 64 676
rect 647 653 673 661
rect 1527 656 1773 664
rect 2107 653 2173 661
rect 2367 656 2613 664
rect 2787 653 2853 661
rect 2916 664 2924 736
rect 3747 736 4313 744
rect 4527 736 4973 744
rect 5127 736 5293 744
rect 5587 736 6233 744
rect 6307 736 6813 744
rect 6947 736 7213 744
rect 7267 736 7653 744
rect 7887 736 8293 744
rect 8316 736 9473 744
rect 5027 716 5453 724
rect 6787 716 6833 724
rect 8316 724 8324 736
rect 10247 736 11313 744
rect 7747 716 8324 724
rect 9527 716 9693 724
rect 10947 716 11113 724
rect 11127 716 11193 724
rect 11247 716 11393 724
rect 11867 716 11893 724
rect 2947 696 2964 704
rect 2956 667 2964 696
rect 2987 696 3173 704
rect 3647 699 3693 707
rect 3827 696 3993 704
rect 4387 699 4433 707
rect 4567 696 4593 704
rect 4927 700 5633 708
rect 5787 696 6273 704
rect 7147 699 7173 707
rect 7216 696 7873 704
rect 3716 676 3793 684
rect 2867 653 2873 661
rect 3127 653 3193 661
rect 3716 664 3724 676
rect 4127 676 5273 684
rect 6256 676 6653 684
rect 3387 656 3433 664
rect 3447 653 3613 661
rect 3767 653 3813 661
rect 4107 656 4273 664
rect 4347 654 4412 662
rect 4447 656 4633 664
rect 4947 654 5012 662
rect 5047 656 5213 664
rect 5227 656 5593 664
rect 6256 664 6264 676
rect 7216 684 7224 696
rect 7967 696 8033 704
rect 8347 699 8493 707
rect 8507 696 8553 704
rect 8707 707 9033 708
rect 8707 700 8733 707
rect 8747 700 8813 707
rect 8827 700 9033 707
rect 9287 696 9713 704
rect 10787 696 10893 704
rect 12007 696 12053 704
rect 7087 676 7224 684
rect 6487 653 6533 661
rect 6907 654 6993 662
rect 7196 664 7204 676
rect 9587 676 10613 684
rect 7507 653 7573 661
rect 7787 656 7813 664
rect 8467 656 8593 664
rect 9776 664 9784 676
rect 11007 679 11413 687
rect 11527 673 11673 681
rect 11807 676 11973 684
rect 9007 656 9433 664
rect 9447 653 9493 661
rect 10267 653 10313 661
rect 10327 656 10393 664
rect 10507 653 10573 661
rect 12076 664 12084 713
rect 10767 656 11093 664
rect 11267 653 11373 661
rect 56 636 57 647
rect 1027 636 1053 644
rect 4547 636 4613 644
rect 4847 636 6193 644
rect 6587 636 6753 644
rect 6767 636 7233 644
rect 7867 636 8053 644
rect 9047 636 9933 644
rect 9947 636 10933 644
rect 11967 636 12053 644
rect 1307 616 2053 624
rect 2067 616 2353 624
rect 2547 616 2973 624
rect 3147 616 3233 624
rect 3347 616 3473 624
rect 4867 616 5913 624
rect 6647 616 6793 624
rect 6807 616 7653 624
rect 7667 616 7893 624
rect 8367 616 8413 624
rect 8427 616 8993 624
rect 9207 616 9533 624
rect 9547 616 10193 624
rect 10207 616 10533 624
rect 47 596 513 604
rect 3627 596 4713 604
rect 4107 576 5073 584
rect 5087 576 5113 584
rect 5127 576 6273 584
rect 6287 576 6993 584
rect 8447 576 10873 584
rect 10887 576 11833 584
rect 11733 567 11747 576
rect 1787 556 2313 564
rect 2587 556 4853 564
rect 5287 556 6833 564
rect 8027 556 8473 564
rect 8487 556 8753 564
rect 8927 556 8953 564
rect 9027 556 10233 564
rect 11027 556 11333 564
rect 1807 536 2653 544
rect 2667 536 4113 544
rect 4307 536 5173 544
rect 7247 536 7933 544
rect 8507 536 9473 544
rect 5427 516 6453 524
rect 6696 516 7133 524
rect 147 496 353 504
rect 467 496 513 504
rect 1087 496 1233 504
rect 1827 496 2033 504
rect 2047 496 2573 504
rect 3787 496 3973 504
rect 3987 496 4293 504
rect 6696 504 6704 516
rect 10007 516 10273 524
rect 5847 496 6704 504
rect 6747 496 8313 504
rect 9787 476 10033 484
rect 10047 476 10213 484
rect 11287 476 11813 484
rect 707 456 1173 464
rect 1767 456 2073 464
rect 2087 456 2153 464
rect 2347 456 4493 464
rect 4547 456 4793 464
rect 5207 456 5613 464
rect 9827 456 10013 464
rect 10027 456 10373 464
rect 907 436 953 444
rect 1367 436 1513 444
rect 4587 436 4613 444
rect 5227 436 6313 444
rect 6607 436 6813 444
rect 6827 436 6933 444
rect 7007 436 8124 444
rect 1227 416 1273 424
rect 2207 416 2393 424
rect 8116 427 8124 436
rect 8487 436 8673 444
rect 8687 436 8913 444
rect 8967 436 9073 444
rect 9087 436 9193 444
rect 9427 436 9713 444
rect 11247 436 11413 444
rect 11427 436 11993 444
rect 12187 436 12253 444
rect 2707 416 2793 424
rect 4687 416 4744 424
rect 967 396 1352 404
rect 1387 396 1453 404
rect 2247 396 2333 404
rect 3067 396 3413 404
rect 3427 396 3633 404
rect 4187 396 4353 404
rect 4367 396 4513 404
rect 107 373 133 381
rect 307 379 392 387
rect 427 376 493 384
rect 1196 376 1604 384
rect 2567 379 2693 387
rect 1196 364 1204 376
rect 1596 364 1604 376
rect 3687 373 3773 381
rect 3947 379 4133 387
rect 4573 384 4587 393
rect 4636 384 4644 396
rect 4573 380 4624 384
rect 4576 376 4624 380
rect 4636 376 4713 384
rect 907 353 933 361
rect 987 356 1193 364
rect 1547 353 1573 361
rect 1596 356 2053 364
rect 2107 353 2233 361
rect 2287 356 2753 364
rect 2827 356 2993 364
rect 3007 353 3033 361
rect 4616 364 4624 376
rect 4736 384 4744 416
rect 8127 416 8433 424
rect 11207 416 11293 424
rect 11316 416 12193 424
rect 5387 396 5553 404
rect 5727 396 5893 404
rect 6107 399 6173 407
rect 7547 399 7913 407
rect 9187 399 9293 407
rect 4736 376 4753 384
rect 4807 379 4953 387
rect 5087 376 5153 384
rect 5936 384 5944 395
rect 5827 376 6053 384
rect 6216 384 6224 396
rect 9587 396 9773 404
rect 9967 399 9993 407
rect 10107 396 10753 404
rect 10807 396 11013 404
rect 11316 404 11324 416
rect 11147 396 11324 404
rect 11807 396 11973 404
rect 6147 376 6224 384
rect 6307 379 6433 387
rect 6887 376 7033 384
rect 8196 376 8273 384
rect 7156 364 7164 376
rect 3267 356 3293 364
rect 3427 353 3553 361
rect 4307 353 4333 361
rect 4616 356 4653 364
rect 5307 353 5333 361
rect 5667 353 5713 361
rect 6247 353 6593 361
rect 7116 356 7164 364
rect 407 336 753 344
rect 2367 336 3133 344
rect 6707 336 6733 344
rect 6747 336 6913 344
rect 1287 316 1773 324
rect 2767 316 3124 324
rect 1507 296 1753 304
rect 1807 296 2273 304
rect 3116 304 3124 316
rect 4567 316 4693 324
rect 5647 316 5753 324
rect 5767 316 5873 324
rect 5927 316 6093 324
rect 6207 316 6293 324
rect 7116 324 7124 356
rect 7427 356 7453 364
rect 7467 356 7633 364
rect 7867 353 7893 361
rect 7907 356 8013 364
rect 8196 364 8204 376
rect 8107 356 8204 364
rect 8707 353 8733 361
rect 8947 356 9133 364
rect 9947 356 10013 364
rect 10227 353 10273 361
rect 10387 353 10513 361
rect 10787 353 10813 361
rect 11007 356 11064 364
rect 9467 336 9533 344
rect 11056 344 11064 356
rect 11056 336 11313 344
rect 11327 336 11413 344
rect 11576 344 11584 376
rect 11707 376 11773 384
rect 11927 353 11993 361
rect 12187 356 12233 364
rect 11576 336 11793 344
rect 6687 316 7124 324
rect 7947 316 8093 324
rect 9107 316 9193 324
rect 9747 316 9813 324
rect 9907 316 10073 324
rect 10307 316 10733 324
rect 10747 316 10833 324
rect 10847 316 11033 324
rect 11187 316 11293 324
rect 11307 316 11373 324
rect 3116 296 3733 304
rect 4547 296 4613 304
rect 5567 296 5813 304
rect 6647 296 7353 304
rect 11107 296 12153 304
rect 47 276 193 284
rect 1896 276 2113 284
rect 1267 256 1733 264
rect 1896 264 1904 276
rect 2447 276 2493 284
rect 5556 284 5564 293
rect 4727 276 5564 284
rect 6707 276 6753 284
rect 7567 276 8273 284
rect 9307 276 10093 284
rect 11627 276 12313 284
rect 1747 256 1904 264
rect 2367 256 2593 264
rect 6527 256 6673 264
rect 6787 256 6993 264
rect 7667 256 7833 264
rect 7847 256 8073 264
rect 8087 256 8173 264
rect 11347 256 12333 264
rect 547 236 713 244
rect 767 236 1173 244
rect 2127 236 2773 244
rect 5927 236 5973 244
rect 10347 236 10993 244
rect 1347 216 1484 224
rect 1127 196 1373 204
rect 487 176 673 184
rect 727 179 813 187
rect 1047 176 1213 184
rect 1476 184 1484 216
rect 2027 216 2093 224
rect 3487 216 3913 224
rect 4087 216 5673 224
rect 5687 216 5833 224
rect 6567 216 6793 224
rect 10336 224 10344 233
rect 10127 216 10344 224
rect 3607 196 3633 204
rect 3647 196 3673 204
rect 5747 196 5793 204
rect 9227 196 9293 204
rect 10656 196 10893 204
rect 1476 176 1584 184
rect 2007 179 2053 187
rect 2107 176 2344 184
rect 2987 179 3053 187
rect 3867 176 4033 184
rect 1267 156 1453 164
rect 1576 164 1584 176
rect 2180 164 2193 167
rect 2176 153 2193 164
rect 2336 164 2344 176
rect 4247 179 4633 187
rect 4967 179 5193 187
rect 5356 176 5413 184
rect 227 136 733 144
rect 927 133 1053 141
rect 1276 140 1353 144
rect 1273 136 1353 140
rect 1273 127 1287 136
rect 2027 133 2073 141
rect 507 116 533 124
rect 2176 124 2184 153
rect 2547 159 2753 167
rect 5356 164 5364 176
rect 5487 176 5513 184
rect 5727 176 5953 184
rect 5967 176 6113 184
rect 6247 176 6453 184
rect 6476 176 6544 184
rect 4507 156 5364 164
rect 5436 156 5504 164
rect 5436 144 5444 156
rect 5496 144 5504 156
rect 6476 164 6484 176
rect 6147 156 6484 164
rect 2787 136 2833 144
rect 3687 133 3833 141
rect 3927 133 4153 141
rect 4167 136 4393 144
rect 5496 136 5633 144
rect 6256 144 6264 156
rect 6536 144 6544 176
rect 6727 176 6753 184
rect 7307 176 7344 184
rect 7336 164 7344 176
rect 7367 176 7653 184
rect 9547 179 9613 187
rect 10056 176 10112 184
rect 7336 156 7593 164
rect 7707 153 7853 161
rect 7987 156 8053 164
rect 8256 156 8473 164
rect 5747 133 5773 141
rect 6127 133 6213 141
rect 6467 133 6493 141
rect 8256 144 8264 156
rect 6707 136 6773 144
rect 7287 136 7513 144
rect 8307 136 8513 144
rect 8527 136 8733 144
rect 9007 133 9073 141
rect 9227 133 9253 141
rect 9307 136 9553 144
rect 9627 136 9793 144
rect 9807 136 9953 144
rect 10056 144 10064 176
rect 10147 176 10293 184
rect 10467 159 10493 167
rect 10656 164 10664 196
rect 11167 179 11373 187
rect 11687 176 11873 184
rect 12147 179 12173 187
rect 10787 156 10853 164
rect 10207 136 10313 144
rect 11047 133 11133 141
rect 11207 133 11353 141
rect 11647 133 11673 141
rect 11827 133 11853 141
rect 12067 136 12153 144
rect 1427 116 2173 124
rect 8027 113 8113 121
rect 9047 116 9293 124
rect 687 96 773 104
rect 827 96 1013 104
rect 1027 96 1113 104
rect 1747 96 2113 104
rect 2847 96 4073 104
rect 4247 96 4433 104
rect 5527 96 5693 104
rect 5707 96 5813 104
rect 9036 104 9044 113
rect 10827 113 10873 121
rect 11407 116 11953 124
rect 8787 96 9044 104
rect 11607 96 11813 104
rect 12047 96 12213 104
rect 4767 56 6633 64
rect 8187 56 10493 64
rect 10507 56 11293 64
rect 11907 56 12293 64
rect 1187 36 5573 44
rect 5467 16 5493 24
rect 5727 16 5793 24
rect 6727 16 6773 24
rect 7527 16 7553 24
rect 7567 16 7693 24
use INVX1  _1688_
timestamp 0
transform -1 0 1050 0 1 4430
box -6 -8 66 268
use NAND2X1  _1689_
timestamp 0
transform -1 0 530 0 1 4430
box -6 -8 86 268
use OAI21X1  _1690_
timestamp 0
transform -1 0 810 0 1 4430
box -6 -8 106 268
use INVX1  _1691_
timestamp 0
transform 1 0 190 0 -1 270
box -6 -8 66 268
use NAND2X1  _1692_
timestamp 0
transform -1 0 510 0 -1 270
box -6 -8 86 268
use OAI21X1  _1693_
timestamp 0
transform 1 0 710 0 -1 270
box -6 -8 106 268
use INVX8  _1694_
timestamp 0
transform -1 0 5790 0 1 4950
box -6 -8 126 268
use OR2X2  _1695_
timestamp 0
transform -1 0 550 0 -1 6510
box -6 -8 106 268
use OAI21X1  _1696_
timestamp 0
transform -1 0 550 0 1 6510
box -6 -8 106 268
use INVX1  _1697_
timestamp 0
transform -1 0 1630 0 1 7550
box -6 -8 66 268
use OR2X2  _1698_
timestamp 0
transform -1 0 3610 0 -1 3910
box -6 -8 106 268
use OAI21X1  _1699_
timestamp 0
transform 1 0 2970 0 -1 3910
box -6 -8 106 268
use INVX1  _1700_
timestamp 0
transform -1 0 4050 0 -1 7550
box -6 -8 66 268
use OR2X2  _1701_
timestamp 0
transform -1 0 790 0 -1 5470
box -6 -8 106 268
use OAI21X1  _1702_
timestamp 0
transform -1 0 790 0 1 5470
box -6 -8 106 268
use INVX1  _1703_
timestamp 0
transform 1 0 3350 0 -1 5470
box -6 -8 66 268
use OR2X2  _1704_
timestamp 0
transform -1 0 570 0 -1 4950
box -6 -8 106 268
use OAI21X1  _1705_
timestamp 0
transform 1 0 190 0 -1 4950
box -6 -8 106 268
use INVX1  _1706_
timestamp 0
transform -1 0 4010 0 1 5470
box -6 -8 66 268
use OR2X2  _1707_
timestamp 0
transform -1 0 830 0 1 5990
box -6 -8 106 268
use OAI21X1  _1708_
timestamp 0
transform 1 0 730 0 -1 6510
box -6 -8 106 268
use INVX1  _1709_
timestamp 0
transform 1 0 4250 0 1 5990
box -6 -8 66 268
use MUX2X1  _1710_
timestamp 0
transform -1 0 5830 0 -1 4430
box -6 -8 126 268
use INVX1  _1711_
timestamp 0
transform 1 0 5270 0 1 5470
box -6 -8 66 268
use INVX1  _1712_
timestamp 0
transform 1 0 7410 0 1 4430
box -6 -8 66 268
use INVX1  _1713_
timestamp 0
transform -1 0 9830 0 -1 270
box -6 -8 66 268
use NAND2X1  _1714_
timestamp 0
transform -1 0 10050 0 1 270
box -6 -8 86 268
use INVX1  _1715_
timestamp 0
transform -1 0 8710 0 1 270
box -6 -8 66 268
use NOR2X1  _1716_
timestamp 0
transform 1 0 11430 0 -1 1310
box -6 -8 86 268
use INVX1  _1717_
timestamp 0
transform 1 0 11230 0 1 270
box -6 -8 66 268
use NOR2X1  _1718_
timestamp 0
transform 1 0 12050 0 -1 790
box -6 -8 86 268
use NAND3X1  _1719_
timestamp 0
transform -1 0 9010 0 -1 790
box -6 -8 106 268
use INVX1  _1720_
timestamp 0
transform -1 0 10290 0 1 270
box -6 -8 66 268
use NAND2X1  _1721_
timestamp 0
transform -1 0 10330 0 -1 790
box -6 -8 86 268
use NAND2X1  _1722_
timestamp 0
transform -1 0 10110 0 -1 270
box -6 -8 86 268
use NOR2X1  _1723_
timestamp 0
transform 1 0 10130 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1724_
timestamp 0
transform 1 0 9350 0 1 2350
box -6 -8 86 268
use INVX1  _1725_
timestamp 0
transform 1 0 9190 0 -1 3390
box -6 -8 66 268
use NOR2X1  _1726_
timestamp 0
transform 1 0 10290 0 -1 270
box -6 -8 86 268
use NAND2X1  _1727_
timestamp 0
transform -1 0 8970 0 1 270
box -6 -8 86 268
use INVX2  _1728_
timestamp 0
transform 1 0 11690 0 -1 1310
box -6 -8 66 268
use NAND2X1  _1729_
timestamp 0
transform 1 0 10290 0 -1 3910
box -6 -8 86 268
use NOR2X1  _1730_
timestamp 0
transform 1 0 8470 0 1 4430
box -6 -8 86 268
use NOR2X1  _1731_
timestamp 0
transform 1 0 8710 0 -1 4430
box -6 -8 86 268
use AND2X2  _1732_
timestamp 0
transform -1 0 7990 0 -1 4430
box -6 -8 106 268
use NOR2X1  _1733_
timestamp 0
transform 1 0 9850 0 1 1310
box -6 -8 86 268
use INVX8  _1734_
timestamp 0
transform 1 0 7550 0 -1 3390
box -6 -8 126 268
use INVX1  _1735_
timestamp 0
transform 1 0 10990 0 1 270
box -6 -8 66 268
use NAND2X1  _1736_
timestamp 0
transform -1 0 10850 0 -1 790
box -6 -8 86 268
use NOR2X1  _1737_
timestamp 0
transform -1 0 11130 0 -1 790
box -6 -8 86 268
use INVX2  _1738_
timestamp 0
transform -1 0 10470 0 1 2870
box -6 -8 66 268
use NAND2X1  _1739_
timestamp 0
transform -1 0 10490 0 1 790
box -6 -8 86 268
use NOR2X1  _1740_
timestamp 0
transform 1 0 10650 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1741_
timestamp 0
transform -1 0 8610 0 1 2870
box -6 -8 86 268
use OAI21X1  _1742_
timestamp 0
transform -1 0 8530 0 -1 4430
box -6 -8 106 268
use NAND2X1  _1743_
timestamp 0
transform -1 0 10070 0 -1 790
box -6 -8 86 268
use NOR2X1  _1744_
timestamp 0
transform 1 0 9890 0 1 790
box -6 -8 86 268
use NAND2X1  _1745_
timestamp 0
transform -1 0 9650 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1746_
timestamp 0
transform 1 0 11450 0 1 790
box -6 -8 86 268
use NOR2X1  _1747_
timestamp 0
transform 1 0 10930 0 1 790
box -6 -8 86 268
use INVX1  _1748_
timestamp 0
transform 1 0 7650 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1749_
timestamp 0
transform 1 0 8070 0 1 3910
box -6 -8 106 268
use NOR2X1  _1750_
timestamp 0
transform -1 0 8250 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1751_
timestamp 0
transform 1 0 7610 0 -1 4430
box -6 -8 106 268
use NOR2X1  _1752_
timestamp 0
transform -1 0 9070 0 1 790
box -6 -8 86 268
use NOR2X1  _1753_
timestamp 0
transform 1 0 9870 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1754_
timestamp 0
transform -1 0 8490 0 -1 1830
box -6 -8 106 268
use INVX1  _1755_
timestamp 0
transform -1 0 9030 0 -1 8070
box -6 -8 66 268
use NAND2X1  _1756_
timestamp 0
transform -1 0 11390 0 -1 790
box -6 -8 86 268
use NOR2X1  _1757_
timestamp 0
transform 1 0 11190 0 1 790
box -6 -8 86 268
use OAI21X1  _1758_
timestamp 0
transform -1 0 9330 0 1 1830
box -6 -8 106 268
use INVX1  _1759_
timestamp 0
transform -1 0 7530 0 1 7550
box -6 -8 66 268
use AOI21X1  _1760_
timestamp 0
transform 1 0 8990 0 1 7550
box -6 -8 106 268
use AND2X2  _1761_
timestamp 0
transform -1 0 9790 0 1 270
box -6 -8 106 268
use NOR2X1  _1762_
timestamp 0
transform 1 0 10730 0 1 270
box -6 -8 86 268
use NAND2X1  _1763_
timestamp 0
transform -1 0 9230 0 1 270
box -6 -8 86 268
use INVX4  _1764_
timestamp 0
transform 1 0 11430 0 1 1310
box -6 -8 86 268
use NAND2X1  _1765_
timestamp 0
transform 1 0 8250 0 1 2350
box -6 -8 86 268
use NOR2X1  _1766_
timestamp 0
transform 1 0 8650 0 -1 5990
box -6 -8 86 268
use INVX1  _1767_
timestamp 0
transform 1 0 9330 0 -1 10150
box -6 -8 66 268
use NAND2X1  _1768_
timestamp 0
transform 1 0 8190 0 1 7550
box -6 -8 86 268
use OAI21X1  _1769_
timestamp 0
transform 1 0 8710 0 1 7550
box -6 -8 106 268
use OAI21X1  _1770_
timestamp 0
transform 1 0 9150 0 -1 7550
box -6 -8 106 268
use OAI21X1  _1771_
timestamp 0
transform 1 0 9110 0 1 7030
box -6 -8 106 268
use OAI21X1  _1772_
timestamp 0
transform 1 0 8830 0 1 7030
box -6 -8 106 268
use NOR2X1  _1773_
timestamp 0
transform 1 0 10910 0 1 1310
box -6 -8 86 268
use NOR2X1  _1774_
timestamp 0
transform 1 0 10910 0 -1 1310
box -6 -8 86 268
use NOR2X1  _1775_
timestamp 0
transform 1 0 10150 0 1 790
box -6 -8 86 268
use OAI21X1  _1776_
timestamp 0
transform -1 0 8230 0 1 1830
box -6 -8 106 268
use NAND3X1  _1777_
timestamp 0
transform 1 0 8190 0 1 4430
box -6 -8 106 268
use OR2X2  _1778_
timestamp 0
transform -1 0 7750 0 1 4430
box -6 -8 106 268
use INVX2  _1779_
timestamp 0
transform 1 0 5810 0 -1 2350
box -6 -8 66 268
use INVX1  _1780_
timestamp 0
transform -1 0 4250 0 1 5470
box -6 -8 66 268
use NAND2X1  _1781_
timestamp 0
transform -1 0 11010 0 1 2870
box -6 -8 86 268
use NAND2X1  _1782_
timestamp 0
transform 1 0 8410 0 1 1830
box -6 -8 86 268
use NOR2X1  _1783_
timestamp 0
transform 1 0 10650 0 1 1310
box -6 -8 86 268
use INVX2  _1784_
timestamp 0
transform -1 0 10170 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1785_
timestamp 0
transform -1 0 9970 0 1 2870
box -6 -8 106 268
use NAND2X1  _1786_
timestamp 0
transform 1 0 10310 0 1 3390
box -6 -8 86 268
use OAI21X1  _1787_
timestamp 0
transform -1 0 9330 0 1 3390
box -6 -8 106 268
use OR2X2  _1788_
timestamp 0
transform -1 0 8750 0 -1 3390
box -6 -8 106 268
use INVX1  _1789_
timestamp 0
transform 1 0 10110 0 1 2350
box -6 -8 66 268
use NOR2X1  _1790_
timestamp 0
transform -1 0 10230 0 1 2870
box -6 -8 86 268
use INVX1  _1791_
timestamp 0
transform -1 0 10290 0 1 5470
box -6 -8 66 268
use NOR2X1  _1792_
timestamp 0
transform -1 0 9850 0 -1 5990
box -6 -8 86 268
use NOR2X1  _1793_
timestamp 0
transform -1 0 9590 0 -1 270
box -6 -8 86 268
use NAND2X1  _1794_
timestamp 0
transform 1 0 9250 0 -1 270
box -6 -8 86 268
use OAI21X1  _1795_
timestamp 0
transform -1 0 8530 0 1 3390
box -6 -8 106 268
use NOR2X1  _1796_
timestamp 0
transform -1 0 8470 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1797_
timestamp 0
transform 1 0 7230 0 1 2870
box -6 -8 86 268
use INVX1  _1798_
timestamp 0
transform 1 0 7490 0 1 2870
box -6 -8 66 268
use NOR2X1  _1799_
timestamp 0
transform -1 0 9570 0 -1 4430
box -6 -8 86 268
use INVX1  _1800_
timestamp 0
transform 1 0 11390 0 1 1830
box -6 -8 66 268
use AND2X2  _1801_
timestamp 0
transform 1 0 9410 0 1 270
box -6 -8 106 268
use NAND2X1  _1802_
timestamp 0
transform -1 0 9130 0 -1 2350
box -6 -8 86 268
use NOR2X1  _1803_
timestamp 0
transform 1 0 10670 0 1 790
box -6 -8 86 268
use OAI21X1  _1804_
timestamp 0
transform -1 0 8770 0 -1 1830
box -6 -8 106 268
use NAND3X1  _1805_
timestamp 0
transform -1 0 8870 0 -1 2350
box -6 -8 106 268
use NOR2X1  _1806_
timestamp 0
transform 1 0 7730 0 1 2870
box -6 -8 86 268
use INVX1  _1807_
timestamp 0
transform -1 0 8230 0 -1 3910
box -6 -8 66 268
use INVX1  _1808_
timestamp 0
transform -1 0 8550 0 -1 270
box -6 -8 66 268
use NAND2X1  _1809_
timestamp 0
transform 1 0 8730 0 -1 270
box -6 -8 86 268
use OAI21X1  _1810_
timestamp 0
transform 1 0 8150 0 1 3390
box -6 -8 106 268
use OR2X2  _1811_
timestamp 0
transform -1 0 7950 0 1 3390
box -6 -8 106 268
use OAI21X1  _1812_
timestamp 0
transform -1 0 8590 0 -1 2870
box -6 -8 106 268
use OAI21X1  _1813_
timestamp 0
transform -1 0 8310 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1814_
timestamp 0
transform -1 0 8030 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1815_
timestamp 0
transform 1 0 7990 0 1 2870
box -6 -8 106 268
use OAI22X1  _1816_
timestamp 0
transform -1 0 4090 0 1 6510
box -6 -8 126 268
use INVX2  _1817_
timestamp 0
transform 1 0 1470 0 -1 1310
box -6 -8 66 268
use INVX2  _1818_
timestamp 0
transform -1 0 6330 0 -1 4430
box -6 -8 66 268
use OAI22X1  _1819_
timestamp 0
transform -1 0 1150 0 1 6510
box -6 -8 126 268
use INVX1  _1820_
timestamp 0
transform 1 0 490 0 -1 1830
box -6 -8 66 268
use OAI22X1  _1821_
timestamp 0
transform 1 0 1010 0 -1 7030
box -6 -8 126 268
use INVX2  _1822_
timestamp 0
transform -1 0 510 0 1 2350
box -6 -8 66 268
use OAI22X1  _1823_
timestamp 0
transform 1 0 1830 0 -1 7030
box -6 -8 126 268
use INVX1  _1824_
timestamp 0
transform 1 0 1410 0 -1 4430
box -6 -8 66 268
use OAI22X1  _1825_
timestamp 0
transform -1 0 1370 0 -1 5990
box -6 -8 126 268
use INVX2  _1826_
timestamp 0
transform -1 0 550 0 -1 3910
box -6 -8 66 268
use OAI22X1  _1827_
timestamp 0
transform 1 0 1010 0 -1 6510
box -6 -8 126 268
use INVX2  _1828_
timestamp 0
transform -1 0 1650 0 -1 3390
box -6 -8 66 268
use OAI22X1  _1829_
timestamp 0
transform -1 0 850 0 1 6510
box -6 -8 126 268
use INVX2  _1830_
timestamp 0
transform -1 0 1590 0 -1 2870
box -6 -8 66 268
use OAI22X1  _1831_
timestamp 0
transform 1 0 2130 0 -1 7030
box -6 -8 126 268
use OAI21X1  _1832_
timestamp 0
transform -1 0 8210 0 -1 1830
box -6 -8 106 268
use NAND2X1  _1833_
timestamp 0
transform 1 0 9770 0 1 1830
box -6 -8 86 268
use NAND2X1  _1834_
timestamp 0
transform 1 0 9350 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1835_
timestamp 0
transform -1 0 7950 0 1 1830
box -6 -8 106 268
use INVX1  _1836_
timestamp 0
transform -1 0 6570 0 1 5470
box -6 -8 66 268
use NAND2X1  _1837_
timestamp 0
transform -1 0 7930 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1838_
timestamp 0
transform -1 0 7390 0 -1 5470
box -6 -8 106 268
use INVX1  _1839_
timestamp 0
transform -1 0 6330 0 1 5470
box -6 -8 66 268
use NAND2X1  _1840_
timestamp 0
transform 1 0 8690 0 1 1830
box -6 -8 86 268
use NAND2X1  _1841_
timestamp 0
transform -1 0 8350 0 1 2870
box -6 -8 86 268
use INVX1  _1842_
timestamp 0
transform -1 0 7090 0 1 5470
box -6 -8 66 268
use NAND3X1  _1843_
timestamp 0
transform -1 0 6850 0 1 5470
box -6 -8 106 268
use NAND2X1  _1844_
timestamp 0
transform 1 0 9190 0 -1 790
box -6 -8 86 268
use NAND2X1  _1845_
timestamp 0
transform 1 0 9730 0 -1 790
box -6 -8 86 268
use NAND2X1  _1846_
timestamp 0
transform -1 0 9390 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1847_
timestamp 0
transform -1 0 8570 0 -1 4950
box -6 -8 106 268
use NAND2X1  _1848_
timestamp 0
transform 1 0 11330 0 -1 1830
box -6 -8 86 268
use NOR2X1  _1849_
timestamp 0
transform -1 0 11710 0 1 1830
box -6 -8 86 268
use INVX1  _1850_
timestamp 0
transform -1 0 11150 0 -1 1830
box -6 -8 66 268
use NOR2X1  _1851_
timestamp 0
transform 1 0 10470 0 1 270
box -6 -8 86 268
use NAND2X1  _1852_
timestamp 0
transform -1 0 10590 0 -1 790
box -6 -8 86 268
use OAI21X1  _1853_
timestamp 0
transform -1 0 10630 0 -1 1830
box -6 -8 106 268
use NOR2X1  _1854_
timestamp 0
transform -1 0 7610 0 1 6510
box -6 -8 86 268
use OAI21X1  _1855_
timestamp 0
transform 1 0 7510 0 1 5990
box -6 -8 106 268
use NOR2X1  _1856_
timestamp 0
transform 1 0 7790 0 1 5990
box -6 -8 86 268
use INVX1  _1857_
timestamp 0
transform -1 0 8970 0 -1 12230
box -6 -8 66 268
use NAND3X1  _1858_
timestamp 0
transform -1 0 9550 0 -1 790
box -6 -8 106 268
use OAI21X1  _1859_
timestamp 0
transform -1 0 9010 0 -1 11710
box -6 -8 106 268
use AOI21X1  _1860_
timestamp 0
transform 1 0 9190 0 1 11710
box -6 -8 106 268
use NOR3X1  _1861_
timestamp 0
transform 1 0 6930 0 -1 5470
box -6 -8 186 268
use NAND3X1  _1862_
timestamp 0
transform -1 0 8510 0 1 11190
box -6 -8 106 268
use OAI21X1  _1863_
timestamp 0
transform 1 0 7790 0 1 6510
box -6 -8 106 268
use INVX2  _1864_
timestamp 0
transform -1 0 6470 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1865_
timestamp 0
transform -1 0 7930 0 1 11190
box -6 -8 86 268
use NAND3X1  _1866_
timestamp 0
transform -1 0 7410 0 -1 11710
box -6 -8 106 268
use MUX2X1  _1867_
timestamp 0
transform -1 0 8210 0 1 11710
box -6 -8 126 268
use NOR2X1  _1868_
timestamp 0
transform 1 0 7830 0 1 11710
box -6 -8 86 268
use NAND2X1  _1869_
timestamp 0
transform -1 0 6210 0 1 10150
box -6 -8 86 268
use INVX1  _1870_
timestamp 0
transform 1 0 9470 0 1 11710
box -6 -8 66 268
use INVX1  _1871_
timestamp 0
transform 1 0 8950 0 1 11710
box -6 -8 66 268
use OAI21X1  _1872_
timestamp 0
transform -1 0 8770 0 1 11710
box -6 -8 106 268
use AND2X2  _1873_
timestamp 0
transform -1 0 7970 0 -1 11710
box -6 -8 106 268
use NAND3X1  _1874_
timestamp 0
transform -1 0 7690 0 -1 11710
box -6 -8 106 268
use OR2X2  _1875_
timestamp 0
transform -1 0 8490 0 1 11710
box -6 -8 106 268
use AOI21X1  _1876_
timestamp 0
transform -1 0 7130 0 -1 11710
box -6 -8 106 268
use NAND2X1  _1877_
timestamp 0
transform -1 0 5950 0 -1 9630
box -6 -8 86 268
use NOR2X1  _1878_
timestamp 0
transform 1 0 6770 0 -1 11710
box -6 -8 86 268
use AOI21X1  _1879_
timestamp 0
transform -1 0 7650 0 1 11710
box -6 -8 106 268
use AOI22X1  _1880_
timestamp 0
transform 1 0 6090 0 -1 10150
box -6 -8 126 268
use NAND3X1  _1881_
timestamp 0
transform 1 0 6090 0 1 9630
box -6 -8 106 268
use INVX1  _1882_
timestamp 0
transform -1 0 5090 0 -1 7550
box -6 -8 66 268
use INVX1  _1883_
timestamp 0
transform -1 0 7990 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1884_
timestamp 0
transform -1 0 8290 0 -1 4950
box -6 -8 106 268
use INVX1  _1885_
timestamp 0
transform -1 0 8790 0 1 4430
box -6 -8 66 268
use NOR2X1  _1886_
timestamp 0
transform 1 0 8590 0 1 5990
box -6 -8 86 268
use INVX1  _1887_
timestamp 0
transform -1 0 8610 0 1 6510
box -6 -8 66 268
use NAND2X1  _1888_
timestamp 0
transform 1 0 11710 0 1 790
box -6 -8 86 268
use OAI22X1  _1889_
timestamp 0
transform -1 0 8670 0 -1 6510
box -6 -8 126 268
use OAI21X1  _1890_
timestamp 0
transform 1 0 9830 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1891_
timestamp 0
transform 1 0 8990 0 -1 270
box -6 -8 86 268
use NOR2X1  _1892_
timestamp 0
transform -1 0 8770 0 -1 3910
box -6 -8 86 268
use INVX2  _1893_
timestamp 0
transform 1 0 12230 0 1 1310
box -6 -8 66 268
use NAND2X1  _1894_
timestamp 0
transform 1 0 12210 0 -1 2870
box -6 -8 86 268
use INVX1  _1895_
timestamp 0
transform 1 0 12230 0 1 2870
box -6 -8 66 268
use NOR2X1  _1896_
timestamp 0
transform -1 0 10910 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1897_
timestamp 0
transform -1 0 9310 0 -1 3910
box -6 -8 86 268
use NOR2X1  _1898_
timestamp 0
transform 1 0 9130 0 1 5990
box -6 -8 86 268
use INVX1  _1899_
timestamp 0
transform 1 0 7590 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1900_
timestamp 0
transform 1 0 9770 0 1 3390
box -6 -8 86 268
use NOR2X1  _1901_
timestamp 0
transform 1 0 8110 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1902_
timestamp 0
transform -1 0 8410 0 1 5990
box -6 -8 106 268
use NOR2X1  _1903_
timestamp 0
transform 1 0 8050 0 1 5990
box -6 -8 86 268
use NOR2X1  _1904_
timestamp 0
transform 1 0 11970 0 1 2870
box -6 -8 86 268
use INVX1  _1905_
timestamp 0
transform 1 0 11730 0 1 2870
box -6 -8 66 268
use INVX1  _1906_
timestamp 0
transform -1 0 6650 0 -1 3910
box -6 -8 66 268
use NAND2X1  _1907_
timestamp 0
transform -1 0 7210 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1908_
timestamp 0
transform -1 0 7150 0 1 3390
box -6 -8 106 268
use INVX1  _1909_
timestamp 0
transform -1 0 6870 0 1 3390
box -6 -8 66 268
use NAND3X1  _1910_
timestamp 0
transform -1 0 6410 0 -1 3910
box -6 -8 106 268
use INVX1  _1911_
timestamp 0
transform 1 0 6910 0 1 270
box -6 -8 66 268
use NOR2X1  _1912_
timestamp 0
transform 1 0 6370 0 -1 1310
box -6 -8 86 268
use INVX1  _1913_
timestamp 0
transform 1 0 6330 0 1 1310
box -6 -8 66 268
use OAI21X1  _1914_
timestamp 0
transform 1 0 5810 0 -1 4950
box -6 -8 106 268
use AOI21X1  _1915_
timestamp 0
transform 1 0 5330 0 -1 5470
box -6 -8 106 268
use OAI21X1  _1916_
timestamp 0
transform 1 0 5330 0 1 7030
box -6 -8 106 268
use NAND2X1  _1917_
timestamp 0
transform -1 0 3890 0 -1 9110
box -6 -8 86 268
use AOI22X1  _1918_
timestamp 0
transform 1 0 3710 0 1 10670
box -6 -8 126 268
use NAND2X1  _1919_
timestamp 0
transform -1 0 4050 0 1 8590
box -6 -8 86 268
use NAND3X1  _1920_
timestamp 0
transform -1 0 3790 0 1 8590
box -6 -8 106 268
use INVX1  _1921_
timestamp 0
transform -1 0 1870 0 1 7550
box -6 -8 66 268
use INVX1  _1922_
timestamp 0
transform 1 0 7630 0 1 270
box -6 -8 66 268
use NOR2X1  _1923_
timestamp 0
transform 1 0 7890 0 1 790
box -6 -8 86 268
use INVX1  _1924_
timestamp 0
transform -1 0 6530 0 1 2870
box -6 -8 66 268
use OAI21X1  _1925_
timestamp 0
transform -1 0 4810 0 1 5470
box -6 -8 106 268
use AOI21X1  _1926_
timestamp 0
transform -1 0 4170 0 -1 6510
box -6 -8 106 268
use OAI21X1  _1927_
timestamp 0
transform 1 0 2130 0 -1 7550
box -6 -8 106 268
use NAND2X1  _1928_
timestamp 0
transform -1 0 3370 0 -1 9110
box -6 -8 86 268
use AOI22X1  _1929_
timestamp 0
transform 1 0 4670 0 1 9630
box -6 -8 126 268
use NAND2X1  _1930_
timestamp 0
transform 1 0 3230 0 1 9110
box -6 -8 86 268
use NAND3X1  _1931_
timestamp 0
transform -1 0 3090 0 -1 9110
box -6 -8 106 268
use INVX1  _1932_
timestamp 0
transform -1 0 1650 0 -1 7030
box -6 -8 66 268
use NOR3X1  _1933_
timestamp 0
transform -1 0 8730 0 -1 790
box -6 -8 186 268
use NAND2X1  _1934_
timestamp 0
transform 1 0 3970 0 -1 790
box -6 -8 86 268
use OAI21X1  _1935_
timestamp 0
transform -1 0 4070 0 1 5990
box -6 -8 106 268
use AOI21X1  _1936_
timestamp 0
transform -1 0 2750 0 1 6510
box -6 -8 106 268
use OAI21X1  _1937_
timestamp 0
transform -1 0 1410 0 -1 7030
box -6 -8 106 268
use NAND2X1  _1938_
timestamp 0
transform -1 0 3750 0 -1 11710
box -6 -8 86 268
use AOI22X1  _1939_
timestamp 0
transform -1 0 4350 0 -1 11710
box -6 -8 126 268
use NAND2X1  _1940_
timestamp 0
transform -1 0 3530 0 1 11710
box -6 -8 86 268
use NAND3X1  _1941_
timestamp 0
transform -1 0 3490 0 -1 11710
box -6 -8 106 268
use INVX1  _1942_
timestamp 0
transform -1 0 1950 0 -1 7550
box -6 -8 66 268
use NAND2X1  _1943_
timestamp 0
transform -1 0 3790 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1944_
timestamp 0
transform -1 0 3890 0 -1 3910
box -6 -8 106 268
use AOI21X1  _1945_
timestamp 0
transform -1 0 3150 0 1 4950
box -6 -8 106 268
use OAI21X1  _1946_
timestamp 0
transform -1 0 1710 0 -1 7550
box -6 -8 106 268
use NAND2X1  _1947_
timestamp 0
transform -1 0 5110 0 -1 9110
box -6 -8 86 268
use AOI22X1  _1948_
timestamp 0
transform 1 0 5250 0 1 9630
box -6 -8 126 268
use NAND2X1  _1949_
timestamp 0
transform 1 0 5310 0 1 8590
box -6 -8 86 268
use NAND3X1  _1950_
timestamp 0
transform -1 0 5130 0 1 8590
box -6 -8 106 268
use INVX1  _1951_
timestamp 0
transform -1 0 2130 0 -1 6510
box -6 -8 66 268
use NAND2X1  _1952_
timestamp 0
transform 1 0 4210 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1953_
timestamp 0
transform 1 0 4150 0 -1 5470
box -6 -8 106 268
use AOI21X1  _1954_
timestamp 0
transform 1 0 4290 0 -1 5990
box -6 -8 106 268
use OAI21X1  _1955_
timestamp 0
transform -1 0 1890 0 -1 6510
box -6 -8 106 268
use NAND2X1  _1956_
timestamp 0
transform -1 0 4490 0 -1 11190
box -6 -8 86 268
use AOI22X1  _1957_
timestamp 0
transform 1 0 5010 0 -1 10670
box -6 -8 126 268
use NAND2X1  _1958_
timestamp 0
transform -1 0 5370 0 1 11190
box -6 -8 86 268
use NAND3X1  _1959_
timestamp 0
transform -1 0 4350 0 1 10670
box -6 -8 106 268
use INVX1  _1960_
timestamp 0
transform -1 0 2470 0 1 6510
box -6 -8 66 268
use NAND2X1  _1961_
timestamp 0
transform 1 0 4250 0 1 1310
box -6 -8 86 268
use OAI21X1  _1962_
timestamp 0
transform 1 0 4010 0 -1 5990
box -6 -8 106 268
use AOI21X1  _1963_
timestamp 0
transform 1 0 3790 0 -1 6510
box -6 -8 106 268
use OAI21X1  _1964_
timestamp 0
transform 1 0 2130 0 1 6510
box -6 -8 106 268
use NAND2X1  _1965_
timestamp 0
transform 1 0 6510 0 -1 11710
box -6 -8 86 268
use AOI22X1  _1966_
timestamp 0
transform 1 0 6450 0 1 11710
box -6 -8 126 268
use NAND2X1  _1967_
timestamp 0
transform 1 0 7290 0 1 11710
box -6 -8 86 268
use NAND3X1  _1968_
timestamp 0
transform 1 0 6750 0 1 11710
box -6 -8 106 268
use INVX1  _1969_
timestamp 0
transform -1 0 3450 0 1 7030
box -6 -8 66 268
use INVX1  _1970_
timestamp 0
transform 1 0 2950 0 1 2350
box -6 -8 66 268
use NOR2X1  _1971_
timestamp 0
transform -1 0 4890 0 1 2350
box -6 -8 86 268
use INVX1  _1972_
timestamp 0
transform 1 0 3710 0 1 5470
box -6 -8 66 268
use OAI21X1  _1973_
timestamp 0
transform -1 0 3790 0 1 5990
box -6 -8 106 268
use AOI21X1  _1974_
timestamp 0
transform -1 0 3290 0 1 6510
box -6 -8 106 268
use OAI21X1  _1975_
timestamp 0
transform 1 0 3110 0 1 7030
box -6 -8 106 268
use NAND2X1  _1976_
timestamp 0
transform -1 0 3270 0 1 11190
box -6 -8 86 268
use AOI22X1  _1977_
timestamp 0
transform 1 0 4490 0 1 11190
box -6 -8 126 268
use NAND2X1  _1978_
timestamp 0
transform 1 0 3190 0 1 11710
box -6 -8 86 268
use NAND3X1  _1979_
timestamp 0
transform -1 0 3010 0 1 11190
box -6 -8 106 268
use INVX1  _1980_
timestamp 0
transform -1 0 2490 0 -1 7030
box -6 -8 66 268
use INVX1  _1981_
timestamp 0
transform 1 0 6070 0 1 1310
box -6 -8 66 268
use NOR2X1  _1982_
timestamp 0
transform 1 0 6190 0 1 1830
box -6 -8 86 268
use INVX1  _1983_
timestamp 0
transform 1 0 6390 0 1 2350
box -6 -8 66 268
use OAI21X1  _1984_
timestamp 0
transform 1 0 5390 0 1 4950
box -6 -8 106 268
use AOI21X1  _1985_
timestamp 0
transform -1 0 4970 0 -1 6510
box -6 -8 106 268
use OAI21X1  _1986_
timestamp 0
transform 1 0 2670 0 -1 7030
box -6 -8 106 268
use NAND2X1  _1987_
timestamp 0
transform -1 0 7470 0 -1 3910
box -6 -8 86 268
use INVX1  _1988_
timestamp 0
transform 1 0 7690 0 -1 4950
box -6 -8 66 268
use OR2X2  _1989_
timestamp 0
transform 1 0 7750 0 -1 6510
box -6 -8 106 268
use AND2X2  _1990_
timestamp 0
transform -1 0 7630 0 1 5470
box -6 -8 106 268
use AOI22X1  _1991_
timestamp 0
transform -1 0 7930 0 1 5470
box -6 -8 126 268
use OR2X2  _1992_
timestamp 0
transform 1 0 10570 0 -1 5990
box -6 -8 106 268
use NOR2X1  _1993_
timestamp 0
transform 1 0 9690 0 -1 8070
box -6 -8 86 268
use INVX1  _1994_
timestamp 0
transform -1 0 6410 0 -1 8590
box -6 -8 66 268
use INVX1  _1995_
timestamp 0
transform 1 0 6750 0 -1 270
box -6 -8 66 268
use INVX1  _1996_
timestamp 0
transform -1 0 6930 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1997_
timestamp 0
transform 1 0 6590 0 -1 2870
box -6 -8 106 268
use AOI21X1  _1998_
timestamp 0
transform 1 0 6590 0 -1 8590
box -6 -8 106 268
use OAI21X1  _1999_
timestamp 0
transform 1 0 7650 0 1 8590
box -6 -8 106 268
use INVX1  _2000_
timestamp 0
transform 1 0 6570 0 1 8590
box -6 -8 66 268
use AOI21X1  _2001_
timestamp 0
transform 1 0 6810 0 1 8590
box -6 -8 106 268
use OAI21X1  _2002_
timestamp 0
transform 1 0 6790 0 -1 9110
box -6 -8 106 268
use NAND2X1  _2003_
timestamp 0
transform 1 0 9650 0 1 10150
box -6 -8 86 268
use INVX1  _2004_
timestamp 0
transform 1 0 7590 0 -1 9110
box -6 -8 66 268
use AOI21X1  _2005_
timestamp 0
transform -1 0 7470 0 1 8590
box -6 -8 106 268
use OAI21X1  _2006_
timestamp 0
transform 1 0 6870 0 -1 8590
box -6 -8 106 268
use INVX1  _2007_
timestamp 0
transform 1 0 6710 0 1 2870
box -6 -8 66 268
use NAND2X1  _2008_
timestamp 0
transform -1 0 6410 0 -1 2870
box -6 -8 86 268
use OAI21X1  _2009_
timestamp 0
transform 1 0 6950 0 1 2870
box -6 -8 106 268
use NAND2X1  _2010_
timestamp 0
transform -1 0 7230 0 1 9110
box -6 -8 86 268
use OAI21X1  _2011_
timestamp 0
transform 1 0 7410 0 1 9110
box -6 -8 106 268
use NAND2X1  _2012_
timestamp 0
transform -1 0 9610 0 1 9110
box -6 -8 86 268
use NAND2X1  _2013_
timestamp 0
transform 1 0 10690 0 1 10150
box -6 -8 86 268
use NOR2X1  _2014_
timestamp 0
transform -1 0 11010 0 -1 9630
box -6 -8 86 268
use NAND2X1  _2015_
timestamp 0
transform -1 0 6450 0 1 9110
box -6 -8 86 268
use OAI21X1  _2016_
timestamp 0
transform -1 0 7530 0 1 9630
box -6 -8 106 268
use NAND2X1  _2017_
timestamp 0
transform -1 0 7270 0 -1 10150
box -6 -8 86 268
use OAI21X1  _2018_
timestamp 0
transform 1 0 7450 0 -1 10150
box -6 -8 106 268
use OAI21X1  _2019_
timestamp 0
transform 1 0 9530 0 1 9630
box -6 -8 106 268
use INVX1  _2020_
timestamp 0
transform -1 0 10470 0 -1 9630
box -6 -8 66 268
use NAND2X1  _2021_
timestamp 0
transform -1 0 7530 0 -1 9630
box -6 -8 86 268
use OAI21X1  _2022_
timestamp 0
transform 1 0 7710 0 -1 9630
box -6 -8 106 268
use NAND2X1  _2023_
timestamp 0
transform -1 0 8070 0 -1 9630
box -6 -8 86 268
use NAND2X1  _2024_
timestamp 0
transform 1 0 6230 0 -1 9110
box -6 -8 86 268
use OAI21X1  _2025_
timestamp 0
transform -1 0 6190 0 1 9110
box -6 -8 106 268
use AND2X2  _2026_
timestamp 0
transform 1 0 9810 0 1 9630
box -6 -8 106 268
use NAND2X1  _2027_
timestamp 0
transform 1 0 10350 0 1 9630
box -6 -8 86 268
use NOR2X1  _2028_
timestamp 0
transform -1 0 10410 0 1 9110
box -6 -8 86 268
use NAND3X1  _2029_
timestamp 0
transform -1 0 11310 0 -1 8070
box -6 -8 106 268
use NAND3X1  _2030_
timestamp 0
transform 1 0 10850 0 -1 5990
box -6 -8 106 268
use INVX1  _2031_
timestamp 0
transform -1 0 11210 0 -1 5990
box -6 -8 66 268
use NAND2X1  _2032_
timestamp 0
transform 1 0 9070 0 -1 9630
box -6 -8 86 268
use INVX1  _2033_
timestamp 0
transform 1 0 8530 0 -1 10150
box -6 -8 66 268
use OAI21X1  _2034_
timestamp 0
transform 1 0 8770 0 -1 10150
box -6 -8 106 268
use AOI21X1  _2035_
timestamp 0
transform 1 0 8730 0 1 9630
box -6 -8 106 268
use NAND2X1  _2036_
timestamp 0
transform 1 0 11690 0 1 9630
box -6 -8 86 268
use INVX1  _2037_
timestamp 0
transform 1 0 11890 0 1 11190
box -6 -8 66 268
use INVX1  _2038_
timestamp 0
transform -1 0 7770 0 -1 10670
box -6 -8 66 268
use NOR2X1  _2039_
timestamp 0
transform -1 0 6870 0 1 10670
box -6 -8 86 268
use NAND2X1  _2040_
timestamp 0
transform 1 0 11070 0 1 10670
box -6 -8 86 268
use NAND2X1  _2041_
timestamp 0
transform 1 0 11150 0 -1 9110
box -6 -8 86 268
use INVX1  _2042_
timestamp 0
transform -1 0 10270 0 -1 11190
box -6 -8 66 268
use NAND2X1  _2043_
timestamp 0
transform -1 0 10670 0 1 9110
box -6 -8 86 268
use OAI21X1  _2044_
timestamp 0
transform -1 0 11210 0 1 9110
box -6 -8 106 268
use NAND3X1  _2045_
timestamp 0
transform -1 0 11550 0 1 8590
box -6 -8 106 268
use NOR2X1  _2046_
timestamp 0
transform 1 0 8970 0 -1 3910
box -6 -8 86 268
use INVX1  _2047_
timestamp 0
transform -1 0 9550 0 -1 3910
box -6 -8 66 268
use NAND2X1  _2048_
timestamp 0
transform 1 0 9310 0 -1 2870
box -6 -8 86 268
use INVX1  _2049_
timestamp 0
transform 1 0 9450 0 1 3910
box -6 -8 66 268
use NAND2X1  _2050_
timestamp 0
transform 1 0 9210 0 -1 1830
box -6 -8 86 268
use OAI21X1  _2051_
timestamp 0
transform 1 0 8910 0 1 3910
box -6 -8 106 268
use NOR2X1  _2052_
timestamp 0
transform 1 0 9190 0 1 3910
box -6 -8 86 268
use OAI21X1  _2053_
timestamp 0
transform -1 0 9830 0 -1 3910
box -6 -8 106 268
use INVX1  _2054_
timestamp 0
transform 1 0 9970 0 1 5990
box -6 -8 66 268
use NOR2X1  _2055_
timestamp 0
transform -1 0 6670 0 -1 4950
box -6 -8 86 268
use INVX1  _2056_
timestamp 0
transform -1 0 6230 0 -1 5470
box -6 -8 66 268
use NOR2X1  _2057_
timestamp 0
transform 1 0 10390 0 -1 1310
box -6 -8 86 268
use OAI21X1  _2058_
timestamp 0
transform -1 0 10210 0 -1 2350
box -6 -8 106 268
use OAI21X1  _2059_
timestamp 0
transform -1 0 10350 0 -1 3390
box -6 -8 106 268
use NAND3X1  _2060_
timestamp 0
transform -1 0 10110 0 -1 3910
box -6 -8 106 268
use NAND3X1  _2061_
timestamp 0
transform 1 0 10230 0 1 5990
box -6 -8 106 268
use NOR2X1  _2062_
timestamp 0
transform -1 0 9350 0 1 6510
box -6 -8 86 268
use NAND2X1  _2063_
timestamp 0
transform 1 0 8370 0 -1 5990
box -6 -8 86 268
use NOR2X1  _2064_
timestamp 0
transform -1 0 8110 0 -1 6510
box -6 -8 86 268
use NAND3X1  _2065_
timestamp 0
transform -1 0 8950 0 -1 6510
box -6 -8 106 268
use OAI21X1  _2066_
timestamp 0
transform 1 0 8850 0 1 5990
box -6 -8 106 268
use OAI21X1  _2067_
timestamp 0
transform -1 0 8190 0 1 4950
box -6 -8 106 268
use OAI21X1  _2068_
timestamp 0
transform -1 0 8470 0 1 4950
box -6 -8 106 268
use OAI21X1  _2069_
timestamp 0
transform 1 0 8110 0 1 5470
box -6 -8 106 268
use OAI21X1  _2070_
timestamp 0
transform -1 0 8490 0 1 5470
box -6 -8 106 268
use NAND2X1  _2071_
timestamp 0
transform -1 0 8750 0 1 5470
box -6 -8 86 268
use NAND2X1  _2072_
timestamp 0
transform 1 0 8910 0 -1 5990
box -6 -8 86 268
use NAND3X1  _2073_
timestamp 0
transform 1 0 9170 0 -1 5990
box -6 -8 106 268
use OR2X2  _2074_
timestamp 0
transform 1 0 9390 0 1 5990
box -6 -8 106 268
use AOI21X1  _2075_
timestamp 0
transform -1 0 9790 0 1 5990
box -6 -8 106 268
use AND2X2  _2076_
timestamp 0
transform 1 0 11350 0 1 5990
box -6 -8 106 268
use NAND3X1  _2077_
timestamp 0
transform -1 0 11490 0 -1 5990
box -6 -8 106 268
use INVX1  _2078_
timestamp 0
transform -1 0 11250 0 1 10150
box -6 -8 66 268
use NAND2X1  _2079_
timestamp 0
transform 1 0 11350 0 1 11190
box -6 -8 86 268
use NAND2X1  _2080_
timestamp 0
transform -1 0 11250 0 1 9630
box -6 -8 86 268
use NOR2X1  _2081_
timestamp 0
transform 1 0 11190 0 -1 9630
box -6 -8 86 268
use AOI22X1  _2082_
timestamp 0
transform 1 0 10450 0 -1 7030
box -6 -8 126 268
use INVX8  _2083_
timestamp 0
transform 1 0 9710 0 1 11190
box -6 -8 126 268
use INVX2  _2084_
timestamp 0
transform 1 0 11730 0 -1 9630
box -6 -8 66 268
use NAND2X1  _2085_
timestamp 0
transform 1 0 11150 0 1 8070
box -6 -8 86 268
use NOR2X1  _2086_
timestamp 0
transform 1 0 11650 0 1 7550
box -6 -8 86 268
use AOI21X1  _2087_
timestamp 0
transform 1 0 11670 0 -1 5990
box -6 -8 106 268
use NOR2X1  _2088_
timestamp 0
transform -1 0 12290 0 -1 4430
box -6 -8 86 268
use OAI21X1  _2089_
timestamp 0
transform 1 0 11950 0 1 4430
box -6 -8 106 268
use OAI21X1  _2090_
timestamp 0
transform 1 0 12150 0 -1 4950
box -6 -8 106 268
use NAND2X1  _2091_
timestamp 0
transform 1 0 10030 0 1 1830
box -6 -8 86 268
use NOR2X1  _2092_
timestamp 0
transform 1 0 10650 0 1 2870
box -6 -8 86 268
use NAND2X1  _2093_
timestamp 0
transform -1 0 11270 0 1 2870
box -6 -8 86 268
use OAI21X1  _2094_
timestamp 0
transform 1 0 11450 0 1 2870
box -6 -8 106 268
use NAND2X1  _2095_
timestamp 0
transform -1 0 11170 0 -1 3910
box -6 -8 86 268
use OAI21X1  _2096_
timestamp 0
transform 1 0 11630 0 -1 3910
box -6 -8 106 268
use NOR2X1  _2097_
timestamp 0
transform -1 0 12030 0 1 3910
box -6 -8 86 268
use AND2X2  _2098_
timestamp 0
transform -1 0 12230 0 -1 270
box -6 -8 106 268
use NAND2X1  _2099_
timestamp 0
transform -1 0 11510 0 -1 2870
box -6 -8 86 268
use NAND2X1  _2100_
timestamp 0
transform 1 0 11410 0 1 3390
box -6 -8 86 268
use OAI21X1  _2101_
timestamp 0
transform -1 0 11450 0 -1 3910
box -6 -8 106 268
use NAND2X1  _2102_
timestamp 0
transform -1 0 11810 0 1 2350
box -6 -8 86 268
use NAND2X1  _2103_
timestamp 0
transform 1 0 12230 0 -1 2350
box -6 -8 86 268
use INVX1  _2104_
timestamp 0
transform 1 0 12230 0 -1 12230
box -6 -8 66 268
use NAND2X1  _2105_
timestamp 0
transform -1 0 11770 0 1 3390
box -6 -8 86 268
use OAI21X1  _2106_
timestamp 0
transform -1 0 11750 0 -1 3390
box -6 -8 106 268
use NOR2X1  _2107_
timestamp 0
transform -1 0 12290 0 1 3910
box -6 -8 86 268
use NOR2X1  _2108_
timestamp 0
transform 1 0 8970 0 1 3390
box -6 -8 86 268
use OAI21X1  _2109_
timestamp 0
transform 1 0 12230 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2110_
timestamp 0
transform -1 0 12330 0 1 3390
box -6 -8 106 268
use AND2X2  _2111_
timestamp 0
transform -1 0 12330 0 1 4430
box -6 -8 106 268
use AND2X2  _2112_
timestamp 0
transform -1 0 12230 0 -1 11710
box -6 -8 106 268
use NAND3X1  _2113_
timestamp 0
transform 1 0 11910 0 -1 5470
box -6 -8 106 268
use INVX1  _2114_
timestamp 0
transform 1 0 10690 0 -1 7550
box -6 -8 66 268
use OAI21X1  _2115_
timestamp 0
transform -1 0 9510 0 -1 6510
box -6 -8 106 268
use OAI21X1  _2116_
timestamp 0
transform -1 0 10390 0 -1 5990
box -6 -8 106 268
use NOR2X1  _2117_
timestamp 0
transform -1 0 10970 0 -1 9110
box -6 -8 86 268
use NOR2X1  _2118_
timestamp 0
transform -1 0 10930 0 1 7550
box -6 -8 86 268
use AOI22X1  _2119_
timestamp 0
transform 1 0 10790 0 -1 6510
box -6 -8 126 268
use OAI21X1  _2120_
timestamp 0
transform 1 0 10810 0 1 3910
box -6 -8 106 268
use OAI21X1  _2121_
timestamp 0
transform -1 0 10630 0 1 3910
box -6 -8 106 268
use NAND2X1  _2122_
timestamp 0
transform 1 0 10750 0 -1 5470
box -6 -8 86 268
use NAND2X1  _2123_
timestamp 0
transform -1 0 8310 0 -1 270
box -6 -8 86 268
use NOR2X1  _2124_
timestamp 0
transform -1 0 8010 0 1 4430
box -6 -8 86 268
use OAI21X1  _2125_
timestamp 0
transform -1 0 10390 0 -1 4430
box -6 -8 106 268
use OAI21X1  _2126_
timestamp 0
transform 1 0 10710 0 -1 4950
box -6 -8 106 268
use OAI21X1  _2127_
timestamp 0
transform -1 0 7210 0 -1 2870
box -6 -8 106 268
use NOR3X1  _2128_
timestamp 0
transform -1 0 9430 0 1 790
box -6 -8 186 268
use OAI21X1  _2129_
timestamp 0
transform 1 0 7390 0 -1 2870
box -6 -8 106 268
use NAND2X1  _2130_
timestamp 0
transform -1 0 11070 0 -1 4950
box -6 -8 86 268
use NAND2X1  _2131_
timestamp 0
transform -1 0 8110 0 -1 1310
box -6 -8 86 268
use XOR2X1  _2132_
timestamp 0
transform 1 0 6830 0 1 4430
box -6 -8 126 268
use NAND2X1  _2133_
timestamp 0
transform -1 0 7190 0 -1 4950
box -6 -8 86 268
use OAI22X1  _2134_
timestamp 0
transform -1 0 7510 0 -1 4950
box -6 -8 126 268
use NOR3X1  _2135_
timestamp 0
transform -1 0 11430 0 -1 4950
box -6 -8 186 268
use OAI21X1  _2136_
timestamp 0
transform -1 0 11510 0 1 3910
box -6 -8 106 268
use OAI21X1  _2137_
timestamp 0
transform 1 0 11410 0 1 4430
box -6 -8 106 268
use INVX1  _2138_
timestamp 0
transform 1 0 11490 0 1 2350
box -6 -8 66 268
use OAI21X1  _2139_
timestamp 0
transform -1 0 11490 0 -1 4430
box -6 -8 106 268
use OAI21X1  _2140_
timestamp 0
transform -1 0 11210 0 -1 4430
box -6 -8 106 268
use INVX1  _2141_
timestamp 0
transform 1 0 10050 0 1 4430
box -6 -8 66 268
use OAI21X1  _2142_
timestamp 0
transform 1 0 10850 0 1 4430
box -6 -8 106 268
use OAI21X1  _2143_
timestamp 0
transform -1 0 10670 0 1 4430
box -6 -8 106 268
use NAND3X1  _2144_
timestamp 0
transform -1 0 11230 0 1 4430
box -6 -8 106 268
use INVX4  _2145_
timestamp 0
transform -1 0 5210 0 1 4950
box -6 -8 86 268
use OAI21X1  _2146_
timestamp 0
transform 1 0 9870 0 -1 4950
box -6 -8 106 268
use OAI21X1  _2147_
timestamp 0
transform 1 0 10430 0 -1 4950
box -6 -8 106 268
use INVX2  _2148_
timestamp 0
transform -1 0 6410 0 -1 4950
box -6 -8 66 268
use NAND2X1  _2149_
timestamp 0
transform 1 0 10170 0 -1 4950
box -6 -8 86 268
use OAI21X1  _2150_
timestamp 0
transform 1 0 8930 0 1 4950
box -6 -8 106 268
use NOR2X1  _2151_
timestamp 0
transform 1 0 7550 0 1 4950
box -6 -8 86 268
use NAND2X1  _2152_
timestamp 0
transform 1 0 8630 0 -1 5470
box -6 -8 86 268
use OAI21X1  _2153_
timestamp 0
transform 1 0 8890 0 -1 5470
box -6 -8 106 268
use NOR2X1  _2154_
timestamp 0
transform 1 0 9170 0 -1 5470
box -6 -8 86 268
use NAND2X1  _2155_
timestamp 0
transform -1 0 10310 0 -1 5470
box -6 -8 86 268
use NOR2X1  _2156_
timestamp 0
transform -1 0 11090 0 -1 5470
box -6 -8 86 268
use NAND3X1  _2157_
timestamp 0
transform 1 0 11270 0 1 5470
box -6 -8 106 268
use NOR3X1  _2158_
timestamp 0
transform -1 0 12010 0 1 5470
box -6 -8 186 268
use INVX1  _2159_
timestamp 0
transform -1 0 12010 0 1 270
box -6 -8 66 268
use INVX1  _2160_
timestamp 0
transform -1 0 11550 0 -1 8070
box -6 -8 66 268
use OAI21X1  _2161_
timestamp 0
transform 1 0 8250 0 -1 9630
box -6 -8 106 268
use NAND2X1  _2162_
timestamp 0
transform 1 0 9010 0 1 9630
box -6 -8 86 268
use NOR2X1  _2163_
timestamp 0
transform -1 0 10170 0 1 9630
box -6 -8 86 268
use NAND2X1  _2164_
timestamp 0
transform 1 0 9890 0 -1 9630
box -6 -8 86 268
use NOR2X1  _2165_
timestamp 0
transform 1 0 11110 0 1 7550
box -6 -8 86 268
use AOI22X1  _2166_
timestamp 0
transform 1 0 10930 0 -1 7550
box -6 -8 126 268
use INVX1  _2167_
timestamp 0
transform 1 0 9310 0 -1 7030
box -6 -8 66 268
use NAND2X1  _2168_
timestamp 0
transform 1 0 10130 0 -1 10150
box -6 -8 86 268
use NOR2X1  _2169_
timestamp 0
transform -1 0 8930 0 -1 9110
box -6 -8 86 268
use NAND2X1  _2170_
timestamp 0
transform -1 0 9350 0 -1 8590
box -6 -8 86 268
use NOR2X1  _2171_
timestamp 0
transform 1 0 10430 0 -1 8070
box -6 -8 86 268
use AOI22X1  _2172_
timestamp 0
transform 1 0 9850 0 -1 7030
box -6 -8 126 268
use NAND2X1  _2173_
timestamp 0
transform 1 0 9970 0 -1 6510
box -6 -8 86 268
use OAI21X1  _2174_
timestamp 0
transform -1 0 9690 0 -1 4950
box -6 -8 106 268
use NAND3X1  _2175_
timestamp 0
transform 1 0 9690 0 1 3910
box -6 -8 106 268
use NOR2X1  _2176_
timestamp 0
transform -1 0 9870 0 1 4430
box -6 -8 86 268
use NAND2X1  _2177_
timestamp 0
transform -1 0 9570 0 1 4950
box -6 -8 86 268
use NAND3X1  _2178_
timestamp 0
transform -1 0 11210 0 -1 3390
box -6 -8 106 268
use AND2X2  _2179_
timestamp 0
transform 1 0 9590 0 -1 9110
box -6 -8 106 268
use NAND2X1  _2180_
timestamp 0
transform 1 0 11950 0 1 9630
box -6 -8 86 268
use NOR2X1  _2181_
timestamp 0
transform 1 0 11930 0 1 10150
box -6 -8 86 268
use NAND2X1  _2182_
timestamp 0
transform 1 0 12010 0 1 8590
box -6 -8 86 268
use OR2X2  _2183_
timestamp 0
transform -1 0 11470 0 1 7550
box -6 -8 106 268
use NAND3X1  _2184_
timestamp 0
transform 1 0 11130 0 1 4950
box -6 -8 106 268
use INVX1  _2185_
timestamp 0
transform -1 0 10410 0 1 8590
box -6 -8 66 268
use NOR2X1  _2186_
timestamp 0
transform 1 0 10310 0 -1 8590
box -6 -8 86 268
use INVX1  _2187_
timestamp 0
transform -1 0 10750 0 -1 8070
box -6 -8 66 268
use NOR2X1  _2188_
timestamp 0
transform 1 0 11670 0 1 10150
box -6 -8 86 268
use NAND2X1  _2189_
timestamp 0
transform 1 0 10050 0 -1 8590
box -6 -8 86 268
use OAI22X1  _2190_
timestamp 0
transform 1 0 10610 0 1 7030
box -6 -8 126 268
use INVX1  _2191_
timestamp 0
transform 1 0 11230 0 -1 7550
box -6 -8 66 268
use NOR2X1  _2192_
timestamp 0
transform 1 0 11170 0 -1 1310
box -6 -8 86 268
use MUX2X1  _2193_
timestamp 0
transform -1 0 11230 0 1 3910
box -6 -8 126 268
use INVX1  _2194_
timestamp 0
transform -1 0 10710 0 -1 9110
box -6 -8 66 268
use NAND2X1  _2195_
timestamp 0
transform -1 0 9610 0 -1 8590
box -6 -8 86 268
use OAI21X1  _2196_
timestamp 0
transform -1 0 11270 0 1 7030
box -6 -8 106 268
use NOR2X1  _2197_
timestamp 0
transform 1 0 11450 0 1 7030
box -6 -8 86 268
use NAND3X1  _2198_
timestamp 0
transform -1 0 10070 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2199_
timestamp 0
transform -1 0 10130 0 1 3390
box -6 -8 106 268
use AND2X2  _2200_
timestamp 0
transform -1 0 5990 0 1 6510
box -6 -8 106 268
use INVX1  _2201_
timestamp 0
transform 1 0 6430 0 -1 6510
box -6 -8 66 268
use NOR2X1  _2202_
timestamp 0
transform 1 0 6170 0 -1 6510
box -6 -8 86 268
use OAI21X1  _2203_
timestamp 0
transform 1 0 6170 0 1 6510
box -6 -8 106 268
use MUX2X1  _2204_
timestamp 0
transform 1 0 6910 0 -1 7030
box -6 -8 126 268
use OAI21X1  _2205_
timestamp 0
transform 1 0 7210 0 -1 7030
box -6 -8 106 268
use XOR2X1  _2206_
timestamp 0
transform 1 0 9550 0 -1 7030
box -6 -8 126 268
use NAND2X1  _2207_
timestamp 0
transform -1 0 10110 0 -1 5990
box -6 -8 86 268
use OAI22X1  _2208_
timestamp 0
transform -1 0 9590 0 -1 5990
box -6 -8 126 268
use NOR2X1  _2209_
timestamp 0
transform 1 0 10510 0 1 5990
box -6 -8 86 268
use NAND2X1  _2210_
timestamp 0
transform 1 0 10510 0 -1 6510
box -6 -8 86 268
use NOR3X1  _2211_
timestamp 0
transform 1 0 11350 0 -1 6510
box -6 -8 186 268
use NOR2X1  _2212_
timestamp 0
transform -1 0 11770 0 1 4430
box -6 -8 86 268
use NOR2X1  _2213_
timestamp 0
transform -1 0 11810 0 -1 7550
box -6 -8 86 268
use AOI22X1  _2214_
timestamp 0
transform 1 0 11710 0 1 7030
box -6 -8 126 268
use INVX1  _2215_
timestamp 0
transform 1 0 11810 0 -1 11190
box -6 -8 66 268
use OAI21X1  _2216_
timestamp 0
transform 1 0 12190 0 1 10150
box -6 -8 106 268
use NOR2X1  _2217_
timestamp 0
transform 1 0 11470 0 -1 7550
box -6 -8 86 268
use NOR2X1  _2218_
timestamp 0
transform 1 0 9750 0 -1 4430
box -6 -8 86 268
use OAI21X1  _2219_
timestamp 0
transform -1 0 10070 0 1 3910
box -6 -8 106 268
use OAI21X1  _2220_
timestamp 0
transform -1 0 10110 0 -1 4430
box -6 -8 106 268
use OAI21X1  _2221_
timestamp 0
transform -1 0 12050 0 1 3390
box -6 -8 106 268
use OAI21X1  _2222_
timestamp 0
transform 1 0 11910 0 -1 3910
box -6 -8 106 268
use NAND3X1  _2223_
timestamp 0
transform -1 0 12050 0 -1 3390
box -6 -8 106 268
use NAND3X1  _2224_
timestamp 0
transform 1 0 11930 0 -1 4430
box -6 -8 106 268
use AOI21X1  _2225_
timestamp 0
transform 1 0 11030 0 -1 270
box -6 -8 106 268
use AND2X2  _2226_
timestamp 0
transform 1 0 11990 0 -1 7550
box -6 -8 106 268
use NAND2X1  _2227_
timestamp 0
transform 1 0 11710 0 -1 6510
box -6 -8 86 268
use OR2X2  _2228_
timestamp 0
transform -1 0 11650 0 1 5470
box -6 -8 106 268
use INVX1  _2229_
timestamp 0
transform -1 0 10690 0 -1 2870
box -6 -8 66 268
use OAI21X1  _2230_
timestamp 0
transform -1 0 10450 0 -1 2870
box -6 -8 106 268
use NAND2X1  _2231_
timestamp 0
transform -1 0 8630 0 -1 1310
box -6 -8 86 268
use OAI21X1  _2232_
timestamp 0
transform 1 0 8810 0 -1 1310
box -6 -8 106 268
use NOR2X1  _2233_
timestamp 0
transform 1 0 9590 0 1 1310
box -6 -8 86 268
use NAND3X1  _2234_
timestamp 0
transform -1 0 9930 0 -1 2870
box -6 -8 106 268
use NAND3X1  _2235_
timestamp 0
transform -1 0 10050 0 1 5470
box -6 -8 106 268
use OAI21X1  _2236_
timestamp 0
transform 1 0 7270 0 1 4950
box -6 -8 106 268
use NOR2X1  _2237_
timestamp 0
transform -1 0 6830 0 1 4950
box -6 -8 86 268
use NAND2X1  _2238_
timestamp 0
transform -1 0 7090 0 1 4950
box -6 -8 86 268
use OAI21X1  _2239_
timestamp 0
transform -1 0 9130 0 -1 4950
box -6 -8 106 268
use OAI21X1  _2240_
timestamp 0
transform -1 0 8850 0 -1 4950
box -6 -8 106 268
use INVX1  _2241_
timestamp 0
transform -1 0 8450 0 -1 5470
box -6 -8 66 268
use OAI21X1  _2242_
timestamp 0
transform -1 0 7670 0 -1 5470
box -6 -8 106 268
use OAI21X1  _2243_
timestamp 0
transform 1 0 7850 0 -1 5470
box -6 -8 106 268
use NOR2X1  _2244_
timestamp 0
transform 1 0 8130 0 -1 5470
box -6 -8 86 268
use NAND3X1  _2245_
timestamp 0
transform -1 0 7910 0 1 4950
box -6 -8 106 268
use AOI21X1  _2246_
timestamp 0
transform 1 0 9210 0 1 4950
box -6 -8 106 268
use NAND2X1  _2247_
timestamp 0
transform -1 0 12270 0 1 270
box -6 -8 86 268
use INVX1  _2248_
timestamp 0
transform 1 0 11410 0 -1 10670
box -6 -8 66 268
use NOR2X1  _2249_
timestamp 0
transform -1 0 9630 0 -1 10670
box -6 -8 86 268
use NAND2X1  _2250_
timestamp 0
transform 1 0 11090 0 1 11190
box -6 -8 86 268
use OAI21X1  _2251_
timestamp 0
transform 1 0 10650 0 -1 9630
box -6 -8 106 268
use AOI21X1  _2252_
timestamp 0
transform 1 0 11410 0 1 9110
box -6 -8 106 268
use NAND2X1  _2253_
timestamp 0
transform -1 0 12050 0 1 9110
box -6 -8 86 268
use INVX1  _2254_
timestamp 0
transform 1 0 12230 0 1 9110
box -6 -8 66 268
use OAI21X1  _2255_
timestamp 0
transform -1 0 10670 0 -1 8590
box -6 -8 106 268
use NOR2X1  _2256_
timestamp 0
transform -1 0 10930 0 -1 8590
box -6 -8 86 268
use NAND3X1  _2257_
timestamp 0
transform 1 0 11110 0 -1 8590
box -6 -8 106 268
use INVX1  _2258_
timestamp 0
transform 1 0 12270 0 1 8590
box -6 -8 66 268
use OR2X2  _2259_
timestamp 0
transform -1 0 12030 0 -1 8590
box -6 -8 106 268
use NAND2X1  _2260_
timestamp 0
transform 1 0 10130 0 -1 9110
box -6 -8 86 268
use NOR2X1  _2261_
timestamp 0
transform 1 0 10390 0 -1 9110
box -6 -8 86 268
use NAND2X1  _2262_
timestamp 0
transform -1 0 10970 0 1 8070
box -6 -8 86 268
use NAND3X1  _2263_
timestamp 0
transform 1 0 11390 0 -1 8590
box -6 -8 106 268
use NOR2X1  _2264_
timestamp 0
transform 1 0 12210 0 -1 8590
box -6 -8 86 268
use OAI21X1  _2265_
timestamp 0
transform -1 0 11550 0 -1 9630
box -6 -8 106 268
use INVX1  _2266_
timestamp 0
transform -1 0 10870 0 -1 11710
box -6 -8 66 268
use NAND2X1  _2267_
timestamp 0
transform 1 0 12070 0 -1 11190
box -6 -8 86 268
use NOR2X1  _2268_
timestamp 0
transform 1 0 12210 0 1 9630
box -6 -8 86 268
use AOI22X1  _2269_
timestamp 0
transform -1 0 12090 0 -1 9630
box -6 -8 126 268
use AOI21X1  _2270_
timestamp 0
transform 1 0 11410 0 -1 9110
box -6 -8 106 268
use NAND3X1  _2271_
timestamp 0
transform -1 0 11790 0 -1 9110
box -6 -8 106 268
use INVX1  _2272_
timestamp 0
transform 1 0 11970 0 -1 9110
box -6 -8 66 268
use NAND3X1  _2273_
timestamp 0
transform -1 0 12310 0 -1 9110
box -6 -8 106 268
use AOI22X1  _2274_
timestamp 0
transform 1 0 10150 0 -1 7030
box -6 -8 126 268
use NOR2X1  _2275_
timestamp 0
transform -1 0 8370 0 -1 6510
box -6 -8 86 268
use OAI21X1  _2276_
timestamp 0
transform 1 0 8970 0 1 4430
box -6 -8 106 268
use OAI21X1  _2277_
timestamp 0
transform 1 0 9250 0 1 4430
box -6 -8 106 268
use OAI21X1  _2278_
timestamp 0
transform -1 0 9410 0 -1 4950
box -6 -8 106 268
use AOI21X1  _2279_
timestamp 0
transform 1 0 9130 0 -1 6510
box -6 -8 106 268
use AND2X2  _2280_
timestamp 0
transform 1 0 10290 0 1 6510
box -6 -8 106 268
use NAND3X1  _2281_
timestamp 0
transform 1 0 12190 0 1 6510
box -6 -8 106 268
use INVX1  _2282_
timestamp 0
transform 1 0 12230 0 -1 5990
box -6 -8 66 268
use NOR2X1  _2283_
timestamp 0
transform -1 0 11170 0 -1 6510
box -6 -8 86 268
use AND2X2  _2284_
timestamp 0
transform 1 0 12190 0 -1 5470
box -6 -8 106 268
use AND2X2  _2285_
timestamp 0
transform 1 0 12190 0 1 5470
box -6 -8 106 268
use NAND3X1  _2286_
timestamp 0
transform -1 0 12050 0 -1 5990
box -6 -8 106 268
use OR2X2  _2287_
timestamp 0
transform 1 0 11910 0 1 5990
box -6 -8 106 268
use AOI22X1  _2288_
timestamp 0
transform -1 0 11170 0 1 5990
box -6 -8 126 268
use MUX2X1  _2289_
timestamp 0
transform -1 0 10950 0 1 3390
box -6 -8 126 268
use NAND2X1  _2290_
timestamp 0
transform -1 0 11090 0 1 5470
box -6 -8 86 268
use NAND2X1  _2291_
timestamp 0
transform 1 0 11390 0 -1 3390
box -6 -8 86 268
use OAI21X1  _2292_
timestamp 0
transform 1 0 10530 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2293_
timestamp 0
transform 1 0 10810 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2294_
timestamp 0
transform 1 0 11130 0 1 3390
box -6 -8 106 268
use NOR2X1  _2295_
timestamp 0
transform 1 0 11010 0 -1 7030
box -6 -8 86 268
use NAND2X1  _2296_
timestamp 0
transform 1 0 11290 0 -1 7030
box -6 -8 86 268
use NOR2X1  _2297_
timestamp 0
transform 1 0 11930 0 1 8070
box -6 -8 86 268
use AOI22X1  _2298_
timestamp 0
transform -1 0 12130 0 1 7030
box -6 -8 126 268
use OAI21X1  _2299_
timestamp 0
transform -1 0 10670 0 -1 4430
box -6 -8 106 268
use OAI21X1  _2300_
timestamp 0
transform 1 0 10290 0 1 4430
box -6 -8 106 268
use OR2X2  _2301_
timestamp 0
transform 1 0 11910 0 1 7550
box -6 -8 106 268
use NAND3X1  _2302_
timestamp 0
transform 1 0 11850 0 -1 270
box -6 -8 106 268
use NOR2X1  _2303_
timestamp 0
transform -1 0 11890 0 -1 7030
box -6 -8 86 268
use NAND3X1  _2304_
timestamp 0
transform 1 0 11970 0 -1 6510
box -6 -8 106 268
use NOR2X1  _2305_
timestamp 0
transform 1 0 10850 0 1 9110
box -6 -8 86 268
use NAND3X1  _2306_
timestamp 0
transform -1 0 11790 0 1 9110
box -6 -8 106 268
use NAND2X1  _2307_
timestamp 0
transform 1 0 11410 0 1 8070
box -6 -8 86 268
use NOR2X1  _2308_
timestamp 0
transform 1 0 12190 0 1 8070
box -6 -8 86 268
use OAI21X1  _2309_
timestamp 0
transform -1 0 11830 0 1 8590
box -6 -8 106 268
use NAND2X1  _2310_
timestamp 0
transform -1 0 11750 0 -1 8590
box -6 -8 86 268
use INVX1  _2311_
timestamp 0
transform 1 0 11690 0 1 8070
box -6 -8 66 268
use OAI21X1  _2312_
timestamp 0
transform 1 0 11730 0 -1 8070
box -6 -8 106 268
use NOR2X1  _2313_
timestamp 0
transform 1 0 12010 0 -1 8070
box -6 -8 86 268
use NAND3X1  _2314_
timestamp 0
transform -1 0 11410 0 -1 270
box -6 -8 106 268
use OAI21X1  _2315_
timestamp 0
transform 1 0 12190 0 1 7550
box -6 -8 106 268
use NAND2X1  _2316_
timestamp 0
transform 1 0 11590 0 -1 270
box -6 -8 86 268
use INVX1  _2317_
timestamp 0
transform -1 0 12130 0 -1 7030
box -6 -8 66 268
use NAND3X1  _2318_
timestamp 0
transform 1 0 11630 0 1 5990
box -6 -8 106 268
use OR2X2  _2319_
timestamp 0
transform 1 0 11270 0 -1 5470
box -6 -8 106 268
use NAND3X1  _2320_
timestamp 0
transform 1 0 11690 0 1 4950
box -6 -8 106 268
use NOR3X1  _2321_
timestamp 0
transform 1 0 11550 0 -1 5470
box -6 -8 186 268
use INVX1  _2322_
timestamp 0
transform -1 0 11450 0 1 6510
box -6 -8 66 268
use NOR2X1  _2323_
timestamp 0
transform -1 0 11710 0 1 6510
box -6 -8 86 268
use NAND3X1  _2324_
timestamp 0
transform 1 0 11890 0 1 6510
box -6 -8 106 268
use NOR2X1  _2325_
timestamp 0
transform -1 0 12330 0 -1 6510
box -6 -8 86 268
use OAI21X1  _2326_
timestamp 0
transform 1 0 12210 0 1 5990
box -6 -8 106 268
use NAND2X1  _2327_
timestamp 0
transform 1 0 11550 0 -1 7030
box -6 -8 86 268
use NOR2X1  _2328_
timestamp 0
transform 1 0 11130 0 1 6510
box -6 -8 86 268
use NAND3X1  _2329_
timestamp 0
transform 1 0 8650 0 1 4950
box -6 -8 106 268
use AND2X2  _2330_
timestamp 0
transform -1 0 10410 0 1 4950
box -6 -8 106 268
use NAND3X1  _2331_
timestamp 0
transform -1 0 9850 0 1 4950
box -6 -8 106 268
use NAND3X1  _2332_
timestamp 0
transform -1 0 12070 0 1 4950
box -6 -8 106 268
use OR2X2  _2333_
timestamp 0
transform -1 0 10950 0 1 4950
box -6 -8 106 268
use NOR2X1  _2334_
timestamp 0
transform 1 0 10590 0 1 4950
box -6 -8 86 268
use AND2X2  _2335_
timestamp 0
transform 1 0 10570 0 1 6510
box -6 -8 106 268
use NOR2X1  _2336_
timestamp 0
transform 1 0 10750 0 -1 7030
box -6 -8 86 268
use NAND3X1  _2337_
timestamp 0
transform -1 0 10950 0 1 6510
box -6 -8 106 268
use AND2X2  _2338_
timestamp 0
transform -1 0 10870 0 1 5990
box -6 -8 106 268
use NAND3X1  _2339_
timestamp 0
transform -1 0 9790 0 -1 6510
box -6 -8 106 268
use INVX1  _2340_
timestamp 0
transform -1 0 10050 0 -1 5470
box -6 -8 66 268
use OAI21X1  _2341_
timestamp 0
transform 1 0 9690 0 -1 5470
box -6 -8 106 268
use OAI21X1  _2342_
timestamp 0
transform -1 0 10650 0 -1 3910
box -6 -8 106 268
use NOR2X1  _2343_
timestamp 0
transform -1 0 10570 0 -1 5470
box -6 -8 86 268
use NAND3X1  _2344_
timestamp 0
transform -1 0 10830 0 1 5470
box -6 -8 106 268
use NAND2X1  _2345_
timestamp 0
transform 1 0 11870 0 -1 4950
box -6 -8 86 268
use NOR2X1  _2346_
timestamp 0
transform 1 0 11610 0 -1 4950
box -6 -8 86 268
use AOI21X1  _2347_
timestamp 0
transform -1 0 9030 0 1 5470
box -6 -8 106 268
use AND2X2  _2348_
timestamp 0
transform -1 0 10130 0 1 4950
box -6 -8 106 268
use NOR2X1  _2349_
timestamp 0
transform -1 0 11770 0 1 3910
box -6 -8 86 268
use NAND3X1  _2350_
timestamp 0
transform -1 0 11510 0 1 4950
box -6 -8 106 268
use NOR2X1  _2351_
timestamp 0
transform -1 0 10550 0 1 5470
box -6 -8 86 268
use NAND3X1  _2352_
timestamp 0
transform -1 0 10330 0 -1 6510
box -6 -8 106 268
use OR2X2  _2353_
timestamp 0
transform -1 0 9630 0 1 6510
box -6 -8 106 268
use INVX1  _2354_
timestamp 0
transform 1 0 7950 0 -1 10670
box -6 -8 66 268
use OAI21X1  _2355_
timestamp 0
transform -1 0 7130 0 -1 5990
box -6 -8 106 268
use INVX2  _2356_
timestamp 0
transform -1 0 7010 0 -1 6510
box -6 -8 66 268
use INVX1  _2357_
timestamp 0
transform -1 0 7670 0 1 3390
box -6 -8 66 268
use NAND3X1  _2358_
timestamp 0
transform -1 0 7290 0 -1 6510
box -6 -8 106 268
use OAI21X1  _2359_
timestamp 0
transform 1 0 7430 0 -1 10670
box -6 -8 106 268
use INVX1  _2360_
timestamp 0
transform -1 0 8150 0 -1 11190
box -6 -8 66 268
use OAI21X1  _2361_
timestamp 0
transform -1 0 7250 0 -1 10670
box -6 -8 106 268
use INVX1  _2362_
timestamp 0
transform 1 0 8890 0 1 10150
box -6 -8 66 268
use NOR2X1  _2363_
timestamp 0
transform -1 0 7630 0 1 3910
box -6 -8 86 268
use INVX1  _2364_
timestamp 0
transform 1 0 7310 0 1 3910
box -6 -8 66 268
use OAI21X1  _2365_
timestamp 0
transform 1 0 7030 0 1 3910
box -6 -8 106 268
use INVX2  _2366_
timestamp 0
transform 1 0 6510 0 1 3910
box -6 -8 66 268
use NOR2X1  _2367_
timestamp 0
transform -1 0 7410 0 -1 4430
box -6 -8 86 268
use NAND3X1  _2368_
timestamp 0
transform 1 0 6750 0 1 3910
box -6 -8 106 268
use AOI21X1  _2369_
timestamp 0
transform 1 0 7130 0 1 4430
box -6 -8 106 268
use OAI21X1  _2370_
timestamp 0
transform -1 0 7490 0 1 10150
box -6 -8 106 268
use INVX1  _2371_
timestamp 0
transform 1 0 7330 0 -1 11190
box -6 -8 66 268
use NOR2X1  _2372_
timestamp 0
transform -1 0 6970 0 -1 10670
box -6 -8 86 268
use NOR2X1  _2373_
timestamp 0
transform 1 0 6850 0 -1 4950
box -6 -8 86 268
use OAI21X1  _2374_
timestamp 0
transform 1 0 8350 0 1 3910
box -6 -8 106 268
use OAI21X1  _2375_
timestamp 0
transform 1 0 8410 0 -1 3910
box -6 -8 106 268
use NAND2X1  _2376_
timestamp 0
transform -1 0 6910 0 -1 3910
box -6 -8 86 268
use NAND2X1  _2377_
timestamp 0
transform 1 0 5550 0 -1 4950
box -6 -8 86 268
use OAI21X1  _2378_
timestamp 0
transform -1 0 3950 0 -1 4950
box -6 -8 106 268
use NAND2X1  _2379_
timestamp 0
transform -1 0 8190 0 -1 3390
box -6 -8 86 268
use OAI21X1  _2380_
timestamp 0
transform -1 0 5850 0 1 5470
box -6 -8 106 268
use INVX1  _2381_
timestamp 0
transform -1 0 6090 0 1 5470
box -6 -8 66 268
use OAI21X1  _2382_
timestamp 0
transform -1 0 5990 0 -1 5470
box -6 -8 106 268
use NAND2X1  _2383_
timestamp 0
transform 1 0 4830 0 1 6510
box -6 -8 86 268
use OAI21X1  _2384_
timestamp 0
transform 1 0 4770 0 1 5990
box -6 -8 106 268
use AOI21X1  _2385_
timestamp 0
transform 1 0 4990 0 1 5470
box -6 -8 106 268
use NAND3X1  _2386_
timestamp 0
transform 1 0 5270 0 -1 4950
box -6 -8 106 268
use NAND2X1  _2387_
timestamp 0
transform 1 0 1790 0 1 5470
box -6 -8 86 268
use OAI21X1  _2388_
timestamp 0
transform 1 0 1730 0 -1 5470
box -6 -8 106 268
use NAND2X1  _2389_
timestamp 0
transform 1 0 5310 0 1 5990
box -6 -8 86 268
use OAI21X1  _2390_
timestamp 0
transform 1 0 2590 0 1 5990
box -6 -8 106 268
use AOI21X1  _2391_
timestamp 0
transform -1 0 2470 0 -1 5990
box -6 -8 106 268
use NAND3X1  _2392_
timestamp 0
transform -1 0 2190 0 -1 5990
box -6 -8 106 268
use NAND2X1  _2393_
timestamp 0
transform -1 0 2730 0 -1 5990
box -6 -8 86 268
use OAI21X1  _2394_
timestamp 0
transform -1 0 3170 0 -1 5470
box -6 -8 106 268
use NAND2X1  _2395_
timestamp 0
transform 1 0 4490 0 1 5990
box -6 -8 86 268
use OAI21X1  _2396_
timestamp 0
transform 1 0 3130 0 1 5990
box -6 -8 106 268
use AOI21X1  _2397_
timestamp 0
transform -1 0 3290 0 -1 5990
box -6 -8 106 268
use NAND3X1  _2398_
timestamp 0
transform -1 0 3010 0 -1 5990
box -6 -8 106 268
use NAND2X1  _2399_
timestamp 0
transform 1 0 2050 0 1 5990
box -6 -8 86 268
use OAI21X1  _2400_
timestamp 0
transform -1 0 1550 0 -1 5470
box -6 -8 106 268
use NAND2X1  _2401_
timestamp 0
transform -1 0 3010 0 1 6510
box -6 -8 86 268
use OAI21X1  _2402_
timestamp 0
transform 1 0 2690 0 -1 6510
box -6 -8 106 268
use AOI21X1  _2403_
timestamp 0
transform -1 0 2410 0 1 5990
box -6 -8 106 268
use NAND3X1  _2404_
timestamp 0
transform -1 0 1850 0 1 5990
box -6 -8 106 268
use INVX1  _2405_
timestamp 0
transform -1 0 1670 0 1 6510
box -6 -8 66 268
use OAI22X1  _2406_
timestamp 0
transform 1 0 6010 0 -1 3910
box -6 -8 126 268
use AOI21X1  _2407_
timestamp 0
transform -1 0 4450 0 -1 3910
box -6 -8 106 268
use OAI21X1  _2408_
timestamp 0
transform -1 0 5810 0 1 3390
box -6 -8 106 268
use OAI21X1  _2409_
timestamp 0
transform -1 0 6630 0 1 3390
box -6 -8 106 268
use AOI22X1  _2410_
timestamp 0
transform -1 0 4430 0 1 3390
box -6 -8 126 268
use AND2X2  _2411_
timestamp 0
transform -1 0 4170 0 -1 3910
box -6 -8 106 268
use OAI21X1  _2412_
timestamp 0
transform -1 0 1430 0 1 6510
box -6 -8 106 268
use AOI22X1  _2413_
timestamp 0
transform -1 0 4730 0 1 3390
box -6 -8 126 268
use OAI21X1  _2414_
timestamp 0
transform 1 0 3170 0 1 5470
box -6 -8 106 268
use NOR2X1  _2415_
timestamp 0
transform -1 0 2950 0 1 5990
box -6 -8 86 268
use OAI21X1  _2416_
timestamp 0
transform 1 0 1850 0 1 6510
box -6 -8 106 268
use NAND2X1  _2417_
timestamp 0
transform -1 0 2410 0 1 5470
box -6 -8 86 268
use OAI21X1  _2418_
timestamp 0
transform -1 0 2310 0 1 4950
box -6 -8 106 268
use NAND2X1  _2419_
timestamp 0
transform -1 0 3610 0 -1 6510
box -6 -8 86 268
use OAI21X1  _2420_
timestamp 0
transform 1 0 2970 0 -1 6510
box -6 -8 106 268
use AOI21X1  _2421_
timestamp 0
transform -1 0 2970 0 1 5470
box -6 -8 106 268
use NAND3X1  _2422_
timestamp 0
transform -1 0 2150 0 1 5470
box -6 -8 106 268
use NAND2X1  _2423_
timestamp 0
transform -1 0 3830 0 -1 5990
box -6 -8 86 268
use OAI21X1  _2424_
timestamp 0
transform -1 0 3690 0 -1 5470
box -6 -8 106 268
use NAND2X1  _2425_
timestamp 0
transform -1 0 3550 0 1 6510
box -6 -8 86 268
use OAI21X1  _2426_
timestamp 0
transform 1 0 3250 0 -1 6510
box -6 -8 106 268
use AOI21X1  _2427_
timestamp 0
transform 1 0 3410 0 1 5990
box -6 -8 106 268
use NAND3X1  _2428_
timestamp 0
transform -1 0 3570 0 -1 5990
box -6 -8 106 268
use INVX1  _2429_
timestamp 0
transform -1 0 5270 0 -1 3910
box -6 -8 66 268
use OAI21X1  _2430_
timestamp 0
transform -1 0 7990 0 -1 3910
box -6 -8 106 268
use OR2X2  _2431_
timestamp 0
transform -1 0 5550 0 -1 3910
box -6 -8 106 268
use NAND2X1  _2432_
timestamp 0
transform -1 0 9650 0 -1 2350
box -6 -8 86 268
use NOR2X1  _2433_
timestamp 0
transform 1 0 11690 0 -1 2870
box -6 -8 86 268
use NAND3X1  _2434_
timestamp 0
transform 1 0 10870 0 -1 2870
box -6 -8 106 268
use OR2X2  _2435_
timestamp 0
transform -1 0 7430 0 1 3390
box -6 -8 106 268
use NOR2X1  _2436_
timestamp 0
transform -1 0 7090 0 -1 3390
box -6 -8 86 268
use NAND3X1  _2437_
timestamp 0
transform -1 0 9790 0 -1 3390
box -6 -8 106 268
use NOR2X1  _2438_
timestamp 0
transform -1 0 9510 0 -1 3390
box -6 -8 86 268
use NAND2X1  _2439_
timestamp 0
transform -1 0 6290 0 -1 3390
box -6 -8 86 268
use NAND2X1  _2440_
timestamp 0
transform 1 0 7850 0 -1 1830
box -6 -8 86 268
use NAND3X1  _2441_
timestamp 0
transform -1 0 7770 0 -1 2870
box -6 -8 106 268
use NOR2X1  _2442_
timestamp 0
transform 1 0 10390 0 1 1310
box -6 -8 86 268
use NAND2X1  _2443_
timestamp 0
transform -1 0 7370 0 -1 1830
box -6 -8 86 268
use NAND3X1  _2444_
timestamp 0
transform -1 0 7370 0 -1 3390
box -6 -8 106 268
use NOR2X1  _2445_
timestamp 0
transform 1 0 5390 0 -1 3390
box -6 -8 86 268
use OAI21X1  _2446_
timestamp 0
transform 1 0 6510 0 -1 4430
box -6 -8 106 268
use NOR2X1  _2447_
timestamp 0
transform -1 0 4950 0 -1 4430
box -6 -8 86 268
use OAI21X1  _2448_
timestamp 0
transform -1 0 6570 0 -1 3390
box -6 -8 106 268
use NAND3X1  _2449_
timestamp 0
transform -1 0 7190 0 -1 3910
box -6 -8 106 268
use NOR2X1  _2450_
timestamp 0
transform 1 0 4250 0 1 3910
box -6 -8 86 268
use INVX2  _2451_
timestamp 0
transform -1 0 4170 0 -1 4430
box -6 -8 66 268
use INVX1  _2452_
timestamp 0
transform 1 0 4770 0 1 4430
box -6 -8 66 268
use OAI21X1  _2453_
timestamp 0
transform 1 0 8630 0 1 3910
box -6 -8 106 268
use INVX1  _2454_
timestamp 0
transform 1 0 4510 0 1 3910
box -6 -8 66 268
use NAND2X1  _2455_
timestamp 0
transform 1 0 4510 0 1 4430
box -6 -8 86 268
use NOR2X1  _2456_
timestamp 0
transform -1 0 4430 0 -1 4430
box -6 -8 86 268
use NAND2X1  _2457_
timestamp 0
transform -1 0 4690 0 -1 4430
box -6 -8 86 268
use OAI21X1  _2458_
timestamp 0
transform -1 0 5090 0 -1 4950
box -6 -8 106 268
use AOI22X1  _2459_
timestamp 0
transform 1 0 5130 0 -1 4430
box -6 -8 126 268
use AND2X2  _2460_
timestamp 0
transform 1 0 5010 0 1 4430
box -6 -8 106 268
use OAI21X1  _2461_
timestamp 0
transform 1 0 5290 0 1 4430
box -6 -8 106 268
use AOI21X1  _2462_
timestamp 0
transform 1 0 5430 0 -1 4430
box -6 -8 106 268
use INVX1  _2463_
timestamp 0
transform 1 0 6370 0 1 790
box -6 -8 66 268
use OAI21X1  _2464_
timestamp 0
transform -1 0 3390 0 -1 4950
box -6 -8 106 268
use AOI22X1  _2465_
timestamp 0
transform -1 0 3130 0 -1 4430
box -6 -8 126 268
use AND2X2  _2466_
timestamp 0
transform -1 0 3110 0 -1 4950
box -6 -8 106 268
use OAI21X1  _2467_
timestamp 0
transform 1 0 2170 0 -1 4950
box -6 -8 106 268
use AOI21X1  _2468_
timestamp 0
transform -1 0 1810 0 1 4430
box -6 -8 106 268
use INVX1  _2469_
timestamp 0
transform 1 0 690 0 -1 4430
box -6 -8 66 268
use OAI21X1  _2470_
timestamp 0
transform -1 0 2870 0 1 4950
box -6 -8 106 268
use AOI22X1  _2471_
timestamp 0
transform -1 0 2910 0 1 4430
box -6 -8 126 268
use AND2X2  _2472_
timestamp 0
transform -1 0 2590 0 1 4950
box -6 -8 106 268
use OAI21X1  _2473_
timestamp 0
transform 1 0 2030 0 -1 5470
box -6 -8 106 268
use AOI21X1  _2474_
timestamp 0
transform -1 0 1610 0 1 5470
box -6 -8 106 268
use INVX1  _2475_
timestamp 0
transform -1 0 510 0 1 5470
box -6 -8 66 268
use INVX1  _2476_
timestamp 0
transform -1 0 3930 0 -1 4430
box -6 -8 66 268
use OR2X2  _2477_
timestamp 0
transform -1 0 5210 0 -1 3390
box -6 -8 106 268
use NOR2X1  _2478_
timestamp 0
transform 1 0 3990 0 1 3910
box -6 -8 86 268
use NAND2X1  _2479_
timestamp 0
transform -1 0 3690 0 -1 4430
box -6 -8 86 268
use INVX1  _2480_
timestamp 0
transform 1 0 1870 0 1 3390
box -6 -8 66 268
use OAI22X1  _2481_
timestamp 0
transform -1 0 3530 0 1 3910
box -6 -8 126 268
use AOI21X1  _2482_
timestamp 0
transform 1 0 3710 0 1 3910
box -6 -8 106 268
use OAI21X1  _2483_
timestamp 0
transform 1 0 3130 0 1 3910
box -6 -8 106 268
use AOI21X1  _2484_
timestamp 0
transform 1 0 2850 0 1 3910
box -6 -8 106 268
use INVX1  _2485_
timestamp 0
transform -1 0 510 0 1 3910
box -6 -8 66 268
use OAI21X1  _2486_
timestamp 0
transform -1 0 2830 0 -1 4950
box -6 -8 106 268
use AOI22X1  _2487_
timestamp 0
transform 1 0 2490 0 1 4430
box -6 -8 126 268
use AND2X2  _2488_
timestamp 0
transform -1 0 2550 0 -1 4950
box -6 -8 106 268
use OAI21X1  _2489_
timestamp 0
transform -1 0 1990 0 -1 4950
box -6 -8 106 268
use AOI21X1  _2490_
timestamp 0
transform -1 0 1550 0 1 4950
box -6 -8 106 268
use INVX1  _2491_
timestamp 0
transform -1 0 510 0 1 4950
box -6 -8 66 268
use OAI21X1  _2492_
timestamp 0
transform 1 0 4690 0 -1 4950
box -6 -8 106 268
use INVX1  _2493_
timestamp 0
transform 1 0 3690 0 1 4430
box -6 -8 66 268
use INVX2  _2494_
timestamp 0
transform 1 0 6270 0 1 3910
box -6 -8 66 268
use OAI22X1  _2495_
timestamp 0
transform 1 0 3930 0 1 4430
box -6 -8 126 268
use AOI21X1  _2496_
timestamp 0
transform 1 0 4230 0 1 4430
box -6 -8 106 268
use AND2X2  _2497_
timestamp 0
transform -1 0 4230 0 -1 4950
box -6 -8 106 268
use OAI21X1  _2498_
timestamp 0
transform 1 0 3610 0 1 4950
box -6 -8 106 268
use AOI21X1  _2499_
timestamp 0
transform 1 0 3870 0 -1 5470
box -6 -8 106 268
use INVX1  _2500_
timestamp 0
transform -1 0 510 0 -1 5470
box -6 -8 66 268
use INVX1  _2501_
timestamp 0
transform -1 0 3510 0 1 5470
box -6 -8 66 268
use AOI22X1  _2502_
timestamp 0
transform -1 0 3230 0 1 4430
box -6 -8 126 268
use OAI21X1  _2503_
timestamp 0
transform -1 0 3670 0 -1 4950
box -6 -8 106 268
use AOI21X1  _2504_
timestamp 0
transform -1 0 3430 0 1 4950
box -6 -8 106 268
use OAI21X1  _2505_
timestamp 0
transform 1 0 2790 0 -1 5470
box -6 -8 106 268
use AOI21X1  _2506_
timestamp 0
transform -1 0 2690 0 1 5470
box -6 -8 106 268
use INVX1  _2507_
timestamp 0
transform 1 0 730 0 -1 5990
box -6 -8 66 268
use NAND2X1  _2508_
timestamp 0
transform 1 0 3230 0 1 3390
box -6 -8 86 268
use INVX1  _2509_
timestamp 0
transform 1 0 2770 0 -1 4430
box -6 -8 66 268
use OAI22X1  _2510_
timestamp 0
transform -1 0 3430 0 -1 4430
box -6 -8 126 268
use AOI21X1  _2511_
timestamp 0
transform 1 0 3410 0 1 4430
box -6 -8 106 268
use NAND2X1  _2512_
timestamp 0
transform 1 0 3250 0 -1 3910
box -6 -8 86 268
use INVX1  _2513_
timestamp 0
transform -1 0 2550 0 -1 3910
box -6 -8 66 268
use OAI21X1  _2514_
timestamp 0
transform 1 0 2210 0 -1 3910
box -6 -8 106 268
use AOI21X1  _2515_
timestamp 0
transform -1 0 2310 0 -1 4430
box -6 -8 106 268
use INVX1  _2516_
timestamp 0
transform -1 0 510 0 -1 4430
box -6 -8 66 268
use INVX1  _2517_
timestamp 0
transform -1 0 2370 0 1 270
box -6 -8 66 268
use NOR2X1  _2518_
timestamp 0
transform 1 0 5410 0 -1 270
box -6 -8 86 268
use AOI21X1  _2519_
timestamp 0
transform -1 0 6030 0 -1 3390
box -6 -8 106 268
use INVX1  _2520_
timestamp 0
transform -1 0 6090 0 1 3910
box -6 -8 66 268
use OAI21X1  _2521_
timestamp 0
transform 1 0 5750 0 1 3910
box -6 -8 106 268
use AOI21X1  _2522_
timestamp 0
transform -1 0 5830 0 -1 3910
box -6 -8 106 268
use NAND3X1  _2523_
timestamp 0
transform -1 0 5750 0 -1 3390
box -6 -8 106 268
use OR2X2  _2524_
timestamp 0
transform -1 0 5690 0 1 270
box -6 -8 106 268
use INVX1  _2525_
timestamp 0
transform -1 0 2870 0 -1 270
box -6 -8 66 268
use INVX2  _2526_
timestamp 0
transform 1 0 6230 0 1 2870
box -6 -8 66 268
use AOI21X1  _2527_
timestamp 0
transform 1 0 6630 0 -1 1310
box -6 -8 106 268
use OAI21X1  _2528_
timestamp 0
transform 1 0 6610 0 1 790
box -6 -8 106 268
use AOI21X1  _2529_
timestamp 0
transform 1 0 6210 0 -1 790
box -6 -8 106 268
use OAI21X1  _2530_
timestamp 0
transform 1 0 5670 0 -1 270
box -6 -8 106 268
use INVX1  _2531_
timestamp 0
transform 1 0 3030 0 1 270
box -6 -8 66 268
use INVX1  _2532_
timestamp 0
transform 1 0 4330 0 1 270
box -6 -8 66 268
use AOI22X1  _2533_
timestamp 0
transform 1 0 5250 0 1 790
box -6 -8 126 268
use OAI21X1  _2534_
timestamp 0
transform 1 0 4970 0 1 790
box -6 -8 106 268
use AOI21X1  _2535_
timestamp 0
transform -1 0 4790 0 1 790
box -6 -8 106 268
use OAI21X1  _2536_
timestamp 0
transform 1 0 3550 0 1 270
box -6 -8 106 268
use INVX1  _2537_
timestamp 0
transform 1 0 2190 0 -1 1310
box -6 -8 66 268
use NAND2X1  _2538_
timestamp 0
transform 1 0 4590 0 1 2870
box -6 -8 86 268
use AOI22X1  _2539_
timestamp 0
transform 1 0 3970 0 -1 3390
box -6 -8 126 268
use AND2X2  _2540_
timestamp 0
transform 1 0 4310 0 1 2870
box -6 -8 106 268
use OAI21X1  _2541_
timestamp 0
transform -1 0 4370 0 -1 3390
box -6 -8 106 268
use INVX1  _2542_
timestamp 0
transform -1 0 3850 0 -1 1310
box -6 -8 66 268
use OAI21X1  _2543_
timestamp 0
transform 1 0 3570 0 1 790
box -6 -8 106 268
use INVX1  _2544_
timestamp 0
transform 1 0 4290 0 -1 1830
box -6 -8 66 268
use INVX1  _2545_
timestamp 0
transform 1 0 4550 0 -1 1310
box -6 -8 66 268
use INVX1  _2546_
timestamp 0
transform 1 0 4930 0 1 3390
box -6 -8 66 268
use OAI21X1  _2547_
timestamp 0
transform -1 0 4930 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2548_
timestamp 0
transform -1 0 4650 0 -1 3390
box -6 -8 106 268
use AOI21X1  _2549_
timestamp 0
transform 1 0 4790 0 1 1830
box -6 -8 106 268
use OAI21X1  _2550_
timestamp 0
transform 1 0 4790 0 -1 1830
box -6 -8 106 268
use INVX1  _2551_
timestamp 0
transform 1 0 5310 0 1 1310
box -6 -8 66 268
use OAI21X1  _2552_
timestamp 0
transform 1 0 5550 0 1 1310
box -6 -8 106 268
use INVX1  _2553_
timestamp 0
transform 1 0 2450 0 1 1310
box -6 -8 66 268
use INVX1  _2554_
timestamp 0
transform 1 0 4590 0 -1 790
box -6 -8 66 268
use INVX1  _2555_
timestamp 0
transform -1 0 4810 0 1 3910
box -6 -8 66 268
use OAI21X1  _2556_
timestamp 0
transform -1 0 5090 0 -1 2870
box -6 -8 106 268
use OAI21X1  _2557_
timestamp 0
transform 1 0 4710 0 -1 2870
box -6 -8 106 268
use AOI21X1  _2558_
timestamp 0
transform 1 0 4790 0 1 1310
box -6 -8 106 268
use OAI21X1  _2559_
timestamp 0
transform 1 0 4510 0 1 1310
box -6 -8 106 268
use INVX1  _2560_
timestamp 0
transform 1 0 4010 0 1 1310
box -6 -8 66 268
use OAI21X1  _2561_
timestamp 0
transform 1 0 3730 0 1 1310
box -6 -8 106 268
use INVX1  _2562_
timestamp 0
transform 1 0 2330 0 -1 2350
box -6 -8 66 268
use AOI21X1  _2563_
timestamp 0
transform -1 0 4630 0 1 2350
box -6 -8 106 268
use OAI21X1  _2564_
timestamp 0
transform 1 0 4470 0 -1 2350
box -6 -8 106 268
use AOI21X1  _2565_
timestamp 0
transform -1 0 4030 0 -1 2350
box -6 -8 106 268
use OAI21X1  _2566_
timestamp 0
transform 1 0 2550 0 1 1830
box -6 -8 106 268
use INVX1  _2567_
timestamp 0
transform 1 0 4030 0 -1 1310
box -6 -8 66 268
use INVX1  _2568_
timestamp 0
transform -1 0 5870 0 -1 2870
box -6 -8 66 268
use OAI21X1  _2569_
timestamp 0
transform -1 0 6050 0 1 2870
box -6 -8 106 268
use OAI21X1  _2570_
timestamp 0
transform 1 0 6050 0 -1 2870
box -6 -8 106 268
use NOR2X1  _2571_
timestamp 0
transform 1 0 6050 0 -1 2350
box -6 -8 86 268
use OAI21X1  _2572_
timestamp 0
transform 1 0 5910 0 1 1830
box -6 -8 106 268
use INVX1  _2573_
timestamp 0
transform 1 0 5830 0 1 1310
box -6 -8 66 268
use OAI21X1  _2574_
timestamp 0
transform 1 0 5810 0 -1 1310
box -6 -8 106 268
use AND2X2  _2575_
timestamp 0
transform -1 0 4930 0 1 7550
box -6 -8 106 268
use INVX1  _2576_
timestamp 0
transform -1 0 4390 0 1 7550
box -6 -8 66 268
use NOR2X1  _2577_
timestamp 0
transform -1 0 4650 0 1 7550
box -6 -8 86 268
use INVX1  _2578_
timestamp 0
transform 1 0 7090 0 -1 11190
box -6 -8 66 268
use NOR2X1  _2579_
timestamp 0
transform 1 0 7110 0 1 10150
box -6 -8 86 268
use INVX8  _2580_
timestamp 0
transform 1 0 8110 0 1 11190
box -6 -8 126 268
use OAI21X1  _2581_
timestamp 0
transform -1 0 9050 0 1 1830
box -6 -8 106 268
use OAI21X1  _2582_
timestamp 0
transform 1 0 7010 0 1 1830
box -6 -8 106 268
use AOI21X1  _2583_
timestamp 0
transform -1 0 7090 0 -1 1830
box -6 -8 106 268
use OAI21X1  _2584_
timestamp 0
transform 1 0 7430 0 1 1310
box -6 -8 106 268
use OAI21X1  _2585_
timestamp 0
transform 1 0 7470 0 -1 1310
box -6 -8 106 268
use NAND3X1  _2586_
timestamp 0
transform -1 0 8630 0 1 1310
box -6 -8 106 268
use NOR2X1  _2587_
timestamp 0
transform -1 0 6950 0 1 1310
box -6 -8 86 268
use NAND2X1  _2588_
timestamp 0
transform -1 0 5990 0 -1 1830
box -6 -8 86 268
use OAI22X1  _2589_
timestamp 0
transform 1 0 7550 0 -1 1830
box -6 -8 126 268
use NAND3X1  _2590_
timestamp 0
transform -1 0 6410 0 -1 2350
box -6 -8 106 268
use NAND3X1  _2591_
timestamp 0
transform 1 0 6590 0 1 1310
box -6 -8 106 268
use NOR2X1  _2592_
timestamp 0
transform -1 0 4610 0 -1 1830
box -6 -8 86 268
use INVX2  _2593_
timestamp 0
transform 1 0 5070 0 1 1310
box -6 -8 66 268
use NOR3X1  _2594_
timestamp 0
transform -1 0 8810 0 1 790
box -6 -8 186 268
use AOI22X1  _2595_
timestamp 0
transform -1 0 5470 0 1 1830
box -6 -8 126 268
use AND2X2  _2596_
timestamp 0
transform 1 0 5370 0 1 2870
box -6 -8 106 268
use NOR2X1  _2597_
timestamp 0
transform 1 0 5550 0 -1 2870
box -6 -8 86 268
use OAI21X1  _2598_
timestamp 0
transform -1 0 5370 0 -1 2870
box -6 -8 106 268
use NAND3X1  _2599_
timestamp 0
transform -1 0 5170 0 1 1830
box -6 -8 106 268
use NAND2X1  _2600_
timestamp 0
transform -1 0 5150 0 -1 1830
box -6 -8 86 268
use AOI21X1  _2601_
timestamp 0
transform -1 0 5430 0 -1 1830
box -6 -8 106 268
use NAND3X1  _2602_
timestamp 0
transform -1 0 8370 0 -1 790
box -6 -8 106 268
use OAI21X1  _2603_
timestamp 0
transform -1 0 6810 0 -1 1830
box -6 -8 106 268
use INVX1  _2604_
timestamp 0
transform -1 0 6530 0 -1 1830
box -6 -8 66 268
use OAI21X1  _2605_
timestamp 0
transform 1 0 6190 0 -1 1830
box -6 -8 106 268
use NAND2X1  _2606_
timestamp 0
transform -1 0 5730 0 1 1830
box -6 -8 86 268
use NOR2X1  _2607_
timestamp 0
transform 1 0 5830 0 1 2350
box -6 -8 86 268
use AOI22X1  _2608_
timestamp 0
transform 1 0 5650 0 1 2870
box -6 -8 126 268
use AOI22X1  _2609_
timestamp 0
transform -1 0 5730 0 -1 1830
box -6 -8 126 268
use INVX1  _2610_
timestamp 0
transform 1 0 5010 0 -1 2350
box -6 -8 66 268
use NAND2X1  _2611_
timestamp 0
transform -1 0 5330 0 -1 2350
box -6 -8 86 268
use OAI22X1  _2612_
timestamp 0
transform -1 0 5630 0 -1 2350
box -6 -8 126 268
use INVX2  _2613_
timestamp 0
transform -1 0 1390 0 -1 2350
box -6 -8 66 268
use NAND2X1  _2614_
timestamp 0
transform 1 0 2330 0 1 2870
box -6 -8 86 268
use OAI21X1  _2615_
timestamp 0
transform -1 0 2690 0 -1 2870
box -6 -8 106 268
use AOI21X1  _2616_
timestamp 0
transform -1 0 2670 0 -1 2350
box -6 -8 106 268
use OAI21X1  _2617_
timestamp 0
transform 1 0 1570 0 -1 2350
box -6 -8 106 268
use NOR2X1  _2618_
timestamp 0
transform 1 0 990 0 -1 1830
box -6 -8 86 268
use NAND2X1  _2619_
timestamp 0
transform -1 0 550 0 1 1830
box -6 -8 86 268
use NAND2X1  _2620_
timestamp 0
transform -1 0 810 0 -1 1310
box -6 -8 86 268
use OAI22X1  _2621_
timestamp 0
transform 1 0 1050 0 1 1310
box -6 -8 126 268
use NAND2X1  _2622_
timestamp 0
transform 1 0 490 0 1 1310
box -6 -8 86 268
use NOR2X1  _2623_
timestamp 0
transform 1 0 2870 0 -1 2870
box -6 -8 86 268
use NAND2X1  _2624_
timestamp 0
transform 1 0 2070 0 1 2870
box -6 -8 86 268
use OAI21X1  _2625_
timestamp 0
transform -1 0 2410 0 -1 2870
box -6 -8 106 268
use AOI21X1  _2626_
timestamp 0
transform -1 0 2130 0 -1 2870
box -6 -8 106 268
use OAI21X1  _2627_
timestamp 0
transform 1 0 190 0 1 1830
box -6 -8 106 268
use XOR2X1  _2628_
timestamp 0
transform 1 0 190 0 1 1310
box -6 -8 126 268
use OAI21X1  _2629_
timestamp 0
transform -1 0 530 0 -1 1310
box -6 -8 106 268
use INVX1  _2630_
timestamp 0
transform 1 0 190 0 -1 1310
box -6 -8 66 268
use INVX2  _2631_
timestamp 0
transform 1 0 5130 0 1 2870
box -6 -8 66 268
use OAI21X1  _2632_
timestamp 0
transform 1 0 2370 0 -1 3390
box -6 -8 106 268
use AOI21X1  _2633_
timestamp 0
transform -1 0 2750 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2634_
timestamp 0
transform -1 0 290 0 -1 2870
box -6 -8 106 268
use AOI21X1  _2635_
timestamp 0
transform 1 0 210 0 -1 1830
box -6 -8 106 268
use NAND2X1  _2636_
timestamp 0
transform 1 0 730 0 -1 1830
box -6 -8 86 268
use NAND2X1  _2637_
timestamp 0
transform 1 0 1070 0 -1 2350
box -6 -8 86 268
use AOI22X1  _2638_
timestamp 0
transform 1 0 490 0 -1 2350
box -6 -8 126 268
use NAND3X1  _2639_
timestamp 0
transform -1 0 890 0 -1 2350
box -6 -8 106 268
use NAND2X1  _2640_
timestamp 0
transform -1 0 270 0 1 2350
box -6 -8 86 268
use OAI22X1  _2641_
timestamp 0
transform -1 0 310 0 -1 2350
box -6 -8 126 268
use NAND2X1  _2642_
timestamp 0
transform 1 0 1450 0 1 3910
box -6 -8 86 268
use INVX1  _2643_
timestamp 0
transform -1 0 2030 0 -1 3910
box -6 -8 66 268
use OAI21X1  _2644_
timestamp 0
transform 1 0 2390 0 1 3390
box -6 -8 106 268
use AOI21X1  _2645_
timestamp 0
transform -1 0 2210 0 1 3390
box -6 -8 106 268
use OAI21X1  _2646_
timestamp 0
transform -1 0 1410 0 -1 3390
box -6 -8 106 268
use XOR2X1  _2647_
timestamp 0
transform 1 0 190 0 -1 3910
box -6 -8 126 268
use OAI21X1  _2648_
timestamp 0
transform 1 0 690 0 1 3910
box -6 -8 106 268
use INVX1  _2649_
timestamp 0
transform 1 0 210 0 -1 3390
box -6 -8 66 268
use OAI21X1  _2650_
timestamp 0
transform -1 0 3870 0 1 3390
box -6 -8 106 268
use AOI21X1  _2651_
timestamp 0
transform -1 0 3590 0 1 3390
box -6 -8 106 268
use OAI21X1  _2652_
timestamp 0
transform 1 0 730 0 -1 3390
box -6 -8 106 268
use AOI21X1  _2653_
timestamp 0
transform 1 0 450 0 -1 3390
box -6 -8 106 268
use NAND2X1  _2654_
timestamp 0
transform 1 0 1330 0 1 3390
box -6 -8 86 268
use NAND2X1  _2655_
timestamp 0
transform 1 0 770 0 1 3390
box -6 -8 86 268
use AOI22X1  _2656_
timestamp 0
transform -1 0 1150 0 1 3390
box -6 -8 126 268
use INVX1  _2657_
timestamp 0
transform 1 0 190 0 1 2870
box -6 -8 66 268
use OAI21X1  _2658_
timestamp 0
transform 1 0 190 0 1 3390
box -6 -8 106 268
use OAI22X1  _2659_
timestamp 0
transform -1 0 590 0 1 3390
box -6 -8 126 268
use NOR2X1  _2660_
timestamp 0
transform 1 0 430 0 1 2870
box -6 -8 86 268
use INVX1  _2661_
timestamp 0
transform -1 0 2790 0 -1 3910
box -6 -8 66 268
use OAI21X1  _2662_
timestamp 0
transform -1 0 2770 0 1 3390
box -6 -8 106 268
use AOI21X1  _2663_
timestamp 0
transform -1 0 2190 0 -1 3390
box -6 -8 106 268
use OAI21X1  _2664_
timestamp 0
transform 1 0 1030 0 -1 3390
box -6 -8 106 268
use NOR2X1  _2665_
timestamp 0
transform -1 0 1030 0 1 2870
box -6 -8 86 268
use NAND2X1  _2666_
timestamp 0
transform -1 0 550 0 -1 2870
box -6 -8 86 268
use NAND2X1  _2667_
timestamp 0
transform -1 0 770 0 1 2870
box -6 -8 86 268
use OAI22X1  _2668_
timestamp 0
transform 1 0 1210 0 1 2870
box -6 -8 126 268
use OAI21X1  _2669_
timestamp 0
transform -1 0 3050 0 1 3390
box -6 -8 106 268
use AOI21X1  _2670_
timestamp 0
transform -1 0 3170 0 1 2870
box -6 -8 106 268
use OAI21X1  _2671_
timestamp 0
transform 1 0 1250 0 -1 2870
box -6 -8 106 268
use INVX1  _2672_
timestamp 0
transform -1 0 790 0 -1 2870
box -6 -8 66 268
use NAND2X1  _2673_
timestamp 0
transform -1 0 770 0 1 2350
box -6 -8 86 268
use NAND3X1  _2674_
timestamp 0
transform 1 0 970 0 -1 2870
box -6 -8 106 268
use NAND3X1  _2675_
timestamp 0
transform 1 0 950 0 1 2350
box -6 -8 106 268
use OAI21X1  _2676_
timestamp 0
transform -1 0 1330 0 1 2350
box -6 -8 106 268
use AOI21X1  _2677_
timestamp 0
transform 1 0 6590 0 -1 2350
box -6 -8 106 268
use OAI22X1  _2678_
timestamp 0
transform -1 0 6610 0 -1 790
box -6 -8 126 268
use NAND3X1  _2679_
timestamp 0
transform 1 0 7150 0 1 1310
box -6 -8 106 268
use NAND3X1  _2680_
timestamp 0
transform -1 0 7010 0 -1 1310
box -6 -8 106 268
use NAND3X1  _2681_
timestamp 0
transform 1 0 7190 0 -1 1310
box -6 -8 106 268
use NOR3X1  _2682_
timestamp 0
transform -1 0 7070 0 1 790
box -6 -8 186 268
use OAI21X1  _2683_
timestamp 0
transform -1 0 2110 0 1 270
box -6 -8 106 268
use NAND2X1  _2684_
timestamp 0
transform -1 0 1910 0 -1 3390
box -6 -8 86 268
use NAND2X1  _2685_
timestamp 0
transform 1 0 1770 0 -1 2870
box -6 -8 86 268
use AOI22X1  _2686_
timestamp 0
transform 1 0 1770 0 1 2870
box -6 -8 126 268
use NAND2X1  _2687_
timestamp 0
transform 1 0 1510 0 1 2870
box -6 -8 86 268
use OR2X2  _2688_
timestamp 0
transform -1 0 1030 0 -1 790
box -6 -8 106 268
use NOR2X1  _2689_
timestamp 0
transform -1 0 990 0 1 270
box -6 -8 86 268
use AOI22X1  _2690_
timestamp 0
transform 1 0 7430 0 1 2350
box -6 -8 126 268
use NOR3X1  _2691_
timestamp 0
transform -1 0 7430 0 1 790
box -6 -8 186 268
use INVX1  _2692_
timestamp 0
transform -1 0 5250 0 -1 790
box -6 -8 66 268
use NAND3X1  _2693_
timestamp 0
transform -1 0 3250 0 -1 790
box -6 -8 106 268
use NOR2X1  _2694_
timestamp 0
transform -1 0 1550 0 -1 790
box -6 -8 86 268
use AOI21X1  _2695_
timestamp 0
transform -1 0 1830 0 -1 790
box -6 -8 106 268
use OAI21X1  _2696_
timestamp 0
transform -1 0 1550 0 1 270
box -6 -8 106 268
use OAI21X1  _2697_
timestamp 0
transform 1 0 2050 0 -1 270
box -6 -8 106 268
use INVX1  _2698_
timestamp 0
transform -1 0 730 0 1 270
box -6 -8 66 268
use AOI21X1  _2699_
timestamp 0
transform 1 0 6450 0 1 1830
box -6 -8 106 268
use OAI22X1  _2700_
timestamp 0
transform -1 0 7270 0 -1 790
box -6 -8 126 268
use NAND3X1  _2701_
timestamp 0
transform 1 0 7750 0 -1 1310
box -6 -8 106 268
use NAND3X1  _2702_
timestamp 0
transform 1 0 7450 0 -1 790
box -6 -8 106 268
use NAND3X1  _2703_
timestamp 0
transform 1 0 7610 0 1 790
box -6 -8 106 268
use NOR3X1  _2704_
timestamp 0
transform -1 0 6970 0 -1 790
box -6 -8 186 268
use OAI21X1  _2705_
timestamp 0
transform 1 0 1730 0 1 270
box -6 -8 106 268
use AOI21X1  _2706_
timestamp 0
transform 1 0 1170 0 1 270
box -6 -8 106 268
use NAND3X1  _2707_
timestamp 0
transform 1 0 2870 0 -1 790
box -6 -8 106 268
use AOI22X1  _2708_
timestamp 0
transform 1 0 2570 0 -1 790
box -6 -8 126 268
use INVX1  _2709_
timestamp 0
transform -1 0 1270 0 -1 790
box -6 -8 66 268
use OAI21X1  _2710_
timestamp 0
transform -1 0 1090 0 -1 270
box -6 -8 106 268
use OAI22X1  _2711_
timestamp 0
transform -1 0 1390 0 -1 270
box -6 -8 126 268
use NAND2X1  _2712_
timestamp 0
transform 1 0 3030 0 1 790
box -6 -8 86 268
use OAI21X1  _2713_
timestamp 0
transform -1 0 4510 0 1 790
box -6 -8 106 268
use NOR3X1  _2714_
timestamp 0
transform -1 0 5010 0 -1 790
box -6 -8 186 268
use OAI21X1  _2715_
timestamp 0
transform 1 0 3690 0 -1 790
box -6 -8 106 268
use INVX1  _2716_
timestamp 0
transform -1 0 4490 0 -1 5470
box -6 -8 66 268
use OAI21X1  _2717_
timestamp 0
transform -1 0 6090 0 1 3390
box -6 -8 106 268
use NOR3X1  _2718_
timestamp 0
transform -1 0 4410 0 -1 790
box -6 -8 186 268
use NAND3X1  _2719_
timestamp 0
transform 1 0 3850 0 1 790
box -6 -8 106 268
use NAND3X1  _2720_
timestamp 0
transform -1 0 4230 0 1 790
box -6 -8 106 268
use NAND2X1  _2721_
timestamp 0
transform -1 0 2370 0 -1 790
box -6 -8 86 268
use XOR2X1  _2722_
timestamp 0
transform 1 0 2430 0 1 790
box -6 -8 126 268
use OAI21X1  _2723_
timestamp 0
transform 1 0 2750 0 1 790
box -6 -8 106 268
use NOR2X1  _2724_
timestamp 0
transform -1 0 1030 0 1 790
box -6 -8 86 268
use AOI22X1  _2725_
timestamp 0
transform -1 0 5670 0 1 790
box -6 -8 126 268
use OAI21X1  _2726_
timestamp 0
transform -1 0 6830 0 1 1830
box -6 -8 106 268
use AOI22X1  _2727_
timestamp 0
transform 1 0 4010 0 1 2870
box -6 -8 126 268
use NAND3X1  _2728_
timestamp 0
transform 1 0 3730 0 1 2870
box -6 -8 106 268
use AOI21X1  _2729_
timestamp 0
transform -1 0 3770 0 1 2350
box -6 -8 106 268
use OAI21X1  _2730_
timestamp 0
transform 1 0 3290 0 1 790
box -6 -8 106 268
use AOI21X1  _2731_
timestamp 0
transform 1 0 2150 0 1 790
box -6 -8 106 268
use NAND3X1  _2732_
timestamp 0
transform -1 0 2110 0 -1 790
box -6 -8 106 268
use OAI21X1  _2733_
timestamp 0
transform 1 0 1570 0 1 790
box -6 -8 106 268
use OAI22X1  _2734_
timestamp 0
transform -1 0 1970 0 1 790
box -6 -8 126 268
use OAI21X1  _2735_
timestamp 0
transform -1 0 4110 0 -1 1830
box -6 -8 106 268
use AOI21X1  _2736_
timestamp 0
transform -1 0 4250 0 -1 2870
box -6 -8 106 268
use OAI21X1  _2737_
timestamp 0
transform -1 0 4330 0 1 1830
box -6 -8 106 268
use OR2X2  _2738_
timestamp 0
transform -1 0 4050 0 1 1830
box -6 -8 106 268
use AOI21X1  _2739_
timestamp 0
transform -1 0 3470 0 1 1830
box -6 -8 106 268
use OAI21X1  _2740_
timestamp 0
transform -1 0 3550 0 -1 1830
box -6 -8 106 268
use NOR3X1  _2741_
timestamp 0
transform -1 0 1390 0 1 790
box -6 -8 186 268
use XOR2X1  _2742_
timestamp 0
transform 1 0 1530 0 -1 1830
box -6 -8 126 268
use NAND2X1  _2743_
timestamp 0
transform 1 0 1470 0 1 1830
box -6 -8 86 268
use OAI21X1  _2744_
timestamp 0
transform 1 0 2010 0 1 1830
box -6 -8 106 268
use NAND2X1  _2745_
timestamp 0
transform 1 0 670 0 -1 790
box -6 -8 86 268
use OAI21X1  _2746_
timestamp 0
transform 1 0 3730 0 -1 1830
box -6 -8 106 268
use AOI21X1  _2747_
timestamp 0
transform 1 0 4850 0 1 2870
box -6 -8 106 268
use OAI21X1  _2748_
timestamp 0
transform 1 0 4510 0 1 1830
box -6 -8 106 268
use OR2X2  _2749_
timestamp 0
transform -1 0 3750 0 1 1830
box -6 -8 106 268
use AOI21X1  _2750_
timestamp 0
transform -1 0 3190 0 1 1830
box -6 -8 106 268
use OAI21X1  _2751_
timestamp 0
transform 1 0 2950 0 1 1310
box -6 -8 106 268
use NAND2X1  _2752_
timestamp 0
transform 1 0 1270 0 -1 1830
box -6 -8 86 268
use XOR2X1  _2753_
timestamp 0
transform 1 0 750 0 1 1310
box -6 -8 126 268
use OAI21X1  _2754_
timestamp 0
transform -1 0 770 0 1 790
box -6 -8 106 268
use NAND2X1  _2755_
timestamp 0
transform -1 0 3270 0 -1 1830
box -6 -8 86 268
use NAND2X1  _2756_
timestamp 0
transform -1 0 2710 0 -1 1830
box -6 -8 86 268
use AOI22X1  _2757_
timestamp 0
transform 1 0 2890 0 -1 1830
box -6 -8 126 268
use NOR2X1  _2758_
timestamp 0
transform 1 0 2370 0 -1 1830
box -6 -8 86 268
use OAI21X1  _2759_
timestamp 0
transform -1 0 4530 0 -1 2870
box -6 -8 106 268
use NOR2X1  _2760_
timestamp 0
transform 1 0 3890 0 -1 2870
box -6 -8 86 268
use AOI22X1  _2761_
timestamp 0
transform 1 0 4230 0 1 2350
box -6 -8 126 268
use NAND3X1  _2762_
timestamp 0
transform -1 0 4050 0 1 2350
box -6 -8 106 268
use NOR2X1  _2763_
timestamp 0
transform -1 0 2270 0 1 1310
box -6 -8 86 268
use NAND3X1  _2764_
timestamp 0
transform -1 0 2010 0 1 1310
box -6 -8 106 268
use NAND2X1  _2765_
timestamp 0
transform -1 0 1910 0 -1 1830
box -6 -8 86 268
use OAI21X1  _2766_
timestamp 0
transform -1 0 2190 0 -1 1830
box -6 -8 106 268
use NAND3X1  _2767_
timestamp 0
transform -1 0 1730 0 1 1310
box -6 -8 106 268
use NAND2X1  _2768_
timestamp 0
transform 1 0 2290 0 1 1830
box -6 -8 86 268
use AND2X2  _2769_
timestamp 0
transform 1 0 1730 0 1 1830
box -6 -8 106 268
use AOI22X1  _2770_
timestamp 0
transform 1 0 6090 0 1 2350
box -6 -8 126 268
use NAND3X1  _2771_
timestamp 0
transform 1 0 6630 0 1 2350
box -6 -8 106 268
use AOI21X1  _2772_
timestamp 0
transform 1 0 5070 0 1 2350
box -6 -8 106 268
use OAI21X1  _2773_
timestamp 0
transform 1 0 4270 0 -1 1310
box -6 -8 106 268
use INVX1  _2774_
timestamp 0
transform 1 0 2430 0 -1 1310
box -6 -8 66 268
use NAND3X1  _2775_
timestamp 0
transform 1 0 2670 0 -1 1310
box -6 -8 106 268
use XOR2X1  _2776_
timestamp 0
transform 1 0 3490 0 -1 1310
box -6 -8 126 268
use NAND2X1  _2777_
timestamp 0
transform -1 0 3030 0 -1 1310
box -6 -8 86 268
use OAI21X1  _2778_
timestamp 0
transform -1 0 3310 0 -1 1310
box -6 -8 106 268
use INVX1  _2779_
timestamp 0
transform -1 0 7310 0 -1 270
box -6 -8 66 268
use NAND2X1  _2780_
timestamp 0
transform -1 0 7570 0 -1 270
box -6 -8 86 268
use OAI21X1  _2781_
timestamp 0
transform 1 0 7990 0 -1 790
box -6 -8 106 268
use OAI21X1  _2782_
timestamp 0
transform 1 0 7890 0 1 270
box -6 -8 106 268
use INVX1  _2783_
timestamp 0
transform 1 0 9810 0 1 7550
box -6 -8 66 268
use INVX2  _2784_
timestamp 0
transform 1 0 10950 0 1 10150
box -6 -8 66 268
use NAND2X1  _2785_
timestamp 0
transform 1 0 10330 0 1 7550
box -6 -8 86 268
use OAI21X1  _2786_
timestamp 0
transform 1 0 10050 0 1 7550
box -6 -8 106 268
use NAND2X1  _2787_
timestamp 0
transform 1 0 8510 0 -1 7030
box -6 -8 86 268
use OAI21X1  _2788_
timestamp 0
transform 1 0 8770 0 -1 7030
box -6 -8 106 268
use NAND2X1  _2789_
timestamp 0
transform 1 0 8290 0 1 7030
box -6 -8 86 268
use OAI21X1  _2790_
timestamp 0
transform -1 0 8110 0 1 7030
box -6 -8 106 268
use INVX1  _2791_
timestamp 0
transform 1 0 6290 0 -1 7550
box -6 -8 66 268
use OAI22X1  _2792_
timestamp 0
transform 1 0 9910 0 -1 7550
box -6 -8 126 268
use INVX1  _2793_
timestamp 0
transform 1 0 10110 0 1 7030
box -6 -8 66 268
use NAND2X1  _2794_
timestamp 0
transform -1 0 10430 0 1 7030
box -6 -8 86 268
use OAI21X1  _2795_
timestamp 0
transform 1 0 8550 0 1 7030
box -6 -8 106 268
use OAI21X1  _2796_
timestamp 0
transform 1 0 8530 0 -1 9630
box -6 -8 106 268
use NAND2X1  _2797_
timestamp 0
transform 1 0 10950 0 -1 8070
box -6 -8 86 268
use OR2X2  _2798_
timestamp 0
transform -1 0 10150 0 1 9110
box -6 -8 106 268
use OAI21X1  _2799_
timestamp 0
transform -1 0 8530 0 1 9110
box -6 -8 106 268
use INVX1  _2800_
timestamp 0
transform -1 0 7890 0 -1 9110
box -6 -8 66 268
use NOR2X1  _2801_
timestamp 0
transform 1 0 9790 0 -1 8590
box -6 -8 86 268
use NAND2X1  _2802_
timestamp 0
transform -1 0 10170 0 1 8590
box -6 -8 86 268
use OAI22X1  _2803_
timestamp 0
transform 1 0 8550 0 -1 9110
box -6 -8 126 268
use OAI21X1  _2804_
timestamp 0
transform -1 0 8530 0 -1 8590
box -6 -8 106 268
use NOR2X1  _2805_
timestamp 0
transform -1 0 10250 0 1 10150
box -6 -8 86 268
use NAND2X1  _2806_
timestamp 0
transform 1 0 9870 0 -1 9110
box -6 -8 86 268
use OAI21X1  _2807_
timestamp 0
transform -1 0 8570 0 1 8590
box -6 -8 106 268
use INVX1  _2808_
timestamp 0
transform -1 0 6770 0 1 8070
box -6 -8 66 268
use OAI22X1  _2809_
timestamp 0
transform 1 0 8250 0 1 8070
box -6 -8 126 268
use INVX1  _2810_
timestamp 0
transform -1 0 7710 0 -1 8070
box -6 -8 66 268
use INVX1  _2811_
timestamp 0
transform 1 0 10170 0 -1 9630
box -6 -8 66 268
use NAND2X1  _2812_
timestamp 0
transform 1 0 9790 0 1 9110
box -6 -8 86 268
use OAI22X1  _2813_
timestamp 0
transform 1 0 8370 0 -1 8070
box -6 -8 126 268
use OAI21X1  _2814_
timestamp 0
transform -1 0 8330 0 -1 7030
box -6 -8 106 268
use OAI21X1  _2815_
timestamp 0
transform -1 0 8410 0 -1 7550
box -6 -8 106 268
use OAI21X1  _2816_
timestamp 0
transform 1 0 9590 0 1 8070
box -6 -8 106 268
use NOR2X1  _2817_
timestamp 0
transform -1 0 10510 0 1 10150
box -6 -8 86 268
use NAND2X1  _2818_
timestamp 0
transform 1 0 11270 0 -1 11190
box -6 -8 86 268
use NOR2X1  _2819_
timestamp 0
transform 1 0 10250 0 1 11190
box -6 -8 86 268
use INVX1  _2820_
timestamp 0
transform -1 0 10070 0 1 11190
box -6 -8 66 268
use OAI21X1  _2821_
timestamp 0
transform -1 0 9970 0 1 8070
box -6 -8 106 268
use INVX1  _2822_
timestamp 0
transform -1 0 7650 0 -1 7550
box -6 -8 66 268
use NAND3X1  _2823_
timestamp 0
transform -1 0 9690 0 -1 9630
box -6 -8 106 268
use NOR2X1  _2824_
timestamp 0
transform -1 0 9410 0 -1 9630
box -6 -8 86 268
use NOR2X1  _2825_
timestamp 0
transform 1 0 8810 0 -1 9630
box -6 -8 86 268
use AOI21X1  _2826_
timestamp 0
transform 1 0 8870 0 -1 7550
box -6 -8 106 268
use NOR2X1  _2827_
timestamp 0
transform 1 0 9270 0 1 9630
box -6 -8 86 268
use AND2X2  _2828_
timestamp 0
transform 1 0 10390 0 -1 10150
box -6 -8 106 268
use INVX1  _2829_
timestamp 0
transform -1 0 9370 0 -1 10670
box -6 -8 66 268
use NOR2X1  _2830_
timestamp 0
transform 1 0 9950 0 -1 11190
box -6 -8 86 268
use NOR2X1  _2831_
timestamp 0
transform 1 0 9130 0 1 10150
box -6 -8 86 268
use OAI21X1  _2832_
timestamp 0
transform -1 0 9130 0 -1 10670
box -6 -8 106 268
use INVX1  _2833_
timestamp 0
transform -1 0 8850 0 -1 10670
box -6 -8 66 268
use INVX1  _2834_
timestamp 0
transform -1 0 8430 0 1 10670
box -6 -8 66 268
use NOR2X1  _2835_
timestamp 0
transform -1 0 9470 0 1 10150
box -6 -8 86 268
use AOI21X1  _2836_
timestamp 0
transform -1 0 8190 0 1 10670
box -6 -8 106 268
use AOI22X1  _2837_
timestamp 0
transform 1 0 8190 0 -1 10670
box -6 -8 126 268
use NAND2X1  _2838_
timestamp 0
transform 1 0 9430 0 1 10670
box -6 -8 86 268
use NOR2X1  _2839_
timestamp 0
transform 1 0 9690 0 -1 11190
box -6 -8 86 268
use OAI21X1  _2840_
timestamp 0
transform -1 0 9510 0 -1 11190
box -6 -8 106 268
use AOI22X1  _2841_
timestamp 0
transform 1 0 8350 0 -1 11190
box -6 -8 126 268
use NAND2X1  _2842_
timestamp 0
transform 1 0 11650 0 -1 10670
box -6 -8 86 268
use OAI21X1  _2843_
timestamp 0
transform -1 0 11230 0 -1 10670
box -6 -8 106 268
use NAND2X1  _2844_
timestamp 0
transform 1 0 10870 0 -1 10670
box -6 -8 86 268
use NAND2X1  _2845_
timestamp 0
transform 1 0 10610 0 -1 10670
box -6 -8 86 268
use OAI21X1  _2846_
timestamp 0
transform -1 0 10330 0 1 10670
box -6 -8 106 268
use NAND2X1  _2847_
timestamp 0
transform 1 0 10450 0 -1 11190
box -6 -8 86 268
use NAND2X1  _2848_
timestamp 0
transform -1 0 9790 0 -1 11710
box -6 -8 86 268
use NOR2X1  _2849_
timestamp 0
transform 1 0 11030 0 1 11710
box -6 -8 86 268
use INVX1  _2850_
timestamp 0
transform 1 0 11190 0 -1 12230
box -6 -8 66 268
use INVX1  _2851_
timestamp 0
transform 1 0 11430 0 1 10150
box -6 -8 66 268
use NOR2X1  _2852_
timestamp 0
transform 1 0 12130 0 1 11190
box -6 -8 86 268
use NAND2X1  _2853_
timestamp 0
transform 1 0 12190 0 -1 10670
box -6 -8 86 268
use NAND3X1  _2854_
timestamp 0
transform 1 0 11870 0 1 10670
box -6 -8 106 268
use OAI21X1  _2855_
timestamp 0
transform 1 0 12150 0 1 10670
box -6 -8 106 268
use INVX1  _2856_
timestamp 0
transform -1 0 9250 0 1 10670
box -6 -8 66 268
use OAI21X1  _2857_
timestamp 0
transform 1 0 9690 0 1 10670
box -6 -8 106 268
use NOR2X1  _2858_
timestamp 0
transform -1 0 10050 0 1 10670
box -6 -8 86 268
use AOI21X1  _2859_
timestamp 0
transform 1 0 10930 0 -1 10150
box -6 -8 106 268
use AND2X2  _2860_
timestamp 0
transform 1 0 7810 0 1 10670
box -6 -8 106 268
use AOI22X1  _2861_
timestamp 0
transform 1 0 8490 0 -1 10670
box -6 -8 126 268
use INVX1  _2862_
timestamp 0
transform -1 0 7910 0 -1 11190
box -6 -8 66 268
use OAI21X1  _2863_
timestamp 0
transform 1 0 7570 0 -1 11190
box -6 -8 106 268
use OAI21X1  _2864_
timestamp 0
transform 1 0 9810 0 1 8590
box -6 -8 106 268
use OAI22X1  _2865_
timestamp 0
transform 1 0 8970 0 -1 8590
box -6 -8 126 268
use AOI21X1  _2866_
timestamp 0
transform -1 0 7150 0 1 10670
box -6 -8 106 268
use AND2X2  _2867_
timestamp 0
transform -1 0 8990 0 1 10670
box -6 -8 106 268
use OAI21X1  _2868_
timestamp 0
transform -1 0 8710 0 1 10670
box -6 -8 106 268
use OAI21X1  _2869_
timestamp 0
transform -1 0 9150 0 -1 10150
box -6 -8 106 268
use NAND2X1  _2870_
timestamp 0
transform 1 0 8730 0 1 9110
box -6 -8 86 268
use OAI22X1  _2871_
timestamp 0
transform 1 0 8670 0 -1 8070
box -6 -8 126 268
use OAI21X1  _2872_
timestamp 0
transform 1 0 5610 0 -1 5470
box -6 -8 106 268
use INVX1  _2873_
timestamp 0
transform -1 0 5670 0 1 7030
box -6 -8 66 268
use NAND2X1  _2874_
timestamp 0
transform 1 0 5550 0 -1 7550
box -6 -8 86 268
use NAND3X1  _2875_
timestamp 0
transform -1 0 5990 0 1 8070
box -6 -8 106 268
use OAI22X1  _2876_
timestamp 0
transform 1 0 5590 0 1 7550
box -6 -8 126 268
use INVX1  _2877_
timestamp 0
transform 1 0 6170 0 1 7550
box -6 -8 66 268
use OAI21X1  _2878_
timestamp 0
transform -1 0 5990 0 1 7550
box -6 -8 106 268
use OAI21X1  _2879_
timestamp 0
transform -1 0 9130 0 1 8070
box -6 -8 106 268
use NOR2X1  _2880_
timestamp 0
transform -1 0 12110 0 -1 10150
box -6 -8 86 268
use AOI22X1  _2881_
timestamp 0
transform 1 0 11730 0 -1 10150
box -6 -8 126 268
use OAI21X1  _2882_
timestamp 0
transform -1 0 9410 0 1 8070
box -6 -8 106 268
use OAI21X1  _2883_
timestamp 0
transform 1 0 9130 0 -1 11190
box -6 -8 106 268
use OAI21X1  _2884_
timestamp 0
transform -1 0 9530 0 1 11190
box -6 -8 106 268
use OR2X2  _2885_
timestamp 0
transform -1 0 10730 0 1 9630
box -6 -8 106 268
use OAI22X1  _2886_
timestamp 0
transform 1 0 10590 0 1 8590
box -6 -8 126 268
use NAND2X1  _2887_
timestamp 0
transform -1 0 9070 0 1 9110
box -6 -8 86 268
use OAI21X1  _2888_
timestamp 0
transform -1 0 9370 0 1 8590
box -6 -8 106 268
use OAI21X1  _2889_
timestamp 0
transform 1 0 9570 0 -1 10150
box -6 -8 106 268
use NOR2X1  _2890_
timestamp 0
transform -1 0 9990 0 1 10150
box -6 -8 86 268
use OAI21X1  _2891_
timestamp 0
transform -1 0 9950 0 -1 10150
box -6 -8 106 268
use OAI21X1  _2892_
timestamp 0
transform 1 0 9250 0 1 9110
box -6 -8 106 268
use INVX1  _2893_
timestamp 0
transform -1 0 9450 0 1 7030
box -6 -8 66 268
use NAND2X1  _2894_
timestamp 0
transform -1 0 11290 0 -1 10150
box -6 -8 86 268
use NOR2X1  _2895_
timestamp 0
transform 1 0 10910 0 1 9630
box -6 -8 86 268
use OAI21X1  _2896_
timestamp 0
transform -1 0 11270 0 1 8590
box -6 -8 106 268
use OAI21X1  _2897_
timestamp 0
transform -1 0 10990 0 1 8590
box -6 -8 106 268
use OAI21X1  _2898_
timestamp 0
transform 1 0 9530 0 1 7550
box -6 -8 106 268
use NAND2X1  _2899_
timestamp 0
transform -1 0 9890 0 -1 10670
box -6 -8 86 268
use OAI21X1  _2900_
timestamp 0
transform 1 0 10530 0 1 11190
box -6 -8 106 268
use OR2X2  _2901_
timestamp 0
transform -1 0 10610 0 1 10670
box -6 -8 106 268
use OAI21X1  _2902_
timestamp 0
transform 1 0 10710 0 -1 11190
box -6 -8 106 268
use AOI21X1  _2903_
timestamp 0
transform -1 0 10910 0 1 11190
box -6 -8 106 268
use OAI21X1  _2904_
timestamp 0
transform -1 0 10070 0 -1 11710
box -6 -8 106 268
use INVX1  _2905_
timestamp 0
transform -1 0 9530 0 -1 11710
box -6 -8 66 268
use OAI21X1  _2906_
timestamp 0
transform -1 0 8730 0 -1 11710
box -6 -8 106 268
use OAI21X1  _2907_
timestamp 0
transform -1 0 9290 0 -1 11710
box -6 -8 106 268
use OAI21X1  _2908_
timestamp 0
transform -1 0 10630 0 -1 11710
box -6 -8 106 268
use NAND3X1  _2909_
timestamp 0
transform 1 0 11910 0 -1 10670
box -6 -8 106 268
use NAND3X1  _2910_
timestamp 0
transform 1 0 10990 0 -1 11190
box -6 -8 106 268
use OAI21X1  _2911_
timestamp 0
transform 1 0 11850 0 -1 11710
box -6 -8 106 268
use NOR2X1  _2912_
timestamp 0
transform 1 0 12130 0 1 11710
box -6 -8 86 268
use AOI22X1  _2913_
timestamp 0
transform 1 0 10730 0 1 11710
box -6 -8 126 268
use INVX1  _2914_
timestamp 0
transform -1 0 7970 0 -1 12230
box -6 -8 66 268
use OAI21X1  _2915_
timestamp 0
transform 1 0 11050 0 -1 11710
box -6 -8 106 268
use OAI21X1  _2916_
timestamp 0
transform 1 0 11290 0 1 11710
box -6 -8 106 268
use OAI21X1  _2917_
timestamp 0
transform 1 0 10790 0 1 10670
box -6 -8 106 268
use NOR2X1  _2918_
timestamp 0
transform -1 0 11010 0 -1 12230
box -6 -8 86 268
use AOI21X1  _2919_
timestamp 0
transform 1 0 8630 0 -1 12230
box -6 -8 106 268
use INVX1  _2920_
timestamp 0
transform 1 0 11330 0 -1 11710
box -6 -8 66 268
use AOI21X1  _2921_
timestamp 0
transform 1 0 11850 0 1 11710
box -6 -8 106 268
use OAI21X1  _2922_
timestamp 0
transform -1 0 12050 0 -1 12230
box -6 -8 106 268
use NOR2X1  _2923_
timestamp 0
transform 1 0 11430 0 -1 12230
box -6 -8 86 268
use AOI21X1  _2924_
timestamp 0
transform 1 0 10350 0 -1 12230
box -6 -8 106 268
use INVX1  _2925_
timestamp 0
transform 1 0 10110 0 -1 12230
box -6 -8 66 268
use OAI21X1  _2926_
timestamp 0
transform 1 0 10250 0 -1 11710
box -6 -8 106 268
use NAND2X1  _2927_
timestamp 0
transform -1 0 10150 0 -1 10670
box -6 -8 86 268
use OAI21X1  _2928_
timestamp 0
transform -1 0 10430 0 -1 10670
box -6 -8 106 268
use NOR2X1  _2929_
timestamp 0
transform -1 0 10550 0 1 11710
box -6 -8 86 268
use NOR2X1  _2930_
timestamp 0
transform -1 0 11410 0 1 10670
box -6 -8 86 268
use NAND3X1  _2931_
timestamp 0
transform -1 0 11690 0 1 10670
box -6 -8 106 268
use NAND3X1  _2932_
timestamp 0
transform 1 0 11570 0 -1 11710
box -6 -8 106 268
use OAI21X1  _2933_
timestamp 0
transform 1 0 11530 0 -1 11190
box -6 -8 106 268
use NAND3X1  _2934_
timestamp 0
transform 1 0 11610 0 1 11190
box -6 -8 106 268
use NOR2X1  _2935_
timestamp 0
transform 1 0 11690 0 -1 12230
box -6 -8 86 268
use AOI22X1  _2936_
timestamp 0
transform 1 0 10630 0 -1 12230
box -6 -8 126 268
use AND2X2  _2937_
timestamp 0
transform -1 0 3710 0 -1 2870
box -6 -8 106 268
use OAI21X1  _2938_
timestamp 0
transform -1 0 7930 0 -1 5990
box -6 -8 106 268
use NOR2X1  _2939_
timestamp 0
transform 1 0 6610 0 1 9630
box -6 -8 86 268
use INVX2  _2940_
timestamp 0
transform -1 0 6430 0 1 9630
box -6 -8 66 268
use OAI21X1  _2941_
timestamp 0
transform -1 0 6390 0 1 8590
box -6 -8 106 268
use OAI21X1  _2942_
timestamp 0
transform 1 0 5210 0 -1 8590
box -6 -8 106 268
use OAI21X1  _2943_
timestamp 0
transform -1 0 7190 0 1 8590
box -6 -8 106 268
use OAI21X1  _2944_
timestamp 0
transform 1 0 5510 0 -1 8590
box -6 -8 106 268
use OAI21X1  _2945_
timestamp 0
transform -1 0 6970 0 1 9110
box -6 -8 106 268
use OAI21X1  _2946_
timestamp 0
transform 1 0 6490 0 -1 9110
box -6 -8 106 268
use OAI21X1  _2947_
timestamp 0
transform 1 0 7970 0 -1 10150
box -6 -8 106 268
use OAI21X1  _2948_
timestamp 0
transform 1 0 7710 0 1 9630
box -6 -8 106 268
use OAI21X1  _2949_
timestamp 0
transform 1 0 5810 0 1 9110
box -6 -8 106 268
use OAI21X1  _2950_
timestamp 0
transform -1 0 6230 0 -1 9630
box -6 -8 106 268
use OAI21X1  _2951_
timestamp 0
transform 1 0 6910 0 -1 10150
box -6 -8 106 268
use OAI21X1  _2952_
timestamp 0
transform 1 0 6630 0 -1 10150
box -6 -8 106 268
use OAI21X1  _2953_
timestamp 0
transform 1 0 5790 0 -1 8590
box -6 -8 106 268
use OAI21X1  _2954_
timestamp 0
transform -1 0 6170 0 -1 8590
box -6 -8 106 268
use OAI21X1  _2955_
timestamp 0
transform 1 0 7170 0 -1 9630
box -6 -8 106 268
use OAI21X1  _2956_
timestamp 0
transform 1 0 6650 0 -1 9630
box -6 -8 106 268
use OAI21X1  _2957_
timestamp 0
transform -1 0 8350 0 -1 10150
box -6 -8 106 268
use OAI21X1  _2958_
timestamp 0
transform 1 0 6650 0 -1 5470
box -6 -8 106 268
use INVX1  _2959_
timestamp 0
transform 1 0 6410 0 -1 7030
box -6 -8 66 268
use OAI21X1  _2960_
timestamp 0
transform -1 0 7350 0 1 7030
box -6 -8 106 268
use NOR2X1  _2961_
timestamp 0
transform 1 0 6650 0 -1 7030
box -6 -8 86 268
use INVX1  _2962_
timestamp 0
transform -1 0 6470 0 1 7550
box -6 -8 66 268
use NOR2X1  _2963_
timestamp 0
transform -1 0 6790 0 -1 8070
box -6 -8 86 268
use INVX1  _2964_
timestamp 0
transform 1 0 4790 0 -1 7550
box -6 -8 66 268
use OAI21X1  _2965_
timestamp 0
transform 1 0 5850 0 1 7030
box -6 -8 106 268
use OAI21X1  _2966_
timestamp 0
transform -1 0 6830 0 -1 5990
box -6 -8 106 268
use NAND2X1  _2967_
timestamp 0
transform -1 0 5230 0 -1 6510
box -6 -8 86 268
use OAI21X1  _2968_
timestamp 0
transform -1 0 5510 0 -1 6510
box -6 -8 106 268
use AOI21X1  _2969_
timestamp 0
transform 1 0 4510 0 -1 7550
box -6 -8 106 268
use NAND2X1  _2970_
timestamp 0
transform 1 0 4870 0 -1 7030
box -6 -8 86 268
use OAI21X1  _2971_
timestamp 0
transform 1 0 4750 0 1 7030
box -6 -8 106 268
use NOR2X1  _2972_
timestamp 0
transform -1 0 6250 0 1 8070
box -6 -8 86 268
use NAND2X1  _2973_
timestamp 0
transform -1 0 6530 0 1 8070
box -6 -8 86 268
use OAI21X1  _2974_
timestamp 0
transform -1 0 6530 0 -1 8070
box -6 -8 106 268
use NAND2X1  _2975_
timestamp 0
transform 1 0 5910 0 -1 8070
box -6 -8 86 268
use NAND2X1  _2976_
timestamp 0
transform -1 0 4890 0 1 8070
box -6 -8 86 268
use OAI21X1  _2977_
timestamp 0
transform -1 0 5170 0 1 8070
box -6 -8 106 268
use MUX2X1  _2978_
timestamp 0
transform 1 0 5350 0 1 8070
box -6 -8 126 268
use OAI21X1  _2979_
timestamp 0
transform 1 0 5630 0 -1 8070
box -6 -8 106 268
use NAND2X1  _2980_
timestamp 0
transform -1 0 7570 0 -1 7030
box -6 -8 86 268
use AOI21X1  _2981_
timestamp 0
transform -1 0 6550 0 1 6510
box -6 -8 106 268
use OAI22X1  _2982_
timestamp 0
transform -1 0 6850 0 1 6510
box -6 -8 126 268
use INVX1  _2983_
timestamp 0
transform 1 0 7270 0 1 5990
box -6 -8 66 268
use OAI21X1  _2984_
timestamp 0
transform 1 0 6670 0 -1 6510
box -6 -8 106 268
use OAI21X1  _2985_
timestamp 0
transform -1 0 7090 0 1 5990
box -6 -8 106 268
use AOI21X1  _2986_
timestamp 0
transform 1 0 6710 0 1 5990
box -6 -8 106 268
use NAND2X1  _2987_
timestamp 0
transform 1 0 6150 0 1 5990
box -6 -8 86 268
use OAI21X1  _2988_
timestamp 0
transform -1 0 6530 0 1 5990
box -6 -8 106 268
use NOR2X1  _2989_
timestamp 0
transform -1 0 8070 0 1 9630
box -6 -8 86 268
use OAI21X1  _2990_
timestamp 0
transform 1 0 7130 0 1 9630
box -6 -8 106 268
use OAI21X1  _2991_
timestamp 0
transform -1 0 7070 0 1 7030
box -6 -8 106 268
use OAI21X1  _2992_
timestamp 0
transform -1 0 5370 0 -1 7550
box -6 -8 106 268
use OAI21X1  _2993_
timestamp 0
transform -1 0 6230 0 1 7030
box -6 -8 106 268
use INVX1  _2994_
timestamp 0
transform 1 0 5610 0 -1 7030
box -6 -8 66 268
use OAI21X1  _2995_
timestamp 0
transform 1 0 6690 0 1 7030
box -6 -8 106 268
use OAI21X1  _2996_
timestamp 0
transform 1 0 6410 0 1 7030
box -6 -8 106 268
use NAND2X1  _2997_
timestamp 0
transform 1 0 6130 0 -1 7030
box -6 -8 86 268
use OAI21X1  _2998_
timestamp 0
transform -1 0 5950 0 -1 7030
box -6 -8 106 268
use OAI22X1  _2999_
timestamp 0
transform 1 0 6530 0 -1 7550
box -6 -8 126 268
use MUX2X1  _3000_
timestamp 0
transform -1 0 5970 0 1 5990
box -6 -8 126 268
use NAND2X1  _3001_
timestamp 0
transform 1 0 5090 0 1 6510
box -6 -8 86 268
use OAI21X1  _3002_
timestamp 0
transform -1 0 5670 0 1 5990
box -6 -8 106 268
use MUX2X1  _3003_
timestamp 0
transform -1 0 6070 0 -1 5990
box -6 -8 126 268
use NAND2X1  _3004_
timestamp 0
transform -1 0 5430 0 1 6510
box -6 -8 86 268
use OAI21X1  _3005_
timestamp 0
transform -1 0 5710 0 1 6510
box -6 -8 106 268
use NOR2X1  _3006_
timestamp 0
transform -1 0 7590 0 1 8070
box -6 -8 86 268
use NAND3X1  _3007_
timestamp 0
transform 1 0 6950 0 1 8070
box -6 -8 106 268
use NOR2X1  _3008_
timestamp 0
transform 1 0 8750 0 1 8590
box -6 -8 86 268
use NAND2X1  _3009_
timestamp 0
transform 1 0 8210 0 1 8590
box -6 -8 86 268
use OAI21X1  _3010_
timestamp 0
transform 1 0 7230 0 1 8070
box -6 -8 106 268
use AOI21X1  _3011_
timestamp 0
transform -1 0 7410 0 -1 7550
box -6 -8 106 268
use AND2X2  _3012_
timestamp 0
transform -1 0 7290 0 1 7550
box -6 -8 106 268
use AOI21X1  _3013_
timestamp 0
transform -1 0 8030 0 1 8590
box -6 -8 106 268
use NAND2X1  _3014_
timestamp 0
transform 1 0 7150 0 -1 8590
box -6 -8 86 268
use OAI21X1  _3015_
timestamp 0
transform -1 0 7510 0 -1 8590
box -6 -8 106 268
use NAND2X1  _3016_
timestamp 0
transform -1 0 6250 0 -1 8070
box -6 -8 86 268
use OAI21X1  _3017_
timestamp 0
transform -1 0 7090 0 -1 8070
box -6 -8 106 268
use NAND2X1  _3018_
timestamp 0
transform -1 0 6730 0 1 7550
box -6 -8 86 268
use OAI21X1  _3019_
timestamp 0
transform -1 0 7010 0 1 7550
box -6 -8 106 268
use INVX1  _3020_
timestamp 0
transform 1 0 5570 0 1 4430
box -6 -8 66 268
use NAND2X1  _3021_
timestamp 0
transform 1 0 6010 0 -1 4430
box -6 -8 86 268
use OAI21X1  _3022_
timestamp 0
transform 1 0 5810 0 1 4430
box -6 -8 106 268
use NOR2X1  _3023_
timestamp 0
transform -1 0 6950 0 1 9630
box -6 -8 86 268
use OAI21X1  _3024_
timestamp 0
transform -1 0 6890 0 -1 4430
box -6 -8 106 268
use NOR2X1  _3025_
timestamp 0
transform 1 0 6090 0 1 4430
box -6 -8 86 268
use INVX1  _3026_
timestamp 0
transform 1 0 5510 0 1 5470
box -6 -8 66 268
use OAI21X1  _3027_
timestamp 0
transform -1 0 5690 0 -1 9630
box -6 -8 106 268
use INVX1  _3028_
timestamp 0
transform 1 0 6090 0 1 11190
box -6 -8 66 268
use NAND2X1  _3029_
timestamp 0
transform 1 0 6850 0 1 11190
box -6 -8 86 268
use OAI21X1  _3030_
timestamp 0
transform 1 0 4990 0 1 3910
box -6 -8 106 268
use OAI21X1  _3031_
timestamp 0
transform 1 0 4530 0 1 8070
box -6 -8 106 268
use NAND2X1  _3032_
timestamp 0
transform -1 0 5390 0 -1 9110
box -6 -8 86 268
use OAI21X1  _3033_
timestamp 0
transform 1 0 5570 0 -1 9110
box -6 -8 106 268
use NAND3X1  _3034_
timestamp 0
transform -1 0 3590 0 1 7550
box -6 -8 106 268
use NAND2X1  _3035_
timestamp 0
transform -1 0 4130 0 1 7550
box -6 -8 86 268
use OAI21X1  _3036_
timestamp 0
transform -1 0 3650 0 -1 8070
box -6 -8 106 268
use INVX1  _3037_
timestamp 0
transform -1 0 3490 0 1 8070
box -6 -8 66 268
use NOR2X1  _3038_
timestamp 0
transform 1 0 3670 0 1 8070
box -6 -8 86 268
use OAI21X1  _3039_
timestamp 0
transform -1 0 3250 0 1 8070
box -6 -8 106 268
use INVX1  _3040_
timestamp 0
transform 1 0 3050 0 -1 8070
box -6 -8 66 268
use NOR2X1  _3041_
timestamp 0
transform 1 0 3290 0 -1 8070
box -6 -8 86 268
use OAI21X1  _3042_
timestamp 0
transform -1 0 3930 0 -1 8070
box -6 -8 106 268
use OAI21X1  _3043_
timestamp 0
transform -1 0 4030 0 -1 8590
box -6 -8 106 268
use INVX1  _3044_
timestamp 0
transform -1 0 3750 0 -1 8590
box -6 -8 66 268
use NAND2X1  _3045_
timestamp 0
transform 1 0 4510 0 1 8590
box -6 -8 86 268
use OAI21X1  _3046_
timestamp 0
transform 1 0 4230 0 1 8590
box -6 -8 106 268
use XNOR2X1  _3047_
timestamp 0
transform -1 0 3310 0 1 7550
box -6 -8 126 268
use INVX1  _3048_
timestamp 0
transform 1 0 3230 0 -1 7550
box -6 -8 66 268
use NAND2X1  _3049_
timestamp 0
transform -1 0 2990 0 1 7550
box -6 -8 86 268
use NOR2X1  _3050_
timestamp 0
transform 1 0 2970 0 -1 7550
box -6 -8 86 268
use NOR2X1  _3051_
timestamp 0
transform 1 0 2710 0 -1 7550
box -6 -8 86 268
use AOI22X1  _3052_
timestamp 0
transform 1 0 2610 0 1 7550
box -6 -8 126 268
use NAND2X1  _3053_
timestamp 0
transform 1 0 3370 0 1 9630
box -6 -8 86 268
use OAI21X1  _3054_
timestamp 0
transform -1 0 3730 0 1 9630
box -6 -8 106 268
use INVX1  _3055_
timestamp 0
transform 1 0 3470 0 -1 7550
box -6 -8 66 268
use OAI21X1  _3056_
timestamp 0
transform -1 0 3810 0 -1 7550
box -6 -8 106 268
use XNOR2X1  _3057_
timestamp 0
transform 1 0 3930 0 1 8070
box -6 -8 126 268
use AND2X2  _3058_
timestamp 0
transform 1 0 4110 0 -1 8070
box -6 -8 106 268
use OAI21X1  _3059_
timestamp 0
transform 1 0 4390 0 -1 8070
box -6 -8 106 268
use OAI22X1  _3060_
timestamp 0
transform 1 0 4230 0 1 8070
box -6 -8 126 268
use NAND2X1  _3061_
timestamp 0
transform 1 0 3710 0 1 11710
box -6 -8 86 268
use OAI21X1  _3062_
timestamp 0
transform -1 0 4050 0 -1 11710
box -6 -8 106 268
use OAI21X1  _3063_
timestamp 0
transform -1 0 5270 0 1 3390
box -6 -8 106 268
use OAI21X1  _3064_
timestamp 0
transform 1 0 5050 0 -1 5470
box -6 -8 106 268
use NAND2X1  _3065_
timestamp 0
transform -1 0 4850 0 1 8590
box -6 -8 86 268
use OAI21X1  _3066_
timestamp 0
transform 1 0 4690 0 -1 8590
box -6 -8 106 268
use NAND3X1  _3067_
timestamp 0
transform -1 0 3870 0 1 7550
box -6 -8 106 268
use OAI21X1  _3068_
timestamp 0
transform -1 0 3610 0 -1 7030
box -6 -8 106 268
use INVX1  _3069_
timestamp 0
transform 1 0 3730 0 1 6510
box -6 -8 66 268
use NAND2X1  _3070_
timestamp 0
transform -1 0 4690 0 -1 6510
box -6 -8 86 268
use NOR2X1  _3071_
timestamp 0
transform 1 0 4350 0 -1 6510
box -6 -8 86 268
use NOR2X1  _3072_
timestamp 0
transform -1 0 4350 0 1 6510
box -6 -8 86 268
use AOI22X1  _3073_
timestamp 0
transform -1 0 4650 0 1 6510
box -6 -8 126 268
use NAND2X1  _3074_
timestamp 0
transform 1 0 5830 0 1 11190
box -6 -8 86 268
use OAI21X1  _3075_
timestamp 0
transform 1 0 5550 0 1 11190
box -6 -8 106 268
use XNOR2X1  _3076_
timestamp 0
transform 1 0 3810 0 -1 7030
box -6 -8 126 268
use AOI21X1  _3077_
timestamp 0
transform 1 0 4110 0 -1 7030
box -6 -8 106 268
use OAI21X1  _3078_
timestamp 0
transform 1 0 4170 0 1 7030
box -6 -8 106 268
use OAI21X1  _3079_
timestamp 0
transform -1 0 4330 0 -1 7550
box -6 -8 106 268
use INVX1  _3080_
timestamp 0
transform 1 0 6390 0 -1 10150
box -6 -8 66 268
use NAND2X1  _3081_
timestamp 0
transform -1 0 7110 0 1 11710
box -6 -8 86 268
use OAI21X1  _3082_
timestamp 0
transform 1 0 6750 0 -1 12230
box -6 -8 106 268
use NAND2X1  _3083_
timestamp 0
transform -1 0 3990 0 1 7030
box -6 -8 86 268
use OAI21X1  _3084_
timestamp 0
transform 1 0 3630 0 1 7030
box -6 -8 106 268
use NOR2X1  _3085_
timestamp 0
transform 1 0 3250 0 -1 7030
box -6 -8 86 268
use XOR2X1  _3086_
timestamp 0
transform -1 0 3070 0 -1 7030
box -6 -8 126 268
use XOR2X1  _3087_
timestamp 0
transform 1 0 4450 0 1 7030
box -6 -8 126 268
use MUX2X1  _3088_
timestamp 0
transform -1 0 5150 0 1 7030
box -6 -8 126 268
use NAND2X1  _3089_
timestamp 0
transform 1 0 3530 0 -1 12230
box -6 -8 86 268
use OAI21X1  _3090_
timestamp 0
transform -1 0 3890 0 -1 12230
box -6 -8 106 268
use NAND2X1  _3091_
timestamp 0
transform -1 0 6430 0 -1 11190
box -6 -8 86 268
use INVX2  _3092_
timestamp 0
transform 1 0 5570 0 1 9110
box -6 -8 66 268
use OAI21X1  _3093_
timestamp 0
transform 1 0 5830 0 1 10150
box -6 -8 106 268
use OAI21X1  _3094_
timestamp 0
transform 1 0 5550 0 1 10150
box -6 -8 106 268
use OAI21X1  _3095_
timestamp 0
transform -1 0 4830 0 1 9110
box -6 -8 106 268
use OAI21X1  _3096_
timestamp 0
transform 1 0 4450 0 1 9110
box -6 -8 106 268
use OAI21X1  _3097_
timestamp 0
transform -1 0 4290 0 -1 9630
box -6 -8 106 268
use OAI21X1  _3098_
timestamp 0
transform 1 0 3910 0 -1 9630
box -6 -8 106 268
use OAI21X1  _3099_
timestamp 0
transform -1 0 4050 0 1 10150
box -6 -8 106 268
use OAI21X1  _3100_
timestamp 0
transform -1 0 3870 0 -1 10150
box -6 -8 106 268
use OAI21X1  _3101_
timestamp 0
transform 1 0 5010 0 1 9110
box -6 -8 106 268
use OAI21X1  _3102_
timestamp 0
transform -1 0 5390 0 1 9110
box -6 -8 106 268
use OAI21X1  _3103_
timestamp 0
transform -1 0 4770 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3104_
timestamp 0
transform -1 0 5050 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3105_
timestamp 0
transform 1 0 5750 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3106_
timestamp 0
transform -1 0 6150 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3107_
timestamp 0
transform -1 0 4230 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3108_
timestamp 0
transform 1 0 3850 0 -1 11190
box -6 -8 106 268
use NAND2X1  _3109_
timestamp 0
transform 1 0 6330 0 1 11190
box -6 -8 86 268
use INVX2  _3110_
timestamp 0
transform 1 0 4010 0 1 10670
box -6 -8 66 268
use OAI21X1  _3111_
timestamp 0
transform 1 0 5870 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3112_
timestamp 0
transform -1 0 5370 0 1 10670
box -6 -8 106 268
use OAI21X1  _3113_
timestamp 0
transform -1 0 4830 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3114_
timestamp 0
transform 1 0 4450 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3115_
timestamp 0
transform 1 0 4970 0 1 9630
box -6 -8 106 268
use OAI21X1  _3116_
timestamp 0
transform 1 0 3910 0 1 9630
box -6 -8 106 268
use OAI21X1  _3117_
timestamp 0
transform 1 0 4530 0 -1 11710
box -6 -8 106 268
use OAI21X1  _3118_
timestamp 0
transform -1 0 4910 0 -1 11710
box -6 -8 106 268
use OAI21X1  _3119_
timestamp 0
transform 1 0 5010 0 1 10150
box -6 -8 106 268
use OAI21X1  _3120_
timestamp 0
transform 1 0 4730 0 1 10150
box -6 -8 106 268
use OAI21X1  _3121_
timestamp 0
transform 1 0 5310 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3122_
timestamp 0
transform 1 0 5590 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3123_
timestamp 0
transform 1 0 5570 0 -1 11710
box -6 -8 106 268
use OAI21X1  _3124_
timestamp 0
transform -1 0 5950 0 -1 11710
box -6 -8 106 268
use OAI21X1  _3125_
timestamp 0
transform -1 0 4310 0 1 11190
box -6 -8 106 268
use OAI21X1  _3126_
timestamp 0
transform 1 0 3930 0 1 11190
box -6 -8 106 268
use NAND2X1  _3127_
timestamp 0
transform 1 0 6590 0 1 11190
box -6 -8 86 268
use NAND2X1  _3128_
timestamp 0
transform 1 0 6150 0 -1 10670
box -6 -8 86 268
use OAI21X1  _3129_
timestamp 0
transform 1 0 5550 0 1 10670
box -6 -8 106 268
use NAND2X1  _3130_
timestamp 0
transform -1 0 3530 0 1 10670
box -6 -8 86 268
use OAI21X1  _3131_
timestamp 0
transform -1 0 3790 0 -1 10670
box -6 -8 106 268
use NAND2X1  _3132_
timestamp 0
transform 1 0 4810 0 -1 10150
box -6 -8 86 268
use OAI21X1  _3133_
timestamp 0
transform 1 0 4050 0 -1 10150
box -6 -8 106 268
use NAND2X1  _3134_
timestamp 0
transform 1 0 5230 0 1 11710
box -6 -8 86 268
use OAI21X1  _3135_
timestamp 0
transform 1 0 4950 0 1 11710
box -6 -8 106 268
use NAND2X1  _3136_
timestamp 0
transform 1 0 5830 0 1 9630
box -6 -8 86 268
use OAI21X1  _3137_
timestamp 0
transform 1 0 5550 0 1 9630
box -6 -8 106 268
use NAND2X1  _3138_
timestamp 0
transform 1 0 5830 0 -1 10150
box -6 -8 86 268
use OAI21X1  _3139_
timestamp 0
transform 1 0 5550 0 -1 10150
box -6 -8 106 268
use NAND2X1  _3140_
timestamp 0
transform -1 0 5810 0 -1 12230
box -6 -8 86 268
use OAI21X1  _3141_
timestamp 0
transform -1 0 6090 0 -1 12230
box -6 -8 106 268
use NAND2X1  _3142_
timestamp 0
transform -1 0 4410 0 -1 12230
box -6 -8 86 268
use OAI21X1  _3143_
timestamp 0
transform -1 0 4690 0 -1 12230
box -6 -8 106 268
use AOI21X1  _3144_
timestamp 0
transform 1 0 11690 0 1 1310
box -6 -8 106 268
use OAI21X1  _3145_
timestamp 0
transform 1 0 11930 0 -1 1310
box -6 -8 106 268
use NOR2X1  _3146_
timestamp 0
transform -1 0 12050 0 1 1310
box -6 -8 86 268
use OAI21X1  _3147_
timestamp 0
transform 1 0 9610 0 1 790
box -6 -8 106 268
use NOR2X1  _3148_
timestamp 0
transform -1 0 12050 0 1 790
box -6 -8 86 268
use OAI21X1  _3149_
timestamp 0
transform -1 0 11690 0 -1 1830
box -6 -8 106 268
use NAND3X1  _3150_
timestamp 0
transform -1 0 11990 0 -1 1830
box -6 -8 106 268
use OAI21X1  _3151_
timestamp 0
transform -1 0 10910 0 -1 1830
box -6 -8 106 268
use OAI21X1  _3152_
timestamp 0
transform 1 0 9470 0 -1 1830
box -6 -8 106 268
use NAND3X1  _3153_
timestamp 0
transform -1 0 9850 0 -1 1830
box -6 -8 106 268
use NOR2X1  _3154_
timestamp 0
transform -1 0 10350 0 -1 1830
box -6 -8 86 268
use INVX1  _3155_
timestamp 0
transform -1 0 10450 0 -1 2350
box -6 -8 66 268
use OAI21X1  _3156_
timestamp 0
transform -1 0 9130 0 -1 2870
box -6 -8 106 268
use AOI21X1  _3157_
timestamp 0
transform -1 0 9170 0 1 2870
box -6 -8 106 268
use NAND3X1  _3158_
timestamp 0
transform -1 0 8890 0 1 2870
box -6 -8 106 268
use NOR2X1  _3159_
timestamp 0
transform -1 0 8850 0 -1 2870
box -6 -8 86 268
use OAI21X1  _3160_
timestamp 0
transform 1 0 10630 0 1 2350
box -6 -8 106 268
use OAI21X1  _3161_
timestamp 0
transform 1 0 10350 0 1 2350
box -6 -8 106 268
use INVX1  _3162_
timestamp 0
transform -1 0 9930 0 1 2350
box -6 -8 66 268
use NOR2X1  _3163_
timestamp 0
transform 1 0 9610 0 1 2350
box -6 -8 86 268
use AND2X2  _3164_
timestamp 0
transform -1 0 9170 0 1 2350
box -6 -8 106 268
use NAND2X1  _3165_
timestamp 0
transform -1 0 7390 0 1 1830
box -6 -8 86 268
use AOI22X1  _3166_
timestamp 0
transform 1 0 7710 0 1 1310
box -6 -8 126 268
use NAND3X1  _3167_
timestamp 0
transform 1 0 7570 0 1 1830
box -6 -8 106 268
use NOR2X1  _3168_
timestamp 0
transform 1 0 7730 0 1 2350
box -6 -8 86 268
use NAND3X1  _3169_
timestamp 0
transform -1 0 8890 0 1 2350
box -6 -8 106 268
use NOR2X1  _3170_
timestamp 0
transform -1 0 8590 0 -1 2350
box -6 -8 86 268
use NOR2X1  _3171_
timestamp 0
transform -1 0 9310 0 -1 4430
box -6 -8 86 268
use AND2X2  _3172_
timestamp 0
transform -1 0 8330 0 -1 2350
box -6 -8 106 268
use OAI21X1  _3173_
timestamp 0
transform 1 0 8510 0 1 2350
box -6 -8 106 268
use NOR2X1  _3174_
timestamp 0
transform 1 0 7990 0 1 2350
box -6 -8 86 268
use AND2X2  _3175_
timestamp 0
transform -1 0 8050 0 -1 2350
box -6 -8 106 268
use NAND3X1  _3176_
timestamp 0
transform -1 0 7770 0 -1 2350
box -6 -8 106 268
use NOR2X1  _3177_
timestamp 0
transform -1 0 12030 0 -1 2870
box -6 -8 86 268
use AND2X2  _3178_
timestamp 0
transform -1 0 11990 0 1 1830
box -6 -8 106 268
use NAND3X1  _3179_
timestamp 0
transform 1 0 12190 0 -1 1830
box -6 -8 106 268
use INVX1  _3180_
timestamp 0
transform 1 0 12230 0 1 790
box -6 -8 66 268
use NAND2X1  _3181_
timestamp 0
transform 1 0 12210 0 -1 1310
box -6 -8 86 268
use OAI21X1  _3182_
timestamp 0
transform -1 0 11510 0 -1 2350
box -6 -8 106 268
use OAI21X1  _3183_
timestamp 0
transform 1 0 11690 0 -1 2350
box -6 -8 106 268
use NOR2X1  _3184_
timestamp 0
transform 1 0 11970 0 -1 2350
box -6 -8 86 268
use NAND3X1  _3185_
timestamp 0
transform 1 0 11990 0 1 2350
box -6 -8 106 268
use OAI21X1  _3186_
timestamp 0
transform 1 0 12170 0 1 1830
box -6 -8 106 268
use INVX1  _3187_
timestamp 0
transform 1 0 10030 0 -1 1830
box -6 -8 66 268
use INVX1  _3188_
timestamp 0
transform 1 0 10910 0 -1 2350
box -6 -8 66 268
use OAI21X1  _3189_
timestamp 0
transform -1 0 11250 0 -1 2870
box -6 -8 106 268
use OR2X2  _3190_
timestamp 0
transform 1 0 11210 0 1 2350
box -6 -8 106 268
use NOR2X1  _3191_
timestamp 0
transform 1 0 11150 0 -1 2350
box -6 -8 86 268
use NAND3X1  _3192_
timestamp 0
transform -1 0 10950 0 1 1830
box -6 -8 106 268
use NOR2X1  _3193_
timestamp 0
transform 1 0 10290 0 1 1830
box -6 -8 86 268
use OAI21X1  _3194_
timestamp 0
transform 1 0 10930 0 1 2350
box -6 -8 106 268
use AND2X2  _3195_
timestamp 0
transform -1 0 10730 0 -1 2350
box -6 -8 106 268
use AOI22X1  _3196_
timestamp 0
transform 1 0 10550 0 1 1830
box -6 -8 126 268
use OAI21X1  _3197_
timestamp 0
transform -1 0 7490 0 -1 2350
box -6 -8 106 268
use NOR2X1  _3198_
timestamp 0
transform -1 0 4830 0 -1 2350
box -6 -8 86 268
use INVX2  _3199_
timestamp 0
transform 1 0 2930 0 -1 3390
box -6 -8 66 268
use OAI21X1  _3200_
timestamp 0
transform 1 0 4910 0 -1 3910
box -6 -8 106 268
use OAI21X1  _3201_
timestamp 0
transform 1 0 4630 0 -1 3910
box -6 -8 106 268
use OAI21X1  _3202_
timestamp 0
transform 1 0 1690 0 -1 3910
box -6 -8 106 268
use OAI21X1  _3203_
timestamp 0
transform 1 0 1650 0 -1 4430
box -6 -8 106 268
use OAI21X1  _3204_
timestamp 0
transform 1 0 1610 0 -1 4950
box -6 -8 106 268
use OAI21X1  _3205_
timestamp 0
transform 1 0 1170 0 1 4950
box -6 -8 106 268
use OAI21X1  _3206_
timestamp 0
transform 1 0 1590 0 1 3390
box -6 -8 106 268
use OAI21X1  _3207_
timestamp 0
transform -1 0 1810 0 1 3910
box -6 -8 106 268
use OAI21X1  _3208_
timestamp 0
transform -1 0 1150 0 -1 4950
box -6 -8 106 268
use OAI21X1  _3209_
timestamp 0
transform -1 0 870 0 -1 4950
box -6 -8 106 268
use OAI21X1  _3210_
timestamp 0
transform -1 0 4510 0 -1 4950
box -6 -8 106 268
use OAI21X1  _3211_
timestamp 0
transform 1 0 4370 0 1 4950
box -6 -8 106 268
use OAI21X1  _3212_
timestamp 0
transform 1 0 1330 0 -1 4950
box -6 -8 106 268
use OAI21X1  _3213_
timestamp 0
transform 1 0 1230 0 1 5470
box -6 -8 106 268
use OAI21X1  _3214_
timestamp 0
transform -1 0 2590 0 -1 4430
box -6 -8 106 268
use OAI21X1  _3215_
timestamp 0
transform 1 0 1930 0 -1 4430
box -6 -8 106 268
use OAI21X1  _3216_
timestamp 0
transform 1 0 5870 0 1 270
box -6 -8 106 268
use OAI21X1  _3217_
timestamp 0
transform -1 0 6250 0 1 270
box -6 -8 106 268
use NAND2X1  _3218_
timestamp 0
transform 1 0 6210 0 -1 270
box -6 -8 86 268
use OAI21X1  _3219_
timestamp 0
transform -1 0 6570 0 -1 270
box -6 -8 106 268
use NAND2X1  _3220_
timestamp 0
transform 1 0 3830 0 -1 270
box -6 -8 86 268
use OAI21X1  _3221_
timestamp 0
transform -1 0 4190 0 -1 270
box -6 -8 106 268
use INVX1  _3222_
timestamp 0
transform -1 0 3750 0 -1 2350
box -6 -8 66 268
use NAND2X1  _3223_
timestamp 0
transform 1 0 3430 0 -1 790
box -6 -8 86 268
use OAI21X1  _3224_
timestamp 0
transform -1 0 3510 0 -1 2350
box -6 -8 106 268
use NAND2X1  _3225_
timestamp 0
transform 1 0 5550 0 -1 1310
box -6 -8 86 268
use OAI21X1  _3226_
timestamp 0
transform 1 0 5270 0 -1 1310
box -6 -8 106 268
use NAND2X1  _3227_
timestamp 0
transform -1 0 4450 0 -1 270
box -6 -8 86 268
use OAI21X1  _3228_
timestamp 0
transform -1 0 4670 0 1 270
box -6 -8 106 268
use NAND2X1  _3229_
timestamp 0
transform 1 0 2830 0 1 1830
box -6 -8 86 268
use OAI21X1  _3230_
timestamp 0
transform -1 0 2950 0 -1 2350
box -6 -8 106 268
use NAND2X1  _3231_
timestamp 0
transform 1 0 6110 0 1 790
box -6 -8 86 268
use OAI21X1  _3232_
timestamp 0
transform 1 0 6090 0 -1 1310
box -6 -8 106 268
use DFFSR  _3233_
timestamp 0
transform -1 0 11770 0 1 270
box -6 -8 486 268
use DFFSR  _3234_
timestamp 0
transform -1 0 11870 0 -1 790
box -6 -8 486 268
use DFFSR  _3235_
timestamp 0
transform -1 0 10850 0 -1 270
box -6 -8 486 268
use DFFSR  _3236_
timestamp 0
transform -1 0 9510 0 1 5470
box -6 -8 486 268
use DFFSR  _3237_
timestamp 0
transform -1 0 9090 0 1 6510
box -6 -8 486 268
use DFFSR  _3238_
timestamp 0
transform 1 0 9630 0 1 6510
box -6 -8 486 268
use DFFSR  _3239_
timestamp 0
transform 1 0 5170 0 1 2350
box -6 -8 486 268
use DFFSR  _3240_
timestamp 0
transform 1 0 810 0 -1 1310
box -6 -8 486 268
use DFFSR  _3241_
timestamp 0
transform 1 0 10 0 1 790
box -6 -8 486 268
use DFFSR  _3242_
timestamp 0
transform 1 0 810 0 1 1830
box -6 -8 486 268
use DFFSR  _3243_
timestamp 0
transform 1 0 790 0 1 3910
box -6 -8 486 268
use DFFSR  _3244_
timestamp 0
transform -1 0 1030 0 -1 3910
box -6 -8 486 268
use DFFSR  _3245_
timestamp 0
transform 1 0 2410 0 1 2870
box -6 -8 486 268
use DFFSR  _3246_
timestamp 0
transform 1 0 1330 0 1 2350
box -6 -8 486 268
use DFFSR  _3247_
timestamp 0
transform 1 0 2150 0 -1 270
box -6 -8 486 268
use DFFSR  _3248_
timestamp 0
transform 1 0 1390 0 -1 270
box -6 -8 486 268
use DFFSR  _3249_
timestamp 0
transform 1 0 2370 0 1 270
box -6 -8 486 268
use DFFSR  _3250_
timestamp 0
transform 1 0 1530 0 -1 1310
box -6 -8 486 268
use DFFSR  _3251_
timestamp 0
transform 1 0 1810 0 1 2350
box -6 -8 486 268
use DFFSR  _3252_
timestamp 0
transform 1 0 10 0 -1 790
box -6 -8 486 268
use DFFSR  _3253_
timestamp 0
transform 1 0 1670 0 -1 2350
box -6 -8 486 268
use DFFSR  _3254_
timestamp 0
transform -1 0 3530 0 1 1310
box -6 -8 486 268
use DFFSR  _3255_
timestamp 0
transform -1 0 8050 0 -1 270
box -6 -8 486 268
use DFFSR  _3256_
timestamp 0
transform -1 0 8470 0 1 270
box -6 -8 486 268
use DFFSR  _3257_
timestamp 0
transform -1 0 10510 0 -1 7550
box -6 -8 486 268
use DFFSR  _3258_
timestamp 0
transform -1 0 8370 0 1 6510
box -6 -8 486 268
use DFFSR  _3259_
timestamp 0
transform -1 0 7830 0 1 7030
box -6 -8 486 268
use DFFSR  _3260_
timestamp 0
transform -1 0 9730 0 -1 7550
box -6 -8 486 268
use DFFSR  _3261_
timestamp 0
transform -1 0 8050 0 -1 7030
box -6 -8 486 268
use DFFSR  _3262_
timestamp 0
transform 1 0 7770 0 1 9110
box -6 -8 486 268
use DFFSR  _3263_
timestamp 0
transform -1 0 8370 0 -1 9110
box -6 -8 486 268
use DFFSR  _3264_
timestamp 0
transform -1 0 8250 0 -1 8590
box -6 -8 486 268
use DFFSR  _3265_
timestamp 0
transform -1 0 8070 0 1 8070
box -6 -8 486 268
use DFFSR  _3266_
timestamp 0
transform -1 0 8190 0 -1 8070
box -6 -8 486 268
use DFFSR  _3267_
timestamp 0
transform 1 0 6850 0 1 6510
box -6 -8 486 268
use DFFSR  _3268_
timestamp 0
transform -1 0 10250 0 -1 8070
box -6 -8 486 268
use DFFSR  _3269_
timestamp 0
transform -1 0 8130 0 -1 7550
box -6 -8 486 268
use DFFSR  _3270_
timestamp 0
transform 1 0 7150 0 1 10670
box -6 -8 486 268
use DFFSR  _3271_
timestamp 0
transform -1 0 8950 0 -1 11190
box -6 -8 486 268
use DFFSR  _3272_
timestamp 0
transform 1 0 8230 0 1 10150
box -6 -8 486 268
use DFFSR  _3273_
timestamp 0
transform -1 0 7670 0 1 11190
box -6 -8 486 268
use DFFSR  _3274_
timestamp 0
transform -1 0 9510 0 -1 8070
box -6 -8 486 268
use DFFSR  _3275_
timestamp 0
transform 1 0 6130 0 1 10670
box -6 -8 486 268
use DFFSR  _3276_
timestamp 0
transform -1 0 8550 0 1 9630
box -6 -8 486 268
use DFFSR  _3277_
timestamp 0
transform -1 0 8010 0 1 7550
box -6 -8 486 268
use DFFSR  _3278_
timestamp 0
transform -1 0 5410 0 1 7550
box -6 -8 486 268
use DFFSR  _3279_
timestamp 0
transform -1 0 6110 0 -1 7550
box -6 -8 486 268
use DFFSR  _3280_
timestamp 0
transform 1 0 8370 0 1 8070
box -6 -8 486 268
use DFFSR  _3281_
timestamp 0
transform -1 0 9250 0 1 11190
box -6 -8 486 268
use DFFSR  _3282_
timestamp 0
transform -1 0 10450 0 1 8070
box -6 -8 486 268
use DFFSR  _3283_
timestamp 0
transform -1 0 9410 0 -1 9110
box -6 -8 486 268
use DFFSR  _3284_
timestamp 0
transform -1 0 9930 0 1 7030
box -6 -8 486 268
use DFFSR  _3285_
timestamp 0
transform -1 0 8450 0 -1 11710
box -6 -8 486 268
use DFFSR  _3286_
timestamp 0
transform -1 0 10010 0 1 11710
box -6 -8 486 268
use DFFSR  _3287_
timestamp 0
transform -1 0 8450 0 -1 12230
box -6 -8 486 268
use DFFSR  _3288_
timestamp 0
transform -1 0 9450 0 -1 12230
box -6 -8 486 268
use DFFSR  _3289_
timestamp 0
transform 1 0 9450 0 -1 12230
box -6 -8 486 268
use DFFSR  _3290_
timestamp 0
transform -1 0 1230 0 -1 4430
box -6 -8 486 268
use DFFSR  _3291_
timestamp 0
transform -1 0 490 0 1 270
box -6 -8 486 268
use DFFSR  _3292_
timestamp 0
transform -1 0 1610 0 -1 6510
box -6 -8 486 268
use DFFSR  _3293_
timestamp 0
transform -1 0 4950 0 1 4950
box -6 -8 486 268
use DFFSR  _3294_
timestamp 0
transform 1 0 2130 0 -1 5470
box -6 -8 486 268
use DFFSR  _3295_
timestamp 0
transform -1 0 990 0 1 4950
box -6 -8 486 268
use DFFSR  _3296_
timestamp 0
transform -1 0 1570 0 1 5990
box -6 -8 486 268
use DFFSR  _3297_
timestamp 0
transform 1 0 5790 0 1 4950
box -6 -8 486 268
use DFFSR  _3298_
timestamp 0
transform -1 0 3430 0 -1 2870
box -6 -8 486 268
use DFFPOSX1  _3299_
timestamp 0
transform 1 0 4790 0 -1 8590
box -6 -8 246 268
use DFFPOSX1  _3300_
timestamp 0
transform 1 0 5470 0 1 8070
box -6 -8 246 268
use DFFPOSX1  _3301_
timestamp 0
transform 1 0 6450 0 1 9110
box -6 -8 246 268
use DFFPOSX1  _3302_
timestamp 0
transform 1 0 7550 0 -1 10150
box -6 -8 246 268
use DFFPOSX1  _3303_
timestamp 0
transform -1 0 6470 0 -1 9630
box -6 -8 246 268
use DFFPOSX1  _3304_
timestamp 0
transform 1 0 6690 0 1 10150
box -6 -8 246 268
use DFFPOSX1  _3305_
timestamp 0
transform -1 0 6110 0 1 8590
box -6 -8 246 268
use DFFPOSX1  _3306_
timestamp 0
transform 1 0 6750 0 -1 9630
box -6 -8 246 268
use DFFSR  _3307_
timestamp 0
transform -1 0 8230 0 1 10150
box -6 -8 486 268
use DFFSR  _3308_
timestamp 0
transform -1 0 4690 0 -1 7030
box -6 -8 486 268
use DFFSR  _3309_
timestamp 0
transform -1 0 5450 0 -1 8070
box -6 -8 486 268
use DFFSR  _3310_
timestamp 0
transform -1 0 6550 0 -1 5990
box -6 -8 486 268
use DFFSR  _3311_
timestamp 0
transform -1 0 5430 0 -1 7030
box -6 -8 486 268
use DFFSR  _3312_
timestamp 0
transform -1 0 5990 0 -1 6510
box -6 -8 486 268
use DFFSR  _3313_
timestamp 0
transform 1 0 6650 0 -1 7550
box -6 -8 486 268
use DFFSR  _3314_
timestamp 0
transform -1 0 6650 0 1 4430
box -6 -8 486 268
use DFFSR  _3315_
timestamp 0
transform -1 0 5870 0 1 8590
box -6 -8 486 268
use DFFSR  _3316_
timestamp 0
transform -1 0 4370 0 -1 9110
box -6 -8 486 268
use DFFSR  _3317_
timestamp 0
transform -1 0 3590 0 -1 10150
box -6 -8 486 268
use DFFSR  _3318_
timestamp 0
transform -1 0 4270 0 1 11710
box -6 -8 486 268
use DFFSR  _3319_
timestamp 0
transform 1 0 4030 0 -1 8590
box -6 -8 486 268
use DFFSR  _3320_
timestamp 0
transform 1 0 4910 0 -1 11710
box -6 -8 486 268
use DFFSR  _3321_
timestamp 0
transform 1 0 6850 0 -1 12230
box -6 -8 486 268
use DFFSR  _3322_
timestamp 0
transform -1 0 3350 0 -1 12230
box -6 -8 486 268
use DFFSR  _3323_
timestamp 0
transform -1 0 6690 0 1 10150
box -6 -8 486 268
use DFFSR  _3324_
timestamp 0
transform -1 0 4270 0 1 9110
box -6 -8 486 268
use DFFSR  _3325_
timestamp 0
transform -1 0 3790 0 1 9110
box -6 -8 486 268
use DFFSR  _3326_
timestamp 0
transform 1 0 3290 0 1 10150
box -6 -8 486 268
use DFFSR  _3327_
timestamp 0
transform 1 0 4370 0 -1 9110
box -6 -8 486 268
use DFFSR  _3328_
timestamp 0
transform -1 0 5090 0 1 11190
box -6 -8 486 268
use DFFSR  _3329_
timestamp 0
transform -1 0 6910 0 -1 11190
box -6 -8 486 268
use DFFSR  _3330_
timestamp 0
transform -1 0 3670 0 -1 11190
box -6 -8 486 268
use DFFSR  _3331_
timestamp 0
transform -1 0 6710 0 -1 10670
box -6 -8 486 268
use DFFSR  _3332_
timestamp 0
transform -1 0 3270 0 1 10670
box -6 -8 486 268
use DFFSR  _3333_
timestamp 0
transform 1 0 4010 0 1 9630
box -6 -8 486 268
use DFFSR  _3334_
timestamp 0
transform 1 0 5310 0 1 11710
box -6 -8 486 268
use DFFSR  _3335_
timestamp 0
transform 1 0 4050 0 1 10150
box -6 -8 486 268
use DFFSR  _3336_
timestamp 0
transform 1 0 4350 0 1 10670
box -6 -8 486 268
use DFFSR  _3337_
timestamp 0
transform -1 0 6270 0 1 11710
box -6 -8 486 268
use DFFSR  _3338_
timestamp 0
transform 1 0 3270 0 1 11190
box -6 -8 486 268
use DFFSR  _3339_
timestamp 0
transform -1 0 4970 0 -1 8070
box -6 -8 486 268
use DFFSR  _3340_
timestamp 0
transform 1 0 5650 0 1 10670
box -6 -8 486 268
use DFFSR  _3341_
timestamp 0
transform -1 0 4270 0 -1 10670
box -6 -8 486 268
use DFFSR  _3342_
timestamp 0
transform 1 0 4150 0 -1 10150
box -6 -8 486 268
use DFFSR  _3343_
timestamp 0
transform -1 0 4750 0 1 11710
box -6 -8 486 268
use DFFSR  _3344_
timestamp 0
transform 1 0 4930 0 -1 9630
box -6 -8 486 268
use DFFSR  _3345_
timestamp 0
transform 1 0 4890 0 -1 10150
box -6 -8 486 268
use DFFSR  _3346_
timestamp 0
transform -1 0 6570 0 -1 12230
box -6 -8 486 268
use DFFSR  _3347_
timestamp 0
transform -1 0 5170 0 -1 12230
box -6 -8 486 268
use DFFSR  _3348_
timestamp 0
transform 1 0 5090 0 1 3910
box -6 -8 486 268
use DFFSR  _3349_
timestamp 0
transform 1 0 1810 0 1 3910
box -6 -8 486 268
use DFFSR  _3350_
timestamp 0
transform 1 0 1550 0 1 4950
box -6 -8 486 268
use DFFSR  _3351_
timestamp 0
transform 1 0 1030 0 -1 3910
box -6 -8 486 268
use DFFSR  _3352_
timestamp 0
transform 1 0 1050 0 1 4430
box -6 -8 486 268
use DFFSR  _3353_
timestamp 0
transform -1 0 4190 0 1 4950
box -6 -8 486 268
use DFFSR  _3354_
timestamp 0
transform 1 0 790 0 -1 5470
box -6 -8 486 268
use DFFSR  _3355_
timestamp 0
transform 1 0 1810 0 1 4430
box -6 -8 486 268
use DFFSR  _3356_
timestamp 0
transform 1 0 6250 0 1 270
box -6 -8 486 268
use DFFSR  _3357_
timestamp 0
transform 1 0 6970 0 1 270
box -6 -8 486 268
use DFFSR  _3358_
timestamp 0
transform -1 0 4130 0 1 270
box -6 -8 486 268
use DFFSR  _3359_
timestamp 0
transform 1 0 3010 0 1 2350
box -6 -8 486 268
use DFFSR  _3360_
timestamp 0
transform -1 0 5090 0 -1 1310
box -6 -8 486 268
use DFFSR  _3361_
timestamp 0
transform -1 0 5150 0 1 270
box -6 -8 486 268
use DFFSR  _3362_
timestamp 0
transform 1 0 2290 0 1 2350
box -6 -8 486 268
use DFFSR  _3363_
timestamp 0
transform -1 0 8450 0 1 790
box -6 -8 486 268
use OR2X2  _3364_
timestamp 0
transform 1 0 5370 0 -1 5990
box -6 -8 106 268
use NOR2X1  _3365_
timestamp 0
transform 1 0 4570 0 -1 5990
box -6 -8 86 268
use NOR2X1  _3366_
timestamp 0
transform 1 0 5050 0 1 5990
box -6 -8 86 268
use NOR2X1  _3367_
timestamp 0
transform -1 0 4910 0 -1 5990
box -6 -8 86 268
use NAND3X1  _3368_
timestamp 0
transform -1 0 5190 0 -1 5990
box -6 -8 106 268
use NOR2X1  _3369_
timestamp 0
transform -1 0 5750 0 -1 5990
box -6 -8 86 268
use XOR2X1  _3370_
timestamp 0
transform 1 0 2810 0 1 7030
box -6 -8 126 268
use XNOR2X1  _3371_
timestamp 0
transform 1 0 2310 0 1 7550
box -6 -8 126 268
use XNOR2X1  _3372_
timestamp 0
transform -1 0 2530 0 -1 7550
box -6 -8 126 268
use INVX4  _3373_
timestamp 0
transform -1 0 4150 0 -1 12230
box -6 -8 86 268
use INVX4  _3374_
timestamp 0
transform -1 0 2470 0 1 11190
box -6 -8 86 268
use NAND2X1  _3375_
timestamp 0
transform 1 0 2410 0 -1 8590
box -6 -8 86 268
use INVX2  _3376_
timestamp 0
transform -1 0 3110 0 -1 10150
box -6 -8 66 268
use NAND2X1  _3377_
timestamp 0
transform 1 0 2530 0 -1 10150
box -6 -8 86 268
use INVX2  _3378_
timestamp 0
transform -1 0 2430 0 -1 9630
box -6 -8 66 268
use AND2X2  _3379_
timestamp 0
transform -1 0 1630 0 -1 8070
box -6 -8 106 268
use NAND2X1  _3380_
timestamp 0
transform 1 0 1330 0 1 8070
box -6 -8 86 268
use AOI22X1  _3381_
timestamp 0
transform -1 0 1690 0 -1 8590
box -6 -8 126 268
use INVX2  _3382_
timestamp 0
transform -1 0 2090 0 -1 10150
box -6 -8 66 268
use OAI21X1  _3383_
timestamp 0
transform -1 0 1690 0 1 8070
box -6 -8 106 268
use OAI21X1  _3384_
timestamp 0
transform 1 0 1890 0 -1 8590
box -6 -8 106 268
use INVX4  _3385_
timestamp 0
transform 1 0 1570 0 1 10150
box -6 -8 86 268
use OAI21X1  _3386_
timestamp 0
transform -1 0 2230 0 -1 9110
box -6 -8 106 268
use AOI21X1  _3387_
timestamp 0
transform 1 0 2410 0 -1 9110
box -6 -8 106 268
use NOR2X1  _3388_
timestamp 0
transform -1 0 810 0 -1 11190
box -6 -8 86 268
use AOI21X1  _3389_
timestamp 0
transform 1 0 2610 0 -1 9630
box -6 -8 106 268
use NAND2X1  _3390_
timestamp 0
transform 1 0 3430 0 -1 10670
box -6 -8 86 268
use OAI21X1  _3391_
timestamp 0
transform 1 0 3150 0 -1 10670
box -6 -8 106 268
use INVX1  _3392_
timestamp 0
transform -1 0 3030 0 -1 8590
box -6 -8 66 268
use OAI21X1  _3393_
timestamp 0
transform 1 0 2390 0 1 9110
box -6 -8 106 268
use NAND2X1  _3394_
timestamp 0
transform 1 0 790 0 1 8070
box -6 -8 86 268
use AND2X2  _3395_
timestamp 0
transform -1 0 830 0 -1 8070
box -6 -8 106 268
use NAND2X1  _3396_
timestamp 0
transform -1 0 550 0 -1 8070
box -6 -8 86 268
use AOI22X1  _3397_
timestamp 0
transform -1 0 610 0 1 8070
box -6 -8 126 268
use OAI21X1  _3398_
timestamp 0
transform -1 0 290 0 -1 8070
box -6 -8 106 268
use OAI21X1  _3399_
timestamp 0
transform 1 0 210 0 1 8070
box -6 -8 106 268
use NAND2X1  _3400_
timestamp 0
transform -1 0 1050 0 1 9630
box -6 -8 86 268
use INVX2  _3401_
timestamp 0
transform -1 0 1610 0 -1 10670
box -6 -8 66 268
use OAI21X1  _3402_
timestamp 0
transform 1 0 1550 0 -1 9630
box -6 -8 106 268
use OAI21X1  _3403_
timestamp 0
transform 1 0 1270 0 -1 9630
box -6 -8 106 268
use NAND2X1  _3404_
timestamp 0
transform -1 0 270 0 -1 7550
box -6 -8 86 268
use AND2X2  _3405_
timestamp 0
transform -1 0 550 0 -1 7030
box -6 -8 106 268
use NAND2X1  _3406_
timestamp 0
transform -1 0 270 0 -1 7030
box -6 -8 86 268
use AOI22X1  _3407_
timestamp 0
transform -1 0 590 0 1 7550
box -6 -8 126 268
use OAI21X1  _3408_
timestamp 0
transform -1 0 290 0 1 7030
box -6 -8 106 268
use OAI21X1  _3409_
timestamp 0
transform -1 0 290 0 1 7550
box -6 -8 106 268
use OAI21X1  _3410_
timestamp 0
transform 1 0 1530 0 1 9110
box -6 -8 106 268
use OAI21X1  _3411_
timestamp 0
transform 1 0 1250 0 1 9110
box -6 -8 106 268
use NAND2X1  _3412_
timestamp 0
transform -1 0 790 0 1 9110
box -6 -8 86 268
use NAND2X1  _3413_
timestamp 0
transform 1 0 490 0 1 7030
box -6 -8 86 268
use AND2X2  _3414_
timestamp 0
transform 1 0 730 0 -1 7030
box -6 -8 106 268
use NAND2X1  _3415_
timestamp 0
transform -1 0 1110 0 1 7030
box -6 -8 86 268
use AOI22X1  _3416_
timestamp 0
transform 1 0 730 0 -1 7550
box -6 -8 126 268
use OAI21X1  _3417_
timestamp 0
transform -1 0 850 0 1 7030
box -6 -8 106 268
use OAI21X1  _3418_
timestamp 0
transform -1 0 550 0 -1 7550
box -6 -8 106 268
use OAI21X1  _3419_
timestamp 0
transform -1 0 1370 0 -1 9110
box -6 -8 106 268
use OAI21X1  _3420_
timestamp 0
transform 1 0 990 0 -1 9110
box -6 -8 106 268
use NAND2X1  _3421_
timestamp 0
transform 1 0 1290 0 1 7030
box -6 -8 86 268
use AND2X2  _3422_
timestamp 0
transform 1 0 1010 0 -1 8070
box -6 -8 106 268
use NAND2X1  _3423_
timestamp 0
transform 1 0 1310 0 1 7550
box -6 -8 86 268
use AOI22X1  _3424_
timestamp 0
transform -1 0 1430 0 -1 7550
box -6 -8 126 268
use OAI21X1  _3425_
timestamp 0
transform -1 0 1130 0 1 7550
box -6 -8 106 268
use OAI21X1  _3426_
timestamp 0
transform 1 0 1030 0 -1 7550
box -6 -8 106 268
use OAI21X1  _3427_
timestamp 0
transform -1 0 1630 0 1 9630
box -6 -8 106 268
use OAI21X1  _3428_
timestamp 0
transform 1 0 1250 0 1 9630
box -6 -8 106 268
use NAND2X1  _3429_
timestamp 0
transform -1 0 1070 0 -1 10150
box -6 -8 86 268
use INVX1  _3430_
timestamp 0
transform 1 0 1530 0 -1 10150
box -6 -8 66 268
use AND2X2  _3431_
timestamp 0
transform 1 0 1250 0 -1 10150
box -6 -8 106 268
use OAI21X1  _3432_
timestamp 0
transform -1 0 1130 0 1 10150
box -6 -8 106 268
use INVX1  _3433_
timestamp 0
transform -1 0 250 0 -1 11190
box -6 -8 66 268
use NAND2X1  _3434_
timestamp 0
transform -1 0 850 0 1 7550
box -6 -8 86 268
use NAND3X1  _3435_
timestamp 0
transform -1 0 1150 0 1 8070
box -6 -8 106 268
use AOI22X1  _3436_
timestamp 0
transform -1 0 1110 0 -1 8590
box -6 -8 126 268
use INVX1  _3437_
timestamp 0
transform 1 0 1830 0 1 8590
box -6 -8 66 268
use INVX1  _3438_
timestamp 0
transform 1 0 1290 0 -1 8070
box -6 -8 66 268
use OAI21X1  _3439_
timestamp 0
transform -1 0 1650 0 1 8590
box -6 -8 106 268
use NAND2X1  _3440_
timestamp 0
transform 1 0 1290 0 1 8590
box -6 -8 86 268
use OAI21X1  _3441_
timestamp 0
transform -1 0 810 0 -1 8590
box -6 -8 106 268
use NOR2X1  _3442_
timestamp 0
transform 1 0 1310 0 1 10150
box -6 -8 86 268
use XOR2X1  _3443_
timestamp 0
transform 1 0 1250 0 -1 10670
box -6 -8 126 268
use NAND3X1  _3444_
timestamp 0
transform -1 0 2210 0 1 9110
box -6 -8 106 268
use AOI22X1  _3445_
timestamp 0
transform 1 0 1810 0 1 9110
box -6 -8 126 268
use INVX1  _3446_
timestamp 0
transform 1 0 2170 0 -1 8590
box -6 -8 66 268
use NOR2X1  _3447_
timestamp 0
transform 1 0 2070 0 1 8590
box -6 -8 86 268
use OAI21X1  _3448_
timestamp 0
transform -1 0 1950 0 -1 9110
box -6 -8 106 268
use OAI22X1  _3449_
timestamp 0
transform 1 0 1550 0 -1 9110
box -6 -8 126 268
use OAI21X1  _3450_
timestamp 0
transform -1 0 1090 0 -1 11190
box -6 -8 106 268
use AOI21X1  _3451_
timestamp 0
transform 1 0 1270 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3452_
timestamp 0
transform 1 0 970 0 1 11190
box -6 -8 106 268
use NAND2X1  _3453_
timestamp 0
transform -1 0 2350 0 -1 10150
box -6 -8 86 268
use NAND2X1  _3454_
timestamp 0
transform 1 0 3210 0 1 10150
box -6 -8 86 268
use AOI22X1  _3455_
timestamp 0
transform -1 0 2250 0 1 10150
box -6 -8 126 268
use INVX1  _3456_
timestamp 0
transform -1 0 1850 0 -1 10670
box -6 -8 66 268
use INVX1  _3457_
timestamp 0
transform -1 0 3030 0 1 10150
box -6 -8 66 268
use OAI21X1  _3458_
timestamp 0
transform -1 0 1950 0 1 10150
box -6 -8 106 268
use NAND2X1  _3459_
timestamp 0
transform -1 0 1850 0 -1 10150
box -6 -8 86 268
use NAND2X1  _3460_
timestamp 0
transform 1 0 1830 0 -1 9630
box -6 -8 86 268
use OAI21X1  _3461_
timestamp 0
transform -1 0 2130 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3462_
timestamp 0
transform -1 0 1890 0 -1 11190
box -6 -8 106 268
use INVX1  _3463_
timestamp 0
transform -1 0 1610 0 -1 11190
box -6 -8 66 268
use OAI21X1  _3464_
timestamp 0
transform 1 0 1290 0 1 10670
box -6 -8 106 268
use OAI21X1  _3465_
timestamp 0
transform -1 0 1630 0 1 11190
box -6 -8 106 268
use OAI21X1  _3466_
timestamp 0
transform 1 0 2090 0 -1 9630
box -6 -8 106 268
use NOR2X1  _3467_
timestamp 0
transform 1 0 2090 0 1 9630
box -6 -8 86 268
use MUX2X1  _3468_
timestamp 0
transform 1 0 2850 0 -1 10670
box -6 -8 126 268
use NAND2X1  _3469_
timestamp 0
transform 1 0 2710 0 1 10150
box -6 -8 86 268
use NAND2X1  _3470_
timestamp 0
transform -1 0 2670 0 -1 10670
box -6 -8 86 268
use AOI21X1  _3471_
timestamp 0
transform 1 0 2430 0 1 10150
box -6 -8 106 268
use NAND2X1  _3472_
timestamp 0
transform -1 0 2410 0 -1 10670
box -6 -8 86 268
use NAND3X1  _3473_
timestamp 0
transform 1 0 1570 0 1 10670
box -6 -8 106 268
use AOI22X1  _3474_
timestamp 0
transform -1 0 1930 0 1 11190
box -6 -8 126 268
use NOR2X1  _3475_
timestamp 0
transform 1 0 1310 0 -1 11710
box -6 -8 86 268
use OAI21X1  _3476_
timestamp 0
transform -1 0 1130 0 -1 11710
box -6 -8 106 268
use NAND2X1  _3477_
timestamp 0
transform 1 0 470 0 -1 11710
box -6 -8 86 268
use NAND2X1  _3478_
timestamp 0
transform -1 0 510 0 1 11190
box -6 -8 86 268
use INVX1  _3479_
timestamp 0
transform -1 0 250 0 1 11190
box -6 -8 66 268
use OAI21X1  _3480_
timestamp 0
transform -1 0 290 0 -1 11710
box -6 -8 106 268
use INVX1  _3481_
timestamp 0
transform -1 0 250 0 -1 12230
box -6 -8 66 268
use AOI22X1  _3482_
timestamp 0
transform 1 0 730 0 -1 11710
box -6 -8 126 268
use XOR2X1  _3483_
timestamp 0
transform -1 0 550 0 -1 11190
box -6 -8 126 268
use AOI21X1  _3484_
timestamp 0
transform 1 0 2070 0 -1 11190
box -6 -8 106 268
use OAI21X1  _3485_
timestamp 0
transform -1 0 2210 0 1 11190
box -6 -8 106 268
use INVX1  _3486_
timestamp 0
transform -1 0 1550 0 -1 12230
box -6 -8 66 268
use NOR2X1  _3487_
timestamp 0
transform -1 0 1910 0 -1 11710
box -6 -8 86 268
use OAI21X1  _3488_
timestamp 0
transform -1 0 1710 0 1 11710
box -6 -8 106 268
use INVX1  _3489_
timestamp 0
transform 1 0 1570 0 -1 11710
box -6 -8 66 268
use OAI21X1  _3490_
timestamp 0
transform 1 0 1250 0 1 11190
box -6 -8 106 268
use MUX2X1  _3491_
timestamp 0
transform -1 0 1430 0 1 11710
box -6 -8 126 268
use NAND2X1  _3492_
timestamp 0
transform 1 0 1230 0 -1 12230
box -6 -8 86 268
use OAI21X1  _3493_
timestamp 0
transform -1 0 1130 0 1 11710
box -6 -8 106 268
use NAND2X1  _3494_
timestamp 0
transform 1 0 970 0 -1 12230
box -6 -8 86 268
use NAND2X1  _3495_
timestamp 0
transform -1 0 790 0 -1 12230
box -6 -8 86 268
use NAND2X1  _3496_
timestamp 0
transform 1 0 490 0 1 11710
box -6 -8 86 268
use NAND3X1  _3497_
timestamp 0
transform -1 0 530 0 -1 12230
box -6 -8 106 268
use NAND3X1  _3498_
timestamp 0
transform 1 0 750 0 1 11710
box -6 -8 106 268
use NAND2X1  _3499_
timestamp 0
transform -1 0 870 0 1 10670
box -6 -8 86 268
use OAI21X1  _3500_
timestamp 0
transform 1 0 750 0 1 10150
box -6 -8 106 268
use INVX1  _3501_
timestamp 0
transform 1 0 990 0 -1 10670
box -6 -8 66 268
use OAI21X1  _3502_
timestamp 0
transform -1 0 610 0 1 10670
box -6 -8 106 268
use NAND2X1  _3503_
timestamp 0
transform -1 0 550 0 1 8590
box -6 -8 86 268
use OAI21X1  _3504_
timestamp 0
transform -1 0 810 0 -1 9110
box -6 -8 106 268
use INVX1  _3505_
timestamp 0
transform -1 0 530 0 -1 9110
box -6 -8 66 268
use OAI21X1  _3506_
timestamp 0
transform -1 0 290 0 1 8590
box -6 -8 106 268
use INVX1  _3507_
timestamp 0
transform -1 0 250 0 -1 8590
box -6 -8 66 268
use AOI22X1  _3508_
timestamp 0
transform 1 0 730 0 1 8590
box -6 -8 126 268
use OAI21X1  _3509_
timestamp 0
transform -1 0 1070 0 1 9110
box -6 -8 106 268
use INVX1  _3510_
timestamp 0
transform -1 0 530 0 1 9110
box -6 -8 66 268
use OAI21X1  _3511_
timestamp 0
transform -1 0 290 0 1 9110
box -6 -8 106 268
use OAI21X1  _3512_
timestamp 0
transform 1 0 690 0 -1 9630
box -6 -8 106 268
use NAND2X1  _3513_
timestamp 0
transform -1 0 570 0 1 10150
box -6 -8 86 268
use OAI21X1  _3514_
timestamp 0
transform -1 0 530 0 -1 10670
box -6 -8 106 268
use INVX1  _3515_
timestamp 0
transform -1 0 250 0 -1 10670
box -6 -8 66 268
use OAI21X1  _3516_
timestamp 0
transform -1 0 310 0 1 10150
box -6 -8 106 268
use INVX1  _3517_
timestamp 0
transform 1 0 750 0 -1 10150
box -6 -8 66 268
use AOI22X1  _3518_
timestamp 0
transform 1 0 970 0 -1 9630
box -6 -8 126 268
use OAI21X1  _3519_
timestamp 0
transform 1 0 2670 0 1 9110
box -6 -8 106 268
use OAI21X1  _3520_
timestamp 0
transform 1 0 2950 0 1 9110
box -6 -8 106 268
use NAND2X1  _3521_
timestamp 0
transform 1 0 3430 0 1 8590
box -6 -8 86 268
use XOR2X1  _3522_
timestamp 0
transform 1 0 3130 0 1 8590
box -6 -8 126 268
use XOR2X1  _3523_
timestamp 0
transform 1 0 2690 0 -1 9110
box -6 -8 126 268
use INVX1  _3524_
timestamp 0
transform -1 0 1110 0 1 10670
box -6 -8 66 268
use XOR2X1  _3525_
timestamp 0
transform -1 0 310 0 1 10670
box -6 -8 126 268
use XOR2X1  _3526_
timestamp 0
transform -1 0 310 0 1 11710
box -6 -8 126 268
use AOI21X1  _3527_
timestamp 0
transform -1 0 790 0 1 11190
box -6 -8 106 268
use AOI21X1  _3528_
timestamp 0
transform -1 0 810 0 -1 10670
box -6 -8 106 268
use OAI21X1  _3529_
timestamp 0
transform -1 0 290 0 -1 9110
box -6 -8 106 268
use INVX1  _3530_
timestamp 0
transform -1 0 250 0 -1 9630
box -6 -8 66 268
use NAND2X1  _3531_
timestamp 0
transform 1 0 210 0 -1 10150
box -6 -8 86 268
use NAND2X1  _3532_
timestamp 0
transform 1 0 430 0 -1 9630
box -6 -8 86 268
use NAND2X1  _3533_
timestamp 0
transform -1 0 270 0 1 9630
box -6 -8 86 268
use NAND2X1  _3534_
timestamp 0
transform -1 0 790 0 1 9630
box -6 -8 86 268
use NAND3X1  _3535_
timestamp 0
transform -1 0 570 0 -1 10150
box -6 -8 106 268
use NAND2X1  _3536_
timestamp 0
transform -1 0 530 0 1 9630
box -6 -8 86 268
use AOI21X1  _3537_
timestamp 0
transform -1 0 1910 0 1 9630
box -6 -8 106 268
use AOI21X1  _3538_
timestamp 0
transform 1 0 2590 0 1 8590
box -6 -8 106 268
use AOI22X1  _3539_
timestamp 0
transform -1 0 2790 0 -1 8590
box -6 -8 126 268
use NAND2X1  _3540_
timestamp 0
transform -1 0 2490 0 1 8070
box -6 -8 86 268
use OAI21X1  _3541_
timestamp 0
transform -1 0 2230 0 1 8070
box -6 -8 106 268
use NAND2X1  _3542_
timestamp 0
transform -1 0 2390 0 -1 12230
box -6 -8 86 268
use AOI21X1  _3543_
timestamp 0
transform 1 0 1730 0 -1 12230
box -6 -8 106 268
use OAI21X1  _3544_
timestamp 0
transform 1 0 2090 0 -1 11710
box -6 -8 106 268
use OAI21X1  _3545_
timestamp 0
transform 1 0 1890 0 1 11710
box -6 -8 106 268
use OAI21X1  _3546_
timestamp 0
transform 1 0 2030 0 -1 12230
box -6 -8 106 268
use NAND2X1  _3547_
timestamp 0
transform -1 0 2730 0 -1 11710
box -6 -8 86 268
use OAI21X1  _3548_
timestamp 0
transform 1 0 2370 0 -1 11710
box -6 -8 106 268
use NAND2X1  _3549_
timestamp 0
transform -1 0 2530 0 1 11710
box -6 -8 86 268
use OAI21X1  _3550_
timestamp 0
transform 1 0 2170 0 1 11710
box -6 -8 106 268
use NAND2X1  _3551_
timestamp 0
transform -1 0 2710 0 -1 11190
box -6 -8 86 268
use OAI21X1  _3552_
timestamp 0
transform 1 0 2350 0 -1 11190
box -6 -8 106 268
use NAND2X1  _3553_
timestamp 0
transform -1 0 1950 0 1 8070
box -6 -8 86 268
use NOR2X1  _3554_
timestamp 0
transform 1 0 1030 0 1 8590
box -6 -8 86 268
use OAI21X1  _3555_
timestamp 0
transform 1 0 430 0 -1 8590
box -6 -8 106 268
use OAI21X1  _3556_
timestamp 0
transform 1 0 1290 0 -1 8590
box -6 -8 106 268
use NAND2X1  _3557_
timestamp 0
transform -1 0 3250 0 -1 9630
box -6 -8 86 268
use OAI21X1  _3558_
timestamp 0
transform 1 0 2890 0 -1 9630
box -6 -8 106 268
use NAND2X1  _3559_
timestamp 0
transform -1 0 2710 0 1 9630
box -6 -8 86 268
use OAI21X1  _3560_
timestamp 0
transform 1 0 2350 0 1 9630
box -6 -8 106 268
use INVX1  _3561_
timestamp 0
transform -1 0 2130 0 1 7550
box -6 -8 66 268
use NAND2X1  _3562_
timestamp 0
transform -1 0 2950 0 1 8590
box -6 -8 86 268
use OAI21X1  _3563_
timestamp 0
transform 1 0 2290 0 -1 8070
box -6 -8 106 268
use INVX1  _3564_
timestamp 0
transform 1 0 2570 0 1 7030
box -6 -8 66 268
use NAND2X1  _3565_
timestamp 0
transform -1 0 1630 0 1 7030
box -6 -8 86 268
use OAI21X1  _3566_
timestamp 0
transform -1 0 1910 0 1 7030
box -6 -8 106 268
use DFFSR  _3567_
timestamp 0
transform 1 0 1670 0 1 10670
box -6 -8 486 268
use DFFSR  _3568_
timestamp 0
transform 1 0 3030 0 -1 8590
box -6 -8 486 268
use DFFSR  _3569_
timestamp 0
transform 1 0 2490 0 1 8070
box -6 -8 486 268
use DFFSR  _3570_
timestamp 0
transform 1 0 2390 0 -1 12230
box -6 -8 486 268
use DFFSR  _3571_
timestamp 0
transform 1 0 2730 0 -1 11710
box -6 -8 486 268
use DFFSR  _3572_
timestamp 0
transform 1 0 2530 0 1 11710
box -6 -8 486 268
use DFFSR  _3573_
timestamp 0
transform 1 0 2710 0 -1 11190
box -6 -8 486 268
use DFFSR  _3574_
timestamp 0
transform 1 0 1630 0 -1 8070
box -6 -8 486 268
use DFFSR  _3575_
timestamp 0
transform 1 0 3250 0 -1 9630
box -6 -8 486 268
use DFFSR  _3576_
timestamp 0
transform 1 0 2710 0 1 9630
box -6 -8 486 268
use DFFSR  _3577_
timestamp 0
transform 1 0 2390 0 -1 8070
box -6 -8 486 268
use DFFSR  _3578_
timestamp 0
transform 1 0 1910 0 1 7030
box -6 -8 486 268
use BUFX2  _3579_
timestamp 0
transform -1 0 5230 0 -1 270
box -6 -8 86 268
use BUFX2  _3580_
timestamp 0
transform -1 0 270 0 -1 4430
box -6 -8 86 268
use BUFX2  _3581_
timestamp 0
transform -1 0 3650 0 -1 270
box -6 -8 86 268
use BUFX2  _3582_
timestamp 0
transform -1 0 3390 0 -1 270
box -6 -8 86 268
use BUFX2  _3583_
timestamp 0
transform -1 0 5510 0 -1 790
box -6 -8 86 268
use BUFX2  _3584_
timestamp 0
transform 1 0 4630 0 -1 270
box -6 -8 86 268
use BUFX2  _3585_
timestamp 0
transform 1 0 3050 0 -1 270
box -6 -8 86 268
use BUFX2  _3586_
timestamp 0
transform -1 0 6030 0 -1 790
box -6 -8 86 268
use BUFX2  _3587_
timestamp 0
transform 1 0 210 0 -1 5990
box -6 -8 86 268
use BUFX2  _3588_
timestamp 0
transform -1 0 270 0 1 3910
box -6 -8 86 268
use BUFX2  _3589_
timestamp 0
transform -1 0 270 0 1 4950
box -6 -8 86 268
use BUFX2  _3590_
timestamp 0
transform -1 0 270 0 -1 5470
box -6 -8 86 268
use BUFX2  _3591_
timestamp 0
transform -1 0 550 0 -1 5990
box -6 -8 86 268
use BUFX2  _3592_
timestamp 0
transform -1 0 270 0 1 4430
box -6 -8 86 268
use BUFX2  _3593_
timestamp 0
transform -1 0 4970 0 -1 270
box -6 -8 86 268
use BUFX2  _3594_
timestamp 0
transform 1 0 5950 0 -1 270
box -6 -8 86 268
use BUFX2  _3595_
timestamp 0
transform 1 0 5690 0 -1 790
box -6 -8 86 268
use BUFX2  _3596_
timestamp 0
transform -1 0 1050 0 -1 5990
box -6 -8 86 268
use BUFX2  _3597_
timestamp 0
transform -1 0 270 0 1 5990
box -6 -8 86 268
use BUFX2  _3598_
timestamp 0
transform -1 0 530 0 1 5990
box -6 -8 86 268
use BUFX2  _3599_
timestamp 0
transform -1 0 270 0 1 6510
box -6 -8 86 268
use BUFX2  _3600_
timestamp 0
transform -1 0 270 0 -1 6510
box -6 -8 86 268
use BUFX2  _3601_
timestamp 0
transform -1 0 270 0 1 5470
box -6 -8 86 268
use BUFX2  _3602_
timestamp 0
transform -1 0 1910 0 -1 5990
box -6 -8 86 268
use BUFX2  _3603_
timestamp 0
transform 1 0 6990 0 -1 270
box -6 -8 86 268
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 8010 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 9510 0 1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 8270 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 11130 0 1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert4
timestamp 0
transform 1 0 730 0 1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert5
timestamp 0
transform -1 0 12270 0 -1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 9770 0 1 5470
box -6 -8 86 268
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 7170 0 1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 1050 0 1 5470
box -6 -8 86 268
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 10270 0 1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert10
timestamp 0
transform -1 0 1090 0 1 5990
box -6 -8 86 268
use BUFX2  BUFX2_insert11
timestamp 0
transform -1 0 6170 0 -1 4950
box -6 -8 86 268
use BUFX2  BUFX2_insert12
timestamp 0
transform 1 0 11670 0 -1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert13
timestamp 0
transform -1 0 6350 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert14
timestamp 0
transform 1 0 6910 0 1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert15
timestamp 0
transform -1 0 3510 0 -1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert16
timestamp 0
transform -1 0 4130 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert17
timestamp 0
transform 1 0 7310 0 -1 5990
box -6 -8 86 268
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 7190 0 1 11190
box -6 -8 86 268
use BUFX2  BUFX2_insert19
timestamp 0
transform 1 0 5450 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 8690 0 1 11190
box -6 -8 86 268
use BUFX2  BUFX2_insert21
timestamp 0
transform -1 0 8670 0 -1 7550
box -6 -8 86 268
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 1630 0 -1 5990
box -6 -8 86 268
use BUFX2  BUFX2_insert23
timestamp 0
transform 1 0 3550 0 -1 9110
box -6 -8 86 268
use BUFX2  BUFX2_insert24
timestamp 0
transform -1 0 4530 0 1 5470
box -6 -8 86 268
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 8290 0 -1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert26
timestamp 0
transform 1 0 5230 0 -1 11190
box -6 -8 86 268
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 1430 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert39
timestamp 0
transform 1 0 6470 0 1 4950
box -6 -8 86 268
use BUFX2  BUFX2_insert40
timestamp 0
transform 1 0 7810 0 1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert41
timestamp 0
transform -1 0 9010 0 -1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert42
timestamp 0
transform -1 0 7150 0 -1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert43
timestamp 0
transform -1 0 9050 0 -1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert44
timestamp 0
transform -1 0 9170 0 -1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert45
timestamp 0
transform 1 0 11170 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert46
timestamp 0
transform 1 0 9610 0 -1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert47
timestamp 0
transform 1 0 9330 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert48
timestamp 0
transform 1 0 7070 0 -1 9110
box -6 -8 86 268
use BUFX2  BUFX2_insert49
timestamp 0
transform 1 0 7330 0 -1 9110
box -6 -8 86 268
use BUFX2  BUFX2_insert50
timestamp 0
transform -1 0 7770 0 1 9110
box -6 -8 86 268
use BUFX2  BUFX2_insert51
timestamp 0
transform 1 0 7670 0 1 10150
box -6 -8 86 268
use BUFX2  BUFX2_insert52
timestamp 0
transform 1 0 9070 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert53
timestamp 0
transform 1 0 10130 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert54
timestamp 0
transform 1 0 8950 0 -1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert55
timestamp 0
transform 1 0 8810 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert56
timestamp 0
transform -1 0 2410 0 1 8590
box -6 -8 86 268
use BUFX2  BUFX2_insert57
timestamp 0
transform 1 0 2650 0 1 11190
box -6 -8 86 268
use BUFX2  BUFX2_insert58
timestamp 0
transform 1 0 2790 0 -1 10150
box -6 -8 86 268
use BUFX2  BUFX2_insert59
timestamp 0
transform -1 0 2410 0 1 10670
box -6 -8 86 268
use BUFX2  BUFX2_insert60
timestamp 0
transform -1 0 10670 0 1 7550
box -6 -8 86 268
use BUFX2  BUFX2_insert61
timestamp 0
transform 1 0 10670 0 -1 10150
box -6 -8 86 268
use BUFX2  BUFX2_insert62
timestamp 0
transform 1 0 10630 0 1 8070
box -6 -8 86 268
use BUFX2  BUFX2_insert63
timestamp 0
transform -1 0 9350 0 1 7550
box -6 -8 86 268
use BUFX2  BUFX2_insert64
timestamp 0
transform -1 0 8790 0 -1 8590
box -6 -8 86 268
use BUFX2  BUFX2_insert65
timestamp 0
transform 1 0 5330 0 1 270
box -6 -8 86 268
use BUFX2  BUFX2_insert66
timestamp 0
transform 1 0 5850 0 1 790
box -6 -8 86 268
use BUFX2  BUFX2_insert67
timestamp 0
transform -1 0 3210 0 -1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert68
timestamp 0
transform 1 0 3290 0 1 270
box -6 -8 86 268
use BUFX2  BUFX2_insert69
timestamp 0
transform -1 0 6830 0 -1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert70
timestamp 0
transform 1 0 8710 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert71
timestamp 0
transform -1 0 9430 0 1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert72
timestamp 0
transform -1 0 6950 0 -1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert73
timestamp 0
transform 1 0 9050 0 -1 7030
box -6 -8 86 268
use BUFX2  BUFX2_insert74
timestamp 0
transform 1 0 10910 0 1 7030
box -6 -8 86 268
use BUFX2  BUFX2_insert75
timestamp 0
transform 1 0 2690 0 1 1310
box -6 -8 86 268
use BUFX2  BUFX2_insert76
timestamp 0
transform -1 0 3250 0 -1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert77
timestamp 0
transform 1 0 10570 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert78
timestamp 0
transform 1 0 9430 0 -1 5470
box -6 -8 86 268
use BUFX2  BUFX2_insert79
timestamp 0
transform -1 0 8530 0 1 7550
box -6 -8 86 268
use BUFX2  BUFX2_insert80
timestamp 0
transform 1 0 7270 0 1 5470
box -6 -8 86 268
use BUFX2  BUFX2_insert81
timestamp 0
transform 1 0 7730 0 -1 790
box -6 -8 86 268
use BUFX2  BUFX2_insert82
timestamp 0
transform -1 0 7770 0 -1 8590
box -6 -8 86 268
use BUFX2  BUFX2_insert83
timestamp 0
transform -1 0 7570 0 -1 6510
box -6 -8 86 268
use BUFX2  BUFX2_insert84
timestamp 0
transform 1 0 9550 0 1 8590
box -6 -8 86 268
use BUFX2  BUFX2_insert85
timestamp 0
transform -1 0 9090 0 1 8590
box -6 -8 86 268
use BUFX2  BUFX2_insert86
timestamp 0
transform -1 0 9690 0 1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert87
timestamp 0
transform 1 0 9530 0 1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert88
timestamp 0
transform -1 0 10930 0 -1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert89
timestamp 0
transform 1 0 9510 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert90
timestamp 0
transform 1 0 5490 0 -1 11190
box -6 -8 86 268
use BUFX2  BUFX2_insert91
timestamp 0
transform -1 0 5090 0 1 10670
box -6 -8 86 268
use BUFX2  BUFX2_insert92
timestamp 0
transform -1 0 4930 0 -1 9630
box -6 -8 86 268
use BUFX2  BUFX2_insert93
timestamp 0
transform 1 0 5290 0 1 10150
box -6 -8 86 268
use BUFX2  BUFX2_insert94
timestamp 0
transform -1 0 11510 0 1 9630
box -6 -8 86 268
use BUFX2  BUFX2_insert95
timestamp 0
transform -1 0 11550 0 -1 10150
box -6 -8 86 268
use BUFX2  BUFX2_insert96
timestamp 0
transform -1 0 10270 0 1 11710
box -6 -8 86 268
use BUFX2  BUFX2_insert97
timestamp 0
transform 1 0 11590 0 1 11710
box -6 -8 86 268
use CLKBUF1  CLKBUF1_insert28
timestamp 0
transform -1 0 6330 0 -1 11710
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert29
timestamp 0
transform -1 0 2510 0 -1 6510
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert30
timestamp 0
transform 1 0 4670 0 -1 5470
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert31
timestamp 0
transform -1 0 3550 0 1 2870
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert32
timestamp 0
transform 1 0 7270 0 -1 8070
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert33
timestamp 0
transform 1 0 5850 0 -1 9110
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert34
timestamp 0
transform -1 0 2790 0 1 10670
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert35
timestamp 0
transform -1 0 5550 0 -1 12230
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert36
timestamp 0
transform -1 0 2670 0 1 3910
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert37
timestamp 0
transform 1 0 7510 0 -1 12230
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert38
timestamp 0
transform -1 0 4670 0 -1 9630
box -6 -8 206 268
use FILL  FILL181050x74250
timestamp 0
transform 1 0 12070 0 1 4950
box -6 -8 26 268
use FILL  FILL181350x35250
timestamp 0
transform 1 0 12090 0 1 2350
box -6 -8 26 268
use FILL  FILL181350x74250
timestamp 0
transform 1 0 12090 0 1 4950
box -6 -8 26 268
use FILL  FILL181350x109350
timestamp 0
transform -1 0 12110 0 -1 7550
box -6 -8 26 268
use FILL  FILL181350x117150
timestamp 0
transform -1 0 12110 0 -1 8070
box -6 -8 26 268
use FILL  FILL181350x140550
timestamp 0
transform -1 0 12110 0 -1 9630
box -6 -8 26 268
use FILL  FILL181650x35250
timestamp 0
transform 1 0 12110 0 1 2350
box -6 -8 26 268
use FILL  FILL181650x74250
timestamp 0
transform 1 0 12110 0 1 4950
box -6 -8 26 268
use FILL  FILL181650x109350
timestamp 0
transform -1 0 12130 0 -1 7550
box -6 -8 26 268
use FILL  FILL181650x117150
timestamp 0
transform -1 0 12130 0 -1 8070
box -6 -8 26 268
use FILL  FILL181650x140550
timestamp 0
transform -1 0 12130 0 -1 9630
box -6 -8 26 268
use FILL  FILL181650x148350
timestamp 0
transform -1 0 12130 0 -1 10150
box -6 -8 26 268
use FILL  FILL181950x7950
timestamp 0
transform -1 0 12150 0 -1 790
box -6 -8 26 268
use FILL  FILL181950x35250
timestamp 0
transform 1 0 12130 0 1 2350
box -6 -8 26 268
use FILL  FILL181950x74250
timestamp 0
transform 1 0 12130 0 1 4950
box -6 -8 26 268
use FILL  FILL181950x101550
timestamp 0
transform -1 0 12150 0 -1 7030
box -6 -8 26 268
use FILL  FILL181950x105450
timestamp 0
transform 1 0 12130 0 1 7030
box -6 -8 26 268
use FILL  FILL181950x109350
timestamp 0
transform -1 0 12150 0 -1 7550
box -6 -8 26 268
use FILL  FILL181950x117150
timestamp 0
transform -1 0 12150 0 -1 8070
box -6 -8 26 268
use FILL  FILL181950x140550
timestamp 0
transform -1 0 12150 0 -1 9630
box -6 -8 26 268
use FILL  FILL181950x148350
timestamp 0
transform -1 0 12150 0 -1 10150
box -6 -8 26 268
use FILL  FILL182250x7950
timestamp 0
transform -1 0 12170 0 -1 790
box -6 -8 26 268
use FILL  FILL182250x35250
timestamp 0
transform 1 0 12150 0 1 2350
box -6 -8 26 268
use FILL  FILL182250x74250
timestamp 0
transform 1 0 12150 0 1 4950
box -6 -8 26 268
use FILL  FILL182250x101550
timestamp 0
transform -1 0 12170 0 -1 7030
box -6 -8 26 268
use FILL  FILL182250x105450
timestamp 0
transform 1 0 12150 0 1 7030
box -6 -8 26 268
use FILL  FILL182250x109350
timestamp 0
transform -1 0 12170 0 -1 7550
box -6 -8 26 268
use FILL  FILL182250x117150
timestamp 0
transform -1 0 12170 0 -1 8070
box -6 -8 26 268
use FILL  FILL182250x140550
timestamp 0
transform -1 0 12170 0 -1 9630
box -6 -8 26 268
use FILL  FILL182250x148350
timestamp 0
transform -1 0 12170 0 -1 10150
box -6 -8 26 268
use FILL  FILL182250x163950
timestamp 0
transform -1 0 12170 0 -1 11190
box -6 -8 26 268
use FILL  FILL182550x7950
timestamp 0
transform -1 0 12190 0 -1 790
box -6 -8 26 268
use FILL  FILL182550x35250
timestamp 0
transform 1 0 12170 0 1 2350
box -6 -8 26 268
use FILL  FILL182550x74250
timestamp 0
transform 1 0 12170 0 1 4950
box -6 -8 26 268
use FILL  FILL182550x101550
timestamp 0
transform -1 0 12190 0 -1 7030
box -6 -8 26 268
use FILL  FILL182550x105450
timestamp 0
transform 1 0 12170 0 1 7030
box -6 -8 26 268
use FILL  FILL182550x109350
timestamp 0
transform -1 0 12190 0 -1 7550
box -6 -8 26 268
use FILL  FILL182550x117150
timestamp 0
transform -1 0 12190 0 -1 8070
box -6 -8 26 268
use FILL  FILL182550x140550
timestamp 0
transform -1 0 12190 0 -1 9630
box -6 -8 26 268
use FILL  FILL182550x148350
timestamp 0
transform -1 0 12190 0 -1 10150
box -6 -8 26 268
use FILL  FILL182550x163950
timestamp 0
transform -1 0 12190 0 -1 11190
box -6 -8 26 268
use FILL  FILL182850x7950
timestamp 0
transform -1 0 12210 0 -1 790
box -6 -8 26 268
use FILL  FILL182850x35250
timestamp 0
transform 1 0 12190 0 1 2350
box -6 -8 26 268
use FILL  FILL182850x74250
timestamp 0
transform 1 0 12190 0 1 4950
box -6 -8 26 268
use FILL  FILL182850x101550
timestamp 0
transform -1 0 12210 0 -1 7030
box -6 -8 26 268
use FILL  FILL182850x105450
timestamp 0
transform 1 0 12190 0 1 7030
box -6 -8 26 268
use FILL  FILL182850x109350
timestamp 0
transform -1 0 12210 0 -1 7550
box -6 -8 26 268
use FILL  FILL182850x117150
timestamp 0
transform -1 0 12210 0 -1 8070
box -6 -8 26 268
use FILL  FILL182850x140550
timestamp 0
transform -1 0 12210 0 -1 9630
box -6 -8 26 268
use FILL  FILL182850x148350
timestamp 0
transform -1 0 12210 0 -1 10150
box -6 -8 26 268
use FILL  FILL182850x163950
timestamp 0
transform -1 0 12210 0 -1 11190
box -6 -8 26 268
use FILL  FILL183150x7950
timestamp 0
transform -1 0 12230 0 -1 790
box -6 -8 26 268
use FILL  FILL183150x35250
timestamp 0
transform 1 0 12210 0 1 2350
box -6 -8 26 268
use FILL  FILL183150x74250
timestamp 0
transform 1 0 12210 0 1 4950
box -6 -8 26 268
use FILL  FILL183150x101550
timestamp 0
transform -1 0 12230 0 -1 7030
box -6 -8 26 268
use FILL  FILL183150x105450
timestamp 0
transform 1 0 12210 0 1 7030
box -6 -8 26 268
use FILL  FILL183150x109350
timestamp 0
transform -1 0 12230 0 -1 7550
box -6 -8 26 268
use FILL  FILL183150x117150
timestamp 0
transform -1 0 12230 0 -1 8070
box -6 -8 26 268
use FILL  FILL183150x140550
timestamp 0
transform -1 0 12230 0 -1 9630
box -6 -8 26 268
use FILL  FILL183150x148350
timestamp 0
transform -1 0 12230 0 -1 10150
box -6 -8 26 268
use FILL  FILL183150x163950
timestamp 0
transform -1 0 12230 0 -1 11190
box -6 -8 26 268
use FILL  FILL183150x167850
timestamp 0
transform 1 0 12210 0 1 11190
box -6 -8 26 268
use FILL  FILL183150x175650
timestamp 0
transform 1 0 12210 0 1 11710
box -6 -8 26 268
use FILL  FILL183450x150
timestamp 0
transform -1 0 12250 0 -1 270
box -6 -8 26 268
use FILL  FILL183450x7950
timestamp 0
transform -1 0 12250 0 -1 790
box -6 -8 26 268
use FILL  FILL183450x35250
timestamp 0
transform 1 0 12230 0 1 2350
box -6 -8 26 268
use FILL  FILL183450x74250
timestamp 0
transform 1 0 12230 0 1 4950
box -6 -8 26 268
use FILL  FILL183450x101550
timestamp 0
transform -1 0 12250 0 -1 7030
box -6 -8 26 268
use FILL  FILL183450x105450
timestamp 0
transform 1 0 12230 0 1 7030
box -6 -8 26 268
use FILL  FILL183450x109350
timestamp 0
transform -1 0 12250 0 -1 7550
box -6 -8 26 268
use FILL  FILL183450x117150
timestamp 0
transform -1 0 12250 0 -1 8070
box -6 -8 26 268
use FILL  FILL183450x140550
timestamp 0
transform -1 0 12250 0 -1 9630
box -6 -8 26 268
use FILL  FILL183450x148350
timestamp 0
transform -1 0 12250 0 -1 10150
box -6 -8 26 268
use FILL  FILL183450x163950
timestamp 0
transform -1 0 12250 0 -1 11190
box -6 -8 26 268
use FILL  FILL183450x167850
timestamp 0
transform 1 0 12230 0 1 11190
box -6 -8 26 268
use FILL  FILL183450x171750
timestamp 0
transform -1 0 12250 0 -1 11710
box -6 -8 26 268
use FILL  FILL183450x175650
timestamp 0
transform 1 0 12230 0 1 11710
box -6 -8 26 268
use FILL  FILL183750x150
timestamp 0
transform -1 0 12270 0 -1 270
box -6 -8 26 268
use FILL  FILL183750x7950
timestamp 0
transform -1 0 12270 0 -1 790
box -6 -8 26 268
use FILL  FILL183750x35250
timestamp 0
transform 1 0 12250 0 1 2350
box -6 -8 26 268
use FILL  FILL183750x70350
timestamp 0
transform -1 0 12270 0 -1 4950
box -6 -8 26 268
use FILL  FILL183750x74250
timestamp 0
transform 1 0 12250 0 1 4950
box -6 -8 26 268
use FILL  FILL183750x101550
timestamp 0
transform -1 0 12270 0 -1 7030
box -6 -8 26 268
use FILL  FILL183750x105450
timestamp 0
transform 1 0 12250 0 1 7030
box -6 -8 26 268
use FILL  FILL183750x109350
timestamp 0
transform -1 0 12270 0 -1 7550
box -6 -8 26 268
use FILL  FILL183750x117150
timestamp 0
transform -1 0 12270 0 -1 8070
box -6 -8 26 268
use FILL  FILL183750x140550
timestamp 0
transform -1 0 12270 0 -1 9630
box -6 -8 26 268
use FILL  FILL183750x148350
timestamp 0
transform -1 0 12270 0 -1 10150
box -6 -8 26 268
use FILL  FILL183750x160050
timestamp 0
transform 1 0 12250 0 1 10670
box -6 -8 26 268
use FILL  FILL183750x163950
timestamp 0
transform -1 0 12270 0 -1 11190
box -6 -8 26 268
use FILL  FILL183750x167850
timestamp 0
transform 1 0 12250 0 1 11190
box -6 -8 26 268
use FILL  FILL183750x171750
timestamp 0
transform -1 0 12270 0 -1 11710
box -6 -8 26 268
use FILL  FILL183750x175650
timestamp 0
transform 1 0 12250 0 1 11710
box -6 -8 26 268
use FILL  FILL184050x150
timestamp 0
transform -1 0 12290 0 -1 270
box -6 -8 26 268
use FILL  FILL184050x4050
timestamp 0
transform 1 0 12270 0 1 270
box -6 -8 26 268
use FILL  FILL184050x7950
timestamp 0
transform -1 0 12290 0 -1 790
box -6 -8 26 268
use FILL  FILL184050x27450
timestamp 0
transform 1 0 12270 0 1 1830
box -6 -8 26 268
use FILL  FILL184050x35250
timestamp 0
transform 1 0 12270 0 1 2350
box -6 -8 26 268
use FILL  FILL184050x54750
timestamp 0
transform -1 0 12290 0 -1 3910
box -6 -8 26 268
use FILL  FILL184050x70350
timestamp 0
transform -1 0 12290 0 -1 4950
box -6 -8 26 268
use FILL  FILL184050x74250
timestamp 0
transform 1 0 12270 0 1 4950
box -6 -8 26 268
use FILL  FILL184050x101550
timestamp 0
transform -1 0 12290 0 -1 7030
box -6 -8 26 268
use FILL  FILL184050x105450
timestamp 0
transform 1 0 12270 0 1 7030
box -6 -8 26 268
use FILL  FILL184050x109350
timestamp 0
transform -1 0 12290 0 -1 7550
box -6 -8 26 268
use FILL  FILL184050x117150
timestamp 0
transform -1 0 12290 0 -1 8070
box -6 -8 26 268
use FILL  FILL184050x121050
timestamp 0
transform 1 0 12270 0 1 8070
box -6 -8 26 268
use FILL  FILL184050x140550
timestamp 0
transform -1 0 12290 0 -1 9630
box -6 -8 26 268
use FILL  FILL184050x148350
timestamp 0
transform -1 0 12290 0 -1 10150
box -6 -8 26 268
use FILL  FILL184050x156150
timestamp 0
transform -1 0 12290 0 -1 10670
box -6 -8 26 268
use FILL  FILL184050x160050
timestamp 0
transform 1 0 12270 0 1 10670
box -6 -8 26 268
use FILL  FILL184050x163950
timestamp 0
transform -1 0 12290 0 -1 11190
box -6 -8 26 268
use FILL  FILL184050x167850
timestamp 0
transform 1 0 12270 0 1 11190
box -6 -8 26 268
use FILL  FILL184050x171750
timestamp 0
transform -1 0 12290 0 -1 11710
box -6 -8 26 268
use FILL  FILL184050x175650
timestamp 0
transform 1 0 12270 0 1 11710
box -6 -8 26 268
use FILL  FILL184350x150
timestamp 0
transform -1 0 12310 0 -1 270
box -6 -8 26 268
use FILL  FILL184350x4050
timestamp 0
transform 1 0 12290 0 1 270
box -6 -8 26 268
use FILL  FILL184350x7950
timestamp 0
transform -1 0 12310 0 -1 790
box -6 -8 26 268
use FILL  FILL184350x11850
timestamp 0
transform 1 0 12290 0 1 790
box -6 -8 26 268
use FILL  FILL184350x15750
timestamp 0
transform -1 0 12310 0 -1 1310
box -6 -8 26 268
use FILL  FILL184350x19650
timestamp 0
transform 1 0 12290 0 1 1310
box -6 -8 26 268
use FILL  FILL184350x23550
timestamp 0
transform -1 0 12310 0 -1 1830
box -6 -8 26 268
use FILL  FILL184350x27450
timestamp 0
transform 1 0 12290 0 1 1830
box -6 -8 26 268
use FILL  FILL184350x35250
timestamp 0
transform 1 0 12290 0 1 2350
box -6 -8 26 268
use FILL  FILL184350x39150
timestamp 0
transform -1 0 12310 0 -1 2870
box -6 -8 26 268
use FILL  FILL184350x43050
timestamp 0
transform 1 0 12290 0 1 2870
box -6 -8 26 268
use FILL  FILL184350x54750
timestamp 0
transform -1 0 12310 0 -1 3910
box -6 -8 26 268
use FILL  FILL184350x58650
timestamp 0
transform 1 0 12290 0 1 3910
box -6 -8 26 268
use FILL  FILL184350x62550
timestamp 0
transform -1 0 12310 0 -1 4430
box -6 -8 26 268
use FILL  FILL184350x70350
timestamp 0
transform -1 0 12310 0 -1 4950
box -6 -8 26 268
use FILL  FILL184350x74250
timestamp 0
transform 1 0 12290 0 1 4950
box -6 -8 26 268
use FILL  FILL184350x78150
timestamp 0
transform -1 0 12310 0 -1 5470
box -6 -8 26 268
use FILL  FILL184350x82050
timestamp 0
transform 1 0 12290 0 1 5470
box -6 -8 26 268
use FILL  FILL184350x85950
timestamp 0
transform -1 0 12310 0 -1 5990
box -6 -8 26 268
use FILL  FILL184350x97650
timestamp 0
transform 1 0 12290 0 1 6510
box -6 -8 26 268
use FILL  FILL184350x101550
timestamp 0
transform -1 0 12310 0 -1 7030
box -6 -8 26 268
use FILL  FILL184350x105450
timestamp 0
transform 1 0 12290 0 1 7030
box -6 -8 26 268
use FILL  FILL184350x109350
timestamp 0
transform -1 0 12310 0 -1 7550
box -6 -8 26 268
use FILL  FILL184350x113250
timestamp 0
transform 1 0 12290 0 1 7550
box -6 -8 26 268
use FILL  FILL184350x117150
timestamp 0
transform -1 0 12310 0 -1 8070
box -6 -8 26 268
use FILL  FILL184350x121050
timestamp 0
transform 1 0 12290 0 1 8070
box -6 -8 26 268
use FILL  FILL184350x124950
timestamp 0
transform -1 0 12310 0 -1 8590
box -6 -8 26 268
use FILL  FILL184350x136650
timestamp 0
transform 1 0 12290 0 1 9110
box -6 -8 26 268
use FILL  FILL184350x140550
timestamp 0
transform -1 0 12310 0 -1 9630
box -6 -8 26 268
use FILL  FILL184350x144450
timestamp 0
transform 1 0 12290 0 1 9630
box -6 -8 26 268
use FILL  FILL184350x148350
timestamp 0
transform -1 0 12310 0 -1 10150
box -6 -8 26 268
use FILL  FILL184350x152250
timestamp 0
transform 1 0 12290 0 1 10150
box -6 -8 26 268
use FILL  FILL184350x156150
timestamp 0
transform -1 0 12310 0 -1 10670
box -6 -8 26 268
use FILL  FILL184350x160050
timestamp 0
transform 1 0 12290 0 1 10670
box -6 -8 26 268
use FILL  FILL184350x163950
timestamp 0
transform -1 0 12310 0 -1 11190
box -6 -8 26 268
use FILL  FILL184350x167850
timestamp 0
transform 1 0 12290 0 1 11190
box -6 -8 26 268
use FILL  FILL184350x171750
timestamp 0
transform -1 0 12310 0 -1 11710
box -6 -8 26 268
use FILL  FILL184350x175650
timestamp 0
transform 1 0 12290 0 1 11710
box -6 -8 26 268
use FILL  FILL184350x179550
timestamp 0
transform -1 0 12310 0 -1 12230
box -6 -8 26 268
use FILL  FILL184650x150
timestamp 0
transform -1 0 12330 0 -1 270
box -6 -8 26 268
use FILL  FILL184650x4050
timestamp 0
transform 1 0 12310 0 1 270
box -6 -8 26 268
use FILL  FILL184650x7950
timestamp 0
transform -1 0 12330 0 -1 790
box -6 -8 26 268
use FILL  FILL184650x11850
timestamp 0
transform 1 0 12310 0 1 790
box -6 -8 26 268
use FILL  FILL184650x15750
timestamp 0
transform -1 0 12330 0 -1 1310
box -6 -8 26 268
use FILL  FILL184650x19650
timestamp 0
transform 1 0 12310 0 1 1310
box -6 -8 26 268
use FILL  FILL184650x23550
timestamp 0
transform -1 0 12330 0 -1 1830
box -6 -8 26 268
use FILL  FILL184650x27450
timestamp 0
transform 1 0 12310 0 1 1830
box -6 -8 26 268
use FILL  FILL184650x31350
timestamp 0
transform -1 0 12330 0 -1 2350
box -6 -8 26 268
use FILL  FILL184650x35250
timestamp 0
transform 1 0 12310 0 1 2350
box -6 -8 26 268
use FILL  FILL184650x39150
timestamp 0
transform -1 0 12330 0 -1 2870
box -6 -8 26 268
use FILL  FILL184650x43050
timestamp 0
transform 1 0 12310 0 1 2870
box -6 -8 26 268
use FILL  FILL184650x54750
timestamp 0
transform -1 0 12330 0 -1 3910
box -6 -8 26 268
use FILL  FILL184650x58650
timestamp 0
transform 1 0 12310 0 1 3910
box -6 -8 26 268
use FILL  FILL184650x62550
timestamp 0
transform -1 0 12330 0 -1 4430
box -6 -8 26 268
use FILL  FILL184650x70350
timestamp 0
transform -1 0 12330 0 -1 4950
box -6 -8 26 268
use FILL  FILL184650x74250
timestamp 0
transform 1 0 12310 0 1 4950
box -6 -8 26 268
use FILL  FILL184650x78150
timestamp 0
transform -1 0 12330 0 -1 5470
box -6 -8 26 268
use FILL  FILL184650x82050
timestamp 0
transform 1 0 12310 0 1 5470
box -6 -8 26 268
use FILL  FILL184650x85950
timestamp 0
transform -1 0 12330 0 -1 5990
box -6 -8 26 268
use FILL  FILL184650x89850
timestamp 0
transform 1 0 12310 0 1 5990
box -6 -8 26 268
use FILL  FILL184650x97650
timestamp 0
transform 1 0 12310 0 1 6510
box -6 -8 26 268
use FILL  FILL184650x101550
timestamp 0
transform -1 0 12330 0 -1 7030
box -6 -8 26 268
use FILL  FILL184650x105450
timestamp 0
transform 1 0 12310 0 1 7030
box -6 -8 26 268
use FILL  FILL184650x109350
timestamp 0
transform -1 0 12330 0 -1 7550
box -6 -8 26 268
use FILL  FILL184650x113250
timestamp 0
transform 1 0 12310 0 1 7550
box -6 -8 26 268
use FILL  FILL184650x117150
timestamp 0
transform -1 0 12330 0 -1 8070
box -6 -8 26 268
use FILL  FILL184650x121050
timestamp 0
transform 1 0 12310 0 1 8070
box -6 -8 26 268
use FILL  FILL184650x124950
timestamp 0
transform -1 0 12330 0 -1 8590
box -6 -8 26 268
use FILL  FILL184650x132750
timestamp 0
transform -1 0 12330 0 -1 9110
box -6 -8 26 268
use FILL  FILL184650x136650
timestamp 0
transform 1 0 12310 0 1 9110
box -6 -8 26 268
use FILL  FILL184650x140550
timestamp 0
transform -1 0 12330 0 -1 9630
box -6 -8 26 268
use FILL  FILL184650x144450
timestamp 0
transform 1 0 12310 0 1 9630
box -6 -8 26 268
use FILL  FILL184650x148350
timestamp 0
transform -1 0 12330 0 -1 10150
box -6 -8 26 268
use FILL  FILL184650x152250
timestamp 0
transform 1 0 12310 0 1 10150
box -6 -8 26 268
use FILL  FILL184650x156150
timestamp 0
transform -1 0 12330 0 -1 10670
box -6 -8 26 268
use FILL  FILL184650x160050
timestamp 0
transform 1 0 12310 0 1 10670
box -6 -8 26 268
use FILL  FILL184650x163950
timestamp 0
transform -1 0 12330 0 -1 11190
box -6 -8 26 268
use FILL  FILL184650x167850
timestamp 0
transform 1 0 12310 0 1 11190
box -6 -8 26 268
use FILL  FILL184650x171750
timestamp 0
transform -1 0 12330 0 -1 11710
box -6 -8 26 268
use FILL  FILL184650x175650
timestamp 0
transform 1 0 12310 0 1 11710
box -6 -8 26 268
use FILL  FILL184650x179550
timestamp 0
transform -1 0 12330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__1688_
timestamp 0
transform -1 0 830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1689_
timestamp 0
transform -1 0 290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1690_
timestamp 0
transform -1 0 550 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1691_
timestamp 0
transform 1 0 10 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1692_
timestamp 0
transform -1 0 270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1693_
timestamp 0
transform 1 0 510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1694_
timestamp 0
transform -1 0 5510 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1695_
timestamp 0
transform -1 0 290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1696_
timestamp 0
transform -1 0 290 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1697_
timestamp 0
transform -1 0 1410 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__1698_
timestamp 0
transform -1 0 3350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1699_
timestamp 0
transform 1 0 2790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1700_
timestamp 0
transform -1 0 3830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__1701_
timestamp 0
transform -1 0 530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1702_
timestamp 0
transform -1 0 530 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1703_
timestamp 0
transform 1 0 3170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1704_
timestamp 0
transform -1 0 310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1705_
timestamp 0
transform 1 0 10 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1706_
timestamp 0
transform -1 0 3790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1707_
timestamp 0
transform -1 0 550 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1708_
timestamp 0
transform 1 0 550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1709_
timestamp 0
transform 1 0 4070 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1710_
timestamp 0
transform -1 0 5550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1711_
timestamp 0
transform 1 0 5090 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1712_
timestamp 0
transform 1 0 7230 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 9610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1714_
timestamp 0
transform -1 0 9810 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1715_
timestamp 0
transform -1 0 8490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1716_
timestamp 0
transform 1 0 11250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1717_
timestamp 0
transform 1 0 11050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1718_
timestamp 0
transform 1 0 11870 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1719_
timestamp 0
transform -1 0 8750 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 10070 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1721_
timestamp 0
transform -1 0 10090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1722_
timestamp 0
transform -1 0 9850 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1723_
timestamp 0
transform 1 0 9950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1724_
timestamp 0
transform 1 0 9170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1725_
timestamp 0
transform 1 0 9010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1726_
timestamp 0
transform 1 0 10110 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1727_
timestamp 0
transform -1 0 8730 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1728_
timestamp 0
transform 1 0 11510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1729_
timestamp 0
transform 1 0 10110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1730_
timestamp 0
transform 1 0 8290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1731_
timestamp 0
transform 1 0 8530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1732_
timestamp 0
transform -1 0 7730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1733_
timestamp 0
transform 1 0 9670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1734_
timestamp 0
transform 1 0 7370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1735_
timestamp 0
transform 1 0 10810 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1736_
timestamp 0
transform -1 0 10610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1737_
timestamp 0
transform -1 0 10870 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1738_
timestamp 0
transform -1 0 10250 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1739_
timestamp 0
transform -1 0 10250 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1740_
timestamp 0
transform 1 0 10470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1741_
timestamp 0
transform -1 0 8370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1742_
timestamp 0
transform -1 0 8270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1743_
timestamp 0
transform -1 0 9830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1744_
timestamp 0
transform 1 0 9710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1745_
timestamp 0
transform -1 0 9410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1746_
timestamp 0
transform 1 0 11270 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1747_
timestamp 0
transform 1 0 10750 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1748_
timestamp 0
transform 1 0 7470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1749_
timestamp 0
transform 1 0 7890 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1750_
timestamp 0
transform -1 0 8010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1751_
timestamp 0
transform 1 0 7410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1752_
timestamp 0
transform -1 0 8830 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1753_
timestamp 0
transform 1 0 9690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1754_
timestamp 0
transform -1 0 8230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1755_
timestamp 0
transform -1 0 8810 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__1756_
timestamp 0
transform -1 0 11150 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1757_
timestamp 0
transform 1 0 11010 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1758_
timestamp 0
transform -1 0 9070 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1759_
timestamp 0
transform -1 0 7310 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__1760_
timestamp 0
transform 1 0 8810 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__1761_
timestamp 0
transform -1 0 9530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1762_
timestamp 0
transform 1 0 10550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1763_
timestamp 0
transform -1 0 8990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1764_
timestamp 0
transform 1 0 11250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1765_
timestamp 0
transform 1 0 8070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1766_
timestamp 0
transform 1 0 8450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1767_
timestamp 0
transform 1 0 9150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__1768_
timestamp 0
transform 1 0 8010 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__1769_
timestamp 0
transform 1 0 8530 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__1770_
timestamp 0
transform 1 0 8970 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__1771_
timestamp 0
transform 1 0 8930 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__1772_
timestamp 0
transform 1 0 8650 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__1773_
timestamp 0
transform 1 0 10730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1774_
timestamp 0
transform 1 0 10730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1775_
timestamp 0
transform 1 0 9970 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1776_
timestamp 0
transform -1 0 7970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1777_
timestamp 0
transform 1 0 8010 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1778_
timestamp 0
transform -1 0 7490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1779_
timestamp 0
transform 1 0 5630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1780_
timestamp 0
transform -1 0 4030 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1781_
timestamp 0
transform -1 0 10750 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1782_
timestamp 0
transform 1 0 8230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1783_
timestamp 0
transform 1 0 10470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1784_
timestamp 0
transform -1 0 9950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1785_
timestamp 0
transform -1 0 9710 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1786_
timestamp 0
transform 1 0 10130 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1787_
timestamp 0
transform -1 0 9070 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1788_
timestamp 0
transform -1 0 8490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1789_
timestamp 0
transform 1 0 9930 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1790_
timestamp 0
transform -1 0 9990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1791_
timestamp 0
transform -1 0 10070 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1792_
timestamp 0
transform -1 0 9610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1793_
timestamp 0
transform -1 0 9350 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1794_
timestamp 0
transform 1 0 9070 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1795_
timestamp 0
transform -1 0 8270 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1796_
timestamp 0
transform -1 0 8210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1797_
timestamp 0
transform 1 0 7050 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1798_
timestamp 0
transform 1 0 7310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1799_
timestamp 0
transform -1 0 9330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1800_
timestamp 0
transform 1 0 11210 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1801_
timestamp 0
transform 1 0 9230 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1802_
timestamp 0
transform -1 0 8890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1803_
timestamp 0
transform 1 0 10490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1804_
timestamp 0
transform -1 0 8510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1805_
timestamp 0
transform -1 0 8610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1806_
timestamp 0
transform 1 0 7550 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1807_
timestamp 0
transform -1 0 8010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1808_
timestamp 0
transform -1 0 8330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1809_
timestamp 0
transform 1 0 8550 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1810_
timestamp 0
transform 1 0 7950 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1811_
timestamp 0
transform -1 0 7690 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1812_
timestamp 0
transform -1 0 8330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1813_
timestamp 0
transform -1 0 8050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1814_
timestamp 0
transform -1 0 7790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1815_
timestamp 0
transform 1 0 7810 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1816_
timestamp 0
transform -1 0 3810 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1817_
timestamp 0
transform 1 0 1290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1818_
timestamp 0
transform -1 0 6110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1819_
timestamp 0
transform -1 0 870 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1820_
timestamp 0
transform 1 0 310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1821_
timestamp 0
transform 1 0 830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1822_
timestamp 0
transform -1 0 290 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1823_
timestamp 0
transform 1 0 1650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1824_
timestamp 0
transform 1 0 1230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1825_
timestamp 0
transform -1 0 1070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1826_
timestamp 0
transform -1 0 330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1827_
timestamp 0
transform 1 0 830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1828_
timestamp 0
transform -1 0 1430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1829_
timestamp 0
transform -1 0 570 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1830_
timestamp 0
transform -1 0 1370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1831_
timestamp 0
transform 1 0 1950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1832_
timestamp 0
transform -1 0 7950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1833_
timestamp 0
transform 1 0 9590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1834_
timestamp 0
transform 1 0 9170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1835_
timestamp 0
transform -1 0 7690 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1836_
timestamp 0
transform -1 0 6350 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1837_
timestamp 0
transform -1 0 7690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1838_
timestamp 0
transform -1 0 7130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1839_
timestamp 0
transform -1 0 6110 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1840_
timestamp 0
transform 1 0 8490 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1841_
timestamp 0
transform -1 0 8110 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1842_
timestamp 0
transform -1 0 6870 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1843_
timestamp 0
transform -1 0 6590 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1844_
timestamp 0
transform 1 0 9010 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1845_
timestamp 0
transform 1 0 9550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1846_
timestamp 0
transform -1 0 9150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1847_
timestamp 0
transform -1 0 8310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1848_
timestamp 0
transform 1 0 11150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1849_
timestamp 0
transform -1 0 11470 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1850_
timestamp 0
transform -1 0 10930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1851_
timestamp 0
transform 1 0 10290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1852_
timestamp 0
transform -1 0 10350 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1853_
timestamp 0
transform -1 0 10370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1854_
timestamp 0
transform -1 0 7350 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1855_
timestamp 0
transform 1 0 7330 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1856_
timestamp 0
transform 1 0 7610 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1857_
timestamp 0
transform -1 0 8750 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__1858_
timestamp 0
transform -1 0 9290 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1859_
timestamp 0
transform -1 0 8750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1860_
timestamp 0
transform 1 0 9010 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1861_
timestamp 0
transform 1 0 6750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1862_
timestamp 0
transform -1 0 8250 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__1863_
timestamp 0
transform 1 0 7610 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1864_
timestamp 0
transform -1 0 6250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1865_
timestamp 0
transform -1 0 7690 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__1866_
timestamp 0
transform -1 0 7150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1867_
timestamp 0
transform -1 0 7930 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1868_
timestamp 0
transform 1 0 7650 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1869_
timestamp 0
transform -1 0 5950 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__1870_
timestamp 0
transform 1 0 9290 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1871_
timestamp 0
transform 1 0 8770 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1872_
timestamp 0
transform -1 0 8510 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1873_
timestamp 0
transform -1 0 7710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1874_
timestamp 0
transform -1 0 7430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1875_
timestamp 0
transform -1 0 8230 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1876_
timestamp 0
transform -1 0 6870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1877_
timestamp 0
transform -1 0 5710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__1878_
timestamp 0
transform 1 0 6590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1879_
timestamp 0
transform -1 0 7390 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1880_
timestamp 0
transform 1 0 5910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__1881_
timestamp 0
transform 1 0 5910 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__1882_
timestamp 0
transform -1 0 4870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__1883_
timestamp 0
transform -1 0 7770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1884_
timestamp 0
transform -1 0 8010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1885_
timestamp 0
transform -1 0 8570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1886_
timestamp 0
transform 1 0 8410 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1887_
timestamp 0
transform -1 0 8390 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1888_
timestamp 0
transform 1 0 11530 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1889_
timestamp 0
transform -1 0 8390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1890_
timestamp 0
transform 1 0 9650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1891_
timestamp 0
transform 1 0 8810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1892_
timestamp 0
transform -1 0 8530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1893_
timestamp 0
transform 1 0 12050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1894_
timestamp 0
transform 1 0 12030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1895_
timestamp 0
transform 1 0 12050 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1896_
timestamp 0
transform -1 0 10670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1897_
timestamp 0
transform -1 0 9070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1898_
timestamp 0
transform 1 0 8950 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1899_
timestamp 0
transform 1 0 7390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1900_
timestamp 0
transform 1 0 9590 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1901_
timestamp 0
transform 1 0 7930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1902_
timestamp 0
transform -1 0 8150 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1903_
timestamp 0
transform 1 0 7870 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1904_
timestamp 0
transform 1 0 11790 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1905_
timestamp 0
transform 1 0 11550 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1906_
timestamp 0
transform -1 0 6430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1907_
timestamp 0
transform -1 0 6970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1908_
timestamp 0
transform -1 0 6890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1909_
timestamp 0
transform -1 0 6650 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1910_
timestamp 0
transform -1 0 6150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1911_
timestamp 0
transform 1 0 6730 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1912_
timestamp 0
transform 1 0 6190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1913_
timestamp 0
transform 1 0 6130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1914_
timestamp 0
transform 1 0 5630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1915_
timestamp 0
transform 1 0 5150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1916_
timestamp 0
transform 1 0 5150 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__1917_
timestamp 0
transform -1 0 3650 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__1918_
timestamp 0
transform 1 0 3530 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__1919_
timestamp 0
transform -1 0 3810 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__1920_
timestamp 0
transform -1 0 3530 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__1921_
timestamp 0
transform -1 0 1650 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__1922_
timestamp 0
transform 1 0 7450 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1923_
timestamp 0
transform 1 0 7710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1924_
timestamp 0
transform -1 0 6310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1925_
timestamp 0
transform -1 0 4550 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1926_
timestamp 0
transform -1 0 3910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1927_
timestamp 0
transform 1 0 1950 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__1928_
timestamp 0
transform -1 0 3110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__1929_
timestamp 0
transform 1 0 4490 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__1930_
timestamp 0
transform 1 0 3050 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__1931_
timestamp 0
transform -1 0 2830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__1932_
timestamp 0
transform -1 0 1430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1933_
timestamp 0
transform -1 0 8390 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1934_
timestamp 0
transform 1 0 3790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1935_
timestamp 0
transform -1 0 3810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1936_
timestamp 0
transform -1 0 2490 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1937_
timestamp 0
transform -1 0 1150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1938_
timestamp 0
transform -1 0 3510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1939_
timestamp 0
transform -1 0 4070 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1940_
timestamp 0
transform -1 0 3290 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1941_
timestamp 0
transform -1 0 3230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1942_
timestamp 0
transform -1 0 1730 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__1943_
timestamp 0
transform -1 0 3530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1944_
timestamp 0
transform -1 0 3630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1945_
timestamp 0
transform -1 0 2890 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1946_
timestamp 0
transform -1 0 1450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__1947_
timestamp 0
transform -1 0 4870 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__1948_
timestamp 0
transform 1 0 5070 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__1949_
timestamp 0
transform 1 0 5130 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__1950_
timestamp 0
transform -1 0 4870 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__1951_
timestamp 0
transform -1 0 1910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1952_
timestamp 0
transform 1 0 4030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1953_
timestamp 0
transform 1 0 3970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1954_
timestamp 0
transform 1 0 4110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1955_
timestamp 0
transform -1 0 1630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1956_
timestamp 0
transform -1 0 4250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__1957_
timestamp 0
transform 1 0 4830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__1958_
timestamp 0
transform -1 0 5110 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__1959_
timestamp 0
transform -1 0 4090 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__1960_
timestamp 0
transform -1 0 2250 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1961_
timestamp 0
transform 1 0 4070 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1962_
timestamp 0
transform 1 0 3830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1963_
timestamp 0
transform 1 0 3610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1964_
timestamp 0
transform 1 0 1950 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1965_
timestamp 0
transform 1 0 6330 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__1966_
timestamp 0
transform 1 0 6270 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1967_
timestamp 0
transform 1 0 7110 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1968_
timestamp 0
transform 1 0 6570 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1969_
timestamp 0
transform -1 0 3230 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__1970_
timestamp 0
transform 1 0 2770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1971_
timestamp 0
transform -1 0 4650 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1972_
timestamp 0
transform 1 0 3510 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1973_
timestamp 0
transform -1 0 3530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1974_
timestamp 0
transform -1 0 3030 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__1975_
timestamp 0
transform 1 0 2930 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__1976_
timestamp 0
transform -1 0 3030 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__1977_
timestamp 0
transform 1 0 4310 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__1978_
timestamp 0
transform 1 0 3010 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__1979_
timestamp 0
transform -1 0 2750 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__1980_
timestamp 0
transform -1 0 2270 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1981_
timestamp 0
transform 1 0 5890 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1982_
timestamp 0
transform 1 0 6010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1983_
timestamp 0
transform 1 0 6210 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1984_
timestamp 0
transform 1 0 5210 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1985_
timestamp 0
transform -1 0 4710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1986_
timestamp 0
transform 1 0 2490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__1987_
timestamp 0
transform -1 0 7210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1988_
timestamp 0
transform 1 0 7510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1989_
timestamp 0
transform 1 0 7570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1990_
timestamp 0
transform -1 0 7370 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1991_
timestamp 0
transform -1 0 7650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1992_
timestamp 0
transform 1 0 10390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1993_
timestamp 0
transform 1 0 9510 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__1994_
timestamp 0
transform -1 0 6190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__1995_
timestamp 0
transform 1 0 6570 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1996_
timestamp 0
transform -1 0 6710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1997_
timestamp 0
transform 1 0 6410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1998_
timestamp 0
transform 1 0 6410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__1999_
timestamp 0
transform 1 0 7470 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2000_
timestamp 0
transform 1 0 6390 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2001_
timestamp 0
transform 1 0 6630 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2002_
timestamp 0
transform 1 0 6590 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2003_
timestamp 0
transform 1 0 9470 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2004_
timestamp 0
transform 1 0 7410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2005_
timestamp 0
transform -1 0 7210 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2006_
timestamp 0
transform 1 0 6690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2007_
timestamp 0
transform 1 0 6530 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2008_
timestamp 0
transform -1 0 6170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2009_
timestamp 0
transform 1 0 6770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2010_
timestamp 0
transform -1 0 6990 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2011_
timestamp 0
transform 1 0 7230 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2012_
timestamp 0
transform -1 0 9370 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2013_
timestamp 0
transform 1 0 10510 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2014_
timestamp 0
transform -1 0 10770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2015_
timestamp 0
transform -1 0 6210 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2016_
timestamp 0
transform -1 0 7250 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2017_
timestamp 0
transform -1 0 7030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2018_
timestamp 0
transform 1 0 7270 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2019_
timestamp 0
transform 1 0 9350 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2020_
timestamp 0
transform -1 0 10250 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2021_
timestamp 0
transform -1 0 7290 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2022_
timestamp 0
transform 1 0 7530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2023_
timestamp 0
transform -1 0 7830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2024_
timestamp 0
transform 1 0 6050 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2025_
timestamp 0
transform -1 0 5930 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2026_
timestamp 0
transform 1 0 9630 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2027_
timestamp 0
transform 1 0 10170 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2028_
timestamp 0
transform -1 0 10170 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2029_
timestamp 0
transform -1 0 11050 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2030_
timestamp 0
transform 1 0 10670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2031_
timestamp 0
transform -1 0 10970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2032_
timestamp 0
transform 1 0 8890 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2033_
timestamp 0
transform 1 0 8350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2034_
timestamp 0
transform 1 0 8590 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2035_
timestamp 0
transform 1 0 8550 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2036_
timestamp 0
transform 1 0 11510 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2037_
timestamp 0
transform 1 0 11710 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2038_
timestamp 0
transform -1 0 7550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2039_
timestamp 0
transform -1 0 6630 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2040_
timestamp 0
transform 1 0 10890 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2041_
timestamp 0
transform 1 0 10970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2042_
timestamp 0
transform -1 0 10050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2043_
timestamp 0
transform -1 0 10430 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2044_
timestamp 0
transform -1 0 10950 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2045_
timestamp 0
transform -1 0 11290 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2046_
timestamp 0
transform 1 0 8770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2047_
timestamp 0
transform -1 0 9330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2048_
timestamp 0
transform 1 0 9130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2049_
timestamp 0
transform 1 0 9270 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2050_
timestamp 0
transform 1 0 9030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2051_
timestamp 0
transform 1 0 8730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2052_
timestamp 0
transform 1 0 9010 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2053_
timestamp 0
transform -1 0 9570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2054_
timestamp 0
transform 1 0 9790 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2055_
timestamp 0
transform -1 0 6430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2056_
timestamp 0
transform -1 0 6010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2057_
timestamp 0
transform 1 0 10210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2058_
timestamp 0
transform -1 0 9950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2059_
timestamp 0
transform -1 0 10090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2060_
timestamp 0
transform -1 0 9850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2061_
timestamp 0
transform 1 0 10030 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2062_
timestamp 0
transform -1 0 9110 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2063_
timestamp 0
transform 1 0 8190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2064_
timestamp 0
transform -1 0 7870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2065_
timestamp 0
transform -1 0 8690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2066_
timestamp 0
transform 1 0 8670 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2067_
timestamp 0
transform -1 0 7930 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2068_
timestamp 0
transform -1 0 8210 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2069_
timestamp 0
transform 1 0 7930 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2070_
timestamp 0
transform -1 0 8230 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2071_
timestamp 0
transform -1 0 8510 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2072_
timestamp 0
transform 1 0 8730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2073_
timestamp 0
transform 1 0 8990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2074_
timestamp 0
transform 1 0 9210 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2075_
timestamp 0
transform -1 0 9510 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2076_
timestamp 0
transform 1 0 11170 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2077_
timestamp 0
transform -1 0 11230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2078_
timestamp 0
transform -1 0 11030 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2079_
timestamp 0
transform 1 0 11170 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2080_
timestamp 0
transform -1 0 11010 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2081_
timestamp 0
transform 1 0 11010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2082_
timestamp 0
transform 1 0 10270 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2083_
timestamp 0
transform 1 0 9530 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2084_
timestamp 0
transform 1 0 11550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2085_
timestamp 0
transform 1 0 10970 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2086_
timestamp 0
transform 1 0 11470 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2087_
timestamp 0
transform 1 0 11490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2088_
timestamp 0
transform -1 0 12050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2089_
timestamp 0
transform 1 0 11770 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2090_
timestamp 0
transform 1 0 11950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2091_
timestamp 0
transform 1 0 9850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2092_
timestamp 0
transform 1 0 10470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2093_
timestamp 0
transform -1 0 11030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2094_
timestamp 0
transform 1 0 11270 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2095_
timestamp 0
transform -1 0 10930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2096_
timestamp 0
transform 1 0 11450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2097_
timestamp 0
transform -1 0 11790 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2098_
timestamp 0
transform -1 0 11970 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2099_
timestamp 0
transform -1 0 11270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2100_
timestamp 0
transform 1 0 11230 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2101_
timestamp 0
transform -1 0 11190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2102_
timestamp 0
transform -1 0 11570 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2103_
timestamp 0
transform 1 0 12050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2104_
timestamp 0
transform 1 0 12050 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2105_
timestamp 0
transform -1 0 11510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2106_
timestamp 0
transform -1 0 11490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2107_
timestamp 0
transform -1 0 12050 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2108_
timestamp 0
transform 1 0 8790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2109_
timestamp 0
transform 1 0 12050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2110_
timestamp 0
transform -1 0 12070 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2111_
timestamp 0
transform -1 0 12070 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2112_
timestamp 0
transform -1 0 11970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2113_
timestamp 0
transform 1 0 11730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2114_
timestamp 0
transform 1 0 10510 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2115_
timestamp 0
transform -1 0 9250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2116_
timestamp 0
transform -1 0 10130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2117_
timestamp 0
transform -1 0 10730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2118_
timestamp 0
transform -1 0 10690 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2119_
timestamp 0
transform 1 0 10590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2120_
timestamp 0
transform 1 0 10630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2121_
timestamp 0
transform -1 0 10370 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2122_
timestamp 0
transform 1 0 10570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2123_
timestamp 0
transform -1 0 8070 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2124_
timestamp 0
transform -1 0 7770 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2125_
timestamp 0
transform -1 0 10130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2126_
timestamp 0
transform 1 0 10530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2127_
timestamp 0
transform -1 0 6950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2128_
timestamp 0
transform -1 0 9090 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2129_
timestamp 0
transform 1 0 7210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2130_
timestamp 0
transform -1 0 10830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2131_
timestamp 0
transform -1 0 7870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2132_
timestamp 0
transform 1 0 6650 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2133_
timestamp 0
transform -1 0 6950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2134_
timestamp 0
transform -1 0 7210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2135_
timestamp 0
transform -1 0 11090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2136_
timestamp 0
transform -1 0 11250 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2137_
timestamp 0
transform 1 0 11230 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2138_
timestamp 0
transform 1 0 11310 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2139_
timestamp 0
transform -1 0 11230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2140_
timestamp 0
transform -1 0 10950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2141_
timestamp 0
transform 1 0 9870 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2142_
timestamp 0
transform 1 0 10670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2143_
timestamp 0
transform -1 0 10410 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2144_
timestamp 0
transform -1 0 10970 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2145_
timestamp 0
transform -1 0 4970 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2146_
timestamp 0
transform 1 0 9690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2147_
timestamp 0
transform 1 0 10250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2148_
timestamp 0
transform -1 0 6190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2149_
timestamp 0
transform 1 0 9970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2150_
timestamp 0
transform 1 0 8750 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2151_
timestamp 0
transform 1 0 7370 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2152_
timestamp 0
transform 1 0 8450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2153_
timestamp 0
transform 1 0 8710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2154_
timestamp 0
transform 1 0 8990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2155_
timestamp 0
transform -1 0 10070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2156_
timestamp 0
transform -1 0 10850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2157_
timestamp 0
transform 1 0 11090 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2158_
timestamp 0
transform -1 0 11670 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2159_
timestamp 0
transform -1 0 11790 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2160_
timestamp 0
transform -1 0 11330 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2161_
timestamp 0
transform 1 0 8070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2162_
timestamp 0
transform 1 0 8830 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2163_
timestamp 0
transform -1 0 9930 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2164_
timestamp 0
transform 1 0 9690 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2165_
timestamp 0
transform 1 0 10930 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2166_
timestamp 0
transform 1 0 10750 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2167_
timestamp 0
transform 1 0 9130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2168_
timestamp 0
transform 1 0 9950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2169_
timestamp 0
transform -1 0 8690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2170_
timestamp 0
transform -1 0 9110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2171_
timestamp 0
transform 1 0 10250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2172_
timestamp 0
transform 1 0 9670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2173_
timestamp 0
transform 1 0 9790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2174_
timestamp 0
transform -1 0 9430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2175_
timestamp 0
transform 1 0 9510 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2176_
timestamp 0
transform -1 0 9630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2177_
timestamp 0
transform -1 0 9330 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2178_
timestamp 0
transform -1 0 10930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2179_
timestamp 0
transform 1 0 9410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2180_
timestamp 0
transform 1 0 11770 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2181_
timestamp 0
transform 1 0 11750 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2182_
timestamp 0
transform 1 0 11830 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2183_
timestamp 0
transform -1 0 11210 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2184_
timestamp 0
transform 1 0 10950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2185_
timestamp 0
transform -1 0 10190 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2186_
timestamp 0
transform 1 0 10130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2187_
timestamp 0
transform -1 0 10530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2188_
timestamp 0
transform 1 0 11490 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2189_
timestamp 0
transform 1 0 9870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2190_
timestamp 0
transform 1 0 10430 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2191_
timestamp 0
transform 1 0 11050 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2192_
timestamp 0
transform 1 0 10990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2193_
timestamp 0
transform -1 0 10930 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2194_
timestamp 0
transform -1 0 10490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2195_
timestamp 0
transform -1 0 9370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2196_
timestamp 0
transform -1 0 11010 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2197_
timestamp 0
transform 1 0 11270 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2198_
timestamp 0
transform -1 0 9810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2199_
timestamp 0
transform -1 0 9870 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2200_
timestamp 0
transform -1 0 5730 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2201_
timestamp 0
transform 1 0 6250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2202_
timestamp 0
transform 1 0 5990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2203_
timestamp 0
transform 1 0 5990 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2204_
timestamp 0
transform 1 0 6730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2205_
timestamp 0
transform 1 0 7030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2206_
timestamp 0
transform 1 0 9370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2207_
timestamp 0
transform -1 0 9870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2208_
timestamp 0
transform -1 0 9290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2209_
timestamp 0
transform 1 0 10330 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2210_
timestamp 0
transform 1 0 10330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2211_
timestamp 0
transform 1 0 11170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2212_
timestamp 0
transform -1 0 11530 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2213_
timestamp 0
transform -1 0 11570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2214_
timestamp 0
transform 1 0 11530 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2215_
timestamp 0
transform 1 0 11630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2216_
timestamp 0
transform 1 0 12010 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2217_
timestamp 0
transform 1 0 11290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2218_
timestamp 0
transform 1 0 9570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2219_
timestamp 0
transform -1 0 9810 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2220_
timestamp 0
transform -1 0 9850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2221_
timestamp 0
transform -1 0 11790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2222_
timestamp 0
transform 1 0 11730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2223_
timestamp 0
transform -1 0 11770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2224_
timestamp 0
transform 1 0 11750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2225_
timestamp 0
transform 1 0 10850 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2226_
timestamp 0
transform 1 0 11810 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2227_
timestamp 0
transform 1 0 11530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2228_
timestamp 0
transform -1 0 11390 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2229_
timestamp 0
transform -1 0 10470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2230_
timestamp 0
transform -1 0 10190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2231_
timestamp 0
transform -1 0 8390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2232_
timestamp 0
transform 1 0 8630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2233_
timestamp 0
transform 1 0 9410 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2234_
timestamp 0
transform -1 0 9670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2235_
timestamp 0
transform -1 0 9790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2236_
timestamp 0
transform 1 0 7090 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2237_
timestamp 0
transform -1 0 6570 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2238_
timestamp 0
transform -1 0 6850 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2239_
timestamp 0
transform -1 0 8870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2240_
timestamp 0
transform -1 0 8590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2241_
timestamp 0
transform -1 0 8230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2242_
timestamp 0
transform -1 0 7410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2243_
timestamp 0
transform 1 0 7670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2244_
timestamp 0
transform 1 0 7950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2245_
timestamp 0
transform -1 0 7650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2246_
timestamp 0
transform 1 0 9030 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2247_
timestamp 0
transform -1 0 12030 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2248_
timestamp 0
transform 1 0 11230 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2249_
timestamp 0
transform -1 0 9390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2250_
timestamp 0
transform 1 0 10910 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2251_
timestamp 0
transform 1 0 10470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2252_
timestamp 0
transform 1 0 11210 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2253_
timestamp 0
transform -1 0 11810 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2254_
timestamp 0
transform 1 0 12050 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2255_
timestamp 0
transform -1 0 10410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2256_
timestamp 0
transform -1 0 10690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2257_
timestamp 0
transform 1 0 10930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2258_
timestamp 0
transform 1 0 12090 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2259_
timestamp 0
transform -1 0 11770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2260_
timestamp 0
transform 1 0 9950 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2261_
timestamp 0
transform 1 0 10210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2262_
timestamp 0
transform -1 0 10730 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2263_
timestamp 0
transform 1 0 11210 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2264_
timestamp 0
transform 1 0 12030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2265_
timestamp 0
transform -1 0 11290 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2266_
timestamp 0
transform -1 0 10650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2267_
timestamp 0
transform 1 0 11870 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2268_
timestamp 0
transform 1 0 12030 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2269_
timestamp 0
transform -1 0 11810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2270_
timestamp 0
transform 1 0 11230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2271_
timestamp 0
transform -1 0 11530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2272_
timestamp 0
transform 1 0 11790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2273_
timestamp 0
transform -1 0 12050 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2274_
timestamp 0
transform 1 0 9970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2275_
timestamp 0
transform -1 0 8130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2276_
timestamp 0
transform 1 0 8790 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2277_
timestamp 0
transform 1 0 9070 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2278_
timestamp 0
transform -1 0 9150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2279_
timestamp 0
transform 1 0 8950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2280_
timestamp 0
transform 1 0 10110 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2281_
timestamp 0
transform 1 0 11990 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2282_
timestamp 0
transform 1 0 12050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2283_
timestamp 0
transform -1 0 10930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2284_
timestamp 0
transform 1 0 12010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2285_
timestamp 0
transform 1 0 12010 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2286_
timestamp 0
transform -1 0 11790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2287_
timestamp 0
transform 1 0 11730 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2288_
timestamp 0
transform -1 0 10890 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2289_
timestamp 0
transform -1 0 10670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2290_
timestamp 0
transform -1 0 10850 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2291_
timestamp 0
transform 1 0 11210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2292_
timestamp 0
transform 1 0 10350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2293_
timestamp 0
transform 1 0 10630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2294_
timestamp 0
transform 1 0 10950 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2295_
timestamp 0
transform 1 0 10830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2296_
timestamp 0
transform 1 0 11090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2297_
timestamp 0
transform 1 0 11750 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2298_
timestamp 0
transform -1 0 11850 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2299_
timestamp 0
transform -1 0 10410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2300_
timestamp 0
transform 1 0 10110 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2301_
timestamp 0
transform 1 0 11730 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2302_
timestamp 0
transform 1 0 11670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2303_
timestamp 0
transform -1 0 11650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2304_
timestamp 0
transform 1 0 11790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2305_
timestamp 0
transform 1 0 10670 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2306_
timestamp 0
transform -1 0 11530 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2307_
timestamp 0
transform 1 0 11230 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2308_
timestamp 0
transform 1 0 12010 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2309_
timestamp 0
transform -1 0 11570 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2310_
timestamp 0
transform -1 0 11510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2311_
timestamp 0
transform 1 0 11490 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2312_
timestamp 0
transform 1 0 11550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2313_
timestamp 0
transform 1 0 11830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2314_
timestamp 0
transform -1 0 11150 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2315_
timestamp 0
transform 1 0 12010 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2316_
timestamp 0
transform 1 0 11410 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2317_
timestamp 0
transform -1 0 11910 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2318_
timestamp 0
transform 1 0 11450 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2319_
timestamp 0
transform 1 0 11090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2320_
timestamp 0
transform 1 0 11510 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2321_
timestamp 0
transform 1 0 11370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2322_
timestamp 0
transform -1 0 11230 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2323_
timestamp 0
transform -1 0 11470 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2324_
timestamp 0
transform 1 0 11710 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2325_
timestamp 0
transform -1 0 12090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2326_
timestamp 0
transform 1 0 12010 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2327_
timestamp 0
transform 1 0 11370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2328_
timestamp 0
transform 1 0 10950 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2329_
timestamp 0
transform 1 0 8470 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2330_
timestamp 0
transform -1 0 10150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2331_
timestamp 0
transform -1 0 9590 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2332_
timestamp 0
transform -1 0 11810 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2333_
timestamp 0
transform -1 0 10690 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2334_
timestamp 0
transform 1 0 10410 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2335_
timestamp 0
transform 1 0 10390 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2336_
timestamp 0
transform 1 0 10570 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2337_
timestamp 0
transform -1 0 10690 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2338_
timestamp 0
transform -1 0 10610 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2339_
timestamp 0
transform -1 0 9530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2340_
timestamp 0
transform -1 0 9810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2341_
timestamp 0
transform 1 0 9510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2342_
timestamp 0
transform -1 0 10390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2343_
timestamp 0
transform -1 0 10330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2344_
timestamp 0
transform -1 0 10570 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2345_
timestamp 0
transform 1 0 11690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2346_
timestamp 0
transform 1 0 11430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2347_
timestamp 0
transform -1 0 8770 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2348_
timestamp 0
transform -1 0 9870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2349_
timestamp 0
transform -1 0 11530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2350_
timestamp 0
transform -1 0 11250 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2351_
timestamp 0
transform -1 0 10310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2352_
timestamp 0
transform -1 0 10070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2353_
timestamp 0
transform -1 0 9370 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2354_
timestamp 0
transform 1 0 7770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2355_
timestamp 0
transform -1 0 6850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2356_
timestamp 0
transform -1 0 6790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2357_
timestamp 0
transform -1 0 7450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2358_
timestamp 0
transform -1 0 7030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2359_
timestamp 0
transform 1 0 7250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2360_
timestamp 0
transform -1 0 7930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2361_
timestamp 0
transform -1 0 6990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2362_
timestamp 0
transform 1 0 8710 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2363_
timestamp 0
transform -1 0 7390 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2364_
timestamp 0
transform 1 0 7130 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2365_
timestamp 0
transform 1 0 6850 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2366_
timestamp 0
transform 1 0 6330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2367_
timestamp 0
transform -1 0 7170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2368_
timestamp 0
transform 1 0 6570 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2369_
timestamp 0
transform 1 0 6950 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2370_
timestamp 0
transform -1 0 7210 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2371_
timestamp 0
transform 1 0 7150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2372_
timestamp 0
transform -1 0 6730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2373_
timestamp 0
transform 1 0 6670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2374_
timestamp 0
transform 1 0 8170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2375_
timestamp 0
transform 1 0 8230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2376_
timestamp 0
transform -1 0 6670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2377_
timestamp 0
transform 1 0 5370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2378_
timestamp 0
transform -1 0 3690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2379_
timestamp 0
transform -1 0 7950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2380_
timestamp 0
transform -1 0 5590 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2381_
timestamp 0
transform -1 0 5870 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2382_
timestamp 0
transform -1 0 5730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2383_
timestamp 0
transform 1 0 4650 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2384_
timestamp 0
transform 1 0 4570 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2385_
timestamp 0
transform 1 0 4810 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2386_
timestamp 0
transform 1 0 5090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2387_
timestamp 0
transform 1 0 1610 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2388_
timestamp 0
transform 1 0 1550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2389_
timestamp 0
transform 1 0 5130 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2390_
timestamp 0
transform 1 0 2410 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2391_
timestamp 0
transform -1 0 2210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2392_
timestamp 0
transform -1 0 1930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2393_
timestamp 0
transform -1 0 2490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2394_
timestamp 0
transform -1 0 2910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2395_
timestamp 0
transform 1 0 4310 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2396_
timestamp 0
transform 1 0 2950 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2397_
timestamp 0
transform -1 0 3030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2398_
timestamp 0
transform -1 0 2750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2399_
timestamp 0
transform 1 0 1850 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2400_
timestamp 0
transform -1 0 1290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2401_
timestamp 0
transform -1 0 2770 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2402_
timestamp 0
transform 1 0 2510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2403_
timestamp 0
transform -1 0 2150 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2404_
timestamp 0
transform -1 0 1590 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2405_
timestamp 0
transform -1 0 1450 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2406_
timestamp 0
transform 1 0 5830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2407_
timestamp 0
transform -1 0 4190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2408_
timestamp 0
transform -1 0 5550 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2409_
timestamp 0
transform -1 0 6370 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2410_
timestamp 0
transform -1 0 4150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2411_
timestamp 0
transform -1 0 3910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2412_
timestamp 0
transform -1 0 1170 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2413_
timestamp 0
transform -1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2414_
timestamp 0
transform 1 0 2970 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2415_
timestamp 0
transform -1 0 2710 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2416_
timestamp 0
transform 1 0 1670 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2417_
timestamp 0
transform -1 0 2170 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2418_
timestamp 0
transform -1 0 2050 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2419_
timestamp 0
transform -1 0 3370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2420_
timestamp 0
transform 1 0 2790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2421_
timestamp 0
transform -1 0 2710 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2422_
timestamp 0
transform -1 0 1890 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2423_
timestamp 0
transform -1 0 3590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2424_
timestamp 0
transform -1 0 3430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2425_
timestamp 0
transform -1 0 3310 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2426_
timestamp 0
transform 1 0 3070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2427_
timestamp 0
transform 1 0 3230 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2428_
timestamp 0
transform -1 0 3310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2429_
timestamp 0
transform -1 0 5030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2430_
timestamp 0
transform -1 0 7730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2431_
timestamp 0
transform -1 0 5290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2432_
timestamp 0
transform -1 0 9410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2433_
timestamp 0
transform 1 0 11510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2434_
timestamp 0
transform 1 0 10690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2435_
timestamp 0
transform -1 0 7170 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2436_
timestamp 0
transform -1 0 6850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2437_
timestamp 0
transform -1 0 9530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2438_
timestamp 0
transform -1 0 9270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2439_
timestamp 0
transform -1 0 6050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2440_
timestamp 0
transform 1 0 7670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2441_
timestamp 0
transform -1 0 7510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2442_
timestamp 0
transform 1 0 10210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2443_
timestamp 0
transform -1 0 7110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2444_
timestamp 0
transform -1 0 7110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2445_
timestamp 0
transform 1 0 5210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2446_
timestamp 0
transform 1 0 6330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2447_
timestamp 0
transform -1 0 4710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2448_
timestamp 0
transform -1 0 6310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2449_
timestamp 0
transform -1 0 6930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2450_
timestamp 0
transform 1 0 4070 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2451_
timestamp 0
transform -1 0 3950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2452_
timestamp 0
transform 1 0 4590 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2453_
timestamp 0
transform 1 0 8450 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2454_
timestamp 0
transform 1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2455_
timestamp 0
transform 1 0 4330 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2456_
timestamp 0
transform -1 0 4190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2457_
timestamp 0
transform -1 0 4450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2458_
timestamp 0
transform -1 0 4810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2459_
timestamp 0
transform 1 0 4950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2460_
timestamp 0
transform 1 0 4830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2461_
timestamp 0
transform 1 0 5110 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2462_
timestamp 0
transform 1 0 5250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2463_
timestamp 0
transform 1 0 6190 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2464_
timestamp 0
transform -1 0 3130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2465_
timestamp 0
transform -1 0 2850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2466_
timestamp 0
transform -1 0 2850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2467_
timestamp 0
transform 1 0 1990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2468_
timestamp 0
transform -1 0 1550 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2469_
timestamp 0
transform 1 0 510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2470_
timestamp 0
transform -1 0 2610 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2471_
timestamp 0
transform -1 0 2630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2472_
timestamp 0
transform -1 0 2330 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2473_
timestamp 0
transform 1 0 1830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2474_
timestamp 0
transform -1 0 1350 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2475_
timestamp 0
transform -1 0 290 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2476_
timestamp 0
transform -1 0 3710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2477_
timestamp 0
transform -1 0 4950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2478_
timestamp 0
transform 1 0 3810 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2479_
timestamp 0
transform -1 0 3450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2480_
timestamp 0
transform 1 0 1690 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2481_
timestamp 0
transform -1 0 3250 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2482_
timestamp 0
transform 1 0 3530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2483_
timestamp 0
transform 1 0 2950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2484_
timestamp 0
transform 1 0 2670 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2485_
timestamp 0
transform -1 0 290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2486_
timestamp 0
transform -1 0 2570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2487_
timestamp 0
transform 1 0 2290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2488_
timestamp 0
transform -1 0 2290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2489_
timestamp 0
transform -1 0 1730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2490_
timestamp 0
transform -1 0 1290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2491_
timestamp 0
transform -1 0 290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2492_
timestamp 0
transform 1 0 4510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2493_
timestamp 0
transform 1 0 3510 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2494_
timestamp 0
transform 1 0 6090 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2495_
timestamp 0
transform 1 0 3750 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2496_
timestamp 0
transform 1 0 4050 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2497_
timestamp 0
transform -1 0 3970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2498_
timestamp 0
transform 1 0 3430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2499_
timestamp 0
transform 1 0 3690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2500_
timestamp 0
transform -1 0 290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2501_
timestamp 0
transform -1 0 3290 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2502_
timestamp 0
transform -1 0 2930 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2503_
timestamp 0
transform -1 0 3410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__2504_
timestamp 0
transform -1 0 3170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__2505_
timestamp 0
transform 1 0 2610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2506_
timestamp 0
transform -1 0 2430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__2507_
timestamp 0
transform 1 0 550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2508_
timestamp 0
transform 1 0 3050 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2509_
timestamp 0
transform 1 0 2590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2510_
timestamp 0
transform -1 0 3150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2511_
timestamp 0
transform 1 0 3230 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__2512_
timestamp 0
transform 1 0 3070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2513_
timestamp 0
transform -1 0 2330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2514_
timestamp 0
transform 1 0 2030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2515_
timestamp 0
transform -1 0 2050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2516_
timestamp 0
transform -1 0 290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__2517_
timestamp 0
transform -1 0 2130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2518_
timestamp 0
transform 1 0 5230 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2519_
timestamp 0
transform -1 0 5770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2520_
timestamp 0
transform -1 0 5870 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2521_
timestamp 0
transform 1 0 5570 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2522_
timestamp 0
transform -1 0 5570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2523_
timestamp 0
transform -1 0 5490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2524_
timestamp 0
transform -1 0 5430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2525_
timestamp 0
transform -1 0 2650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2526_
timestamp 0
transform 1 0 6050 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2527_
timestamp 0
transform 1 0 6450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2528_
timestamp 0
transform 1 0 6430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2529_
timestamp 0
transform 1 0 6030 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2530_
timestamp 0
transform 1 0 5490 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2531_
timestamp 0
transform 1 0 2850 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2532_
timestamp 0
transform 1 0 4130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2533_
timestamp 0
transform 1 0 5070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2534_
timestamp 0
transform 1 0 4790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2535_
timestamp 0
transform -1 0 4530 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2536_
timestamp 0
transform 1 0 3370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2537_
timestamp 0
transform 1 0 2010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2538_
timestamp 0
transform 1 0 4410 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2539_
timestamp 0
transform 1 0 3790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2540_
timestamp 0
transform 1 0 4130 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2541_
timestamp 0
transform -1 0 4110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2542_
timestamp 0
transform -1 0 3630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2543_
timestamp 0
transform 1 0 3390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2544_
timestamp 0
transform 1 0 4110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2545_
timestamp 0
transform 1 0 4370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2546_
timestamp 0
transform 1 0 4730 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2547_
timestamp 0
transform -1 0 4670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2548_
timestamp 0
transform -1 0 4390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2549_
timestamp 0
transform 1 0 4610 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2550_
timestamp 0
transform 1 0 4610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2551_
timestamp 0
transform 1 0 5130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2552_
timestamp 0
transform 1 0 5370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2553_
timestamp 0
transform 1 0 2270 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2554_
timestamp 0
transform 1 0 4410 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2555_
timestamp 0
transform -1 0 4590 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2556_
timestamp 0
transform -1 0 4830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2557_
timestamp 0
transform 1 0 4530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2558_
timestamp 0
transform 1 0 4610 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2559_
timestamp 0
transform 1 0 4330 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2560_
timestamp 0
transform 1 0 3830 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2561_
timestamp 0
transform 1 0 3530 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2562_
timestamp 0
transform 1 0 2150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2563_
timestamp 0
transform -1 0 4370 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2564_
timestamp 0
transform 1 0 4290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2565_
timestamp 0
transform -1 0 3770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2566_
timestamp 0
transform 1 0 2370 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2567_
timestamp 0
transform 1 0 3850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2568_
timestamp 0
transform -1 0 5650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2569_
timestamp 0
transform -1 0 5790 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2570_
timestamp 0
transform 1 0 5870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2571_
timestamp 0
transform 1 0 5870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2572_
timestamp 0
transform 1 0 5730 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2573_
timestamp 0
transform 1 0 5650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2574_
timestamp 0
transform 1 0 5630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2575_
timestamp 0
transform -1 0 4670 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2576_
timestamp 0
transform -1 0 4150 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2577_
timestamp 0
transform -1 0 4410 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2578_
timestamp 0
transform 1 0 6910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2579_
timestamp 0
transform 1 0 6930 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2580_
timestamp 0
transform 1 0 7930 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2581_
timestamp 0
transform -1 0 8790 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2582_
timestamp 0
transform 1 0 6830 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2583_
timestamp 0
transform -1 0 6830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2584_
timestamp 0
transform 1 0 7250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2585_
timestamp 0
transform 1 0 7290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2586_
timestamp 0
transform -1 0 8370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2587_
timestamp 0
transform -1 0 6710 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2588_
timestamp 0
transform -1 0 5750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2589_
timestamp 0
transform 1 0 7370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2590_
timestamp 0
transform -1 0 6150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2591_
timestamp 0
transform 1 0 6390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2592_
timestamp 0
transform -1 0 4370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2593_
timestamp 0
transform 1 0 4890 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2594_
timestamp 0
transform -1 0 8470 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2595_
timestamp 0
transform -1 0 5190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2596_
timestamp 0
transform 1 0 5190 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2597_
timestamp 0
transform 1 0 5370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2598_
timestamp 0
transform -1 0 5110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2599_
timestamp 0
transform -1 0 4910 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2600_
timestamp 0
transform -1 0 4910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2601_
timestamp 0
transform -1 0 5170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2602_
timestamp 0
transform -1 0 8110 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2603_
timestamp 0
transform -1 0 6550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2604_
timestamp 0
transform -1 0 6310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2605_
timestamp 0
transform 1 0 5990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2606_
timestamp 0
transform -1 0 5490 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2607_
timestamp 0
transform 1 0 5650 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2608_
timestamp 0
transform 1 0 5470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2609_
timestamp 0
transform -1 0 5450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2610_
timestamp 0
transform 1 0 4830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2611_
timestamp 0
transform -1 0 5090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2612_
timestamp 0
transform -1 0 5350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2613_
timestamp 0
transform -1 0 1170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2614_
timestamp 0
transform 1 0 2150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2615_
timestamp 0
transform -1 0 2430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2616_
timestamp 0
transform -1 0 2410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2617_
timestamp 0
transform 1 0 1390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2618_
timestamp 0
transform 1 0 810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2619_
timestamp 0
transform -1 0 310 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2620_
timestamp 0
transform -1 0 550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2621_
timestamp 0
transform 1 0 870 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2622_
timestamp 0
transform 1 0 310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2623_
timestamp 0
transform 1 0 2690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2624_
timestamp 0
transform 1 0 1890 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2625_
timestamp 0
transform -1 0 2150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2626_
timestamp 0
transform -1 0 1870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2627_
timestamp 0
transform 1 0 10 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2628_
timestamp 0
transform 1 0 10 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2629_
timestamp 0
transform -1 0 270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2630_
timestamp 0
transform 1 0 10 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2631_
timestamp 0
transform 1 0 4950 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2632_
timestamp 0
transform 1 0 2190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2633_
timestamp 0
transform -1 0 2490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2634_
timestamp 0
transform -1 0 30 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2635_
timestamp 0
transform 1 0 10 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2636_
timestamp 0
transform 1 0 550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2637_
timestamp 0
transform 1 0 890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2638_
timestamp 0
transform 1 0 310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2639_
timestamp 0
transform -1 0 630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2640_
timestamp 0
transform -1 0 30 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2641_
timestamp 0
transform -1 0 30 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2642_
timestamp 0
transform 1 0 1270 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2643_
timestamp 0
transform -1 0 1810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2644_
timestamp 0
transform 1 0 2210 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2645_
timestamp 0
transform -1 0 1950 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2646_
timestamp 0
transform -1 0 1150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2647_
timestamp 0
transform 1 0 10 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2648_
timestamp 0
transform 1 0 510 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__2649_
timestamp 0
transform 1 0 10 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2650_
timestamp 0
transform -1 0 3610 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2651_
timestamp 0
transform -1 0 3330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2652_
timestamp 0
transform 1 0 550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2653_
timestamp 0
transform 1 0 270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2654_
timestamp 0
transform 1 0 1150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2655_
timestamp 0
transform 1 0 590 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2656_
timestamp 0
transform -1 0 870 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2657_
timestamp 0
transform 1 0 10 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2658_
timestamp 0
transform 1 0 10 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2659_
timestamp 0
transform -1 0 310 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2660_
timestamp 0
transform 1 0 250 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2661_
timestamp 0
transform -1 0 2570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__2662_
timestamp 0
transform -1 0 2510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2663_
timestamp 0
transform -1 0 1930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2664_
timestamp 0
transform 1 0 830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2665_
timestamp 0
transform -1 0 790 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2666_
timestamp 0
transform -1 0 310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2667_
timestamp 0
transform -1 0 530 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2668_
timestamp 0
transform 1 0 1030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2669_
timestamp 0
transform -1 0 2790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2670_
timestamp 0
transform -1 0 2910 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2671_
timestamp 0
transform 1 0 1070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2672_
timestamp 0
transform -1 0 570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2673_
timestamp 0
transform -1 0 530 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2674_
timestamp 0
transform 1 0 790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2675_
timestamp 0
transform 1 0 770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2676_
timestamp 0
transform -1 0 1070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2677_
timestamp 0
transform 1 0 6410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__2678_
timestamp 0
transform -1 0 6330 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2679_
timestamp 0
transform 1 0 6950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2680_
timestamp 0
transform -1 0 6750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2681_
timestamp 0
transform 1 0 7010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2682_
timestamp 0
transform -1 0 6730 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2683_
timestamp 0
transform -1 0 1850 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2684_
timestamp 0
transform -1 0 1670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__2685_
timestamp 0
transform 1 0 1590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2686_
timestamp 0
transform 1 0 1590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2687_
timestamp 0
transform 1 0 1330 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2688_
timestamp 0
transform -1 0 770 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2689_
timestamp 0
transform -1 0 750 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2690_
timestamp 0
transform 1 0 7250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2691_
timestamp 0
transform -1 0 7090 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2692_
timestamp 0
transform -1 0 5030 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2693_
timestamp 0
transform -1 0 2990 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2694_
timestamp 0
transform -1 0 1290 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2695_
timestamp 0
transform -1 0 1570 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2696_
timestamp 0
transform -1 0 1290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2697_
timestamp 0
transform 1 0 1870 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2698_
timestamp 0
transform -1 0 510 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2699_
timestamp 0
transform 1 0 6270 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2700_
timestamp 0
transform -1 0 6990 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2701_
timestamp 0
transform 1 0 7570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2702_
timestamp 0
transform 1 0 7270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2703_
timestamp 0
transform 1 0 7430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2704_
timestamp 0
transform -1 0 6630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2705_
timestamp 0
transform 1 0 1550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2706_
timestamp 0
transform 1 0 990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2707_
timestamp 0
transform 1 0 2690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2708_
timestamp 0
transform 1 0 2370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2709_
timestamp 0
transform -1 0 1050 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2710_
timestamp 0
transform -1 0 830 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2711_
timestamp 0
transform -1 0 1110 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2712_
timestamp 0
transform 1 0 2850 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2713_
timestamp 0
transform -1 0 4250 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2714_
timestamp 0
transform -1 0 4670 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2715_
timestamp 0
transform 1 0 3510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2716_
timestamp 0
transform -1 0 4270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2717_
timestamp 0
transform -1 0 5830 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__2718_
timestamp 0
transform -1 0 4070 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2719_
timestamp 0
transform 1 0 3670 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2720_
timestamp 0
transform -1 0 3970 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2721_
timestamp 0
transform -1 0 2130 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2722_
timestamp 0
transform 1 0 2250 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2723_
timestamp 0
transform 1 0 2550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2724_
timestamp 0
transform -1 0 790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2725_
timestamp 0
transform -1 0 5390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2726_
timestamp 0
transform -1 0 6570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2727_
timestamp 0
transform 1 0 3830 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2728_
timestamp 0
transform 1 0 3550 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2729_
timestamp 0
transform -1 0 3510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2730_
timestamp 0
transform 1 0 3110 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2731_
timestamp 0
transform 1 0 1970 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2732_
timestamp 0
transform -1 0 1850 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2733_
timestamp 0
transform 1 0 1390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2734_
timestamp 0
transform -1 0 1690 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2735_
timestamp 0
transform -1 0 3850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2736_
timestamp 0
transform -1 0 3990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2737_
timestamp 0
transform -1 0 4070 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2738_
timestamp 0
transform -1 0 3770 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2739_
timestamp 0
transform -1 0 3210 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2740_
timestamp 0
transform -1 0 3290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2741_
timestamp 0
transform -1 0 1050 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2742_
timestamp 0
transform 1 0 1350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2743_
timestamp 0
transform 1 0 1290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2744_
timestamp 0
transform 1 0 1830 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2745_
timestamp 0
transform 1 0 490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2746_
timestamp 0
transform 1 0 3550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2747_
timestamp 0
transform 1 0 4670 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__2748_
timestamp 0
transform 1 0 4330 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2749_
timestamp 0
transform -1 0 3490 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2750_
timestamp 0
transform -1 0 2930 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2751_
timestamp 0
transform 1 0 2770 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2752_
timestamp 0
transform 1 0 1070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2753_
timestamp 0
transform 1 0 570 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2754_
timestamp 0
transform -1 0 510 0 1 790
box -6 -8 26 268
use FILL  FILL_0__2755_
timestamp 0
transform -1 0 3030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2756_
timestamp 0
transform -1 0 2470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2757_
timestamp 0
transform 1 0 2710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2758_
timestamp 0
transform 1 0 2190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2759_
timestamp 0
transform -1 0 4270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2760_
timestamp 0
transform 1 0 3710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2761_
timestamp 0
transform 1 0 4050 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2762_
timestamp 0
transform -1 0 3790 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2763_
timestamp 0
transform -1 0 2030 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2764_
timestamp 0
transform -1 0 1750 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2765_
timestamp 0
transform -1 0 1670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2766_
timestamp 0
transform -1 0 1930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__2767_
timestamp 0
transform -1 0 1450 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__2768_
timestamp 0
transform 1 0 2110 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2769_
timestamp 0
transform 1 0 1550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__2770_
timestamp 0
transform 1 0 5910 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2771_
timestamp 0
transform 1 0 6450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2772_
timestamp 0
transform 1 0 4890 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__2773_
timestamp 0
transform 1 0 4090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2774_
timestamp 0
transform 1 0 2250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2775_
timestamp 0
transform 1 0 2490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2776_
timestamp 0
transform 1 0 3310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2777_
timestamp 0
transform -1 0 2790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2778_
timestamp 0
transform -1 0 3050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__2779_
timestamp 0
transform -1 0 7090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2780_
timestamp 0
transform -1 0 7330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__2781_
timestamp 0
transform 1 0 7810 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__2782_
timestamp 0
transform 1 0 7690 0 1 270
box -6 -8 26 268
use FILL  FILL_0__2783_
timestamp 0
transform 1 0 9630 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2784_
timestamp 0
transform 1 0 10770 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2785_
timestamp 0
transform 1 0 10150 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2786_
timestamp 0
transform 1 0 9870 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2787_
timestamp 0
transform 1 0 8330 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2788_
timestamp 0
transform 1 0 8590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2789_
timestamp 0
transform 1 0 8110 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2790_
timestamp 0
transform -1 0 7850 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2791_
timestamp 0
transform 1 0 6110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2792_
timestamp 0
transform 1 0 9730 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2793_
timestamp 0
transform 1 0 9930 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2794_
timestamp 0
transform -1 0 10190 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2795_
timestamp 0
transform 1 0 8370 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2796_
timestamp 0
transform 1 0 8350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2797_
timestamp 0
transform 1 0 10750 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2798_
timestamp 0
transform -1 0 9890 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2799_
timestamp 0
transform -1 0 8270 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2800_
timestamp 0
transform -1 0 7670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2801_
timestamp 0
transform 1 0 9610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2802_
timestamp 0
transform -1 0 9930 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2803_
timestamp 0
transform 1 0 8370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2804_
timestamp 0
transform -1 0 8270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2805_
timestamp 0
transform -1 0 10010 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2806_
timestamp 0
transform 1 0 9690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2807_
timestamp 0
transform -1 0 8310 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2808_
timestamp 0
transform -1 0 6550 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2809_
timestamp 0
transform 1 0 8070 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2810_
timestamp 0
transform -1 0 7490 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2811_
timestamp 0
transform 1 0 9970 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2812_
timestamp 0
transform 1 0 9610 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2813_
timestamp 0
transform 1 0 8190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2814_
timestamp 0
transform -1 0 8070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2815_
timestamp 0
transform -1 0 8150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2816_
timestamp 0
transform 1 0 9410 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2817_
timestamp 0
transform -1 0 10270 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2818_
timestamp 0
transform 1 0 11090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2819_
timestamp 0
transform 1 0 10070 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2820_
timestamp 0
transform -1 0 9850 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2821_
timestamp 0
transform -1 0 9710 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2822_
timestamp 0
transform -1 0 7430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2823_
timestamp 0
transform -1 0 9430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2824_
timestamp 0
transform -1 0 9170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2825_
timestamp 0
transform 1 0 8630 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2826_
timestamp 0
transform 1 0 8670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2827_
timestamp 0
transform 1 0 9090 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2828_
timestamp 0
transform 1 0 10210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2829_
timestamp 0
transform -1 0 9150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2830_
timestamp 0
transform 1 0 9770 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2831_
timestamp 0
transform 1 0 8950 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2832_
timestamp 0
transform -1 0 8870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2833_
timestamp 0
transform -1 0 8630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2834_
timestamp 0
transform -1 0 8210 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2835_
timestamp 0
transform -1 0 9230 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2836_
timestamp 0
transform -1 0 7930 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2837_
timestamp 0
transform 1 0 8010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2838_
timestamp 0
transform 1 0 9250 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2839_
timestamp 0
transform 1 0 9510 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2840_
timestamp 0
transform -1 0 9250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2841_
timestamp 0
transform 1 0 8150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2842_
timestamp 0
transform 1 0 11470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2843_
timestamp 0
transform -1 0 10970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2844_
timestamp 0
transform 1 0 10690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2845_
timestamp 0
transform 1 0 10430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2846_
timestamp 0
transform -1 0 10070 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2847_
timestamp 0
transform 1 0 10270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2848_
timestamp 0
transform -1 0 9550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2849_
timestamp 0
transform 1 0 10850 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__2850_
timestamp 0
transform 1 0 11010 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2851_
timestamp 0
transform 1 0 11250 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2852_
timestamp 0
transform 1 0 11950 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2853_
timestamp 0
transform 1 0 12010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2854_
timestamp 0
transform 1 0 11690 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2855_
timestamp 0
transform 1 0 11970 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2856_
timestamp 0
transform -1 0 9010 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2857_
timestamp 0
transform 1 0 9510 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2858_
timestamp 0
transform -1 0 9810 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2859_
timestamp 0
transform 1 0 10750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2860_
timestamp 0
transform 1 0 7630 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2861_
timestamp 0
transform 1 0 8310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2862_
timestamp 0
transform -1 0 7690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2863_
timestamp 0
transform 1 0 7390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2864_
timestamp 0
transform 1 0 9630 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2865_
timestamp 0
transform 1 0 8790 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2866_
timestamp 0
transform -1 0 6890 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2867_
timestamp 0
transform -1 0 8730 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2868_
timestamp 0
transform -1 0 8450 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2869_
timestamp 0
transform -1 0 8890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2870_
timestamp 0
transform 1 0 8530 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2871_
timestamp 0
transform 1 0 8490 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2872_
timestamp 0
transform 1 0 5430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2873_
timestamp 0
transform -1 0 5450 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2874_
timestamp 0
transform 1 0 5370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2875_
timestamp 0
transform -1 0 5730 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2876_
timestamp 0
transform 1 0 5410 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2877_
timestamp 0
transform 1 0 5990 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2878_
timestamp 0
transform -1 0 5730 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2879_
timestamp 0
transform -1 0 8870 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2880_
timestamp 0
transform -1 0 11870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2881_
timestamp 0
transform 1 0 11550 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2882_
timestamp 0
transform -1 0 9150 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2883_
timestamp 0
transform 1 0 8950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2884_
timestamp 0
transform -1 0 9270 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2885_
timestamp 0
transform -1 0 10450 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2886_
timestamp 0
transform 1 0 10410 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2887_
timestamp 0
transform -1 0 8830 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2888_
timestamp 0
transform -1 0 9110 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2889_
timestamp 0
transform 1 0 9390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2890_
timestamp 0
transform -1 0 9750 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__2891_
timestamp 0
transform -1 0 9690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2892_
timestamp 0
transform 1 0 9070 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2893_
timestamp 0
transform -1 0 9230 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2894_
timestamp 0
transform -1 0 11050 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2895_
timestamp 0
transform 1 0 10730 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2896_
timestamp 0
transform -1 0 11010 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2897_
timestamp 0
transform -1 0 10730 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2898_
timestamp 0
transform 1 0 9350 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2899_
timestamp 0
transform -1 0 9650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2900_
timestamp 0
transform 1 0 10330 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2901_
timestamp 0
transform -1 0 10350 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2902_
timestamp 0
transform 1 0 10530 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2903_
timestamp 0
transform -1 0 10650 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2904_
timestamp 0
transform -1 0 9810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2905_
timestamp 0
transform -1 0 9310 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2906_
timestamp 0
transform -1 0 8470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2907_
timestamp 0
transform -1 0 9030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2908_
timestamp 0
transform -1 0 10370 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2909_
timestamp 0
transform 1 0 11730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2910_
timestamp 0
transform 1 0 10810 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2911_
timestamp 0
transform 1 0 11670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2912_
timestamp 0
transform 1 0 11950 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__2913_
timestamp 0
transform 1 0 10550 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__2914_
timestamp 0
transform -1 0 7730 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2915_
timestamp 0
transform 1 0 10870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2916_
timestamp 0
transform 1 0 11110 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__2917_
timestamp 0
transform 1 0 10610 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2918_
timestamp 0
transform -1 0 10770 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2919_
timestamp 0
transform 1 0 8450 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2920_
timestamp 0
transform 1 0 11150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2921_
timestamp 0
transform 1 0 11670 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__2922_
timestamp 0
transform -1 0 11790 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2923_
timestamp 0
transform 1 0 11250 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2924_
timestamp 0
transform 1 0 10170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2925_
timestamp 0
transform 1 0 9930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2926_
timestamp 0
transform 1 0 10070 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2927_
timestamp 0
transform -1 0 9910 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2928_
timestamp 0
transform -1 0 10170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__2929_
timestamp 0
transform -1 0 10290 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__2930_
timestamp 0
transform -1 0 11170 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2931_
timestamp 0
transform -1 0 11430 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__2932_
timestamp 0
transform 1 0 11390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__2933_
timestamp 0
transform 1 0 11350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__2934_
timestamp 0
transform 1 0 11430 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__2935_
timestamp 0
transform 1 0 11510 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2936_
timestamp 0
transform 1 0 10450 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__2937_
timestamp 0
transform -1 0 3450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__2938_
timestamp 0
transform -1 0 7670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2939_
timestamp 0
transform 1 0 6430 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2940_
timestamp 0
transform -1 0 6210 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2941_
timestamp 0
transform -1 0 6130 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2942_
timestamp 0
transform 1 0 5030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2943_
timestamp 0
transform -1 0 6930 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__2944_
timestamp 0
transform 1 0 5310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2945_
timestamp 0
transform -1 0 6710 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2946_
timestamp 0
transform 1 0 6310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__2947_
timestamp 0
transform 1 0 7790 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2948_
timestamp 0
transform 1 0 7530 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2949_
timestamp 0
transform 1 0 5630 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__2950_
timestamp 0
transform -1 0 5970 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2951_
timestamp 0
transform 1 0 6730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2952_
timestamp 0
transform 1 0 6450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2953_
timestamp 0
transform 1 0 5610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2954_
timestamp 0
transform -1 0 5910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__2955_
timestamp 0
transform 1 0 6990 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2956_
timestamp 0
transform 1 0 6470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__2957_
timestamp 0
transform -1 0 8090 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__2958_
timestamp 0
transform 1 0 6470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__2959_
timestamp 0
transform 1 0 6210 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2960_
timestamp 0
transform -1 0 7090 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2961_
timestamp 0
transform 1 0 6470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2962_
timestamp 0
transform -1 0 6250 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__2963_
timestamp 0
transform -1 0 6550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2964_
timestamp 0
transform 1 0 4610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2965_
timestamp 0
transform 1 0 5670 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2966_
timestamp 0
transform -1 0 6570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__2967_
timestamp 0
transform -1 0 4990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2968_
timestamp 0
transform -1 0 5250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2969_
timestamp 0
transform 1 0 4330 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2970_
timestamp 0
transform 1 0 4690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2971_
timestamp 0
transform 1 0 4570 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2972_
timestamp 0
transform -1 0 6010 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2973_
timestamp 0
transform -1 0 6270 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2974_
timestamp 0
transform -1 0 6270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2975_
timestamp 0
transform 1 0 5730 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2976_
timestamp 0
transform -1 0 4650 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2977_
timestamp 0
transform -1 0 4910 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2978_
timestamp 0
transform 1 0 5170 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__2979_
timestamp 0
transform 1 0 5450 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__2980_
timestamp 0
transform -1 0 7330 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2981_
timestamp 0
transform -1 0 6290 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2982_
timestamp 0
transform -1 0 6570 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__2983_
timestamp 0
transform 1 0 7090 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2984_
timestamp 0
transform 1 0 6490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__2985_
timestamp 0
transform -1 0 6830 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2986_
timestamp 0
transform 1 0 6530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2987_
timestamp 0
transform 1 0 5970 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2988_
timestamp 0
transform -1 0 6250 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__2989_
timestamp 0
transform -1 0 7830 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2990_
timestamp 0
transform 1 0 6950 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__2991_
timestamp 0
transform -1 0 6810 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2992_
timestamp 0
transform -1 0 5110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__2993_
timestamp 0
transform -1 0 5970 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2994_
timestamp 0
transform 1 0 5430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2995_
timestamp 0
transform 1 0 6510 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2996_
timestamp 0
transform 1 0 6230 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__2997_
timestamp 0
transform 1 0 5950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2998_
timestamp 0
transform -1 0 5690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__2999_
timestamp 0
transform 1 0 6350 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3000_
timestamp 0
transform -1 0 5690 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__3001_
timestamp 0
transform 1 0 4910 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3002_
timestamp 0
transform -1 0 5410 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__3003_
timestamp 0
transform -1 0 5770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3004_
timestamp 0
transform -1 0 5190 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3005_
timestamp 0
transform -1 0 5450 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3006_
timestamp 0
transform -1 0 7350 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3007_
timestamp 0
transform 1 0 6770 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3008_
timestamp 0
transform 1 0 8570 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3009_
timestamp 0
transform 1 0 8030 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3010_
timestamp 0
transform 1 0 7050 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3011_
timestamp 0
transform -1 0 7150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3012_
timestamp 0
transform -1 0 7030 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3013_
timestamp 0
transform -1 0 7770 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3014_
timestamp 0
transform 1 0 6970 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3015_
timestamp 0
transform -1 0 7250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3016_
timestamp 0
transform -1 0 6010 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3017_
timestamp 0
transform -1 0 6810 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3018_
timestamp 0
transform -1 0 6490 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3019_
timestamp 0
transform -1 0 6750 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3020_
timestamp 0
transform 1 0 5390 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__3021_
timestamp 0
transform 1 0 5830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3022_
timestamp 0
transform 1 0 5630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__3023_
timestamp 0
transform -1 0 6710 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3024_
timestamp 0
transform -1 0 6630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3025_
timestamp 0
transform 1 0 5910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__3026_
timestamp 0
transform 1 0 5330 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__3027_
timestamp 0
transform -1 0 5430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3028_
timestamp 0
transform 1 0 5910 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3029_
timestamp 0
transform 1 0 6670 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3030_
timestamp 0
transform 1 0 4810 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__3031_
timestamp 0
transform 1 0 4350 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3032_
timestamp 0
transform -1 0 5130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3033_
timestamp 0
transform 1 0 5390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3034_
timestamp 0
transform -1 0 3330 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3035_
timestamp 0
transform -1 0 3890 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3036_
timestamp 0
transform -1 0 3390 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3037_
timestamp 0
transform -1 0 3270 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3038_
timestamp 0
transform 1 0 3490 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3039_
timestamp 0
transform -1 0 2990 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3040_
timestamp 0
transform 1 0 2870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3041_
timestamp 0
transform 1 0 3110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3042_
timestamp 0
transform -1 0 3670 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3043_
timestamp 0
transform -1 0 3770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3044_
timestamp 0
transform -1 0 3530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3045_
timestamp 0
transform 1 0 4330 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3046_
timestamp 0
transform 1 0 4050 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3047_
timestamp 0
transform -1 0 3010 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3048_
timestamp 0
transform 1 0 3050 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3049_
timestamp 0
transform -1 0 2750 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3050_
timestamp 0
transform 1 0 2790 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3051_
timestamp 0
transform 1 0 2530 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3052_
timestamp 0
transform 1 0 2430 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3053_
timestamp 0
transform 1 0 3190 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3054_
timestamp 0
transform -1 0 3470 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3055_
timestamp 0
transform 1 0 3290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3056_
timestamp 0
transform -1 0 3550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3057_
timestamp 0
transform 1 0 3750 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3058_
timestamp 0
transform 1 0 3930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3059_
timestamp 0
transform 1 0 4210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3060_
timestamp 0
transform 1 0 4050 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3061_
timestamp 0
transform 1 0 3530 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3062_
timestamp 0
transform -1 0 3770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3063_
timestamp 0
transform -1 0 5010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__3064_
timestamp 0
transform 1 0 4870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__3065_
timestamp 0
transform -1 0 4610 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3066_
timestamp 0
transform 1 0 4510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3067_
timestamp 0
transform -1 0 3610 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3068_
timestamp 0
transform -1 0 3350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3069_
timestamp 0
transform 1 0 3550 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3070_
timestamp 0
transform -1 0 4450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__3071_
timestamp 0
transform 1 0 4170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__3072_
timestamp 0
transform -1 0 4110 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3073_
timestamp 0
transform -1 0 4370 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3074_
timestamp 0
transform 1 0 5650 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3075_
timestamp 0
transform 1 0 5370 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3076_
timestamp 0
transform 1 0 3610 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3077_
timestamp 0
transform 1 0 3930 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3078_
timestamp 0
transform 1 0 3990 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3079_
timestamp 0
transform -1 0 4070 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3080_
timestamp 0
transform 1 0 6210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3081_
timestamp 0
transform -1 0 6870 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3082_
timestamp 0
transform 1 0 6570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3083_
timestamp 0
transform -1 0 3750 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3084_
timestamp 0
transform 1 0 3450 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3085_
timestamp 0
transform 1 0 3070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3086_
timestamp 0
transform -1 0 2790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3087_
timestamp 0
transform 1 0 4270 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3088_
timestamp 0
transform -1 0 4870 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3089_
timestamp 0
transform 1 0 3350 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3090_
timestamp 0
transform -1 0 3630 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3091_
timestamp 0
transform -1 0 6170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3092_
timestamp 0
transform 1 0 5390 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3093_
timestamp 0
transform 1 0 5650 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3094_
timestamp 0
transform 1 0 5370 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3095_
timestamp 0
transform -1 0 4570 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3096_
timestamp 0
transform 1 0 4270 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3097_
timestamp 0
transform -1 0 4030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3098_
timestamp 0
transform 1 0 3730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3099_
timestamp 0
transform -1 0 3790 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3100_
timestamp 0
transform -1 0 3610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3101_
timestamp 0
transform 1 0 4830 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3102_
timestamp 0
transform -1 0 5130 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3103_
timestamp 0
transform -1 0 4510 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3104_
timestamp 0
transform -1 0 4790 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3105_
timestamp 0
transform 1 0 5570 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3106_
timestamp 0
transform -1 0 5870 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3107_
timestamp 0
transform -1 0 3970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3108_
timestamp 0
transform 1 0 3670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3109_
timestamp 0
transform 1 0 6150 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3110_
timestamp 0
transform 1 0 3830 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3111_
timestamp 0
transform 1 0 5690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3112_
timestamp 0
transform -1 0 5110 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3113_
timestamp 0
transform -1 0 4570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3114_
timestamp 0
transform 1 0 4270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3115_
timestamp 0
transform 1 0 4790 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3116_
timestamp 0
transform 1 0 3730 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3117_
timestamp 0
transform 1 0 4350 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3118_
timestamp 0
transform -1 0 4650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3119_
timestamp 0
transform 1 0 4830 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3120_
timestamp 0
transform 1 0 4530 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3121_
timestamp 0
transform 1 0 5130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3122_
timestamp 0
transform 1 0 5410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3123_
timestamp 0
transform 1 0 5390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3124_
timestamp 0
transform -1 0 5690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3125_
timestamp 0
transform -1 0 4050 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3126_
timestamp 0
transform 1 0 3750 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3127_
timestamp 0
transform 1 0 6410 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3128_
timestamp 0
transform 1 0 5970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3129_
timestamp 0
transform 1 0 5370 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3130_
timestamp 0
transform -1 0 3290 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3131_
timestamp 0
transform -1 0 3530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3132_
timestamp 0
transform 1 0 4630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3133_
timestamp 0
transform 1 0 3870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3134_
timestamp 0
transform 1 0 5050 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3135_
timestamp 0
transform 1 0 4750 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3136_
timestamp 0
transform 1 0 5650 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3137_
timestamp 0
transform 1 0 5370 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3138_
timestamp 0
transform 1 0 5650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3139_
timestamp 0
transform 1 0 5370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3140_
timestamp 0
transform -1 0 5570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3141_
timestamp 0
transform -1 0 5830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3142_
timestamp 0
transform -1 0 4170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3143_
timestamp 0
transform -1 0 4430 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3144_
timestamp 0
transform 1 0 11510 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__3145_
timestamp 0
transform 1 0 11750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__3146_
timestamp 0
transform -1 0 11810 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__3147_
timestamp 0
transform 1 0 9430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__3148_
timestamp 0
transform -1 0 11810 0 1 790
box -6 -8 26 268
use FILL  FILL_0__3149_
timestamp 0
transform -1 0 11430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3150_
timestamp 0
transform -1 0 11710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3151_
timestamp 0
transform -1 0 10650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3152_
timestamp 0
transform 1 0 9290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3153_
timestamp 0
transform -1 0 9590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3154_
timestamp 0
transform -1 0 10110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3155_
timestamp 0
transform -1 0 10230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3156_
timestamp 0
transform -1 0 8870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__3157_
timestamp 0
transform -1 0 8910 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__3158_
timestamp 0
transform -1 0 8630 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__3159_
timestamp 0
transform -1 0 8610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__3160_
timestamp 0
transform 1 0 10450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3161_
timestamp 0
transform 1 0 10170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3162_
timestamp 0
transform -1 0 9710 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3163_
timestamp 0
transform 1 0 9430 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3164_
timestamp 0
transform -1 0 8910 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3165_
timestamp 0
transform -1 0 7130 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3166_
timestamp 0
transform 1 0 7530 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__3167_
timestamp 0
transform 1 0 7390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3168_
timestamp 0
transform 1 0 7550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3169_
timestamp 0
transform -1 0 8630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3170_
timestamp 0
transform -1 0 8350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3171_
timestamp 0
transform -1 0 9070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3172_
timestamp 0
transform -1 0 8070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3173_
timestamp 0
transform 1 0 8330 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3174_
timestamp 0
transform 1 0 7810 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3175_
timestamp 0
transform -1 0 7790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3176_
timestamp 0
transform -1 0 7510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3177_
timestamp 0
transform -1 0 11790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__3178_
timestamp 0
transform -1 0 11730 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3179_
timestamp 0
transform 1 0 11990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3180_
timestamp 0
transform 1 0 12050 0 1 790
box -6 -8 26 268
use FILL  FILL_0__3181_
timestamp 0
transform 1 0 12030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__3182_
timestamp 0
transform -1 0 11250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3183_
timestamp 0
transform 1 0 11510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3184_
timestamp 0
transform 1 0 11790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3185_
timestamp 0
transform 1 0 11810 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3186_
timestamp 0
transform 1 0 11990 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3187_
timestamp 0
transform 1 0 9850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__3188_
timestamp 0
transform 1 0 10730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3189_
timestamp 0
transform -1 0 10990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__3190_
timestamp 0
transform 1 0 11030 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3191_
timestamp 0
transform 1 0 10970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3192_
timestamp 0
transform -1 0 10690 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3193_
timestamp 0
transform 1 0 10110 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3194_
timestamp 0
transform 1 0 10730 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__3195_
timestamp 0
transform -1 0 10470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3196_
timestamp 0
transform 1 0 10370 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3197_
timestamp 0
transform -1 0 7230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3198_
timestamp 0
transform -1 0 4590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3199_
timestamp 0
transform 1 0 2750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__3200_
timestamp 0
transform 1 0 4730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__3201_
timestamp 0
transform 1 0 4450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__3202_
timestamp 0
transform 1 0 1510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__3203_
timestamp 0
transform 1 0 1470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3204_
timestamp 0
transform 1 0 1430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__3205_
timestamp 0
transform 1 0 990 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__3206_
timestamp 0
transform 1 0 1410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__3207_
timestamp 0
transform -1 0 1550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__3208_
timestamp 0
transform -1 0 890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__3209_
timestamp 0
transform -1 0 590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__3210_
timestamp 0
transform -1 0 4250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__3211_
timestamp 0
transform 1 0 4190 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__3212_
timestamp 0
transform 1 0 1150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__3213_
timestamp 0
transform 1 0 1050 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__3214_
timestamp 0
transform -1 0 2330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3215_
timestamp 0
transform 1 0 1750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3216_
timestamp 0
transform 1 0 5690 0 1 270
box -6 -8 26 268
use FILL  FILL_0__3217_
timestamp 0
transform -1 0 5990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__3218_
timestamp 0
transform 1 0 6030 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3219_
timestamp 0
transform -1 0 6310 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3220_
timestamp 0
transform 1 0 3650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3221_
timestamp 0
transform -1 0 3930 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3222_
timestamp 0
transform -1 0 3530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3223_
timestamp 0
transform 1 0 3250 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__3224_
timestamp 0
transform -1 0 3230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3225_
timestamp 0
transform 1 0 5370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__3226_
timestamp 0
transform 1 0 5090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__3227_
timestamp 0
transform -1 0 4210 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3228_
timestamp 0
transform -1 0 4410 0 1 270
box -6 -8 26 268
use FILL  FILL_0__3229_
timestamp 0
transform 1 0 2650 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__3230_
timestamp 0
transform -1 0 2690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__3231_
timestamp 0
transform 1 0 5930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__3232_
timestamp 0
transform 1 0 5910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__3364_
timestamp 0
transform 1 0 5190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3365_
timestamp 0
transform 1 0 4390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3366_
timestamp 0
transform 1 0 4870 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__3367_
timestamp 0
transform -1 0 4670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3368_
timestamp 0
transform -1 0 4930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3369_
timestamp 0
transform -1 0 5490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3370_
timestamp 0
transform 1 0 2630 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3371_
timestamp 0
transform 1 0 2130 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3372_
timestamp 0
transform -1 0 2250 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3373_
timestamp 0
transform -1 0 3910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3374_
timestamp 0
transform -1 0 2230 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3375_
timestamp 0
transform 1 0 2230 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3376_
timestamp 0
transform -1 0 2890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3377_
timestamp 0
transform 1 0 2350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3378_
timestamp 0
transform -1 0 2210 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3379_
timestamp 0
transform -1 0 1370 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3380_
timestamp 0
transform 1 0 1150 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3381_
timestamp 0
transform -1 0 1410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3382_
timestamp 0
transform -1 0 1870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3383_
timestamp 0
transform -1 0 1430 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3384_
timestamp 0
transform 1 0 1690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3385_
timestamp 0
transform 1 0 1390 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3386_
timestamp 0
transform -1 0 1970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3387_
timestamp 0
transform 1 0 2230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3388_
timestamp 0
transform -1 0 570 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3389_
timestamp 0
transform 1 0 2430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3390_
timestamp 0
transform 1 0 3250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3391_
timestamp 0
transform 1 0 2970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3392_
timestamp 0
transform -1 0 2810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3393_
timestamp 0
transform 1 0 2210 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3394_
timestamp 0
transform 1 0 610 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3395_
timestamp 0
transform -1 0 570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3396_
timestamp 0
transform -1 0 310 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3397_
timestamp 0
transform -1 0 330 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3398_
timestamp 0
transform -1 0 30 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3399_
timestamp 0
transform 1 0 10 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3400_
timestamp 0
transform -1 0 810 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3401_
timestamp 0
transform -1 0 1390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3402_
timestamp 0
transform 1 0 1370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3403_
timestamp 0
transform 1 0 1090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3404_
timestamp 0
transform -1 0 30 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3405_
timestamp 0
transform -1 0 290 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3406_
timestamp 0
transform -1 0 30 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3407_
timestamp 0
transform -1 0 310 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3408_
timestamp 0
transform -1 0 30 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3409_
timestamp 0
transform -1 0 30 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3410_
timestamp 0
transform 1 0 1350 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3411_
timestamp 0
transform 1 0 1070 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3412_
timestamp 0
transform -1 0 550 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3413_
timestamp 0
transform 1 0 290 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3414_
timestamp 0
transform 1 0 550 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0__3415_
timestamp 0
transform -1 0 870 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3416_
timestamp 0
transform 1 0 550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3417_
timestamp 0
transform -1 0 590 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3418_
timestamp 0
transform -1 0 290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3419_
timestamp 0
transform -1 0 1110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3420_
timestamp 0
transform 1 0 810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3421_
timestamp 0
transform 1 0 1110 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3422_
timestamp 0
transform 1 0 830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3423_
timestamp 0
transform 1 0 1130 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3424_
timestamp 0
transform -1 0 1150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3425_
timestamp 0
transform -1 0 870 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3426_
timestamp 0
transform 1 0 850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0__3427_
timestamp 0
transform -1 0 1370 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3428_
timestamp 0
transform 1 0 1050 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3429_
timestamp 0
transform -1 0 830 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3430_
timestamp 0
transform 1 0 1350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3431_
timestamp 0
transform 1 0 1070 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3432_
timestamp 0
transform -1 0 870 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3433_
timestamp 0
transform -1 0 30 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3434_
timestamp 0
transform -1 0 610 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3435_
timestamp 0
transform -1 0 890 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3436_
timestamp 0
transform -1 0 830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3437_
timestamp 0
transform 1 0 1650 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3438_
timestamp 0
transform 1 0 1110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3439_
timestamp 0
transform -1 0 1390 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3440_
timestamp 0
transform 1 0 1110 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3441_
timestamp 0
transform -1 0 550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3442_
timestamp 0
transform 1 0 1130 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3443_
timestamp 0
transform 1 0 1050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3444_
timestamp 0
transform -1 0 1950 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3445_
timestamp 0
transform 1 0 1630 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3446_
timestamp 0
transform 1 0 1990 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3447_
timestamp 0
transform 1 0 1890 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3448_
timestamp 0
transform -1 0 1690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3449_
timestamp 0
transform 1 0 1370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3450_
timestamp 0
transform -1 0 830 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3451_
timestamp 0
transform 1 0 1090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3452_
timestamp 0
transform 1 0 790 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3453_
timestamp 0
transform -1 0 2110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3454_
timestamp 0
transform 1 0 3030 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3455_
timestamp 0
transform -1 0 1970 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3456_
timestamp 0
transform -1 0 1630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3457_
timestamp 0
transform -1 0 2810 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3458_
timestamp 0
transform -1 0 1670 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3459_
timestamp 0
transform -1 0 1610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3460_
timestamp 0
transform 1 0 1650 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3461_
timestamp 0
transform -1 0 1870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3462_
timestamp 0
transform -1 0 1630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3463_
timestamp 0
transform -1 0 1390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3464_
timestamp 0
transform 1 0 1110 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3465_
timestamp 0
transform -1 0 1370 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3466_
timestamp 0
transform 1 0 1910 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3467_
timestamp 0
transform 1 0 1910 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3468_
timestamp 0
transform 1 0 2670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3469_
timestamp 0
transform 1 0 2530 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3470_
timestamp 0
transform -1 0 2430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3471_
timestamp 0
transform 1 0 2250 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3472_
timestamp 0
transform -1 0 2150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3473_
timestamp 0
transform 1 0 1390 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3474_
timestamp 0
transform -1 0 1650 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3475_
timestamp 0
transform 1 0 1130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3476_
timestamp 0
transform -1 0 870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3477_
timestamp 0
transform 1 0 290 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3478_
timestamp 0
transform -1 0 270 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3479_
timestamp 0
transform -1 0 30 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3480_
timestamp 0
transform -1 0 30 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3481_
timestamp 0
transform -1 0 30 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3482_
timestamp 0
transform 1 0 550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3483_
timestamp 0
transform -1 0 270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3484_
timestamp 0
transform 1 0 1890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3485_
timestamp 0
transform -1 0 1950 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3486_
timestamp 0
transform -1 0 1330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3487_
timestamp 0
transform -1 0 1650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3488_
timestamp 0
transform -1 0 1450 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3489_
timestamp 0
transform 1 0 1390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3490_
timestamp 0
transform 1 0 1070 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3491_
timestamp 0
transform -1 0 1150 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3492_
timestamp 0
transform 1 0 1050 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3493_
timestamp 0
transform -1 0 870 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3494_
timestamp 0
transform 1 0 790 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3495_
timestamp 0
transform -1 0 550 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3496_
timestamp 0
transform 1 0 310 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3497_
timestamp 0
transform -1 0 270 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3498_
timestamp 0
transform 1 0 570 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3499_
timestamp 0
transform -1 0 630 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3500_
timestamp 0
transform 1 0 570 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3501_
timestamp 0
transform 1 0 810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3502_
timestamp 0
transform -1 0 330 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3503_
timestamp 0
transform -1 0 310 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3504_
timestamp 0
transform -1 0 550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3505_
timestamp 0
transform -1 0 310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3506_
timestamp 0
transform -1 0 30 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3507_
timestamp 0
transform -1 0 30 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3508_
timestamp 0
transform 1 0 550 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3509_
timestamp 0
transform -1 0 810 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3510_
timestamp 0
transform -1 0 310 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3511_
timestamp 0
transform -1 0 30 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3512_
timestamp 0
transform 1 0 510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3513_
timestamp 0
transform -1 0 330 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3514_
timestamp 0
transform -1 0 270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3515_
timestamp 0
transform -1 0 30 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3516_
timestamp 0
transform -1 0 30 0 1 10150
box -6 -8 26 268
use FILL  FILL_0__3517_
timestamp 0
transform 1 0 570 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3518_
timestamp 0
transform 1 0 790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3519_
timestamp 0
transform 1 0 2490 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3520_
timestamp 0
transform 1 0 2770 0 1 9110
box -6 -8 26 268
use FILL  FILL_0__3521_
timestamp 0
transform 1 0 3250 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3522_
timestamp 0
transform 1 0 2950 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3523_
timestamp 0
transform 1 0 2510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3524_
timestamp 0
transform -1 0 890 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3525_
timestamp 0
transform -1 0 30 0 1 10670
box -6 -8 26 268
use FILL  FILL_0__3526_
timestamp 0
transform -1 0 30 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3527_
timestamp 0
transform -1 0 530 0 1 11190
box -6 -8 26 268
use FILL  FILL_0__3528_
timestamp 0
transform -1 0 550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_0__3529_
timestamp 0
transform -1 0 30 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0__3530_
timestamp 0
transform -1 0 30 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3531_
timestamp 0
transform 1 0 10 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3532_
timestamp 0
transform 1 0 250 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3533_
timestamp 0
transform -1 0 30 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3534_
timestamp 0
transform -1 0 550 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3535_
timestamp 0
transform -1 0 310 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0__3536_
timestamp 0
transform -1 0 290 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3537_
timestamp 0
transform -1 0 1650 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3538_
timestamp 0
transform 1 0 2410 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3539_
timestamp 0
transform -1 0 2510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3540_
timestamp 0
transform -1 0 2250 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3541_
timestamp 0
transform -1 0 1970 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3542_
timestamp 0
transform -1 0 2150 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3543_
timestamp 0
transform 1 0 1550 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3544_
timestamp 0
transform 1 0 1910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3545_
timestamp 0
transform 1 0 1710 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3546_
timestamp 0
transform 1 0 1830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0__3547_
timestamp 0
transform -1 0 2490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3548_
timestamp 0
transform 1 0 2190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0__3549_
timestamp 0
transform -1 0 2290 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3550_
timestamp 0
transform 1 0 1990 0 1 11710
box -6 -8 26 268
use FILL  FILL_0__3551_
timestamp 0
transform -1 0 2470 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3552_
timestamp 0
transform 1 0 2170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0__3553_
timestamp 0
transform -1 0 1710 0 1 8070
box -6 -8 26 268
use FILL  FILL_0__3554_
timestamp 0
transform 1 0 850 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3555_
timestamp 0
transform 1 0 250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3556_
timestamp 0
transform 1 0 1110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0__3557_
timestamp 0
transform -1 0 3010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3558_
timestamp 0
transform 1 0 2710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0__3559_
timestamp 0
transform -1 0 2470 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3560_
timestamp 0
transform 1 0 2170 0 1 9630
box -6 -8 26 268
use FILL  FILL_0__3561_
timestamp 0
transform -1 0 1890 0 1 7550
box -6 -8 26 268
use FILL  FILL_0__3562_
timestamp 0
transform -1 0 2710 0 1 8590
box -6 -8 26 268
use FILL  FILL_0__3563_
timestamp 0
transform 1 0 2110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0__3564_
timestamp 0
transform 1 0 2390 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3565_
timestamp 0
transform -1 0 1390 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3566_
timestamp 0
transform -1 0 1650 0 1 7030
box -6 -8 26 268
use FILL  FILL_0__3579_
timestamp 0
transform -1 0 4990 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3580_
timestamp 0
transform -1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__3581_
timestamp 0
transform -1 0 3410 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3582_
timestamp 0
transform -1 0 3150 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3583_
timestamp 0
transform -1 0 5270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__3584_
timestamp 0
transform 1 0 4450 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3585_
timestamp 0
transform 1 0 2870 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3586_
timestamp 0
transform -1 0 5790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__3587_
timestamp 0
transform 1 0 10 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3588_
timestamp 0
transform -1 0 30 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__3589_
timestamp 0
transform -1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__3590_
timestamp 0
transform -1 0 30 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__3591_
timestamp 0
transform -1 0 310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3592_
timestamp 0
transform -1 0 30 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__3593_
timestamp 0
transform -1 0 4730 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3594_
timestamp 0
transform 1 0 5770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__3595_
timestamp 0
transform 1 0 5510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__3596_
timestamp 0
transform -1 0 810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3597_
timestamp 0
transform -1 0 30 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__3598_
timestamp 0
transform -1 0 290 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__3599_
timestamp 0
transform -1 0 30 0 1 6510
box -6 -8 26 268
use FILL  FILL_0__3600_
timestamp 0
transform -1 0 30 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__3601_
timestamp 0
transform -1 0 30 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__3602_
timestamp 0
transform -1 0 1650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__3603_
timestamp 0
transform 1 0 6810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 7830 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 9330 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 8090 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 10950 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform 1 0 550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform -1 0 12030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 9530 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 6990 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 810 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 10070 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform -1 0 850 0 1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform -1 0 5930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform 1 0 11490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform -1 0 6110 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform 1 0 6730 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform -1 0 3270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform -1 0 3890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform 1 0 7130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform -1 0 6950 0 1 11190
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform 1 0 5270 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 8510 0 1 11190
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform -1 0 8430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 1390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform 1 0 3370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform -1 0 4270 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform 1 0 8110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform 1 0 5050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 1190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert39
timestamp 0
transform 1 0 6270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert40
timestamp 0
transform 1 0 7630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert41
timestamp 0
transform -1 0 8770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert42
timestamp 0
transform -1 0 6910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert43
timestamp 0
transform -1 0 8810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert44
timestamp 0
transform -1 0 8930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert45
timestamp 0
transform 1 0 10990 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert46
timestamp 0
transform 1 0 9430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert47
timestamp 0
transform 1 0 9150 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert48
timestamp 0
transform 1 0 6890 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert49
timestamp 0
transform 1 0 7150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert50
timestamp 0
transform -1 0 7530 0 1 9110
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert51
timestamp 0
transform 1 0 7490 0 1 10150
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert52
timestamp 0
transform 1 0 8890 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert53
timestamp 0
transform 1 0 9930 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert54
timestamp 0
transform 1 0 8770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert55
timestamp 0
transform 1 0 8630 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert56
timestamp 0
transform -1 0 2170 0 1 8590
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert57
timestamp 0
transform 1 0 2470 0 1 11190
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert58
timestamp 0
transform 1 0 2610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert59
timestamp 0
transform -1 0 2170 0 1 10670
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert60
timestamp 0
transform -1 0 10430 0 1 7550
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert61
timestamp 0
transform 1 0 10490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert62
timestamp 0
transform 1 0 10450 0 1 8070
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert63
timestamp 0
transform -1 0 9110 0 1 7550
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert64
timestamp 0
transform -1 0 8550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert65
timestamp 0
transform 1 0 5150 0 1 270
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert66
timestamp 0
transform 1 0 5670 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert67
timestamp 0
transform -1 0 2970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert68
timestamp 0
transform 1 0 3090 0 1 270
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert69
timestamp 0
transform -1 0 6590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert70
timestamp 0
transform 1 0 8530 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert71
timestamp 0
transform -1 0 9190 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert72
timestamp 0
transform -1 0 6710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert73
timestamp 0
transform 1 0 8870 0 -1 7030
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert74
timestamp 0
transform 1 0 10730 0 1 7030
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert75
timestamp 0
transform 1 0 2510 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert76
timestamp 0
transform -1 0 3010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert77
timestamp 0
transform 1 0 10390 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert78
timestamp 0
transform 1 0 9250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert79
timestamp 0
transform -1 0 8290 0 1 7550
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert80
timestamp 0
transform 1 0 7090 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert81
timestamp 0
transform 1 0 7550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert82
timestamp 0
transform -1 0 7530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert83
timestamp 0
transform -1 0 7310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert84
timestamp 0
transform 1 0 9370 0 1 8590
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert85
timestamp 0
transform -1 0 8850 0 1 8590
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert86
timestamp 0
transform -1 0 9450 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert87
timestamp 0
transform 1 0 9350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert88
timestamp 0
transform -1 0 10690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert89
timestamp 0
transform 1 0 9330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert90
timestamp 0
transform 1 0 5310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert91
timestamp 0
transform -1 0 4850 0 1 10670
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert92
timestamp 0
transform -1 0 4690 0 -1 9630
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert93
timestamp 0
transform 1 0 5110 0 1 10150
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert94
timestamp 0
transform -1 0 11270 0 1 9630
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert95
timestamp 0
transform -1 0 11310 0 -1 10150
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert96
timestamp 0
transform -1 0 10030 0 1 11710
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert97
timestamp 0
transform 1 0 11390 0 1 11710
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert28
timestamp 0
transform -1 0 5970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert29
timestamp 0
transform -1 0 2150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert30
timestamp 0
transform 1 0 4490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert31
timestamp 0
transform -1 0 3190 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert32
timestamp 0
transform 1 0 7090 0 -1 8070
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert33
timestamp 0
transform 1 0 5670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert34
timestamp 0
transform -1 0 2430 0 1 10670
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert35
timestamp 0
transform -1 0 5190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert36
timestamp 0
transform -1 0 2310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert37
timestamp 0
transform 1 0 7330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert38
timestamp 0
transform -1 0 4310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__1688_
timestamp 0
transform -1 0 850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1689_
timestamp 0
transform -1 0 310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1690_
timestamp 0
transform -1 0 570 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1691_
timestamp 0
transform 1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1692_
timestamp 0
transform -1 0 290 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1693_
timestamp 0
transform 1 0 530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1694_
timestamp 0
transform -1 0 5530 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1695_
timestamp 0
transform -1 0 310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1696_
timestamp 0
transform -1 0 310 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1697_
timestamp 0
transform -1 0 1430 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__1698_
timestamp 0
transform -1 0 3370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1699_
timestamp 0
transform 1 0 2810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1700_
timestamp 0
transform -1 0 3850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__1701_
timestamp 0
transform -1 0 550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1702_
timestamp 0
transform -1 0 550 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1703_
timestamp 0
transform 1 0 3190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1704_
timestamp 0
transform -1 0 330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1705_
timestamp 0
transform 1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1706_
timestamp 0
transform -1 0 3810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1707_
timestamp 0
transform -1 0 570 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1708_
timestamp 0
transform 1 0 570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1709_
timestamp 0
transform 1 0 4090 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1710_
timestamp 0
transform -1 0 5570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1711_
timestamp 0
transform 1 0 5110 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1712_
timestamp 0
transform 1 0 7250 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1713_
timestamp 0
transform -1 0 9630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1714_
timestamp 0
transform -1 0 9830 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1715_
timestamp 0
transform -1 0 8510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1716_
timestamp 0
transform 1 0 11270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1717_
timestamp 0
transform 1 0 11070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1718_
timestamp 0
transform 1 0 11890 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1719_
timestamp 0
transform -1 0 8770 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1720_
timestamp 0
transform -1 0 10090 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1721_
timestamp 0
transform -1 0 10110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1722_
timestamp 0
transform -1 0 9870 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1723_
timestamp 0
transform 1 0 9970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1724_
timestamp 0
transform 1 0 9190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1725_
timestamp 0
transform 1 0 9030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1726_
timestamp 0
transform 1 0 10130 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1727_
timestamp 0
transform -1 0 8750 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1728_
timestamp 0
transform 1 0 11530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1729_
timestamp 0
transform 1 0 10130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1730_
timestamp 0
transform 1 0 8310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1731_
timestamp 0
transform 1 0 8550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1732_
timestamp 0
transform -1 0 7750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1733_
timestamp 0
transform 1 0 9690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1734_
timestamp 0
transform 1 0 7390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1735_
timestamp 0
transform 1 0 10830 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1736_
timestamp 0
transform -1 0 10630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1737_
timestamp 0
transform -1 0 10890 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1738_
timestamp 0
transform -1 0 10270 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1739_
timestamp 0
transform -1 0 10270 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1740_
timestamp 0
transform 1 0 10490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1741_
timestamp 0
transform -1 0 8390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1742_
timestamp 0
transform -1 0 8290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1743_
timestamp 0
transform -1 0 9850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1744_
timestamp 0
transform 1 0 9730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1745_
timestamp 0
transform -1 0 9430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1746_
timestamp 0
transform 1 0 11290 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1747_
timestamp 0
transform 1 0 10770 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1748_
timestamp 0
transform 1 0 7490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1749_
timestamp 0
transform 1 0 7910 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1750_
timestamp 0
transform -1 0 8030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1751_
timestamp 0
transform 1 0 7430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1752_
timestamp 0
transform -1 0 8850 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1753_
timestamp 0
transform 1 0 9710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1754_
timestamp 0
transform -1 0 8250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1755_
timestamp 0
transform -1 0 8830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__1756_
timestamp 0
transform -1 0 11170 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1757_
timestamp 0
transform 1 0 11030 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1758_
timestamp 0
transform -1 0 9090 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1759_
timestamp 0
transform -1 0 7330 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__1760_
timestamp 0
transform 1 0 8830 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__1761_
timestamp 0
transform -1 0 9550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1762_
timestamp 0
transform 1 0 10570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1763_
timestamp 0
transform -1 0 9010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1764_
timestamp 0
transform 1 0 11270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1765_
timestamp 0
transform 1 0 8090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1766_
timestamp 0
transform 1 0 8470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1767_
timestamp 0
transform 1 0 9170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__1768_
timestamp 0
transform 1 0 8030 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__1769_
timestamp 0
transform 1 0 8550 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__1770_
timestamp 0
transform 1 0 8990 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__1771_
timestamp 0
transform 1 0 8950 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__1772_
timestamp 0
transform 1 0 8670 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__1773_
timestamp 0
transform 1 0 10750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1774_
timestamp 0
transform 1 0 10750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1775_
timestamp 0
transform 1 0 9990 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1776_
timestamp 0
transform -1 0 7990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1777_
timestamp 0
transform 1 0 8030 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1778_
timestamp 0
transform -1 0 7510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1779_
timestamp 0
transform 1 0 5650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1780_
timestamp 0
transform -1 0 4050 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1781_
timestamp 0
transform -1 0 10770 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1782_
timestamp 0
transform 1 0 8250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1783_
timestamp 0
transform 1 0 10490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1784_
timestamp 0
transform -1 0 9970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1785_
timestamp 0
transform -1 0 9730 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1786_
timestamp 0
transform 1 0 10150 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1787_
timestamp 0
transform -1 0 9090 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1788_
timestamp 0
transform -1 0 8510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1789_
timestamp 0
transform 1 0 9950 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1790_
timestamp 0
transform -1 0 10010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1791_
timestamp 0
transform -1 0 10090 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1792_
timestamp 0
transform -1 0 9630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1793_
timestamp 0
transform -1 0 9370 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1794_
timestamp 0
transform 1 0 9090 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1795_
timestamp 0
transform -1 0 8290 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1796_
timestamp 0
transform -1 0 8230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1797_
timestamp 0
transform 1 0 7070 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1798_
timestamp 0
transform 1 0 7330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1799_
timestamp 0
transform -1 0 9350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1800_
timestamp 0
transform 1 0 11230 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1801_
timestamp 0
transform 1 0 9250 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1802_
timestamp 0
transform -1 0 8910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1803_
timestamp 0
transform 1 0 10510 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1804_
timestamp 0
transform -1 0 8530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1805_
timestamp 0
transform -1 0 8630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1806_
timestamp 0
transform 1 0 7570 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1807_
timestamp 0
transform -1 0 8030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1808_
timestamp 0
transform -1 0 8350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1809_
timestamp 0
transform 1 0 8570 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1810_
timestamp 0
transform 1 0 7970 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1811_
timestamp 0
transform -1 0 7710 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1812_
timestamp 0
transform -1 0 8350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1813_
timestamp 0
transform -1 0 8070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1814_
timestamp 0
transform -1 0 7810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1815_
timestamp 0
transform 1 0 7830 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1816_
timestamp 0
transform -1 0 3830 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1817_
timestamp 0
transform 1 0 1310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1818_
timestamp 0
transform -1 0 6130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1819_
timestamp 0
transform -1 0 890 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1820_
timestamp 0
transform 1 0 330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1821_
timestamp 0
transform 1 0 850 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1822_
timestamp 0
transform -1 0 310 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1823_
timestamp 0
transform 1 0 1670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1824_
timestamp 0
transform 1 0 1250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1825_
timestamp 0
transform -1 0 1090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1826_
timestamp 0
transform -1 0 350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1827_
timestamp 0
transform 1 0 850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1828_
timestamp 0
transform -1 0 1450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1829_
timestamp 0
transform -1 0 590 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1830_
timestamp 0
transform -1 0 1390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1831_
timestamp 0
transform 1 0 1970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1832_
timestamp 0
transform -1 0 7970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1833_
timestamp 0
transform 1 0 9610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1834_
timestamp 0
transform 1 0 9190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1835_
timestamp 0
transform -1 0 7710 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1836_
timestamp 0
transform -1 0 6370 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1837_
timestamp 0
transform -1 0 7710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1838_
timestamp 0
transform -1 0 7150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1839_
timestamp 0
transform -1 0 6130 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1840_
timestamp 0
transform 1 0 8510 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1841_
timestamp 0
transform -1 0 8130 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1842_
timestamp 0
transform -1 0 6890 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1843_
timestamp 0
transform -1 0 6610 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1844_
timestamp 0
transform 1 0 9030 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1845_
timestamp 0
transform 1 0 9570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1846_
timestamp 0
transform -1 0 9170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1847_
timestamp 0
transform -1 0 8330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1848_
timestamp 0
transform 1 0 11170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1849_
timestamp 0
transform -1 0 11490 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1850_
timestamp 0
transform -1 0 10950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1851_
timestamp 0
transform 1 0 10310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1852_
timestamp 0
transform -1 0 10370 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1853_
timestamp 0
transform -1 0 10390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1854_
timestamp 0
transform -1 0 7370 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1855_
timestamp 0
transform 1 0 7350 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1856_
timestamp 0
transform 1 0 7630 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1857_
timestamp 0
transform -1 0 8770 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__1858_
timestamp 0
transform -1 0 9310 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1859_
timestamp 0
transform -1 0 8770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1860_
timestamp 0
transform 1 0 9030 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1861_
timestamp 0
transform 1 0 6770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1862_
timestamp 0
transform -1 0 8270 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__1863_
timestamp 0
transform 1 0 7630 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1864_
timestamp 0
transform -1 0 6270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1865_
timestamp 0
transform -1 0 7710 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__1866_
timestamp 0
transform -1 0 7170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1867_
timestamp 0
transform -1 0 7950 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1868_
timestamp 0
transform 1 0 7670 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1869_
timestamp 0
transform -1 0 5970 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__1870_
timestamp 0
transform 1 0 9310 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1871_
timestamp 0
transform 1 0 8790 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1872_
timestamp 0
transform -1 0 8530 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1873_
timestamp 0
transform -1 0 7730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1874_
timestamp 0
transform -1 0 7450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1875_
timestamp 0
transform -1 0 8250 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1876_
timestamp 0
transform -1 0 6890 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1877_
timestamp 0
transform -1 0 5730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__1878_
timestamp 0
transform 1 0 6610 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1879_
timestamp 0
transform -1 0 7410 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1880_
timestamp 0
transform 1 0 5930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__1881_
timestamp 0
transform 1 0 5930 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__1882_
timestamp 0
transform -1 0 4890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__1883_
timestamp 0
transform -1 0 7790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1884_
timestamp 0
transform -1 0 8030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1885_
timestamp 0
transform -1 0 8590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1886_
timestamp 0
transform 1 0 8430 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1887_
timestamp 0
transform -1 0 8410 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1888_
timestamp 0
transform 1 0 11550 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1889_
timestamp 0
transform -1 0 8410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1890_
timestamp 0
transform 1 0 9670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1891_
timestamp 0
transform 1 0 8830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1892_
timestamp 0
transform -1 0 8550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1893_
timestamp 0
transform 1 0 12070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1894_
timestamp 0
transform 1 0 12050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1895_
timestamp 0
transform 1 0 12070 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1896_
timestamp 0
transform -1 0 10690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1897_
timestamp 0
transform -1 0 9090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1898_
timestamp 0
transform 1 0 8970 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1899_
timestamp 0
transform 1 0 7410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1900_
timestamp 0
transform 1 0 9610 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1901_
timestamp 0
transform 1 0 7950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1902_
timestamp 0
transform -1 0 8170 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1903_
timestamp 0
transform 1 0 7890 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1904_
timestamp 0
transform 1 0 11810 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1905_
timestamp 0
transform 1 0 11570 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1906_
timestamp 0
transform -1 0 6450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1907_
timestamp 0
transform -1 0 6990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1908_
timestamp 0
transform -1 0 6910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1909_
timestamp 0
transform -1 0 6670 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1910_
timestamp 0
transform -1 0 6170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1911_
timestamp 0
transform 1 0 6750 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1912_
timestamp 0
transform 1 0 6210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1913_
timestamp 0
transform 1 0 6150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1914_
timestamp 0
transform 1 0 5650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1915_
timestamp 0
transform 1 0 5170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1916_
timestamp 0
transform 1 0 5170 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__1917_
timestamp 0
transform -1 0 3670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__1918_
timestamp 0
transform 1 0 3550 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__1919_
timestamp 0
transform -1 0 3830 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__1920_
timestamp 0
transform -1 0 3550 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__1921_
timestamp 0
transform -1 0 1670 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__1922_
timestamp 0
transform 1 0 7470 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1923_
timestamp 0
transform 1 0 7730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1924_
timestamp 0
transform -1 0 6330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1925_
timestamp 0
transform -1 0 4570 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1926_
timestamp 0
transform -1 0 3930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1927_
timestamp 0
transform 1 0 1970 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__1928_
timestamp 0
transform -1 0 3130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__1929_
timestamp 0
transform 1 0 4510 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__1930_
timestamp 0
transform 1 0 3070 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__1931_
timestamp 0
transform -1 0 2850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__1932_
timestamp 0
transform -1 0 1450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1933_
timestamp 0
transform -1 0 8410 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1934_
timestamp 0
transform 1 0 3810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1935_
timestamp 0
transform -1 0 3830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1936_
timestamp 0
transform -1 0 2510 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1937_
timestamp 0
transform -1 0 1170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1938_
timestamp 0
transform -1 0 3530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1939_
timestamp 0
transform -1 0 4090 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1940_
timestamp 0
transform -1 0 3310 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1941_
timestamp 0
transform -1 0 3250 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1942_
timestamp 0
transform -1 0 1750 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__1943_
timestamp 0
transform -1 0 3550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1944_
timestamp 0
transform -1 0 3650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1945_
timestamp 0
transform -1 0 2910 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1946_
timestamp 0
transform -1 0 1470 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__1947_
timestamp 0
transform -1 0 4890 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__1948_
timestamp 0
transform 1 0 5090 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__1949_
timestamp 0
transform 1 0 5150 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__1950_
timestamp 0
transform -1 0 4890 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__1951_
timestamp 0
transform -1 0 1930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1952_
timestamp 0
transform 1 0 4050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1953_
timestamp 0
transform 1 0 3990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1954_
timestamp 0
transform 1 0 4130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1955_
timestamp 0
transform -1 0 1650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1956_
timestamp 0
transform -1 0 4270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__1957_
timestamp 0
transform 1 0 4850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__1958_
timestamp 0
transform -1 0 5130 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__1959_
timestamp 0
transform -1 0 4110 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__1960_
timestamp 0
transform -1 0 2270 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1961_
timestamp 0
transform 1 0 4090 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1962_
timestamp 0
transform 1 0 3850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1963_
timestamp 0
transform 1 0 3630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1964_
timestamp 0
transform 1 0 1970 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1965_
timestamp 0
transform 1 0 6350 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__1966_
timestamp 0
transform 1 0 6290 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1967_
timestamp 0
transform 1 0 7130 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1968_
timestamp 0
transform 1 0 6590 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1969_
timestamp 0
transform -1 0 3250 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__1970_
timestamp 0
transform 1 0 2790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1971_
timestamp 0
transform -1 0 4670 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1972_
timestamp 0
transform 1 0 3530 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1973_
timestamp 0
transform -1 0 3550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1974_
timestamp 0
transform -1 0 3050 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__1975_
timestamp 0
transform 1 0 2950 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__1976_
timestamp 0
transform -1 0 3050 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__1977_
timestamp 0
transform 1 0 4330 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__1978_
timestamp 0
transform 1 0 3030 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__1979_
timestamp 0
transform -1 0 2770 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__1980_
timestamp 0
transform -1 0 2290 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1981_
timestamp 0
transform 1 0 5910 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1982_
timestamp 0
transform 1 0 6030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1983_
timestamp 0
transform 1 0 6230 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1984_
timestamp 0
transform 1 0 5230 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1985_
timestamp 0
transform -1 0 4730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1986_
timestamp 0
transform 1 0 2510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__1987_
timestamp 0
transform -1 0 7230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1988_
timestamp 0
transform 1 0 7530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1989_
timestamp 0
transform 1 0 7590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1990_
timestamp 0
transform -1 0 7390 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1991_
timestamp 0
transform -1 0 7670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1992_
timestamp 0
transform 1 0 10410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1993_
timestamp 0
transform 1 0 9530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__1994_
timestamp 0
transform -1 0 6210 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__1995_
timestamp 0
transform 1 0 6590 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1996_
timestamp 0
transform -1 0 6730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1997_
timestamp 0
transform 1 0 6430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1998_
timestamp 0
transform 1 0 6430 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__1999_
timestamp 0
transform 1 0 7490 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2000_
timestamp 0
transform 1 0 6410 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2001_
timestamp 0
transform 1 0 6650 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2002_
timestamp 0
transform 1 0 6610 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2003_
timestamp 0
transform 1 0 9490 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2004_
timestamp 0
transform 1 0 7430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2005_
timestamp 0
transform -1 0 7230 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2006_
timestamp 0
transform 1 0 6710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2007_
timestamp 0
transform 1 0 6550 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2008_
timestamp 0
transform -1 0 6190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2009_
timestamp 0
transform 1 0 6790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2010_
timestamp 0
transform -1 0 7010 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2011_
timestamp 0
transform 1 0 7250 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2012_
timestamp 0
transform -1 0 9390 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2013_
timestamp 0
transform 1 0 10530 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2014_
timestamp 0
transform -1 0 10790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2015_
timestamp 0
transform -1 0 6230 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2016_
timestamp 0
transform -1 0 7270 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2017_
timestamp 0
transform -1 0 7050 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2018_
timestamp 0
transform 1 0 7290 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2019_
timestamp 0
transform 1 0 9370 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2020_
timestamp 0
transform -1 0 10270 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2021_
timestamp 0
transform -1 0 7310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2022_
timestamp 0
transform 1 0 7550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2023_
timestamp 0
transform -1 0 7850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2024_
timestamp 0
transform 1 0 6070 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2025_
timestamp 0
transform -1 0 5950 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2026_
timestamp 0
transform 1 0 9650 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2027_
timestamp 0
transform 1 0 10190 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2028_
timestamp 0
transform -1 0 10190 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2029_
timestamp 0
transform -1 0 11070 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2030_
timestamp 0
transform 1 0 10690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2031_
timestamp 0
transform -1 0 10990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2032_
timestamp 0
transform 1 0 8910 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2033_
timestamp 0
transform 1 0 8370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2034_
timestamp 0
transform 1 0 8610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2035_
timestamp 0
transform 1 0 8570 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2036_
timestamp 0
transform 1 0 11530 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2037_
timestamp 0
transform 1 0 11730 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2038_
timestamp 0
transform -1 0 7570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2039_
timestamp 0
transform -1 0 6650 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2040_
timestamp 0
transform 1 0 10910 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2041_
timestamp 0
transform 1 0 10990 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2042_
timestamp 0
transform -1 0 10070 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2043_
timestamp 0
transform -1 0 10450 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2044_
timestamp 0
transform -1 0 10970 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2045_
timestamp 0
transform -1 0 11310 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2046_
timestamp 0
transform 1 0 8790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2047_
timestamp 0
transform -1 0 9350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2048_
timestamp 0
transform 1 0 9150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2049_
timestamp 0
transform 1 0 9290 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2050_
timestamp 0
transform 1 0 9050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2051_
timestamp 0
transform 1 0 8750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2052_
timestamp 0
transform 1 0 9030 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2053_
timestamp 0
transform -1 0 9590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2054_
timestamp 0
transform 1 0 9810 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2055_
timestamp 0
transform -1 0 6450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2056_
timestamp 0
transform -1 0 6030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2057_
timestamp 0
transform 1 0 10230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2058_
timestamp 0
transform -1 0 9970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2059_
timestamp 0
transform -1 0 10110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2060_
timestamp 0
transform -1 0 9870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2061_
timestamp 0
transform 1 0 10050 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2062_
timestamp 0
transform -1 0 9130 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2063_
timestamp 0
transform 1 0 8210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2064_
timestamp 0
transform -1 0 7890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2065_
timestamp 0
transform -1 0 8710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2066_
timestamp 0
transform 1 0 8690 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2067_
timestamp 0
transform -1 0 7950 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2068_
timestamp 0
transform -1 0 8230 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2069_
timestamp 0
transform 1 0 7950 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2070_
timestamp 0
transform -1 0 8250 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2071_
timestamp 0
transform -1 0 8530 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2072_
timestamp 0
transform 1 0 8750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2073_
timestamp 0
transform 1 0 9010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2074_
timestamp 0
transform 1 0 9230 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2075_
timestamp 0
transform -1 0 9530 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2076_
timestamp 0
transform 1 0 11190 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2077_
timestamp 0
transform -1 0 11250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2078_
timestamp 0
transform -1 0 11050 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2079_
timestamp 0
transform 1 0 11190 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2080_
timestamp 0
transform -1 0 11030 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2081_
timestamp 0
transform 1 0 11030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2082_
timestamp 0
transform 1 0 10290 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2083_
timestamp 0
transform 1 0 9550 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2084_
timestamp 0
transform 1 0 11570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2085_
timestamp 0
transform 1 0 10990 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2086_
timestamp 0
transform 1 0 11490 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2087_
timestamp 0
transform 1 0 11510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2088_
timestamp 0
transform -1 0 12070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2089_
timestamp 0
transform 1 0 11790 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2090_
timestamp 0
transform 1 0 11970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2091_
timestamp 0
transform 1 0 9870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2092_
timestamp 0
transform 1 0 10490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2093_
timestamp 0
transform -1 0 11050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2094_
timestamp 0
transform 1 0 11290 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2095_
timestamp 0
transform -1 0 10950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2096_
timestamp 0
transform 1 0 11470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2097_
timestamp 0
transform -1 0 11810 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2098_
timestamp 0
transform -1 0 11990 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2099_
timestamp 0
transform -1 0 11290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2100_
timestamp 0
transform 1 0 11250 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2101_
timestamp 0
transform -1 0 11210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2102_
timestamp 0
transform -1 0 11590 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2103_
timestamp 0
transform 1 0 12070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2104_
timestamp 0
transform 1 0 12070 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2105_
timestamp 0
transform -1 0 11530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2106_
timestamp 0
transform -1 0 11510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2107_
timestamp 0
transform -1 0 12070 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2108_
timestamp 0
transform 1 0 8810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2109_
timestamp 0
transform 1 0 12070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2110_
timestamp 0
transform -1 0 12090 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2111_
timestamp 0
transform -1 0 12090 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2112_
timestamp 0
transform -1 0 11990 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2113_
timestamp 0
transform 1 0 11750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2114_
timestamp 0
transform 1 0 10530 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2115_
timestamp 0
transform -1 0 9270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2116_
timestamp 0
transform -1 0 10150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2117_
timestamp 0
transform -1 0 10750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2118_
timestamp 0
transform -1 0 10710 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2119_
timestamp 0
transform 1 0 10610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2120_
timestamp 0
transform 1 0 10650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2121_
timestamp 0
transform -1 0 10390 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2122_
timestamp 0
transform 1 0 10590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2123_
timestamp 0
transform -1 0 8090 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2124_
timestamp 0
transform -1 0 7790 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2125_
timestamp 0
transform -1 0 10150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2126_
timestamp 0
transform 1 0 10550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2127_
timestamp 0
transform -1 0 6970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2128_
timestamp 0
transform -1 0 9110 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2129_
timestamp 0
transform 1 0 7230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2130_
timestamp 0
transform -1 0 10850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2131_
timestamp 0
transform -1 0 7890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2132_
timestamp 0
transform 1 0 6670 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2133_
timestamp 0
transform -1 0 6970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2134_
timestamp 0
transform -1 0 7230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2135_
timestamp 0
transform -1 0 11110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2136_
timestamp 0
transform -1 0 11270 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2137_
timestamp 0
transform 1 0 11250 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2138_
timestamp 0
transform 1 0 11330 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2139_
timestamp 0
transform -1 0 11250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2140_
timestamp 0
transform -1 0 10970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2141_
timestamp 0
transform 1 0 9890 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2142_
timestamp 0
transform 1 0 10690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2143_
timestamp 0
transform -1 0 10430 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2144_
timestamp 0
transform -1 0 10990 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2145_
timestamp 0
transform -1 0 4990 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2146_
timestamp 0
transform 1 0 9710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2147_
timestamp 0
transform 1 0 10270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2148_
timestamp 0
transform -1 0 6210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2149_
timestamp 0
transform 1 0 9990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2150_
timestamp 0
transform 1 0 8770 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2151_
timestamp 0
transform 1 0 7390 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2152_
timestamp 0
transform 1 0 8470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2153_
timestamp 0
transform 1 0 8730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2154_
timestamp 0
transform 1 0 9010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2155_
timestamp 0
transform -1 0 10090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2156_
timestamp 0
transform -1 0 10870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2157_
timestamp 0
transform 1 0 11110 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2158_
timestamp 0
transform -1 0 11690 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2159_
timestamp 0
transform -1 0 11810 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2160_
timestamp 0
transform -1 0 11350 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2161_
timestamp 0
transform 1 0 8090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2162_
timestamp 0
transform 1 0 8850 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2163_
timestamp 0
transform -1 0 9950 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2164_
timestamp 0
transform 1 0 9710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2165_
timestamp 0
transform 1 0 10950 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2166_
timestamp 0
transform 1 0 10770 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2167_
timestamp 0
transform 1 0 9150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2168_
timestamp 0
transform 1 0 9970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2169_
timestamp 0
transform -1 0 8710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2170_
timestamp 0
transform -1 0 9130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2171_
timestamp 0
transform 1 0 10270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2172_
timestamp 0
transform 1 0 9690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2173_
timestamp 0
transform 1 0 9810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2174_
timestamp 0
transform -1 0 9450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2175_
timestamp 0
transform 1 0 9530 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2176_
timestamp 0
transform -1 0 9650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2177_
timestamp 0
transform -1 0 9350 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2178_
timestamp 0
transform -1 0 10950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2179_
timestamp 0
transform 1 0 9430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2180_
timestamp 0
transform 1 0 11790 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2181_
timestamp 0
transform 1 0 11770 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2182_
timestamp 0
transform 1 0 11850 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2183_
timestamp 0
transform -1 0 11230 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2184_
timestamp 0
transform 1 0 10970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2185_
timestamp 0
transform -1 0 10210 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2186_
timestamp 0
transform 1 0 10150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2187_
timestamp 0
transform -1 0 10550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2188_
timestamp 0
transform 1 0 11510 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2189_
timestamp 0
transform 1 0 9890 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2190_
timestamp 0
transform 1 0 10450 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2191_
timestamp 0
transform 1 0 11070 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2192_
timestamp 0
transform 1 0 11010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2193_
timestamp 0
transform -1 0 10950 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2194_
timestamp 0
transform -1 0 10510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2195_
timestamp 0
transform -1 0 9390 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2196_
timestamp 0
transform -1 0 11030 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2197_
timestamp 0
transform 1 0 11290 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2198_
timestamp 0
transform -1 0 9830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2199_
timestamp 0
transform -1 0 9890 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2200_
timestamp 0
transform -1 0 5750 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2201_
timestamp 0
transform 1 0 6270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2202_
timestamp 0
transform 1 0 6010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2203_
timestamp 0
transform 1 0 6010 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2204_
timestamp 0
transform 1 0 6750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2205_
timestamp 0
transform 1 0 7050 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2206_
timestamp 0
transform 1 0 9390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2207_
timestamp 0
transform -1 0 9890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2208_
timestamp 0
transform -1 0 9310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2209_
timestamp 0
transform 1 0 10350 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2210_
timestamp 0
transform 1 0 10350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2211_
timestamp 0
transform 1 0 11190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2212_
timestamp 0
transform -1 0 11550 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2213_
timestamp 0
transform -1 0 11590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2214_
timestamp 0
transform 1 0 11550 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2215_
timestamp 0
transform 1 0 11650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2216_
timestamp 0
transform 1 0 12030 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2217_
timestamp 0
transform 1 0 11310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2218_
timestamp 0
transform 1 0 9590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2219_
timestamp 0
transform -1 0 9830 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2220_
timestamp 0
transform -1 0 9870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2221_
timestamp 0
transform -1 0 11810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2222_
timestamp 0
transform 1 0 11750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2223_
timestamp 0
transform -1 0 11790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2224_
timestamp 0
transform 1 0 11770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2225_
timestamp 0
transform 1 0 10870 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2226_
timestamp 0
transform 1 0 11830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2227_
timestamp 0
transform 1 0 11550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2228_
timestamp 0
transform -1 0 11410 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2229_
timestamp 0
transform -1 0 10490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2230_
timestamp 0
transform -1 0 10210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2231_
timestamp 0
transform -1 0 8410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2232_
timestamp 0
transform 1 0 8650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2233_
timestamp 0
transform 1 0 9430 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2234_
timestamp 0
transform -1 0 9690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2235_
timestamp 0
transform -1 0 9810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2236_
timestamp 0
transform 1 0 7110 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2237_
timestamp 0
transform -1 0 6590 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2238_
timestamp 0
transform -1 0 6870 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2239_
timestamp 0
transform -1 0 8890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2240_
timestamp 0
transform -1 0 8610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2241_
timestamp 0
transform -1 0 8250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2242_
timestamp 0
transform -1 0 7430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2243_
timestamp 0
transform 1 0 7690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2244_
timestamp 0
transform 1 0 7970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2245_
timestamp 0
transform -1 0 7670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2246_
timestamp 0
transform 1 0 9050 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2247_
timestamp 0
transform -1 0 12050 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2248_
timestamp 0
transform 1 0 11250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2249_
timestamp 0
transform -1 0 9410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2250_
timestamp 0
transform 1 0 10930 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2251_
timestamp 0
transform 1 0 10490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2252_
timestamp 0
transform 1 0 11230 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2253_
timestamp 0
transform -1 0 11830 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2254_
timestamp 0
transform 1 0 12070 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2255_
timestamp 0
transform -1 0 10430 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2256_
timestamp 0
transform -1 0 10710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2257_
timestamp 0
transform 1 0 10950 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2258_
timestamp 0
transform 1 0 12110 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2259_
timestamp 0
transform -1 0 11790 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2260_
timestamp 0
transform 1 0 9970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2261_
timestamp 0
transform 1 0 10230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2262_
timestamp 0
transform -1 0 10750 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2263_
timestamp 0
transform 1 0 11230 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2264_
timestamp 0
transform 1 0 12050 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2265_
timestamp 0
transform -1 0 11310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2266_
timestamp 0
transform -1 0 10670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2267_
timestamp 0
transform 1 0 11890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2268_
timestamp 0
transform 1 0 12050 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2269_
timestamp 0
transform -1 0 11830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2270_
timestamp 0
transform 1 0 11250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2271_
timestamp 0
transform -1 0 11550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2272_
timestamp 0
transform 1 0 11810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2273_
timestamp 0
transform -1 0 12070 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2274_
timestamp 0
transform 1 0 9990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2275_
timestamp 0
transform -1 0 8150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2276_
timestamp 0
transform 1 0 8810 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2277_
timestamp 0
transform 1 0 9090 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2278_
timestamp 0
transform -1 0 9170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2279_
timestamp 0
transform 1 0 8970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2280_
timestamp 0
transform 1 0 10130 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2281_
timestamp 0
transform 1 0 12010 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2282_
timestamp 0
transform 1 0 12070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2283_
timestamp 0
transform -1 0 10950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2284_
timestamp 0
transform 1 0 12030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2285_
timestamp 0
transform 1 0 12030 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2286_
timestamp 0
transform -1 0 11810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2287_
timestamp 0
transform 1 0 11750 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2288_
timestamp 0
transform -1 0 10910 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2289_
timestamp 0
transform -1 0 10690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2290_
timestamp 0
transform -1 0 10870 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2291_
timestamp 0
transform 1 0 11230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2292_
timestamp 0
transform 1 0 10370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2293_
timestamp 0
transform 1 0 10650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2294_
timestamp 0
transform 1 0 10970 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2295_
timestamp 0
transform 1 0 10850 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2296_
timestamp 0
transform 1 0 11110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2297_
timestamp 0
transform 1 0 11770 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2298_
timestamp 0
transform -1 0 11870 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2299_
timestamp 0
transform -1 0 10430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2300_
timestamp 0
transform 1 0 10130 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2301_
timestamp 0
transform 1 0 11750 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2302_
timestamp 0
transform 1 0 11690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2303_
timestamp 0
transform -1 0 11670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2304_
timestamp 0
transform 1 0 11810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2305_
timestamp 0
transform 1 0 10690 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2306_
timestamp 0
transform -1 0 11550 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2307_
timestamp 0
transform 1 0 11250 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2308_
timestamp 0
transform 1 0 12030 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2309_
timestamp 0
transform -1 0 11590 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2310_
timestamp 0
transform -1 0 11530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2311_
timestamp 0
transform 1 0 11510 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2312_
timestamp 0
transform 1 0 11570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2313_
timestamp 0
transform 1 0 11850 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2314_
timestamp 0
transform -1 0 11170 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2315_
timestamp 0
transform 1 0 12030 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2316_
timestamp 0
transform 1 0 11430 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2317_
timestamp 0
transform -1 0 11930 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2318_
timestamp 0
transform 1 0 11470 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2319_
timestamp 0
transform 1 0 11110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2320_
timestamp 0
transform 1 0 11530 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2321_
timestamp 0
transform 1 0 11390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2322_
timestamp 0
transform -1 0 11250 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2323_
timestamp 0
transform -1 0 11490 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2324_
timestamp 0
transform 1 0 11730 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2325_
timestamp 0
transform -1 0 12110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2326_
timestamp 0
transform 1 0 12030 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2327_
timestamp 0
transform 1 0 11390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2328_
timestamp 0
transform 1 0 10970 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2329_
timestamp 0
transform 1 0 8490 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2330_
timestamp 0
transform -1 0 10170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2331_
timestamp 0
transform -1 0 9610 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2332_
timestamp 0
transform -1 0 11830 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2333_
timestamp 0
transform -1 0 10710 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2334_
timestamp 0
transform 1 0 10430 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2335_
timestamp 0
transform 1 0 10410 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2336_
timestamp 0
transform 1 0 10590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2337_
timestamp 0
transform -1 0 10710 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2338_
timestamp 0
transform -1 0 10630 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2339_
timestamp 0
transform -1 0 9550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2340_
timestamp 0
transform -1 0 9830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2341_
timestamp 0
transform 1 0 9530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2342_
timestamp 0
transform -1 0 10410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2343_
timestamp 0
transform -1 0 10350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2344_
timestamp 0
transform -1 0 10590 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2345_
timestamp 0
transform 1 0 11710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2346_
timestamp 0
transform 1 0 11450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2347_
timestamp 0
transform -1 0 8790 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2348_
timestamp 0
transform -1 0 9890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2349_
timestamp 0
transform -1 0 11550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2350_
timestamp 0
transform -1 0 11270 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2351_
timestamp 0
transform -1 0 10330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2352_
timestamp 0
transform -1 0 10090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2353_
timestamp 0
transform -1 0 9390 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2354_
timestamp 0
transform 1 0 7790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2355_
timestamp 0
transform -1 0 6870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2356_
timestamp 0
transform -1 0 6810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2357_
timestamp 0
transform -1 0 7470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2358_
timestamp 0
transform -1 0 7050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2359_
timestamp 0
transform 1 0 7270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2360_
timestamp 0
transform -1 0 7950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2361_
timestamp 0
transform -1 0 7010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2362_
timestamp 0
transform 1 0 8730 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2363_
timestamp 0
transform -1 0 7410 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2364_
timestamp 0
transform 1 0 7150 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2365_
timestamp 0
transform 1 0 6870 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2366_
timestamp 0
transform 1 0 6350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2367_
timestamp 0
transform -1 0 7190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2368_
timestamp 0
transform 1 0 6590 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2369_
timestamp 0
transform 1 0 6970 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2370_
timestamp 0
transform -1 0 7230 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2371_
timestamp 0
transform 1 0 7170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2372_
timestamp 0
transform -1 0 6750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2373_
timestamp 0
transform 1 0 6690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2374_
timestamp 0
transform 1 0 8190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2375_
timestamp 0
transform 1 0 8250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2376_
timestamp 0
transform -1 0 6690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2377_
timestamp 0
transform 1 0 5390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2378_
timestamp 0
transform -1 0 3710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2379_
timestamp 0
transform -1 0 7970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2380_
timestamp 0
transform -1 0 5610 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2381_
timestamp 0
transform -1 0 5890 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2382_
timestamp 0
transform -1 0 5750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2383_
timestamp 0
transform 1 0 4670 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2384_
timestamp 0
transform 1 0 4590 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2385_
timestamp 0
transform 1 0 4830 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2386_
timestamp 0
transform 1 0 5110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2387_
timestamp 0
transform 1 0 1630 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2388_
timestamp 0
transform 1 0 1570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2389_
timestamp 0
transform 1 0 5150 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2390_
timestamp 0
transform 1 0 2430 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2391_
timestamp 0
transform -1 0 2230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2392_
timestamp 0
transform -1 0 1950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2393_
timestamp 0
transform -1 0 2510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2394_
timestamp 0
transform -1 0 2930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2395_
timestamp 0
transform 1 0 4330 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2396_
timestamp 0
transform 1 0 2970 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2397_
timestamp 0
transform -1 0 3050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2398_
timestamp 0
transform -1 0 2770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2399_
timestamp 0
transform 1 0 1870 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2400_
timestamp 0
transform -1 0 1310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2401_
timestamp 0
transform -1 0 2790 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2402_
timestamp 0
transform 1 0 2530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2403_
timestamp 0
transform -1 0 2170 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2404_
timestamp 0
transform -1 0 1610 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2405_
timestamp 0
transform -1 0 1470 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2406_
timestamp 0
transform 1 0 5850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2407_
timestamp 0
transform -1 0 4210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2408_
timestamp 0
transform -1 0 5570 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2409_
timestamp 0
transform -1 0 6390 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2410_
timestamp 0
transform -1 0 4170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2411_
timestamp 0
transform -1 0 3930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2412_
timestamp 0
transform -1 0 1190 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2413_
timestamp 0
transform -1 0 4470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2414_
timestamp 0
transform 1 0 2990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2415_
timestamp 0
transform -1 0 2730 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2416_
timestamp 0
transform 1 0 1690 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2417_
timestamp 0
transform -1 0 2190 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2418_
timestamp 0
transform -1 0 2070 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2419_
timestamp 0
transform -1 0 3390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2420_
timestamp 0
transform 1 0 2810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2421_
timestamp 0
transform -1 0 2730 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2422_
timestamp 0
transform -1 0 1910 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2423_
timestamp 0
transform -1 0 3610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2424_
timestamp 0
transform -1 0 3450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2425_
timestamp 0
transform -1 0 3330 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2426_
timestamp 0
transform 1 0 3090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2427_
timestamp 0
transform 1 0 3250 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2428_
timestamp 0
transform -1 0 3330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2429_
timestamp 0
transform -1 0 5050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2430_
timestamp 0
transform -1 0 7750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2431_
timestamp 0
transform -1 0 5310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2432_
timestamp 0
transform -1 0 9430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2433_
timestamp 0
transform 1 0 11530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2434_
timestamp 0
transform 1 0 10710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2435_
timestamp 0
transform -1 0 7190 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2436_
timestamp 0
transform -1 0 6870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2437_
timestamp 0
transform -1 0 9550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2438_
timestamp 0
transform -1 0 9290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2439_
timestamp 0
transform -1 0 6070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2440_
timestamp 0
transform 1 0 7690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2441_
timestamp 0
transform -1 0 7530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2442_
timestamp 0
transform 1 0 10230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2443_
timestamp 0
transform -1 0 7130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2444_
timestamp 0
transform -1 0 7130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2445_
timestamp 0
transform 1 0 5230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2446_
timestamp 0
transform 1 0 6350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2447_
timestamp 0
transform -1 0 4730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2448_
timestamp 0
transform -1 0 6330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2449_
timestamp 0
transform -1 0 6950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2450_
timestamp 0
transform 1 0 4090 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2451_
timestamp 0
transform -1 0 3970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2452_
timestamp 0
transform 1 0 4610 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2453_
timestamp 0
transform 1 0 8470 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2454_
timestamp 0
transform 1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2455_
timestamp 0
transform 1 0 4350 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2456_
timestamp 0
transform -1 0 4210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2457_
timestamp 0
transform -1 0 4470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2458_
timestamp 0
transform -1 0 4830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2459_
timestamp 0
transform 1 0 4970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2460_
timestamp 0
transform 1 0 4850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2461_
timestamp 0
transform 1 0 5130 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2462_
timestamp 0
transform 1 0 5270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2463_
timestamp 0
transform 1 0 6210 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2464_
timestamp 0
transform -1 0 3150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2465_
timestamp 0
transform -1 0 2870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2466_
timestamp 0
transform -1 0 2870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2467_
timestamp 0
transform 1 0 2010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2468_
timestamp 0
transform -1 0 1570 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2469_
timestamp 0
transform 1 0 530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2470_
timestamp 0
transform -1 0 2630 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2471_
timestamp 0
transform -1 0 2650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2472_
timestamp 0
transform -1 0 2350 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2473_
timestamp 0
transform 1 0 1850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2474_
timestamp 0
transform -1 0 1370 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2475_
timestamp 0
transform -1 0 310 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2476_
timestamp 0
transform -1 0 3730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2477_
timestamp 0
transform -1 0 4970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2478_
timestamp 0
transform 1 0 3830 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2479_
timestamp 0
transform -1 0 3470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2480_
timestamp 0
transform 1 0 1710 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2481_
timestamp 0
transform -1 0 3270 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2482_
timestamp 0
transform 1 0 3550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2483_
timestamp 0
transform 1 0 2970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2484_
timestamp 0
transform 1 0 2690 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2485_
timestamp 0
transform -1 0 310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2486_
timestamp 0
transform -1 0 2590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2487_
timestamp 0
transform 1 0 2310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2488_
timestamp 0
transform -1 0 2310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2489_
timestamp 0
transform -1 0 1750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2490_
timestamp 0
transform -1 0 1310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2491_
timestamp 0
transform -1 0 310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2492_
timestamp 0
transform 1 0 4530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2493_
timestamp 0
transform 1 0 3530 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2494_
timestamp 0
transform 1 0 6110 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2495_
timestamp 0
transform 1 0 3770 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2496_
timestamp 0
transform 1 0 4070 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2497_
timestamp 0
transform -1 0 3990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2498_
timestamp 0
transform 1 0 3450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2499_
timestamp 0
transform 1 0 3710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2500_
timestamp 0
transform -1 0 310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2501_
timestamp 0
transform -1 0 3310 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2502_
timestamp 0
transform -1 0 2950 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2503_
timestamp 0
transform -1 0 3430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__2504_
timestamp 0
transform -1 0 3190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__2505_
timestamp 0
transform 1 0 2630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2506_
timestamp 0
transform -1 0 2450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__2507_
timestamp 0
transform 1 0 570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2508_
timestamp 0
transform 1 0 3070 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2509_
timestamp 0
transform 1 0 2610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2510_
timestamp 0
transform -1 0 3170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2511_
timestamp 0
transform 1 0 3250 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__2512_
timestamp 0
transform 1 0 3090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2513_
timestamp 0
transform -1 0 2350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2514_
timestamp 0
transform 1 0 2050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2515_
timestamp 0
transform -1 0 2070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2516_
timestamp 0
transform -1 0 310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__2517_
timestamp 0
transform -1 0 2150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2518_
timestamp 0
transform 1 0 5250 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2519_
timestamp 0
transform -1 0 5790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2520_
timestamp 0
transform -1 0 5890 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2521_
timestamp 0
transform 1 0 5590 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2522_
timestamp 0
transform -1 0 5590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2523_
timestamp 0
transform -1 0 5510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2524_
timestamp 0
transform -1 0 5450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2525_
timestamp 0
transform -1 0 2670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2526_
timestamp 0
transform 1 0 6070 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2527_
timestamp 0
transform 1 0 6470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2528_
timestamp 0
transform 1 0 6450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2529_
timestamp 0
transform 1 0 6050 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2530_
timestamp 0
transform 1 0 5510 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2531_
timestamp 0
transform 1 0 2870 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2532_
timestamp 0
transform 1 0 4150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2533_
timestamp 0
transform 1 0 5090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2534_
timestamp 0
transform 1 0 4810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2535_
timestamp 0
transform -1 0 4550 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2536_
timestamp 0
transform 1 0 3390 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2537_
timestamp 0
transform 1 0 2030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2538_
timestamp 0
transform 1 0 4430 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2539_
timestamp 0
transform 1 0 3810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2540_
timestamp 0
transform 1 0 4150 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2541_
timestamp 0
transform -1 0 4130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2542_
timestamp 0
transform -1 0 3650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2543_
timestamp 0
transform 1 0 3410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2544_
timestamp 0
transform 1 0 4130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2545_
timestamp 0
transform 1 0 4390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2546_
timestamp 0
transform 1 0 4750 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2547_
timestamp 0
transform -1 0 4690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2548_
timestamp 0
transform -1 0 4410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2549_
timestamp 0
transform 1 0 4630 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2550_
timestamp 0
transform 1 0 4630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2551_
timestamp 0
transform 1 0 5150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2552_
timestamp 0
transform 1 0 5390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2553_
timestamp 0
transform 1 0 2290 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2554_
timestamp 0
transform 1 0 4430 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2555_
timestamp 0
transform -1 0 4610 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2556_
timestamp 0
transform -1 0 4850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2557_
timestamp 0
transform 1 0 4550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2558_
timestamp 0
transform 1 0 4630 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2559_
timestamp 0
transform 1 0 4350 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2560_
timestamp 0
transform 1 0 3850 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2561_
timestamp 0
transform 1 0 3550 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2562_
timestamp 0
transform 1 0 2170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2563_
timestamp 0
transform -1 0 4390 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2564_
timestamp 0
transform 1 0 4310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2565_
timestamp 0
transform -1 0 3790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2566_
timestamp 0
transform 1 0 2390 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2567_
timestamp 0
transform 1 0 3870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2568_
timestamp 0
transform -1 0 5670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2569_
timestamp 0
transform -1 0 5810 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2570_
timestamp 0
transform 1 0 5890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2571_
timestamp 0
transform 1 0 5890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2572_
timestamp 0
transform 1 0 5750 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2573_
timestamp 0
transform 1 0 5670 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2574_
timestamp 0
transform 1 0 5650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2575_
timestamp 0
transform -1 0 4690 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2576_
timestamp 0
transform -1 0 4170 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2577_
timestamp 0
transform -1 0 4430 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2578_
timestamp 0
transform 1 0 6930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2579_
timestamp 0
transform 1 0 6950 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2580_
timestamp 0
transform 1 0 7950 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2581_
timestamp 0
transform -1 0 8810 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2582_
timestamp 0
transform 1 0 6850 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2583_
timestamp 0
transform -1 0 6850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2584_
timestamp 0
transform 1 0 7270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2585_
timestamp 0
transform 1 0 7310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2586_
timestamp 0
transform -1 0 8390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2587_
timestamp 0
transform -1 0 6730 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2588_
timestamp 0
transform -1 0 5770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2589_
timestamp 0
transform 1 0 7390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2590_
timestamp 0
transform -1 0 6170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2591_
timestamp 0
transform 1 0 6410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2592_
timestamp 0
transform -1 0 4390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2593_
timestamp 0
transform 1 0 4910 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2594_
timestamp 0
transform -1 0 8490 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2595_
timestamp 0
transform -1 0 5210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2596_
timestamp 0
transform 1 0 5210 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2597_
timestamp 0
transform 1 0 5390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2598_
timestamp 0
transform -1 0 5130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2599_
timestamp 0
transform -1 0 4930 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2600_
timestamp 0
transform -1 0 4930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2601_
timestamp 0
transform -1 0 5190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2602_
timestamp 0
transform -1 0 8130 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2603_
timestamp 0
transform -1 0 6570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2604_
timestamp 0
transform -1 0 6330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2605_
timestamp 0
transform 1 0 6010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2606_
timestamp 0
transform -1 0 5510 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2607_
timestamp 0
transform 1 0 5670 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2608_
timestamp 0
transform 1 0 5490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2609_
timestamp 0
transform -1 0 5470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2610_
timestamp 0
transform 1 0 4850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2611_
timestamp 0
transform -1 0 5110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2612_
timestamp 0
transform -1 0 5370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2613_
timestamp 0
transform -1 0 1190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2614_
timestamp 0
transform 1 0 2170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2615_
timestamp 0
transform -1 0 2450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2616_
timestamp 0
transform -1 0 2430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2617_
timestamp 0
transform 1 0 1410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2618_
timestamp 0
transform 1 0 830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2619_
timestamp 0
transform -1 0 330 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2620_
timestamp 0
transform -1 0 570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2621_
timestamp 0
transform 1 0 890 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2622_
timestamp 0
transform 1 0 330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2623_
timestamp 0
transform 1 0 2710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2624_
timestamp 0
transform 1 0 1910 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2625_
timestamp 0
transform -1 0 2170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2626_
timestamp 0
transform -1 0 1890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2627_
timestamp 0
transform 1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2628_
timestamp 0
transform 1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2629_
timestamp 0
transform -1 0 290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2630_
timestamp 0
transform 1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2631_
timestamp 0
transform 1 0 4970 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2632_
timestamp 0
transform 1 0 2210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2633_
timestamp 0
transform -1 0 2510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2634_
timestamp 0
transform -1 0 50 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2635_
timestamp 0
transform 1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2636_
timestamp 0
transform 1 0 570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2637_
timestamp 0
transform 1 0 910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2638_
timestamp 0
transform 1 0 330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2639_
timestamp 0
transform -1 0 650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2640_
timestamp 0
transform -1 0 50 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2641_
timestamp 0
transform -1 0 50 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2642_
timestamp 0
transform 1 0 1290 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2643_
timestamp 0
transform -1 0 1830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2644_
timestamp 0
transform 1 0 2230 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2645_
timestamp 0
transform -1 0 1970 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2646_
timestamp 0
transform -1 0 1170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2647_
timestamp 0
transform 1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2648_
timestamp 0
transform 1 0 530 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__2649_
timestamp 0
transform 1 0 30 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2650_
timestamp 0
transform -1 0 3630 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2651_
timestamp 0
transform -1 0 3350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2652_
timestamp 0
transform 1 0 570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2653_
timestamp 0
transform 1 0 290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2654_
timestamp 0
transform 1 0 1170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2655_
timestamp 0
transform 1 0 610 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2656_
timestamp 0
transform -1 0 890 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2657_
timestamp 0
transform 1 0 30 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2658_
timestamp 0
transform 1 0 30 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2659_
timestamp 0
transform -1 0 330 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2660_
timestamp 0
transform 1 0 270 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2661_
timestamp 0
transform -1 0 2590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__2662_
timestamp 0
transform -1 0 2530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2663_
timestamp 0
transform -1 0 1950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2664_
timestamp 0
transform 1 0 850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2665_
timestamp 0
transform -1 0 810 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2666_
timestamp 0
transform -1 0 330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2667_
timestamp 0
transform -1 0 550 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2668_
timestamp 0
transform 1 0 1050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2669_
timestamp 0
transform -1 0 2810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2670_
timestamp 0
transform -1 0 2930 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2671_
timestamp 0
transform 1 0 1090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2672_
timestamp 0
transform -1 0 590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2673_
timestamp 0
transform -1 0 550 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2674_
timestamp 0
transform 1 0 810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2675_
timestamp 0
transform 1 0 790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2676_
timestamp 0
transform -1 0 1090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2677_
timestamp 0
transform 1 0 6430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__2678_
timestamp 0
transform -1 0 6350 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2679_
timestamp 0
transform 1 0 6970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2680_
timestamp 0
transform -1 0 6770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2681_
timestamp 0
transform 1 0 7030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2682_
timestamp 0
transform -1 0 6750 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2683_
timestamp 0
transform -1 0 1870 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2684_
timestamp 0
transform -1 0 1690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__2685_
timestamp 0
transform 1 0 1610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2686_
timestamp 0
transform 1 0 1610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2687_
timestamp 0
transform 1 0 1350 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2688_
timestamp 0
transform -1 0 790 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2689_
timestamp 0
transform -1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2690_
timestamp 0
transform 1 0 7270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2691_
timestamp 0
transform -1 0 7110 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2692_
timestamp 0
transform -1 0 5050 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2693_
timestamp 0
transform -1 0 3010 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2694_
timestamp 0
transform -1 0 1310 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2695_
timestamp 0
transform -1 0 1590 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2696_
timestamp 0
transform -1 0 1310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2697_
timestamp 0
transform 1 0 1890 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2698_
timestamp 0
transform -1 0 530 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2699_
timestamp 0
transform 1 0 6290 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2700_
timestamp 0
transform -1 0 7010 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2701_
timestamp 0
transform 1 0 7590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2702_
timestamp 0
transform 1 0 7290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2703_
timestamp 0
transform 1 0 7450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2704_
timestamp 0
transform -1 0 6650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2705_
timestamp 0
transform 1 0 1570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2706_
timestamp 0
transform 1 0 1010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2707_
timestamp 0
transform 1 0 2710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2708_
timestamp 0
transform 1 0 2390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2709_
timestamp 0
transform -1 0 1070 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2710_
timestamp 0
transform -1 0 850 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2711_
timestamp 0
transform -1 0 1130 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2712_
timestamp 0
transform 1 0 2870 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2713_
timestamp 0
transform -1 0 4270 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2714_
timestamp 0
transform -1 0 4690 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2715_
timestamp 0
transform 1 0 3530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2716_
timestamp 0
transform -1 0 4290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2717_
timestamp 0
transform -1 0 5850 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__2718_
timestamp 0
transform -1 0 4090 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2719_
timestamp 0
transform 1 0 3690 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2720_
timestamp 0
transform -1 0 3990 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2721_
timestamp 0
transform -1 0 2150 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2722_
timestamp 0
transform 1 0 2270 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2723_
timestamp 0
transform 1 0 2570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2724_
timestamp 0
transform -1 0 810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2725_
timestamp 0
transform -1 0 5410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2726_
timestamp 0
transform -1 0 6590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2727_
timestamp 0
transform 1 0 3850 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2728_
timestamp 0
transform 1 0 3570 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2729_
timestamp 0
transform -1 0 3530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2730_
timestamp 0
transform 1 0 3130 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2731_
timestamp 0
transform 1 0 1990 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2732_
timestamp 0
transform -1 0 1870 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2733_
timestamp 0
transform 1 0 1410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2734_
timestamp 0
transform -1 0 1710 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2735_
timestamp 0
transform -1 0 3870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2736_
timestamp 0
transform -1 0 4010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2737_
timestamp 0
transform -1 0 4090 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2738_
timestamp 0
transform -1 0 3790 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2739_
timestamp 0
transform -1 0 3230 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2740_
timestamp 0
transform -1 0 3310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2741_
timestamp 0
transform -1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2742_
timestamp 0
transform 1 0 1370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2743_
timestamp 0
transform 1 0 1310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2744_
timestamp 0
transform 1 0 1850 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2745_
timestamp 0
transform 1 0 510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2746_
timestamp 0
transform 1 0 3570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2747_
timestamp 0
transform 1 0 4690 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__2748_
timestamp 0
transform 1 0 4350 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2749_
timestamp 0
transform -1 0 3510 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2750_
timestamp 0
transform -1 0 2950 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2751_
timestamp 0
transform 1 0 2790 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2752_
timestamp 0
transform 1 0 1090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2753_
timestamp 0
transform 1 0 590 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2754_
timestamp 0
transform -1 0 530 0 1 790
box -6 -8 26 268
use FILL  FILL_1__2755_
timestamp 0
transform -1 0 3050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2756_
timestamp 0
transform -1 0 2490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2757_
timestamp 0
transform 1 0 2730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2758_
timestamp 0
transform 1 0 2210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2759_
timestamp 0
transform -1 0 4290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2760_
timestamp 0
transform 1 0 3730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2761_
timestamp 0
transform 1 0 4070 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2762_
timestamp 0
transform -1 0 3810 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2763_
timestamp 0
transform -1 0 2050 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2764_
timestamp 0
transform -1 0 1770 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2765_
timestamp 0
transform -1 0 1690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2766_
timestamp 0
transform -1 0 1950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__2767_
timestamp 0
transform -1 0 1470 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__2768_
timestamp 0
transform 1 0 2130 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2769_
timestamp 0
transform 1 0 1570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__2770_
timestamp 0
transform 1 0 5930 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2771_
timestamp 0
transform 1 0 6470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2772_
timestamp 0
transform 1 0 4910 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__2773_
timestamp 0
transform 1 0 4110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2774_
timestamp 0
transform 1 0 2270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2775_
timestamp 0
transform 1 0 2510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2776_
timestamp 0
transform 1 0 3330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2777_
timestamp 0
transform -1 0 2810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2778_
timestamp 0
transform -1 0 3070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__2779_
timestamp 0
transform -1 0 7110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2780_
timestamp 0
transform -1 0 7350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__2781_
timestamp 0
transform 1 0 7830 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__2782_
timestamp 0
transform 1 0 7710 0 1 270
box -6 -8 26 268
use FILL  FILL_1__2783_
timestamp 0
transform 1 0 9650 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2784_
timestamp 0
transform 1 0 10790 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2785_
timestamp 0
transform 1 0 10170 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2786_
timestamp 0
transform 1 0 9890 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2787_
timestamp 0
transform 1 0 8350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2788_
timestamp 0
transform 1 0 8610 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2789_
timestamp 0
transform 1 0 8130 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2790_
timestamp 0
transform -1 0 7870 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2791_
timestamp 0
transform 1 0 6130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2792_
timestamp 0
transform 1 0 9750 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2793_
timestamp 0
transform 1 0 9950 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2794_
timestamp 0
transform -1 0 10210 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2795_
timestamp 0
transform 1 0 8390 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2796_
timestamp 0
transform 1 0 8370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2797_
timestamp 0
transform 1 0 10770 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2798_
timestamp 0
transform -1 0 9910 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2799_
timestamp 0
transform -1 0 8290 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2800_
timestamp 0
transform -1 0 7690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2801_
timestamp 0
transform 1 0 9630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2802_
timestamp 0
transform -1 0 9950 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2803_
timestamp 0
transform 1 0 8390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2804_
timestamp 0
transform -1 0 8290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2805_
timestamp 0
transform -1 0 10030 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2806_
timestamp 0
transform 1 0 9710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2807_
timestamp 0
transform -1 0 8330 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2808_
timestamp 0
transform -1 0 6570 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2809_
timestamp 0
transform 1 0 8090 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2810_
timestamp 0
transform -1 0 7510 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2811_
timestamp 0
transform 1 0 9990 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2812_
timestamp 0
transform 1 0 9630 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2813_
timestamp 0
transform 1 0 8210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2814_
timestamp 0
transform -1 0 8090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2815_
timestamp 0
transform -1 0 8170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2816_
timestamp 0
transform 1 0 9430 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2817_
timestamp 0
transform -1 0 10290 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2818_
timestamp 0
transform 1 0 11110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2819_
timestamp 0
transform 1 0 10090 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2820_
timestamp 0
transform -1 0 9870 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2821_
timestamp 0
transform -1 0 9730 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2822_
timestamp 0
transform -1 0 7450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2823_
timestamp 0
transform -1 0 9450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2824_
timestamp 0
transform -1 0 9190 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2825_
timestamp 0
transform 1 0 8650 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2826_
timestamp 0
transform 1 0 8690 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2827_
timestamp 0
transform 1 0 9110 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2828_
timestamp 0
transform 1 0 10230 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2829_
timestamp 0
transform -1 0 9170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2830_
timestamp 0
transform 1 0 9790 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2831_
timestamp 0
transform 1 0 8970 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2832_
timestamp 0
transform -1 0 8890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2833_
timestamp 0
transform -1 0 8650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2834_
timestamp 0
transform -1 0 8230 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2835_
timestamp 0
transform -1 0 9250 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2836_
timestamp 0
transform -1 0 7950 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2837_
timestamp 0
transform 1 0 8030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2838_
timestamp 0
transform 1 0 9270 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2839_
timestamp 0
transform 1 0 9530 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2840_
timestamp 0
transform -1 0 9270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2841_
timestamp 0
transform 1 0 8170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2842_
timestamp 0
transform 1 0 11490 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2843_
timestamp 0
transform -1 0 10990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2844_
timestamp 0
transform 1 0 10710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2845_
timestamp 0
transform 1 0 10450 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2846_
timestamp 0
transform -1 0 10090 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2847_
timestamp 0
transform 1 0 10290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2848_
timestamp 0
transform -1 0 9570 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2849_
timestamp 0
transform 1 0 10870 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__2850_
timestamp 0
transform 1 0 11030 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2851_
timestamp 0
transform 1 0 11270 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2852_
timestamp 0
transform 1 0 11970 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2853_
timestamp 0
transform 1 0 12030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2854_
timestamp 0
transform 1 0 11710 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2855_
timestamp 0
transform 1 0 11990 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2856_
timestamp 0
transform -1 0 9030 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2857_
timestamp 0
transform 1 0 9530 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2858_
timestamp 0
transform -1 0 9830 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2859_
timestamp 0
transform 1 0 10770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2860_
timestamp 0
transform 1 0 7650 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2861_
timestamp 0
transform 1 0 8330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2862_
timestamp 0
transform -1 0 7710 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2863_
timestamp 0
transform 1 0 7410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2864_
timestamp 0
transform 1 0 9650 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2865_
timestamp 0
transform 1 0 8810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2866_
timestamp 0
transform -1 0 6910 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2867_
timestamp 0
transform -1 0 8750 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2868_
timestamp 0
transform -1 0 8470 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2869_
timestamp 0
transform -1 0 8910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2870_
timestamp 0
transform 1 0 8550 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2871_
timestamp 0
transform 1 0 8510 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2872_
timestamp 0
transform 1 0 5450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2873_
timestamp 0
transform -1 0 5470 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2874_
timestamp 0
transform 1 0 5390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2875_
timestamp 0
transform -1 0 5750 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2876_
timestamp 0
transform 1 0 5430 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2877_
timestamp 0
transform 1 0 6010 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2878_
timestamp 0
transform -1 0 5750 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2879_
timestamp 0
transform -1 0 8890 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2880_
timestamp 0
transform -1 0 11890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2881_
timestamp 0
transform 1 0 11570 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2882_
timestamp 0
transform -1 0 9170 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2883_
timestamp 0
transform 1 0 8970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2884_
timestamp 0
transform -1 0 9290 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2885_
timestamp 0
transform -1 0 10470 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2886_
timestamp 0
transform 1 0 10430 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2887_
timestamp 0
transform -1 0 8850 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2888_
timestamp 0
transform -1 0 9130 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2889_
timestamp 0
transform 1 0 9410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2890_
timestamp 0
transform -1 0 9770 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__2891_
timestamp 0
transform -1 0 9710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2892_
timestamp 0
transform 1 0 9090 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2893_
timestamp 0
transform -1 0 9250 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2894_
timestamp 0
transform -1 0 11070 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2895_
timestamp 0
transform 1 0 10750 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2896_
timestamp 0
transform -1 0 11030 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2897_
timestamp 0
transform -1 0 10750 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2898_
timestamp 0
transform 1 0 9370 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2899_
timestamp 0
transform -1 0 9670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2900_
timestamp 0
transform 1 0 10350 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2901_
timestamp 0
transform -1 0 10370 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2902_
timestamp 0
transform 1 0 10550 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2903_
timestamp 0
transform -1 0 10670 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2904_
timestamp 0
transform -1 0 9830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2905_
timestamp 0
transform -1 0 9330 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2906_
timestamp 0
transform -1 0 8490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2907_
timestamp 0
transform -1 0 9050 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2908_
timestamp 0
transform -1 0 10390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2909_
timestamp 0
transform 1 0 11750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2910_
timestamp 0
transform 1 0 10830 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2911_
timestamp 0
transform 1 0 11690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2912_
timestamp 0
transform 1 0 11970 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__2913_
timestamp 0
transform 1 0 10570 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__2914_
timestamp 0
transform -1 0 7750 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2915_
timestamp 0
transform 1 0 10890 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2916_
timestamp 0
transform 1 0 11130 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__2917_
timestamp 0
transform 1 0 10630 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2918_
timestamp 0
transform -1 0 10790 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2919_
timestamp 0
transform 1 0 8470 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2920_
timestamp 0
transform 1 0 11170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2921_
timestamp 0
transform 1 0 11690 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__2922_
timestamp 0
transform -1 0 11810 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2923_
timestamp 0
transform 1 0 11270 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2924_
timestamp 0
transform 1 0 10190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2925_
timestamp 0
transform 1 0 9950 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2926_
timestamp 0
transform 1 0 10090 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2927_
timestamp 0
transform -1 0 9930 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2928_
timestamp 0
transform -1 0 10190 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__2929_
timestamp 0
transform -1 0 10310 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__2930_
timestamp 0
transform -1 0 11190 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2931_
timestamp 0
transform -1 0 11450 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__2932_
timestamp 0
transform 1 0 11410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__2933_
timestamp 0
transform 1 0 11370 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__2934_
timestamp 0
transform 1 0 11450 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__2935_
timestamp 0
transform 1 0 11530 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2936_
timestamp 0
transform 1 0 10470 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__2937_
timestamp 0
transform -1 0 3470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__2938_
timestamp 0
transform -1 0 7690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2939_
timestamp 0
transform 1 0 6450 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2940_
timestamp 0
transform -1 0 6230 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2941_
timestamp 0
transform -1 0 6150 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2942_
timestamp 0
transform 1 0 5050 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2943_
timestamp 0
transform -1 0 6950 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__2944_
timestamp 0
transform 1 0 5330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2945_
timestamp 0
transform -1 0 6730 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2946_
timestamp 0
transform 1 0 6330 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__2947_
timestamp 0
transform 1 0 7810 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2948_
timestamp 0
transform 1 0 7550 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2949_
timestamp 0
transform 1 0 5650 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__2950_
timestamp 0
transform -1 0 5990 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2951_
timestamp 0
transform 1 0 6750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2952_
timestamp 0
transform 1 0 6470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2953_
timestamp 0
transform 1 0 5630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2954_
timestamp 0
transform -1 0 5930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__2955_
timestamp 0
transform 1 0 7010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2956_
timestamp 0
transform 1 0 6490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__2957_
timestamp 0
transform -1 0 8110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__2958_
timestamp 0
transform 1 0 6490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__2959_
timestamp 0
transform 1 0 6230 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2960_
timestamp 0
transform -1 0 7110 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2961_
timestamp 0
transform 1 0 6490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2962_
timestamp 0
transform -1 0 6270 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__2963_
timestamp 0
transform -1 0 6570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2964_
timestamp 0
transform 1 0 4630 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2965_
timestamp 0
transform 1 0 5690 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2966_
timestamp 0
transform -1 0 6590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__2967_
timestamp 0
transform -1 0 5010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2968_
timestamp 0
transform -1 0 5270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2969_
timestamp 0
transform 1 0 4350 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2970_
timestamp 0
transform 1 0 4710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2971_
timestamp 0
transform 1 0 4590 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2972_
timestamp 0
transform -1 0 6030 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2973_
timestamp 0
transform -1 0 6290 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2974_
timestamp 0
transform -1 0 6290 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2975_
timestamp 0
transform 1 0 5750 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2976_
timestamp 0
transform -1 0 4670 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2977_
timestamp 0
transform -1 0 4930 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2978_
timestamp 0
transform 1 0 5190 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__2979_
timestamp 0
transform 1 0 5470 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__2980_
timestamp 0
transform -1 0 7350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2981_
timestamp 0
transform -1 0 6310 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2982_
timestamp 0
transform -1 0 6590 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__2983_
timestamp 0
transform 1 0 7110 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2984_
timestamp 0
transform 1 0 6510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__2985_
timestamp 0
transform -1 0 6850 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2986_
timestamp 0
transform 1 0 6550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2987_
timestamp 0
transform 1 0 5990 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2988_
timestamp 0
transform -1 0 6270 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__2989_
timestamp 0
transform -1 0 7850 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2990_
timestamp 0
transform 1 0 6970 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__2991_
timestamp 0
transform -1 0 6830 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2992_
timestamp 0
transform -1 0 5130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__2993_
timestamp 0
transform -1 0 5990 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2994_
timestamp 0
transform 1 0 5450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2995_
timestamp 0
transform 1 0 6530 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2996_
timestamp 0
transform 1 0 6250 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__2997_
timestamp 0
transform 1 0 5970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2998_
timestamp 0
transform -1 0 5710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__2999_
timestamp 0
transform 1 0 6370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3000_
timestamp 0
transform -1 0 5710 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__3001_
timestamp 0
transform 1 0 4930 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3002_
timestamp 0
transform -1 0 5430 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__3003_
timestamp 0
transform -1 0 5790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3004_
timestamp 0
transform -1 0 5210 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3005_
timestamp 0
transform -1 0 5470 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3006_
timestamp 0
transform -1 0 7370 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3007_
timestamp 0
transform 1 0 6790 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3008_
timestamp 0
transform 1 0 8590 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3009_
timestamp 0
transform 1 0 8050 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3010_
timestamp 0
transform 1 0 7070 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3011_
timestamp 0
transform -1 0 7170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3012_
timestamp 0
transform -1 0 7050 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3013_
timestamp 0
transform -1 0 7790 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3014_
timestamp 0
transform 1 0 6990 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3015_
timestamp 0
transform -1 0 7270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3016_
timestamp 0
transform -1 0 6030 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3017_
timestamp 0
transform -1 0 6830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3018_
timestamp 0
transform -1 0 6510 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3019_
timestamp 0
transform -1 0 6770 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3020_
timestamp 0
transform 1 0 5410 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__3021_
timestamp 0
transform 1 0 5850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3022_
timestamp 0
transform 1 0 5650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__3023_
timestamp 0
transform -1 0 6730 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3024_
timestamp 0
transform -1 0 6650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3025_
timestamp 0
transform 1 0 5930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__3026_
timestamp 0
transform 1 0 5350 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__3027_
timestamp 0
transform -1 0 5450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3028_
timestamp 0
transform 1 0 5930 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3029_
timestamp 0
transform 1 0 6690 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3030_
timestamp 0
transform 1 0 4830 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__3031_
timestamp 0
transform 1 0 4370 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3032_
timestamp 0
transform -1 0 5150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3033_
timestamp 0
transform 1 0 5410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3034_
timestamp 0
transform -1 0 3350 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3035_
timestamp 0
transform -1 0 3910 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3036_
timestamp 0
transform -1 0 3410 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3037_
timestamp 0
transform -1 0 3290 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3038_
timestamp 0
transform 1 0 3510 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3039_
timestamp 0
transform -1 0 3010 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3040_
timestamp 0
transform 1 0 2890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3041_
timestamp 0
transform 1 0 3130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3042_
timestamp 0
transform -1 0 3690 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3043_
timestamp 0
transform -1 0 3790 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3044_
timestamp 0
transform -1 0 3550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3045_
timestamp 0
transform 1 0 4350 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3046_
timestamp 0
transform 1 0 4070 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3047_
timestamp 0
transform -1 0 3030 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3048_
timestamp 0
transform 1 0 3070 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3049_
timestamp 0
transform -1 0 2770 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3050_
timestamp 0
transform 1 0 2810 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3051_
timestamp 0
transform 1 0 2550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3052_
timestamp 0
transform 1 0 2450 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3053_
timestamp 0
transform 1 0 3210 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3054_
timestamp 0
transform -1 0 3490 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3055_
timestamp 0
transform 1 0 3310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3056_
timestamp 0
transform -1 0 3570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3057_
timestamp 0
transform 1 0 3770 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3058_
timestamp 0
transform 1 0 3950 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3059_
timestamp 0
transform 1 0 4230 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3060_
timestamp 0
transform 1 0 4070 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3061_
timestamp 0
transform 1 0 3550 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3062_
timestamp 0
transform -1 0 3790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3063_
timestamp 0
transform -1 0 5030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__3064_
timestamp 0
transform 1 0 4890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__3065_
timestamp 0
transform -1 0 4630 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3066_
timestamp 0
transform 1 0 4530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3067_
timestamp 0
transform -1 0 3630 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3068_
timestamp 0
transform -1 0 3370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3069_
timestamp 0
transform 1 0 3570 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3070_
timestamp 0
transform -1 0 4470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__3071_
timestamp 0
transform 1 0 4190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__3072_
timestamp 0
transform -1 0 4130 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3073_
timestamp 0
transform -1 0 4390 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3074_
timestamp 0
transform 1 0 5670 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3075_
timestamp 0
transform 1 0 5390 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3076_
timestamp 0
transform 1 0 3630 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3077_
timestamp 0
transform 1 0 3950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3078_
timestamp 0
transform 1 0 4010 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3079_
timestamp 0
transform -1 0 4090 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3080_
timestamp 0
transform 1 0 6230 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3081_
timestamp 0
transform -1 0 6890 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3082_
timestamp 0
transform 1 0 6590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3083_
timestamp 0
transform -1 0 3770 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3084_
timestamp 0
transform 1 0 3470 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3085_
timestamp 0
transform 1 0 3090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3086_
timestamp 0
transform -1 0 2810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3087_
timestamp 0
transform 1 0 4290 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3088_
timestamp 0
transform -1 0 4890 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3089_
timestamp 0
transform 1 0 3370 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3090_
timestamp 0
transform -1 0 3650 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3091_
timestamp 0
transform -1 0 6190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3092_
timestamp 0
transform 1 0 5410 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3093_
timestamp 0
transform 1 0 5670 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3094_
timestamp 0
transform 1 0 5390 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3095_
timestamp 0
transform -1 0 4590 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3096_
timestamp 0
transform 1 0 4290 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3097_
timestamp 0
transform -1 0 4050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3098_
timestamp 0
transform 1 0 3750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3099_
timestamp 0
transform -1 0 3810 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3100_
timestamp 0
transform -1 0 3630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3101_
timestamp 0
transform 1 0 4850 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3102_
timestamp 0
transform -1 0 5150 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3103_
timestamp 0
transform -1 0 4530 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3104_
timestamp 0
transform -1 0 4810 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3105_
timestamp 0
transform 1 0 5590 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3106_
timestamp 0
transform -1 0 5890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3107_
timestamp 0
transform -1 0 3990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3108_
timestamp 0
transform 1 0 3690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3109_
timestamp 0
transform 1 0 6170 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3110_
timestamp 0
transform 1 0 3850 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3111_
timestamp 0
transform 1 0 5710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3112_
timestamp 0
transform -1 0 5130 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3113_
timestamp 0
transform -1 0 4590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3114_
timestamp 0
transform 1 0 4290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3115_
timestamp 0
transform 1 0 4810 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3116_
timestamp 0
transform 1 0 3750 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3117_
timestamp 0
transform 1 0 4370 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3118_
timestamp 0
transform -1 0 4670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3119_
timestamp 0
transform 1 0 4850 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3120_
timestamp 0
transform 1 0 4550 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3121_
timestamp 0
transform 1 0 5150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3122_
timestamp 0
transform 1 0 5430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3123_
timestamp 0
transform 1 0 5410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3124_
timestamp 0
transform -1 0 5710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3125_
timestamp 0
transform -1 0 4070 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3126_
timestamp 0
transform 1 0 3770 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3127_
timestamp 0
transform 1 0 6430 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3128_
timestamp 0
transform 1 0 5990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3129_
timestamp 0
transform 1 0 5390 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3130_
timestamp 0
transform -1 0 3310 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3131_
timestamp 0
transform -1 0 3550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3132_
timestamp 0
transform 1 0 4650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3133_
timestamp 0
transform 1 0 3890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3134_
timestamp 0
transform 1 0 5070 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3135_
timestamp 0
transform 1 0 4770 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3136_
timestamp 0
transform 1 0 5670 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3137_
timestamp 0
transform 1 0 5390 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3138_
timestamp 0
transform 1 0 5670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3139_
timestamp 0
transform 1 0 5390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3140_
timestamp 0
transform -1 0 5590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3141_
timestamp 0
transform -1 0 5850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3142_
timestamp 0
transform -1 0 4190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3143_
timestamp 0
transform -1 0 4450 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3144_
timestamp 0
transform 1 0 11530 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__3145_
timestamp 0
transform 1 0 11770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__3146_
timestamp 0
transform -1 0 11830 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__3147_
timestamp 0
transform 1 0 9450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__3148_
timestamp 0
transform -1 0 11830 0 1 790
box -6 -8 26 268
use FILL  FILL_1__3149_
timestamp 0
transform -1 0 11450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3150_
timestamp 0
transform -1 0 11730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3151_
timestamp 0
transform -1 0 10670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3152_
timestamp 0
transform 1 0 9310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3153_
timestamp 0
transform -1 0 9610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3154_
timestamp 0
transform -1 0 10130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3155_
timestamp 0
transform -1 0 10250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3156_
timestamp 0
transform -1 0 8890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__3157_
timestamp 0
transform -1 0 8930 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__3158_
timestamp 0
transform -1 0 8650 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__3159_
timestamp 0
transform -1 0 8630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__3160_
timestamp 0
transform 1 0 10470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3161_
timestamp 0
transform 1 0 10190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3162_
timestamp 0
transform -1 0 9730 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3163_
timestamp 0
transform 1 0 9450 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3164_
timestamp 0
transform -1 0 8930 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3165_
timestamp 0
transform -1 0 7150 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3166_
timestamp 0
transform 1 0 7550 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__3167_
timestamp 0
transform 1 0 7410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3168_
timestamp 0
transform 1 0 7570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3169_
timestamp 0
transform -1 0 8650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3170_
timestamp 0
transform -1 0 8370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3171_
timestamp 0
transform -1 0 9090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3172_
timestamp 0
transform -1 0 8090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3173_
timestamp 0
transform 1 0 8350 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3174_
timestamp 0
transform 1 0 7830 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3175_
timestamp 0
transform -1 0 7810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3176_
timestamp 0
transform -1 0 7530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3177_
timestamp 0
transform -1 0 11810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__3178_
timestamp 0
transform -1 0 11750 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3179_
timestamp 0
transform 1 0 12010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3180_
timestamp 0
transform 1 0 12070 0 1 790
box -6 -8 26 268
use FILL  FILL_1__3181_
timestamp 0
transform 1 0 12050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__3182_
timestamp 0
transform -1 0 11270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3183_
timestamp 0
transform 1 0 11530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3184_
timestamp 0
transform 1 0 11810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3185_
timestamp 0
transform 1 0 11830 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3186_
timestamp 0
transform 1 0 12010 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3187_
timestamp 0
transform 1 0 9870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__3188_
timestamp 0
transform 1 0 10750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3189_
timestamp 0
transform -1 0 11010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__3190_
timestamp 0
transform 1 0 11050 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3191_
timestamp 0
transform 1 0 10990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3192_
timestamp 0
transform -1 0 10710 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3193_
timestamp 0
transform 1 0 10130 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3194_
timestamp 0
transform 1 0 10750 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__3195_
timestamp 0
transform -1 0 10490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3196_
timestamp 0
transform 1 0 10390 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3197_
timestamp 0
transform -1 0 7250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3198_
timestamp 0
transform -1 0 4610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3199_
timestamp 0
transform 1 0 2770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__3200_
timestamp 0
transform 1 0 4750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__3201_
timestamp 0
transform 1 0 4470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__3202_
timestamp 0
transform 1 0 1530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__3203_
timestamp 0
transform 1 0 1490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3204_
timestamp 0
transform 1 0 1450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__3205_
timestamp 0
transform 1 0 1010 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__3206_
timestamp 0
transform 1 0 1430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__3207_
timestamp 0
transform -1 0 1570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__3208_
timestamp 0
transform -1 0 910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__3209_
timestamp 0
transform -1 0 610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__3210_
timestamp 0
transform -1 0 4270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__3211_
timestamp 0
transform 1 0 4210 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__3212_
timestamp 0
transform 1 0 1170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__3213_
timestamp 0
transform 1 0 1070 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__3214_
timestamp 0
transform -1 0 2350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3215_
timestamp 0
transform 1 0 1770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3216_
timestamp 0
transform 1 0 5710 0 1 270
box -6 -8 26 268
use FILL  FILL_1__3217_
timestamp 0
transform -1 0 6010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__3218_
timestamp 0
transform 1 0 6050 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3219_
timestamp 0
transform -1 0 6330 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3220_
timestamp 0
transform 1 0 3670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3221_
timestamp 0
transform -1 0 3950 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3222_
timestamp 0
transform -1 0 3550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3223_
timestamp 0
transform 1 0 3270 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__3224_
timestamp 0
transform -1 0 3250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3225_
timestamp 0
transform 1 0 5390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__3226_
timestamp 0
transform 1 0 5110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__3227_
timestamp 0
transform -1 0 4230 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3228_
timestamp 0
transform -1 0 4430 0 1 270
box -6 -8 26 268
use FILL  FILL_1__3229_
timestamp 0
transform 1 0 2670 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__3230_
timestamp 0
transform -1 0 2710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__3231_
timestamp 0
transform 1 0 5950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__3232_
timestamp 0
transform 1 0 5930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__3364_
timestamp 0
transform 1 0 5210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3365_
timestamp 0
transform 1 0 4410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3366_
timestamp 0
transform 1 0 4890 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__3367_
timestamp 0
transform -1 0 4690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3368_
timestamp 0
transform -1 0 4950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3369_
timestamp 0
transform -1 0 5510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3370_
timestamp 0
transform 1 0 2650 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3371_
timestamp 0
transform 1 0 2150 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3372_
timestamp 0
transform -1 0 2270 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3373_
timestamp 0
transform -1 0 3930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3374_
timestamp 0
transform -1 0 2250 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3375_
timestamp 0
transform 1 0 2250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3376_
timestamp 0
transform -1 0 2910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3377_
timestamp 0
transform 1 0 2370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3378_
timestamp 0
transform -1 0 2230 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3379_
timestamp 0
transform -1 0 1390 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3380_
timestamp 0
transform 1 0 1170 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3381_
timestamp 0
transform -1 0 1430 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3382_
timestamp 0
transform -1 0 1890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3383_
timestamp 0
transform -1 0 1450 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3384_
timestamp 0
transform 1 0 1710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3385_
timestamp 0
transform 1 0 1410 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3386_
timestamp 0
transform -1 0 1990 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3387_
timestamp 0
transform 1 0 2250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3388_
timestamp 0
transform -1 0 590 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3389_
timestamp 0
transform 1 0 2450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3390_
timestamp 0
transform 1 0 3270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3391_
timestamp 0
transform 1 0 2990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3392_
timestamp 0
transform -1 0 2830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3393_
timestamp 0
transform 1 0 2230 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3394_
timestamp 0
transform 1 0 630 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3395_
timestamp 0
transform -1 0 590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3396_
timestamp 0
transform -1 0 330 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3397_
timestamp 0
transform -1 0 350 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3398_
timestamp 0
transform -1 0 50 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3399_
timestamp 0
transform 1 0 30 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3400_
timestamp 0
transform -1 0 830 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3401_
timestamp 0
transform -1 0 1410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3402_
timestamp 0
transform 1 0 1390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3403_
timestamp 0
transform 1 0 1110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3404_
timestamp 0
transform -1 0 50 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3405_
timestamp 0
transform -1 0 310 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3406_
timestamp 0
transform -1 0 50 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3407_
timestamp 0
transform -1 0 330 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3408_
timestamp 0
transform -1 0 50 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3409_
timestamp 0
transform -1 0 50 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3410_
timestamp 0
transform 1 0 1370 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3411_
timestamp 0
transform 1 0 1090 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3412_
timestamp 0
transform -1 0 570 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3413_
timestamp 0
transform 1 0 310 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3414_
timestamp 0
transform 1 0 570 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1__3415_
timestamp 0
transform -1 0 890 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3416_
timestamp 0
transform 1 0 570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3417_
timestamp 0
transform -1 0 610 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3418_
timestamp 0
transform -1 0 310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3419_
timestamp 0
transform -1 0 1130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3420_
timestamp 0
transform 1 0 830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3421_
timestamp 0
transform 1 0 1130 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3422_
timestamp 0
transform 1 0 850 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3423_
timestamp 0
transform 1 0 1150 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3424_
timestamp 0
transform -1 0 1170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3425_
timestamp 0
transform -1 0 890 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3426_
timestamp 0
transform 1 0 870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1__3427_
timestamp 0
transform -1 0 1390 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3428_
timestamp 0
transform 1 0 1070 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3429_
timestamp 0
transform -1 0 850 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3430_
timestamp 0
transform 1 0 1370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3431_
timestamp 0
transform 1 0 1090 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3432_
timestamp 0
transform -1 0 890 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3433_
timestamp 0
transform -1 0 50 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3434_
timestamp 0
transform -1 0 630 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3435_
timestamp 0
transform -1 0 910 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3436_
timestamp 0
transform -1 0 850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3437_
timestamp 0
transform 1 0 1670 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3438_
timestamp 0
transform 1 0 1130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3439_
timestamp 0
transform -1 0 1410 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3440_
timestamp 0
transform 1 0 1130 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3441_
timestamp 0
transform -1 0 570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3442_
timestamp 0
transform 1 0 1150 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3443_
timestamp 0
transform 1 0 1070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3444_
timestamp 0
transform -1 0 1970 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3445_
timestamp 0
transform 1 0 1650 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3446_
timestamp 0
transform 1 0 2010 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3447_
timestamp 0
transform 1 0 1910 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3448_
timestamp 0
transform -1 0 1710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3449_
timestamp 0
transform 1 0 1390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3450_
timestamp 0
transform -1 0 850 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3451_
timestamp 0
transform 1 0 1110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3452_
timestamp 0
transform 1 0 810 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3453_
timestamp 0
transform -1 0 2130 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3454_
timestamp 0
transform 1 0 3050 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3455_
timestamp 0
transform -1 0 1990 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3456_
timestamp 0
transform -1 0 1650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3457_
timestamp 0
transform -1 0 2830 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3458_
timestamp 0
transform -1 0 1690 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3459_
timestamp 0
transform -1 0 1630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3460_
timestamp 0
transform 1 0 1670 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3461_
timestamp 0
transform -1 0 1890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3462_
timestamp 0
transform -1 0 1650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3463_
timestamp 0
transform -1 0 1410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3464_
timestamp 0
transform 1 0 1130 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3465_
timestamp 0
transform -1 0 1390 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3466_
timestamp 0
transform 1 0 1930 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3467_
timestamp 0
transform 1 0 1930 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3468_
timestamp 0
transform 1 0 2690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3469_
timestamp 0
transform 1 0 2550 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3470_
timestamp 0
transform -1 0 2450 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3471_
timestamp 0
transform 1 0 2270 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3472_
timestamp 0
transform -1 0 2170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3473_
timestamp 0
transform 1 0 1410 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3474_
timestamp 0
transform -1 0 1670 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3475_
timestamp 0
transform 1 0 1150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3476_
timestamp 0
transform -1 0 890 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3477_
timestamp 0
transform 1 0 310 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3478_
timestamp 0
transform -1 0 290 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3479_
timestamp 0
transform -1 0 50 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3480_
timestamp 0
transform -1 0 50 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3481_
timestamp 0
transform -1 0 50 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3482_
timestamp 0
transform 1 0 570 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3483_
timestamp 0
transform -1 0 290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3484_
timestamp 0
transform 1 0 1910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3485_
timestamp 0
transform -1 0 1970 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3486_
timestamp 0
transform -1 0 1350 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3487_
timestamp 0
transform -1 0 1670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3488_
timestamp 0
transform -1 0 1470 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3489_
timestamp 0
transform 1 0 1410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3490_
timestamp 0
transform 1 0 1090 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3491_
timestamp 0
transform -1 0 1170 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3492_
timestamp 0
transform 1 0 1070 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3493_
timestamp 0
transform -1 0 890 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3494_
timestamp 0
transform 1 0 810 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3495_
timestamp 0
transform -1 0 570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3496_
timestamp 0
transform 1 0 330 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3497_
timestamp 0
transform -1 0 290 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3498_
timestamp 0
transform 1 0 590 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3499_
timestamp 0
transform -1 0 650 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3500_
timestamp 0
transform 1 0 590 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3501_
timestamp 0
transform 1 0 830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3502_
timestamp 0
transform -1 0 350 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3503_
timestamp 0
transform -1 0 330 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3504_
timestamp 0
transform -1 0 570 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3505_
timestamp 0
transform -1 0 330 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3506_
timestamp 0
transform -1 0 50 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3507_
timestamp 0
transform -1 0 50 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3508_
timestamp 0
transform 1 0 570 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3509_
timestamp 0
transform -1 0 830 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3510_
timestamp 0
transform -1 0 330 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3511_
timestamp 0
transform -1 0 50 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3512_
timestamp 0
transform 1 0 530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3513_
timestamp 0
transform -1 0 350 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3514_
timestamp 0
transform -1 0 290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3515_
timestamp 0
transform -1 0 50 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3516_
timestamp 0
transform -1 0 50 0 1 10150
box -6 -8 26 268
use FILL  FILL_1__3517_
timestamp 0
transform 1 0 590 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3518_
timestamp 0
transform 1 0 810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3519_
timestamp 0
transform 1 0 2510 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3520_
timestamp 0
transform 1 0 2790 0 1 9110
box -6 -8 26 268
use FILL  FILL_1__3521_
timestamp 0
transform 1 0 3270 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3522_
timestamp 0
transform 1 0 2970 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3523_
timestamp 0
transform 1 0 2530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3524_
timestamp 0
transform -1 0 910 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3525_
timestamp 0
transform -1 0 50 0 1 10670
box -6 -8 26 268
use FILL  FILL_1__3526_
timestamp 0
transform -1 0 50 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3527_
timestamp 0
transform -1 0 550 0 1 11190
box -6 -8 26 268
use FILL  FILL_1__3528_
timestamp 0
transform -1 0 570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_1__3529_
timestamp 0
transform -1 0 50 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1__3530_
timestamp 0
transform -1 0 50 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3531_
timestamp 0
transform 1 0 30 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3532_
timestamp 0
transform 1 0 270 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3533_
timestamp 0
transform -1 0 50 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3534_
timestamp 0
transform -1 0 570 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3535_
timestamp 0
transform -1 0 330 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1__3536_
timestamp 0
transform -1 0 310 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3537_
timestamp 0
transform -1 0 1670 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3538_
timestamp 0
transform 1 0 2430 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3539_
timestamp 0
transform -1 0 2530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3540_
timestamp 0
transform -1 0 2270 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3541_
timestamp 0
transform -1 0 1990 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3542_
timestamp 0
transform -1 0 2170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3543_
timestamp 0
transform 1 0 1570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3544_
timestamp 0
transform 1 0 1930 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3545_
timestamp 0
transform 1 0 1730 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3546_
timestamp 0
transform 1 0 1850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1__3547_
timestamp 0
transform -1 0 2510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3548_
timestamp 0
transform 1 0 2210 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1__3549_
timestamp 0
transform -1 0 2310 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3550_
timestamp 0
transform 1 0 2010 0 1 11710
box -6 -8 26 268
use FILL  FILL_1__3551_
timestamp 0
transform -1 0 2490 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3552_
timestamp 0
transform 1 0 2190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1__3553_
timestamp 0
transform -1 0 1730 0 1 8070
box -6 -8 26 268
use FILL  FILL_1__3554_
timestamp 0
transform 1 0 870 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3555_
timestamp 0
transform 1 0 270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3556_
timestamp 0
transform 1 0 1130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1__3557_
timestamp 0
transform -1 0 3030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3558_
timestamp 0
transform 1 0 2730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1__3559_
timestamp 0
transform -1 0 2490 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3560_
timestamp 0
transform 1 0 2190 0 1 9630
box -6 -8 26 268
use FILL  FILL_1__3561_
timestamp 0
transform -1 0 1910 0 1 7550
box -6 -8 26 268
use FILL  FILL_1__3562_
timestamp 0
transform -1 0 2730 0 1 8590
box -6 -8 26 268
use FILL  FILL_1__3563_
timestamp 0
transform 1 0 2130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1__3564_
timestamp 0
transform 1 0 2410 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3565_
timestamp 0
transform -1 0 1410 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3566_
timestamp 0
transform -1 0 1670 0 1 7030
box -6 -8 26 268
use FILL  FILL_1__3579_
timestamp 0
transform -1 0 5010 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3580_
timestamp 0
transform -1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__3581_
timestamp 0
transform -1 0 3430 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3582_
timestamp 0
transform -1 0 3170 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3583_
timestamp 0
transform -1 0 5290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__3584_
timestamp 0
transform 1 0 4470 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3585_
timestamp 0
transform 1 0 2890 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3586_
timestamp 0
transform -1 0 5810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__3587_
timestamp 0
transform 1 0 30 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3588_
timestamp 0
transform -1 0 50 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__3589_
timestamp 0
transform -1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__3590_
timestamp 0
transform -1 0 50 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__3591_
timestamp 0
transform -1 0 330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3592_
timestamp 0
transform -1 0 50 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__3593_
timestamp 0
transform -1 0 4750 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3594_
timestamp 0
transform 1 0 5790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__3595_
timestamp 0
transform 1 0 5530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__3596_
timestamp 0
transform -1 0 830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3597_
timestamp 0
transform -1 0 50 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__3598_
timestamp 0
transform -1 0 310 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__3599_
timestamp 0
transform -1 0 50 0 1 6510
box -6 -8 26 268
use FILL  FILL_1__3600_
timestamp 0
transform -1 0 50 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__3601_
timestamp 0
transform -1 0 50 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__3602_
timestamp 0
transform -1 0 1670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__3603_
timestamp 0
transform 1 0 6830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform 1 0 7850 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 9350 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 8110 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 10970 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform 1 0 570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform -1 0 12050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 9550 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 7010 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 830 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 10090 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform -1 0 870 0 1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform -1 0 5950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform 1 0 11510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform -1 0 6130 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform 1 0 6750 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform -1 0 3290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform -1 0 3910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform 1 0 7150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform -1 0 6970 0 1 11190
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform 1 0 5290 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 8530 0 1 11190
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform -1 0 8450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 1410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform 1 0 3390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform -1 0 4290 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform 1 0 8130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform 1 0 5070 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform -1 0 1210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert39
timestamp 0
transform 1 0 6290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert40
timestamp 0
transform 1 0 7650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert41
timestamp 0
transform -1 0 8790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert42
timestamp 0
transform -1 0 6930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert43
timestamp 0
transform -1 0 8830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert44
timestamp 0
transform -1 0 8950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert45
timestamp 0
transform 1 0 11010 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert46
timestamp 0
transform 1 0 9450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert47
timestamp 0
transform 1 0 9170 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert48
timestamp 0
transform 1 0 6910 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert49
timestamp 0
transform 1 0 7170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert50
timestamp 0
transform -1 0 7550 0 1 9110
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert51
timestamp 0
transform 1 0 7510 0 1 10150
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert52
timestamp 0
transform 1 0 8910 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert53
timestamp 0
transform 1 0 9950 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert54
timestamp 0
transform 1 0 8790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert55
timestamp 0
transform 1 0 8650 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert56
timestamp 0
transform -1 0 2190 0 1 8590
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert57
timestamp 0
transform 1 0 2490 0 1 11190
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert58
timestamp 0
transform 1 0 2630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert59
timestamp 0
transform -1 0 2190 0 1 10670
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert60
timestamp 0
transform -1 0 10450 0 1 7550
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert61
timestamp 0
transform 1 0 10510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert62
timestamp 0
transform 1 0 10470 0 1 8070
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert63
timestamp 0
transform -1 0 9130 0 1 7550
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert64
timestamp 0
transform -1 0 8570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert65
timestamp 0
transform 1 0 5170 0 1 270
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert66
timestamp 0
transform 1 0 5690 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert67
timestamp 0
transform -1 0 2990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert68
timestamp 0
transform 1 0 3110 0 1 270
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert69
timestamp 0
transform -1 0 6610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert70
timestamp 0
transform 1 0 8550 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert71
timestamp 0
transform -1 0 9210 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert72
timestamp 0
transform -1 0 6730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert73
timestamp 0
transform 1 0 8890 0 -1 7030
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert74
timestamp 0
transform 1 0 10750 0 1 7030
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert75
timestamp 0
transform 1 0 2530 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert76
timestamp 0
transform -1 0 3030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert77
timestamp 0
transform 1 0 10410 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert78
timestamp 0
transform 1 0 9270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert79
timestamp 0
transform -1 0 8310 0 1 7550
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert80
timestamp 0
transform 1 0 7110 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert81
timestamp 0
transform 1 0 7570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert82
timestamp 0
transform -1 0 7550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert83
timestamp 0
transform -1 0 7330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert84
timestamp 0
transform 1 0 9390 0 1 8590
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert85
timestamp 0
transform -1 0 8870 0 1 8590
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert86
timestamp 0
transform -1 0 9470 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert87
timestamp 0
transform 1 0 9370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert88
timestamp 0
transform -1 0 10710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert89
timestamp 0
transform 1 0 9350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert90
timestamp 0
transform 1 0 5330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert91
timestamp 0
transform -1 0 4870 0 1 10670
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert92
timestamp 0
transform -1 0 4710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert93
timestamp 0
transform 1 0 5130 0 1 10150
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert94
timestamp 0
transform -1 0 11290 0 1 9630
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert95
timestamp 0
transform -1 0 11330 0 -1 10150
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert96
timestamp 0
transform -1 0 10050 0 1 11710
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert97
timestamp 0
transform 1 0 11410 0 1 11710
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert28
timestamp 0
transform -1 0 5990 0 -1 11710
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert29
timestamp 0
transform -1 0 2170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert30
timestamp 0
transform 1 0 4510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert31
timestamp 0
transform -1 0 3210 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert32
timestamp 0
transform 1 0 7110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert33
timestamp 0
transform 1 0 5690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert34
timestamp 0
transform -1 0 2450 0 1 10670
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert35
timestamp 0
transform -1 0 5210 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert36
timestamp 0
transform -1 0 2330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert37
timestamp 0
transform 1 0 7350 0 -1 12230
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert38
timestamp 0
transform -1 0 4330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__1688_
timestamp 0
transform -1 0 870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1689_
timestamp 0
transform -1 0 330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1690_
timestamp 0
transform -1 0 590 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1691_
timestamp 0
transform 1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1692_
timestamp 0
transform -1 0 310 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1693_
timestamp 0
transform 1 0 550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1694_
timestamp 0
transform -1 0 5550 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1695_
timestamp 0
transform -1 0 330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1696_
timestamp 0
transform -1 0 330 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1697_
timestamp 0
transform -1 0 1450 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__1698_
timestamp 0
transform -1 0 3390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1699_
timestamp 0
transform 1 0 2830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1700_
timestamp 0
transform -1 0 3870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__1701_
timestamp 0
transform -1 0 570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1702_
timestamp 0
transform -1 0 570 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1703_
timestamp 0
transform 1 0 3210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1704_
timestamp 0
transform -1 0 350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1705_
timestamp 0
transform 1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1706_
timestamp 0
transform -1 0 3830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1707_
timestamp 0
transform -1 0 590 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1708_
timestamp 0
transform 1 0 590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1709_
timestamp 0
transform 1 0 4110 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1710_
timestamp 0
transform -1 0 5590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1711_
timestamp 0
transform 1 0 5130 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1712_
timestamp 0
transform 1 0 7270 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1713_
timestamp 0
transform -1 0 9650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1714_
timestamp 0
transform -1 0 9850 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1715_
timestamp 0
transform -1 0 8530 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1716_
timestamp 0
transform 1 0 11290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1717_
timestamp 0
transform 1 0 11090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1718_
timestamp 0
transform 1 0 11910 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1719_
timestamp 0
transform -1 0 8790 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1720_
timestamp 0
transform -1 0 10110 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1721_
timestamp 0
transform -1 0 10130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1722_
timestamp 0
transform -1 0 9890 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1723_
timestamp 0
transform 1 0 9990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1724_
timestamp 0
transform 1 0 9210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1725_
timestamp 0
transform 1 0 9050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1726_
timestamp 0
transform 1 0 10150 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1727_
timestamp 0
transform -1 0 8770 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1728_
timestamp 0
transform 1 0 11550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1729_
timestamp 0
transform 1 0 10150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1730_
timestamp 0
transform 1 0 8330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1731_
timestamp 0
transform 1 0 8570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1732_
timestamp 0
transform -1 0 7770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1733_
timestamp 0
transform 1 0 9710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1734_
timestamp 0
transform 1 0 7410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1735_
timestamp 0
transform 1 0 10850 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1736_
timestamp 0
transform -1 0 10650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1737_
timestamp 0
transform -1 0 10910 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1738_
timestamp 0
transform -1 0 10290 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1739_
timestamp 0
transform -1 0 10290 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1740_
timestamp 0
transform 1 0 10510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1741_
timestamp 0
transform -1 0 8410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1742_
timestamp 0
transform -1 0 8310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1743_
timestamp 0
transform -1 0 9870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1744_
timestamp 0
transform 1 0 9750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1745_
timestamp 0
transform -1 0 9450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1746_
timestamp 0
transform 1 0 11310 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1747_
timestamp 0
transform 1 0 10790 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1748_
timestamp 0
transform 1 0 7510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1749_
timestamp 0
transform 1 0 7930 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1750_
timestamp 0
transform -1 0 8050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1751_
timestamp 0
transform 1 0 7450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1752_
timestamp 0
transform -1 0 8870 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1753_
timestamp 0
transform 1 0 9730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1754_
timestamp 0
transform -1 0 8270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1755_
timestamp 0
transform -1 0 8850 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__1756_
timestamp 0
transform -1 0 11190 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1757_
timestamp 0
transform 1 0 11050 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1758_
timestamp 0
transform -1 0 9110 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1759_
timestamp 0
transform -1 0 7350 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__1760_
timestamp 0
transform 1 0 8850 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__1761_
timestamp 0
transform -1 0 9570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1762_
timestamp 0
transform 1 0 10590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1763_
timestamp 0
transform -1 0 9030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1764_
timestamp 0
transform 1 0 11290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1765_
timestamp 0
transform 1 0 8110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1766_
timestamp 0
transform 1 0 8490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1767_
timestamp 0
transform 1 0 9190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__1768_
timestamp 0
transform 1 0 8050 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__1769_
timestamp 0
transform 1 0 8570 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__1770_
timestamp 0
transform 1 0 9010 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__1771_
timestamp 0
transform 1 0 8970 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__1772_
timestamp 0
transform 1 0 8690 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__1773_
timestamp 0
transform 1 0 10770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1774_
timestamp 0
transform 1 0 10770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1775_
timestamp 0
transform 1 0 10010 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1776_
timestamp 0
transform -1 0 8010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1777_
timestamp 0
transform 1 0 8050 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1778_
timestamp 0
transform -1 0 7530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1779_
timestamp 0
transform 1 0 5670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1780_
timestamp 0
transform -1 0 4070 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1781_
timestamp 0
transform -1 0 10790 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1782_
timestamp 0
transform 1 0 8270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1783_
timestamp 0
transform 1 0 10510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1784_
timestamp 0
transform -1 0 9990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1785_
timestamp 0
transform -1 0 9750 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1786_
timestamp 0
transform 1 0 10170 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1787_
timestamp 0
transform -1 0 9110 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1788_
timestamp 0
transform -1 0 8530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1789_
timestamp 0
transform 1 0 9970 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1790_
timestamp 0
transform -1 0 10030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1791_
timestamp 0
transform -1 0 10110 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1792_
timestamp 0
transform -1 0 9650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1793_
timestamp 0
transform -1 0 9390 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1794_
timestamp 0
transform 1 0 9110 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1795_
timestamp 0
transform -1 0 8310 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1796_
timestamp 0
transform -1 0 8250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1797_
timestamp 0
transform 1 0 7090 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1798_
timestamp 0
transform 1 0 7350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1799_
timestamp 0
transform -1 0 9370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1800_
timestamp 0
transform 1 0 11250 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1801_
timestamp 0
transform 1 0 9270 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1802_
timestamp 0
transform -1 0 8930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1803_
timestamp 0
transform 1 0 10530 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1804_
timestamp 0
transform -1 0 8550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1805_
timestamp 0
transform -1 0 8650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1806_
timestamp 0
transform 1 0 7590 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1807_
timestamp 0
transform -1 0 8050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1808_
timestamp 0
transform -1 0 8370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1809_
timestamp 0
transform 1 0 8590 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1810_
timestamp 0
transform 1 0 7990 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1811_
timestamp 0
transform -1 0 7730 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1812_
timestamp 0
transform -1 0 8370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1813_
timestamp 0
transform -1 0 8090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1814_
timestamp 0
transform -1 0 7830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1815_
timestamp 0
transform 1 0 7850 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1816_
timestamp 0
transform -1 0 3850 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1817_
timestamp 0
transform 1 0 1330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1818_
timestamp 0
transform -1 0 6150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1819_
timestamp 0
transform -1 0 910 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1820_
timestamp 0
transform 1 0 350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1821_
timestamp 0
transform 1 0 870 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1822_
timestamp 0
transform -1 0 330 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1823_
timestamp 0
transform 1 0 1690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1824_
timestamp 0
transform 1 0 1270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1825_
timestamp 0
transform -1 0 1110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1826_
timestamp 0
transform -1 0 370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1827_
timestamp 0
transform 1 0 870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1828_
timestamp 0
transform -1 0 1470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1829_
timestamp 0
transform -1 0 610 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1830_
timestamp 0
transform -1 0 1410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1831_
timestamp 0
transform 1 0 1990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1832_
timestamp 0
transform -1 0 7990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1833_
timestamp 0
transform 1 0 9630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1834_
timestamp 0
transform 1 0 9210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1835_
timestamp 0
transform -1 0 7730 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1836_
timestamp 0
transform -1 0 6390 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1837_
timestamp 0
transform -1 0 7730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1838_
timestamp 0
transform -1 0 7170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1839_
timestamp 0
transform -1 0 6150 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1840_
timestamp 0
transform 1 0 8530 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1841_
timestamp 0
transform -1 0 8150 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1842_
timestamp 0
transform -1 0 6910 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1843_
timestamp 0
transform -1 0 6630 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1844_
timestamp 0
transform 1 0 9050 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1845_
timestamp 0
transform 1 0 9590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1846_
timestamp 0
transform -1 0 9190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1847_
timestamp 0
transform -1 0 8350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1848_
timestamp 0
transform 1 0 11190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1849_
timestamp 0
transform -1 0 11510 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1850_
timestamp 0
transform -1 0 10970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1851_
timestamp 0
transform 1 0 10330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1852_
timestamp 0
transform -1 0 10390 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1853_
timestamp 0
transform -1 0 10410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1854_
timestamp 0
transform -1 0 7390 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1855_
timestamp 0
transform 1 0 7370 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1856_
timestamp 0
transform 1 0 7650 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1857_
timestamp 0
transform -1 0 8790 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__1858_
timestamp 0
transform -1 0 9330 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1859_
timestamp 0
transform -1 0 8790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1860_
timestamp 0
transform 1 0 9050 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1861_
timestamp 0
transform 1 0 6790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1862_
timestamp 0
transform -1 0 8290 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__1863_
timestamp 0
transform 1 0 7650 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1864_
timestamp 0
transform -1 0 6290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1865_
timestamp 0
transform -1 0 7730 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__1866_
timestamp 0
transform -1 0 7190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1867_
timestamp 0
transform -1 0 7970 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1868_
timestamp 0
transform 1 0 7690 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1869_
timestamp 0
transform -1 0 5990 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__1870_
timestamp 0
transform 1 0 9330 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1871_
timestamp 0
transform 1 0 8810 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1872_
timestamp 0
transform -1 0 8550 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1873_
timestamp 0
transform -1 0 7750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1874_
timestamp 0
transform -1 0 7470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1875_
timestamp 0
transform -1 0 8270 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1876_
timestamp 0
transform -1 0 6910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1877_
timestamp 0
transform -1 0 5750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__1878_
timestamp 0
transform 1 0 6630 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1879_
timestamp 0
transform -1 0 7430 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1880_
timestamp 0
transform 1 0 5950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__1881_
timestamp 0
transform 1 0 5950 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__1882_
timestamp 0
transform -1 0 4910 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__1883_
timestamp 0
transform -1 0 7810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1884_
timestamp 0
transform -1 0 8050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1885_
timestamp 0
transform -1 0 8610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1886_
timestamp 0
transform 1 0 8450 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1887_
timestamp 0
transform -1 0 8430 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1888_
timestamp 0
transform 1 0 11570 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1889_
timestamp 0
transform -1 0 8430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1890_
timestamp 0
transform 1 0 9690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1891_
timestamp 0
transform 1 0 8850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1892_
timestamp 0
transform -1 0 8570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1893_
timestamp 0
transform 1 0 12090 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1894_
timestamp 0
transform 1 0 12070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1895_
timestamp 0
transform 1 0 12090 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1896_
timestamp 0
transform -1 0 10710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1897_
timestamp 0
transform -1 0 9110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1898_
timestamp 0
transform 1 0 8990 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1899_
timestamp 0
transform 1 0 7430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1900_
timestamp 0
transform 1 0 9630 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1901_
timestamp 0
transform 1 0 7970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1902_
timestamp 0
transform -1 0 8190 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1903_
timestamp 0
transform 1 0 7910 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1904_
timestamp 0
transform 1 0 11830 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1905_
timestamp 0
transform 1 0 11590 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1906_
timestamp 0
transform -1 0 6470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1907_
timestamp 0
transform -1 0 7010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1908_
timestamp 0
transform -1 0 6930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1909_
timestamp 0
transform -1 0 6690 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1910_
timestamp 0
transform -1 0 6190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1911_
timestamp 0
transform 1 0 6770 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1912_
timestamp 0
transform 1 0 6230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1913_
timestamp 0
transform 1 0 6170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1914_
timestamp 0
transform 1 0 5670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1915_
timestamp 0
transform 1 0 5190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1916_
timestamp 0
transform 1 0 5190 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__1917_
timestamp 0
transform -1 0 3690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__1918_
timestamp 0
transform 1 0 3570 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__1919_
timestamp 0
transform -1 0 3850 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__1920_
timestamp 0
transform -1 0 3570 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__1921_
timestamp 0
transform -1 0 1690 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__1922_
timestamp 0
transform 1 0 7490 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1923_
timestamp 0
transform 1 0 7750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1924_
timestamp 0
transform -1 0 6350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1925_
timestamp 0
transform -1 0 4590 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1926_
timestamp 0
transform -1 0 3950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1927_
timestamp 0
transform 1 0 1990 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__1928_
timestamp 0
transform -1 0 3150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__1929_
timestamp 0
transform 1 0 4530 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__1930_
timestamp 0
transform 1 0 3090 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__1931_
timestamp 0
transform -1 0 2870 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__1932_
timestamp 0
transform -1 0 1470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1933_
timestamp 0
transform -1 0 8430 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1934_
timestamp 0
transform 1 0 3830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1935_
timestamp 0
transform -1 0 3850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1936_
timestamp 0
transform -1 0 2530 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1937_
timestamp 0
transform -1 0 1190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1938_
timestamp 0
transform -1 0 3550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1939_
timestamp 0
transform -1 0 4110 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1940_
timestamp 0
transform -1 0 3330 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1941_
timestamp 0
transform -1 0 3270 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1942_
timestamp 0
transform -1 0 1770 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__1943_
timestamp 0
transform -1 0 3570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1944_
timestamp 0
transform -1 0 3670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1945_
timestamp 0
transform -1 0 2930 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1946_
timestamp 0
transform -1 0 1490 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__1947_
timestamp 0
transform -1 0 4910 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__1948_
timestamp 0
transform 1 0 5110 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__1949_
timestamp 0
transform 1 0 5170 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__1950_
timestamp 0
transform -1 0 4910 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__1951_
timestamp 0
transform -1 0 1950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1952_
timestamp 0
transform 1 0 4070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1953_
timestamp 0
transform 1 0 4010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1954_
timestamp 0
transform 1 0 4150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1955_
timestamp 0
transform -1 0 1670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1956_
timestamp 0
transform -1 0 4290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__1957_
timestamp 0
transform 1 0 4870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__1958_
timestamp 0
transform -1 0 5150 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__1959_
timestamp 0
transform -1 0 4130 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__1960_
timestamp 0
transform -1 0 2290 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1961_
timestamp 0
transform 1 0 4110 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1962_
timestamp 0
transform 1 0 3870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1963_
timestamp 0
transform 1 0 3650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1964_
timestamp 0
transform 1 0 1990 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1965_
timestamp 0
transform 1 0 6370 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__1966_
timestamp 0
transform 1 0 6310 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1967_
timestamp 0
transform 1 0 7150 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1968_
timestamp 0
transform 1 0 6610 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1969_
timestamp 0
transform -1 0 3270 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__1970_
timestamp 0
transform 1 0 2810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1971_
timestamp 0
transform -1 0 4690 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1972_
timestamp 0
transform 1 0 3550 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1973_
timestamp 0
transform -1 0 3570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1974_
timestamp 0
transform -1 0 3070 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__1975_
timestamp 0
transform 1 0 2970 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__1976_
timestamp 0
transform -1 0 3070 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__1977_
timestamp 0
transform 1 0 4350 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__1978_
timestamp 0
transform 1 0 3050 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__1979_
timestamp 0
transform -1 0 2790 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__1980_
timestamp 0
transform -1 0 2310 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1981_
timestamp 0
transform 1 0 5930 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1982_
timestamp 0
transform 1 0 6050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1983_
timestamp 0
transform 1 0 6250 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1984_
timestamp 0
transform 1 0 5250 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1985_
timestamp 0
transform -1 0 4750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1986_
timestamp 0
transform 1 0 2530 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__1987_
timestamp 0
transform -1 0 7250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1988_
timestamp 0
transform 1 0 7550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1989_
timestamp 0
transform 1 0 7610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1990_
timestamp 0
transform -1 0 7410 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1991_
timestamp 0
transform -1 0 7690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1992_
timestamp 0
transform 1 0 10430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1993_
timestamp 0
transform 1 0 9550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__1994_
timestamp 0
transform -1 0 6230 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__1995_
timestamp 0
transform 1 0 6610 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1996_
timestamp 0
transform -1 0 6750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1997_
timestamp 0
transform 1 0 6450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1998_
timestamp 0
transform 1 0 6450 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__1999_
timestamp 0
transform 1 0 7510 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2000_
timestamp 0
transform 1 0 6430 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2001_
timestamp 0
transform 1 0 6670 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2002_
timestamp 0
transform 1 0 6630 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2003_
timestamp 0
transform 1 0 9510 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2004_
timestamp 0
transform 1 0 7450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2005_
timestamp 0
transform -1 0 7250 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2006_
timestamp 0
transform 1 0 6730 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2007_
timestamp 0
transform 1 0 6570 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2008_
timestamp 0
transform -1 0 6210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2009_
timestamp 0
transform 1 0 6810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2010_
timestamp 0
transform -1 0 7030 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2011_
timestamp 0
transform 1 0 7270 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2012_
timestamp 0
transform -1 0 9410 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2013_
timestamp 0
transform 1 0 10550 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2014_
timestamp 0
transform -1 0 10810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2015_
timestamp 0
transform -1 0 6250 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2016_
timestamp 0
transform -1 0 7290 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2017_
timestamp 0
transform -1 0 7070 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2018_
timestamp 0
transform 1 0 7310 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2019_
timestamp 0
transform 1 0 9390 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2020_
timestamp 0
transform -1 0 10290 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2021_
timestamp 0
transform -1 0 7330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2022_
timestamp 0
transform 1 0 7570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2023_
timestamp 0
transform -1 0 7870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2024_
timestamp 0
transform 1 0 6090 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2025_
timestamp 0
transform -1 0 5970 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2026_
timestamp 0
transform 1 0 9670 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2027_
timestamp 0
transform 1 0 10210 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2028_
timestamp 0
transform -1 0 10210 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2029_
timestamp 0
transform -1 0 11090 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2030_
timestamp 0
transform 1 0 10710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2031_
timestamp 0
transform -1 0 11010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2032_
timestamp 0
transform 1 0 8930 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2033_
timestamp 0
transform 1 0 8390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2034_
timestamp 0
transform 1 0 8630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2035_
timestamp 0
transform 1 0 8590 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2036_
timestamp 0
transform 1 0 11550 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2037_
timestamp 0
transform 1 0 11750 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2038_
timestamp 0
transform -1 0 7590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2039_
timestamp 0
transform -1 0 6670 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2040_
timestamp 0
transform 1 0 10930 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2041_
timestamp 0
transform 1 0 11010 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2042_
timestamp 0
transform -1 0 10090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2043_
timestamp 0
transform -1 0 10470 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2044_
timestamp 0
transform -1 0 10990 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2045_
timestamp 0
transform -1 0 11330 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2046_
timestamp 0
transform 1 0 8810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2047_
timestamp 0
transform -1 0 9370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2048_
timestamp 0
transform 1 0 9170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2049_
timestamp 0
transform 1 0 9310 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2050_
timestamp 0
transform 1 0 9070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2051_
timestamp 0
transform 1 0 8770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2052_
timestamp 0
transform 1 0 9050 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2053_
timestamp 0
transform -1 0 9610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2054_
timestamp 0
transform 1 0 9830 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2055_
timestamp 0
transform -1 0 6470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2056_
timestamp 0
transform -1 0 6050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2057_
timestamp 0
transform 1 0 10250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2058_
timestamp 0
transform -1 0 9990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2059_
timestamp 0
transform -1 0 10130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2060_
timestamp 0
transform -1 0 9890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2061_
timestamp 0
transform 1 0 10070 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2062_
timestamp 0
transform -1 0 9150 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2063_
timestamp 0
transform 1 0 8230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2064_
timestamp 0
transform -1 0 7910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2065_
timestamp 0
transform -1 0 8730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2066_
timestamp 0
transform 1 0 8710 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2067_
timestamp 0
transform -1 0 7970 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2068_
timestamp 0
transform -1 0 8250 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2069_
timestamp 0
transform 1 0 7970 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2070_
timestamp 0
transform -1 0 8270 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2071_
timestamp 0
transform -1 0 8550 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2072_
timestamp 0
transform 1 0 8770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2073_
timestamp 0
transform 1 0 9030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2074_
timestamp 0
transform 1 0 9250 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2075_
timestamp 0
transform -1 0 9550 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2076_
timestamp 0
transform 1 0 11210 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2077_
timestamp 0
transform -1 0 11270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2078_
timestamp 0
transform -1 0 11070 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2079_
timestamp 0
transform 1 0 11210 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2080_
timestamp 0
transform -1 0 11050 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2081_
timestamp 0
transform 1 0 11050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2082_
timestamp 0
transform 1 0 10310 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2083_
timestamp 0
transform 1 0 9570 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2084_
timestamp 0
transform 1 0 11590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2085_
timestamp 0
transform 1 0 11010 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2086_
timestamp 0
transform 1 0 11510 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2087_
timestamp 0
transform 1 0 11530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2088_
timestamp 0
transform -1 0 12090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2089_
timestamp 0
transform 1 0 11810 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2090_
timestamp 0
transform 1 0 11990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2091_
timestamp 0
transform 1 0 9890 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2092_
timestamp 0
transform 1 0 10510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2093_
timestamp 0
transform -1 0 11070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2094_
timestamp 0
transform 1 0 11310 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2095_
timestamp 0
transform -1 0 10970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2096_
timestamp 0
transform 1 0 11490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2097_
timestamp 0
transform -1 0 11830 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2098_
timestamp 0
transform -1 0 12010 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2099_
timestamp 0
transform -1 0 11310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2100_
timestamp 0
transform 1 0 11270 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2101_
timestamp 0
transform -1 0 11230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2102_
timestamp 0
transform -1 0 11610 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2103_
timestamp 0
transform 1 0 12090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2104_
timestamp 0
transform 1 0 12090 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2105_
timestamp 0
transform -1 0 11550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2106_
timestamp 0
transform -1 0 11530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2107_
timestamp 0
transform -1 0 12090 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2108_
timestamp 0
transform 1 0 8830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2109_
timestamp 0
transform 1 0 12090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2110_
timestamp 0
transform -1 0 12110 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2111_
timestamp 0
transform -1 0 12110 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2112_
timestamp 0
transform -1 0 12010 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2113_
timestamp 0
transform 1 0 11770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2114_
timestamp 0
transform 1 0 10550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2115_
timestamp 0
transform -1 0 9290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2116_
timestamp 0
transform -1 0 10170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2117_
timestamp 0
transform -1 0 10770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2118_
timestamp 0
transform -1 0 10730 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2119_
timestamp 0
transform 1 0 10630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2120_
timestamp 0
transform 1 0 10670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2121_
timestamp 0
transform -1 0 10410 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2122_
timestamp 0
transform 1 0 10610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2123_
timestamp 0
transform -1 0 8110 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2124_
timestamp 0
transform -1 0 7810 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2125_
timestamp 0
transform -1 0 10170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2126_
timestamp 0
transform 1 0 10570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2127_
timestamp 0
transform -1 0 6990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2128_
timestamp 0
transform -1 0 9130 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2129_
timestamp 0
transform 1 0 7250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2130_
timestamp 0
transform -1 0 10870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2131_
timestamp 0
transform -1 0 7910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2132_
timestamp 0
transform 1 0 6690 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2133_
timestamp 0
transform -1 0 6990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2134_
timestamp 0
transform -1 0 7250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2135_
timestamp 0
transform -1 0 11130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2136_
timestamp 0
transform -1 0 11290 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2137_
timestamp 0
transform 1 0 11270 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2138_
timestamp 0
transform 1 0 11350 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2139_
timestamp 0
transform -1 0 11270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2140_
timestamp 0
transform -1 0 10990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2141_
timestamp 0
transform 1 0 9910 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2142_
timestamp 0
transform 1 0 10710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2143_
timestamp 0
transform -1 0 10450 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2144_
timestamp 0
transform -1 0 11010 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2145_
timestamp 0
transform -1 0 5010 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2146_
timestamp 0
transform 1 0 9730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2147_
timestamp 0
transform 1 0 10290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2148_
timestamp 0
transform -1 0 6230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2149_
timestamp 0
transform 1 0 10010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2150_
timestamp 0
transform 1 0 8790 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2151_
timestamp 0
transform 1 0 7410 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2152_
timestamp 0
transform 1 0 8490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2153_
timestamp 0
transform 1 0 8750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2154_
timestamp 0
transform 1 0 9030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2155_
timestamp 0
transform -1 0 10110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2156_
timestamp 0
transform -1 0 10890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2157_
timestamp 0
transform 1 0 11130 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2158_
timestamp 0
transform -1 0 11710 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2159_
timestamp 0
transform -1 0 11830 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2160_
timestamp 0
transform -1 0 11370 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2161_
timestamp 0
transform 1 0 8110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2162_
timestamp 0
transform 1 0 8870 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2163_
timestamp 0
transform -1 0 9970 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2164_
timestamp 0
transform 1 0 9730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2165_
timestamp 0
transform 1 0 10970 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2166_
timestamp 0
transform 1 0 10790 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2167_
timestamp 0
transform 1 0 9170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2168_
timestamp 0
transform 1 0 9990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2169_
timestamp 0
transform -1 0 8730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2170_
timestamp 0
transform -1 0 9150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2171_
timestamp 0
transform 1 0 10290 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2172_
timestamp 0
transform 1 0 9710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2173_
timestamp 0
transform 1 0 9830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2174_
timestamp 0
transform -1 0 9470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2175_
timestamp 0
transform 1 0 9550 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2176_
timestamp 0
transform -1 0 9670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2177_
timestamp 0
transform -1 0 9370 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2178_
timestamp 0
transform -1 0 10970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2179_
timestamp 0
transform 1 0 9450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2180_
timestamp 0
transform 1 0 11810 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2181_
timestamp 0
transform 1 0 11790 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2182_
timestamp 0
transform 1 0 11870 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2183_
timestamp 0
transform -1 0 11250 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2184_
timestamp 0
transform 1 0 10990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2185_
timestamp 0
transform -1 0 10230 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2186_
timestamp 0
transform 1 0 10170 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2187_
timestamp 0
transform -1 0 10570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2188_
timestamp 0
transform 1 0 11530 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2189_
timestamp 0
transform 1 0 9910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2190_
timestamp 0
transform 1 0 10470 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2191_
timestamp 0
transform 1 0 11090 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2192_
timestamp 0
transform 1 0 11030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2193_
timestamp 0
transform -1 0 10970 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2194_
timestamp 0
transform -1 0 10530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2195_
timestamp 0
transform -1 0 9410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2196_
timestamp 0
transform -1 0 11050 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2197_
timestamp 0
transform 1 0 11310 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2198_
timestamp 0
transform -1 0 9850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2199_
timestamp 0
transform -1 0 9910 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2200_
timestamp 0
transform -1 0 5770 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2201_
timestamp 0
transform 1 0 6290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2202_
timestamp 0
transform 1 0 6030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2203_
timestamp 0
transform 1 0 6030 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2204_
timestamp 0
transform 1 0 6770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2205_
timestamp 0
transform 1 0 7070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2206_
timestamp 0
transform 1 0 9410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2207_
timestamp 0
transform -1 0 9910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2208_
timestamp 0
transform -1 0 9330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2209_
timestamp 0
transform 1 0 10370 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2210_
timestamp 0
transform 1 0 10370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2211_
timestamp 0
transform 1 0 11210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2212_
timestamp 0
transform -1 0 11570 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2213_
timestamp 0
transform -1 0 11610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2214_
timestamp 0
transform 1 0 11570 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2215_
timestamp 0
transform 1 0 11670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2216_
timestamp 0
transform 1 0 12050 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2217_
timestamp 0
transform 1 0 11330 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2218_
timestamp 0
transform 1 0 9610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2219_
timestamp 0
transform -1 0 9850 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2220_
timestamp 0
transform -1 0 9890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2221_
timestamp 0
transform -1 0 11830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2222_
timestamp 0
transform 1 0 11770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2223_
timestamp 0
transform -1 0 11810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2224_
timestamp 0
transform 1 0 11790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2225_
timestamp 0
transform 1 0 10890 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2226_
timestamp 0
transform 1 0 11850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2227_
timestamp 0
transform 1 0 11570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2228_
timestamp 0
transform -1 0 11430 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2229_
timestamp 0
transform -1 0 10510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2230_
timestamp 0
transform -1 0 10230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2231_
timestamp 0
transform -1 0 8430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2232_
timestamp 0
transform 1 0 8670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2233_
timestamp 0
transform 1 0 9450 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2234_
timestamp 0
transform -1 0 9710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2235_
timestamp 0
transform -1 0 9830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2236_
timestamp 0
transform 1 0 7130 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2237_
timestamp 0
transform -1 0 6610 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2238_
timestamp 0
transform -1 0 6890 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2239_
timestamp 0
transform -1 0 8910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2240_
timestamp 0
transform -1 0 8630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2241_
timestamp 0
transform -1 0 8270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2242_
timestamp 0
transform -1 0 7450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2243_
timestamp 0
transform 1 0 7710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2244_
timestamp 0
transform 1 0 7990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2245_
timestamp 0
transform -1 0 7690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2246_
timestamp 0
transform 1 0 9070 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2247_
timestamp 0
transform -1 0 12070 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2248_
timestamp 0
transform 1 0 11270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2249_
timestamp 0
transform -1 0 9430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2250_
timestamp 0
transform 1 0 10950 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2251_
timestamp 0
transform 1 0 10510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2252_
timestamp 0
transform 1 0 11250 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2253_
timestamp 0
transform -1 0 11850 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2254_
timestamp 0
transform 1 0 12090 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2255_
timestamp 0
transform -1 0 10450 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2256_
timestamp 0
transform -1 0 10730 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2257_
timestamp 0
transform 1 0 10970 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2258_
timestamp 0
transform 1 0 12130 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2259_
timestamp 0
transform -1 0 11810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2260_
timestamp 0
transform 1 0 9990 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2261_
timestamp 0
transform 1 0 10250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2262_
timestamp 0
transform -1 0 10770 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2263_
timestamp 0
transform 1 0 11250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2264_
timestamp 0
transform 1 0 12070 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2265_
timestamp 0
transform -1 0 11330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2266_
timestamp 0
transform -1 0 10690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2267_
timestamp 0
transform 1 0 11910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2268_
timestamp 0
transform 1 0 12070 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2269_
timestamp 0
transform -1 0 11850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2270_
timestamp 0
transform 1 0 11270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2271_
timestamp 0
transform -1 0 11570 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2272_
timestamp 0
transform 1 0 11830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2273_
timestamp 0
transform -1 0 12090 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2274_
timestamp 0
transform 1 0 10010 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2275_
timestamp 0
transform -1 0 8170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2276_
timestamp 0
transform 1 0 8830 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2277_
timestamp 0
transform 1 0 9110 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2278_
timestamp 0
transform -1 0 9190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2279_
timestamp 0
transform 1 0 8990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2280_
timestamp 0
transform 1 0 10150 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2281_
timestamp 0
transform 1 0 12030 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2282_
timestamp 0
transform 1 0 12090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2283_
timestamp 0
transform -1 0 10970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2284_
timestamp 0
transform 1 0 12050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2285_
timestamp 0
transform 1 0 12050 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2286_
timestamp 0
transform -1 0 11830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2287_
timestamp 0
transform 1 0 11770 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2288_
timestamp 0
transform -1 0 10930 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2289_
timestamp 0
transform -1 0 10710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2290_
timestamp 0
transform -1 0 10890 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2291_
timestamp 0
transform 1 0 11250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2292_
timestamp 0
transform 1 0 10390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2293_
timestamp 0
transform 1 0 10670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2294_
timestamp 0
transform 1 0 10990 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2295_
timestamp 0
transform 1 0 10870 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2296_
timestamp 0
transform 1 0 11130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2297_
timestamp 0
transform 1 0 11790 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2298_
timestamp 0
transform -1 0 11890 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2299_
timestamp 0
transform -1 0 10450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2300_
timestamp 0
transform 1 0 10150 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2301_
timestamp 0
transform 1 0 11770 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2302_
timestamp 0
transform 1 0 11710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2303_
timestamp 0
transform -1 0 11690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2304_
timestamp 0
transform 1 0 11830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2305_
timestamp 0
transform 1 0 10710 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2306_
timestamp 0
transform -1 0 11570 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2307_
timestamp 0
transform 1 0 11270 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2308_
timestamp 0
transform 1 0 12050 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2309_
timestamp 0
transform -1 0 11610 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2310_
timestamp 0
transform -1 0 11550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2311_
timestamp 0
transform 1 0 11530 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2312_
timestamp 0
transform 1 0 11590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2313_
timestamp 0
transform 1 0 11870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2314_
timestamp 0
transform -1 0 11190 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2315_
timestamp 0
transform 1 0 12050 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2316_
timestamp 0
transform 1 0 11450 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2317_
timestamp 0
transform -1 0 11950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2318_
timestamp 0
transform 1 0 11490 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2319_
timestamp 0
transform 1 0 11130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2320_
timestamp 0
transform 1 0 11550 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2321_
timestamp 0
transform 1 0 11410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2322_
timestamp 0
transform -1 0 11270 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2323_
timestamp 0
transform -1 0 11510 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2324_
timestamp 0
transform 1 0 11750 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2325_
timestamp 0
transform -1 0 12130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2326_
timestamp 0
transform 1 0 12050 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2327_
timestamp 0
transform 1 0 11410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2328_
timestamp 0
transform 1 0 10990 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2329_
timestamp 0
transform 1 0 8510 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2330_
timestamp 0
transform -1 0 10190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2331_
timestamp 0
transform -1 0 9630 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2332_
timestamp 0
transform -1 0 11850 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2333_
timestamp 0
transform -1 0 10730 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2334_
timestamp 0
transform 1 0 10450 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2335_
timestamp 0
transform 1 0 10430 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2336_
timestamp 0
transform 1 0 10610 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2337_
timestamp 0
transform -1 0 10730 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2338_
timestamp 0
transform -1 0 10650 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2339_
timestamp 0
transform -1 0 9570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2340_
timestamp 0
transform -1 0 9850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2341_
timestamp 0
transform 1 0 9550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2342_
timestamp 0
transform -1 0 10430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2343_
timestamp 0
transform -1 0 10370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2344_
timestamp 0
transform -1 0 10610 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2345_
timestamp 0
transform 1 0 11730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2346_
timestamp 0
transform 1 0 11470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2347_
timestamp 0
transform -1 0 8810 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2348_
timestamp 0
transform -1 0 9910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2349_
timestamp 0
transform -1 0 11570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2350_
timestamp 0
transform -1 0 11290 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2351_
timestamp 0
transform -1 0 10350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2352_
timestamp 0
transform -1 0 10110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2353_
timestamp 0
transform -1 0 9410 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2354_
timestamp 0
transform 1 0 7810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2355_
timestamp 0
transform -1 0 6890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2356_
timestamp 0
transform -1 0 6830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2357_
timestamp 0
transform -1 0 7490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2358_
timestamp 0
transform -1 0 7070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2359_
timestamp 0
transform 1 0 7290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2360_
timestamp 0
transform -1 0 7970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2361_
timestamp 0
transform -1 0 7030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2362_
timestamp 0
transform 1 0 8750 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2363_
timestamp 0
transform -1 0 7430 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2364_
timestamp 0
transform 1 0 7170 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2365_
timestamp 0
transform 1 0 6890 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2366_
timestamp 0
transform 1 0 6370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2367_
timestamp 0
transform -1 0 7210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2368_
timestamp 0
transform 1 0 6610 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2369_
timestamp 0
transform 1 0 6990 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2370_
timestamp 0
transform -1 0 7250 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2371_
timestamp 0
transform 1 0 7190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2372_
timestamp 0
transform -1 0 6770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2373_
timestamp 0
transform 1 0 6710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2374_
timestamp 0
transform 1 0 8210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2375_
timestamp 0
transform 1 0 8270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2376_
timestamp 0
transform -1 0 6710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2377_
timestamp 0
transform 1 0 5410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2378_
timestamp 0
transform -1 0 3730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2379_
timestamp 0
transform -1 0 7990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2380_
timestamp 0
transform -1 0 5630 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2381_
timestamp 0
transform -1 0 5910 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2382_
timestamp 0
transform -1 0 5770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2383_
timestamp 0
transform 1 0 4690 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2384_
timestamp 0
transform 1 0 4610 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2385_
timestamp 0
transform 1 0 4850 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2386_
timestamp 0
transform 1 0 5130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2387_
timestamp 0
transform 1 0 1650 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2388_
timestamp 0
transform 1 0 1590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2389_
timestamp 0
transform 1 0 5170 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2390_
timestamp 0
transform 1 0 2450 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2391_
timestamp 0
transform -1 0 2250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2392_
timestamp 0
transform -1 0 1970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2393_
timestamp 0
transform -1 0 2530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2394_
timestamp 0
transform -1 0 2950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2395_
timestamp 0
transform 1 0 4350 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2396_
timestamp 0
transform 1 0 2990 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2397_
timestamp 0
transform -1 0 3070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2398_
timestamp 0
transform -1 0 2790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2399_
timestamp 0
transform 1 0 1890 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2400_
timestamp 0
transform -1 0 1330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2401_
timestamp 0
transform -1 0 2810 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2402_
timestamp 0
transform 1 0 2550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2403_
timestamp 0
transform -1 0 2190 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2404_
timestamp 0
transform -1 0 1630 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2405_
timestamp 0
transform -1 0 1490 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2406_
timestamp 0
transform 1 0 5870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2407_
timestamp 0
transform -1 0 4230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2408_
timestamp 0
transform -1 0 5590 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2409_
timestamp 0
transform -1 0 6410 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2410_
timestamp 0
transform -1 0 4190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2411_
timestamp 0
transform -1 0 3950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2412_
timestamp 0
transform -1 0 1210 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2413_
timestamp 0
transform -1 0 4490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2414_
timestamp 0
transform 1 0 3010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2415_
timestamp 0
transform -1 0 2750 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2416_
timestamp 0
transform 1 0 1710 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2417_
timestamp 0
transform -1 0 2210 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2418_
timestamp 0
transform -1 0 2090 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2419_
timestamp 0
transform -1 0 3410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2420_
timestamp 0
transform 1 0 2830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2421_
timestamp 0
transform -1 0 2750 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2422_
timestamp 0
transform -1 0 1930 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2423_
timestamp 0
transform -1 0 3630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2424_
timestamp 0
transform -1 0 3470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2425_
timestamp 0
transform -1 0 3350 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2426_
timestamp 0
transform 1 0 3110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2427_
timestamp 0
transform 1 0 3270 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2428_
timestamp 0
transform -1 0 3350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2429_
timestamp 0
transform -1 0 5070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2430_
timestamp 0
transform -1 0 7770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2431_
timestamp 0
transform -1 0 5330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2432_
timestamp 0
transform -1 0 9450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2433_
timestamp 0
transform 1 0 11550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2434_
timestamp 0
transform 1 0 10730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2435_
timestamp 0
transform -1 0 7210 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2436_
timestamp 0
transform -1 0 6890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2437_
timestamp 0
transform -1 0 9570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2438_
timestamp 0
transform -1 0 9310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2439_
timestamp 0
transform -1 0 6090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2440_
timestamp 0
transform 1 0 7710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2441_
timestamp 0
transform -1 0 7550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2442_
timestamp 0
transform 1 0 10250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2443_
timestamp 0
transform -1 0 7150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2444_
timestamp 0
transform -1 0 7150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2445_
timestamp 0
transform 1 0 5250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2446_
timestamp 0
transform 1 0 6370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2447_
timestamp 0
transform -1 0 4750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2448_
timestamp 0
transform -1 0 6350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2449_
timestamp 0
transform -1 0 6970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2450_
timestamp 0
transform 1 0 4110 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2451_
timestamp 0
transform -1 0 3990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2452_
timestamp 0
transform 1 0 4630 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2453_
timestamp 0
transform 1 0 8490 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2454_
timestamp 0
transform 1 0 4370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2455_
timestamp 0
transform 1 0 4370 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2456_
timestamp 0
transform -1 0 4230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2457_
timestamp 0
transform -1 0 4490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2458_
timestamp 0
transform -1 0 4850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2459_
timestamp 0
transform 1 0 4990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2460_
timestamp 0
transform 1 0 4870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2461_
timestamp 0
transform 1 0 5150 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2462_
timestamp 0
transform 1 0 5290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2463_
timestamp 0
transform 1 0 6230 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2464_
timestamp 0
transform -1 0 3170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2465_
timestamp 0
transform -1 0 2890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2466_
timestamp 0
transform -1 0 2890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2467_
timestamp 0
transform 1 0 2030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2468_
timestamp 0
transform -1 0 1590 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2469_
timestamp 0
transform 1 0 550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2470_
timestamp 0
transform -1 0 2650 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2471_
timestamp 0
transform -1 0 2670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2472_
timestamp 0
transform -1 0 2370 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2473_
timestamp 0
transform 1 0 1870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2474_
timestamp 0
transform -1 0 1390 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2475_
timestamp 0
transform -1 0 330 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2476_
timestamp 0
transform -1 0 3750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2477_
timestamp 0
transform -1 0 4990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2478_
timestamp 0
transform 1 0 3850 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2479_
timestamp 0
transform -1 0 3490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2480_
timestamp 0
transform 1 0 1730 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2481_
timestamp 0
transform -1 0 3290 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2482_
timestamp 0
transform 1 0 3570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2483_
timestamp 0
transform 1 0 2990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2484_
timestamp 0
transform 1 0 2710 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2485_
timestamp 0
transform -1 0 330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2486_
timestamp 0
transform -1 0 2610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2487_
timestamp 0
transform 1 0 2330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2488_
timestamp 0
transform -1 0 2330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2489_
timestamp 0
transform -1 0 1770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2490_
timestamp 0
transform -1 0 1330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2491_
timestamp 0
transform -1 0 330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2492_
timestamp 0
transform 1 0 4550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2493_
timestamp 0
transform 1 0 3550 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2494_
timestamp 0
transform 1 0 6130 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2495_
timestamp 0
transform 1 0 3790 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2496_
timestamp 0
transform 1 0 4090 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2497_
timestamp 0
transform -1 0 4010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2498_
timestamp 0
transform 1 0 3470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2499_
timestamp 0
transform 1 0 3730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2500_
timestamp 0
transform -1 0 330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2501_
timestamp 0
transform -1 0 3330 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2502_
timestamp 0
transform -1 0 2970 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2503_
timestamp 0
transform -1 0 3450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__2504_
timestamp 0
transform -1 0 3210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__2505_
timestamp 0
transform 1 0 2650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2506_
timestamp 0
transform -1 0 2470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__2507_
timestamp 0
transform 1 0 590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2508_
timestamp 0
transform 1 0 3090 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2509_
timestamp 0
transform 1 0 2630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2510_
timestamp 0
transform -1 0 3190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2511_
timestamp 0
transform 1 0 3270 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__2512_
timestamp 0
transform 1 0 3110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2513_
timestamp 0
transform -1 0 2370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2514_
timestamp 0
transform 1 0 2070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2515_
timestamp 0
transform -1 0 2090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2516_
timestamp 0
transform -1 0 330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__2517_
timestamp 0
transform -1 0 2170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2518_
timestamp 0
transform 1 0 5270 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2519_
timestamp 0
transform -1 0 5810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2520_
timestamp 0
transform -1 0 5910 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2521_
timestamp 0
transform 1 0 5610 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2522_
timestamp 0
transform -1 0 5610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2523_
timestamp 0
transform -1 0 5530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2524_
timestamp 0
transform -1 0 5470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2525_
timestamp 0
transform -1 0 2690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2526_
timestamp 0
transform 1 0 6090 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2527_
timestamp 0
transform 1 0 6490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2528_
timestamp 0
transform 1 0 6470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2529_
timestamp 0
transform 1 0 6070 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2530_
timestamp 0
transform 1 0 5530 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2531_
timestamp 0
transform 1 0 2890 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2532_
timestamp 0
transform 1 0 4170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2533_
timestamp 0
transform 1 0 5110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2534_
timestamp 0
transform 1 0 4830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2535_
timestamp 0
transform -1 0 4570 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2536_
timestamp 0
transform 1 0 3410 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2537_
timestamp 0
transform 1 0 2050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2538_
timestamp 0
transform 1 0 4450 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2539_
timestamp 0
transform 1 0 3830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2540_
timestamp 0
transform 1 0 4170 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2541_
timestamp 0
transform -1 0 4150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2542_
timestamp 0
transform -1 0 3670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2543_
timestamp 0
transform 1 0 3430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2544_
timestamp 0
transform 1 0 4150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2545_
timestamp 0
transform 1 0 4410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2546_
timestamp 0
transform 1 0 4770 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2547_
timestamp 0
transform -1 0 4710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2548_
timestamp 0
transform -1 0 4430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2549_
timestamp 0
transform 1 0 4650 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2550_
timestamp 0
transform 1 0 4650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2551_
timestamp 0
transform 1 0 5170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2552_
timestamp 0
transform 1 0 5410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2553_
timestamp 0
transform 1 0 2310 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2554_
timestamp 0
transform 1 0 4450 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2555_
timestamp 0
transform -1 0 4630 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2556_
timestamp 0
transform -1 0 4870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2557_
timestamp 0
transform 1 0 4570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2558_
timestamp 0
transform 1 0 4650 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2559_
timestamp 0
transform 1 0 4370 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2560_
timestamp 0
transform 1 0 3870 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2561_
timestamp 0
transform 1 0 3570 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2562_
timestamp 0
transform 1 0 2190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2563_
timestamp 0
transform -1 0 4410 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2564_
timestamp 0
transform 1 0 4330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2565_
timestamp 0
transform -1 0 3810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2566_
timestamp 0
transform 1 0 2410 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2567_
timestamp 0
transform 1 0 3890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2568_
timestamp 0
transform -1 0 5690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2569_
timestamp 0
transform -1 0 5830 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2570_
timestamp 0
transform 1 0 5910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2571_
timestamp 0
transform 1 0 5910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2572_
timestamp 0
transform 1 0 5770 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2573_
timestamp 0
transform 1 0 5690 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2574_
timestamp 0
transform 1 0 5670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2575_
timestamp 0
transform -1 0 4710 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2576_
timestamp 0
transform -1 0 4190 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2577_
timestamp 0
transform -1 0 4450 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2578_
timestamp 0
transform 1 0 6950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2579_
timestamp 0
transform 1 0 6970 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2580_
timestamp 0
transform 1 0 7970 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2581_
timestamp 0
transform -1 0 8830 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2582_
timestamp 0
transform 1 0 6870 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2583_
timestamp 0
transform -1 0 6870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2584_
timestamp 0
transform 1 0 7290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2585_
timestamp 0
transform 1 0 7330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2586_
timestamp 0
transform -1 0 8410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2587_
timestamp 0
transform -1 0 6750 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2588_
timestamp 0
transform -1 0 5790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2589_
timestamp 0
transform 1 0 7410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2590_
timestamp 0
transform -1 0 6190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2591_
timestamp 0
transform 1 0 6430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2592_
timestamp 0
transform -1 0 4410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2593_
timestamp 0
transform 1 0 4930 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2594_
timestamp 0
transform -1 0 8510 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2595_
timestamp 0
transform -1 0 5230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2596_
timestamp 0
transform 1 0 5230 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2597_
timestamp 0
transform 1 0 5410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2598_
timestamp 0
transform -1 0 5150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2599_
timestamp 0
transform -1 0 4950 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2600_
timestamp 0
transform -1 0 4950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2601_
timestamp 0
transform -1 0 5210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2602_
timestamp 0
transform -1 0 8150 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2603_
timestamp 0
transform -1 0 6590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2604_
timestamp 0
transform -1 0 6350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2605_
timestamp 0
transform 1 0 6030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2606_
timestamp 0
transform -1 0 5530 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2607_
timestamp 0
transform 1 0 5690 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2608_
timestamp 0
transform 1 0 5510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2609_
timestamp 0
transform -1 0 5490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2610_
timestamp 0
transform 1 0 4870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2611_
timestamp 0
transform -1 0 5130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2612_
timestamp 0
transform -1 0 5390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2613_
timestamp 0
transform -1 0 1210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2614_
timestamp 0
transform 1 0 2190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2615_
timestamp 0
transform -1 0 2470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2616_
timestamp 0
transform -1 0 2450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2617_
timestamp 0
transform 1 0 1430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2618_
timestamp 0
transform 1 0 850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2619_
timestamp 0
transform -1 0 350 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2620_
timestamp 0
transform -1 0 590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2621_
timestamp 0
transform 1 0 910 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2622_
timestamp 0
transform 1 0 350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2623_
timestamp 0
transform 1 0 2730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2624_
timestamp 0
transform 1 0 1930 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2625_
timestamp 0
transform -1 0 2190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2626_
timestamp 0
transform -1 0 1910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2627_
timestamp 0
transform 1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2628_
timestamp 0
transform 1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2629_
timestamp 0
transform -1 0 310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2630_
timestamp 0
transform 1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2631_
timestamp 0
transform 1 0 4990 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2632_
timestamp 0
transform 1 0 2230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2633_
timestamp 0
transform -1 0 2530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2634_
timestamp 0
transform -1 0 70 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2635_
timestamp 0
transform 1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2636_
timestamp 0
transform 1 0 590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2637_
timestamp 0
transform 1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2638_
timestamp 0
transform 1 0 350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2639_
timestamp 0
transform -1 0 670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2640_
timestamp 0
transform -1 0 70 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2641_
timestamp 0
transform -1 0 70 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2642_
timestamp 0
transform 1 0 1310 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2643_
timestamp 0
transform -1 0 1850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2644_
timestamp 0
transform 1 0 2250 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2645_
timestamp 0
transform -1 0 1990 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2646_
timestamp 0
transform -1 0 1190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2647_
timestamp 0
transform 1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2648_
timestamp 0
transform 1 0 550 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__2649_
timestamp 0
transform 1 0 50 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2650_
timestamp 0
transform -1 0 3650 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2651_
timestamp 0
transform -1 0 3370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2652_
timestamp 0
transform 1 0 590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2653_
timestamp 0
transform 1 0 310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2654_
timestamp 0
transform 1 0 1190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2655_
timestamp 0
transform 1 0 630 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2656_
timestamp 0
transform -1 0 910 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2657_
timestamp 0
transform 1 0 50 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2658_
timestamp 0
transform 1 0 50 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2659_
timestamp 0
transform -1 0 350 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2660_
timestamp 0
transform 1 0 290 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2661_
timestamp 0
transform -1 0 2610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__2662_
timestamp 0
transform -1 0 2550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2663_
timestamp 0
transform -1 0 1970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2664_
timestamp 0
transform 1 0 870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2665_
timestamp 0
transform -1 0 830 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2666_
timestamp 0
transform -1 0 350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2667_
timestamp 0
transform -1 0 570 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2668_
timestamp 0
transform 1 0 1070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2669_
timestamp 0
transform -1 0 2830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2670_
timestamp 0
transform -1 0 2950 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2671_
timestamp 0
transform 1 0 1110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2672_
timestamp 0
transform -1 0 610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2673_
timestamp 0
transform -1 0 570 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2674_
timestamp 0
transform 1 0 830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2675_
timestamp 0
transform 1 0 810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2676_
timestamp 0
transform -1 0 1110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2677_
timestamp 0
transform 1 0 6450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__2678_
timestamp 0
transform -1 0 6370 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2679_
timestamp 0
transform 1 0 6990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2680_
timestamp 0
transform -1 0 6790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2681_
timestamp 0
transform 1 0 7050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2682_
timestamp 0
transform -1 0 6770 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2683_
timestamp 0
transform -1 0 1890 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2684_
timestamp 0
transform -1 0 1710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__2685_
timestamp 0
transform 1 0 1630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2686_
timestamp 0
transform 1 0 1630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2687_
timestamp 0
transform 1 0 1370 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2688_
timestamp 0
transform -1 0 810 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2689_
timestamp 0
transform -1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2690_
timestamp 0
transform 1 0 7290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2691_
timestamp 0
transform -1 0 7130 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2692_
timestamp 0
transform -1 0 5070 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2693_
timestamp 0
transform -1 0 3030 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2694_
timestamp 0
transform -1 0 1330 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2695_
timestamp 0
transform -1 0 1610 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2696_
timestamp 0
transform -1 0 1330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2697_
timestamp 0
transform 1 0 1910 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2698_
timestamp 0
transform -1 0 550 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2699_
timestamp 0
transform 1 0 6310 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2700_
timestamp 0
transform -1 0 7030 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2701_
timestamp 0
transform 1 0 7610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2702_
timestamp 0
transform 1 0 7310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2703_
timestamp 0
transform 1 0 7470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2704_
timestamp 0
transform -1 0 6670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2705_
timestamp 0
transform 1 0 1590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2706_
timestamp 0
transform 1 0 1030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2707_
timestamp 0
transform 1 0 2730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2708_
timestamp 0
transform 1 0 2410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2709_
timestamp 0
transform -1 0 1090 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2710_
timestamp 0
transform -1 0 870 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2711_
timestamp 0
transform -1 0 1150 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2712_
timestamp 0
transform 1 0 2890 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2713_
timestamp 0
transform -1 0 4290 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2714_
timestamp 0
transform -1 0 4710 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2715_
timestamp 0
transform 1 0 3550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2716_
timestamp 0
transform -1 0 4310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2717_
timestamp 0
transform -1 0 5870 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__2718_
timestamp 0
transform -1 0 4110 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2719_
timestamp 0
transform 1 0 3710 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2720_
timestamp 0
transform -1 0 4010 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2721_
timestamp 0
transform -1 0 2170 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2722_
timestamp 0
transform 1 0 2290 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2723_
timestamp 0
transform 1 0 2590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2724_
timestamp 0
transform -1 0 830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2725_
timestamp 0
transform -1 0 5430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2726_
timestamp 0
transform -1 0 6610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2727_
timestamp 0
transform 1 0 3870 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2728_
timestamp 0
transform 1 0 3590 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2729_
timestamp 0
transform -1 0 3550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2730_
timestamp 0
transform 1 0 3150 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2731_
timestamp 0
transform 1 0 2010 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2732_
timestamp 0
transform -1 0 1890 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2733_
timestamp 0
transform 1 0 1430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2734_
timestamp 0
transform -1 0 1730 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2735_
timestamp 0
transform -1 0 3890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2736_
timestamp 0
transform -1 0 4030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2737_
timestamp 0
transform -1 0 4110 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2738_
timestamp 0
transform -1 0 3810 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2739_
timestamp 0
transform -1 0 3250 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2740_
timestamp 0
transform -1 0 3330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2741_
timestamp 0
transform -1 0 1090 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2742_
timestamp 0
transform 1 0 1390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2743_
timestamp 0
transform 1 0 1330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2744_
timestamp 0
transform 1 0 1870 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2745_
timestamp 0
transform 1 0 530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2746_
timestamp 0
transform 1 0 3590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2747_
timestamp 0
transform 1 0 4710 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__2748_
timestamp 0
transform 1 0 4370 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2749_
timestamp 0
transform -1 0 3530 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2750_
timestamp 0
transform -1 0 2970 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2751_
timestamp 0
transform 1 0 2810 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2752_
timestamp 0
transform 1 0 1110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2753_
timestamp 0
transform 1 0 610 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2754_
timestamp 0
transform -1 0 550 0 1 790
box -6 -8 26 268
use FILL  FILL_2__2755_
timestamp 0
transform -1 0 3070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2756_
timestamp 0
transform -1 0 2510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2757_
timestamp 0
transform 1 0 2750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2758_
timestamp 0
transform 1 0 2230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2759_
timestamp 0
transform -1 0 4310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2760_
timestamp 0
transform 1 0 3750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2761_
timestamp 0
transform 1 0 4090 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2762_
timestamp 0
transform -1 0 3830 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2763_
timestamp 0
transform -1 0 2070 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2764_
timestamp 0
transform -1 0 1790 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2765_
timestamp 0
transform -1 0 1710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2766_
timestamp 0
transform -1 0 1970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__2767_
timestamp 0
transform -1 0 1490 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__2768_
timestamp 0
transform 1 0 2150 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2769_
timestamp 0
transform 1 0 1590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__2770_
timestamp 0
transform 1 0 5950 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2771_
timestamp 0
transform 1 0 6490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2772_
timestamp 0
transform 1 0 4930 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__2773_
timestamp 0
transform 1 0 4130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2774_
timestamp 0
transform 1 0 2290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2775_
timestamp 0
transform 1 0 2530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2776_
timestamp 0
transform 1 0 3350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2777_
timestamp 0
transform -1 0 2830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2778_
timestamp 0
transform -1 0 3090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__2779_
timestamp 0
transform -1 0 7130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2780_
timestamp 0
transform -1 0 7370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__2781_
timestamp 0
transform 1 0 7850 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__2782_
timestamp 0
transform 1 0 7730 0 1 270
box -6 -8 26 268
use FILL  FILL_2__2783_
timestamp 0
transform 1 0 9670 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2784_
timestamp 0
transform 1 0 10810 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2785_
timestamp 0
transform 1 0 10190 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2786_
timestamp 0
transform 1 0 9910 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2787_
timestamp 0
transform 1 0 8370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2788_
timestamp 0
transform 1 0 8630 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2789_
timestamp 0
transform 1 0 8150 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2790_
timestamp 0
transform -1 0 7890 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2791_
timestamp 0
transform 1 0 6150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2792_
timestamp 0
transform 1 0 9770 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2793_
timestamp 0
transform 1 0 9970 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2794_
timestamp 0
transform -1 0 10230 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2795_
timestamp 0
transform 1 0 8410 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2796_
timestamp 0
transform 1 0 8390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2797_
timestamp 0
transform 1 0 10790 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2798_
timestamp 0
transform -1 0 9930 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2799_
timestamp 0
transform -1 0 8310 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2800_
timestamp 0
transform -1 0 7710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2801_
timestamp 0
transform 1 0 9650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2802_
timestamp 0
transform -1 0 9970 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2803_
timestamp 0
transform 1 0 8410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2804_
timestamp 0
transform -1 0 8310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2805_
timestamp 0
transform -1 0 10050 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2806_
timestamp 0
transform 1 0 9730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2807_
timestamp 0
transform -1 0 8350 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2808_
timestamp 0
transform -1 0 6590 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2809_
timestamp 0
transform 1 0 8110 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2810_
timestamp 0
transform -1 0 7530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2811_
timestamp 0
transform 1 0 10010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2812_
timestamp 0
transform 1 0 9650 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2813_
timestamp 0
transform 1 0 8230 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2814_
timestamp 0
transform -1 0 8110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2815_
timestamp 0
transform -1 0 8190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2816_
timestamp 0
transform 1 0 9450 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2817_
timestamp 0
transform -1 0 10310 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2818_
timestamp 0
transform 1 0 11130 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2819_
timestamp 0
transform 1 0 10110 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2820_
timestamp 0
transform -1 0 9890 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2821_
timestamp 0
transform -1 0 9750 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2822_
timestamp 0
transform -1 0 7470 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2823_
timestamp 0
transform -1 0 9470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2824_
timestamp 0
transform -1 0 9210 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2825_
timestamp 0
transform 1 0 8670 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2826_
timestamp 0
transform 1 0 8710 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2827_
timestamp 0
transform 1 0 9130 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2828_
timestamp 0
transform 1 0 10250 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2829_
timestamp 0
transform -1 0 9190 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2830_
timestamp 0
transform 1 0 9810 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2831_
timestamp 0
transform 1 0 8990 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2832_
timestamp 0
transform -1 0 8910 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2833_
timestamp 0
transform -1 0 8670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2834_
timestamp 0
transform -1 0 8250 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2835_
timestamp 0
transform -1 0 9270 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2836_
timestamp 0
transform -1 0 7970 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2837_
timestamp 0
transform 1 0 8050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2838_
timestamp 0
transform 1 0 9290 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2839_
timestamp 0
transform 1 0 9550 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2840_
timestamp 0
transform -1 0 9290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2841_
timestamp 0
transform 1 0 8190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2842_
timestamp 0
transform 1 0 11510 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2843_
timestamp 0
transform -1 0 11010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2844_
timestamp 0
transform 1 0 10730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2845_
timestamp 0
transform 1 0 10470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2846_
timestamp 0
transform -1 0 10110 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2847_
timestamp 0
transform 1 0 10310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2848_
timestamp 0
transform -1 0 9590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2849_
timestamp 0
transform 1 0 10890 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__2850_
timestamp 0
transform 1 0 11050 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2851_
timestamp 0
transform 1 0 11290 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2852_
timestamp 0
transform 1 0 11990 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2853_
timestamp 0
transform 1 0 12050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2854_
timestamp 0
transform 1 0 11730 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2855_
timestamp 0
transform 1 0 12010 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2856_
timestamp 0
transform -1 0 9050 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2857_
timestamp 0
transform 1 0 9550 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2858_
timestamp 0
transform -1 0 9850 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2859_
timestamp 0
transform 1 0 10790 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2860_
timestamp 0
transform 1 0 7670 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2861_
timestamp 0
transform 1 0 8350 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2862_
timestamp 0
transform -1 0 7730 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2863_
timestamp 0
transform 1 0 7430 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2864_
timestamp 0
transform 1 0 9670 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2865_
timestamp 0
transform 1 0 8830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2866_
timestamp 0
transform -1 0 6930 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2867_
timestamp 0
transform -1 0 8770 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2868_
timestamp 0
transform -1 0 8490 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2869_
timestamp 0
transform -1 0 8930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2870_
timestamp 0
transform 1 0 8570 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2871_
timestamp 0
transform 1 0 8530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2872_
timestamp 0
transform 1 0 5470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2873_
timestamp 0
transform -1 0 5490 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2874_
timestamp 0
transform 1 0 5410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2875_
timestamp 0
transform -1 0 5770 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2876_
timestamp 0
transform 1 0 5450 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2877_
timestamp 0
transform 1 0 6030 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2878_
timestamp 0
transform -1 0 5770 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2879_
timestamp 0
transform -1 0 8910 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2880_
timestamp 0
transform -1 0 11910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2881_
timestamp 0
transform 1 0 11590 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2882_
timestamp 0
transform -1 0 9190 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2883_
timestamp 0
transform 1 0 8990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2884_
timestamp 0
transform -1 0 9310 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2885_
timestamp 0
transform -1 0 10490 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2886_
timestamp 0
transform 1 0 10450 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2887_
timestamp 0
transform -1 0 8870 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2888_
timestamp 0
transform -1 0 9150 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2889_
timestamp 0
transform 1 0 9430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2890_
timestamp 0
transform -1 0 9790 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__2891_
timestamp 0
transform -1 0 9730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2892_
timestamp 0
transform 1 0 9110 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2893_
timestamp 0
transform -1 0 9270 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2894_
timestamp 0
transform -1 0 11090 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2895_
timestamp 0
transform 1 0 10770 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2896_
timestamp 0
transform -1 0 11050 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2897_
timestamp 0
transform -1 0 10770 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2898_
timestamp 0
transform 1 0 9390 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2899_
timestamp 0
transform -1 0 9690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2900_
timestamp 0
transform 1 0 10370 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2901_
timestamp 0
transform -1 0 10390 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2902_
timestamp 0
transform 1 0 10570 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2903_
timestamp 0
transform -1 0 10690 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2904_
timestamp 0
transform -1 0 9850 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2905_
timestamp 0
transform -1 0 9350 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2906_
timestamp 0
transform -1 0 8510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2907_
timestamp 0
transform -1 0 9070 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2908_
timestamp 0
transform -1 0 10410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2909_
timestamp 0
transform 1 0 11770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2910_
timestamp 0
transform 1 0 10850 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2911_
timestamp 0
transform 1 0 11710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2912_
timestamp 0
transform 1 0 11990 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__2913_
timestamp 0
transform 1 0 10590 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__2914_
timestamp 0
transform -1 0 7770 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2915_
timestamp 0
transform 1 0 10910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2916_
timestamp 0
transform 1 0 11150 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__2917_
timestamp 0
transform 1 0 10650 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2918_
timestamp 0
transform -1 0 10810 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2919_
timestamp 0
transform 1 0 8490 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2920_
timestamp 0
transform 1 0 11190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2921_
timestamp 0
transform 1 0 11710 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__2922_
timestamp 0
transform -1 0 11830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2923_
timestamp 0
transform 1 0 11290 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2924_
timestamp 0
transform 1 0 10210 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2925_
timestamp 0
transform 1 0 9970 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2926_
timestamp 0
transform 1 0 10110 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2927_
timestamp 0
transform -1 0 9950 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2928_
timestamp 0
transform -1 0 10210 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__2929_
timestamp 0
transform -1 0 10330 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__2930_
timestamp 0
transform -1 0 11210 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2931_
timestamp 0
transform -1 0 11470 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__2932_
timestamp 0
transform 1 0 11430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__2933_
timestamp 0
transform 1 0 11390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__2934_
timestamp 0
transform 1 0 11470 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__2935_
timestamp 0
transform 1 0 11550 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2936_
timestamp 0
transform 1 0 10490 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__2937_
timestamp 0
transform -1 0 3490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__2938_
timestamp 0
transform -1 0 7710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2939_
timestamp 0
transform 1 0 6470 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2940_
timestamp 0
transform -1 0 6250 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2941_
timestamp 0
transform -1 0 6170 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2942_
timestamp 0
transform 1 0 5070 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2943_
timestamp 0
transform -1 0 6970 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__2944_
timestamp 0
transform 1 0 5350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2945_
timestamp 0
transform -1 0 6750 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2946_
timestamp 0
transform 1 0 6350 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__2947_
timestamp 0
transform 1 0 7830 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2948_
timestamp 0
transform 1 0 7570 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2949_
timestamp 0
transform 1 0 5670 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__2950_
timestamp 0
transform -1 0 6010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2951_
timestamp 0
transform 1 0 6770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2952_
timestamp 0
transform 1 0 6490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2953_
timestamp 0
transform 1 0 5650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2954_
timestamp 0
transform -1 0 5950 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__2955_
timestamp 0
transform 1 0 7030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2956_
timestamp 0
transform 1 0 6510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__2957_
timestamp 0
transform -1 0 8130 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__2958_
timestamp 0
transform 1 0 6510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__2959_
timestamp 0
transform 1 0 6250 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2960_
timestamp 0
transform -1 0 7130 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2961_
timestamp 0
transform 1 0 6510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2962_
timestamp 0
transform -1 0 6290 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__2963_
timestamp 0
transform -1 0 6590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2964_
timestamp 0
transform 1 0 4650 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2965_
timestamp 0
transform 1 0 5710 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2966_
timestamp 0
transform -1 0 6610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__2967_
timestamp 0
transform -1 0 5030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2968_
timestamp 0
transform -1 0 5290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2969_
timestamp 0
transform 1 0 4370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2970_
timestamp 0
transform 1 0 4730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2971_
timestamp 0
transform 1 0 4610 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2972_
timestamp 0
transform -1 0 6050 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2973_
timestamp 0
transform -1 0 6310 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2974_
timestamp 0
transform -1 0 6310 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2975_
timestamp 0
transform 1 0 5770 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2976_
timestamp 0
transform -1 0 4690 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2977_
timestamp 0
transform -1 0 4950 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2978_
timestamp 0
transform 1 0 5210 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__2979_
timestamp 0
transform 1 0 5490 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__2980_
timestamp 0
transform -1 0 7370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2981_
timestamp 0
transform -1 0 6330 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2982_
timestamp 0
transform -1 0 6610 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__2983_
timestamp 0
transform 1 0 7130 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2984_
timestamp 0
transform 1 0 6530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__2985_
timestamp 0
transform -1 0 6870 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2986_
timestamp 0
transform 1 0 6570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2987_
timestamp 0
transform 1 0 6010 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2988_
timestamp 0
transform -1 0 6290 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__2989_
timestamp 0
transform -1 0 7870 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2990_
timestamp 0
transform 1 0 6990 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__2991_
timestamp 0
transform -1 0 6850 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2992_
timestamp 0
transform -1 0 5150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__2993_
timestamp 0
transform -1 0 6010 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2994_
timestamp 0
transform 1 0 5470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2995_
timestamp 0
transform 1 0 6550 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2996_
timestamp 0
transform 1 0 6270 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__2997_
timestamp 0
transform 1 0 5990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2998_
timestamp 0
transform -1 0 5730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__2999_
timestamp 0
transform 1 0 6390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3000_
timestamp 0
transform -1 0 5730 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__3001_
timestamp 0
transform 1 0 4950 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3002_
timestamp 0
transform -1 0 5450 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__3003_
timestamp 0
transform -1 0 5810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3004_
timestamp 0
transform -1 0 5230 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3005_
timestamp 0
transform -1 0 5490 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3006_
timestamp 0
transform -1 0 7390 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3007_
timestamp 0
transform 1 0 6810 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3008_
timestamp 0
transform 1 0 8610 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3009_
timestamp 0
transform 1 0 8070 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3010_
timestamp 0
transform 1 0 7090 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3011_
timestamp 0
transform -1 0 7190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3012_
timestamp 0
transform -1 0 7070 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3013_
timestamp 0
transform -1 0 7810 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3014_
timestamp 0
transform 1 0 7010 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3015_
timestamp 0
transform -1 0 7290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3016_
timestamp 0
transform -1 0 6050 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3017_
timestamp 0
transform -1 0 6850 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3018_
timestamp 0
transform -1 0 6530 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3019_
timestamp 0
transform -1 0 6790 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3020_
timestamp 0
transform 1 0 5430 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__3021_
timestamp 0
transform 1 0 5870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3022_
timestamp 0
transform 1 0 5670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__3023_
timestamp 0
transform -1 0 6750 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3024_
timestamp 0
transform -1 0 6670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3025_
timestamp 0
transform 1 0 5950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__3026_
timestamp 0
transform 1 0 5370 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__3027_
timestamp 0
transform -1 0 5470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3028_
timestamp 0
transform 1 0 5950 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3029_
timestamp 0
transform 1 0 6710 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3030_
timestamp 0
transform 1 0 4850 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__3031_
timestamp 0
transform 1 0 4390 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3032_
timestamp 0
transform -1 0 5170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3033_
timestamp 0
transform 1 0 5430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3034_
timestamp 0
transform -1 0 3370 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3035_
timestamp 0
transform -1 0 3930 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3036_
timestamp 0
transform -1 0 3430 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3037_
timestamp 0
transform -1 0 3310 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3038_
timestamp 0
transform 1 0 3530 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3039_
timestamp 0
transform -1 0 3030 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3040_
timestamp 0
transform 1 0 2910 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3041_
timestamp 0
transform 1 0 3150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3042_
timestamp 0
transform -1 0 3710 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3043_
timestamp 0
transform -1 0 3810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3044_
timestamp 0
transform -1 0 3570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3045_
timestamp 0
transform 1 0 4370 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3046_
timestamp 0
transform 1 0 4090 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3047_
timestamp 0
transform -1 0 3050 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3048_
timestamp 0
transform 1 0 3090 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3049_
timestamp 0
transform -1 0 2790 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3050_
timestamp 0
transform 1 0 2830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3051_
timestamp 0
transform 1 0 2570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3052_
timestamp 0
transform 1 0 2470 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3053_
timestamp 0
transform 1 0 3230 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3054_
timestamp 0
transform -1 0 3510 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3055_
timestamp 0
transform 1 0 3330 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3056_
timestamp 0
transform -1 0 3590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3057_
timestamp 0
transform 1 0 3790 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3058_
timestamp 0
transform 1 0 3970 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3059_
timestamp 0
transform 1 0 4250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3060_
timestamp 0
transform 1 0 4090 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3061_
timestamp 0
transform 1 0 3570 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3062_
timestamp 0
transform -1 0 3810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3063_
timestamp 0
transform -1 0 5050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__3064_
timestamp 0
transform 1 0 4910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__3065_
timestamp 0
transform -1 0 4650 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3066_
timestamp 0
transform 1 0 4550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3067_
timestamp 0
transform -1 0 3650 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3068_
timestamp 0
transform -1 0 3390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3069_
timestamp 0
transform 1 0 3590 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3070_
timestamp 0
transform -1 0 4490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__3071_
timestamp 0
transform 1 0 4210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__3072_
timestamp 0
transform -1 0 4150 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3073_
timestamp 0
transform -1 0 4410 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3074_
timestamp 0
transform 1 0 5690 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3075_
timestamp 0
transform 1 0 5410 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3076_
timestamp 0
transform 1 0 3650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3077_
timestamp 0
transform 1 0 3970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3078_
timestamp 0
transform 1 0 4030 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3079_
timestamp 0
transform -1 0 4110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3080_
timestamp 0
transform 1 0 6250 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3081_
timestamp 0
transform -1 0 6910 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3082_
timestamp 0
transform 1 0 6610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3083_
timestamp 0
transform -1 0 3790 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3084_
timestamp 0
transform 1 0 3490 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3085_
timestamp 0
transform 1 0 3110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3086_
timestamp 0
transform -1 0 2830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3087_
timestamp 0
transform 1 0 4310 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3088_
timestamp 0
transform -1 0 4910 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3089_
timestamp 0
transform 1 0 3390 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3090_
timestamp 0
transform -1 0 3670 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3091_
timestamp 0
transform -1 0 6210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3092_
timestamp 0
transform 1 0 5430 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3093_
timestamp 0
transform 1 0 5690 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3094_
timestamp 0
transform 1 0 5410 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3095_
timestamp 0
transform -1 0 4610 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3096_
timestamp 0
transform 1 0 4310 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3097_
timestamp 0
transform -1 0 4070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3098_
timestamp 0
transform 1 0 3770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3099_
timestamp 0
transform -1 0 3830 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3100_
timestamp 0
transform -1 0 3650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3101_
timestamp 0
transform 1 0 4870 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3102_
timestamp 0
transform -1 0 5170 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3103_
timestamp 0
transform -1 0 4550 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3104_
timestamp 0
transform -1 0 4830 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3105_
timestamp 0
transform 1 0 5610 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3106_
timestamp 0
transform -1 0 5910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3107_
timestamp 0
transform -1 0 4010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3108_
timestamp 0
transform 1 0 3710 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3109_
timestamp 0
transform 1 0 6190 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3110_
timestamp 0
transform 1 0 3870 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3111_
timestamp 0
transform 1 0 5730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3112_
timestamp 0
transform -1 0 5150 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3113_
timestamp 0
transform -1 0 4610 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3114_
timestamp 0
transform 1 0 4310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3115_
timestamp 0
transform 1 0 4830 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3116_
timestamp 0
transform 1 0 3770 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3117_
timestamp 0
transform 1 0 4390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3118_
timestamp 0
transform -1 0 4690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3119_
timestamp 0
transform 1 0 4870 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3120_
timestamp 0
transform 1 0 4570 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3121_
timestamp 0
transform 1 0 5170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3122_
timestamp 0
transform 1 0 5450 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3123_
timestamp 0
transform 1 0 5430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3124_
timestamp 0
transform -1 0 5730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3125_
timestamp 0
transform -1 0 4090 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3126_
timestamp 0
transform 1 0 3790 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3127_
timestamp 0
transform 1 0 6450 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3128_
timestamp 0
transform 1 0 6010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3129_
timestamp 0
transform 1 0 5410 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3130_
timestamp 0
transform -1 0 3330 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3131_
timestamp 0
transform -1 0 3570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3132_
timestamp 0
transform 1 0 4670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3133_
timestamp 0
transform 1 0 3910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3134_
timestamp 0
transform 1 0 5090 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3135_
timestamp 0
transform 1 0 4790 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3136_
timestamp 0
transform 1 0 5690 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3137_
timestamp 0
transform 1 0 5410 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3138_
timestamp 0
transform 1 0 5690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3139_
timestamp 0
transform 1 0 5410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3140_
timestamp 0
transform -1 0 5610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3141_
timestamp 0
transform -1 0 5870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3142_
timestamp 0
transform -1 0 4210 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3143_
timestamp 0
transform -1 0 4470 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3144_
timestamp 0
transform 1 0 11550 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__3145_
timestamp 0
transform 1 0 11790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__3146_
timestamp 0
transform -1 0 11850 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__3147_
timestamp 0
transform 1 0 9470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__3148_
timestamp 0
transform -1 0 11850 0 1 790
box -6 -8 26 268
use FILL  FILL_2__3149_
timestamp 0
transform -1 0 11470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3150_
timestamp 0
transform -1 0 11750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3151_
timestamp 0
transform -1 0 10690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3152_
timestamp 0
transform 1 0 9330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3153_
timestamp 0
transform -1 0 9630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3154_
timestamp 0
transform -1 0 10150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3155_
timestamp 0
transform -1 0 10270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3156_
timestamp 0
transform -1 0 8910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__3157_
timestamp 0
transform -1 0 8950 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__3158_
timestamp 0
transform -1 0 8670 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__3159_
timestamp 0
transform -1 0 8650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__3160_
timestamp 0
transform 1 0 10490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3161_
timestamp 0
transform 1 0 10210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3162_
timestamp 0
transform -1 0 9750 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3163_
timestamp 0
transform 1 0 9470 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3164_
timestamp 0
transform -1 0 8950 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3165_
timestamp 0
transform -1 0 7170 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3166_
timestamp 0
transform 1 0 7570 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__3167_
timestamp 0
transform 1 0 7430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3168_
timestamp 0
transform 1 0 7590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3169_
timestamp 0
transform -1 0 8670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3170_
timestamp 0
transform -1 0 8390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3171_
timestamp 0
transform -1 0 9110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3172_
timestamp 0
transform -1 0 8110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3173_
timestamp 0
transform 1 0 8370 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3174_
timestamp 0
transform 1 0 7850 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3175_
timestamp 0
transform -1 0 7830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3176_
timestamp 0
transform -1 0 7550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3177_
timestamp 0
transform -1 0 11830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__3178_
timestamp 0
transform -1 0 11770 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3179_
timestamp 0
transform 1 0 12030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3180_
timestamp 0
transform 1 0 12090 0 1 790
box -6 -8 26 268
use FILL  FILL_2__3181_
timestamp 0
transform 1 0 12070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__3182_
timestamp 0
transform -1 0 11290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3183_
timestamp 0
transform 1 0 11550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3184_
timestamp 0
transform 1 0 11830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3185_
timestamp 0
transform 1 0 11850 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3186_
timestamp 0
transform 1 0 12030 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3187_
timestamp 0
transform 1 0 9890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__3188_
timestamp 0
transform 1 0 10770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3189_
timestamp 0
transform -1 0 11030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__3190_
timestamp 0
transform 1 0 11070 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3191_
timestamp 0
transform 1 0 11010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3192_
timestamp 0
transform -1 0 10730 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3193_
timestamp 0
transform 1 0 10150 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3194_
timestamp 0
transform 1 0 10770 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__3195_
timestamp 0
transform -1 0 10510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3196_
timestamp 0
transform 1 0 10410 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3197_
timestamp 0
transform -1 0 7270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3198_
timestamp 0
transform -1 0 4630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3199_
timestamp 0
transform 1 0 2790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__3200_
timestamp 0
transform 1 0 4770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__3201_
timestamp 0
transform 1 0 4490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__3202_
timestamp 0
transform 1 0 1550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__3203_
timestamp 0
transform 1 0 1510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3204_
timestamp 0
transform 1 0 1470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__3205_
timestamp 0
transform 1 0 1030 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__3206_
timestamp 0
transform 1 0 1450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__3207_
timestamp 0
transform -1 0 1590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__3208_
timestamp 0
transform -1 0 930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__3209_
timestamp 0
transform -1 0 630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__3210_
timestamp 0
transform -1 0 4290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__3211_
timestamp 0
transform 1 0 4230 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__3212_
timestamp 0
transform 1 0 1190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__3213_
timestamp 0
transform 1 0 1090 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__3214_
timestamp 0
transform -1 0 2370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3215_
timestamp 0
transform 1 0 1790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3216_
timestamp 0
transform 1 0 5730 0 1 270
box -6 -8 26 268
use FILL  FILL_2__3217_
timestamp 0
transform -1 0 6030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__3218_
timestamp 0
transform 1 0 6070 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3219_
timestamp 0
transform -1 0 6350 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3220_
timestamp 0
transform 1 0 3690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3221_
timestamp 0
transform -1 0 3970 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3222_
timestamp 0
transform -1 0 3570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3223_
timestamp 0
transform 1 0 3290 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__3224_
timestamp 0
transform -1 0 3270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3225_
timestamp 0
transform 1 0 5410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__3226_
timestamp 0
transform 1 0 5130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__3227_
timestamp 0
transform -1 0 4250 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3228_
timestamp 0
transform -1 0 4450 0 1 270
box -6 -8 26 268
use FILL  FILL_2__3229_
timestamp 0
transform 1 0 2690 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__3230_
timestamp 0
transform -1 0 2730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__3231_
timestamp 0
transform 1 0 5970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__3232_
timestamp 0
transform 1 0 5950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__3364_
timestamp 0
transform 1 0 5230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3365_
timestamp 0
transform 1 0 4430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3366_
timestamp 0
transform 1 0 4910 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__3367_
timestamp 0
transform -1 0 4710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3368_
timestamp 0
transform -1 0 4970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3369_
timestamp 0
transform -1 0 5530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3370_
timestamp 0
transform 1 0 2670 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3371_
timestamp 0
transform 1 0 2170 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3372_
timestamp 0
transform -1 0 2290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3373_
timestamp 0
transform -1 0 3950 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3374_
timestamp 0
transform -1 0 2270 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3375_
timestamp 0
transform 1 0 2270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3376_
timestamp 0
transform -1 0 2930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3377_
timestamp 0
transform 1 0 2390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3378_
timestamp 0
transform -1 0 2250 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3379_
timestamp 0
transform -1 0 1410 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3380_
timestamp 0
transform 1 0 1190 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3381_
timestamp 0
transform -1 0 1450 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3382_
timestamp 0
transform -1 0 1910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3383_
timestamp 0
transform -1 0 1470 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3384_
timestamp 0
transform 1 0 1730 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3385_
timestamp 0
transform 1 0 1430 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3386_
timestamp 0
transform -1 0 2010 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3387_
timestamp 0
transform 1 0 2270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3388_
timestamp 0
transform -1 0 610 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3389_
timestamp 0
transform 1 0 2470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3390_
timestamp 0
transform 1 0 3290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3391_
timestamp 0
transform 1 0 3010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3392_
timestamp 0
transform -1 0 2850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3393_
timestamp 0
transform 1 0 2250 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3394_
timestamp 0
transform 1 0 650 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3395_
timestamp 0
transform -1 0 610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3396_
timestamp 0
transform -1 0 350 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3397_
timestamp 0
transform -1 0 370 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3398_
timestamp 0
transform -1 0 70 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3399_
timestamp 0
transform 1 0 50 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3400_
timestamp 0
transform -1 0 850 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3401_
timestamp 0
transform -1 0 1430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3402_
timestamp 0
transform 1 0 1410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3403_
timestamp 0
transform 1 0 1130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3404_
timestamp 0
transform -1 0 70 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3405_
timestamp 0
transform -1 0 330 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3406_
timestamp 0
transform -1 0 70 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3407_
timestamp 0
transform -1 0 350 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3408_
timestamp 0
transform -1 0 70 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3409_
timestamp 0
transform -1 0 70 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3410_
timestamp 0
transform 1 0 1390 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3411_
timestamp 0
transform 1 0 1110 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3412_
timestamp 0
transform -1 0 590 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3413_
timestamp 0
transform 1 0 330 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3414_
timestamp 0
transform 1 0 590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2__3415_
timestamp 0
transform -1 0 910 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3416_
timestamp 0
transform 1 0 590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3417_
timestamp 0
transform -1 0 630 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3418_
timestamp 0
transform -1 0 330 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3419_
timestamp 0
transform -1 0 1150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3420_
timestamp 0
transform 1 0 850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3421_
timestamp 0
transform 1 0 1150 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3422_
timestamp 0
transform 1 0 870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3423_
timestamp 0
transform 1 0 1170 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3424_
timestamp 0
transform -1 0 1190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3425_
timestamp 0
transform -1 0 910 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3426_
timestamp 0
transform 1 0 890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2__3427_
timestamp 0
transform -1 0 1410 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3428_
timestamp 0
transform 1 0 1090 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3429_
timestamp 0
transform -1 0 870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3430_
timestamp 0
transform 1 0 1390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3431_
timestamp 0
transform 1 0 1110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3432_
timestamp 0
transform -1 0 910 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3433_
timestamp 0
transform -1 0 70 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3434_
timestamp 0
transform -1 0 650 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3435_
timestamp 0
transform -1 0 930 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3436_
timestamp 0
transform -1 0 870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3437_
timestamp 0
transform 1 0 1690 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3438_
timestamp 0
transform 1 0 1150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3439_
timestamp 0
transform -1 0 1430 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3440_
timestamp 0
transform 1 0 1150 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3441_
timestamp 0
transform -1 0 590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3442_
timestamp 0
transform 1 0 1170 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3443_
timestamp 0
transform 1 0 1090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3444_
timestamp 0
transform -1 0 1990 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3445_
timestamp 0
transform 1 0 1670 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3446_
timestamp 0
transform 1 0 2030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3447_
timestamp 0
transform 1 0 1930 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3448_
timestamp 0
transform -1 0 1730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3449_
timestamp 0
transform 1 0 1410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3450_
timestamp 0
transform -1 0 870 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3451_
timestamp 0
transform 1 0 1130 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3452_
timestamp 0
transform 1 0 830 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3453_
timestamp 0
transform -1 0 2150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3454_
timestamp 0
transform 1 0 3070 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3455_
timestamp 0
transform -1 0 2010 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3456_
timestamp 0
transform -1 0 1670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3457_
timestamp 0
transform -1 0 2850 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3458_
timestamp 0
transform -1 0 1710 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3459_
timestamp 0
transform -1 0 1650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3460_
timestamp 0
transform 1 0 1690 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3461_
timestamp 0
transform -1 0 1910 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3462_
timestamp 0
transform -1 0 1670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3463_
timestamp 0
transform -1 0 1430 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3464_
timestamp 0
transform 1 0 1150 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3465_
timestamp 0
transform -1 0 1410 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3466_
timestamp 0
transform 1 0 1950 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3467_
timestamp 0
transform 1 0 1950 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3468_
timestamp 0
transform 1 0 2710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3469_
timestamp 0
transform 1 0 2570 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3470_
timestamp 0
transform -1 0 2470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3471_
timestamp 0
transform 1 0 2290 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3472_
timestamp 0
transform -1 0 2190 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3473_
timestamp 0
transform 1 0 1430 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3474_
timestamp 0
transform -1 0 1690 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3475_
timestamp 0
transform 1 0 1170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3476_
timestamp 0
transform -1 0 910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3477_
timestamp 0
transform 1 0 330 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3478_
timestamp 0
transform -1 0 310 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3479_
timestamp 0
transform -1 0 70 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3480_
timestamp 0
transform -1 0 70 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3481_
timestamp 0
transform -1 0 70 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3482_
timestamp 0
transform 1 0 590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3483_
timestamp 0
transform -1 0 310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3484_
timestamp 0
transform 1 0 1930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3485_
timestamp 0
transform -1 0 1990 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3486_
timestamp 0
transform -1 0 1370 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3487_
timestamp 0
transform -1 0 1690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3488_
timestamp 0
transform -1 0 1490 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3489_
timestamp 0
transform 1 0 1430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3490_
timestamp 0
transform 1 0 1110 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3491_
timestamp 0
transform -1 0 1190 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3492_
timestamp 0
transform 1 0 1090 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3493_
timestamp 0
transform -1 0 910 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3494_
timestamp 0
transform 1 0 830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3495_
timestamp 0
transform -1 0 590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3496_
timestamp 0
transform 1 0 350 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3497_
timestamp 0
transform -1 0 310 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3498_
timestamp 0
transform 1 0 610 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3499_
timestamp 0
transform -1 0 670 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3500_
timestamp 0
transform 1 0 610 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3501_
timestamp 0
transform 1 0 850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3502_
timestamp 0
transform -1 0 370 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3503_
timestamp 0
transform -1 0 350 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3504_
timestamp 0
transform -1 0 590 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3505_
timestamp 0
transform -1 0 350 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3506_
timestamp 0
transform -1 0 70 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3507_
timestamp 0
transform -1 0 70 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3508_
timestamp 0
transform 1 0 590 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3509_
timestamp 0
transform -1 0 850 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3510_
timestamp 0
transform -1 0 350 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3511_
timestamp 0
transform -1 0 70 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3512_
timestamp 0
transform 1 0 550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3513_
timestamp 0
transform -1 0 370 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3514_
timestamp 0
transform -1 0 310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3515_
timestamp 0
transform -1 0 70 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3516_
timestamp 0
transform -1 0 70 0 1 10150
box -6 -8 26 268
use FILL  FILL_2__3517_
timestamp 0
transform 1 0 610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3518_
timestamp 0
transform 1 0 830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3519_
timestamp 0
transform 1 0 2530 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3520_
timestamp 0
transform 1 0 2810 0 1 9110
box -6 -8 26 268
use FILL  FILL_2__3521_
timestamp 0
transform 1 0 3290 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3522_
timestamp 0
transform 1 0 2990 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3523_
timestamp 0
transform 1 0 2550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3524_
timestamp 0
transform -1 0 930 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3525_
timestamp 0
transform -1 0 70 0 1 10670
box -6 -8 26 268
use FILL  FILL_2__3526_
timestamp 0
transform -1 0 70 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3527_
timestamp 0
transform -1 0 570 0 1 11190
box -6 -8 26 268
use FILL  FILL_2__3528_
timestamp 0
transform -1 0 590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_2__3529_
timestamp 0
transform -1 0 70 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2__3530_
timestamp 0
transform -1 0 70 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3531_
timestamp 0
transform 1 0 50 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3532_
timestamp 0
transform 1 0 290 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3533_
timestamp 0
transform -1 0 70 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3534_
timestamp 0
transform -1 0 590 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3535_
timestamp 0
transform -1 0 350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2__3536_
timestamp 0
transform -1 0 330 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3537_
timestamp 0
transform -1 0 1690 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3538_
timestamp 0
transform 1 0 2450 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3539_
timestamp 0
transform -1 0 2550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3540_
timestamp 0
transform -1 0 2290 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3541_
timestamp 0
transform -1 0 2010 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3542_
timestamp 0
transform -1 0 2190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3543_
timestamp 0
transform 1 0 1590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3544_
timestamp 0
transform 1 0 1950 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3545_
timestamp 0
transform 1 0 1750 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3546_
timestamp 0
transform 1 0 1870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2__3547_
timestamp 0
transform -1 0 2530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3548_
timestamp 0
transform 1 0 2230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2__3549_
timestamp 0
transform -1 0 2330 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3550_
timestamp 0
transform 1 0 2030 0 1 11710
box -6 -8 26 268
use FILL  FILL_2__3551_
timestamp 0
transform -1 0 2510 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3552_
timestamp 0
transform 1 0 2210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2__3553_
timestamp 0
transform -1 0 1750 0 1 8070
box -6 -8 26 268
use FILL  FILL_2__3554_
timestamp 0
transform 1 0 890 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3555_
timestamp 0
transform 1 0 290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3556_
timestamp 0
transform 1 0 1150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2__3557_
timestamp 0
transform -1 0 3050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3558_
timestamp 0
transform 1 0 2750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2__3559_
timestamp 0
transform -1 0 2510 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3560_
timestamp 0
transform 1 0 2210 0 1 9630
box -6 -8 26 268
use FILL  FILL_2__3561_
timestamp 0
transform -1 0 1930 0 1 7550
box -6 -8 26 268
use FILL  FILL_2__3562_
timestamp 0
transform -1 0 2750 0 1 8590
box -6 -8 26 268
use FILL  FILL_2__3563_
timestamp 0
transform 1 0 2150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2__3564_
timestamp 0
transform 1 0 2430 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3565_
timestamp 0
transform -1 0 1430 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3566_
timestamp 0
transform -1 0 1690 0 1 7030
box -6 -8 26 268
use FILL  FILL_2__3579_
timestamp 0
transform -1 0 5030 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3580_
timestamp 0
transform -1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__3581_
timestamp 0
transform -1 0 3450 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3582_
timestamp 0
transform -1 0 3190 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3583_
timestamp 0
transform -1 0 5310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__3584_
timestamp 0
transform 1 0 4490 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3585_
timestamp 0
transform 1 0 2910 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3586_
timestamp 0
transform -1 0 5830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__3587_
timestamp 0
transform 1 0 50 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3588_
timestamp 0
transform -1 0 70 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__3589_
timestamp 0
transform -1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__3590_
timestamp 0
transform -1 0 70 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__3591_
timestamp 0
transform -1 0 350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3592_
timestamp 0
transform -1 0 70 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__3593_
timestamp 0
transform -1 0 4770 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3594_
timestamp 0
transform 1 0 5810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__3595_
timestamp 0
transform 1 0 5550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__3596_
timestamp 0
transform -1 0 850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3597_
timestamp 0
transform -1 0 70 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__3598_
timestamp 0
transform -1 0 330 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__3599_
timestamp 0
transform -1 0 70 0 1 6510
box -6 -8 26 268
use FILL  FILL_2__3600_
timestamp 0
transform -1 0 70 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__3601_
timestamp 0
transform -1 0 70 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__3602_
timestamp 0
transform -1 0 1690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__3603_
timestamp 0
transform 1 0 6850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform 1 0 7870 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 9370 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform 1 0 8130 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform 1 0 10990 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert4
timestamp 0
transform 1 0 590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert5
timestamp 0
transform -1 0 12070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform -1 0 9570 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert7
timestamp 0
transform 1 0 7030 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 850 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert9
timestamp 0
transform 1 0 10110 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert10
timestamp 0
transform -1 0 890 0 1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform -1 0 5970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform 1 0 11530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform -1 0 6150 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform 1 0 6770 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform -1 0 3310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform -1 0 3930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform 1 0 7170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform -1 0 6990 0 1 11190
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform 1 0 5310 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform 1 0 8550 0 1 11190
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform -1 0 8470 0 -1 7550
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 1430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform 1 0 3410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform -1 0 4310 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform 1 0 8150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert26
timestamp 0
transform 1 0 5090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert27
timestamp 0
transform -1 0 1230 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert39
timestamp 0
transform 1 0 6310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert40
timestamp 0
transform 1 0 7670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert41
timestamp 0
transform -1 0 8810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert42
timestamp 0
transform -1 0 6950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert43
timestamp 0
transform -1 0 8850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert44
timestamp 0
transform -1 0 8970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert45
timestamp 0
transform 1 0 11030 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert46
timestamp 0
transform 1 0 9470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert47
timestamp 0
transform 1 0 9190 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert48
timestamp 0
transform 1 0 6930 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert49
timestamp 0
transform 1 0 7190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert50
timestamp 0
transform -1 0 7570 0 1 9110
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert51
timestamp 0
transform 1 0 7530 0 1 10150
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert52
timestamp 0
transform 1 0 8930 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert53
timestamp 0
transform 1 0 9970 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert54
timestamp 0
transform 1 0 8810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert55
timestamp 0
transform 1 0 8670 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert56
timestamp 0
transform -1 0 2210 0 1 8590
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert57
timestamp 0
transform 1 0 2510 0 1 11190
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert58
timestamp 0
transform 1 0 2650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert59
timestamp 0
transform -1 0 2210 0 1 10670
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert60
timestamp 0
transform -1 0 10470 0 1 7550
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert61
timestamp 0
transform 1 0 10530 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert62
timestamp 0
transform 1 0 10490 0 1 8070
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert63
timestamp 0
transform -1 0 9150 0 1 7550
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert64
timestamp 0
transform -1 0 8590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert65
timestamp 0
transform 1 0 5190 0 1 270
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert66
timestamp 0
transform 1 0 5710 0 1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert67
timestamp 0
transform -1 0 3010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert68
timestamp 0
transform 1 0 3130 0 1 270
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert69
timestamp 0
transform -1 0 6630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert70
timestamp 0
transform 1 0 8570 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert71
timestamp 0
transform -1 0 9230 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert72
timestamp 0
transform -1 0 6750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert73
timestamp 0
transform 1 0 8910 0 -1 7030
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert74
timestamp 0
transform 1 0 10770 0 1 7030
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert75
timestamp 0
transform 1 0 2550 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert76
timestamp 0
transform -1 0 3050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert77
timestamp 0
transform 1 0 10430 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert78
timestamp 0
transform 1 0 9290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert79
timestamp 0
transform -1 0 8330 0 1 7550
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert80
timestamp 0
transform 1 0 7130 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert81
timestamp 0
transform 1 0 7590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert82
timestamp 0
transform -1 0 7570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert83
timestamp 0
transform -1 0 7350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert84
timestamp 0
transform 1 0 9410 0 1 8590
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert85
timestamp 0
transform -1 0 8890 0 1 8590
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert86
timestamp 0
transform -1 0 9490 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert87
timestamp 0
transform 1 0 9390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert88
timestamp 0
transform -1 0 10730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert89
timestamp 0
transform 1 0 9370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert90
timestamp 0
transform 1 0 5350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert91
timestamp 0
transform -1 0 4890 0 1 10670
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert92
timestamp 0
transform -1 0 4730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert93
timestamp 0
transform 1 0 5150 0 1 10150
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert94
timestamp 0
transform -1 0 11310 0 1 9630
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert95
timestamp 0
transform -1 0 11350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert96
timestamp 0
transform -1 0 10070 0 1 11710
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert97
timestamp 0
transform 1 0 11430 0 1 11710
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert28
timestamp 0
transform -1 0 6010 0 -1 11710
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert29
timestamp 0
transform -1 0 2190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert30
timestamp 0
transform 1 0 4530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert31
timestamp 0
transform -1 0 3230 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert32
timestamp 0
transform 1 0 7130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert33
timestamp 0
transform 1 0 5710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert34
timestamp 0
transform -1 0 2470 0 1 10670
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert35
timestamp 0
transform -1 0 5230 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert36
timestamp 0
transform -1 0 2350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert37
timestamp 0
transform 1 0 7370 0 -1 12230
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert38
timestamp 0
transform -1 0 4350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__1688_
timestamp 0
transform -1 0 890 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1689_
timestamp 0
transform -1 0 350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1690_
timestamp 0
transform -1 0 610 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1691_
timestamp 0
transform 1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1692_
timestamp 0
transform -1 0 330 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1693_
timestamp 0
transform 1 0 570 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1694_
timestamp 0
transform -1 0 5570 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1695_
timestamp 0
transform -1 0 350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1696_
timestamp 0
transform -1 0 350 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1697_
timestamp 0
transform -1 0 1470 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__1698_
timestamp 0
transform -1 0 3410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1699_
timestamp 0
transform 1 0 2850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1700_
timestamp 0
transform -1 0 3890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__1701_
timestamp 0
transform -1 0 590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1702_
timestamp 0
transform -1 0 590 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1703_
timestamp 0
transform 1 0 3230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1704_
timestamp 0
transform -1 0 370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1705_
timestamp 0
transform 1 0 70 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1706_
timestamp 0
transform -1 0 3850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1707_
timestamp 0
transform -1 0 610 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1708_
timestamp 0
transform 1 0 610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1709_
timestamp 0
transform 1 0 4130 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1710_
timestamp 0
transform -1 0 5610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1711_
timestamp 0
transform 1 0 5150 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1712_
timestamp 0
transform 1 0 7290 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1713_
timestamp 0
transform -1 0 9670 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1714_
timestamp 0
transform -1 0 9870 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1715_
timestamp 0
transform -1 0 8550 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1716_
timestamp 0
transform 1 0 11310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1717_
timestamp 0
transform 1 0 11110 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1718_
timestamp 0
transform 1 0 11930 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1719_
timestamp 0
transform -1 0 8810 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1720_
timestamp 0
transform -1 0 10130 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1721_
timestamp 0
transform -1 0 10150 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1722_
timestamp 0
transform -1 0 9910 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1723_
timestamp 0
transform 1 0 10010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1724_
timestamp 0
transform 1 0 9230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1725_
timestamp 0
transform 1 0 9070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1726_
timestamp 0
transform 1 0 10170 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1727_
timestamp 0
transform -1 0 8790 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1728_
timestamp 0
transform 1 0 11570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1729_
timestamp 0
transform 1 0 10170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1730_
timestamp 0
transform 1 0 8350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1731_
timestamp 0
transform 1 0 8590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1732_
timestamp 0
transform -1 0 7790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1733_
timestamp 0
transform 1 0 9730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1734_
timestamp 0
transform 1 0 7430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1735_
timestamp 0
transform 1 0 10870 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1736_
timestamp 0
transform -1 0 10670 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1737_
timestamp 0
transform -1 0 10930 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1738_
timestamp 0
transform -1 0 10310 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1739_
timestamp 0
transform -1 0 10310 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1740_
timestamp 0
transform 1 0 10530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1741_
timestamp 0
transform -1 0 8430 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1742_
timestamp 0
transform -1 0 8330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1743_
timestamp 0
transform -1 0 9890 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1744_
timestamp 0
transform 1 0 9770 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1745_
timestamp 0
transform -1 0 9470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1746_
timestamp 0
transform 1 0 11330 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1747_
timestamp 0
transform 1 0 10810 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1748_
timestamp 0
transform 1 0 7530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1749_
timestamp 0
transform 1 0 7950 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1750_
timestamp 0
transform -1 0 8070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1751_
timestamp 0
transform 1 0 7470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1752_
timestamp 0
transform -1 0 8890 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1753_
timestamp 0
transform 1 0 9750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1754_
timestamp 0
transform -1 0 8290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1755_
timestamp 0
transform -1 0 8870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__1756_
timestamp 0
transform -1 0 11210 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1757_
timestamp 0
transform 1 0 11070 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1758_
timestamp 0
transform -1 0 9130 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1759_
timestamp 0
transform -1 0 7370 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__1760_
timestamp 0
transform 1 0 8870 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__1761_
timestamp 0
transform -1 0 9590 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1762_
timestamp 0
transform 1 0 10610 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1763_
timestamp 0
transform -1 0 9050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1764_
timestamp 0
transform 1 0 11310 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1765_
timestamp 0
transform 1 0 8130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1766_
timestamp 0
transform 1 0 8510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1767_
timestamp 0
transform 1 0 9210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__1768_
timestamp 0
transform 1 0 8070 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__1769_
timestamp 0
transform 1 0 8590 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__1770_
timestamp 0
transform 1 0 9030 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__1771_
timestamp 0
transform 1 0 8990 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__1772_
timestamp 0
transform 1 0 8710 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__1773_
timestamp 0
transform 1 0 10790 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1774_
timestamp 0
transform 1 0 10790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1775_
timestamp 0
transform 1 0 10030 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1776_
timestamp 0
transform -1 0 8030 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1777_
timestamp 0
transform 1 0 8070 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1778_
timestamp 0
transform -1 0 7550 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1779_
timestamp 0
transform 1 0 5690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1780_
timestamp 0
transform -1 0 4090 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1781_
timestamp 0
transform -1 0 10810 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1782_
timestamp 0
transform 1 0 8290 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1783_
timestamp 0
transform 1 0 10530 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1784_
timestamp 0
transform -1 0 10010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1785_
timestamp 0
transform -1 0 9770 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1786_
timestamp 0
transform 1 0 10190 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1787_
timestamp 0
transform -1 0 9130 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1788_
timestamp 0
transform -1 0 8550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1789_
timestamp 0
transform 1 0 9990 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1790_
timestamp 0
transform -1 0 10050 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1791_
timestamp 0
transform -1 0 10130 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1792_
timestamp 0
transform -1 0 9670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1793_
timestamp 0
transform -1 0 9410 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1794_
timestamp 0
transform 1 0 9130 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1795_
timestamp 0
transform -1 0 8330 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1796_
timestamp 0
transform -1 0 8270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1797_
timestamp 0
transform 1 0 7110 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1798_
timestamp 0
transform 1 0 7370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1799_
timestamp 0
transform -1 0 9390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1800_
timestamp 0
transform 1 0 11270 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1801_
timestamp 0
transform 1 0 9290 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1802_
timestamp 0
transform -1 0 8950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1803_
timestamp 0
transform 1 0 10550 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1804_
timestamp 0
transform -1 0 8570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1805_
timestamp 0
transform -1 0 8670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1806_
timestamp 0
transform 1 0 7610 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1807_
timestamp 0
transform -1 0 8070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1808_
timestamp 0
transform -1 0 8390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1809_
timestamp 0
transform 1 0 8610 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1810_
timestamp 0
transform 1 0 8010 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1811_
timestamp 0
transform -1 0 7750 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1812_
timestamp 0
transform -1 0 8390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1813_
timestamp 0
transform -1 0 8110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1814_
timestamp 0
transform -1 0 7850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1815_
timestamp 0
transform 1 0 7870 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1816_
timestamp 0
transform -1 0 3870 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1817_
timestamp 0
transform 1 0 1350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1818_
timestamp 0
transform -1 0 6170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1819_
timestamp 0
transform -1 0 930 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1820_
timestamp 0
transform 1 0 370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1821_
timestamp 0
transform 1 0 890 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1822_
timestamp 0
transform -1 0 350 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1823_
timestamp 0
transform 1 0 1710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1824_
timestamp 0
transform 1 0 1290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1825_
timestamp 0
transform -1 0 1130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1826_
timestamp 0
transform -1 0 390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1827_
timestamp 0
transform 1 0 890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1828_
timestamp 0
transform -1 0 1490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1829_
timestamp 0
transform -1 0 630 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1830_
timestamp 0
transform -1 0 1430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1831_
timestamp 0
transform 1 0 2010 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1832_
timestamp 0
transform -1 0 8010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1833_
timestamp 0
transform 1 0 9650 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1834_
timestamp 0
transform 1 0 9230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1835_
timestamp 0
transform -1 0 7750 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1836_
timestamp 0
transform -1 0 6410 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1837_
timestamp 0
transform -1 0 7750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1838_
timestamp 0
transform -1 0 7190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1839_
timestamp 0
transform -1 0 6170 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1840_
timestamp 0
transform 1 0 8550 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1841_
timestamp 0
transform -1 0 8170 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1842_
timestamp 0
transform -1 0 6930 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1843_
timestamp 0
transform -1 0 6650 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1844_
timestamp 0
transform 1 0 9070 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1845_
timestamp 0
transform 1 0 9610 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1846_
timestamp 0
transform -1 0 9210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1847_
timestamp 0
transform -1 0 8370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1848_
timestamp 0
transform 1 0 11210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1849_
timestamp 0
transform -1 0 11530 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1850_
timestamp 0
transform -1 0 10990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1851_
timestamp 0
transform 1 0 10350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1852_
timestamp 0
transform -1 0 10410 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1853_
timestamp 0
transform -1 0 10430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1854_
timestamp 0
transform -1 0 7410 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1855_
timestamp 0
transform 1 0 7390 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1856_
timestamp 0
transform 1 0 7670 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1857_
timestamp 0
transform -1 0 8810 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__1858_
timestamp 0
transform -1 0 9350 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1859_
timestamp 0
transform -1 0 8810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1860_
timestamp 0
transform 1 0 9070 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1861_
timestamp 0
transform 1 0 6810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1862_
timestamp 0
transform -1 0 8310 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__1863_
timestamp 0
transform 1 0 7670 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1864_
timestamp 0
transform -1 0 6310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1865_
timestamp 0
transform -1 0 7750 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__1866_
timestamp 0
transform -1 0 7210 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1867_
timestamp 0
transform -1 0 7990 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1868_
timestamp 0
transform 1 0 7710 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1869_
timestamp 0
transform -1 0 6010 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__1870_
timestamp 0
transform 1 0 9350 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1871_
timestamp 0
transform 1 0 8830 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1872_
timestamp 0
transform -1 0 8570 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1873_
timestamp 0
transform -1 0 7770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1874_
timestamp 0
transform -1 0 7490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1875_
timestamp 0
transform -1 0 8290 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1876_
timestamp 0
transform -1 0 6930 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1877_
timestamp 0
transform -1 0 5770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__1878_
timestamp 0
transform 1 0 6650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1879_
timestamp 0
transform -1 0 7450 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1880_
timestamp 0
transform 1 0 5970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__1881_
timestamp 0
transform 1 0 5970 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__1882_
timestamp 0
transform -1 0 4930 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__1883_
timestamp 0
transform -1 0 7830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1884_
timestamp 0
transform -1 0 8070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1885_
timestamp 0
transform -1 0 8630 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1886_
timestamp 0
transform 1 0 8470 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1887_
timestamp 0
transform -1 0 8450 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1888_
timestamp 0
transform 1 0 11590 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1889_
timestamp 0
transform -1 0 8450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1890_
timestamp 0
transform 1 0 9710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1891_
timestamp 0
transform 1 0 8870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1892_
timestamp 0
transform -1 0 8590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1893_
timestamp 0
transform 1 0 12110 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1894_
timestamp 0
transform 1 0 12090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1895_
timestamp 0
transform 1 0 12110 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1896_
timestamp 0
transform -1 0 10730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1897_
timestamp 0
transform -1 0 9130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1898_
timestamp 0
transform 1 0 9010 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1899_
timestamp 0
transform 1 0 7450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1900_
timestamp 0
transform 1 0 9650 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1901_
timestamp 0
transform 1 0 7990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1902_
timestamp 0
transform -1 0 8210 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1903_
timestamp 0
transform 1 0 7930 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1904_
timestamp 0
transform 1 0 11850 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1905_
timestamp 0
transform 1 0 11610 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1906_
timestamp 0
transform -1 0 6490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1907_
timestamp 0
transform -1 0 7030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1908_
timestamp 0
transform -1 0 6950 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1909_
timestamp 0
transform -1 0 6710 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1910_
timestamp 0
transform -1 0 6210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1911_
timestamp 0
transform 1 0 6790 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1912_
timestamp 0
transform 1 0 6250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1913_
timestamp 0
transform 1 0 6190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1914_
timestamp 0
transform 1 0 5690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1915_
timestamp 0
transform 1 0 5210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1916_
timestamp 0
transform 1 0 5210 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__1917_
timestamp 0
transform -1 0 3710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__1918_
timestamp 0
transform 1 0 3590 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__1919_
timestamp 0
transform -1 0 3870 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__1920_
timestamp 0
transform -1 0 3590 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__1921_
timestamp 0
transform -1 0 1710 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__1922_
timestamp 0
transform 1 0 7510 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1923_
timestamp 0
transform 1 0 7770 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1924_
timestamp 0
transform -1 0 6370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1925_
timestamp 0
transform -1 0 4610 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1926_
timestamp 0
transform -1 0 3970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1927_
timestamp 0
transform 1 0 2010 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__1928_
timestamp 0
transform -1 0 3170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__1929_
timestamp 0
transform 1 0 4550 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__1930_
timestamp 0
transform 1 0 3110 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__1931_
timestamp 0
transform -1 0 2890 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__1932_
timestamp 0
transform -1 0 1490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1933_
timestamp 0
transform -1 0 8450 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1934_
timestamp 0
transform 1 0 3850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1935_
timestamp 0
transform -1 0 3870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1936_
timestamp 0
transform -1 0 2550 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1937_
timestamp 0
transform -1 0 1210 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1938_
timestamp 0
transform -1 0 3570 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1939_
timestamp 0
transform -1 0 4130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1940_
timestamp 0
transform -1 0 3350 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1941_
timestamp 0
transform -1 0 3290 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1942_
timestamp 0
transform -1 0 1790 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__1943_
timestamp 0
transform -1 0 3590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1944_
timestamp 0
transform -1 0 3690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1945_
timestamp 0
transform -1 0 2950 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1946_
timestamp 0
transform -1 0 1510 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__1947_
timestamp 0
transform -1 0 4930 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__1948_
timestamp 0
transform 1 0 5130 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__1949_
timestamp 0
transform 1 0 5190 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__1950_
timestamp 0
transform -1 0 4930 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__1951_
timestamp 0
transform -1 0 1970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1952_
timestamp 0
transform 1 0 4090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1953_
timestamp 0
transform 1 0 4030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1954_
timestamp 0
transform 1 0 4170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1955_
timestamp 0
transform -1 0 1690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1956_
timestamp 0
transform -1 0 4310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__1957_
timestamp 0
transform 1 0 4890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__1958_
timestamp 0
transform -1 0 5170 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__1959_
timestamp 0
transform -1 0 4150 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__1960_
timestamp 0
transform -1 0 2310 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1961_
timestamp 0
transform 1 0 4130 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1962_
timestamp 0
transform 1 0 3890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1963_
timestamp 0
transform 1 0 3670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1964_
timestamp 0
transform 1 0 2010 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1965_
timestamp 0
transform 1 0 6390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__1966_
timestamp 0
transform 1 0 6330 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1967_
timestamp 0
transform 1 0 7170 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1968_
timestamp 0
transform 1 0 6630 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1969_
timestamp 0
transform -1 0 3290 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__1970_
timestamp 0
transform 1 0 2830 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1971_
timestamp 0
transform -1 0 4710 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1972_
timestamp 0
transform 1 0 3570 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1973_
timestamp 0
transform -1 0 3590 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1974_
timestamp 0
transform -1 0 3090 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__1975_
timestamp 0
transform 1 0 2990 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__1976_
timestamp 0
transform -1 0 3090 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__1977_
timestamp 0
transform 1 0 4370 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__1978_
timestamp 0
transform 1 0 3070 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__1979_
timestamp 0
transform -1 0 2810 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__1980_
timestamp 0
transform -1 0 2330 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1981_
timestamp 0
transform 1 0 5950 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1982_
timestamp 0
transform 1 0 6070 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1983_
timestamp 0
transform 1 0 6270 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1984_
timestamp 0
transform 1 0 5270 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1985_
timestamp 0
transform -1 0 4770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1986_
timestamp 0
transform 1 0 2550 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__1987_
timestamp 0
transform -1 0 7270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1988_
timestamp 0
transform 1 0 7570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1989_
timestamp 0
transform 1 0 7630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1990_
timestamp 0
transform -1 0 7430 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1991_
timestamp 0
transform -1 0 7710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1992_
timestamp 0
transform 1 0 10450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1993_
timestamp 0
transform 1 0 9570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__1994_
timestamp 0
transform -1 0 6250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__1995_
timestamp 0
transform 1 0 6630 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1996_
timestamp 0
transform -1 0 6770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1997_
timestamp 0
transform 1 0 6470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1998_
timestamp 0
transform 1 0 6470 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__1999_
timestamp 0
transform 1 0 7530 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2000_
timestamp 0
transform 1 0 6450 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2001_
timestamp 0
transform 1 0 6690 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2002_
timestamp 0
transform 1 0 6650 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2003_
timestamp 0
transform 1 0 9530 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2004_
timestamp 0
transform 1 0 7470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2005_
timestamp 0
transform -1 0 7270 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2006_
timestamp 0
transform 1 0 6750 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2007_
timestamp 0
transform 1 0 6590 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2008_
timestamp 0
transform -1 0 6230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2009_
timestamp 0
transform 1 0 6830 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2010_
timestamp 0
transform -1 0 7050 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2011_
timestamp 0
transform 1 0 7290 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2012_
timestamp 0
transform -1 0 9430 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2013_
timestamp 0
transform 1 0 10570 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2014_
timestamp 0
transform -1 0 10830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2015_
timestamp 0
transform -1 0 6270 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2016_
timestamp 0
transform -1 0 7310 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2017_
timestamp 0
transform -1 0 7090 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2018_
timestamp 0
transform 1 0 7330 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2019_
timestamp 0
transform 1 0 9410 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2020_
timestamp 0
transform -1 0 10310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2021_
timestamp 0
transform -1 0 7350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2022_
timestamp 0
transform 1 0 7590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2023_
timestamp 0
transform -1 0 7890 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2024_
timestamp 0
transform 1 0 6110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2025_
timestamp 0
transform -1 0 5990 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2026_
timestamp 0
transform 1 0 9690 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2027_
timestamp 0
transform 1 0 10230 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2028_
timestamp 0
transform -1 0 10230 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2029_
timestamp 0
transform -1 0 11110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2030_
timestamp 0
transform 1 0 10730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2031_
timestamp 0
transform -1 0 11030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2032_
timestamp 0
transform 1 0 8950 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2033_
timestamp 0
transform 1 0 8410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2034_
timestamp 0
transform 1 0 8650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2035_
timestamp 0
transform 1 0 8610 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2036_
timestamp 0
transform 1 0 11570 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2037_
timestamp 0
transform 1 0 11770 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2038_
timestamp 0
transform -1 0 7610 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2039_
timestamp 0
transform -1 0 6690 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2040_
timestamp 0
transform 1 0 10950 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2041_
timestamp 0
transform 1 0 11030 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2042_
timestamp 0
transform -1 0 10110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2043_
timestamp 0
transform -1 0 10490 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2044_
timestamp 0
transform -1 0 11010 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2045_
timestamp 0
transform -1 0 11350 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2046_
timestamp 0
transform 1 0 8830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2047_
timestamp 0
transform -1 0 9390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2048_
timestamp 0
transform 1 0 9190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2049_
timestamp 0
transform 1 0 9330 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2050_
timestamp 0
transform 1 0 9090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2051_
timestamp 0
transform 1 0 8790 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2052_
timestamp 0
transform 1 0 9070 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2053_
timestamp 0
transform -1 0 9630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2054_
timestamp 0
transform 1 0 9850 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2055_
timestamp 0
transform -1 0 6490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2056_
timestamp 0
transform -1 0 6070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2057_
timestamp 0
transform 1 0 10270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2058_
timestamp 0
transform -1 0 10010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2059_
timestamp 0
transform -1 0 10150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2060_
timestamp 0
transform -1 0 9910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2061_
timestamp 0
transform 1 0 10090 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2062_
timestamp 0
transform -1 0 9170 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2063_
timestamp 0
transform 1 0 8250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2064_
timestamp 0
transform -1 0 7930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2065_
timestamp 0
transform -1 0 8750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2066_
timestamp 0
transform 1 0 8730 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2067_
timestamp 0
transform -1 0 7990 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2068_
timestamp 0
transform -1 0 8270 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2069_
timestamp 0
transform 1 0 7990 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2070_
timestamp 0
transform -1 0 8290 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2071_
timestamp 0
transform -1 0 8570 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2072_
timestamp 0
transform 1 0 8790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2073_
timestamp 0
transform 1 0 9050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2074_
timestamp 0
transform 1 0 9270 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2075_
timestamp 0
transform -1 0 9570 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2076_
timestamp 0
transform 1 0 11230 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2077_
timestamp 0
transform -1 0 11290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2078_
timestamp 0
transform -1 0 11090 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2079_
timestamp 0
transform 1 0 11230 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2080_
timestamp 0
transform -1 0 11070 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2081_
timestamp 0
transform 1 0 11070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2082_
timestamp 0
transform 1 0 10330 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2083_
timestamp 0
transform 1 0 9590 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2084_
timestamp 0
transform 1 0 11610 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2085_
timestamp 0
transform 1 0 11030 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2086_
timestamp 0
transform 1 0 11530 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2087_
timestamp 0
transform 1 0 11550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2088_
timestamp 0
transform -1 0 12110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2089_
timestamp 0
transform 1 0 11830 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2090_
timestamp 0
transform 1 0 12010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2091_
timestamp 0
transform 1 0 9910 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2092_
timestamp 0
transform 1 0 10530 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2093_
timestamp 0
transform -1 0 11090 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2094_
timestamp 0
transform 1 0 11330 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2095_
timestamp 0
transform -1 0 10990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2096_
timestamp 0
transform 1 0 11510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2097_
timestamp 0
transform -1 0 11850 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2098_
timestamp 0
transform -1 0 12030 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2099_
timestamp 0
transform -1 0 11330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2100_
timestamp 0
transform 1 0 11290 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2101_
timestamp 0
transform -1 0 11250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2102_
timestamp 0
transform -1 0 11630 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2103_
timestamp 0
transform 1 0 12110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2104_
timestamp 0
transform 1 0 12110 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2105_
timestamp 0
transform -1 0 11570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2106_
timestamp 0
transform -1 0 11550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2107_
timestamp 0
transform -1 0 12110 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2108_
timestamp 0
transform 1 0 8850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2109_
timestamp 0
transform 1 0 12110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2110_
timestamp 0
transform -1 0 12130 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2111_
timestamp 0
transform -1 0 12130 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2112_
timestamp 0
transform -1 0 12030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2113_
timestamp 0
transform 1 0 11790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2114_
timestamp 0
transform 1 0 10570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2115_
timestamp 0
transform -1 0 9310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2116_
timestamp 0
transform -1 0 10190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2117_
timestamp 0
transform -1 0 10790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2118_
timestamp 0
transform -1 0 10750 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2119_
timestamp 0
transform 1 0 10650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2120_
timestamp 0
transform 1 0 10690 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2121_
timestamp 0
transform -1 0 10430 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2122_
timestamp 0
transform 1 0 10630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2123_
timestamp 0
transform -1 0 8130 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2124_
timestamp 0
transform -1 0 7830 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2125_
timestamp 0
transform -1 0 10190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2126_
timestamp 0
transform 1 0 10590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2127_
timestamp 0
transform -1 0 7010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2128_
timestamp 0
transform -1 0 9150 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2129_
timestamp 0
transform 1 0 7270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2130_
timestamp 0
transform -1 0 10890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2131_
timestamp 0
transform -1 0 7930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2132_
timestamp 0
transform 1 0 6710 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2133_
timestamp 0
transform -1 0 7010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2134_
timestamp 0
transform -1 0 7270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2135_
timestamp 0
transform -1 0 11150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2136_
timestamp 0
transform -1 0 11310 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2137_
timestamp 0
transform 1 0 11290 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2138_
timestamp 0
transform 1 0 11370 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2139_
timestamp 0
transform -1 0 11290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2140_
timestamp 0
transform -1 0 11010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2141_
timestamp 0
transform 1 0 9930 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2142_
timestamp 0
transform 1 0 10730 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2143_
timestamp 0
transform -1 0 10470 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2144_
timestamp 0
transform -1 0 11030 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2145_
timestamp 0
transform -1 0 5030 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2146_
timestamp 0
transform 1 0 9750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2147_
timestamp 0
transform 1 0 10310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2148_
timestamp 0
transform -1 0 6250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2149_
timestamp 0
transform 1 0 10030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2150_
timestamp 0
transform 1 0 8810 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2151_
timestamp 0
transform 1 0 7430 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2152_
timestamp 0
transform 1 0 8510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2153_
timestamp 0
transform 1 0 8770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2154_
timestamp 0
transform 1 0 9050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2155_
timestamp 0
transform -1 0 10130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2156_
timestamp 0
transform -1 0 10910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2157_
timestamp 0
transform 1 0 11150 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2158_
timestamp 0
transform -1 0 11730 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2159_
timestamp 0
transform -1 0 11850 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2160_
timestamp 0
transform -1 0 11390 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2161_
timestamp 0
transform 1 0 8130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2162_
timestamp 0
transform 1 0 8890 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2163_
timestamp 0
transform -1 0 9990 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2164_
timestamp 0
transform 1 0 9750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2165_
timestamp 0
transform 1 0 10990 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2166_
timestamp 0
transform 1 0 10810 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2167_
timestamp 0
transform 1 0 9190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2168_
timestamp 0
transform 1 0 10010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2169_
timestamp 0
transform -1 0 8750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2170_
timestamp 0
transform -1 0 9170 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2171_
timestamp 0
transform 1 0 10310 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2172_
timestamp 0
transform 1 0 9730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2173_
timestamp 0
transform 1 0 9850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2174_
timestamp 0
transform -1 0 9490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2175_
timestamp 0
transform 1 0 9570 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2176_
timestamp 0
transform -1 0 9690 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2177_
timestamp 0
transform -1 0 9390 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2178_
timestamp 0
transform -1 0 10990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2179_
timestamp 0
transform 1 0 9470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2180_
timestamp 0
transform 1 0 11830 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2181_
timestamp 0
transform 1 0 11810 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2182_
timestamp 0
transform 1 0 11890 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2183_
timestamp 0
transform -1 0 11270 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2184_
timestamp 0
transform 1 0 11010 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2185_
timestamp 0
transform -1 0 10250 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2186_
timestamp 0
transform 1 0 10190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2187_
timestamp 0
transform -1 0 10590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2188_
timestamp 0
transform 1 0 11550 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2189_
timestamp 0
transform 1 0 9930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2190_
timestamp 0
transform 1 0 10490 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2191_
timestamp 0
transform 1 0 11110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2192_
timestamp 0
transform 1 0 11050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2193_
timestamp 0
transform -1 0 10990 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2194_
timestamp 0
transform -1 0 10550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2195_
timestamp 0
transform -1 0 9430 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2196_
timestamp 0
transform -1 0 11070 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2197_
timestamp 0
transform 1 0 11330 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2198_
timestamp 0
transform -1 0 9870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2199_
timestamp 0
transform -1 0 9930 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2200_
timestamp 0
transform -1 0 5790 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2201_
timestamp 0
transform 1 0 6310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2202_
timestamp 0
transform 1 0 6050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2203_
timestamp 0
transform 1 0 6050 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2204_
timestamp 0
transform 1 0 6790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2205_
timestamp 0
transform 1 0 7090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2206_
timestamp 0
transform 1 0 9430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2207_
timestamp 0
transform -1 0 9930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2208_
timestamp 0
transform -1 0 9350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2209_
timestamp 0
transform 1 0 10390 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2210_
timestamp 0
transform 1 0 10390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2211_
timestamp 0
transform 1 0 11230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2212_
timestamp 0
transform -1 0 11590 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2213_
timestamp 0
transform -1 0 11630 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2214_
timestamp 0
transform 1 0 11590 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2215_
timestamp 0
transform 1 0 11690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2216_
timestamp 0
transform 1 0 12070 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2217_
timestamp 0
transform 1 0 11350 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2218_
timestamp 0
transform 1 0 9630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2219_
timestamp 0
transform -1 0 9870 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2220_
timestamp 0
transform -1 0 9910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2221_
timestamp 0
transform -1 0 11850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2222_
timestamp 0
transform 1 0 11790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2223_
timestamp 0
transform -1 0 11830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2224_
timestamp 0
transform 1 0 11810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2225_
timestamp 0
transform 1 0 10910 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2226_
timestamp 0
transform 1 0 11870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2227_
timestamp 0
transform 1 0 11590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2228_
timestamp 0
transform -1 0 11450 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2229_
timestamp 0
transform -1 0 10530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2230_
timestamp 0
transform -1 0 10250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2231_
timestamp 0
transform -1 0 8450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2232_
timestamp 0
transform 1 0 8690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2233_
timestamp 0
transform 1 0 9470 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2234_
timestamp 0
transform -1 0 9730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2235_
timestamp 0
transform -1 0 9850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2236_
timestamp 0
transform 1 0 7150 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2237_
timestamp 0
transform -1 0 6630 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2238_
timestamp 0
transform -1 0 6910 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2239_
timestamp 0
transform -1 0 8930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2240_
timestamp 0
transform -1 0 8650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2241_
timestamp 0
transform -1 0 8290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2242_
timestamp 0
transform -1 0 7470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2243_
timestamp 0
transform 1 0 7730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2244_
timestamp 0
transform 1 0 8010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2245_
timestamp 0
transform -1 0 7710 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2246_
timestamp 0
transform 1 0 9090 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2247_
timestamp 0
transform -1 0 12090 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2248_
timestamp 0
transform 1 0 11290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2249_
timestamp 0
transform -1 0 9450 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2250_
timestamp 0
transform 1 0 10970 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2251_
timestamp 0
transform 1 0 10530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2252_
timestamp 0
transform 1 0 11270 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2253_
timestamp 0
transform -1 0 11870 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2254_
timestamp 0
transform 1 0 12110 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2255_
timestamp 0
transform -1 0 10470 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2256_
timestamp 0
transform -1 0 10750 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2257_
timestamp 0
transform 1 0 10990 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2258_
timestamp 0
transform 1 0 12150 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2259_
timestamp 0
transform -1 0 11830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2260_
timestamp 0
transform 1 0 10010 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2261_
timestamp 0
transform 1 0 10270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2262_
timestamp 0
transform -1 0 10790 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2263_
timestamp 0
transform 1 0 11270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2264_
timestamp 0
transform 1 0 12090 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2265_
timestamp 0
transform -1 0 11350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2266_
timestamp 0
transform -1 0 10710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2267_
timestamp 0
transform 1 0 11930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2268_
timestamp 0
transform 1 0 12090 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2269_
timestamp 0
transform -1 0 11870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2270_
timestamp 0
transform 1 0 11290 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2271_
timestamp 0
transform -1 0 11590 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2272_
timestamp 0
transform 1 0 11850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2273_
timestamp 0
transform -1 0 12110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2274_
timestamp 0
transform 1 0 10030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2275_
timestamp 0
transform -1 0 8190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2276_
timestamp 0
transform 1 0 8850 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2277_
timestamp 0
transform 1 0 9130 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2278_
timestamp 0
transform -1 0 9210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2279_
timestamp 0
transform 1 0 9010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2280_
timestamp 0
transform 1 0 10170 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2281_
timestamp 0
transform 1 0 12050 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2282_
timestamp 0
transform 1 0 12110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2283_
timestamp 0
transform -1 0 10990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2284_
timestamp 0
transform 1 0 12070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2285_
timestamp 0
transform 1 0 12070 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2286_
timestamp 0
transform -1 0 11850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2287_
timestamp 0
transform 1 0 11790 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2288_
timestamp 0
transform -1 0 10950 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2289_
timestamp 0
transform -1 0 10730 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2290_
timestamp 0
transform -1 0 10910 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2291_
timestamp 0
transform 1 0 11270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2292_
timestamp 0
transform 1 0 10410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2293_
timestamp 0
transform 1 0 10690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2294_
timestamp 0
transform 1 0 11010 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2295_
timestamp 0
transform 1 0 10890 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2296_
timestamp 0
transform 1 0 11150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2297_
timestamp 0
transform 1 0 11810 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2298_
timestamp 0
transform -1 0 11910 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2299_
timestamp 0
transform -1 0 10470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2300_
timestamp 0
transform 1 0 10170 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2301_
timestamp 0
transform 1 0 11790 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2302_
timestamp 0
transform 1 0 11730 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2303_
timestamp 0
transform -1 0 11710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2304_
timestamp 0
transform 1 0 11850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2305_
timestamp 0
transform 1 0 10730 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2306_
timestamp 0
transform -1 0 11590 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2307_
timestamp 0
transform 1 0 11290 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2308_
timestamp 0
transform 1 0 12070 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2309_
timestamp 0
transform -1 0 11630 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2310_
timestamp 0
transform -1 0 11570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2311_
timestamp 0
transform 1 0 11550 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2312_
timestamp 0
transform 1 0 11610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2313_
timestamp 0
transform 1 0 11890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2314_
timestamp 0
transform -1 0 11210 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2315_
timestamp 0
transform 1 0 12070 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2316_
timestamp 0
transform 1 0 11470 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2317_
timestamp 0
transform -1 0 11970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2318_
timestamp 0
transform 1 0 11510 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2319_
timestamp 0
transform 1 0 11150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2320_
timestamp 0
transform 1 0 11570 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2321_
timestamp 0
transform 1 0 11430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2322_
timestamp 0
transform -1 0 11290 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2323_
timestamp 0
transform -1 0 11530 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2324_
timestamp 0
transform 1 0 11770 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2325_
timestamp 0
transform -1 0 12150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2326_
timestamp 0
transform 1 0 12070 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2327_
timestamp 0
transform 1 0 11430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2328_
timestamp 0
transform 1 0 11010 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2329_
timestamp 0
transform 1 0 8530 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2330_
timestamp 0
transform -1 0 10210 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2331_
timestamp 0
transform -1 0 9650 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2332_
timestamp 0
transform -1 0 11870 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2333_
timestamp 0
transform -1 0 10750 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2334_
timestamp 0
transform 1 0 10470 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2335_
timestamp 0
transform 1 0 10450 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2336_
timestamp 0
transform 1 0 10630 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2337_
timestamp 0
transform -1 0 10750 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2338_
timestamp 0
transform -1 0 10670 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2339_
timestamp 0
transform -1 0 9590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2340_
timestamp 0
transform -1 0 9870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2341_
timestamp 0
transform 1 0 9570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2342_
timestamp 0
transform -1 0 10450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2343_
timestamp 0
transform -1 0 10390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2344_
timestamp 0
transform -1 0 10630 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2345_
timestamp 0
transform 1 0 11750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2346_
timestamp 0
transform 1 0 11490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2347_
timestamp 0
transform -1 0 8830 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2348_
timestamp 0
transform -1 0 9930 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2349_
timestamp 0
transform -1 0 11590 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2350_
timestamp 0
transform -1 0 11310 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2351_
timestamp 0
transform -1 0 10370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2352_
timestamp 0
transform -1 0 10130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2353_
timestamp 0
transform -1 0 9430 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2354_
timestamp 0
transform 1 0 7830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2355_
timestamp 0
transform -1 0 6910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2356_
timestamp 0
transform -1 0 6850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2357_
timestamp 0
transform -1 0 7510 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2358_
timestamp 0
transform -1 0 7090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2359_
timestamp 0
transform 1 0 7310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2360_
timestamp 0
transform -1 0 7990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2361_
timestamp 0
transform -1 0 7050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2362_
timestamp 0
transform 1 0 8770 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2363_
timestamp 0
transform -1 0 7450 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2364_
timestamp 0
transform 1 0 7190 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2365_
timestamp 0
transform 1 0 6910 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2366_
timestamp 0
transform 1 0 6390 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2367_
timestamp 0
transform -1 0 7230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2368_
timestamp 0
transform 1 0 6630 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2369_
timestamp 0
transform 1 0 7010 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2370_
timestamp 0
transform -1 0 7270 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2371_
timestamp 0
transform 1 0 7210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2372_
timestamp 0
transform -1 0 6790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2373_
timestamp 0
transform 1 0 6730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2374_
timestamp 0
transform 1 0 8230 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2375_
timestamp 0
transform 1 0 8290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2376_
timestamp 0
transform -1 0 6730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2377_
timestamp 0
transform 1 0 5430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2378_
timestamp 0
transform -1 0 3750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2379_
timestamp 0
transform -1 0 8010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2380_
timestamp 0
transform -1 0 5650 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2381_
timestamp 0
transform -1 0 5930 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2382_
timestamp 0
transform -1 0 5790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2383_
timestamp 0
transform 1 0 4710 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2384_
timestamp 0
transform 1 0 4630 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2385_
timestamp 0
transform 1 0 4870 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2386_
timestamp 0
transform 1 0 5150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2387_
timestamp 0
transform 1 0 1670 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2388_
timestamp 0
transform 1 0 1610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2389_
timestamp 0
transform 1 0 5190 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2390_
timestamp 0
transform 1 0 2470 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2391_
timestamp 0
transform -1 0 2270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2392_
timestamp 0
transform -1 0 1990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2393_
timestamp 0
transform -1 0 2550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2394_
timestamp 0
transform -1 0 2970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2395_
timestamp 0
transform 1 0 4370 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2396_
timestamp 0
transform 1 0 3010 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2397_
timestamp 0
transform -1 0 3090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2398_
timestamp 0
transform -1 0 2810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2399_
timestamp 0
transform 1 0 1910 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2400_
timestamp 0
transform -1 0 1350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2401_
timestamp 0
transform -1 0 2830 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2402_
timestamp 0
transform 1 0 2570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2403_
timestamp 0
transform -1 0 2210 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2404_
timestamp 0
transform -1 0 1650 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2405_
timestamp 0
transform -1 0 1510 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2406_
timestamp 0
transform 1 0 5890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2407_
timestamp 0
transform -1 0 4250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2408_
timestamp 0
transform -1 0 5610 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2409_
timestamp 0
transform -1 0 6430 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2410_
timestamp 0
transform -1 0 4210 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2411_
timestamp 0
transform -1 0 3970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2412_
timestamp 0
transform -1 0 1230 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2413_
timestamp 0
transform -1 0 4510 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2414_
timestamp 0
transform 1 0 3030 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2415_
timestamp 0
transform -1 0 2770 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2416_
timestamp 0
transform 1 0 1730 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2417_
timestamp 0
transform -1 0 2230 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2418_
timestamp 0
transform -1 0 2110 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2419_
timestamp 0
transform -1 0 3430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2420_
timestamp 0
transform 1 0 2850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2421_
timestamp 0
transform -1 0 2770 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2422_
timestamp 0
transform -1 0 1950 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2423_
timestamp 0
transform -1 0 3650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2424_
timestamp 0
transform -1 0 3490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2425_
timestamp 0
transform -1 0 3370 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2426_
timestamp 0
transform 1 0 3130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2427_
timestamp 0
transform 1 0 3290 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2428_
timestamp 0
transform -1 0 3370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2429_
timestamp 0
transform -1 0 5090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2430_
timestamp 0
transform -1 0 7790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2431_
timestamp 0
transform -1 0 5350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2432_
timestamp 0
transform -1 0 9470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2433_
timestamp 0
transform 1 0 11570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2434_
timestamp 0
transform 1 0 10750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2435_
timestamp 0
transform -1 0 7230 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2436_
timestamp 0
transform -1 0 6910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2437_
timestamp 0
transform -1 0 9590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2438_
timestamp 0
transform -1 0 9330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2439_
timestamp 0
transform -1 0 6110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2440_
timestamp 0
transform 1 0 7730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2441_
timestamp 0
transform -1 0 7570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2442_
timestamp 0
transform 1 0 10270 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2443_
timestamp 0
transform -1 0 7170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2444_
timestamp 0
transform -1 0 7170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2445_
timestamp 0
transform 1 0 5270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2446_
timestamp 0
transform 1 0 6390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2447_
timestamp 0
transform -1 0 4770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2448_
timestamp 0
transform -1 0 6370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2449_
timestamp 0
transform -1 0 6990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2450_
timestamp 0
transform 1 0 4130 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2451_
timestamp 0
transform -1 0 4010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2452_
timestamp 0
transform 1 0 4650 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2453_
timestamp 0
transform 1 0 8510 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2454_
timestamp 0
transform 1 0 4390 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2455_
timestamp 0
transform 1 0 4390 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2456_
timestamp 0
transform -1 0 4250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2457_
timestamp 0
transform -1 0 4510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2458_
timestamp 0
transform -1 0 4870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2459_
timestamp 0
transform 1 0 5010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2460_
timestamp 0
transform 1 0 4890 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2461_
timestamp 0
transform 1 0 5170 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2462_
timestamp 0
transform 1 0 5310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2463_
timestamp 0
transform 1 0 6250 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2464_
timestamp 0
transform -1 0 3190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2465_
timestamp 0
transform -1 0 2910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2466_
timestamp 0
transform -1 0 2910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2467_
timestamp 0
transform 1 0 2050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2468_
timestamp 0
transform -1 0 1610 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2469_
timestamp 0
transform 1 0 570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2470_
timestamp 0
transform -1 0 2670 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2471_
timestamp 0
transform -1 0 2690 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2472_
timestamp 0
transform -1 0 2390 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2473_
timestamp 0
transform 1 0 1890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2474_
timestamp 0
transform -1 0 1410 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2475_
timestamp 0
transform -1 0 350 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2476_
timestamp 0
transform -1 0 3770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2477_
timestamp 0
transform -1 0 5010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2478_
timestamp 0
transform 1 0 3870 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2479_
timestamp 0
transform -1 0 3510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2480_
timestamp 0
transform 1 0 1750 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2481_
timestamp 0
transform -1 0 3310 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2482_
timestamp 0
transform 1 0 3590 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2483_
timestamp 0
transform 1 0 3010 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2484_
timestamp 0
transform 1 0 2730 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2485_
timestamp 0
transform -1 0 350 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2486_
timestamp 0
transform -1 0 2630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2487_
timestamp 0
transform 1 0 2350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2488_
timestamp 0
transform -1 0 2350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2489_
timestamp 0
transform -1 0 1790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2490_
timestamp 0
transform -1 0 1350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2491_
timestamp 0
transform -1 0 350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2492_
timestamp 0
transform 1 0 4570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2493_
timestamp 0
transform 1 0 3570 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2494_
timestamp 0
transform 1 0 6150 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2495_
timestamp 0
transform 1 0 3810 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2496_
timestamp 0
transform 1 0 4110 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2497_
timestamp 0
transform -1 0 4030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2498_
timestamp 0
transform 1 0 3490 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2499_
timestamp 0
transform 1 0 3750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2500_
timestamp 0
transform -1 0 350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2501_
timestamp 0
transform -1 0 3350 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2502_
timestamp 0
transform -1 0 2990 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2503_
timestamp 0
transform -1 0 3470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__2504_
timestamp 0
transform -1 0 3230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__2505_
timestamp 0
transform 1 0 2670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2506_
timestamp 0
transform -1 0 2490 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__2507_
timestamp 0
transform 1 0 610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2508_
timestamp 0
transform 1 0 3110 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2509_
timestamp 0
transform 1 0 2650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2510_
timestamp 0
transform -1 0 3210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2511_
timestamp 0
transform 1 0 3290 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__2512_
timestamp 0
transform 1 0 3130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2513_
timestamp 0
transform -1 0 2390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2514_
timestamp 0
transform 1 0 2090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2515_
timestamp 0
transform -1 0 2110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2516_
timestamp 0
transform -1 0 350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__2517_
timestamp 0
transform -1 0 2190 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2518_
timestamp 0
transform 1 0 5290 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2519_
timestamp 0
transform -1 0 5830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2520_
timestamp 0
transform -1 0 5930 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2521_
timestamp 0
transform 1 0 5630 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2522_
timestamp 0
transform -1 0 5630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2523_
timestamp 0
transform -1 0 5550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2524_
timestamp 0
transform -1 0 5490 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2525_
timestamp 0
transform -1 0 2710 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2526_
timestamp 0
transform 1 0 6110 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2527_
timestamp 0
transform 1 0 6510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2528_
timestamp 0
transform 1 0 6490 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2529_
timestamp 0
transform 1 0 6090 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2530_
timestamp 0
transform 1 0 5550 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2531_
timestamp 0
transform 1 0 2910 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2532_
timestamp 0
transform 1 0 4190 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2533_
timestamp 0
transform 1 0 5130 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2534_
timestamp 0
transform 1 0 4850 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2535_
timestamp 0
transform -1 0 4590 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2536_
timestamp 0
transform 1 0 3430 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2537_
timestamp 0
transform 1 0 2070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2538_
timestamp 0
transform 1 0 4470 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2539_
timestamp 0
transform 1 0 3850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2540_
timestamp 0
transform 1 0 4190 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2541_
timestamp 0
transform -1 0 4170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2542_
timestamp 0
transform -1 0 3690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2543_
timestamp 0
transform 1 0 3450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2544_
timestamp 0
transform 1 0 4170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2545_
timestamp 0
transform 1 0 4430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2546_
timestamp 0
transform 1 0 4790 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2547_
timestamp 0
transform -1 0 4730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2548_
timestamp 0
transform -1 0 4450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2549_
timestamp 0
transform 1 0 4670 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2550_
timestamp 0
transform 1 0 4670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2551_
timestamp 0
transform 1 0 5190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2552_
timestamp 0
transform 1 0 5430 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2553_
timestamp 0
transform 1 0 2330 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2554_
timestamp 0
transform 1 0 4470 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2555_
timestamp 0
transform -1 0 4650 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2556_
timestamp 0
transform -1 0 4890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2557_
timestamp 0
transform 1 0 4590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2558_
timestamp 0
transform 1 0 4670 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2559_
timestamp 0
transform 1 0 4390 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2560_
timestamp 0
transform 1 0 3890 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2561_
timestamp 0
transform 1 0 3590 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2562_
timestamp 0
transform 1 0 2210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2563_
timestamp 0
transform -1 0 4430 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2564_
timestamp 0
transform 1 0 4350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2565_
timestamp 0
transform -1 0 3830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2566_
timestamp 0
transform 1 0 2430 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2567_
timestamp 0
transform 1 0 3910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2568_
timestamp 0
transform -1 0 5710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2569_
timestamp 0
transform -1 0 5850 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2570_
timestamp 0
transform 1 0 5930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2571_
timestamp 0
transform 1 0 5930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2572_
timestamp 0
transform 1 0 5790 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2573_
timestamp 0
transform 1 0 5710 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2574_
timestamp 0
transform 1 0 5690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2575_
timestamp 0
transform -1 0 4730 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2576_
timestamp 0
transform -1 0 4210 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2577_
timestamp 0
transform -1 0 4470 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2578_
timestamp 0
transform 1 0 6970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2579_
timestamp 0
transform 1 0 6990 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2580_
timestamp 0
transform 1 0 7990 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2581_
timestamp 0
transform -1 0 8850 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2582_
timestamp 0
transform 1 0 6890 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2583_
timestamp 0
transform -1 0 6890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2584_
timestamp 0
transform 1 0 7310 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2585_
timestamp 0
transform 1 0 7350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2586_
timestamp 0
transform -1 0 8430 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2587_
timestamp 0
transform -1 0 6770 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2588_
timestamp 0
transform -1 0 5810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2589_
timestamp 0
transform 1 0 7430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2590_
timestamp 0
transform -1 0 6210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2591_
timestamp 0
transform 1 0 6450 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2592_
timestamp 0
transform -1 0 4430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2593_
timestamp 0
transform 1 0 4950 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2594_
timestamp 0
transform -1 0 8530 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2595_
timestamp 0
transform -1 0 5250 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2596_
timestamp 0
transform 1 0 5250 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2597_
timestamp 0
transform 1 0 5430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2598_
timestamp 0
transform -1 0 5170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2599_
timestamp 0
transform -1 0 4970 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2600_
timestamp 0
transform -1 0 4970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2601_
timestamp 0
transform -1 0 5230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2602_
timestamp 0
transform -1 0 8170 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2603_
timestamp 0
transform -1 0 6610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2604_
timestamp 0
transform -1 0 6370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2605_
timestamp 0
transform 1 0 6050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2606_
timestamp 0
transform -1 0 5550 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2607_
timestamp 0
transform 1 0 5710 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2608_
timestamp 0
transform 1 0 5530 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2609_
timestamp 0
transform -1 0 5510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2610_
timestamp 0
transform 1 0 4890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2611_
timestamp 0
transform -1 0 5150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2612_
timestamp 0
transform -1 0 5410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2613_
timestamp 0
transform -1 0 1230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2614_
timestamp 0
transform 1 0 2210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2615_
timestamp 0
transform -1 0 2490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2616_
timestamp 0
transform -1 0 2470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2617_
timestamp 0
transform 1 0 1450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2618_
timestamp 0
transform 1 0 870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2619_
timestamp 0
transform -1 0 370 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2620_
timestamp 0
transform -1 0 610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2621_
timestamp 0
transform 1 0 930 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2622_
timestamp 0
transform 1 0 370 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2623_
timestamp 0
transform 1 0 2750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2624_
timestamp 0
transform 1 0 1950 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2625_
timestamp 0
transform -1 0 2210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2626_
timestamp 0
transform -1 0 1930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2627_
timestamp 0
transform 1 0 70 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2628_
timestamp 0
transform 1 0 70 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2629_
timestamp 0
transform -1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2630_
timestamp 0
transform 1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2631_
timestamp 0
transform 1 0 5010 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2632_
timestamp 0
transform 1 0 2250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2633_
timestamp 0
transform -1 0 2550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2634_
timestamp 0
transform -1 0 90 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2635_
timestamp 0
transform 1 0 70 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2636_
timestamp 0
transform 1 0 610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2637_
timestamp 0
transform 1 0 950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2638_
timestamp 0
transform 1 0 370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2639_
timestamp 0
transform -1 0 690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2640_
timestamp 0
transform -1 0 90 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2641_
timestamp 0
transform -1 0 90 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2642_
timestamp 0
transform 1 0 1330 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2643_
timestamp 0
transform -1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2644_
timestamp 0
transform 1 0 2270 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2645_
timestamp 0
transform -1 0 2010 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2646_
timestamp 0
transform -1 0 1210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2647_
timestamp 0
transform 1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2648_
timestamp 0
transform 1 0 570 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__2649_
timestamp 0
transform 1 0 70 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2650_
timestamp 0
transform -1 0 3670 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2651_
timestamp 0
transform -1 0 3390 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2652_
timestamp 0
transform 1 0 610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2653_
timestamp 0
transform 1 0 330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2654_
timestamp 0
transform 1 0 1210 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2655_
timestamp 0
transform 1 0 650 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2656_
timestamp 0
transform -1 0 930 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2657_
timestamp 0
transform 1 0 70 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2658_
timestamp 0
transform 1 0 70 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2659_
timestamp 0
transform -1 0 370 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2660_
timestamp 0
transform 1 0 310 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2661_
timestamp 0
transform -1 0 2630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__2662_
timestamp 0
transform -1 0 2570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2663_
timestamp 0
transform -1 0 1990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2664_
timestamp 0
transform 1 0 890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2665_
timestamp 0
transform -1 0 850 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2666_
timestamp 0
transform -1 0 370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2667_
timestamp 0
transform -1 0 590 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2668_
timestamp 0
transform 1 0 1090 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2669_
timestamp 0
transform -1 0 2850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2670_
timestamp 0
transform -1 0 2970 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2671_
timestamp 0
transform 1 0 1130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2672_
timestamp 0
transform -1 0 630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2673_
timestamp 0
transform -1 0 590 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2674_
timestamp 0
transform 1 0 850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2675_
timestamp 0
transform 1 0 830 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2676_
timestamp 0
transform -1 0 1130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2677_
timestamp 0
transform 1 0 6470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__2678_
timestamp 0
transform -1 0 6390 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2679_
timestamp 0
transform 1 0 7010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2680_
timestamp 0
transform -1 0 6810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2681_
timestamp 0
transform 1 0 7070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2682_
timestamp 0
transform -1 0 6790 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2683_
timestamp 0
transform -1 0 1910 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2684_
timestamp 0
transform -1 0 1730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__2685_
timestamp 0
transform 1 0 1650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2686_
timestamp 0
transform 1 0 1650 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2687_
timestamp 0
transform 1 0 1390 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2688_
timestamp 0
transform -1 0 830 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2689_
timestamp 0
transform -1 0 810 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2690_
timestamp 0
transform 1 0 7310 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2691_
timestamp 0
transform -1 0 7150 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2692_
timestamp 0
transform -1 0 5090 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2693_
timestamp 0
transform -1 0 3050 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2694_
timestamp 0
transform -1 0 1350 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2695_
timestamp 0
transform -1 0 1630 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2696_
timestamp 0
transform -1 0 1350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2697_
timestamp 0
transform 1 0 1930 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2698_
timestamp 0
transform -1 0 570 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2699_
timestamp 0
transform 1 0 6330 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2700_
timestamp 0
transform -1 0 7050 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2701_
timestamp 0
transform 1 0 7630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2702_
timestamp 0
transform 1 0 7330 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2703_
timestamp 0
transform 1 0 7490 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2704_
timestamp 0
transform -1 0 6690 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2705_
timestamp 0
transform 1 0 1610 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2706_
timestamp 0
transform 1 0 1050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2707_
timestamp 0
transform 1 0 2750 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2708_
timestamp 0
transform 1 0 2430 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2709_
timestamp 0
transform -1 0 1110 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2710_
timestamp 0
transform -1 0 890 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2711_
timestamp 0
transform -1 0 1170 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2712_
timestamp 0
transform 1 0 2910 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2713_
timestamp 0
transform -1 0 4310 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2714_
timestamp 0
transform -1 0 4730 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2715_
timestamp 0
transform 1 0 3570 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2716_
timestamp 0
transform -1 0 4330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2717_
timestamp 0
transform -1 0 5890 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__2718_
timestamp 0
transform -1 0 4130 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2719_
timestamp 0
transform 1 0 3730 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2720_
timestamp 0
transform -1 0 4030 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2721_
timestamp 0
transform -1 0 2190 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2722_
timestamp 0
transform 1 0 2310 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2723_
timestamp 0
transform 1 0 2610 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2724_
timestamp 0
transform -1 0 850 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2725_
timestamp 0
transform -1 0 5450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2726_
timestamp 0
transform -1 0 6630 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2727_
timestamp 0
transform 1 0 3890 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2728_
timestamp 0
transform 1 0 3610 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2729_
timestamp 0
transform -1 0 3570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2730_
timestamp 0
transform 1 0 3170 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2731_
timestamp 0
transform 1 0 2030 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2732_
timestamp 0
transform -1 0 1910 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2733_
timestamp 0
transform 1 0 1450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2734_
timestamp 0
transform -1 0 1750 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2735_
timestamp 0
transform -1 0 3910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2736_
timestamp 0
transform -1 0 4050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2737_
timestamp 0
transform -1 0 4130 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2738_
timestamp 0
transform -1 0 3830 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2739_
timestamp 0
transform -1 0 3270 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2740_
timestamp 0
transform -1 0 3350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2741_
timestamp 0
transform -1 0 1110 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2742_
timestamp 0
transform 1 0 1410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2743_
timestamp 0
transform 1 0 1350 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2744_
timestamp 0
transform 1 0 1890 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2745_
timestamp 0
transform 1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2746_
timestamp 0
transform 1 0 3610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2747_
timestamp 0
transform 1 0 4730 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__2748_
timestamp 0
transform 1 0 4390 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2749_
timestamp 0
transform -1 0 3550 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2750_
timestamp 0
transform -1 0 2990 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2751_
timestamp 0
transform 1 0 2830 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2752_
timestamp 0
transform 1 0 1130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2753_
timestamp 0
transform 1 0 630 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2754_
timestamp 0
transform -1 0 570 0 1 790
box -6 -8 26 268
use FILL  FILL_3__2755_
timestamp 0
transform -1 0 3090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2756_
timestamp 0
transform -1 0 2530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2757_
timestamp 0
transform 1 0 2770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2758_
timestamp 0
transform 1 0 2250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2759_
timestamp 0
transform -1 0 4330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2760_
timestamp 0
transform 1 0 3770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2761_
timestamp 0
transform 1 0 4110 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2762_
timestamp 0
transform -1 0 3850 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2763_
timestamp 0
transform -1 0 2090 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2764_
timestamp 0
transform -1 0 1810 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2765_
timestamp 0
transform -1 0 1730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2766_
timestamp 0
transform -1 0 1990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__2767_
timestamp 0
transform -1 0 1510 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__2768_
timestamp 0
transform 1 0 2170 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2769_
timestamp 0
transform 1 0 1610 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__2770_
timestamp 0
transform 1 0 5970 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2771_
timestamp 0
transform 1 0 6510 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2772_
timestamp 0
transform 1 0 4950 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__2773_
timestamp 0
transform 1 0 4150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2774_
timestamp 0
transform 1 0 2310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2775_
timestamp 0
transform 1 0 2550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2776_
timestamp 0
transform 1 0 3370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2777_
timestamp 0
transform -1 0 2850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2778_
timestamp 0
transform -1 0 3110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__2779_
timestamp 0
transform -1 0 7150 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2780_
timestamp 0
transform -1 0 7390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__2781_
timestamp 0
transform 1 0 7870 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__2782_
timestamp 0
transform 1 0 7750 0 1 270
box -6 -8 26 268
use FILL  FILL_3__2783_
timestamp 0
transform 1 0 9690 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2784_
timestamp 0
transform 1 0 10830 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2785_
timestamp 0
transform 1 0 10210 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2786_
timestamp 0
transform 1 0 9930 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2787_
timestamp 0
transform 1 0 8390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2788_
timestamp 0
transform 1 0 8650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2789_
timestamp 0
transform 1 0 8170 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2790_
timestamp 0
transform -1 0 7910 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2791_
timestamp 0
transform 1 0 6170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2792_
timestamp 0
transform 1 0 9790 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2793_
timestamp 0
transform 1 0 9990 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2794_
timestamp 0
transform -1 0 10250 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2795_
timestamp 0
transform 1 0 8430 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2796_
timestamp 0
transform 1 0 8410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2797_
timestamp 0
transform 1 0 10810 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2798_
timestamp 0
transform -1 0 9950 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2799_
timestamp 0
transform -1 0 8330 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2800_
timestamp 0
transform -1 0 7730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2801_
timestamp 0
transform 1 0 9670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2802_
timestamp 0
transform -1 0 9990 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2803_
timestamp 0
transform 1 0 8430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2804_
timestamp 0
transform -1 0 8330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2805_
timestamp 0
transform -1 0 10070 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2806_
timestamp 0
transform 1 0 9750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2807_
timestamp 0
transform -1 0 8370 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2808_
timestamp 0
transform -1 0 6610 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2809_
timestamp 0
transform 1 0 8130 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2810_
timestamp 0
transform -1 0 7550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2811_
timestamp 0
transform 1 0 10030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2812_
timestamp 0
transform 1 0 9670 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2813_
timestamp 0
transform 1 0 8250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2814_
timestamp 0
transform -1 0 8130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2815_
timestamp 0
transform -1 0 8210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2816_
timestamp 0
transform 1 0 9470 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2817_
timestamp 0
transform -1 0 10330 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2818_
timestamp 0
transform 1 0 11150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2819_
timestamp 0
transform 1 0 10130 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2820_
timestamp 0
transform -1 0 9910 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2821_
timestamp 0
transform -1 0 9770 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2822_
timestamp 0
transform -1 0 7490 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2823_
timestamp 0
transform -1 0 9490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2824_
timestamp 0
transform -1 0 9230 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2825_
timestamp 0
transform 1 0 8690 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2826_
timestamp 0
transform 1 0 8730 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2827_
timestamp 0
transform 1 0 9150 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2828_
timestamp 0
transform 1 0 10270 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2829_
timestamp 0
transform -1 0 9210 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2830_
timestamp 0
transform 1 0 9830 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2831_
timestamp 0
transform 1 0 9010 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2832_
timestamp 0
transform -1 0 8930 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2833_
timestamp 0
transform -1 0 8690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2834_
timestamp 0
transform -1 0 8270 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2835_
timestamp 0
transform -1 0 9290 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2836_
timestamp 0
transform -1 0 7990 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2837_
timestamp 0
transform 1 0 8070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2838_
timestamp 0
transform 1 0 9310 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2839_
timestamp 0
transform 1 0 9570 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2840_
timestamp 0
transform -1 0 9310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2841_
timestamp 0
transform 1 0 8210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2842_
timestamp 0
transform 1 0 11530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2843_
timestamp 0
transform -1 0 11030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2844_
timestamp 0
transform 1 0 10750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2845_
timestamp 0
transform 1 0 10490 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2846_
timestamp 0
transform -1 0 10130 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2847_
timestamp 0
transform 1 0 10330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2848_
timestamp 0
transform -1 0 9610 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2849_
timestamp 0
transform 1 0 10910 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__2850_
timestamp 0
transform 1 0 11070 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2851_
timestamp 0
transform 1 0 11310 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2852_
timestamp 0
transform 1 0 12010 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2853_
timestamp 0
transform 1 0 12070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2854_
timestamp 0
transform 1 0 11750 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2855_
timestamp 0
transform 1 0 12030 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2856_
timestamp 0
transform -1 0 9070 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2857_
timestamp 0
transform 1 0 9570 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2858_
timestamp 0
transform -1 0 9870 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2859_
timestamp 0
transform 1 0 10810 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2860_
timestamp 0
transform 1 0 7690 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2861_
timestamp 0
transform 1 0 8370 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2862_
timestamp 0
transform -1 0 7750 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2863_
timestamp 0
transform 1 0 7450 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2864_
timestamp 0
transform 1 0 9690 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2865_
timestamp 0
transform 1 0 8850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2866_
timestamp 0
transform -1 0 6950 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2867_
timestamp 0
transform -1 0 8790 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2868_
timestamp 0
transform -1 0 8510 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2869_
timestamp 0
transform -1 0 8950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2870_
timestamp 0
transform 1 0 8590 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2871_
timestamp 0
transform 1 0 8550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2872_
timestamp 0
transform 1 0 5490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2873_
timestamp 0
transform -1 0 5510 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2874_
timestamp 0
transform 1 0 5430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2875_
timestamp 0
transform -1 0 5790 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2876_
timestamp 0
transform 1 0 5470 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2877_
timestamp 0
transform 1 0 6050 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2878_
timestamp 0
transform -1 0 5790 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2879_
timestamp 0
transform -1 0 8930 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2880_
timestamp 0
transform -1 0 11930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2881_
timestamp 0
transform 1 0 11610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2882_
timestamp 0
transform -1 0 9210 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2883_
timestamp 0
transform 1 0 9010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2884_
timestamp 0
transform -1 0 9330 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2885_
timestamp 0
transform -1 0 10510 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2886_
timestamp 0
transform 1 0 10470 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2887_
timestamp 0
transform -1 0 8890 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2888_
timestamp 0
transform -1 0 9170 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2889_
timestamp 0
transform 1 0 9450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2890_
timestamp 0
transform -1 0 9810 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__2891_
timestamp 0
transform -1 0 9750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2892_
timestamp 0
transform 1 0 9130 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2893_
timestamp 0
transform -1 0 9290 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2894_
timestamp 0
transform -1 0 11110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2895_
timestamp 0
transform 1 0 10790 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2896_
timestamp 0
transform -1 0 11070 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2897_
timestamp 0
transform -1 0 10790 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2898_
timestamp 0
transform 1 0 9410 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2899_
timestamp 0
transform -1 0 9710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2900_
timestamp 0
transform 1 0 10390 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2901_
timestamp 0
transform -1 0 10410 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2902_
timestamp 0
transform 1 0 10590 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2903_
timestamp 0
transform -1 0 10710 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2904_
timestamp 0
transform -1 0 9870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2905_
timestamp 0
transform -1 0 9370 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2906_
timestamp 0
transform -1 0 8530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2907_
timestamp 0
transform -1 0 9090 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2908_
timestamp 0
transform -1 0 10430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2909_
timestamp 0
transform 1 0 11790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2910_
timestamp 0
transform 1 0 10870 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2911_
timestamp 0
transform 1 0 11730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2912_
timestamp 0
transform 1 0 12010 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__2913_
timestamp 0
transform 1 0 10610 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__2914_
timestamp 0
transform -1 0 7790 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2915_
timestamp 0
transform 1 0 10930 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2916_
timestamp 0
transform 1 0 11170 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__2917_
timestamp 0
transform 1 0 10670 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2918_
timestamp 0
transform -1 0 10830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2919_
timestamp 0
transform 1 0 8510 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2920_
timestamp 0
transform 1 0 11210 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2921_
timestamp 0
transform 1 0 11730 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__2922_
timestamp 0
transform -1 0 11850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2923_
timestamp 0
transform 1 0 11310 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2924_
timestamp 0
transform 1 0 10230 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2925_
timestamp 0
transform 1 0 9990 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2926_
timestamp 0
transform 1 0 10130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2927_
timestamp 0
transform -1 0 9970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2928_
timestamp 0
transform -1 0 10230 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__2929_
timestamp 0
transform -1 0 10350 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__2930_
timestamp 0
transform -1 0 11230 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2931_
timestamp 0
transform -1 0 11490 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__2932_
timestamp 0
transform 1 0 11450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__2933_
timestamp 0
transform 1 0 11410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__2934_
timestamp 0
transform 1 0 11490 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__2935_
timestamp 0
transform 1 0 11570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2936_
timestamp 0
transform 1 0 10510 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__2937_
timestamp 0
transform -1 0 3510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__2938_
timestamp 0
transform -1 0 7730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2939_
timestamp 0
transform 1 0 6490 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2940_
timestamp 0
transform -1 0 6270 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2941_
timestamp 0
transform -1 0 6190 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2942_
timestamp 0
transform 1 0 5090 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2943_
timestamp 0
transform -1 0 6990 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__2944_
timestamp 0
transform 1 0 5370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2945_
timestamp 0
transform -1 0 6770 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2946_
timestamp 0
transform 1 0 6370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__2947_
timestamp 0
transform 1 0 7850 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2948_
timestamp 0
transform 1 0 7590 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2949_
timestamp 0
transform 1 0 5690 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__2950_
timestamp 0
transform -1 0 6030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2951_
timestamp 0
transform 1 0 6790 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2952_
timestamp 0
transform 1 0 6510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2953_
timestamp 0
transform 1 0 5670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2954_
timestamp 0
transform -1 0 5970 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__2955_
timestamp 0
transform 1 0 7050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2956_
timestamp 0
transform 1 0 6530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__2957_
timestamp 0
transform -1 0 8150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__2958_
timestamp 0
transform 1 0 6530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__2959_
timestamp 0
transform 1 0 6270 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2960_
timestamp 0
transform -1 0 7150 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2961_
timestamp 0
transform 1 0 6530 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2962_
timestamp 0
transform -1 0 6310 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__2963_
timestamp 0
transform -1 0 6610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2964_
timestamp 0
transform 1 0 4670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2965_
timestamp 0
transform 1 0 5730 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2966_
timestamp 0
transform -1 0 6630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__2967_
timestamp 0
transform -1 0 5050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2968_
timestamp 0
transform -1 0 5310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2969_
timestamp 0
transform 1 0 4390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2970_
timestamp 0
transform 1 0 4750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2971_
timestamp 0
transform 1 0 4630 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2972_
timestamp 0
transform -1 0 6070 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2973_
timestamp 0
transform -1 0 6330 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2974_
timestamp 0
transform -1 0 6330 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2975_
timestamp 0
transform 1 0 5790 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2976_
timestamp 0
transform -1 0 4710 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2977_
timestamp 0
transform -1 0 4970 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2978_
timestamp 0
transform 1 0 5230 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__2979_
timestamp 0
transform 1 0 5510 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__2980_
timestamp 0
transform -1 0 7390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2981_
timestamp 0
transform -1 0 6350 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2982_
timestamp 0
transform -1 0 6630 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__2983_
timestamp 0
transform 1 0 7150 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2984_
timestamp 0
transform 1 0 6550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__2985_
timestamp 0
transform -1 0 6890 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2986_
timestamp 0
transform 1 0 6590 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2987_
timestamp 0
transform 1 0 6030 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2988_
timestamp 0
transform -1 0 6310 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__2989_
timestamp 0
transform -1 0 7890 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2990_
timestamp 0
transform 1 0 7010 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__2991_
timestamp 0
transform -1 0 6870 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2992_
timestamp 0
transform -1 0 5170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__2993_
timestamp 0
transform -1 0 6030 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2994_
timestamp 0
transform 1 0 5490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2995_
timestamp 0
transform 1 0 6570 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2996_
timestamp 0
transform 1 0 6290 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__2997_
timestamp 0
transform 1 0 6010 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2998_
timestamp 0
transform -1 0 5750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__2999_
timestamp 0
transform 1 0 6410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3000_
timestamp 0
transform -1 0 5750 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__3001_
timestamp 0
transform 1 0 4970 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3002_
timestamp 0
transform -1 0 5470 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__3003_
timestamp 0
transform -1 0 5830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3004_
timestamp 0
transform -1 0 5250 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3005_
timestamp 0
transform -1 0 5510 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3006_
timestamp 0
transform -1 0 7410 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3007_
timestamp 0
transform 1 0 6830 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3008_
timestamp 0
transform 1 0 8630 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3009_
timestamp 0
transform 1 0 8090 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3010_
timestamp 0
transform 1 0 7110 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3011_
timestamp 0
transform -1 0 7210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3012_
timestamp 0
transform -1 0 7090 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3013_
timestamp 0
transform -1 0 7830 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3014_
timestamp 0
transform 1 0 7030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3015_
timestamp 0
transform -1 0 7310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3016_
timestamp 0
transform -1 0 6070 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3017_
timestamp 0
transform -1 0 6870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3018_
timestamp 0
transform -1 0 6550 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3019_
timestamp 0
transform -1 0 6810 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3020_
timestamp 0
transform 1 0 5450 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__3021_
timestamp 0
transform 1 0 5890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3022_
timestamp 0
transform 1 0 5690 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__3023_
timestamp 0
transform -1 0 6770 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3024_
timestamp 0
transform -1 0 6690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3025_
timestamp 0
transform 1 0 5970 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__3026_
timestamp 0
transform 1 0 5390 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__3027_
timestamp 0
transform -1 0 5490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3028_
timestamp 0
transform 1 0 5970 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3029_
timestamp 0
transform 1 0 6730 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3030_
timestamp 0
transform 1 0 4870 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__3031_
timestamp 0
transform 1 0 4410 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3032_
timestamp 0
transform -1 0 5190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3033_
timestamp 0
transform 1 0 5450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3034_
timestamp 0
transform -1 0 3390 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3035_
timestamp 0
transform -1 0 3950 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3036_
timestamp 0
transform -1 0 3450 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3037_
timestamp 0
transform -1 0 3330 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3038_
timestamp 0
transform 1 0 3550 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3039_
timestamp 0
transform -1 0 3050 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3040_
timestamp 0
transform 1 0 2930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3041_
timestamp 0
transform 1 0 3170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3042_
timestamp 0
transform -1 0 3730 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3043_
timestamp 0
transform -1 0 3830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3044_
timestamp 0
transform -1 0 3590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3045_
timestamp 0
transform 1 0 4390 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3046_
timestamp 0
transform 1 0 4110 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3047_
timestamp 0
transform -1 0 3070 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3048_
timestamp 0
transform 1 0 3110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3049_
timestamp 0
transform -1 0 2810 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3050_
timestamp 0
transform 1 0 2850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3051_
timestamp 0
transform 1 0 2590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3052_
timestamp 0
transform 1 0 2490 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3053_
timestamp 0
transform 1 0 3250 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3054_
timestamp 0
transform -1 0 3530 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3055_
timestamp 0
transform 1 0 3350 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3056_
timestamp 0
transform -1 0 3610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3057_
timestamp 0
transform 1 0 3810 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3058_
timestamp 0
transform 1 0 3990 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3059_
timestamp 0
transform 1 0 4270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3060_
timestamp 0
transform 1 0 4110 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3061_
timestamp 0
transform 1 0 3590 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3062_
timestamp 0
transform -1 0 3830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3063_
timestamp 0
transform -1 0 5070 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__3064_
timestamp 0
transform 1 0 4930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__3065_
timestamp 0
transform -1 0 4670 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3066_
timestamp 0
transform 1 0 4570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3067_
timestamp 0
transform -1 0 3670 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3068_
timestamp 0
transform -1 0 3410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3069_
timestamp 0
transform 1 0 3610 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3070_
timestamp 0
transform -1 0 4510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__3071_
timestamp 0
transform 1 0 4230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__3072_
timestamp 0
transform -1 0 4170 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3073_
timestamp 0
transform -1 0 4430 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3074_
timestamp 0
transform 1 0 5710 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3075_
timestamp 0
transform 1 0 5430 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3076_
timestamp 0
transform 1 0 3670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3077_
timestamp 0
transform 1 0 3990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3078_
timestamp 0
transform 1 0 4050 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3079_
timestamp 0
transform -1 0 4130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3080_
timestamp 0
transform 1 0 6270 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3081_
timestamp 0
transform -1 0 6930 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3082_
timestamp 0
transform 1 0 6630 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3083_
timestamp 0
transform -1 0 3810 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3084_
timestamp 0
transform 1 0 3510 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3085_
timestamp 0
transform 1 0 3130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3086_
timestamp 0
transform -1 0 2850 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3087_
timestamp 0
transform 1 0 4330 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3088_
timestamp 0
transform -1 0 4930 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3089_
timestamp 0
transform 1 0 3410 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3090_
timestamp 0
transform -1 0 3690 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3091_
timestamp 0
transform -1 0 6230 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3092_
timestamp 0
transform 1 0 5450 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3093_
timestamp 0
transform 1 0 5710 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3094_
timestamp 0
transform 1 0 5430 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3095_
timestamp 0
transform -1 0 4630 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3096_
timestamp 0
transform 1 0 4330 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3097_
timestamp 0
transform -1 0 4090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3098_
timestamp 0
transform 1 0 3790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3099_
timestamp 0
transform -1 0 3850 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3100_
timestamp 0
transform -1 0 3670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3101_
timestamp 0
transform 1 0 4890 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3102_
timestamp 0
transform -1 0 5190 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3103_
timestamp 0
transform -1 0 4570 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3104_
timestamp 0
transform -1 0 4850 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3105_
timestamp 0
transform 1 0 5630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3106_
timestamp 0
transform -1 0 5930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3107_
timestamp 0
transform -1 0 4030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3108_
timestamp 0
transform 1 0 3730 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3109_
timestamp 0
transform 1 0 6210 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3110_
timestamp 0
transform 1 0 3890 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3111_
timestamp 0
transform 1 0 5750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3112_
timestamp 0
transform -1 0 5170 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3113_
timestamp 0
transform -1 0 4630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3114_
timestamp 0
transform 1 0 4330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3115_
timestamp 0
transform 1 0 4850 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3116_
timestamp 0
transform 1 0 3790 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3117_
timestamp 0
transform 1 0 4410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3118_
timestamp 0
transform -1 0 4710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3119_
timestamp 0
transform 1 0 4890 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3120_
timestamp 0
transform 1 0 4590 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3121_
timestamp 0
transform 1 0 5190 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3122_
timestamp 0
transform 1 0 5470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3123_
timestamp 0
transform 1 0 5450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3124_
timestamp 0
transform -1 0 5750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3125_
timestamp 0
transform -1 0 4110 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3126_
timestamp 0
transform 1 0 3810 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3127_
timestamp 0
transform 1 0 6470 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3128_
timestamp 0
transform 1 0 6030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3129_
timestamp 0
transform 1 0 5430 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3130_
timestamp 0
transform -1 0 3350 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3131_
timestamp 0
transform -1 0 3590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3132_
timestamp 0
transform 1 0 4690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3133_
timestamp 0
transform 1 0 3930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3134_
timestamp 0
transform 1 0 5110 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3135_
timestamp 0
transform 1 0 4810 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3136_
timestamp 0
transform 1 0 5710 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3137_
timestamp 0
transform 1 0 5430 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3138_
timestamp 0
transform 1 0 5710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3139_
timestamp 0
transform 1 0 5430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3140_
timestamp 0
transform -1 0 5630 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3141_
timestamp 0
transform -1 0 5890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3142_
timestamp 0
transform -1 0 4230 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3143_
timestamp 0
transform -1 0 4490 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3144_
timestamp 0
transform 1 0 11570 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__3145_
timestamp 0
transform 1 0 11810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__3146_
timestamp 0
transform -1 0 11870 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__3147_
timestamp 0
transform 1 0 9490 0 1 790
box -6 -8 26 268
use FILL  FILL_3__3148_
timestamp 0
transform -1 0 11870 0 1 790
box -6 -8 26 268
use FILL  FILL_3__3149_
timestamp 0
transform -1 0 11490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3150_
timestamp 0
transform -1 0 11770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3151_
timestamp 0
transform -1 0 10710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3152_
timestamp 0
transform 1 0 9350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3153_
timestamp 0
transform -1 0 9650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3154_
timestamp 0
transform -1 0 10170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3155_
timestamp 0
transform -1 0 10290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3156_
timestamp 0
transform -1 0 8930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__3157_
timestamp 0
transform -1 0 8970 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__3158_
timestamp 0
transform -1 0 8690 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__3159_
timestamp 0
transform -1 0 8670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__3160_
timestamp 0
transform 1 0 10510 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3161_
timestamp 0
transform 1 0 10230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3162_
timestamp 0
transform -1 0 9770 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3163_
timestamp 0
transform 1 0 9490 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3164_
timestamp 0
transform -1 0 8970 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3165_
timestamp 0
transform -1 0 7190 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3166_
timestamp 0
transform 1 0 7590 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__3167_
timestamp 0
transform 1 0 7450 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3168_
timestamp 0
transform 1 0 7610 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3169_
timestamp 0
transform -1 0 8690 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3170_
timestamp 0
transform -1 0 8410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3171_
timestamp 0
transform -1 0 9130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3172_
timestamp 0
transform -1 0 8130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3173_
timestamp 0
transform 1 0 8390 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3174_
timestamp 0
transform 1 0 7870 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3175_
timestamp 0
transform -1 0 7850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3176_
timestamp 0
transform -1 0 7570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3177_
timestamp 0
transform -1 0 11850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__3178_
timestamp 0
transform -1 0 11790 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3179_
timestamp 0
transform 1 0 12050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3180_
timestamp 0
transform 1 0 12110 0 1 790
box -6 -8 26 268
use FILL  FILL_3__3181_
timestamp 0
transform 1 0 12090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__3182_
timestamp 0
transform -1 0 11310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3183_
timestamp 0
transform 1 0 11570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3184_
timestamp 0
transform 1 0 11850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3185_
timestamp 0
transform 1 0 11870 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3186_
timestamp 0
transform 1 0 12050 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3187_
timestamp 0
transform 1 0 9910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__3188_
timestamp 0
transform 1 0 10790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3189_
timestamp 0
transform -1 0 11050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__3190_
timestamp 0
transform 1 0 11090 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3191_
timestamp 0
transform 1 0 11030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3192_
timestamp 0
transform -1 0 10750 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3193_
timestamp 0
transform 1 0 10170 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3194_
timestamp 0
transform 1 0 10790 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__3195_
timestamp 0
transform -1 0 10530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3196_
timestamp 0
transform 1 0 10430 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3197_
timestamp 0
transform -1 0 7290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3198_
timestamp 0
transform -1 0 4650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3199_
timestamp 0
transform 1 0 2810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__3200_
timestamp 0
transform 1 0 4790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__3201_
timestamp 0
transform 1 0 4510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__3202_
timestamp 0
transform 1 0 1570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__3203_
timestamp 0
transform 1 0 1530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3204_
timestamp 0
transform 1 0 1490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__3205_
timestamp 0
transform 1 0 1050 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__3206_
timestamp 0
transform 1 0 1470 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__3207_
timestamp 0
transform -1 0 1610 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__3208_
timestamp 0
transform -1 0 950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__3209_
timestamp 0
transform -1 0 650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__3210_
timestamp 0
transform -1 0 4310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__3211_
timestamp 0
transform 1 0 4250 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__3212_
timestamp 0
transform 1 0 1210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__3213_
timestamp 0
transform 1 0 1110 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__3214_
timestamp 0
transform -1 0 2390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3215_
timestamp 0
transform 1 0 1810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3216_
timestamp 0
transform 1 0 5750 0 1 270
box -6 -8 26 268
use FILL  FILL_3__3217_
timestamp 0
transform -1 0 6050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__3218_
timestamp 0
transform 1 0 6090 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3219_
timestamp 0
transform -1 0 6370 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3220_
timestamp 0
transform 1 0 3710 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3221_
timestamp 0
transform -1 0 3990 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3222_
timestamp 0
transform -1 0 3590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3223_
timestamp 0
transform 1 0 3310 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__3224_
timestamp 0
transform -1 0 3290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3225_
timestamp 0
transform 1 0 5430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__3226_
timestamp 0
transform 1 0 5150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__3227_
timestamp 0
transform -1 0 4270 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3228_
timestamp 0
transform -1 0 4470 0 1 270
box -6 -8 26 268
use FILL  FILL_3__3229_
timestamp 0
transform 1 0 2710 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__3230_
timestamp 0
transform -1 0 2750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__3231_
timestamp 0
transform 1 0 5990 0 1 790
box -6 -8 26 268
use FILL  FILL_3__3232_
timestamp 0
transform 1 0 5970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__3364_
timestamp 0
transform 1 0 5250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3365_
timestamp 0
transform 1 0 4450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3366_
timestamp 0
transform 1 0 4930 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__3367_
timestamp 0
transform -1 0 4730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3368_
timestamp 0
transform -1 0 4990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3369_
timestamp 0
transform -1 0 5550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3370_
timestamp 0
transform 1 0 2690 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3371_
timestamp 0
transform 1 0 2190 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3372_
timestamp 0
transform -1 0 2310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3373_
timestamp 0
transform -1 0 3970 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3374_
timestamp 0
transform -1 0 2290 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3375_
timestamp 0
transform 1 0 2290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3376_
timestamp 0
transform -1 0 2950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3377_
timestamp 0
transform 1 0 2410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3378_
timestamp 0
transform -1 0 2270 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3379_
timestamp 0
transform -1 0 1430 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3380_
timestamp 0
transform 1 0 1210 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3381_
timestamp 0
transform -1 0 1470 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3382_
timestamp 0
transform -1 0 1930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3383_
timestamp 0
transform -1 0 1490 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3384_
timestamp 0
transform 1 0 1750 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3385_
timestamp 0
transform 1 0 1450 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3386_
timestamp 0
transform -1 0 2030 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3387_
timestamp 0
transform 1 0 2290 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3388_
timestamp 0
transform -1 0 630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3389_
timestamp 0
transform 1 0 2490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3390_
timestamp 0
transform 1 0 3310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3391_
timestamp 0
transform 1 0 3030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3392_
timestamp 0
transform -1 0 2870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3393_
timestamp 0
transform 1 0 2270 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3394_
timestamp 0
transform 1 0 670 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3395_
timestamp 0
transform -1 0 630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3396_
timestamp 0
transform -1 0 370 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3397_
timestamp 0
transform -1 0 390 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3398_
timestamp 0
transform -1 0 90 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3399_
timestamp 0
transform 1 0 70 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3400_
timestamp 0
transform -1 0 870 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3401_
timestamp 0
transform -1 0 1450 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3402_
timestamp 0
transform 1 0 1430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3403_
timestamp 0
transform 1 0 1150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3404_
timestamp 0
transform -1 0 90 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3405_
timestamp 0
transform -1 0 350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3406_
timestamp 0
transform -1 0 90 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3407_
timestamp 0
transform -1 0 370 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3408_
timestamp 0
transform -1 0 90 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3409_
timestamp 0
transform -1 0 90 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3410_
timestamp 0
transform 1 0 1410 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3411_
timestamp 0
transform 1 0 1130 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3412_
timestamp 0
transform -1 0 610 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3413_
timestamp 0
transform 1 0 350 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3414_
timestamp 0
transform 1 0 610 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3__3415_
timestamp 0
transform -1 0 930 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3416_
timestamp 0
transform 1 0 610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3417_
timestamp 0
transform -1 0 650 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3418_
timestamp 0
transform -1 0 350 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3419_
timestamp 0
transform -1 0 1170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3420_
timestamp 0
transform 1 0 870 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3421_
timestamp 0
transform 1 0 1170 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3422_
timestamp 0
transform 1 0 890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3423_
timestamp 0
transform 1 0 1190 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3424_
timestamp 0
transform -1 0 1210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3425_
timestamp 0
transform -1 0 930 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3426_
timestamp 0
transform 1 0 910 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3__3427_
timestamp 0
transform -1 0 1430 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3428_
timestamp 0
transform 1 0 1110 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3429_
timestamp 0
transform -1 0 890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3430_
timestamp 0
transform 1 0 1410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3431_
timestamp 0
transform 1 0 1130 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3432_
timestamp 0
transform -1 0 930 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3433_
timestamp 0
transform -1 0 90 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3434_
timestamp 0
transform -1 0 670 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3435_
timestamp 0
transform -1 0 950 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3436_
timestamp 0
transform -1 0 890 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3437_
timestamp 0
transform 1 0 1710 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3438_
timestamp 0
transform 1 0 1170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3439_
timestamp 0
transform -1 0 1450 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3440_
timestamp 0
transform 1 0 1170 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3441_
timestamp 0
transform -1 0 610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3442_
timestamp 0
transform 1 0 1190 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3443_
timestamp 0
transform 1 0 1110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3444_
timestamp 0
transform -1 0 2010 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3445_
timestamp 0
transform 1 0 1690 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3446_
timestamp 0
transform 1 0 2050 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3447_
timestamp 0
transform 1 0 1950 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3448_
timestamp 0
transform -1 0 1750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3449_
timestamp 0
transform 1 0 1430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3450_
timestamp 0
transform -1 0 890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3451_
timestamp 0
transform 1 0 1150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3452_
timestamp 0
transform 1 0 850 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3453_
timestamp 0
transform -1 0 2170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3454_
timestamp 0
transform 1 0 3090 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3455_
timestamp 0
transform -1 0 2030 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3456_
timestamp 0
transform -1 0 1690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3457_
timestamp 0
transform -1 0 2870 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3458_
timestamp 0
transform -1 0 1730 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3459_
timestamp 0
transform -1 0 1670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3460_
timestamp 0
transform 1 0 1710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3461_
timestamp 0
transform -1 0 1930 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3462_
timestamp 0
transform -1 0 1690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3463_
timestamp 0
transform -1 0 1450 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3464_
timestamp 0
transform 1 0 1170 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3465_
timestamp 0
transform -1 0 1430 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3466_
timestamp 0
transform 1 0 1970 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3467_
timestamp 0
transform 1 0 1970 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3468_
timestamp 0
transform 1 0 2730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3469_
timestamp 0
transform 1 0 2590 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3470_
timestamp 0
transform -1 0 2490 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3471_
timestamp 0
transform 1 0 2310 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3472_
timestamp 0
transform -1 0 2210 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3473_
timestamp 0
transform 1 0 1450 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3474_
timestamp 0
transform -1 0 1710 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3475_
timestamp 0
transform 1 0 1190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3476_
timestamp 0
transform -1 0 930 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3477_
timestamp 0
transform 1 0 350 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3478_
timestamp 0
transform -1 0 330 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3479_
timestamp 0
transform -1 0 90 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3480_
timestamp 0
transform -1 0 90 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3481_
timestamp 0
transform -1 0 90 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3482_
timestamp 0
transform 1 0 610 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3483_
timestamp 0
transform -1 0 330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3484_
timestamp 0
transform 1 0 1950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3485_
timestamp 0
transform -1 0 2010 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3486_
timestamp 0
transform -1 0 1390 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3487_
timestamp 0
transform -1 0 1710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3488_
timestamp 0
transform -1 0 1510 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3489_
timestamp 0
transform 1 0 1450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3490_
timestamp 0
transform 1 0 1130 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3491_
timestamp 0
transform -1 0 1210 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3492_
timestamp 0
transform 1 0 1110 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3493_
timestamp 0
transform -1 0 930 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3494_
timestamp 0
transform 1 0 850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3495_
timestamp 0
transform -1 0 610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3496_
timestamp 0
transform 1 0 370 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3497_
timestamp 0
transform -1 0 330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3498_
timestamp 0
transform 1 0 630 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3499_
timestamp 0
transform -1 0 690 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3500_
timestamp 0
transform 1 0 630 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3501_
timestamp 0
transform 1 0 870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3502_
timestamp 0
transform -1 0 390 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3503_
timestamp 0
transform -1 0 370 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3504_
timestamp 0
transform -1 0 610 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3505_
timestamp 0
transform -1 0 370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3506_
timestamp 0
transform -1 0 90 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3507_
timestamp 0
transform -1 0 90 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3508_
timestamp 0
transform 1 0 610 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3509_
timestamp 0
transform -1 0 870 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3510_
timestamp 0
transform -1 0 370 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3511_
timestamp 0
transform -1 0 90 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3512_
timestamp 0
transform 1 0 570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3513_
timestamp 0
transform -1 0 390 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3514_
timestamp 0
transform -1 0 330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3515_
timestamp 0
transform -1 0 90 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3516_
timestamp 0
transform -1 0 90 0 1 10150
box -6 -8 26 268
use FILL  FILL_3__3517_
timestamp 0
transform 1 0 630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3518_
timestamp 0
transform 1 0 850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3519_
timestamp 0
transform 1 0 2550 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3520_
timestamp 0
transform 1 0 2830 0 1 9110
box -6 -8 26 268
use FILL  FILL_3__3521_
timestamp 0
transform 1 0 3310 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3522_
timestamp 0
transform 1 0 3010 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3523_
timestamp 0
transform 1 0 2570 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3524_
timestamp 0
transform -1 0 950 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3525_
timestamp 0
transform -1 0 90 0 1 10670
box -6 -8 26 268
use FILL  FILL_3__3526_
timestamp 0
transform -1 0 90 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3527_
timestamp 0
transform -1 0 590 0 1 11190
box -6 -8 26 268
use FILL  FILL_3__3528_
timestamp 0
transform -1 0 610 0 -1 10670
box -6 -8 26 268
use FILL  FILL_3__3529_
timestamp 0
transform -1 0 90 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3__3530_
timestamp 0
transform -1 0 90 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3531_
timestamp 0
transform 1 0 70 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3532_
timestamp 0
transform 1 0 310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3533_
timestamp 0
transform -1 0 90 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3534_
timestamp 0
transform -1 0 610 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3535_
timestamp 0
transform -1 0 370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3__3536_
timestamp 0
transform -1 0 350 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3537_
timestamp 0
transform -1 0 1710 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3538_
timestamp 0
transform 1 0 2470 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3539_
timestamp 0
transform -1 0 2570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3540_
timestamp 0
transform -1 0 2310 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3541_
timestamp 0
transform -1 0 2030 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3542_
timestamp 0
transform -1 0 2210 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3543_
timestamp 0
transform 1 0 1610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3544_
timestamp 0
transform 1 0 1970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3545_
timestamp 0
transform 1 0 1770 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3546_
timestamp 0
transform 1 0 1890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3__3547_
timestamp 0
transform -1 0 2550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3548_
timestamp 0
transform 1 0 2250 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3__3549_
timestamp 0
transform -1 0 2350 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3550_
timestamp 0
transform 1 0 2050 0 1 11710
box -6 -8 26 268
use FILL  FILL_3__3551_
timestamp 0
transform -1 0 2530 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3552_
timestamp 0
transform 1 0 2230 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3__3553_
timestamp 0
transform -1 0 1770 0 1 8070
box -6 -8 26 268
use FILL  FILL_3__3554_
timestamp 0
transform 1 0 910 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3555_
timestamp 0
transform 1 0 310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3556_
timestamp 0
transform 1 0 1170 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3__3557_
timestamp 0
transform -1 0 3070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3558_
timestamp 0
transform 1 0 2770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3__3559_
timestamp 0
transform -1 0 2530 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3560_
timestamp 0
transform 1 0 2230 0 1 9630
box -6 -8 26 268
use FILL  FILL_3__3561_
timestamp 0
transform -1 0 1950 0 1 7550
box -6 -8 26 268
use FILL  FILL_3__3562_
timestamp 0
transform -1 0 2770 0 1 8590
box -6 -8 26 268
use FILL  FILL_3__3563_
timestamp 0
transform 1 0 2170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3__3564_
timestamp 0
transform 1 0 2450 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3565_
timestamp 0
transform -1 0 1450 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3566_
timestamp 0
transform -1 0 1710 0 1 7030
box -6 -8 26 268
use FILL  FILL_3__3579_
timestamp 0
transform -1 0 5050 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3580_
timestamp 0
transform -1 0 90 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__3581_
timestamp 0
transform -1 0 3470 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3582_
timestamp 0
transform -1 0 3210 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3583_
timestamp 0
transform -1 0 5330 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__3584_
timestamp 0
transform 1 0 4510 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3585_
timestamp 0
transform 1 0 2930 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3586_
timestamp 0
transform -1 0 5850 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__3587_
timestamp 0
transform 1 0 70 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3588_
timestamp 0
transform -1 0 90 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__3589_
timestamp 0
transform -1 0 90 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__3590_
timestamp 0
transform -1 0 90 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__3591_
timestamp 0
transform -1 0 370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3592_
timestamp 0
transform -1 0 90 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__3593_
timestamp 0
transform -1 0 4790 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3594_
timestamp 0
transform 1 0 5830 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__3595_
timestamp 0
transform 1 0 5570 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__3596_
timestamp 0
transform -1 0 870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3597_
timestamp 0
transform -1 0 90 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__3598_
timestamp 0
transform -1 0 350 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__3599_
timestamp 0
transform -1 0 90 0 1 6510
box -6 -8 26 268
use FILL  FILL_3__3600_
timestamp 0
transform -1 0 90 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__3601_
timestamp 0
transform -1 0 90 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__3602_
timestamp 0
transform -1 0 1710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__3603_
timestamp 0
transform 1 0 6870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert0
timestamp 0
transform 1 0 7890 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert1
timestamp 0
transform 1 0 9390 0 1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert2
timestamp 0
transform 1 0 8150 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert3
timestamp 0
transform 1 0 11010 0 1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert4
timestamp 0
transform 1 0 610 0 1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert5
timestamp 0
transform -1 0 12090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert6
timestamp 0
transform -1 0 9590 0 1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert7
timestamp 0
transform 1 0 7050 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert8
timestamp 0
transform -1 0 870 0 1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert9
timestamp 0
transform 1 0 10130 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert10
timestamp 0
transform -1 0 910 0 1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert11
timestamp 0
transform -1 0 5990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform 1 0 11550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform -1 0 6170 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform 1 0 6790 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform -1 0 3330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform -1 0 3950 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform 1 0 7190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert18
timestamp 0
transform -1 0 7010 0 1 11190
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform 1 0 5330 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert20
timestamp 0
transform 1 0 8570 0 1 11190
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert21
timestamp 0
transform -1 0 8490 0 -1 7550
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert22
timestamp 0
transform -1 0 1450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert23
timestamp 0
transform 1 0 3430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert24
timestamp 0
transform -1 0 4330 0 1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert25
timestamp 0
transform 1 0 8170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert26
timestamp 0
transform 1 0 5110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert27
timestamp 0
transform -1 0 1250 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert39
timestamp 0
transform 1 0 6330 0 1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert40
timestamp 0
transform 1 0 7690 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert41
timestamp 0
transform -1 0 8830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert42
timestamp 0
transform -1 0 6970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert43
timestamp 0
transform -1 0 8870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert44
timestamp 0
transform -1 0 8990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert45
timestamp 0
transform 1 0 11050 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert46
timestamp 0
transform 1 0 9490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert47
timestamp 0
transform 1 0 9210 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert48
timestamp 0
transform 1 0 6950 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert49
timestamp 0
transform 1 0 7210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert50
timestamp 0
transform -1 0 7590 0 1 9110
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert51
timestamp 0
transform 1 0 7550 0 1 10150
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert52
timestamp 0
transform 1 0 8950 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert53
timestamp 0
transform 1 0 9990 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert54
timestamp 0
transform 1 0 8830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert55
timestamp 0
transform 1 0 8690 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert56
timestamp 0
transform -1 0 2230 0 1 8590
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert57
timestamp 0
transform 1 0 2530 0 1 11190
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert58
timestamp 0
transform 1 0 2670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert59
timestamp 0
transform -1 0 2230 0 1 10670
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert60
timestamp 0
transform -1 0 10490 0 1 7550
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert61
timestamp 0
transform 1 0 10550 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert62
timestamp 0
transform 1 0 10510 0 1 8070
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert63
timestamp 0
transform -1 0 9170 0 1 7550
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert64
timestamp 0
transform -1 0 8610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert65
timestamp 0
transform 1 0 5210 0 1 270
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert66
timestamp 0
transform 1 0 5730 0 1 790
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert67
timestamp 0
transform -1 0 3030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert68
timestamp 0
transform 1 0 3150 0 1 270
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert69
timestamp 0
transform -1 0 6650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert70
timestamp 0
transform 1 0 8590 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert71
timestamp 0
transform -1 0 9250 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert72
timestamp 0
transform -1 0 6770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert73
timestamp 0
transform 1 0 8930 0 -1 7030
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert74
timestamp 0
transform 1 0 10790 0 1 7030
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert75
timestamp 0
transform 1 0 2570 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert76
timestamp 0
transform -1 0 3070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert77
timestamp 0
transform 1 0 10450 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert78
timestamp 0
transform 1 0 9310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert79
timestamp 0
transform -1 0 8350 0 1 7550
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert80
timestamp 0
transform 1 0 7150 0 1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert81
timestamp 0
transform 1 0 7610 0 -1 790
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert82
timestamp 0
transform -1 0 7590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert83
timestamp 0
transform -1 0 7370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert84
timestamp 0
transform 1 0 9430 0 1 8590
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert85
timestamp 0
transform -1 0 8910 0 1 8590
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert86
timestamp 0
transform -1 0 9510 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert87
timestamp 0
transform 1 0 9410 0 1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert88
timestamp 0
transform -1 0 10750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert89
timestamp 0
transform 1 0 9390 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert90
timestamp 0
transform 1 0 5370 0 -1 11190
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert91
timestamp 0
transform -1 0 4910 0 1 10670
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert92
timestamp 0
transform -1 0 4750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert93
timestamp 0
transform 1 0 5170 0 1 10150
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert94
timestamp 0
transform -1 0 11330 0 1 9630
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert95
timestamp 0
transform -1 0 11370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert96
timestamp 0
transform -1 0 10090 0 1 11710
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert97
timestamp 0
transform 1 0 11450 0 1 11710
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert28
timestamp 0
transform -1 0 6030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert29
timestamp 0
transform -1 0 2210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert30
timestamp 0
transform 1 0 4550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert31
timestamp 0
transform -1 0 3250 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert32
timestamp 0
transform 1 0 7150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert33
timestamp 0
transform 1 0 5730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert34
timestamp 0
transform -1 0 2490 0 1 10670
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert35
timestamp 0
transform -1 0 5250 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert36
timestamp 0
transform -1 0 2370 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert37
timestamp 0
transform 1 0 7390 0 -1 12230
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert38
timestamp 0
transform -1 0 4370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__1688_
timestamp 0
transform -1 0 910 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1689_
timestamp 0
transform -1 0 370 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1690_
timestamp 0
transform -1 0 630 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1691_
timestamp 0
transform 1 0 90 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1692_
timestamp 0
transform -1 0 350 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1693_
timestamp 0
transform 1 0 590 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1694_
timestamp 0
transform -1 0 5590 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1695_
timestamp 0
transform -1 0 370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1696_
timestamp 0
transform -1 0 370 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1697_
timestamp 0
transform -1 0 1490 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__1698_
timestamp 0
transform -1 0 3430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1699_
timestamp 0
transform 1 0 2870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1700_
timestamp 0
transform -1 0 3910 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__1701_
timestamp 0
transform -1 0 610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1702_
timestamp 0
transform -1 0 610 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1703_
timestamp 0
transform 1 0 3250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1704_
timestamp 0
transform -1 0 390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1705_
timestamp 0
transform 1 0 90 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1706_
timestamp 0
transform -1 0 3870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1707_
timestamp 0
transform -1 0 630 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1708_
timestamp 0
transform 1 0 630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1709_
timestamp 0
transform 1 0 4150 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1710_
timestamp 0
transform -1 0 5630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1711_
timestamp 0
transform 1 0 5170 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1712_
timestamp 0
transform 1 0 7310 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1713_
timestamp 0
transform -1 0 9690 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1714_
timestamp 0
transform -1 0 9890 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1715_
timestamp 0
transform -1 0 8570 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1716_
timestamp 0
transform 1 0 11330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1717_
timestamp 0
transform 1 0 11130 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1718_
timestamp 0
transform 1 0 11950 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1719_
timestamp 0
transform -1 0 8830 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1720_
timestamp 0
transform -1 0 10150 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1721_
timestamp 0
transform -1 0 10170 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1722_
timestamp 0
transform -1 0 9930 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1723_
timestamp 0
transform 1 0 10030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1724_
timestamp 0
transform 1 0 9250 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1725_
timestamp 0
transform 1 0 9090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1726_
timestamp 0
transform 1 0 10190 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1727_
timestamp 0
transform -1 0 8810 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1728_
timestamp 0
transform 1 0 11590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1729_
timestamp 0
transform 1 0 10190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1730_
timestamp 0
transform 1 0 8370 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1731_
timestamp 0
transform 1 0 8610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1732_
timestamp 0
transform -1 0 7810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1733_
timestamp 0
transform 1 0 9750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1734_
timestamp 0
transform 1 0 7450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1735_
timestamp 0
transform 1 0 10890 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1736_
timestamp 0
transform -1 0 10690 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1737_
timestamp 0
transform -1 0 10950 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1738_
timestamp 0
transform -1 0 10330 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1739_
timestamp 0
transform -1 0 10330 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1740_
timestamp 0
transform 1 0 10550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1741_
timestamp 0
transform -1 0 8450 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1742_
timestamp 0
transform -1 0 8350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1743_
timestamp 0
transform -1 0 9910 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1744_
timestamp 0
transform 1 0 9790 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1745_
timestamp 0
transform -1 0 9490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1746_
timestamp 0
transform 1 0 11350 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1747_
timestamp 0
transform 1 0 10830 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1748_
timestamp 0
transform 1 0 7550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1749_
timestamp 0
transform 1 0 7970 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1750_
timestamp 0
transform -1 0 8090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1751_
timestamp 0
transform 1 0 7490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1752_
timestamp 0
transform -1 0 8910 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1753_
timestamp 0
transform 1 0 9770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1754_
timestamp 0
transform -1 0 8310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1755_
timestamp 0
transform -1 0 8890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__1756_
timestamp 0
transform -1 0 11230 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1757_
timestamp 0
transform 1 0 11090 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1758_
timestamp 0
transform -1 0 9150 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1759_
timestamp 0
transform -1 0 7390 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__1760_
timestamp 0
transform 1 0 8890 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__1761_
timestamp 0
transform -1 0 9610 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1762_
timestamp 0
transform 1 0 10630 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1763_
timestamp 0
transform -1 0 9070 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1764_
timestamp 0
transform 1 0 11330 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1765_
timestamp 0
transform 1 0 8150 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1766_
timestamp 0
transform 1 0 8530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1767_
timestamp 0
transform 1 0 9230 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__1768_
timestamp 0
transform 1 0 8090 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__1769_
timestamp 0
transform 1 0 8610 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__1770_
timestamp 0
transform 1 0 9050 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__1771_
timestamp 0
transform 1 0 9010 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__1772_
timestamp 0
transform 1 0 8730 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__1773_
timestamp 0
transform 1 0 10810 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1774_
timestamp 0
transform 1 0 10810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1775_
timestamp 0
transform 1 0 10050 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1776_
timestamp 0
transform -1 0 8050 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1777_
timestamp 0
transform 1 0 8090 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1778_
timestamp 0
transform -1 0 7570 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1779_
timestamp 0
transform 1 0 5710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1780_
timestamp 0
transform -1 0 4110 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1781_
timestamp 0
transform -1 0 10830 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1782_
timestamp 0
transform 1 0 8310 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1783_
timestamp 0
transform 1 0 10550 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1784_
timestamp 0
transform -1 0 10030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1785_
timestamp 0
transform -1 0 9790 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1786_
timestamp 0
transform 1 0 10210 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1787_
timestamp 0
transform -1 0 9150 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1788_
timestamp 0
transform -1 0 8570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1789_
timestamp 0
transform 1 0 10010 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1790_
timestamp 0
transform -1 0 10070 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1791_
timestamp 0
transform -1 0 10150 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1792_
timestamp 0
transform -1 0 9690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1793_
timestamp 0
transform -1 0 9430 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1794_
timestamp 0
transform 1 0 9150 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1795_
timestamp 0
transform -1 0 8350 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1796_
timestamp 0
transform -1 0 8290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1797_
timestamp 0
transform 1 0 7130 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1798_
timestamp 0
transform 1 0 7390 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1799_
timestamp 0
transform -1 0 9410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1800_
timestamp 0
transform 1 0 11290 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1801_
timestamp 0
transform 1 0 9310 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1802_
timestamp 0
transform -1 0 8970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1803_
timestamp 0
transform 1 0 10570 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1804_
timestamp 0
transform -1 0 8590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1805_
timestamp 0
transform -1 0 8690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1806_
timestamp 0
transform 1 0 7630 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1807_
timestamp 0
transform -1 0 8090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1808_
timestamp 0
transform -1 0 8410 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1809_
timestamp 0
transform 1 0 8630 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1810_
timestamp 0
transform 1 0 8030 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1811_
timestamp 0
transform -1 0 7770 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1812_
timestamp 0
transform -1 0 8410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1813_
timestamp 0
transform -1 0 8130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1814_
timestamp 0
transform -1 0 7870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1815_
timestamp 0
transform 1 0 7890 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1816_
timestamp 0
transform -1 0 3890 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1817_
timestamp 0
transform 1 0 1370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1818_
timestamp 0
transform -1 0 6190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1819_
timestamp 0
transform -1 0 950 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1820_
timestamp 0
transform 1 0 390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1821_
timestamp 0
transform 1 0 910 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1822_
timestamp 0
transform -1 0 370 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1823_
timestamp 0
transform 1 0 1730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1824_
timestamp 0
transform 1 0 1310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1825_
timestamp 0
transform -1 0 1150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1826_
timestamp 0
transform -1 0 410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1827_
timestamp 0
transform 1 0 910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1828_
timestamp 0
transform -1 0 1510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1829_
timestamp 0
transform -1 0 650 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1830_
timestamp 0
transform -1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1831_
timestamp 0
transform 1 0 2030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1832_
timestamp 0
transform -1 0 8030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1833_
timestamp 0
transform 1 0 9670 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1834_
timestamp 0
transform 1 0 9250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1835_
timestamp 0
transform -1 0 7770 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1836_
timestamp 0
transform -1 0 6430 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1837_
timestamp 0
transform -1 0 7770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1838_
timestamp 0
transform -1 0 7210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1839_
timestamp 0
transform -1 0 6190 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1840_
timestamp 0
transform 1 0 8570 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1841_
timestamp 0
transform -1 0 8190 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1842_
timestamp 0
transform -1 0 6950 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1843_
timestamp 0
transform -1 0 6670 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1844_
timestamp 0
transform 1 0 9090 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1845_
timestamp 0
transform 1 0 9630 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1846_
timestamp 0
transform -1 0 9230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1847_
timestamp 0
transform -1 0 8390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1848_
timestamp 0
transform 1 0 11230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1849_
timestamp 0
transform -1 0 11550 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1850_
timestamp 0
transform -1 0 11010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1851_
timestamp 0
transform 1 0 10370 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1852_
timestamp 0
transform -1 0 10430 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1853_
timestamp 0
transform -1 0 10450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1854_
timestamp 0
transform -1 0 7430 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1855_
timestamp 0
transform 1 0 7410 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1856_
timestamp 0
transform 1 0 7690 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1857_
timestamp 0
transform -1 0 8830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__1858_
timestamp 0
transform -1 0 9370 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1859_
timestamp 0
transform -1 0 8830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1860_
timestamp 0
transform 1 0 9090 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1861_
timestamp 0
transform 1 0 6830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1862_
timestamp 0
transform -1 0 8330 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__1863_
timestamp 0
transform 1 0 7690 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1864_
timestamp 0
transform -1 0 6330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1865_
timestamp 0
transform -1 0 7770 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__1866_
timestamp 0
transform -1 0 7230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1867_
timestamp 0
transform -1 0 8010 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1868_
timestamp 0
transform 1 0 7730 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1869_
timestamp 0
transform -1 0 6030 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__1870_
timestamp 0
transform 1 0 9370 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1871_
timestamp 0
transform 1 0 8850 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1872_
timestamp 0
transform -1 0 8590 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1873_
timestamp 0
transform -1 0 7790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1874_
timestamp 0
transform -1 0 7510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1875_
timestamp 0
transform -1 0 8310 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1876_
timestamp 0
transform -1 0 6950 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1877_
timestamp 0
transform -1 0 5790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__1878_
timestamp 0
transform 1 0 6670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1879_
timestamp 0
transform -1 0 7470 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1880_
timestamp 0
transform 1 0 5990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__1881_
timestamp 0
transform 1 0 5990 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__1882_
timestamp 0
transform -1 0 4950 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__1883_
timestamp 0
transform -1 0 7850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1884_
timestamp 0
transform -1 0 8090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1885_
timestamp 0
transform -1 0 8650 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1886_
timestamp 0
transform 1 0 8490 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1887_
timestamp 0
transform -1 0 8470 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1888_
timestamp 0
transform 1 0 11610 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1889_
timestamp 0
transform -1 0 8470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1890_
timestamp 0
transform 1 0 9730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1891_
timestamp 0
transform 1 0 8890 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1892_
timestamp 0
transform -1 0 8610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1893_
timestamp 0
transform 1 0 12130 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1894_
timestamp 0
transform 1 0 12110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1895_
timestamp 0
transform 1 0 12130 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1896_
timestamp 0
transform -1 0 10750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1897_
timestamp 0
transform -1 0 9150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1898_
timestamp 0
transform 1 0 9030 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1899_
timestamp 0
transform 1 0 7470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1900_
timestamp 0
transform 1 0 9670 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1901_
timestamp 0
transform 1 0 8010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1902_
timestamp 0
transform -1 0 8230 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1903_
timestamp 0
transform 1 0 7950 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1904_
timestamp 0
transform 1 0 11870 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1905_
timestamp 0
transform 1 0 11630 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1906_
timestamp 0
transform -1 0 6510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1907_
timestamp 0
transform -1 0 7050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1908_
timestamp 0
transform -1 0 6970 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1909_
timestamp 0
transform -1 0 6730 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1910_
timestamp 0
transform -1 0 6230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1911_
timestamp 0
transform 1 0 6810 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1912_
timestamp 0
transform 1 0 6270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1913_
timestamp 0
transform 1 0 6210 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1914_
timestamp 0
transform 1 0 5710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1915_
timestamp 0
transform 1 0 5230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1916_
timestamp 0
transform 1 0 5230 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__1917_
timestamp 0
transform -1 0 3730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__1918_
timestamp 0
transform 1 0 3610 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__1919_
timestamp 0
transform -1 0 3890 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__1920_
timestamp 0
transform -1 0 3610 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__1921_
timestamp 0
transform -1 0 1730 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__1922_
timestamp 0
transform 1 0 7530 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1923_
timestamp 0
transform 1 0 7790 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1924_
timestamp 0
transform -1 0 6390 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1925_
timestamp 0
transform -1 0 4630 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1926_
timestamp 0
transform -1 0 3990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1927_
timestamp 0
transform 1 0 2030 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__1928_
timestamp 0
transform -1 0 3190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__1929_
timestamp 0
transform 1 0 4570 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__1930_
timestamp 0
transform 1 0 3130 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__1931_
timestamp 0
transform -1 0 2910 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__1932_
timestamp 0
transform -1 0 1510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1933_
timestamp 0
transform -1 0 8470 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1934_
timestamp 0
transform 1 0 3870 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1935_
timestamp 0
transform -1 0 3890 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1936_
timestamp 0
transform -1 0 2570 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1937_
timestamp 0
transform -1 0 1230 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1938_
timestamp 0
transform -1 0 3590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1939_
timestamp 0
transform -1 0 4150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1940_
timestamp 0
transform -1 0 3370 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1941_
timestamp 0
transform -1 0 3310 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1942_
timestamp 0
transform -1 0 1810 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__1943_
timestamp 0
transform -1 0 3610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1944_
timestamp 0
transform -1 0 3710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1945_
timestamp 0
transform -1 0 2970 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1946_
timestamp 0
transform -1 0 1530 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__1947_
timestamp 0
transform -1 0 4950 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__1948_
timestamp 0
transform 1 0 5150 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__1949_
timestamp 0
transform 1 0 5210 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__1950_
timestamp 0
transform -1 0 4950 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__1951_
timestamp 0
transform -1 0 1990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1952_
timestamp 0
transform 1 0 4110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1953_
timestamp 0
transform 1 0 4050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1954_
timestamp 0
transform 1 0 4190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1955_
timestamp 0
transform -1 0 1710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1956_
timestamp 0
transform -1 0 4330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__1957_
timestamp 0
transform 1 0 4910 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__1958_
timestamp 0
transform -1 0 5190 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__1959_
timestamp 0
transform -1 0 4170 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__1960_
timestamp 0
transform -1 0 2330 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1961_
timestamp 0
transform 1 0 4150 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1962_
timestamp 0
transform 1 0 3910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1963_
timestamp 0
transform 1 0 3690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1964_
timestamp 0
transform 1 0 2030 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1965_
timestamp 0
transform 1 0 6410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__1966_
timestamp 0
transform 1 0 6350 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1967_
timestamp 0
transform 1 0 7190 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1968_
timestamp 0
transform 1 0 6650 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1969_
timestamp 0
transform -1 0 3310 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__1970_
timestamp 0
transform 1 0 2850 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1971_
timestamp 0
transform -1 0 4730 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1972_
timestamp 0
transform 1 0 3590 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1973_
timestamp 0
transform -1 0 3610 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1974_
timestamp 0
transform -1 0 3110 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__1975_
timestamp 0
transform 1 0 3010 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__1976_
timestamp 0
transform -1 0 3110 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__1977_
timestamp 0
transform 1 0 4390 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__1978_
timestamp 0
transform 1 0 3090 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__1979_
timestamp 0
transform -1 0 2830 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__1980_
timestamp 0
transform -1 0 2350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1981_
timestamp 0
transform 1 0 5970 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1982_
timestamp 0
transform 1 0 6090 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1983_
timestamp 0
transform 1 0 6290 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1984_
timestamp 0
transform 1 0 5290 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1985_
timestamp 0
transform -1 0 4790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1986_
timestamp 0
transform 1 0 2570 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__1987_
timestamp 0
transform -1 0 7290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1988_
timestamp 0
transform 1 0 7590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1989_
timestamp 0
transform 1 0 7650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1990_
timestamp 0
transform -1 0 7450 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1991_
timestamp 0
transform -1 0 7730 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1992_
timestamp 0
transform 1 0 10470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1993_
timestamp 0
transform 1 0 9590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__1994_
timestamp 0
transform -1 0 6270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__1995_
timestamp 0
transform 1 0 6650 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1996_
timestamp 0
transform -1 0 6790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1997_
timestamp 0
transform 1 0 6490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1998_
timestamp 0
transform 1 0 6490 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__1999_
timestamp 0
transform 1 0 7550 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2000_
timestamp 0
transform 1 0 6470 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2001_
timestamp 0
transform 1 0 6710 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2002_
timestamp 0
transform 1 0 6670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2003_
timestamp 0
transform 1 0 9550 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2004_
timestamp 0
transform 1 0 7490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2005_
timestamp 0
transform -1 0 7290 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2006_
timestamp 0
transform 1 0 6770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2007_
timestamp 0
transform 1 0 6610 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2008_
timestamp 0
transform -1 0 6250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2009_
timestamp 0
transform 1 0 6850 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2010_
timestamp 0
transform -1 0 7070 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2011_
timestamp 0
transform 1 0 7310 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2012_
timestamp 0
transform -1 0 9450 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2013_
timestamp 0
transform 1 0 10590 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2014_
timestamp 0
transform -1 0 10850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2015_
timestamp 0
transform -1 0 6290 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2016_
timestamp 0
transform -1 0 7330 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2017_
timestamp 0
transform -1 0 7110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2018_
timestamp 0
transform 1 0 7350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2019_
timestamp 0
transform 1 0 9430 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2020_
timestamp 0
transform -1 0 10330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2021_
timestamp 0
transform -1 0 7370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2022_
timestamp 0
transform 1 0 7610 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2023_
timestamp 0
transform -1 0 7910 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2024_
timestamp 0
transform 1 0 6130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2025_
timestamp 0
transform -1 0 6010 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2026_
timestamp 0
transform 1 0 9710 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2027_
timestamp 0
transform 1 0 10250 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2028_
timestamp 0
transform -1 0 10250 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2029_
timestamp 0
transform -1 0 11130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2030_
timestamp 0
transform 1 0 10750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2031_
timestamp 0
transform -1 0 11050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2032_
timestamp 0
transform 1 0 8970 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2033_
timestamp 0
transform 1 0 8430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2034_
timestamp 0
transform 1 0 8670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2035_
timestamp 0
transform 1 0 8630 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2036_
timestamp 0
transform 1 0 11590 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2037_
timestamp 0
transform 1 0 11790 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2038_
timestamp 0
transform -1 0 7630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2039_
timestamp 0
transform -1 0 6710 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2040_
timestamp 0
transform 1 0 10970 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2041_
timestamp 0
transform 1 0 11050 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2042_
timestamp 0
transform -1 0 10130 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2043_
timestamp 0
transform -1 0 10510 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2044_
timestamp 0
transform -1 0 11030 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2045_
timestamp 0
transform -1 0 11370 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2046_
timestamp 0
transform 1 0 8850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2047_
timestamp 0
transform -1 0 9410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2048_
timestamp 0
transform 1 0 9210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2049_
timestamp 0
transform 1 0 9350 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2050_
timestamp 0
transform 1 0 9110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2051_
timestamp 0
transform 1 0 8810 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2052_
timestamp 0
transform 1 0 9090 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2053_
timestamp 0
transform -1 0 9650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2054_
timestamp 0
transform 1 0 9870 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2055_
timestamp 0
transform -1 0 6510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2056_
timestamp 0
transform -1 0 6090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2057_
timestamp 0
transform 1 0 10290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2058_
timestamp 0
transform -1 0 10030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2059_
timestamp 0
transform -1 0 10170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2060_
timestamp 0
transform -1 0 9930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2061_
timestamp 0
transform 1 0 10110 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2062_
timestamp 0
transform -1 0 9190 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2063_
timestamp 0
transform 1 0 8270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2064_
timestamp 0
transform -1 0 7950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2065_
timestamp 0
transform -1 0 8770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2066_
timestamp 0
transform 1 0 8750 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2067_
timestamp 0
transform -1 0 8010 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2068_
timestamp 0
transform -1 0 8290 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2069_
timestamp 0
transform 1 0 8010 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2070_
timestamp 0
transform -1 0 8310 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2071_
timestamp 0
transform -1 0 8590 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2072_
timestamp 0
transform 1 0 8810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2073_
timestamp 0
transform 1 0 9070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2074_
timestamp 0
transform 1 0 9290 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2075_
timestamp 0
transform -1 0 9590 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2076_
timestamp 0
transform 1 0 11250 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2077_
timestamp 0
transform -1 0 11310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2078_
timestamp 0
transform -1 0 11110 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2079_
timestamp 0
transform 1 0 11250 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2080_
timestamp 0
transform -1 0 11090 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2081_
timestamp 0
transform 1 0 11090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2082_
timestamp 0
transform 1 0 10350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2083_
timestamp 0
transform 1 0 9610 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2084_
timestamp 0
transform 1 0 11630 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2085_
timestamp 0
transform 1 0 11050 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2086_
timestamp 0
transform 1 0 11550 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2087_
timestamp 0
transform 1 0 11570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2088_
timestamp 0
transform -1 0 12130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2089_
timestamp 0
transform 1 0 11850 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2090_
timestamp 0
transform 1 0 12030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2091_
timestamp 0
transform 1 0 9930 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2092_
timestamp 0
transform 1 0 10550 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2093_
timestamp 0
transform -1 0 11110 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2094_
timestamp 0
transform 1 0 11350 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2095_
timestamp 0
transform -1 0 11010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2096_
timestamp 0
transform 1 0 11530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2097_
timestamp 0
transform -1 0 11870 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2098_
timestamp 0
transform -1 0 12050 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2099_
timestamp 0
transform -1 0 11350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2100_
timestamp 0
transform 1 0 11310 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2101_
timestamp 0
transform -1 0 11270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2102_
timestamp 0
transform -1 0 11650 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2103_
timestamp 0
transform 1 0 12130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2104_
timestamp 0
transform 1 0 12130 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2105_
timestamp 0
transform -1 0 11590 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2106_
timestamp 0
transform -1 0 11570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2107_
timestamp 0
transform -1 0 12130 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2108_
timestamp 0
transform 1 0 8870 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2109_
timestamp 0
transform 1 0 12130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2110_
timestamp 0
transform -1 0 12150 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2111_
timestamp 0
transform -1 0 12150 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2112_
timestamp 0
transform -1 0 12050 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2113_
timestamp 0
transform 1 0 11810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2114_
timestamp 0
transform 1 0 10590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2115_
timestamp 0
transform -1 0 9330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2116_
timestamp 0
transform -1 0 10210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2117_
timestamp 0
transform -1 0 10810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2118_
timestamp 0
transform -1 0 10770 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2119_
timestamp 0
transform 1 0 10670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2120_
timestamp 0
transform 1 0 10710 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2121_
timestamp 0
transform -1 0 10450 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2122_
timestamp 0
transform 1 0 10650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2123_
timestamp 0
transform -1 0 8150 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2124_
timestamp 0
transform -1 0 7850 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2125_
timestamp 0
transform -1 0 10210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2126_
timestamp 0
transform 1 0 10610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2127_
timestamp 0
transform -1 0 7030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2128_
timestamp 0
transform -1 0 9170 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2129_
timestamp 0
transform 1 0 7290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2130_
timestamp 0
transform -1 0 10910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2131_
timestamp 0
transform -1 0 7950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2132_
timestamp 0
transform 1 0 6730 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2133_
timestamp 0
transform -1 0 7030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2134_
timestamp 0
transform -1 0 7290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2135_
timestamp 0
transform -1 0 11170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2136_
timestamp 0
transform -1 0 11330 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2137_
timestamp 0
transform 1 0 11310 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2138_
timestamp 0
transform 1 0 11390 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2139_
timestamp 0
transform -1 0 11310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2140_
timestamp 0
transform -1 0 11030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2141_
timestamp 0
transform 1 0 9950 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2142_
timestamp 0
transform 1 0 10750 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2143_
timestamp 0
transform -1 0 10490 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2144_
timestamp 0
transform -1 0 11050 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2145_
timestamp 0
transform -1 0 5050 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2146_
timestamp 0
transform 1 0 9770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2147_
timestamp 0
transform 1 0 10330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2148_
timestamp 0
transform -1 0 6270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2149_
timestamp 0
transform 1 0 10050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2150_
timestamp 0
transform 1 0 8830 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2151_
timestamp 0
transform 1 0 7450 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2152_
timestamp 0
transform 1 0 8530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2153_
timestamp 0
transform 1 0 8790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2154_
timestamp 0
transform 1 0 9070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2155_
timestamp 0
transform -1 0 10150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2156_
timestamp 0
transform -1 0 10930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2157_
timestamp 0
transform 1 0 11170 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2158_
timestamp 0
transform -1 0 11750 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2159_
timestamp 0
transform -1 0 11870 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2160_
timestamp 0
transform -1 0 11410 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2161_
timestamp 0
transform 1 0 8150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2162_
timestamp 0
transform 1 0 8910 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2163_
timestamp 0
transform -1 0 10010 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2164_
timestamp 0
transform 1 0 9770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2165_
timestamp 0
transform 1 0 11010 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2166_
timestamp 0
transform 1 0 10830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2167_
timestamp 0
transform 1 0 9210 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2168_
timestamp 0
transform 1 0 10030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2169_
timestamp 0
transform -1 0 8770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2170_
timestamp 0
transform -1 0 9190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2171_
timestamp 0
transform 1 0 10330 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2172_
timestamp 0
transform 1 0 9750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2173_
timestamp 0
transform 1 0 9870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2174_
timestamp 0
transform -1 0 9510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2175_
timestamp 0
transform 1 0 9590 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2176_
timestamp 0
transform -1 0 9710 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2177_
timestamp 0
transform -1 0 9410 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2178_
timestamp 0
transform -1 0 11010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2179_
timestamp 0
transform 1 0 9490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2180_
timestamp 0
transform 1 0 11850 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2181_
timestamp 0
transform 1 0 11830 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2182_
timestamp 0
transform 1 0 11910 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2183_
timestamp 0
transform -1 0 11290 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2184_
timestamp 0
transform 1 0 11030 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2185_
timestamp 0
transform -1 0 10270 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2186_
timestamp 0
transform 1 0 10210 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2187_
timestamp 0
transform -1 0 10610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2188_
timestamp 0
transform 1 0 11570 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2189_
timestamp 0
transform 1 0 9950 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2190_
timestamp 0
transform 1 0 10510 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2191_
timestamp 0
transform 1 0 11130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2192_
timestamp 0
transform 1 0 11070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2193_
timestamp 0
transform -1 0 11010 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2194_
timestamp 0
transform -1 0 10570 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2195_
timestamp 0
transform -1 0 9450 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2196_
timestamp 0
transform -1 0 11090 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2197_
timestamp 0
transform 1 0 11350 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2198_
timestamp 0
transform -1 0 9890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2199_
timestamp 0
transform -1 0 9950 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2200_
timestamp 0
transform -1 0 5810 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2201_
timestamp 0
transform 1 0 6330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2202_
timestamp 0
transform 1 0 6070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2203_
timestamp 0
transform 1 0 6070 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2204_
timestamp 0
transform 1 0 6810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2205_
timestamp 0
transform 1 0 7110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2206_
timestamp 0
transform 1 0 9450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2207_
timestamp 0
transform -1 0 9950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2208_
timestamp 0
transform -1 0 9370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2209_
timestamp 0
transform 1 0 10410 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2210_
timestamp 0
transform 1 0 10410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2211_
timestamp 0
transform 1 0 11250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2212_
timestamp 0
transform -1 0 11610 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2213_
timestamp 0
transform -1 0 11650 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2214_
timestamp 0
transform 1 0 11610 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2215_
timestamp 0
transform 1 0 11710 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2216_
timestamp 0
transform 1 0 12090 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2217_
timestamp 0
transform 1 0 11370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2218_
timestamp 0
transform 1 0 9650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2219_
timestamp 0
transform -1 0 9890 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2220_
timestamp 0
transform -1 0 9930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2221_
timestamp 0
transform -1 0 11870 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2222_
timestamp 0
transform 1 0 11810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2223_
timestamp 0
transform -1 0 11850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2224_
timestamp 0
transform 1 0 11830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2225_
timestamp 0
transform 1 0 10930 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2226_
timestamp 0
transform 1 0 11890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2227_
timestamp 0
transform 1 0 11610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2228_
timestamp 0
transform -1 0 11470 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2229_
timestamp 0
transform -1 0 10550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2230_
timestamp 0
transform -1 0 10270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2231_
timestamp 0
transform -1 0 8470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2232_
timestamp 0
transform 1 0 8710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2233_
timestamp 0
transform 1 0 9490 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2234_
timestamp 0
transform -1 0 9750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2235_
timestamp 0
transform -1 0 9870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2236_
timestamp 0
transform 1 0 7170 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2237_
timestamp 0
transform -1 0 6650 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2238_
timestamp 0
transform -1 0 6930 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2239_
timestamp 0
transform -1 0 8950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2240_
timestamp 0
transform -1 0 8670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2241_
timestamp 0
transform -1 0 8310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2242_
timestamp 0
transform -1 0 7490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2243_
timestamp 0
transform 1 0 7750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2244_
timestamp 0
transform 1 0 8030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2245_
timestamp 0
transform -1 0 7730 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2246_
timestamp 0
transform 1 0 9110 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2247_
timestamp 0
transform -1 0 12110 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2248_
timestamp 0
transform 1 0 11310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2249_
timestamp 0
transform -1 0 9470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2250_
timestamp 0
transform 1 0 10990 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2251_
timestamp 0
transform 1 0 10550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2252_
timestamp 0
transform 1 0 11290 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2253_
timestamp 0
transform -1 0 11890 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2254_
timestamp 0
transform 1 0 12130 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2255_
timestamp 0
transform -1 0 10490 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2256_
timestamp 0
transform -1 0 10770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2257_
timestamp 0
transform 1 0 11010 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2258_
timestamp 0
transform 1 0 12170 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2259_
timestamp 0
transform -1 0 11850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2260_
timestamp 0
transform 1 0 10030 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2261_
timestamp 0
transform 1 0 10290 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2262_
timestamp 0
transform -1 0 10810 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2263_
timestamp 0
transform 1 0 11290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2264_
timestamp 0
transform 1 0 12110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2265_
timestamp 0
transform -1 0 11370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2266_
timestamp 0
transform -1 0 10730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2267_
timestamp 0
transform 1 0 11950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2268_
timestamp 0
transform 1 0 12110 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2269_
timestamp 0
transform -1 0 11890 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2270_
timestamp 0
transform 1 0 11310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2271_
timestamp 0
transform -1 0 11610 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2272_
timestamp 0
transform 1 0 11870 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2273_
timestamp 0
transform -1 0 12130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2274_
timestamp 0
transform 1 0 10050 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2275_
timestamp 0
transform -1 0 8210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2276_
timestamp 0
transform 1 0 8870 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2277_
timestamp 0
transform 1 0 9150 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2278_
timestamp 0
transform -1 0 9230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2279_
timestamp 0
transform 1 0 9030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2280_
timestamp 0
transform 1 0 10190 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2281_
timestamp 0
transform 1 0 12070 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2282_
timestamp 0
transform 1 0 12130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2283_
timestamp 0
transform -1 0 11010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2284_
timestamp 0
transform 1 0 12090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2285_
timestamp 0
transform 1 0 12090 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2286_
timestamp 0
transform -1 0 11870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2287_
timestamp 0
transform 1 0 11810 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2288_
timestamp 0
transform -1 0 10970 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2289_
timestamp 0
transform -1 0 10750 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2290_
timestamp 0
transform -1 0 10930 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2291_
timestamp 0
transform 1 0 11290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2292_
timestamp 0
transform 1 0 10430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2293_
timestamp 0
transform 1 0 10710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2294_
timestamp 0
transform 1 0 11030 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2295_
timestamp 0
transform 1 0 10910 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2296_
timestamp 0
transform 1 0 11170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2297_
timestamp 0
transform 1 0 11830 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2298_
timestamp 0
transform -1 0 11930 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2299_
timestamp 0
transform -1 0 10490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2300_
timestamp 0
transform 1 0 10190 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2301_
timestamp 0
transform 1 0 11810 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2302_
timestamp 0
transform 1 0 11750 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2303_
timestamp 0
transform -1 0 11730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2304_
timestamp 0
transform 1 0 11870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2305_
timestamp 0
transform 1 0 10750 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2306_
timestamp 0
transform -1 0 11610 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2307_
timestamp 0
transform 1 0 11310 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2308_
timestamp 0
transform 1 0 12090 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2309_
timestamp 0
transform -1 0 11650 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2310_
timestamp 0
transform -1 0 11590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2311_
timestamp 0
transform 1 0 11570 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2312_
timestamp 0
transform 1 0 11630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2313_
timestamp 0
transform 1 0 11910 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2314_
timestamp 0
transform -1 0 11230 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2315_
timestamp 0
transform 1 0 12090 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2316_
timestamp 0
transform 1 0 11490 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2317_
timestamp 0
transform -1 0 11990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2318_
timestamp 0
transform 1 0 11530 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2319_
timestamp 0
transform 1 0 11170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2320_
timestamp 0
transform 1 0 11590 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2321_
timestamp 0
transform 1 0 11450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2322_
timestamp 0
transform -1 0 11310 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2323_
timestamp 0
transform -1 0 11550 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2324_
timestamp 0
transform 1 0 11790 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2325_
timestamp 0
transform -1 0 12170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2326_
timestamp 0
transform 1 0 12090 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2327_
timestamp 0
transform 1 0 11450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2328_
timestamp 0
transform 1 0 11030 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2329_
timestamp 0
transform 1 0 8550 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2330_
timestamp 0
transform -1 0 10230 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2331_
timestamp 0
transform -1 0 9670 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2332_
timestamp 0
transform -1 0 11890 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2333_
timestamp 0
transform -1 0 10770 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2334_
timestamp 0
transform 1 0 10490 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2335_
timestamp 0
transform 1 0 10470 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2336_
timestamp 0
transform 1 0 10650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2337_
timestamp 0
transform -1 0 10770 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2338_
timestamp 0
transform -1 0 10690 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2339_
timestamp 0
transform -1 0 9610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2340_
timestamp 0
transform -1 0 9890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2341_
timestamp 0
transform 1 0 9590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2342_
timestamp 0
transform -1 0 10470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2343_
timestamp 0
transform -1 0 10410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2344_
timestamp 0
transform -1 0 10650 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2345_
timestamp 0
transform 1 0 11770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2346_
timestamp 0
transform 1 0 11510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2347_
timestamp 0
transform -1 0 8850 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2348_
timestamp 0
transform -1 0 9950 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2349_
timestamp 0
transform -1 0 11610 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2350_
timestamp 0
transform -1 0 11330 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2351_
timestamp 0
transform -1 0 10390 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2352_
timestamp 0
transform -1 0 10150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2353_
timestamp 0
transform -1 0 9450 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2354_
timestamp 0
transform 1 0 7850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2355_
timestamp 0
transform -1 0 6930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2356_
timestamp 0
transform -1 0 6870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2357_
timestamp 0
transform -1 0 7530 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2358_
timestamp 0
transform -1 0 7110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2359_
timestamp 0
transform 1 0 7330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2360_
timestamp 0
transform -1 0 8010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2361_
timestamp 0
transform -1 0 7070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2362_
timestamp 0
transform 1 0 8790 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2363_
timestamp 0
transform -1 0 7470 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2364_
timestamp 0
transform 1 0 7210 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2365_
timestamp 0
transform 1 0 6930 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2366_
timestamp 0
transform 1 0 6410 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2367_
timestamp 0
transform -1 0 7250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2368_
timestamp 0
transform 1 0 6650 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2369_
timestamp 0
transform 1 0 7030 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2370_
timestamp 0
transform -1 0 7290 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2371_
timestamp 0
transform 1 0 7230 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2372_
timestamp 0
transform -1 0 6810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2373_
timestamp 0
transform 1 0 6750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2374_
timestamp 0
transform 1 0 8250 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2375_
timestamp 0
transform 1 0 8310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2376_
timestamp 0
transform -1 0 6750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2377_
timestamp 0
transform 1 0 5450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2378_
timestamp 0
transform -1 0 3770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2379_
timestamp 0
transform -1 0 8030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2380_
timestamp 0
transform -1 0 5670 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2381_
timestamp 0
transform -1 0 5950 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2382_
timestamp 0
transform -1 0 5810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2383_
timestamp 0
transform 1 0 4730 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2384_
timestamp 0
transform 1 0 4650 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2385_
timestamp 0
transform 1 0 4890 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2386_
timestamp 0
transform 1 0 5170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2387_
timestamp 0
transform 1 0 1690 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2388_
timestamp 0
transform 1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2389_
timestamp 0
transform 1 0 5210 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2390_
timestamp 0
transform 1 0 2490 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2391_
timestamp 0
transform -1 0 2290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2392_
timestamp 0
transform -1 0 2010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2393_
timestamp 0
transform -1 0 2570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2394_
timestamp 0
transform -1 0 2990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2395_
timestamp 0
transform 1 0 4390 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2396_
timestamp 0
transform 1 0 3030 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2397_
timestamp 0
transform -1 0 3110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2398_
timestamp 0
transform -1 0 2830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2399_
timestamp 0
transform 1 0 1930 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2400_
timestamp 0
transform -1 0 1370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2401_
timestamp 0
transform -1 0 2850 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2402_
timestamp 0
transform 1 0 2590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2403_
timestamp 0
transform -1 0 2230 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2404_
timestamp 0
transform -1 0 1670 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2405_
timestamp 0
transform -1 0 1530 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2406_
timestamp 0
transform 1 0 5910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2407_
timestamp 0
transform -1 0 4270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2408_
timestamp 0
transform -1 0 5630 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2409_
timestamp 0
transform -1 0 6450 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2410_
timestamp 0
transform -1 0 4230 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2411_
timestamp 0
transform -1 0 3990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2412_
timestamp 0
transform -1 0 1250 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2413_
timestamp 0
transform -1 0 4530 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2414_
timestamp 0
transform 1 0 3050 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2415_
timestamp 0
transform -1 0 2790 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2416_
timestamp 0
transform 1 0 1750 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2417_
timestamp 0
transform -1 0 2250 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2418_
timestamp 0
transform -1 0 2130 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2419_
timestamp 0
transform -1 0 3450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2420_
timestamp 0
transform 1 0 2870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2421_
timestamp 0
transform -1 0 2790 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2422_
timestamp 0
transform -1 0 1970 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2423_
timestamp 0
transform -1 0 3670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2424_
timestamp 0
transform -1 0 3510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2425_
timestamp 0
transform -1 0 3390 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2426_
timestamp 0
transform 1 0 3150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2427_
timestamp 0
transform 1 0 3310 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2428_
timestamp 0
transform -1 0 3390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2429_
timestamp 0
transform -1 0 5110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2430_
timestamp 0
transform -1 0 7810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2431_
timestamp 0
transform -1 0 5370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2432_
timestamp 0
transform -1 0 9490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2433_
timestamp 0
transform 1 0 11590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2434_
timestamp 0
transform 1 0 10770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2435_
timestamp 0
transform -1 0 7250 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2436_
timestamp 0
transform -1 0 6930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2437_
timestamp 0
transform -1 0 9610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2438_
timestamp 0
transform -1 0 9350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2439_
timestamp 0
transform -1 0 6130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2440_
timestamp 0
transform 1 0 7750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2441_
timestamp 0
transform -1 0 7590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2442_
timestamp 0
transform 1 0 10290 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2443_
timestamp 0
transform -1 0 7190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2444_
timestamp 0
transform -1 0 7190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2445_
timestamp 0
transform 1 0 5290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2446_
timestamp 0
transform 1 0 6410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2447_
timestamp 0
transform -1 0 4790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2448_
timestamp 0
transform -1 0 6390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2449_
timestamp 0
transform -1 0 7010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2450_
timestamp 0
transform 1 0 4150 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2451_
timestamp 0
transform -1 0 4030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2452_
timestamp 0
transform 1 0 4670 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2453_
timestamp 0
transform 1 0 8530 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2454_
timestamp 0
transform 1 0 4410 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2455_
timestamp 0
transform 1 0 4410 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2456_
timestamp 0
transform -1 0 4270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2457_
timestamp 0
transform -1 0 4530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2458_
timestamp 0
transform -1 0 4890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2459_
timestamp 0
transform 1 0 5030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2460_
timestamp 0
transform 1 0 4910 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2461_
timestamp 0
transform 1 0 5190 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2462_
timestamp 0
transform 1 0 5330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2463_
timestamp 0
transform 1 0 6270 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2464_
timestamp 0
transform -1 0 3210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2465_
timestamp 0
transform -1 0 2930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2466_
timestamp 0
transform -1 0 2930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2467_
timestamp 0
transform 1 0 2070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2468_
timestamp 0
transform -1 0 1630 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2469_
timestamp 0
transform 1 0 590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2470_
timestamp 0
transform -1 0 2690 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2471_
timestamp 0
transform -1 0 2710 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2472_
timestamp 0
transform -1 0 2410 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2473_
timestamp 0
transform 1 0 1910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2474_
timestamp 0
transform -1 0 1430 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2475_
timestamp 0
transform -1 0 370 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2476_
timestamp 0
transform -1 0 3790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2477_
timestamp 0
transform -1 0 5030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2478_
timestamp 0
transform 1 0 3890 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2479_
timestamp 0
transform -1 0 3530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2480_
timestamp 0
transform 1 0 1770 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2481_
timestamp 0
transform -1 0 3330 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2482_
timestamp 0
transform 1 0 3610 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2483_
timestamp 0
transform 1 0 3030 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2484_
timestamp 0
transform 1 0 2750 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2485_
timestamp 0
transform -1 0 370 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2486_
timestamp 0
transform -1 0 2650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2487_
timestamp 0
transform 1 0 2370 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2488_
timestamp 0
transform -1 0 2370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2489_
timestamp 0
transform -1 0 1810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2490_
timestamp 0
transform -1 0 1370 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2491_
timestamp 0
transform -1 0 370 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2492_
timestamp 0
transform 1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2493_
timestamp 0
transform 1 0 3590 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2494_
timestamp 0
transform 1 0 6170 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2495_
timestamp 0
transform 1 0 3830 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2496_
timestamp 0
transform 1 0 4130 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2497_
timestamp 0
transform -1 0 4050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2498_
timestamp 0
transform 1 0 3510 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2499_
timestamp 0
transform 1 0 3770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2500_
timestamp 0
transform -1 0 370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2501_
timestamp 0
transform -1 0 3370 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2502_
timestamp 0
transform -1 0 3010 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2503_
timestamp 0
transform -1 0 3490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__2504_
timestamp 0
transform -1 0 3250 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__2505_
timestamp 0
transform 1 0 2690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2506_
timestamp 0
transform -1 0 2510 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__2507_
timestamp 0
transform 1 0 630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2508_
timestamp 0
transform 1 0 3130 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2509_
timestamp 0
transform 1 0 2670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2510_
timestamp 0
transform -1 0 3230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2511_
timestamp 0
transform 1 0 3310 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__2512_
timestamp 0
transform 1 0 3150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2513_
timestamp 0
transform -1 0 2410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2514_
timestamp 0
transform 1 0 2110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2515_
timestamp 0
transform -1 0 2130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2516_
timestamp 0
transform -1 0 370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__2517_
timestamp 0
transform -1 0 2210 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2518_
timestamp 0
transform 1 0 5310 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2519_
timestamp 0
transform -1 0 5850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2520_
timestamp 0
transform -1 0 5950 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2521_
timestamp 0
transform 1 0 5650 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2522_
timestamp 0
transform -1 0 5650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2523_
timestamp 0
transform -1 0 5570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2524_
timestamp 0
transform -1 0 5510 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2525_
timestamp 0
transform -1 0 2730 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2526_
timestamp 0
transform 1 0 6130 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2527_
timestamp 0
transform 1 0 6530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2528_
timestamp 0
transform 1 0 6510 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2529_
timestamp 0
transform 1 0 6110 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2530_
timestamp 0
transform 1 0 5570 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2531_
timestamp 0
transform 1 0 2930 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2532_
timestamp 0
transform 1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2533_
timestamp 0
transform 1 0 5150 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2534_
timestamp 0
transform 1 0 4870 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2535_
timestamp 0
transform -1 0 4610 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2536_
timestamp 0
transform 1 0 3450 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2537_
timestamp 0
transform 1 0 2090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2538_
timestamp 0
transform 1 0 4490 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2539_
timestamp 0
transform 1 0 3870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2540_
timestamp 0
transform 1 0 4210 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2541_
timestamp 0
transform -1 0 4190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2542_
timestamp 0
transform -1 0 3710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2543_
timestamp 0
transform 1 0 3470 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2544_
timestamp 0
transform 1 0 4190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2545_
timestamp 0
transform 1 0 4450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2546_
timestamp 0
transform 1 0 4810 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2547_
timestamp 0
transform -1 0 4750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2548_
timestamp 0
transform -1 0 4470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2549_
timestamp 0
transform 1 0 4690 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2550_
timestamp 0
transform 1 0 4690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2551_
timestamp 0
transform 1 0 5210 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2552_
timestamp 0
transform 1 0 5450 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2553_
timestamp 0
transform 1 0 2350 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2554_
timestamp 0
transform 1 0 4490 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2555_
timestamp 0
transform -1 0 4670 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2556_
timestamp 0
transform -1 0 4910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2557_
timestamp 0
transform 1 0 4610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2558_
timestamp 0
transform 1 0 4690 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2559_
timestamp 0
transform 1 0 4410 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2560_
timestamp 0
transform 1 0 3910 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2561_
timestamp 0
transform 1 0 3610 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2562_
timestamp 0
transform 1 0 2230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2563_
timestamp 0
transform -1 0 4450 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2564_
timestamp 0
transform 1 0 4370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2565_
timestamp 0
transform -1 0 3850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2566_
timestamp 0
transform 1 0 2450 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2567_
timestamp 0
transform 1 0 3930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2568_
timestamp 0
transform -1 0 5730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2569_
timestamp 0
transform -1 0 5870 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2570_
timestamp 0
transform 1 0 5950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2571_
timestamp 0
transform 1 0 5950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2572_
timestamp 0
transform 1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2573_
timestamp 0
transform 1 0 5730 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2574_
timestamp 0
transform 1 0 5710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2575_
timestamp 0
transform -1 0 4750 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2576_
timestamp 0
transform -1 0 4230 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2577_
timestamp 0
transform -1 0 4490 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2578_
timestamp 0
transform 1 0 6990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2579_
timestamp 0
transform 1 0 7010 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2580_
timestamp 0
transform 1 0 8010 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2581_
timestamp 0
transform -1 0 8870 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2582_
timestamp 0
transform 1 0 6910 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2583_
timestamp 0
transform -1 0 6910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2584_
timestamp 0
transform 1 0 7330 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2585_
timestamp 0
transform 1 0 7370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2586_
timestamp 0
transform -1 0 8450 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2587_
timestamp 0
transform -1 0 6790 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2588_
timestamp 0
transform -1 0 5830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2589_
timestamp 0
transform 1 0 7450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2590_
timestamp 0
transform -1 0 6230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2591_
timestamp 0
transform 1 0 6470 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2592_
timestamp 0
transform -1 0 4450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2593_
timestamp 0
transform 1 0 4970 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2594_
timestamp 0
transform -1 0 8550 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2595_
timestamp 0
transform -1 0 5270 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2596_
timestamp 0
transform 1 0 5270 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2597_
timestamp 0
transform 1 0 5450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2598_
timestamp 0
transform -1 0 5190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2599_
timestamp 0
transform -1 0 4990 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2600_
timestamp 0
transform -1 0 4990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2601_
timestamp 0
transform -1 0 5250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2602_
timestamp 0
transform -1 0 8190 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2603_
timestamp 0
transform -1 0 6630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2604_
timestamp 0
transform -1 0 6390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2605_
timestamp 0
transform 1 0 6070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2606_
timestamp 0
transform -1 0 5570 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2607_
timestamp 0
transform 1 0 5730 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2608_
timestamp 0
transform 1 0 5550 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2609_
timestamp 0
transform -1 0 5530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2610_
timestamp 0
transform 1 0 4910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2611_
timestamp 0
transform -1 0 5170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2612_
timestamp 0
transform -1 0 5430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2613_
timestamp 0
transform -1 0 1250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2614_
timestamp 0
transform 1 0 2230 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2615_
timestamp 0
transform -1 0 2510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2616_
timestamp 0
transform -1 0 2490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2617_
timestamp 0
transform 1 0 1470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2618_
timestamp 0
transform 1 0 890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2619_
timestamp 0
transform -1 0 390 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2620_
timestamp 0
transform -1 0 630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2621_
timestamp 0
transform 1 0 950 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2622_
timestamp 0
transform 1 0 390 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2623_
timestamp 0
transform 1 0 2770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2624_
timestamp 0
transform 1 0 1970 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2625_
timestamp 0
transform -1 0 2230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2626_
timestamp 0
transform -1 0 1950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2627_
timestamp 0
transform 1 0 90 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2628_
timestamp 0
transform 1 0 90 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2629_
timestamp 0
transform -1 0 350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2630_
timestamp 0
transform 1 0 90 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2631_
timestamp 0
transform 1 0 5030 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2632_
timestamp 0
transform 1 0 2270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2633_
timestamp 0
transform -1 0 2570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2634_
timestamp 0
transform -1 0 110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2635_
timestamp 0
transform 1 0 90 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2636_
timestamp 0
transform 1 0 630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2637_
timestamp 0
transform 1 0 970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2638_
timestamp 0
transform 1 0 390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2639_
timestamp 0
transform -1 0 710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2640_
timestamp 0
transform -1 0 110 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2641_
timestamp 0
transform -1 0 110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2642_
timestamp 0
transform 1 0 1350 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2643_
timestamp 0
transform -1 0 1890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2644_
timestamp 0
transform 1 0 2290 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2645_
timestamp 0
transform -1 0 2030 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2646_
timestamp 0
transform -1 0 1230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2647_
timestamp 0
transform 1 0 90 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2648_
timestamp 0
transform 1 0 590 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__2649_
timestamp 0
transform 1 0 90 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2650_
timestamp 0
transform -1 0 3690 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2651_
timestamp 0
transform -1 0 3410 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2652_
timestamp 0
transform 1 0 630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2653_
timestamp 0
transform 1 0 350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2654_
timestamp 0
transform 1 0 1230 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2655_
timestamp 0
transform 1 0 670 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2656_
timestamp 0
transform -1 0 950 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2657_
timestamp 0
transform 1 0 90 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2658_
timestamp 0
transform 1 0 90 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2659_
timestamp 0
transform -1 0 390 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2660_
timestamp 0
transform 1 0 330 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2661_
timestamp 0
transform -1 0 2650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__2662_
timestamp 0
transform -1 0 2590 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2663_
timestamp 0
transform -1 0 2010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2664_
timestamp 0
transform 1 0 910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2665_
timestamp 0
transform -1 0 870 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2666_
timestamp 0
transform -1 0 390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2667_
timestamp 0
transform -1 0 610 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2668_
timestamp 0
transform 1 0 1110 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2669_
timestamp 0
transform -1 0 2870 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2670_
timestamp 0
transform -1 0 2990 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2671_
timestamp 0
transform 1 0 1150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2672_
timestamp 0
transform -1 0 650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2673_
timestamp 0
transform -1 0 610 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2674_
timestamp 0
transform 1 0 870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2675_
timestamp 0
transform 1 0 850 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2676_
timestamp 0
transform -1 0 1150 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2677_
timestamp 0
transform 1 0 6490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__2678_
timestamp 0
transform -1 0 6410 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2679_
timestamp 0
transform 1 0 7030 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2680_
timestamp 0
transform -1 0 6830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2681_
timestamp 0
transform 1 0 7090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2682_
timestamp 0
transform -1 0 6810 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2683_
timestamp 0
transform -1 0 1930 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2684_
timestamp 0
transform -1 0 1750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__2685_
timestamp 0
transform 1 0 1670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2686_
timestamp 0
transform 1 0 1670 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2687_
timestamp 0
transform 1 0 1410 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2688_
timestamp 0
transform -1 0 850 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2689_
timestamp 0
transform -1 0 830 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2690_
timestamp 0
transform 1 0 7330 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2691_
timestamp 0
transform -1 0 7170 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2692_
timestamp 0
transform -1 0 5110 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2693_
timestamp 0
transform -1 0 3070 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2694_
timestamp 0
transform -1 0 1370 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2695_
timestamp 0
transform -1 0 1650 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2696_
timestamp 0
transform -1 0 1370 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2697_
timestamp 0
transform 1 0 1950 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2698_
timestamp 0
transform -1 0 590 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2699_
timestamp 0
transform 1 0 6350 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2700_
timestamp 0
transform -1 0 7070 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2701_
timestamp 0
transform 1 0 7650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2702_
timestamp 0
transform 1 0 7350 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2703_
timestamp 0
transform 1 0 7510 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2704_
timestamp 0
transform -1 0 6710 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2705_
timestamp 0
transform 1 0 1630 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2706_
timestamp 0
transform 1 0 1070 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2707_
timestamp 0
transform 1 0 2770 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2708_
timestamp 0
transform 1 0 2450 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2709_
timestamp 0
transform -1 0 1130 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2710_
timestamp 0
transform -1 0 910 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2711_
timestamp 0
transform -1 0 1190 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2712_
timestamp 0
transform 1 0 2930 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2713_
timestamp 0
transform -1 0 4330 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2714_
timestamp 0
transform -1 0 4750 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2715_
timestamp 0
transform 1 0 3590 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2716_
timestamp 0
transform -1 0 4350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2717_
timestamp 0
transform -1 0 5910 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__2718_
timestamp 0
transform -1 0 4150 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2719_
timestamp 0
transform 1 0 3750 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2720_
timestamp 0
transform -1 0 4050 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2721_
timestamp 0
transform -1 0 2210 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2722_
timestamp 0
transform 1 0 2330 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2723_
timestamp 0
transform 1 0 2630 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2724_
timestamp 0
transform -1 0 870 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2725_
timestamp 0
transform -1 0 5470 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2726_
timestamp 0
transform -1 0 6650 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2727_
timestamp 0
transform 1 0 3910 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2728_
timestamp 0
transform 1 0 3630 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2729_
timestamp 0
transform -1 0 3590 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2730_
timestamp 0
transform 1 0 3190 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2731_
timestamp 0
transform 1 0 2050 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2732_
timestamp 0
transform -1 0 1930 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2733_
timestamp 0
transform 1 0 1470 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2734_
timestamp 0
transform -1 0 1770 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2735_
timestamp 0
transform -1 0 3930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2736_
timestamp 0
transform -1 0 4070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2737_
timestamp 0
transform -1 0 4150 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2738_
timestamp 0
transform -1 0 3850 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2739_
timestamp 0
transform -1 0 3290 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2740_
timestamp 0
transform -1 0 3370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2741_
timestamp 0
transform -1 0 1130 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2742_
timestamp 0
transform 1 0 1430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2743_
timestamp 0
transform 1 0 1370 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2744_
timestamp 0
transform 1 0 1910 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2745_
timestamp 0
transform 1 0 570 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2746_
timestamp 0
transform 1 0 3630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2747_
timestamp 0
transform 1 0 4750 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__2748_
timestamp 0
transform 1 0 4410 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2749_
timestamp 0
transform -1 0 3570 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2750_
timestamp 0
transform -1 0 3010 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2751_
timestamp 0
transform 1 0 2850 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2752_
timestamp 0
transform 1 0 1150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2753_
timestamp 0
transform 1 0 650 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2754_
timestamp 0
transform -1 0 590 0 1 790
box -6 -8 26 268
use FILL  FILL_4__2755_
timestamp 0
transform -1 0 3110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2756_
timestamp 0
transform -1 0 2550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2757_
timestamp 0
transform 1 0 2790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2758_
timestamp 0
transform 1 0 2270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2759_
timestamp 0
transform -1 0 4350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2760_
timestamp 0
transform 1 0 3790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2761_
timestamp 0
transform 1 0 4130 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2762_
timestamp 0
transform -1 0 3870 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2763_
timestamp 0
transform -1 0 2110 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2764_
timestamp 0
transform -1 0 1830 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2765_
timestamp 0
transform -1 0 1750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2766_
timestamp 0
transform -1 0 2010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__2767_
timestamp 0
transform -1 0 1530 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__2768_
timestamp 0
transform 1 0 2190 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2769_
timestamp 0
transform 1 0 1630 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__2770_
timestamp 0
transform 1 0 5990 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2771_
timestamp 0
transform 1 0 6530 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2772_
timestamp 0
transform 1 0 4970 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__2773_
timestamp 0
transform 1 0 4170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2774_
timestamp 0
transform 1 0 2330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2775_
timestamp 0
transform 1 0 2570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2776_
timestamp 0
transform 1 0 3390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2777_
timestamp 0
transform -1 0 2870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2778_
timestamp 0
transform -1 0 3130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__2779_
timestamp 0
transform -1 0 7170 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2780_
timestamp 0
transform -1 0 7410 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__2781_
timestamp 0
transform 1 0 7890 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__2782_
timestamp 0
transform 1 0 7770 0 1 270
box -6 -8 26 268
use FILL  FILL_4__2783_
timestamp 0
transform 1 0 9710 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2784_
timestamp 0
transform 1 0 10850 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2785_
timestamp 0
transform 1 0 10230 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2786_
timestamp 0
transform 1 0 9950 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2787_
timestamp 0
transform 1 0 8410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2788_
timestamp 0
transform 1 0 8670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2789_
timestamp 0
transform 1 0 8190 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2790_
timestamp 0
transform -1 0 7930 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2791_
timestamp 0
transform 1 0 6190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2792_
timestamp 0
transform 1 0 9810 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2793_
timestamp 0
transform 1 0 10010 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2794_
timestamp 0
transform -1 0 10270 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2795_
timestamp 0
transform 1 0 8450 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2796_
timestamp 0
transform 1 0 8430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2797_
timestamp 0
transform 1 0 10830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2798_
timestamp 0
transform -1 0 9970 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2799_
timestamp 0
transform -1 0 8350 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2800_
timestamp 0
transform -1 0 7750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2801_
timestamp 0
transform 1 0 9690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2802_
timestamp 0
transform -1 0 10010 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2803_
timestamp 0
transform 1 0 8450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2804_
timestamp 0
transform -1 0 8350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2805_
timestamp 0
transform -1 0 10090 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2806_
timestamp 0
transform 1 0 9770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2807_
timestamp 0
transform -1 0 8390 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2808_
timestamp 0
transform -1 0 6630 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2809_
timestamp 0
transform 1 0 8150 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2810_
timestamp 0
transform -1 0 7570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2811_
timestamp 0
transform 1 0 10050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2812_
timestamp 0
transform 1 0 9690 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2813_
timestamp 0
transform 1 0 8270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2814_
timestamp 0
transform -1 0 8150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2815_
timestamp 0
transform -1 0 8230 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2816_
timestamp 0
transform 1 0 9490 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2817_
timestamp 0
transform -1 0 10350 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2818_
timestamp 0
transform 1 0 11170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2819_
timestamp 0
transform 1 0 10150 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2820_
timestamp 0
transform -1 0 9930 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2821_
timestamp 0
transform -1 0 9790 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2822_
timestamp 0
transform -1 0 7510 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2823_
timestamp 0
transform -1 0 9510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2824_
timestamp 0
transform -1 0 9250 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2825_
timestamp 0
transform 1 0 8710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2826_
timestamp 0
transform 1 0 8750 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2827_
timestamp 0
transform 1 0 9170 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2828_
timestamp 0
transform 1 0 10290 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2829_
timestamp 0
transform -1 0 9230 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2830_
timestamp 0
transform 1 0 9850 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2831_
timestamp 0
transform 1 0 9030 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2832_
timestamp 0
transform -1 0 8950 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2833_
timestamp 0
transform -1 0 8710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2834_
timestamp 0
transform -1 0 8290 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2835_
timestamp 0
transform -1 0 9310 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2836_
timestamp 0
transform -1 0 8010 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2837_
timestamp 0
transform 1 0 8090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2838_
timestamp 0
transform 1 0 9330 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2839_
timestamp 0
transform 1 0 9590 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2840_
timestamp 0
transform -1 0 9330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2841_
timestamp 0
transform 1 0 8230 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2842_
timestamp 0
transform 1 0 11550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2843_
timestamp 0
transform -1 0 11050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2844_
timestamp 0
transform 1 0 10770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2845_
timestamp 0
transform 1 0 10510 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2846_
timestamp 0
transform -1 0 10150 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2847_
timestamp 0
transform 1 0 10350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2848_
timestamp 0
transform -1 0 9630 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2849_
timestamp 0
transform 1 0 10930 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__2850_
timestamp 0
transform 1 0 11090 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2851_
timestamp 0
transform 1 0 11330 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2852_
timestamp 0
transform 1 0 12030 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2853_
timestamp 0
transform 1 0 12090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2854_
timestamp 0
transform 1 0 11770 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2855_
timestamp 0
transform 1 0 12050 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2856_
timestamp 0
transform -1 0 9090 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2857_
timestamp 0
transform 1 0 9590 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2858_
timestamp 0
transform -1 0 9890 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2859_
timestamp 0
transform 1 0 10830 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2860_
timestamp 0
transform 1 0 7710 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2861_
timestamp 0
transform 1 0 8390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2862_
timestamp 0
transform -1 0 7770 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2863_
timestamp 0
transform 1 0 7470 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2864_
timestamp 0
transform 1 0 9710 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2865_
timestamp 0
transform 1 0 8870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2866_
timestamp 0
transform -1 0 6970 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2867_
timestamp 0
transform -1 0 8810 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2868_
timestamp 0
transform -1 0 8530 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2869_
timestamp 0
transform -1 0 8970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2870_
timestamp 0
transform 1 0 8610 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2871_
timestamp 0
transform 1 0 8570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2872_
timestamp 0
transform 1 0 5510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2873_
timestamp 0
transform -1 0 5530 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2874_
timestamp 0
transform 1 0 5450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2875_
timestamp 0
transform -1 0 5810 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2876_
timestamp 0
transform 1 0 5490 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2877_
timestamp 0
transform 1 0 6070 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2878_
timestamp 0
transform -1 0 5810 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2879_
timestamp 0
transform -1 0 8950 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2880_
timestamp 0
transform -1 0 11950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2881_
timestamp 0
transform 1 0 11630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2882_
timestamp 0
transform -1 0 9230 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2883_
timestamp 0
transform 1 0 9030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2884_
timestamp 0
transform -1 0 9350 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2885_
timestamp 0
transform -1 0 10530 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2886_
timestamp 0
transform 1 0 10490 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2887_
timestamp 0
transform -1 0 8910 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2888_
timestamp 0
transform -1 0 9190 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2889_
timestamp 0
transform 1 0 9470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2890_
timestamp 0
transform -1 0 9830 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__2891_
timestamp 0
transform -1 0 9770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2892_
timestamp 0
transform 1 0 9150 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2893_
timestamp 0
transform -1 0 9310 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2894_
timestamp 0
transform -1 0 11130 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2895_
timestamp 0
transform 1 0 10810 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2896_
timestamp 0
transform -1 0 11090 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2897_
timestamp 0
transform -1 0 10810 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2898_
timestamp 0
transform 1 0 9430 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2899_
timestamp 0
transform -1 0 9730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2900_
timestamp 0
transform 1 0 10410 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2901_
timestamp 0
transform -1 0 10430 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2902_
timestamp 0
transform 1 0 10610 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2903_
timestamp 0
transform -1 0 10730 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2904_
timestamp 0
transform -1 0 9890 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2905_
timestamp 0
transform -1 0 9390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2906_
timestamp 0
transform -1 0 8550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2907_
timestamp 0
transform -1 0 9110 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2908_
timestamp 0
transform -1 0 10450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2909_
timestamp 0
transform 1 0 11810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2910_
timestamp 0
transform 1 0 10890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2911_
timestamp 0
transform 1 0 11750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2912_
timestamp 0
transform 1 0 12030 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__2913_
timestamp 0
transform 1 0 10630 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__2914_
timestamp 0
transform -1 0 7810 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2915_
timestamp 0
transform 1 0 10950 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2916_
timestamp 0
transform 1 0 11190 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__2917_
timestamp 0
transform 1 0 10690 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2918_
timestamp 0
transform -1 0 10850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2919_
timestamp 0
transform 1 0 8530 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2920_
timestamp 0
transform 1 0 11230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2921_
timestamp 0
transform 1 0 11750 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__2922_
timestamp 0
transform -1 0 11870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2923_
timestamp 0
transform 1 0 11330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2924_
timestamp 0
transform 1 0 10250 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2925_
timestamp 0
transform 1 0 10010 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2926_
timestamp 0
transform 1 0 10150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2927_
timestamp 0
transform -1 0 9990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2928_
timestamp 0
transform -1 0 10250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__2929_
timestamp 0
transform -1 0 10370 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__2930_
timestamp 0
transform -1 0 11250 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2931_
timestamp 0
transform -1 0 11510 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__2932_
timestamp 0
transform 1 0 11470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__2933_
timestamp 0
transform 1 0 11430 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__2934_
timestamp 0
transform 1 0 11510 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__2935_
timestamp 0
transform 1 0 11590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2936_
timestamp 0
transform 1 0 10530 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__2937_
timestamp 0
transform -1 0 3530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__2938_
timestamp 0
transform -1 0 7750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2939_
timestamp 0
transform 1 0 6510 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2940_
timestamp 0
transform -1 0 6290 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2941_
timestamp 0
transform -1 0 6210 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2942_
timestamp 0
transform 1 0 5110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2943_
timestamp 0
transform -1 0 7010 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__2944_
timestamp 0
transform 1 0 5390 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2945_
timestamp 0
transform -1 0 6790 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2946_
timestamp 0
transform 1 0 6390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__2947_
timestamp 0
transform 1 0 7870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2948_
timestamp 0
transform 1 0 7610 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2949_
timestamp 0
transform 1 0 5710 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__2950_
timestamp 0
transform -1 0 6050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2951_
timestamp 0
transform 1 0 6810 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2952_
timestamp 0
transform 1 0 6530 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2953_
timestamp 0
transform 1 0 5690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2954_
timestamp 0
transform -1 0 5990 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__2955_
timestamp 0
transform 1 0 7070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2956_
timestamp 0
transform 1 0 6550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__2957_
timestamp 0
transform -1 0 8170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__2958_
timestamp 0
transform 1 0 6550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__2959_
timestamp 0
transform 1 0 6290 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2960_
timestamp 0
transform -1 0 7170 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2961_
timestamp 0
transform 1 0 6550 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2962_
timestamp 0
transform -1 0 6330 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__2963_
timestamp 0
transform -1 0 6630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2964_
timestamp 0
transform 1 0 4690 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2965_
timestamp 0
transform 1 0 5750 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2966_
timestamp 0
transform -1 0 6650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__2967_
timestamp 0
transform -1 0 5070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2968_
timestamp 0
transform -1 0 5330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2969_
timestamp 0
transform 1 0 4410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2970_
timestamp 0
transform 1 0 4770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2971_
timestamp 0
transform 1 0 4650 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2972_
timestamp 0
transform -1 0 6090 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2973_
timestamp 0
transform -1 0 6350 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2974_
timestamp 0
transform -1 0 6350 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2975_
timestamp 0
transform 1 0 5810 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2976_
timestamp 0
transform -1 0 4730 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2977_
timestamp 0
transform -1 0 4990 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2978_
timestamp 0
transform 1 0 5250 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__2979_
timestamp 0
transform 1 0 5530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__2980_
timestamp 0
transform -1 0 7410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2981_
timestamp 0
transform -1 0 6370 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2982_
timestamp 0
transform -1 0 6650 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__2983_
timestamp 0
transform 1 0 7170 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2984_
timestamp 0
transform 1 0 6570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__2985_
timestamp 0
transform -1 0 6910 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2986_
timestamp 0
transform 1 0 6610 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2987_
timestamp 0
transform 1 0 6050 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2988_
timestamp 0
transform -1 0 6330 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__2989_
timestamp 0
transform -1 0 7910 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2990_
timestamp 0
transform 1 0 7030 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__2991_
timestamp 0
transform -1 0 6890 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2992_
timestamp 0
transform -1 0 5190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__2993_
timestamp 0
transform -1 0 6050 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2994_
timestamp 0
transform 1 0 5510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2995_
timestamp 0
transform 1 0 6590 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2996_
timestamp 0
transform 1 0 6310 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__2997_
timestamp 0
transform 1 0 6030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2998_
timestamp 0
transform -1 0 5770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__2999_
timestamp 0
transform 1 0 6430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3000_
timestamp 0
transform -1 0 5770 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__3001_
timestamp 0
transform 1 0 4990 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3002_
timestamp 0
transform -1 0 5490 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__3003_
timestamp 0
transform -1 0 5850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3004_
timestamp 0
transform -1 0 5270 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3005_
timestamp 0
transform -1 0 5530 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3006_
timestamp 0
transform -1 0 7430 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3007_
timestamp 0
transform 1 0 6850 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3008_
timestamp 0
transform 1 0 8650 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3009_
timestamp 0
transform 1 0 8110 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3010_
timestamp 0
transform 1 0 7130 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3011_
timestamp 0
transform -1 0 7230 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3012_
timestamp 0
transform -1 0 7110 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3013_
timestamp 0
transform -1 0 7850 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3014_
timestamp 0
transform 1 0 7050 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3015_
timestamp 0
transform -1 0 7330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3016_
timestamp 0
transform -1 0 6090 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3017_
timestamp 0
transform -1 0 6890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3018_
timestamp 0
transform -1 0 6570 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3019_
timestamp 0
transform -1 0 6830 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3020_
timestamp 0
transform 1 0 5470 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__3021_
timestamp 0
transform 1 0 5910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3022_
timestamp 0
transform 1 0 5710 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__3023_
timestamp 0
transform -1 0 6790 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3024_
timestamp 0
transform -1 0 6710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3025_
timestamp 0
transform 1 0 5990 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__3026_
timestamp 0
transform 1 0 5410 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__3027_
timestamp 0
transform -1 0 5510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3028_
timestamp 0
transform 1 0 5990 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3029_
timestamp 0
transform 1 0 6750 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3030_
timestamp 0
transform 1 0 4890 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__3031_
timestamp 0
transform 1 0 4430 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3032_
timestamp 0
transform -1 0 5210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3033_
timestamp 0
transform 1 0 5470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3034_
timestamp 0
transform -1 0 3410 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3035_
timestamp 0
transform -1 0 3970 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3036_
timestamp 0
transform -1 0 3470 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3037_
timestamp 0
transform -1 0 3350 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3038_
timestamp 0
transform 1 0 3570 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3039_
timestamp 0
transform -1 0 3070 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3040_
timestamp 0
transform 1 0 2950 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3041_
timestamp 0
transform 1 0 3190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3042_
timestamp 0
transform -1 0 3750 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3043_
timestamp 0
transform -1 0 3850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3044_
timestamp 0
transform -1 0 3610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3045_
timestamp 0
transform 1 0 4410 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3046_
timestamp 0
transform 1 0 4130 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3047_
timestamp 0
transform -1 0 3090 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3048_
timestamp 0
transform 1 0 3130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3049_
timestamp 0
transform -1 0 2830 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3050_
timestamp 0
transform 1 0 2870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3051_
timestamp 0
transform 1 0 2610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3052_
timestamp 0
transform 1 0 2510 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3053_
timestamp 0
transform 1 0 3270 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3054_
timestamp 0
transform -1 0 3550 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3055_
timestamp 0
transform 1 0 3370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3056_
timestamp 0
transform -1 0 3630 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3057_
timestamp 0
transform 1 0 3830 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3058_
timestamp 0
transform 1 0 4010 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3059_
timestamp 0
transform 1 0 4290 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3060_
timestamp 0
transform 1 0 4130 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3061_
timestamp 0
transform 1 0 3610 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3062_
timestamp 0
transform -1 0 3850 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3063_
timestamp 0
transform -1 0 5090 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__3064_
timestamp 0
transform 1 0 4950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__3065_
timestamp 0
transform -1 0 4690 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3066_
timestamp 0
transform 1 0 4590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3067_
timestamp 0
transform -1 0 3690 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3068_
timestamp 0
transform -1 0 3430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3069_
timestamp 0
transform 1 0 3630 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3070_
timestamp 0
transform -1 0 4530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__3071_
timestamp 0
transform 1 0 4250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__3072_
timestamp 0
transform -1 0 4190 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3073_
timestamp 0
transform -1 0 4450 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3074_
timestamp 0
transform 1 0 5730 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3075_
timestamp 0
transform 1 0 5450 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3076_
timestamp 0
transform 1 0 3690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3077_
timestamp 0
transform 1 0 4010 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3078_
timestamp 0
transform 1 0 4070 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3079_
timestamp 0
transform -1 0 4150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3080_
timestamp 0
transform 1 0 6290 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3081_
timestamp 0
transform -1 0 6950 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3082_
timestamp 0
transform 1 0 6650 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3083_
timestamp 0
transform -1 0 3830 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3084_
timestamp 0
transform 1 0 3530 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3085_
timestamp 0
transform 1 0 3150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3086_
timestamp 0
transform -1 0 2870 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3087_
timestamp 0
transform 1 0 4350 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3088_
timestamp 0
transform -1 0 4950 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3089_
timestamp 0
transform 1 0 3430 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3090_
timestamp 0
transform -1 0 3710 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3091_
timestamp 0
transform -1 0 6250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3092_
timestamp 0
transform 1 0 5470 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3093_
timestamp 0
transform 1 0 5730 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3094_
timestamp 0
transform 1 0 5450 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3095_
timestamp 0
transform -1 0 4650 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3096_
timestamp 0
transform 1 0 4350 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3097_
timestamp 0
transform -1 0 4110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3098_
timestamp 0
transform 1 0 3810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3099_
timestamp 0
transform -1 0 3870 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3100_
timestamp 0
transform -1 0 3690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3101_
timestamp 0
transform 1 0 4910 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3102_
timestamp 0
transform -1 0 5210 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3103_
timestamp 0
transform -1 0 4590 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3104_
timestamp 0
transform -1 0 4870 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3105_
timestamp 0
transform 1 0 5650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3106_
timestamp 0
transform -1 0 5950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3107_
timestamp 0
transform -1 0 4050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3108_
timestamp 0
transform 1 0 3750 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3109_
timestamp 0
transform 1 0 6230 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3110_
timestamp 0
transform 1 0 3910 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3111_
timestamp 0
transform 1 0 5770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3112_
timestamp 0
transform -1 0 5190 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3113_
timestamp 0
transform -1 0 4650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3114_
timestamp 0
transform 1 0 4350 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3115_
timestamp 0
transform 1 0 4870 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3116_
timestamp 0
transform 1 0 3810 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3117_
timestamp 0
transform 1 0 4430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3118_
timestamp 0
transform -1 0 4730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3119_
timestamp 0
transform 1 0 4910 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3120_
timestamp 0
transform 1 0 4610 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3121_
timestamp 0
transform 1 0 5210 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3122_
timestamp 0
transform 1 0 5490 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3123_
timestamp 0
transform 1 0 5470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3124_
timestamp 0
transform -1 0 5770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3125_
timestamp 0
transform -1 0 4130 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3126_
timestamp 0
transform 1 0 3830 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3127_
timestamp 0
transform 1 0 6490 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3128_
timestamp 0
transform 1 0 6050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3129_
timestamp 0
transform 1 0 5450 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3130_
timestamp 0
transform -1 0 3370 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3131_
timestamp 0
transform -1 0 3610 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3132_
timestamp 0
transform 1 0 4710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3133_
timestamp 0
transform 1 0 3950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3134_
timestamp 0
transform 1 0 5130 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3135_
timestamp 0
transform 1 0 4830 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3136_
timestamp 0
transform 1 0 5730 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3137_
timestamp 0
transform 1 0 5450 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3138_
timestamp 0
transform 1 0 5730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3139_
timestamp 0
transform 1 0 5450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3140_
timestamp 0
transform -1 0 5650 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3141_
timestamp 0
transform -1 0 5910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3142_
timestamp 0
transform -1 0 4250 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3143_
timestamp 0
transform -1 0 4510 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3144_
timestamp 0
transform 1 0 11590 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__3145_
timestamp 0
transform 1 0 11830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__3146_
timestamp 0
transform -1 0 11890 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__3147_
timestamp 0
transform 1 0 9510 0 1 790
box -6 -8 26 268
use FILL  FILL_4__3148_
timestamp 0
transform -1 0 11890 0 1 790
box -6 -8 26 268
use FILL  FILL_4__3149_
timestamp 0
transform -1 0 11510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3150_
timestamp 0
transform -1 0 11790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3151_
timestamp 0
transform -1 0 10730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3152_
timestamp 0
transform 1 0 9370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3153_
timestamp 0
transform -1 0 9670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3154_
timestamp 0
transform -1 0 10190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3155_
timestamp 0
transform -1 0 10310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3156_
timestamp 0
transform -1 0 8950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__3157_
timestamp 0
transform -1 0 8990 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__3158_
timestamp 0
transform -1 0 8710 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__3159_
timestamp 0
transform -1 0 8690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__3160_
timestamp 0
transform 1 0 10530 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3161_
timestamp 0
transform 1 0 10250 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3162_
timestamp 0
transform -1 0 9790 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3163_
timestamp 0
transform 1 0 9510 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3164_
timestamp 0
transform -1 0 8990 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3165_
timestamp 0
transform -1 0 7210 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3166_
timestamp 0
transform 1 0 7610 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__3167_
timestamp 0
transform 1 0 7470 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3168_
timestamp 0
transform 1 0 7630 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3169_
timestamp 0
transform -1 0 8710 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3170_
timestamp 0
transform -1 0 8430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3171_
timestamp 0
transform -1 0 9150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3172_
timestamp 0
transform -1 0 8150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3173_
timestamp 0
transform 1 0 8410 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3174_
timestamp 0
transform 1 0 7890 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3175_
timestamp 0
transform -1 0 7870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3176_
timestamp 0
transform -1 0 7590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3177_
timestamp 0
transform -1 0 11870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__3178_
timestamp 0
transform -1 0 11810 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3179_
timestamp 0
transform 1 0 12070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3180_
timestamp 0
transform 1 0 12130 0 1 790
box -6 -8 26 268
use FILL  FILL_4__3181_
timestamp 0
transform 1 0 12110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__3182_
timestamp 0
transform -1 0 11330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3183_
timestamp 0
transform 1 0 11590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3184_
timestamp 0
transform 1 0 11870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3185_
timestamp 0
transform 1 0 11890 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3186_
timestamp 0
transform 1 0 12070 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3187_
timestamp 0
transform 1 0 9930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__3188_
timestamp 0
transform 1 0 10810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3189_
timestamp 0
transform -1 0 11070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__3190_
timestamp 0
transform 1 0 11110 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3191_
timestamp 0
transform 1 0 11050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3192_
timestamp 0
transform -1 0 10770 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3193_
timestamp 0
transform 1 0 10190 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3194_
timestamp 0
transform 1 0 10810 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__3195_
timestamp 0
transform -1 0 10550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3196_
timestamp 0
transform 1 0 10450 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3197_
timestamp 0
transform -1 0 7310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3198_
timestamp 0
transform -1 0 4670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3199_
timestamp 0
transform 1 0 2830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__3200_
timestamp 0
transform 1 0 4810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__3201_
timestamp 0
transform 1 0 4530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__3202_
timestamp 0
transform 1 0 1590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__3203_
timestamp 0
transform 1 0 1550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3204_
timestamp 0
transform 1 0 1510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__3205_
timestamp 0
transform 1 0 1070 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__3206_
timestamp 0
transform 1 0 1490 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__3207_
timestamp 0
transform -1 0 1630 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__3208_
timestamp 0
transform -1 0 970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__3209_
timestamp 0
transform -1 0 670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__3210_
timestamp 0
transform -1 0 4330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__3211_
timestamp 0
transform 1 0 4270 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__3212_
timestamp 0
transform 1 0 1230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__3213_
timestamp 0
transform 1 0 1130 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__3214_
timestamp 0
transform -1 0 2410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3215_
timestamp 0
transform 1 0 1830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3216_
timestamp 0
transform 1 0 5770 0 1 270
box -6 -8 26 268
use FILL  FILL_4__3217_
timestamp 0
transform -1 0 6070 0 1 270
box -6 -8 26 268
use FILL  FILL_4__3218_
timestamp 0
transform 1 0 6110 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3219_
timestamp 0
transform -1 0 6390 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3220_
timestamp 0
transform 1 0 3730 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3221_
timestamp 0
transform -1 0 4010 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3222_
timestamp 0
transform -1 0 3610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3223_
timestamp 0
transform 1 0 3330 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__3224_
timestamp 0
transform -1 0 3310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3225_
timestamp 0
transform 1 0 5450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__3226_
timestamp 0
transform 1 0 5170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__3227_
timestamp 0
transform -1 0 4290 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3228_
timestamp 0
transform -1 0 4490 0 1 270
box -6 -8 26 268
use FILL  FILL_4__3229_
timestamp 0
transform 1 0 2730 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__3230_
timestamp 0
transform -1 0 2770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__3231_
timestamp 0
transform 1 0 6010 0 1 790
box -6 -8 26 268
use FILL  FILL_4__3232_
timestamp 0
transform 1 0 5990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__3364_
timestamp 0
transform 1 0 5270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3365_
timestamp 0
transform 1 0 4470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3366_
timestamp 0
transform 1 0 4950 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__3367_
timestamp 0
transform -1 0 4750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3368_
timestamp 0
transform -1 0 5010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3369_
timestamp 0
transform -1 0 5570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3370_
timestamp 0
transform 1 0 2710 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3371_
timestamp 0
transform 1 0 2210 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3372_
timestamp 0
transform -1 0 2330 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3373_
timestamp 0
transform -1 0 3990 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3374_
timestamp 0
transform -1 0 2310 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3375_
timestamp 0
transform 1 0 2310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3376_
timestamp 0
transform -1 0 2970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3377_
timestamp 0
transform 1 0 2430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3378_
timestamp 0
transform -1 0 2290 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3379_
timestamp 0
transform -1 0 1450 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3380_
timestamp 0
transform 1 0 1230 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3381_
timestamp 0
transform -1 0 1490 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3382_
timestamp 0
transform -1 0 1950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3383_
timestamp 0
transform -1 0 1510 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3384_
timestamp 0
transform 1 0 1770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3385_
timestamp 0
transform 1 0 1470 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3386_
timestamp 0
transform -1 0 2050 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3387_
timestamp 0
transform 1 0 2310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3388_
timestamp 0
transform -1 0 650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3389_
timestamp 0
transform 1 0 2510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3390_
timestamp 0
transform 1 0 3330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3391_
timestamp 0
transform 1 0 3050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3392_
timestamp 0
transform -1 0 2890 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3393_
timestamp 0
transform 1 0 2290 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3394_
timestamp 0
transform 1 0 690 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3395_
timestamp 0
transform -1 0 650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3396_
timestamp 0
transform -1 0 390 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3397_
timestamp 0
transform -1 0 410 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3398_
timestamp 0
transform -1 0 110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3399_
timestamp 0
transform 1 0 90 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3400_
timestamp 0
transform -1 0 890 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3401_
timestamp 0
transform -1 0 1470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3402_
timestamp 0
transform 1 0 1450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3403_
timestamp 0
transform 1 0 1170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3404_
timestamp 0
transform -1 0 110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3405_
timestamp 0
transform -1 0 370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3406_
timestamp 0
transform -1 0 110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3407_
timestamp 0
transform -1 0 390 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3408_
timestamp 0
transform -1 0 110 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3409_
timestamp 0
transform -1 0 110 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3410_
timestamp 0
transform 1 0 1430 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3411_
timestamp 0
transform 1 0 1150 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3412_
timestamp 0
transform -1 0 630 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3413_
timestamp 0
transform 1 0 370 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3414_
timestamp 0
transform 1 0 630 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4__3415_
timestamp 0
transform -1 0 950 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3416_
timestamp 0
transform 1 0 630 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3417_
timestamp 0
transform -1 0 670 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3418_
timestamp 0
transform -1 0 370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3419_
timestamp 0
transform -1 0 1190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3420_
timestamp 0
transform 1 0 890 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3421_
timestamp 0
transform 1 0 1190 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3422_
timestamp 0
transform 1 0 910 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3423_
timestamp 0
transform 1 0 1210 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3424_
timestamp 0
transform -1 0 1230 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3425_
timestamp 0
transform -1 0 950 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3426_
timestamp 0
transform 1 0 930 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4__3427_
timestamp 0
transform -1 0 1450 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3428_
timestamp 0
transform 1 0 1130 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3429_
timestamp 0
transform -1 0 910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3430_
timestamp 0
transform 1 0 1430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3431_
timestamp 0
transform 1 0 1150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3432_
timestamp 0
transform -1 0 950 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3433_
timestamp 0
transform -1 0 110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3434_
timestamp 0
transform -1 0 690 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3435_
timestamp 0
transform -1 0 970 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3436_
timestamp 0
transform -1 0 910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3437_
timestamp 0
transform 1 0 1730 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3438_
timestamp 0
transform 1 0 1190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3439_
timestamp 0
transform -1 0 1470 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3440_
timestamp 0
transform 1 0 1190 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3441_
timestamp 0
transform -1 0 630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3442_
timestamp 0
transform 1 0 1210 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3443_
timestamp 0
transform 1 0 1130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3444_
timestamp 0
transform -1 0 2030 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3445_
timestamp 0
transform 1 0 1710 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3446_
timestamp 0
transform 1 0 2070 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3447_
timestamp 0
transform 1 0 1970 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3448_
timestamp 0
transform -1 0 1770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3449_
timestamp 0
transform 1 0 1450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3450_
timestamp 0
transform -1 0 910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3451_
timestamp 0
transform 1 0 1170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3452_
timestamp 0
transform 1 0 870 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3453_
timestamp 0
transform -1 0 2190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3454_
timestamp 0
transform 1 0 3110 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3455_
timestamp 0
transform -1 0 2050 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3456_
timestamp 0
transform -1 0 1710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3457_
timestamp 0
transform -1 0 2890 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3458_
timestamp 0
transform -1 0 1750 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3459_
timestamp 0
transform -1 0 1690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3460_
timestamp 0
transform 1 0 1730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3461_
timestamp 0
transform -1 0 1950 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3462_
timestamp 0
transform -1 0 1710 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3463_
timestamp 0
transform -1 0 1470 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3464_
timestamp 0
transform 1 0 1190 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3465_
timestamp 0
transform -1 0 1450 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3466_
timestamp 0
transform 1 0 1990 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3467_
timestamp 0
transform 1 0 1990 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3468_
timestamp 0
transform 1 0 2750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3469_
timestamp 0
transform 1 0 2610 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3470_
timestamp 0
transform -1 0 2510 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3471_
timestamp 0
transform 1 0 2330 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3472_
timestamp 0
transform -1 0 2230 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3473_
timestamp 0
transform 1 0 1470 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3474_
timestamp 0
transform -1 0 1730 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3475_
timestamp 0
transform 1 0 1210 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3476_
timestamp 0
transform -1 0 950 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3477_
timestamp 0
transform 1 0 370 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3478_
timestamp 0
transform -1 0 350 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3479_
timestamp 0
transform -1 0 110 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3480_
timestamp 0
transform -1 0 110 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3481_
timestamp 0
transform -1 0 110 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3482_
timestamp 0
transform 1 0 630 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3483_
timestamp 0
transform -1 0 350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3484_
timestamp 0
transform 1 0 1970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3485_
timestamp 0
transform -1 0 2030 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3486_
timestamp 0
transform -1 0 1410 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3487_
timestamp 0
transform -1 0 1730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3488_
timestamp 0
transform -1 0 1530 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3489_
timestamp 0
transform 1 0 1470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3490_
timestamp 0
transform 1 0 1150 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3491_
timestamp 0
transform -1 0 1230 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3492_
timestamp 0
transform 1 0 1130 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3493_
timestamp 0
transform -1 0 950 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3494_
timestamp 0
transform 1 0 870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3495_
timestamp 0
transform -1 0 630 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3496_
timestamp 0
transform 1 0 390 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3497_
timestamp 0
transform -1 0 350 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3498_
timestamp 0
transform 1 0 650 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3499_
timestamp 0
transform -1 0 710 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3500_
timestamp 0
transform 1 0 650 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3501_
timestamp 0
transform 1 0 890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3502_
timestamp 0
transform -1 0 410 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3503_
timestamp 0
transform -1 0 390 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3504_
timestamp 0
transform -1 0 630 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3505_
timestamp 0
transform -1 0 390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3506_
timestamp 0
transform -1 0 110 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3507_
timestamp 0
transform -1 0 110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3508_
timestamp 0
transform 1 0 630 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3509_
timestamp 0
transform -1 0 890 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3510_
timestamp 0
transform -1 0 390 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3511_
timestamp 0
transform -1 0 110 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3512_
timestamp 0
transform 1 0 590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3513_
timestamp 0
transform -1 0 410 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3514_
timestamp 0
transform -1 0 350 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3515_
timestamp 0
transform -1 0 110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3516_
timestamp 0
transform -1 0 110 0 1 10150
box -6 -8 26 268
use FILL  FILL_4__3517_
timestamp 0
transform 1 0 650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3518_
timestamp 0
transform 1 0 870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3519_
timestamp 0
transform 1 0 2570 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3520_
timestamp 0
transform 1 0 2850 0 1 9110
box -6 -8 26 268
use FILL  FILL_4__3521_
timestamp 0
transform 1 0 3330 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3522_
timestamp 0
transform 1 0 3030 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3523_
timestamp 0
transform 1 0 2590 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3524_
timestamp 0
transform -1 0 970 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3525_
timestamp 0
transform -1 0 110 0 1 10670
box -6 -8 26 268
use FILL  FILL_4__3526_
timestamp 0
transform -1 0 110 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3527_
timestamp 0
transform -1 0 610 0 1 11190
box -6 -8 26 268
use FILL  FILL_4__3528_
timestamp 0
transform -1 0 630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_4__3529_
timestamp 0
transform -1 0 110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4__3530_
timestamp 0
transform -1 0 110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3531_
timestamp 0
transform 1 0 90 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3532_
timestamp 0
transform 1 0 330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3533_
timestamp 0
transform -1 0 110 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3534_
timestamp 0
transform -1 0 630 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3535_
timestamp 0
transform -1 0 390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4__3536_
timestamp 0
transform -1 0 370 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3537_
timestamp 0
transform -1 0 1730 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3538_
timestamp 0
transform 1 0 2490 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3539_
timestamp 0
transform -1 0 2590 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3540_
timestamp 0
transform -1 0 2330 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3541_
timestamp 0
transform -1 0 2050 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3542_
timestamp 0
transform -1 0 2230 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3543_
timestamp 0
transform 1 0 1630 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3544_
timestamp 0
transform 1 0 1990 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3545_
timestamp 0
transform 1 0 1790 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3546_
timestamp 0
transform 1 0 1910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4__3547_
timestamp 0
transform -1 0 2570 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3548_
timestamp 0
transform 1 0 2270 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4__3549_
timestamp 0
transform -1 0 2370 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3550_
timestamp 0
transform 1 0 2070 0 1 11710
box -6 -8 26 268
use FILL  FILL_4__3551_
timestamp 0
transform -1 0 2550 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3552_
timestamp 0
transform 1 0 2250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4__3553_
timestamp 0
transform -1 0 1790 0 1 8070
box -6 -8 26 268
use FILL  FILL_4__3554_
timestamp 0
transform 1 0 930 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3555_
timestamp 0
transform 1 0 330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3556_
timestamp 0
transform 1 0 1190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4__3557_
timestamp 0
transform -1 0 3090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3558_
timestamp 0
transform 1 0 2790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4__3559_
timestamp 0
transform -1 0 2550 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3560_
timestamp 0
transform 1 0 2250 0 1 9630
box -6 -8 26 268
use FILL  FILL_4__3561_
timestamp 0
transform -1 0 1970 0 1 7550
box -6 -8 26 268
use FILL  FILL_4__3562_
timestamp 0
transform -1 0 2790 0 1 8590
box -6 -8 26 268
use FILL  FILL_4__3563_
timestamp 0
transform 1 0 2190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4__3564_
timestamp 0
transform 1 0 2470 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3565_
timestamp 0
transform -1 0 1470 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3566_
timestamp 0
transform -1 0 1730 0 1 7030
box -6 -8 26 268
use FILL  FILL_4__3579_
timestamp 0
transform -1 0 5070 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3580_
timestamp 0
transform -1 0 110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__3581_
timestamp 0
transform -1 0 3490 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3582_
timestamp 0
transform -1 0 3230 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3583_
timestamp 0
transform -1 0 5350 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__3584_
timestamp 0
transform 1 0 4530 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3585_
timestamp 0
transform 1 0 2950 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3586_
timestamp 0
transform -1 0 5870 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__3587_
timestamp 0
transform 1 0 90 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3588_
timestamp 0
transform -1 0 110 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__3589_
timestamp 0
transform -1 0 110 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__3590_
timestamp 0
transform -1 0 110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__3591_
timestamp 0
transform -1 0 390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3592_
timestamp 0
transform -1 0 110 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__3593_
timestamp 0
transform -1 0 4810 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3594_
timestamp 0
transform 1 0 5850 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__3595_
timestamp 0
transform 1 0 5590 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__3596_
timestamp 0
transform -1 0 890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3597_
timestamp 0
transform -1 0 110 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__3598_
timestamp 0
transform -1 0 370 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__3599_
timestamp 0
transform -1 0 110 0 1 6510
box -6 -8 26 268
use FILL  FILL_4__3600_
timestamp 0
transform -1 0 110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__3601_
timestamp 0
transform -1 0 110 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__3602_
timestamp 0
transform -1 0 1730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__3603_
timestamp 0
transform 1 0 6890 0 -1 270
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert0
timestamp 0
transform 1 0 7910 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert1
timestamp 0
transform 1 0 9410 0 1 1830
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert2
timestamp 0
transform 1 0 8170 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert3
timestamp 0
transform 1 0 11030 0 1 1830
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert4
timestamp 0
transform 1 0 630 0 1 1830
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert5
timestamp 0
transform -1 0 12110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert6
timestamp 0
transform -1 0 9610 0 1 5470
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert7
timestamp 0
transform 1 0 7070 0 1 2350
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert8
timestamp 0
transform -1 0 890 0 1 5470
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert9
timestamp 0
transform 1 0 10150 0 1 3910
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert10
timestamp 0
transform -1 0 930 0 1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert11
timestamp 0
transform -1 0 6010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert12
timestamp 0
transform 1 0 11570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert13
timestamp 0
transform -1 0 6190 0 1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert14
timestamp 0
transform 1 0 6810 0 1 2350
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert15
timestamp 0
transform -1 0 3350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert16
timestamp 0
transform -1 0 3970 0 1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert17
timestamp 0
transform 1 0 7210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert18
timestamp 0
transform -1 0 7030 0 1 11190
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert19
timestamp 0
transform 1 0 5350 0 1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert20
timestamp 0
transform 1 0 8590 0 1 11190
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert21
timestamp 0
transform -1 0 8510 0 -1 7550
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert22
timestamp 0
transform -1 0 1470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert23
timestamp 0
transform 1 0 3450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert24
timestamp 0
transform -1 0 4350 0 1 5470
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert25
timestamp 0
transform 1 0 8190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert26
timestamp 0
transform 1 0 5130 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert27
timestamp 0
transform -1 0 1270 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert39
timestamp 0
transform 1 0 6350 0 1 4950
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert40
timestamp 0
transform 1 0 7710 0 1 3910
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert41
timestamp 0
transform -1 0 8850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert42
timestamp 0
transform -1 0 6990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert43
timestamp 0
transform -1 0 8890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert44
timestamp 0
transform -1 0 9010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert45
timestamp 0
transform 1 0 11070 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert46
timestamp 0
transform 1 0 9510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert47
timestamp 0
transform 1 0 9230 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert48
timestamp 0
transform 1 0 6970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert49
timestamp 0
transform 1 0 7230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert50
timestamp 0
transform -1 0 7610 0 1 9110
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert51
timestamp 0
transform 1 0 7570 0 1 10150
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert52
timestamp 0
transform 1 0 8970 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert53
timestamp 0
transform 1 0 10010 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert54
timestamp 0
transform 1 0 8850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert55
timestamp 0
transform 1 0 8710 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert56
timestamp 0
transform -1 0 2250 0 1 8590
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert57
timestamp 0
transform 1 0 2550 0 1 11190
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert58
timestamp 0
transform 1 0 2690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert59
timestamp 0
transform -1 0 2250 0 1 10670
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert60
timestamp 0
transform -1 0 10510 0 1 7550
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert61
timestamp 0
transform 1 0 10570 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert62
timestamp 0
transform 1 0 10530 0 1 8070
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert63
timestamp 0
transform -1 0 9190 0 1 7550
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert64
timestamp 0
transform -1 0 8630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert65
timestamp 0
transform 1 0 5230 0 1 270
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert66
timestamp 0
transform 1 0 5750 0 1 790
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert67
timestamp 0
transform -1 0 3050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert68
timestamp 0
transform 1 0 3170 0 1 270
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert69
timestamp 0
transform -1 0 6670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert70
timestamp 0
transform 1 0 8610 0 1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert71
timestamp 0
transform -1 0 9270 0 1 2870
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert72
timestamp 0
transform -1 0 6790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert73
timestamp 0
transform 1 0 8950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert74
timestamp 0
transform 1 0 10810 0 1 7030
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert75
timestamp 0
transform 1 0 2590 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert76
timestamp 0
transform -1 0 3090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert77
timestamp 0
transform 1 0 10470 0 1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert78
timestamp 0
transform 1 0 9330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert79
timestamp 0
transform -1 0 8370 0 1 7550
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert80
timestamp 0
transform 1 0 7170 0 1 5470
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert81
timestamp 0
transform 1 0 7630 0 -1 790
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert82
timestamp 0
transform -1 0 7610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert83
timestamp 0
transform -1 0 7390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert84
timestamp 0
transform 1 0 9450 0 1 8590
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert85
timestamp 0
transform -1 0 8930 0 1 8590
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert86
timestamp 0
transform -1 0 9530 0 1 2870
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert87
timestamp 0
transform 1 0 9430 0 1 4430
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert88
timestamp 0
transform -1 0 10770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert89
timestamp 0
transform 1 0 9410 0 1 3390
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert90
timestamp 0
transform 1 0 5390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert91
timestamp 0
transform -1 0 4930 0 1 10670
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert92
timestamp 0
transform -1 0 4770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert93
timestamp 0
transform 1 0 5190 0 1 10150
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert94
timestamp 0
transform -1 0 11350 0 1 9630
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert95
timestamp 0
transform -1 0 11390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert96
timestamp 0
transform -1 0 10110 0 1 11710
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert97
timestamp 0
transform 1 0 11470 0 1 11710
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert28
timestamp 0
transform -1 0 6050 0 -1 11710
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert29
timestamp 0
transform -1 0 2230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert30
timestamp 0
transform 1 0 4570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert31
timestamp 0
transform -1 0 3270 0 1 2870
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert32
timestamp 0
transform 1 0 7170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert33
timestamp 0
transform 1 0 5750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert34
timestamp 0
transform -1 0 2510 0 1 10670
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert35
timestamp 0
transform -1 0 5270 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert36
timestamp 0
transform -1 0 2390 0 1 3910
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert37
timestamp 0
transform 1 0 7410 0 -1 12230
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert38
timestamp 0
transform -1 0 4390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__1688_
timestamp 0
transform -1 0 930 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1689_
timestamp 0
transform -1 0 390 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1690_
timestamp 0
transform -1 0 650 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1691_
timestamp 0
transform 1 0 110 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1692_
timestamp 0
transform -1 0 370 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1693_
timestamp 0
transform 1 0 610 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1694_
timestamp 0
transform -1 0 5610 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__1695_
timestamp 0
transform -1 0 390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1696_
timestamp 0
transform -1 0 390 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1697_
timestamp 0
transform -1 0 1510 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__1698_
timestamp 0
transform -1 0 3450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1699_
timestamp 0
transform 1 0 2890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1700_
timestamp 0
transform -1 0 3930 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__1701_
timestamp 0
transform -1 0 630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1702_
timestamp 0
transform -1 0 630 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1703_
timestamp 0
transform 1 0 3270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1704_
timestamp 0
transform -1 0 410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1705_
timestamp 0
transform 1 0 110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1706_
timestamp 0
transform -1 0 3890 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1707_
timestamp 0
transform -1 0 650 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1708_
timestamp 0
transform 1 0 650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1709_
timestamp 0
transform 1 0 4170 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1710_
timestamp 0
transform -1 0 5650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1711_
timestamp 0
transform 1 0 5190 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1712_
timestamp 0
transform 1 0 7330 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1713_
timestamp 0
transform -1 0 9710 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1714_
timestamp 0
transform -1 0 9910 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1715_
timestamp 0
transform -1 0 8590 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1716_
timestamp 0
transform 1 0 11350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1717_
timestamp 0
transform 1 0 11150 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1718_
timestamp 0
transform 1 0 11970 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1719_
timestamp 0
transform -1 0 8850 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1720_
timestamp 0
transform -1 0 10170 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1721_
timestamp 0
transform -1 0 10190 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1722_
timestamp 0
transform -1 0 9950 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1723_
timestamp 0
transform 1 0 10050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1724_
timestamp 0
transform 1 0 9270 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1725_
timestamp 0
transform 1 0 9110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1726_
timestamp 0
transform 1 0 10210 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1727_
timestamp 0
transform -1 0 8830 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1728_
timestamp 0
transform 1 0 11610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1729_
timestamp 0
transform 1 0 10210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1730_
timestamp 0
transform 1 0 8390 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1731_
timestamp 0
transform 1 0 8630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1732_
timestamp 0
transform -1 0 7830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1733_
timestamp 0
transform 1 0 9770 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1734_
timestamp 0
transform 1 0 7470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1735_
timestamp 0
transform 1 0 10910 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1736_
timestamp 0
transform -1 0 10710 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1737_
timestamp 0
transform -1 0 10970 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1738_
timestamp 0
transform -1 0 10350 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1739_
timestamp 0
transform -1 0 10350 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1740_
timestamp 0
transform 1 0 10570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1741_
timestamp 0
transform -1 0 8470 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1742_
timestamp 0
transform -1 0 8370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1743_
timestamp 0
transform -1 0 9930 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1744_
timestamp 0
transform 1 0 9810 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1745_
timestamp 0
transform -1 0 9510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1746_
timestamp 0
transform 1 0 11370 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1747_
timestamp 0
transform 1 0 10850 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1748_
timestamp 0
transform 1 0 7570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1749_
timestamp 0
transform 1 0 7990 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__1750_
timestamp 0
transform -1 0 8110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1751_
timestamp 0
transform 1 0 7510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1752_
timestamp 0
transform -1 0 8930 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1753_
timestamp 0
transform 1 0 9790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1754_
timestamp 0
transform -1 0 8330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1755_
timestamp 0
transform -1 0 8910 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__1756_
timestamp 0
transform -1 0 11250 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1757_
timestamp 0
transform 1 0 11110 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1758_
timestamp 0
transform -1 0 9170 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1759_
timestamp 0
transform -1 0 7410 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__1760_
timestamp 0
transform 1 0 8910 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__1761_
timestamp 0
transform -1 0 9630 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1762_
timestamp 0
transform 1 0 10650 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1763_
timestamp 0
transform -1 0 9090 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1764_
timestamp 0
transform 1 0 11350 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1765_
timestamp 0
transform 1 0 8170 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1766_
timestamp 0
transform 1 0 8550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1767_
timestamp 0
transform 1 0 9250 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__1768_
timestamp 0
transform 1 0 8110 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__1769_
timestamp 0
transform 1 0 8630 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__1770_
timestamp 0
transform 1 0 9070 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__1771_
timestamp 0
transform 1 0 9030 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__1772_
timestamp 0
transform 1 0 8750 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__1773_
timestamp 0
transform 1 0 10830 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1774_
timestamp 0
transform 1 0 10830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1775_
timestamp 0
transform 1 0 10070 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1776_
timestamp 0
transform -1 0 8070 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1777_
timestamp 0
transform 1 0 8110 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1778_
timestamp 0
transform -1 0 7590 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1779_
timestamp 0
transform 1 0 5730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1780_
timestamp 0
transform -1 0 4130 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1781_
timestamp 0
transform -1 0 10850 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1782_
timestamp 0
transform 1 0 8330 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1783_
timestamp 0
transform 1 0 10570 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1784_
timestamp 0
transform -1 0 10050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1785_
timestamp 0
transform -1 0 9810 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1786_
timestamp 0
transform 1 0 10230 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1787_
timestamp 0
transform -1 0 9170 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1788_
timestamp 0
transform -1 0 8590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1789_
timestamp 0
transform 1 0 10030 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1790_
timestamp 0
transform -1 0 10090 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1791_
timestamp 0
transform -1 0 10170 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1792_
timestamp 0
transform -1 0 9710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1793_
timestamp 0
transform -1 0 9450 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1794_
timestamp 0
transform 1 0 9170 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1795_
timestamp 0
transform -1 0 8370 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1796_
timestamp 0
transform -1 0 8310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1797_
timestamp 0
transform 1 0 7150 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1798_
timestamp 0
transform 1 0 7410 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1799_
timestamp 0
transform -1 0 9430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1800_
timestamp 0
transform 1 0 11310 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1801_
timestamp 0
transform 1 0 9330 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1802_
timestamp 0
transform -1 0 8990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1803_
timestamp 0
transform 1 0 10590 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1804_
timestamp 0
transform -1 0 8610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1805_
timestamp 0
transform -1 0 8710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1806_
timestamp 0
transform 1 0 7650 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1807_
timestamp 0
transform -1 0 8110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1808_
timestamp 0
transform -1 0 8430 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1809_
timestamp 0
transform 1 0 8650 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1810_
timestamp 0
transform 1 0 8050 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1811_
timestamp 0
transform -1 0 7790 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1812_
timestamp 0
transform -1 0 8430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1813_
timestamp 0
transform -1 0 8150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1814_
timestamp 0
transform -1 0 7890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1815_
timestamp 0
transform 1 0 7910 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1816_
timestamp 0
transform -1 0 3910 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1817_
timestamp 0
transform 1 0 1390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1818_
timestamp 0
transform -1 0 6210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1819_
timestamp 0
transform -1 0 970 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1820_
timestamp 0
transform 1 0 410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1821_
timestamp 0
transform 1 0 930 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1822_
timestamp 0
transform -1 0 390 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1823_
timestamp 0
transform 1 0 1750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1824_
timestamp 0
transform 1 0 1330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__1825_
timestamp 0
transform -1 0 1170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1826_
timestamp 0
transform -1 0 430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1827_
timestamp 0
transform 1 0 930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1828_
timestamp 0
transform -1 0 1530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1829_
timestamp 0
transform -1 0 670 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1830_
timestamp 0
transform -1 0 1470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1831_
timestamp 0
transform 1 0 2050 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1832_
timestamp 0
transform -1 0 8050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1833_
timestamp 0
transform 1 0 9690 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1834_
timestamp 0
transform 1 0 9270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1835_
timestamp 0
transform -1 0 7790 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1836_
timestamp 0
transform -1 0 6450 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1837_
timestamp 0
transform -1 0 7790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1838_
timestamp 0
transform -1 0 7230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1839_
timestamp 0
transform -1 0 6210 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1840_
timestamp 0
transform 1 0 8590 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1841_
timestamp 0
transform -1 0 8210 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1842_
timestamp 0
transform -1 0 6970 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1843_
timestamp 0
transform -1 0 6690 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1844_
timestamp 0
transform 1 0 9110 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1845_
timestamp 0
transform 1 0 9650 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1846_
timestamp 0
transform -1 0 9250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1847_
timestamp 0
transform -1 0 8410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1848_
timestamp 0
transform 1 0 11250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1849_
timestamp 0
transform -1 0 11570 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1850_
timestamp 0
transform -1 0 11030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1851_
timestamp 0
transform 1 0 10390 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1852_
timestamp 0
transform -1 0 10450 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1853_
timestamp 0
transform -1 0 10470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__1854_
timestamp 0
transform -1 0 7450 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1855_
timestamp 0
transform 1 0 7430 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1856_
timestamp 0
transform 1 0 7710 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1857_
timestamp 0
transform -1 0 8850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__1858_
timestamp 0
transform -1 0 9390 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1859_
timestamp 0
transform -1 0 8850 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1860_
timestamp 0
transform 1 0 9110 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1861_
timestamp 0
transform 1 0 6850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1862_
timestamp 0
transform -1 0 8350 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__1863_
timestamp 0
transform 1 0 7710 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1864_
timestamp 0
transform -1 0 6350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1865_
timestamp 0
transform -1 0 7790 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__1866_
timestamp 0
transform -1 0 7250 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1867_
timestamp 0
transform -1 0 8030 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1868_
timestamp 0
transform 1 0 7750 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1869_
timestamp 0
transform -1 0 6050 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__1870_
timestamp 0
transform 1 0 9390 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1871_
timestamp 0
transform 1 0 8870 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1872_
timestamp 0
transform -1 0 8610 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1873_
timestamp 0
transform -1 0 7810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1874_
timestamp 0
transform -1 0 7530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1875_
timestamp 0
transform -1 0 8330 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1876_
timestamp 0
transform -1 0 6970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1877_
timestamp 0
transform -1 0 5810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__1878_
timestamp 0
transform 1 0 6690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1879_
timestamp 0
transform -1 0 7490 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1880_
timestamp 0
transform 1 0 6010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__1881_
timestamp 0
transform 1 0 6010 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__1882_
timestamp 0
transform -1 0 4970 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__1883_
timestamp 0
transform -1 0 7870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1884_
timestamp 0
transform -1 0 8110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1885_
timestamp 0
transform -1 0 8670 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__1886_
timestamp 0
transform 1 0 8510 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1887_
timestamp 0
transform -1 0 8490 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1888_
timestamp 0
transform 1 0 11630 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1889_
timestamp 0
transform -1 0 8490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1890_
timestamp 0
transform 1 0 9750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1891_
timestamp 0
transform 1 0 8910 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1892_
timestamp 0
transform -1 0 8630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1893_
timestamp 0
transform 1 0 12150 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1894_
timestamp 0
transform 1 0 12130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1895_
timestamp 0
transform 1 0 12150 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1896_
timestamp 0
transform -1 0 10770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1897_
timestamp 0
transform -1 0 9170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1898_
timestamp 0
transform 1 0 9050 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1899_
timestamp 0
transform 1 0 7490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1900_
timestamp 0
transform 1 0 9690 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1901_
timestamp 0
transform 1 0 8030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1902_
timestamp 0
transform -1 0 8250 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1903_
timestamp 0
transform 1 0 7970 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1904_
timestamp 0
transform 1 0 11890 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1905_
timestamp 0
transform 1 0 11650 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1906_
timestamp 0
transform -1 0 6530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1907_
timestamp 0
transform -1 0 7070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1908_
timestamp 0
transform -1 0 6990 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1909_
timestamp 0
transform -1 0 6750 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__1910_
timestamp 0
transform -1 0 6250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1911_
timestamp 0
transform 1 0 6830 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1912_
timestamp 0
transform 1 0 6290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__1913_
timestamp 0
transform 1 0 6230 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1914_
timestamp 0
transform 1 0 5730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1915_
timestamp 0
transform 1 0 5250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1916_
timestamp 0
transform 1 0 5250 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__1917_
timestamp 0
transform -1 0 3750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__1918_
timestamp 0
transform 1 0 3630 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__1919_
timestamp 0
transform -1 0 3910 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__1920_
timestamp 0
transform -1 0 3630 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__1921_
timestamp 0
transform -1 0 1750 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__1922_
timestamp 0
transform 1 0 7550 0 1 270
box -6 -8 26 268
use FILL  FILL_5__1923_
timestamp 0
transform 1 0 7810 0 1 790
box -6 -8 26 268
use FILL  FILL_5__1924_
timestamp 0
transform -1 0 6410 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__1925_
timestamp 0
transform -1 0 4650 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1926_
timestamp 0
transform -1 0 4010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1927_
timestamp 0
transform 1 0 2050 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__1928_
timestamp 0
transform -1 0 3210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__1929_
timestamp 0
transform 1 0 4590 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__1930_
timestamp 0
transform 1 0 3150 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__1931_
timestamp 0
transform -1 0 2930 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__1932_
timestamp 0
transform -1 0 1530 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1933_
timestamp 0
transform -1 0 8490 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1934_
timestamp 0
transform 1 0 3890 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__1935_
timestamp 0
transform -1 0 3910 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1936_
timestamp 0
transform -1 0 2590 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1937_
timestamp 0
transform -1 0 1250 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1938_
timestamp 0
transform -1 0 3610 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1939_
timestamp 0
transform -1 0 4170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1940_
timestamp 0
transform -1 0 3390 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1941_
timestamp 0
transform -1 0 3330 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1942_
timestamp 0
transform -1 0 1830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__1943_
timestamp 0
transform -1 0 3630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__1944_
timestamp 0
transform -1 0 3730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1945_
timestamp 0
transform -1 0 2990 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__1946_
timestamp 0
transform -1 0 1550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__1947_
timestamp 0
transform -1 0 4970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__1948_
timestamp 0
transform 1 0 5170 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__1949_
timestamp 0
transform 1 0 5230 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__1950_
timestamp 0
transform -1 0 4970 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__1951_
timestamp 0
transform -1 0 2010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1952_
timestamp 0
transform 1 0 4130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__1953_
timestamp 0
transform 1 0 4070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__1954_
timestamp 0
transform 1 0 4210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1955_
timestamp 0
transform -1 0 1730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1956_
timestamp 0
transform -1 0 4350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__1957_
timestamp 0
transform 1 0 4930 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__1958_
timestamp 0
transform -1 0 5210 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__1959_
timestamp 0
transform -1 0 4190 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__1960_
timestamp 0
transform -1 0 2350 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1961_
timestamp 0
transform 1 0 4170 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1962_
timestamp 0
transform 1 0 3930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1963_
timestamp 0
transform 1 0 3710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1964_
timestamp 0
transform 1 0 2050 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1965_
timestamp 0
transform 1 0 6430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__1966_
timestamp 0
transform 1 0 6370 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1967_
timestamp 0
transform 1 0 7210 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1968_
timestamp 0
transform 1 0 6670 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1969_
timestamp 0
transform -1 0 3330 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__1970_
timestamp 0
transform 1 0 2870 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1971_
timestamp 0
transform -1 0 4750 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1972_
timestamp 0
transform 1 0 3610 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1973_
timestamp 0
transform -1 0 3630 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__1974_
timestamp 0
transform -1 0 3130 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__1975_
timestamp 0
transform 1 0 3030 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__1976_
timestamp 0
transform -1 0 3130 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__1977_
timestamp 0
transform 1 0 4410 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__1978_
timestamp 0
transform 1 0 3110 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__1979_
timestamp 0
transform -1 0 2850 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__1980_
timestamp 0
transform -1 0 2370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1981_
timestamp 0
transform 1 0 5990 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__1982_
timestamp 0
transform 1 0 6110 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__1983_
timestamp 0
transform 1 0 6310 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__1984_
timestamp 0
transform 1 0 5310 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__1985_
timestamp 0
transform -1 0 4810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1986_
timestamp 0
transform 1 0 2590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__1987_
timestamp 0
transform -1 0 7310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__1988_
timestamp 0
transform 1 0 7610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__1989_
timestamp 0
transform 1 0 7670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__1990_
timestamp 0
transform -1 0 7470 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1991_
timestamp 0
transform -1 0 7750 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__1992_
timestamp 0
transform 1 0 10490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__1993_
timestamp 0
transform 1 0 9610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__1994_
timestamp 0
transform -1 0 6290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__1995_
timestamp 0
transform 1 0 6670 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__1996_
timestamp 0
transform -1 0 6810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1997_
timestamp 0
transform 1 0 6510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__1998_
timestamp 0
transform 1 0 6510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__1999_
timestamp 0
transform 1 0 7570 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2000_
timestamp 0
transform 1 0 6490 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2001_
timestamp 0
transform 1 0 6730 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2002_
timestamp 0
transform 1 0 6690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2003_
timestamp 0
transform 1 0 9570 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2004_
timestamp 0
transform 1 0 7510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2005_
timestamp 0
transform -1 0 7310 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2006_
timestamp 0
transform 1 0 6790 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2007_
timestamp 0
transform 1 0 6630 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2008_
timestamp 0
transform -1 0 6270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2009_
timestamp 0
transform 1 0 6870 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2010_
timestamp 0
transform -1 0 7090 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2011_
timestamp 0
transform 1 0 7330 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2012_
timestamp 0
transform -1 0 9470 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2013_
timestamp 0
transform 1 0 10610 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2014_
timestamp 0
transform -1 0 10870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2015_
timestamp 0
transform -1 0 6310 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2016_
timestamp 0
transform -1 0 7350 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2017_
timestamp 0
transform -1 0 7130 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2018_
timestamp 0
transform 1 0 7370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2019_
timestamp 0
transform 1 0 9450 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2020_
timestamp 0
transform -1 0 10350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2021_
timestamp 0
transform -1 0 7390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2022_
timestamp 0
transform 1 0 7630 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2023_
timestamp 0
transform -1 0 7930 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2024_
timestamp 0
transform 1 0 6150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2025_
timestamp 0
transform -1 0 6030 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2026_
timestamp 0
transform 1 0 9730 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2027_
timestamp 0
transform 1 0 10270 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2028_
timestamp 0
transform -1 0 10270 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2029_
timestamp 0
transform -1 0 11150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2030_
timestamp 0
transform 1 0 10770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2031_
timestamp 0
transform -1 0 11070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2032_
timestamp 0
transform 1 0 8990 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2033_
timestamp 0
transform 1 0 8450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2034_
timestamp 0
transform 1 0 8690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2035_
timestamp 0
transform 1 0 8650 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2036_
timestamp 0
transform 1 0 11610 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2037_
timestamp 0
transform 1 0 11810 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2038_
timestamp 0
transform -1 0 7650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2039_
timestamp 0
transform -1 0 6730 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2040_
timestamp 0
transform 1 0 10990 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2041_
timestamp 0
transform 1 0 11070 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2042_
timestamp 0
transform -1 0 10150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2043_
timestamp 0
transform -1 0 10530 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2044_
timestamp 0
transform -1 0 11050 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2045_
timestamp 0
transform -1 0 11390 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2046_
timestamp 0
transform 1 0 8870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2047_
timestamp 0
transform -1 0 9430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2048_
timestamp 0
transform 1 0 9230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2049_
timestamp 0
transform 1 0 9370 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2050_
timestamp 0
transform 1 0 9130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2051_
timestamp 0
transform 1 0 8830 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2052_
timestamp 0
transform 1 0 9110 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2053_
timestamp 0
transform -1 0 9670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2054_
timestamp 0
transform 1 0 9890 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2055_
timestamp 0
transform -1 0 6530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2056_
timestamp 0
transform -1 0 6110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2057_
timestamp 0
transform 1 0 10310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2058_
timestamp 0
transform -1 0 10050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2059_
timestamp 0
transform -1 0 10190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2060_
timestamp 0
transform -1 0 9950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2061_
timestamp 0
transform 1 0 10130 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2062_
timestamp 0
transform -1 0 9210 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2063_
timestamp 0
transform 1 0 8290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2064_
timestamp 0
transform -1 0 7970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2065_
timestamp 0
transform -1 0 8790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2066_
timestamp 0
transform 1 0 8770 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2067_
timestamp 0
transform -1 0 8030 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2068_
timestamp 0
transform -1 0 8310 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2069_
timestamp 0
transform 1 0 8030 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2070_
timestamp 0
transform -1 0 8330 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2071_
timestamp 0
transform -1 0 8610 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2072_
timestamp 0
transform 1 0 8830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2073_
timestamp 0
transform 1 0 9090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2074_
timestamp 0
transform 1 0 9310 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2075_
timestamp 0
transform -1 0 9610 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2076_
timestamp 0
transform 1 0 11270 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2077_
timestamp 0
transform -1 0 11330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2078_
timestamp 0
transform -1 0 11130 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2079_
timestamp 0
transform 1 0 11270 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2080_
timestamp 0
transform -1 0 11110 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2081_
timestamp 0
transform 1 0 11110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2082_
timestamp 0
transform 1 0 10370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2083_
timestamp 0
transform 1 0 9630 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2084_
timestamp 0
transform 1 0 11650 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2085_
timestamp 0
transform 1 0 11070 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2086_
timestamp 0
transform 1 0 11570 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2087_
timestamp 0
transform 1 0 11590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2088_
timestamp 0
transform -1 0 12150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2089_
timestamp 0
transform 1 0 11870 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2090_
timestamp 0
transform 1 0 12050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2091_
timestamp 0
transform 1 0 9950 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2092_
timestamp 0
transform 1 0 10570 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2093_
timestamp 0
transform -1 0 11130 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2094_
timestamp 0
transform 1 0 11370 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2095_
timestamp 0
transform -1 0 11030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2096_
timestamp 0
transform 1 0 11550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2097_
timestamp 0
transform -1 0 11890 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2098_
timestamp 0
transform -1 0 12070 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2099_
timestamp 0
transform -1 0 11370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2100_
timestamp 0
transform 1 0 11330 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2101_
timestamp 0
transform -1 0 11290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2102_
timestamp 0
transform -1 0 11670 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2103_
timestamp 0
transform 1 0 12150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2104_
timestamp 0
transform 1 0 12150 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2105_
timestamp 0
transform -1 0 11610 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2106_
timestamp 0
transform -1 0 11590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2107_
timestamp 0
transform -1 0 12150 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2108_
timestamp 0
transform 1 0 8890 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2109_
timestamp 0
transform 1 0 12150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2110_
timestamp 0
transform -1 0 12170 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2111_
timestamp 0
transform -1 0 12170 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2112_
timestamp 0
transform -1 0 12070 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2113_
timestamp 0
transform 1 0 11830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2114_
timestamp 0
transform 1 0 10610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2115_
timestamp 0
transform -1 0 9350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2116_
timestamp 0
transform -1 0 10230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2117_
timestamp 0
transform -1 0 10830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2118_
timestamp 0
transform -1 0 10790 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2119_
timestamp 0
transform 1 0 10690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2120_
timestamp 0
transform 1 0 10730 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2121_
timestamp 0
transform -1 0 10470 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2122_
timestamp 0
transform 1 0 10670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2123_
timestamp 0
transform -1 0 8170 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2124_
timestamp 0
transform -1 0 7870 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2125_
timestamp 0
transform -1 0 10230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2126_
timestamp 0
transform 1 0 10630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2127_
timestamp 0
transform -1 0 7050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2128_
timestamp 0
transform -1 0 9190 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2129_
timestamp 0
transform 1 0 7310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2130_
timestamp 0
transform -1 0 10930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2131_
timestamp 0
transform -1 0 7970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2132_
timestamp 0
transform 1 0 6750 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2133_
timestamp 0
transform -1 0 7050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2134_
timestamp 0
transform -1 0 7310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2135_
timestamp 0
transform -1 0 11190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2136_
timestamp 0
transform -1 0 11350 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2137_
timestamp 0
transform 1 0 11330 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2138_
timestamp 0
transform 1 0 11410 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2139_
timestamp 0
transform -1 0 11330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2140_
timestamp 0
transform -1 0 11050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2141_
timestamp 0
transform 1 0 9970 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2142_
timestamp 0
transform 1 0 10770 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2143_
timestamp 0
transform -1 0 10510 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2144_
timestamp 0
transform -1 0 11070 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2145_
timestamp 0
transform -1 0 5070 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2146_
timestamp 0
transform 1 0 9790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2147_
timestamp 0
transform 1 0 10350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2148_
timestamp 0
transform -1 0 6290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2149_
timestamp 0
transform 1 0 10070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2150_
timestamp 0
transform 1 0 8850 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2151_
timestamp 0
transform 1 0 7470 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2152_
timestamp 0
transform 1 0 8550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2153_
timestamp 0
transform 1 0 8810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2154_
timestamp 0
transform 1 0 9090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2155_
timestamp 0
transform -1 0 10170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2156_
timestamp 0
transform -1 0 10950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2157_
timestamp 0
transform 1 0 11190 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2158_
timestamp 0
transform -1 0 11770 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2159_
timestamp 0
transform -1 0 11890 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2160_
timestamp 0
transform -1 0 11430 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2161_
timestamp 0
transform 1 0 8170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2162_
timestamp 0
transform 1 0 8930 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2163_
timestamp 0
transform -1 0 10030 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2164_
timestamp 0
transform 1 0 9790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2165_
timestamp 0
transform 1 0 11030 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2166_
timestamp 0
transform 1 0 10850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2167_
timestamp 0
transform 1 0 9230 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2168_
timestamp 0
transform 1 0 10050 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2169_
timestamp 0
transform -1 0 8790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2170_
timestamp 0
transform -1 0 9210 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2171_
timestamp 0
transform 1 0 10350 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2172_
timestamp 0
transform 1 0 9770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2173_
timestamp 0
transform 1 0 9890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2174_
timestamp 0
transform -1 0 9530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2175_
timestamp 0
transform 1 0 9610 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2176_
timestamp 0
transform -1 0 9730 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2177_
timestamp 0
transform -1 0 9430 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2178_
timestamp 0
transform -1 0 11030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2179_
timestamp 0
transform 1 0 9510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2180_
timestamp 0
transform 1 0 11870 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2181_
timestamp 0
transform 1 0 11850 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2182_
timestamp 0
transform 1 0 11930 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2183_
timestamp 0
transform -1 0 11310 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2184_
timestamp 0
transform 1 0 11050 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2185_
timestamp 0
transform -1 0 10290 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2186_
timestamp 0
transform 1 0 10230 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2187_
timestamp 0
transform -1 0 10630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2188_
timestamp 0
transform 1 0 11590 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2189_
timestamp 0
transform 1 0 9970 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2190_
timestamp 0
transform 1 0 10530 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2191_
timestamp 0
transform 1 0 11150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2192_
timestamp 0
transform 1 0 11090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2193_
timestamp 0
transform -1 0 11030 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2194_
timestamp 0
transform -1 0 10590 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2195_
timestamp 0
transform -1 0 9470 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2196_
timestamp 0
transform -1 0 11110 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2197_
timestamp 0
transform 1 0 11370 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2198_
timestamp 0
transform -1 0 9910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2199_
timestamp 0
transform -1 0 9970 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2200_
timestamp 0
transform -1 0 5830 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2201_
timestamp 0
transform 1 0 6350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2202_
timestamp 0
transform 1 0 6090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2203_
timestamp 0
transform 1 0 6090 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2204_
timestamp 0
transform 1 0 6830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2205_
timestamp 0
transform 1 0 7130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2206_
timestamp 0
transform 1 0 9470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2207_
timestamp 0
transform -1 0 9970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2208_
timestamp 0
transform -1 0 9390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2209_
timestamp 0
transform 1 0 10430 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2210_
timestamp 0
transform 1 0 10430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2211_
timestamp 0
transform 1 0 11270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2212_
timestamp 0
transform -1 0 11630 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2213_
timestamp 0
transform -1 0 11670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2214_
timestamp 0
transform 1 0 11630 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2215_
timestamp 0
transform 1 0 11730 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2216_
timestamp 0
transform 1 0 12110 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2217_
timestamp 0
transform 1 0 11390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2218_
timestamp 0
transform 1 0 9670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2219_
timestamp 0
transform -1 0 9910 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2220_
timestamp 0
transform -1 0 9950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2221_
timestamp 0
transform -1 0 11890 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2222_
timestamp 0
transform 1 0 11830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2223_
timestamp 0
transform -1 0 11870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2224_
timestamp 0
transform 1 0 11850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2225_
timestamp 0
transform 1 0 10950 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2226_
timestamp 0
transform 1 0 11910 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2227_
timestamp 0
transform 1 0 11630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2228_
timestamp 0
transform -1 0 11490 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2229_
timestamp 0
transform -1 0 10570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2230_
timestamp 0
transform -1 0 10290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2231_
timestamp 0
transform -1 0 8490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2232_
timestamp 0
transform 1 0 8730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2233_
timestamp 0
transform 1 0 9510 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2234_
timestamp 0
transform -1 0 9770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2235_
timestamp 0
transform -1 0 9890 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2236_
timestamp 0
transform 1 0 7190 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2237_
timestamp 0
transform -1 0 6670 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2238_
timestamp 0
transform -1 0 6950 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2239_
timestamp 0
transform -1 0 8970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2240_
timestamp 0
transform -1 0 8690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2241_
timestamp 0
transform -1 0 8330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2242_
timestamp 0
transform -1 0 7510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2243_
timestamp 0
transform 1 0 7770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2244_
timestamp 0
transform 1 0 8050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2245_
timestamp 0
transform -1 0 7750 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2246_
timestamp 0
transform 1 0 9130 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2247_
timestamp 0
transform -1 0 12130 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2248_
timestamp 0
transform 1 0 11330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2249_
timestamp 0
transform -1 0 9490 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2250_
timestamp 0
transform 1 0 11010 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2251_
timestamp 0
transform 1 0 10570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2252_
timestamp 0
transform 1 0 11310 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2253_
timestamp 0
transform -1 0 11910 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2254_
timestamp 0
transform 1 0 12150 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2255_
timestamp 0
transform -1 0 10510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2256_
timestamp 0
transform -1 0 10790 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2257_
timestamp 0
transform 1 0 11030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2258_
timestamp 0
transform 1 0 12190 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2259_
timestamp 0
transform -1 0 11870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2260_
timestamp 0
transform 1 0 10050 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2261_
timestamp 0
transform 1 0 10310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2262_
timestamp 0
transform -1 0 10830 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2263_
timestamp 0
transform 1 0 11310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2264_
timestamp 0
transform 1 0 12130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2265_
timestamp 0
transform -1 0 11390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2266_
timestamp 0
transform -1 0 10750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2267_
timestamp 0
transform 1 0 11970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2268_
timestamp 0
transform 1 0 12130 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2269_
timestamp 0
transform -1 0 11910 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2270_
timestamp 0
transform 1 0 11330 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2271_
timestamp 0
transform -1 0 11630 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2272_
timestamp 0
transform 1 0 11890 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2273_
timestamp 0
transform -1 0 12150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2274_
timestamp 0
transform 1 0 10070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2275_
timestamp 0
transform -1 0 8230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2276_
timestamp 0
transform 1 0 8890 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2277_
timestamp 0
transform 1 0 9170 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2278_
timestamp 0
transform -1 0 9250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2279_
timestamp 0
transform 1 0 9050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2280_
timestamp 0
transform 1 0 10210 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2281_
timestamp 0
transform 1 0 12090 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2282_
timestamp 0
transform 1 0 12150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2283_
timestamp 0
transform -1 0 11030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2284_
timestamp 0
transform 1 0 12110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2285_
timestamp 0
transform 1 0 12110 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2286_
timestamp 0
transform -1 0 11890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2287_
timestamp 0
transform 1 0 11830 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2288_
timestamp 0
transform -1 0 10990 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2289_
timestamp 0
transform -1 0 10770 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2290_
timestamp 0
transform -1 0 10950 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2291_
timestamp 0
transform 1 0 11310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2292_
timestamp 0
transform 1 0 10450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2293_
timestamp 0
transform 1 0 10730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2294_
timestamp 0
transform 1 0 11050 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2295_
timestamp 0
transform 1 0 10930 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2296_
timestamp 0
transform 1 0 11190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2297_
timestamp 0
transform 1 0 11850 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2298_
timestamp 0
transform -1 0 11950 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2299_
timestamp 0
transform -1 0 10510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2300_
timestamp 0
transform 1 0 10210 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2301_
timestamp 0
transform 1 0 11830 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2302_
timestamp 0
transform 1 0 11770 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2303_
timestamp 0
transform -1 0 11750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2304_
timestamp 0
transform 1 0 11890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2305_
timestamp 0
transform 1 0 10770 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2306_
timestamp 0
transform -1 0 11630 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2307_
timestamp 0
transform 1 0 11330 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2308_
timestamp 0
transform 1 0 12110 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2309_
timestamp 0
transform -1 0 11670 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2310_
timestamp 0
transform -1 0 11610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2311_
timestamp 0
transform 1 0 11590 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2312_
timestamp 0
transform 1 0 11650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2313_
timestamp 0
transform 1 0 11930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2314_
timestamp 0
transform -1 0 11250 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2315_
timestamp 0
transform 1 0 12110 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2316_
timestamp 0
transform 1 0 11510 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2317_
timestamp 0
transform -1 0 12010 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2318_
timestamp 0
transform 1 0 11550 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2319_
timestamp 0
transform 1 0 11190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2320_
timestamp 0
transform 1 0 11610 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2321_
timestamp 0
transform 1 0 11470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2322_
timestamp 0
transform -1 0 11330 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2323_
timestamp 0
transform -1 0 11570 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2324_
timestamp 0
transform 1 0 11810 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2325_
timestamp 0
transform -1 0 12190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2326_
timestamp 0
transform 1 0 12110 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2327_
timestamp 0
transform 1 0 11470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2328_
timestamp 0
transform 1 0 11050 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2329_
timestamp 0
transform 1 0 8570 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2330_
timestamp 0
transform -1 0 10250 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2331_
timestamp 0
transform -1 0 9690 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2332_
timestamp 0
transform -1 0 11910 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2333_
timestamp 0
transform -1 0 10790 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2334_
timestamp 0
transform 1 0 10510 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2335_
timestamp 0
transform 1 0 10490 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2336_
timestamp 0
transform 1 0 10670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2337_
timestamp 0
transform -1 0 10790 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2338_
timestamp 0
transform -1 0 10710 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2339_
timestamp 0
transform -1 0 9630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2340_
timestamp 0
transform -1 0 9910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2341_
timestamp 0
transform 1 0 9610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2342_
timestamp 0
transform -1 0 10490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2343_
timestamp 0
transform -1 0 10430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2344_
timestamp 0
transform -1 0 10670 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2345_
timestamp 0
transform 1 0 11790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2346_
timestamp 0
transform 1 0 11530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2347_
timestamp 0
transform -1 0 8870 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2348_
timestamp 0
transform -1 0 9970 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2349_
timestamp 0
transform -1 0 11630 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2350_
timestamp 0
transform -1 0 11350 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2351_
timestamp 0
transform -1 0 10410 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2352_
timestamp 0
transform -1 0 10170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2353_
timestamp 0
transform -1 0 9470 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2354_
timestamp 0
transform 1 0 7870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2355_
timestamp 0
transform -1 0 6950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2356_
timestamp 0
transform -1 0 6890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2357_
timestamp 0
transform -1 0 7550 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2358_
timestamp 0
transform -1 0 7130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2359_
timestamp 0
transform 1 0 7350 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2360_
timestamp 0
transform -1 0 8030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2361_
timestamp 0
transform -1 0 7090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2362_
timestamp 0
transform 1 0 8810 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2363_
timestamp 0
transform -1 0 7490 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2364_
timestamp 0
transform 1 0 7230 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2365_
timestamp 0
transform 1 0 6950 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2366_
timestamp 0
transform 1 0 6430 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2367_
timestamp 0
transform -1 0 7270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2368_
timestamp 0
transform 1 0 6670 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2369_
timestamp 0
transform 1 0 7050 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2370_
timestamp 0
transform -1 0 7310 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2371_
timestamp 0
transform 1 0 7250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2372_
timestamp 0
transform -1 0 6830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2373_
timestamp 0
transform 1 0 6770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2374_
timestamp 0
transform 1 0 8270 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2375_
timestamp 0
transform 1 0 8330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2376_
timestamp 0
transform -1 0 6770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2377_
timestamp 0
transform 1 0 5470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2378_
timestamp 0
transform -1 0 3790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2379_
timestamp 0
transform -1 0 8050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2380_
timestamp 0
transform -1 0 5690 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2381_
timestamp 0
transform -1 0 5970 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2382_
timestamp 0
transform -1 0 5830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2383_
timestamp 0
transform 1 0 4750 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2384_
timestamp 0
transform 1 0 4670 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2385_
timestamp 0
transform 1 0 4910 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2386_
timestamp 0
transform 1 0 5190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2387_
timestamp 0
transform 1 0 1710 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2388_
timestamp 0
transform 1 0 1650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2389_
timestamp 0
transform 1 0 5230 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2390_
timestamp 0
transform 1 0 2510 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2391_
timestamp 0
transform -1 0 2310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2392_
timestamp 0
transform -1 0 2030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2393_
timestamp 0
transform -1 0 2590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2394_
timestamp 0
transform -1 0 3010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2395_
timestamp 0
transform 1 0 4410 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2396_
timestamp 0
transform 1 0 3050 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2397_
timestamp 0
transform -1 0 3130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2398_
timestamp 0
transform -1 0 2850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2399_
timestamp 0
transform 1 0 1950 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2400_
timestamp 0
transform -1 0 1390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2401_
timestamp 0
transform -1 0 2870 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2402_
timestamp 0
transform 1 0 2610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2403_
timestamp 0
transform -1 0 2250 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2404_
timestamp 0
transform -1 0 1690 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2405_
timestamp 0
transform -1 0 1550 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2406_
timestamp 0
transform 1 0 5930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2407_
timestamp 0
transform -1 0 4290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2408_
timestamp 0
transform -1 0 5650 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2409_
timestamp 0
transform -1 0 6470 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2410_
timestamp 0
transform -1 0 4250 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2411_
timestamp 0
transform -1 0 4010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2412_
timestamp 0
transform -1 0 1270 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2413_
timestamp 0
transform -1 0 4550 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2414_
timestamp 0
transform 1 0 3070 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2415_
timestamp 0
transform -1 0 2810 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2416_
timestamp 0
transform 1 0 1770 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2417_
timestamp 0
transform -1 0 2270 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2418_
timestamp 0
transform -1 0 2150 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2419_
timestamp 0
transform -1 0 3470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2420_
timestamp 0
transform 1 0 2890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2421_
timestamp 0
transform -1 0 2810 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2422_
timestamp 0
transform -1 0 1990 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2423_
timestamp 0
transform -1 0 3690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2424_
timestamp 0
transform -1 0 3530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2425_
timestamp 0
transform -1 0 3410 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2426_
timestamp 0
transform 1 0 3170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2427_
timestamp 0
transform 1 0 3330 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2428_
timestamp 0
transform -1 0 3410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2429_
timestamp 0
transform -1 0 5130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2430_
timestamp 0
transform -1 0 7830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2431_
timestamp 0
transform -1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2432_
timestamp 0
transform -1 0 9510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2433_
timestamp 0
transform 1 0 11610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2434_
timestamp 0
transform 1 0 10790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2435_
timestamp 0
transform -1 0 7270 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2436_
timestamp 0
transform -1 0 6950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2437_
timestamp 0
transform -1 0 9630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2438_
timestamp 0
transform -1 0 9370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2439_
timestamp 0
transform -1 0 6150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2440_
timestamp 0
transform 1 0 7770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2441_
timestamp 0
transform -1 0 7610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2442_
timestamp 0
transform 1 0 10310 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2443_
timestamp 0
transform -1 0 7210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2444_
timestamp 0
transform -1 0 7210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2445_
timestamp 0
transform 1 0 5310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2446_
timestamp 0
transform 1 0 6430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2447_
timestamp 0
transform -1 0 4810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2448_
timestamp 0
transform -1 0 6410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2449_
timestamp 0
transform -1 0 7030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2450_
timestamp 0
transform 1 0 4170 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2451_
timestamp 0
transform -1 0 4050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2452_
timestamp 0
transform 1 0 4690 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2453_
timestamp 0
transform 1 0 8550 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2454_
timestamp 0
transform 1 0 4430 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2455_
timestamp 0
transform 1 0 4430 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2456_
timestamp 0
transform -1 0 4290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2457_
timestamp 0
transform -1 0 4550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2458_
timestamp 0
transform -1 0 4910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2459_
timestamp 0
transform 1 0 5050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2460_
timestamp 0
transform 1 0 4930 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2461_
timestamp 0
transform 1 0 5210 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2462_
timestamp 0
transform 1 0 5350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2463_
timestamp 0
transform 1 0 6290 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2464_
timestamp 0
transform -1 0 3230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2465_
timestamp 0
transform -1 0 2950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2466_
timestamp 0
transform -1 0 2950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2467_
timestamp 0
transform 1 0 2090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2468_
timestamp 0
transform -1 0 1650 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2469_
timestamp 0
transform 1 0 610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2470_
timestamp 0
transform -1 0 2710 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2471_
timestamp 0
transform -1 0 2730 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2472_
timestamp 0
transform -1 0 2430 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2473_
timestamp 0
transform 1 0 1930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2474_
timestamp 0
transform -1 0 1450 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2475_
timestamp 0
transform -1 0 390 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2476_
timestamp 0
transform -1 0 3810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2477_
timestamp 0
transform -1 0 5050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2478_
timestamp 0
transform 1 0 3910 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2479_
timestamp 0
transform -1 0 3550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2480_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2481_
timestamp 0
transform -1 0 3350 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2482_
timestamp 0
transform 1 0 3630 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2483_
timestamp 0
transform 1 0 3050 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2484_
timestamp 0
transform 1 0 2770 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2485_
timestamp 0
transform -1 0 390 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2486_
timestamp 0
transform -1 0 2670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2487_
timestamp 0
transform 1 0 2390 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2488_
timestamp 0
transform -1 0 2390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2489_
timestamp 0
transform -1 0 1830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2490_
timestamp 0
transform -1 0 1390 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2491_
timestamp 0
transform -1 0 390 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2492_
timestamp 0
transform 1 0 4610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2493_
timestamp 0
transform 1 0 3610 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2494_
timestamp 0
transform 1 0 6190 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2495_
timestamp 0
transform 1 0 3850 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2496_
timestamp 0
transform 1 0 4150 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2497_
timestamp 0
transform -1 0 4070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2498_
timestamp 0
transform 1 0 3530 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2499_
timestamp 0
transform 1 0 3790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2500_
timestamp 0
transform -1 0 390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2501_
timestamp 0
transform -1 0 3390 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2502_
timestamp 0
transform -1 0 3030 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2503_
timestamp 0
transform -1 0 3510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__2504_
timestamp 0
transform -1 0 3270 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__2505_
timestamp 0
transform 1 0 2710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2506_
timestamp 0
transform -1 0 2530 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__2507_
timestamp 0
transform 1 0 650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2508_
timestamp 0
transform 1 0 3150 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2509_
timestamp 0
transform 1 0 2690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2510_
timestamp 0
transform -1 0 3250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2511_
timestamp 0
transform 1 0 3330 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__2512_
timestamp 0
transform 1 0 3170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2513_
timestamp 0
transform -1 0 2430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2514_
timestamp 0
transform 1 0 2130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2515_
timestamp 0
transform -1 0 2150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2516_
timestamp 0
transform -1 0 390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__2517_
timestamp 0
transform -1 0 2230 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2518_
timestamp 0
transform 1 0 5330 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2519_
timestamp 0
transform -1 0 5870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2520_
timestamp 0
transform -1 0 5970 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2521_
timestamp 0
transform 1 0 5670 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2522_
timestamp 0
transform -1 0 5670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2523_
timestamp 0
transform -1 0 5590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2524_
timestamp 0
transform -1 0 5530 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2525_
timestamp 0
transform -1 0 2750 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2526_
timestamp 0
transform 1 0 6150 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2527_
timestamp 0
transform 1 0 6550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2528_
timestamp 0
transform 1 0 6530 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2529_
timestamp 0
transform 1 0 6130 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2530_
timestamp 0
transform 1 0 5590 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2531_
timestamp 0
transform 1 0 2950 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2532_
timestamp 0
transform 1 0 4230 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2533_
timestamp 0
transform 1 0 5170 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2534_
timestamp 0
transform 1 0 4890 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2535_
timestamp 0
transform -1 0 4630 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2536_
timestamp 0
transform 1 0 3470 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2537_
timestamp 0
transform 1 0 2110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2538_
timestamp 0
transform 1 0 4510 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2539_
timestamp 0
transform 1 0 3890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2540_
timestamp 0
transform 1 0 4230 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2541_
timestamp 0
transform -1 0 4210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2542_
timestamp 0
transform -1 0 3730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2543_
timestamp 0
transform 1 0 3490 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2544_
timestamp 0
transform 1 0 4210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2545_
timestamp 0
transform 1 0 4470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2546_
timestamp 0
transform 1 0 4830 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2547_
timestamp 0
transform -1 0 4770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2548_
timestamp 0
transform -1 0 4490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2549_
timestamp 0
transform 1 0 4710 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2550_
timestamp 0
transform 1 0 4710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2551_
timestamp 0
transform 1 0 5230 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2552_
timestamp 0
transform 1 0 5470 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2553_
timestamp 0
transform 1 0 2370 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2554_
timestamp 0
transform 1 0 4510 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2555_
timestamp 0
transform -1 0 4690 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2556_
timestamp 0
transform -1 0 4930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2557_
timestamp 0
transform 1 0 4630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2558_
timestamp 0
transform 1 0 4710 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2559_
timestamp 0
transform 1 0 4430 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2560_
timestamp 0
transform 1 0 3930 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2561_
timestamp 0
transform 1 0 3630 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2562_
timestamp 0
transform 1 0 2250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2563_
timestamp 0
transform -1 0 4470 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2564_
timestamp 0
transform 1 0 4390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2565_
timestamp 0
transform -1 0 3870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2566_
timestamp 0
transform 1 0 2470 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2567_
timestamp 0
transform 1 0 3950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2568_
timestamp 0
transform -1 0 5750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2569_
timestamp 0
transform -1 0 5890 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2570_
timestamp 0
transform 1 0 5970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2571_
timestamp 0
transform 1 0 5970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2572_
timestamp 0
transform 1 0 5830 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2573_
timestamp 0
transform 1 0 5750 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2574_
timestamp 0
transform 1 0 5730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2575_
timestamp 0
transform -1 0 4770 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2576_
timestamp 0
transform -1 0 4250 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2577_
timestamp 0
transform -1 0 4510 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2578_
timestamp 0
transform 1 0 7010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2579_
timestamp 0
transform 1 0 7030 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2580_
timestamp 0
transform 1 0 8030 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2581_
timestamp 0
transform -1 0 8890 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2582_
timestamp 0
transform 1 0 6930 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2583_
timestamp 0
transform -1 0 6930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2584_
timestamp 0
transform 1 0 7350 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2585_
timestamp 0
transform 1 0 7390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2586_
timestamp 0
transform -1 0 8470 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2587_
timestamp 0
transform -1 0 6810 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2588_
timestamp 0
transform -1 0 5850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2589_
timestamp 0
transform 1 0 7470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2590_
timestamp 0
transform -1 0 6250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2591_
timestamp 0
transform 1 0 6490 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2592_
timestamp 0
transform -1 0 4470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2593_
timestamp 0
transform 1 0 4990 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2594_
timestamp 0
transform -1 0 8570 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2595_
timestamp 0
transform -1 0 5290 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2596_
timestamp 0
transform 1 0 5290 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2597_
timestamp 0
transform 1 0 5470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2598_
timestamp 0
transform -1 0 5210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2599_
timestamp 0
transform -1 0 5010 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2600_
timestamp 0
transform -1 0 5010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2601_
timestamp 0
transform -1 0 5270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2602_
timestamp 0
transform -1 0 8210 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2603_
timestamp 0
transform -1 0 6650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2604_
timestamp 0
transform -1 0 6410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2605_
timestamp 0
transform 1 0 6090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2606_
timestamp 0
transform -1 0 5590 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2607_
timestamp 0
transform 1 0 5750 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2608_
timestamp 0
transform 1 0 5570 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2609_
timestamp 0
transform -1 0 5550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2610_
timestamp 0
transform 1 0 4930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2611_
timestamp 0
transform -1 0 5190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2612_
timestamp 0
transform -1 0 5450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2613_
timestamp 0
transform -1 0 1270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2614_
timestamp 0
transform 1 0 2250 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2615_
timestamp 0
transform -1 0 2530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2616_
timestamp 0
transform -1 0 2510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2617_
timestamp 0
transform 1 0 1490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2618_
timestamp 0
transform 1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2619_
timestamp 0
transform -1 0 410 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2620_
timestamp 0
transform -1 0 650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2621_
timestamp 0
transform 1 0 970 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2622_
timestamp 0
transform 1 0 410 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2623_
timestamp 0
transform 1 0 2790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2624_
timestamp 0
transform 1 0 1990 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2625_
timestamp 0
transform -1 0 2250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2626_
timestamp 0
transform -1 0 1970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2627_
timestamp 0
transform 1 0 110 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2628_
timestamp 0
transform 1 0 110 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2629_
timestamp 0
transform -1 0 370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2630_
timestamp 0
transform 1 0 110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2631_
timestamp 0
transform 1 0 5050 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2632_
timestamp 0
transform 1 0 2290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2633_
timestamp 0
transform -1 0 2590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2634_
timestamp 0
transform -1 0 130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2635_
timestamp 0
transform 1 0 110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2636_
timestamp 0
transform 1 0 650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2637_
timestamp 0
transform 1 0 990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2638_
timestamp 0
transform 1 0 410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2639_
timestamp 0
transform -1 0 730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2640_
timestamp 0
transform -1 0 130 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2641_
timestamp 0
transform -1 0 130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2642_
timestamp 0
transform 1 0 1370 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2643_
timestamp 0
transform -1 0 1910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2644_
timestamp 0
transform 1 0 2310 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2645_
timestamp 0
transform -1 0 2050 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2646_
timestamp 0
transform -1 0 1250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2647_
timestamp 0
transform 1 0 110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2648_
timestamp 0
transform 1 0 610 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__2649_
timestamp 0
transform 1 0 110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2650_
timestamp 0
transform -1 0 3710 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2651_
timestamp 0
transform -1 0 3430 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2652_
timestamp 0
transform 1 0 650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2653_
timestamp 0
transform 1 0 370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2654_
timestamp 0
transform 1 0 1250 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2655_
timestamp 0
transform 1 0 690 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2656_
timestamp 0
transform -1 0 970 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2657_
timestamp 0
transform 1 0 110 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2658_
timestamp 0
transform 1 0 110 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2659_
timestamp 0
transform -1 0 410 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2660_
timestamp 0
transform 1 0 350 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2661_
timestamp 0
transform -1 0 2670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__2662_
timestamp 0
transform -1 0 2610 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2663_
timestamp 0
transform -1 0 2030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2664_
timestamp 0
transform 1 0 930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2665_
timestamp 0
transform -1 0 890 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2666_
timestamp 0
transform -1 0 410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2667_
timestamp 0
transform -1 0 630 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2668_
timestamp 0
transform 1 0 1130 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2669_
timestamp 0
transform -1 0 2890 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2670_
timestamp 0
transform -1 0 3010 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2671_
timestamp 0
transform 1 0 1170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2672_
timestamp 0
transform -1 0 670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2673_
timestamp 0
transform -1 0 630 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2674_
timestamp 0
transform 1 0 890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2675_
timestamp 0
transform 1 0 870 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2676_
timestamp 0
transform -1 0 1170 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2677_
timestamp 0
transform 1 0 6510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__2678_
timestamp 0
transform -1 0 6430 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2679_
timestamp 0
transform 1 0 7050 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2680_
timestamp 0
transform -1 0 6850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2681_
timestamp 0
transform 1 0 7110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2682_
timestamp 0
transform -1 0 6830 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2683_
timestamp 0
transform -1 0 1950 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2684_
timestamp 0
transform -1 0 1770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__2685_
timestamp 0
transform 1 0 1690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2686_
timestamp 0
transform 1 0 1690 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2687_
timestamp 0
transform 1 0 1430 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2688_
timestamp 0
transform -1 0 870 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2689_
timestamp 0
transform -1 0 850 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2690_
timestamp 0
transform 1 0 7350 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2691_
timestamp 0
transform -1 0 7190 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2692_
timestamp 0
transform -1 0 5130 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2693_
timestamp 0
transform -1 0 3090 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2694_
timestamp 0
transform -1 0 1390 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2695_
timestamp 0
transform -1 0 1670 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2696_
timestamp 0
transform -1 0 1390 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2697_
timestamp 0
transform 1 0 1970 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2698_
timestamp 0
transform -1 0 610 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2699_
timestamp 0
transform 1 0 6370 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2700_
timestamp 0
transform -1 0 7090 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2701_
timestamp 0
transform 1 0 7670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2702_
timestamp 0
transform 1 0 7370 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2703_
timestamp 0
transform 1 0 7530 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2704_
timestamp 0
transform -1 0 6730 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2705_
timestamp 0
transform 1 0 1650 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2706_
timestamp 0
transform 1 0 1090 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2707_
timestamp 0
transform 1 0 2790 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2708_
timestamp 0
transform 1 0 2470 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2709_
timestamp 0
transform -1 0 1150 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2710_
timestamp 0
transform -1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2711_
timestamp 0
transform -1 0 1210 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2712_
timestamp 0
transform 1 0 2950 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2713_
timestamp 0
transform -1 0 4350 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2714_
timestamp 0
transform -1 0 4770 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2715_
timestamp 0
transform 1 0 3610 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2716_
timestamp 0
transform -1 0 4370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2717_
timestamp 0
transform -1 0 5930 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__2718_
timestamp 0
transform -1 0 4170 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2719_
timestamp 0
transform 1 0 3770 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2720_
timestamp 0
transform -1 0 4070 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2721_
timestamp 0
transform -1 0 2230 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2722_
timestamp 0
transform 1 0 2350 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2723_
timestamp 0
transform 1 0 2650 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2724_
timestamp 0
transform -1 0 890 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2725_
timestamp 0
transform -1 0 5490 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2726_
timestamp 0
transform -1 0 6670 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2727_
timestamp 0
transform 1 0 3930 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2728_
timestamp 0
transform 1 0 3650 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2729_
timestamp 0
transform -1 0 3610 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2730_
timestamp 0
transform 1 0 3210 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2731_
timestamp 0
transform 1 0 2070 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2732_
timestamp 0
transform -1 0 1950 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2733_
timestamp 0
transform 1 0 1490 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2734_
timestamp 0
transform -1 0 1790 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2735_
timestamp 0
transform -1 0 3950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2736_
timestamp 0
transform -1 0 4090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2737_
timestamp 0
transform -1 0 4170 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2738_
timestamp 0
transform -1 0 3870 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2739_
timestamp 0
transform -1 0 3310 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2740_
timestamp 0
transform -1 0 3390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2741_
timestamp 0
transform -1 0 1150 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2742_
timestamp 0
transform 1 0 1450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2743_
timestamp 0
transform 1 0 1390 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2744_
timestamp 0
transform 1 0 1930 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2745_
timestamp 0
transform 1 0 590 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2746_
timestamp 0
transform 1 0 3650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2747_
timestamp 0
transform 1 0 4770 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__2748_
timestamp 0
transform 1 0 4430 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2749_
timestamp 0
transform -1 0 3590 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2750_
timestamp 0
transform -1 0 3030 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2751_
timestamp 0
transform 1 0 2870 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2752_
timestamp 0
transform 1 0 1170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2753_
timestamp 0
transform 1 0 670 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2754_
timestamp 0
transform -1 0 610 0 1 790
box -6 -8 26 268
use FILL  FILL_5__2755_
timestamp 0
transform -1 0 3130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2756_
timestamp 0
transform -1 0 2570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2757_
timestamp 0
transform 1 0 2810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2758_
timestamp 0
transform 1 0 2290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2759_
timestamp 0
transform -1 0 4370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2760_
timestamp 0
transform 1 0 3810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2761_
timestamp 0
transform 1 0 4150 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2762_
timestamp 0
transform -1 0 3890 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2763_
timestamp 0
transform -1 0 2130 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2764_
timestamp 0
transform -1 0 1850 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2765_
timestamp 0
transform -1 0 1770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2766_
timestamp 0
transform -1 0 2030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__2767_
timestamp 0
transform -1 0 1550 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__2768_
timestamp 0
transform 1 0 2210 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2769_
timestamp 0
transform 1 0 1650 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__2770_
timestamp 0
transform 1 0 6010 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2771_
timestamp 0
transform 1 0 6550 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2772_
timestamp 0
transform 1 0 4990 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__2773_
timestamp 0
transform 1 0 4190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2774_
timestamp 0
transform 1 0 2350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2775_
timestamp 0
transform 1 0 2590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2776_
timestamp 0
transform 1 0 3410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2777_
timestamp 0
transform -1 0 2890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2778_
timestamp 0
transform -1 0 3150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__2779_
timestamp 0
transform -1 0 7190 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2780_
timestamp 0
transform -1 0 7430 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__2781_
timestamp 0
transform 1 0 7910 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__2782_
timestamp 0
transform 1 0 7790 0 1 270
box -6 -8 26 268
use FILL  FILL_5__2783_
timestamp 0
transform 1 0 9730 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2784_
timestamp 0
transform 1 0 10870 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2785_
timestamp 0
transform 1 0 10250 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2786_
timestamp 0
transform 1 0 9970 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2787_
timestamp 0
transform 1 0 8430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2788_
timestamp 0
transform 1 0 8690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2789_
timestamp 0
transform 1 0 8210 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2790_
timestamp 0
transform -1 0 7950 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2791_
timestamp 0
transform 1 0 6210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2792_
timestamp 0
transform 1 0 9830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2793_
timestamp 0
transform 1 0 10030 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2794_
timestamp 0
transform -1 0 10290 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2795_
timestamp 0
transform 1 0 8470 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2796_
timestamp 0
transform 1 0 8450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2797_
timestamp 0
transform 1 0 10850 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2798_
timestamp 0
transform -1 0 9990 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2799_
timestamp 0
transform -1 0 8370 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2800_
timestamp 0
transform -1 0 7770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2801_
timestamp 0
transform 1 0 9710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2802_
timestamp 0
transform -1 0 10030 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2803_
timestamp 0
transform 1 0 8470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2804_
timestamp 0
transform -1 0 8370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2805_
timestamp 0
transform -1 0 10110 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2806_
timestamp 0
transform 1 0 9790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2807_
timestamp 0
transform -1 0 8410 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2808_
timestamp 0
transform -1 0 6650 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2809_
timestamp 0
transform 1 0 8170 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2810_
timestamp 0
transform -1 0 7590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2811_
timestamp 0
transform 1 0 10070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2812_
timestamp 0
transform 1 0 9710 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2813_
timestamp 0
transform 1 0 8290 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2814_
timestamp 0
transform -1 0 8170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2815_
timestamp 0
transform -1 0 8250 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2816_
timestamp 0
transform 1 0 9510 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2817_
timestamp 0
transform -1 0 10370 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2818_
timestamp 0
transform 1 0 11190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2819_
timestamp 0
transform 1 0 10170 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2820_
timestamp 0
transform -1 0 9950 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2821_
timestamp 0
transform -1 0 9810 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2822_
timestamp 0
transform -1 0 7530 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2823_
timestamp 0
transform -1 0 9530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2824_
timestamp 0
transform -1 0 9270 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2825_
timestamp 0
transform 1 0 8730 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2826_
timestamp 0
transform 1 0 8770 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2827_
timestamp 0
transform 1 0 9190 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2828_
timestamp 0
transform 1 0 10310 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2829_
timestamp 0
transform -1 0 9250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2830_
timestamp 0
transform 1 0 9870 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2831_
timestamp 0
transform 1 0 9050 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2832_
timestamp 0
transform -1 0 8970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2833_
timestamp 0
transform -1 0 8730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2834_
timestamp 0
transform -1 0 8310 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2835_
timestamp 0
transform -1 0 9330 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2836_
timestamp 0
transform -1 0 8030 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2837_
timestamp 0
transform 1 0 8110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2838_
timestamp 0
transform 1 0 9350 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2839_
timestamp 0
transform 1 0 9610 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2840_
timestamp 0
transform -1 0 9350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2841_
timestamp 0
transform 1 0 8250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2842_
timestamp 0
transform 1 0 11570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2843_
timestamp 0
transform -1 0 11070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2844_
timestamp 0
transform 1 0 10790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2845_
timestamp 0
transform 1 0 10530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2846_
timestamp 0
transform -1 0 10170 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2847_
timestamp 0
transform 1 0 10370 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2848_
timestamp 0
transform -1 0 9650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2849_
timestamp 0
transform 1 0 10950 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__2850_
timestamp 0
transform 1 0 11110 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2851_
timestamp 0
transform 1 0 11350 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2852_
timestamp 0
transform 1 0 12050 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2853_
timestamp 0
transform 1 0 12110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2854_
timestamp 0
transform 1 0 11790 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2855_
timestamp 0
transform 1 0 12070 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2856_
timestamp 0
transform -1 0 9110 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2857_
timestamp 0
transform 1 0 9610 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2858_
timestamp 0
transform -1 0 9910 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2859_
timestamp 0
transform 1 0 10850 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2860_
timestamp 0
transform 1 0 7730 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2861_
timestamp 0
transform 1 0 8410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2862_
timestamp 0
transform -1 0 7790 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2863_
timestamp 0
transform 1 0 7490 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2864_
timestamp 0
transform 1 0 9730 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2865_
timestamp 0
transform 1 0 8890 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2866_
timestamp 0
transform -1 0 6990 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2867_
timestamp 0
transform -1 0 8830 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2868_
timestamp 0
transform -1 0 8550 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2869_
timestamp 0
transform -1 0 8990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2870_
timestamp 0
transform 1 0 8630 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2871_
timestamp 0
transform 1 0 8590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2872_
timestamp 0
transform 1 0 5530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2873_
timestamp 0
transform -1 0 5550 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2874_
timestamp 0
transform 1 0 5470 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2875_
timestamp 0
transform -1 0 5830 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2876_
timestamp 0
transform 1 0 5510 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2877_
timestamp 0
transform 1 0 6090 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2878_
timestamp 0
transform -1 0 5830 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2879_
timestamp 0
transform -1 0 8970 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2880_
timestamp 0
transform -1 0 11970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2881_
timestamp 0
transform 1 0 11650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2882_
timestamp 0
transform -1 0 9250 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2883_
timestamp 0
transform 1 0 9050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2884_
timestamp 0
transform -1 0 9370 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2885_
timestamp 0
transform -1 0 10550 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2886_
timestamp 0
transform 1 0 10510 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2887_
timestamp 0
transform -1 0 8930 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2888_
timestamp 0
transform -1 0 9210 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2889_
timestamp 0
transform 1 0 9490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2890_
timestamp 0
transform -1 0 9850 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__2891_
timestamp 0
transform -1 0 9790 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2892_
timestamp 0
transform 1 0 9170 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2893_
timestamp 0
transform -1 0 9330 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2894_
timestamp 0
transform -1 0 11150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2895_
timestamp 0
transform 1 0 10830 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2896_
timestamp 0
transform -1 0 11110 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2897_
timestamp 0
transform -1 0 10830 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2898_
timestamp 0
transform 1 0 9450 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2899_
timestamp 0
transform -1 0 9750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2900_
timestamp 0
transform 1 0 10430 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2901_
timestamp 0
transform -1 0 10450 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2902_
timestamp 0
transform 1 0 10630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2903_
timestamp 0
transform -1 0 10750 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2904_
timestamp 0
transform -1 0 9910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2905_
timestamp 0
transform -1 0 9410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2906_
timestamp 0
transform -1 0 8570 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2907_
timestamp 0
transform -1 0 9130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2908_
timestamp 0
transform -1 0 10470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2909_
timestamp 0
transform 1 0 11830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2910_
timestamp 0
transform 1 0 10910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2911_
timestamp 0
transform 1 0 11770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2912_
timestamp 0
transform 1 0 12050 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__2913_
timestamp 0
transform 1 0 10650 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__2914_
timestamp 0
transform -1 0 7830 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2915_
timestamp 0
transform 1 0 10970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2916_
timestamp 0
transform 1 0 11210 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__2917_
timestamp 0
transform 1 0 10710 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2918_
timestamp 0
transform -1 0 10870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2919_
timestamp 0
transform 1 0 8550 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2920_
timestamp 0
transform 1 0 11250 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2921_
timestamp 0
transform 1 0 11770 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__2922_
timestamp 0
transform -1 0 11890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2923_
timestamp 0
transform 1 0 11350 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2924_
timestamp 0
transform 1 0 10270 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2925_
timestamp 0
transform 1 0 10030 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2926_
timestamp 0
transform 1 0 10170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2927_
timestamp 0
transform -1 0 10010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2928_
timestamp 0
transform -1 0 10270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__2929_
timestamp 0
transform -1 0 10390 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__2930_
timestamp 0
transform -1 0 11270 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2931_
timestamp 0
transform -1 0 11530 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__2932_
timestamp 0
transform 1 0 11490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__2933_
timestamp 0
transform 1 0 11450 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__2934_
timestamp 0
transform 1 0 11530 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__2935_
timestamp 0
transform 1 0 11610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2936_
timestamp 0
transform 1 0 10550 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__2937_
timestamp 0
transform -1 0 3550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__2938_
timestamp 0
transform -1 0 7770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2939_
timestamp 0
transform 1 0 6530 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2940_
timestamp 0
transform -1 0 6310 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2941_
timestamp 0
transform -1 0 6230 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2942_
timestamp 0
transform 1 0 5130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2943_
timestamp 0
transform -1 0 7030 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__2944_
timestamp 0
transform 1 0 5410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2945_
timestamp 0
transform -1 0 6810 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2946_
timestamp 0
transform 1 0 6410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__2947_
timestamp 0
transform 1 0 7890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2948_
timestamp 0
transform 1 0 7630 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2949_
timestamp 0
transform 1 0 5730 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__2950_
timestamp 0
transform -1 0 6070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2951_
timestamp 0
transform 1 0 6830 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2952_
timestamp 0
transform 1 0 6550 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2953_
timestamp 0
transform 1 0 5710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2954_
timestamp 0
transform -1 0 6010 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__2955_
timestamp 0
transform 1 0 7090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2956_
timestamp 0
transform 1 0 6570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__2957_
timestamp 0
transform -1 0 8190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__2958_
timestamp 0
transform 1 0 6570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__2959_
timestamp 0
transform 1 0 6310 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2960_
timestamp 0
transform -1 0 7190 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2961_
timestamp 0
transform 1 0 6570 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2962_
timestamp 0
transform -1 0 6350 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__2963_
timestamp 0
transform -1 0 6650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2964_
timestamp 0
transform 1 0 4710 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2965_
timestamp 0
transform 1 0 5770 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2966_
timestamp 0
transform -1 0 6670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__2967_
timestamp 0
transform -1 0 5090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2968_
timestamp 0
transform -1 0 5350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2969_
timestamp 0
transform 1 0 4430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2970_
timestamp 0
transform 1 0 4790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2971_
timestamp 0
transform 1 0 4670 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2972_
timestamp 0
transform -1 0 6110 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2973_
timestamp 0
transform -1 0 6370 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2974_
timestamp 0
transform -1 0 6370 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2975_
timestamp 0
transform 1 0 5830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2976_
timestamp 0
transform -1 0 4750 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2977_
timestamp 0
transform -1 0 5010 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2978_
timestamp 0
transform 1 0 5270 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__2979_
timestamp 0
transform 1 0 5550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__2980_
timestamp 0
transform -1 0 7430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2981_
timestamp 0
transform -1 0 6390 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2982_
timestamp 0
transform -1 0 6670 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__2983_
timestamp 0
transform 1 0 7190 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2984_
timestamp 0
transform 1 0 6590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__2985_
timestamp 0
transform -1 0 6930 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2986_
timestamp 0
transform 1 0 6630 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2987_
timestamp 0
transform 1 0 6070 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2988_
timestamp 0
transform -1 0 6350 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__2989_
timestamp 0
transform -1 0 7930 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2990_
timestamp 0
transform 1 0 7050 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__2991_
timestamp 0
transform -1 0 6910 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2992_
timestamp 0
transform -1 0 5210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__2993_
timestamp 0
transform -1 0 6070 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2994_
timestamp 0
transform 1 0 5530 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2995_
timestamp 0
transform 1 0 6610 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2996_
timestamp 0
transform 1 0 6330 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__2997_
timestamp 0
transform 1 0 6050 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2998_
timestamp 0
transform -1 0 5790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__2999_
timestamp 0
transform 1 0 6450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3000_
timestamp 0
transform -1 0 5790 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__3001_
timestamp 0
transform 1 0 5010 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3002_
timestamp 0
transform -1 0 5510 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__3003_
timestamp 0
transform -1 0 5870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3004_
timestamp 0
transform -1 0 5290 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3005_
timestamp 0
transform -1 0 5550 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3006_
timestamp 0
transform -1 0 7450 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3007_
timestamp 0
transform 1 0 6870 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3008_
timestamp 0
transform 1 0 8670 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3009_
timestamp 0
transform 1 0 8130 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3010_
timestamp 0
transform 1 0 7150 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3011_
timestamp 0
transform -1 0 7250 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3012_
timestamp 0
transform -1 0 7130 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3013_
timestamp 0
transform -1 0 7870 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3014_
timestamp 0
transform 1 0 7070 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3015_
timestamp 0
transform -1 0 7350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3016_
timestamp 0
transform -1 0 6110 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3017_
timestamp 0
transform -1 0 6910 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3018_
timestamp 0
transform -1 0 6590 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3019_
timestamp 0
transform -1 0 6850 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3020_
timestamp 0
transform 1 0 5490 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__3021_
timestamp 0
transform 1 0 5930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3022_
timestamp 0
transform 1 0 5730 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__3023_
timestamp 0
transform -1 0 6810 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3024_
timestamp 0
transform -1 0 6730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3025_
timestamp 0
transform 1 0 6010 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__3026_
timestamp 0
transform 1 0 5430 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__3027_
timestamp 0
transform -1 0 5530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3028_
timestamp 0
transform 1 0 6010 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3029_
timestamp 0
transform 1 0 6770 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3030_
timestamp 0
transform 1 0 4910 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__3031_
timestamp 0
transform 1 0 4450 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3032_
timestamp 0
transform -1 0 5230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3033_
timestamp 0
transform 1 0 5490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3034_
timestamp 0
transform -1 0 3430 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3035_
timestamp 0
transform -1 0 3990 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3036_
timestamp 0
transform -1 0 3490 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3037_
timestamp 0
transform -1 0 3370 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3038_
timestamp 0
transform 1 0 3590 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3039_
timestamp 0
transform -1 0 3090 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3040_
timestamp 0
transform 1 0 2970 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3041_
timestamp 0
transform 1 0 3210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3042_
timestamp 0
transform -1 0 3770 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3043_
timestamp 0
transform -1 0 3870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3044_
timestamp 0
transform -1 0 3630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3045_
timestamp 0
transform 1 0 4430 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3046_
timestamp 0
transform 1 0 4150 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3047_
timestamp 0
transform -1 0 3110 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3048_
timestamp 0
transform 1 0 3150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3049_
timestamp 0
transform -1 0 2850 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3050_
timestamp 0
transform 1 0 2890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3051_
timestamp 0
transform 1 0 2630 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3052_
timestamp 0
transform 1 0 2530 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3053_
timestamp 0
transform 1 0 3290 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3054_
timestamp 0
transform -1 0 3570 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3055_
timestamp 0
transform 1 0 3390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3056_
timestamp 0
transform -1 0 3650 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3057_
timestamp 0
transform 1 0 3850 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3058_
timestamp 0
transform 1 0 4030 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3059_
timestamp 0
transform 1 0 4310 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3060_
timestamp 0
transform 1 0 4150 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3061_
timestamp 0
transform 1 0 3630 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3062_
timestamp 0
transform -1 0 3870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3063_
timestamp 0
transform -1 0 5110 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__3064_
timestamp 0
transform 1 0 4970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__3065_
timestamp 0
transform -1 0 4710 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3066_
timestamp 0
transform 1 0 4610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3067_
timestamp 0
transform -1 0 3710 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3068_
timestamp 0
transform -1 0 3450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3069_
timestamp 0
transform 1 0 3650 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3070_
timestamp 0
transform -1 0 4550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__3071_
timestamp 0
transform 1 0 4270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__3072_
timestamp 0
transform -1 0 4210 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3073_
timestamp 0
transform -1 0 4470 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3074_
timestamp 0
transform 1 0 5750 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3075_
timestamp 0
transform 1 0 5470 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3076_
timestamp 0
transform 1 0 3710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3077_
timestamp 0
transform 1 0 4030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3078_
timestamp 0
transform 1 0 4090 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3079_
timestamp 0
transform -1 0 4170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3080_
timestamp 0
transform 1 0 6310 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3081_
timestamp 0
transform -1 0 6970 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3082_
timestamp 0
transform 1 0 6670 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3083_
timestamp 0
transform -1 0 3850 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3084_
timestamp 0
transform 1 0 3550 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3085_
timestamp 0
transform 1 0 3170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3086_
timestamp 0
transform -1 0 2890 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3087_
timestamp 0
transform 1 0 4370 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3088_
timestamp 0
transform -1 0 4970 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3089_
timestamp 0
transform 1 0 3450 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3090_
timestamp 0
transform -1 0 3730 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3091_
timestamp 0
transform -1 0 6270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3092_
timestamp 0
transform 1 0 5490 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3093_
timestamp 0
transform 1 0 5750 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3094_
timestamp 0
transform 1 0 5470 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3095_
timestamp 0
transform -1 0 4670 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3096_
timestamp 0
transform 1 0 4370 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3097_
timestamp 0
transform -1 0 4130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3098_
timestamp 0
transform 1 0 3830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3099_
timestamp 0
transform -1 0 3890 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3100_
timestamp 0
transform -1 0 3710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3101_
timestamp 0
transform 1 0 4930 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3102_
timestamp 0
transform -1 0 5230 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3103_
timestamp 0
transform -1 0 4610 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3104_
timestamp 0
transform -1 0 4890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3105_
timestamp 0
transform 1 0 5670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3106_
timestamp 0
transform -1 0 5970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3107_
timestamp 0
transform -1 0 4070 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3108_
timestamp 0
transform 1 0 3770 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3109_
timestamp 0
transform 1 0 6250 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3110_
timestamp 0
transform 1 0 3930 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3111_
timestamp 0
transform 1 0 5790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3112_
timestamp 0
transform -1 0 5210 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3113_
timestamp 0
transform -1 0 4670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3114_
timestamp 0
transform 1 0 4370 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3115_
timestamp 0
transform 1 0 4890 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3116_
timestamp 0
transform 1 0 3830 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3117_
timestamp 0
transform 1 0 4450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3118_
timestamp 0
transform -1 0 4750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3119_
timestamp 0
transform 1 0 4930 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3120_
timestamp 0
transform 1 0 4630 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3121_
timestamp 0
transform 1 0 5230 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3122_
timestamp 0
transform 1 0 5510 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3123_
timestamp 0
transform 1 0 5490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3124_
timestamp 0
transform -1 0 5790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3125_
timestamp 0
transform -1 0 4150 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3126_
timestamp 0
transform 1 0 3850 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3127_
timestamp 0
transform 1 0 6510 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3128_
timestamp 0
transform 1 0 6070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3129_
timestamp 0
transform 1 0 5470 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3130_
timestamp 0
transform -1 0 3390 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3131_
timestamp 0
transform -1 0 3630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3132_
timestamp 0
transform 1 0 4730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3133_
timestamp 0
transform 1 0 3970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3134_
timestamp 0
transform 1 0 5150 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3135_
timestamp 0
transform 1 0 4850 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3136_
timestamp 0
transform 1 0 5750 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3137_
timestamp 0
transform 1 0 5470 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3138_
timestamp 0
transform 1 0 5750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3139_
timestamp 0
transform 1 0 5470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3140_
timestamp 0
transform -1 0 5670 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3141_
timestamp 0
transform -1 0 5930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3142_
timestamp 0
transform -1 0 4270 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3143_
timestamp 0
transform -1 0 4530 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3144_
timestamp 0
transform 1 0 11610 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__3145_
timestamp 0
transform 1 0 11850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__3146_
timestamp 0
transform -1 0 11910 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__3147_
timestamp 0
transform 1 0 9530 0 1 790
box -6 -8 26 268
use FILL  FILL_5__3148_
timestamp 0
transform -1 0 11910 0 1 790
box -6 -8 26 268
use FILL  FILL_5__3149_
timestamp 0
transform -1 0 11530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3150_
timestamp 0
transform -1 0 11810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3151_
timestamp 0
transform -1 0 10750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3152_
timestamp 0
transform 1 0 9390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3153_
timestamp 0
transform -1 0 9690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3154_
timestamp 0
transform -1 0 10210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3155_
timestamp 0
transform -1 0 10330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3156_
timestamp 0
transform -1 0 8970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__3157_
timestamp 0
transform -1 0 9010 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__3158_
timestamp 0
transform -1 0 8730 0 1 2870
box -6 -8 26 268
use FILL  FILL_5__3159_
timestamp 0
transform -1 0 8710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__3160_
timestamp 0
transform 1 0 10550 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3161_
timestamp 0
transform 1 0 10270 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3162_
timestamp 0
transform -1 0 9810 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3163_
timestamp 0
transform 1 0 9530 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3164_
timestamp 0
transform -1 0 9010 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3165_
timestamp 0
transform -1 0 7230 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3166_
timestamp 0
transform 1 0 7630 0 1 1310
box -6 -8 26 268
use FILL  FILL_5__3167_
timestamp 0
transform 1 0 7490 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3168_
timestamp 0
transform 1 0 7650 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3169_
timestamp 0
transform -1 0 8730 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3170_
timestamp 0
transform -1 0 8450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3171_
timestamp 0
transform -1 0 9170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3172_
timestamp 0
transform -1 0 8170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3173_
timestamp 0
transform 1 0 8430 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3174_
timestamp 0
transform 1 0 7910 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3175_
timestamp 0
transform -1 0 7890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3176_
timestamp 0
transform -1 0 7610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3177_
timestamp 0
transform -1 0 11890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__3178_
timestamp 0
transform -1 0 11830 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3179_
timestamp 0
transform 1 0 12090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3180_
timestamp 0
transform 1 0 12150 0 1 790
box -6 -8 26 268
use FILL  FILL_5__3181_
timestamp 0
transform 1 0 12130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__3182_
timestamp 0
transform -1 0 11350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3183_
timestamp 0
transform 1 0 11610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3184_
timestamp 0
transform 1 0 11890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3185_
timestamp 0
transform 1 0 11910 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3186_
timestamp 0
transform 1 0 12090 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3187_
timestamp 0
transform 1 0 9950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5__3188_
timestamp 0
transform 1 0 10830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3189_
timestamp 0
transform -1 0 11090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_5__3190_
timestamp 0
transform 1 0 11130 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3191_
timestamp 0
transform 1 0 11070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3192_
timestamp 0
transform -1 0 10790 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3193_
timestamp 0
transform 1 0 10210 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3194_
timestamp 0
transform 1 0 10830 0 1 2350
box -6 -8 26 268
use FILL  FILL_5__3195_
timestamp 0
transform -1 0 10570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3196_
timestamp 0
transform 1 0 10470 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3197_
timestamp 0
transform -1 0 7330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3198_
timestamp 0
transform -1 0 4690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3199_
timestamp 0
transform 1 0 2850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5__3200_
timestamp 0
transform 1 0 4830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__3201_
timestamp 0
transform 1 0 4550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__3202_
timestamp 0
transform 1 0 1610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5__3203_
timestamp 0
transform 1 0 1570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3204_
timestamp 0
transform 1 0 1530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__3205_
timestamp 0
transform 1 0 1090 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__3206_
timestamp 0
transform 1 0 1510 0 1 3390
box -6 -8 26 268
use FILL  FILL_5__3207_
timestamp 0
transform -1 0 1650 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__3208_
timestamp 0
transform -1 0 990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__3209_
timestamp 0
transform -1 0 690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__3210_
timestamp 0
transform -1 0 4350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__3211_
timestamp 0
transform 1 0 4290 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__3212_
timestamp 0
transform 1 0 1250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5__3213_
timestamp 0
transform 1 0 1150 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__3214_
timestamp 0
transform -1 0 2430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3215_
timestamp 0
transform 1 0 1850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3216_
timestamp 0
transform 1 0 5790 0 1 270
box -6 -8 26 268
use FILL  FILL_5__3217_
timestamp 0
transform -1 0 6090 0 1 270
box -6 -8 26 268
use FILL  FILL_5__3218_
timestamp 0
transform 1 0 6130 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3219_
timestamp 0
transform -1 0 6410 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3220_
timestamp 0
transform 1 0 3750 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3221_
timestamp 0
transform -1 0 4030 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3222_
timestamp 0
transform -1 0 3630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3223_
timestamp 0
transform 1 0 3350 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__3224_
timestamp 0
transform -1 0 3330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3225_
timestamp 0
transform 1 0 5470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__3226_
timestamp 0
transform 1 0 5190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__3227_
timestamp 0
transform -1 0 4310 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3228_
timestamp 0
transform -1 0 4510 0 1 270
box -6 -8 26 268
use FILL  FILL_5__3229_
timestamp 0
transform 1 0 2750 0 1 1830
box -6 -8 26 268
use FILL  FILL_5__3230_
timestamp 0
transform -1 0 2790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5__3231_
timestamp 0
transform 1 0 6030 0 1 790
box -6 -8 26 268
use FILL  FILL_5__3232_
timestamp 0
transform 1 0 6010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5__3364_
timestamp 0
transform 1 0 5290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3365_
timestamp 0
transform 1 0 4490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3366_
timestamp 0
transform 1 0 4970 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__3367_
timestamp 0
transform -1 0 4770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3368_
timestamp 0
transform -1 0 5030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3369_
timestamp 0
transform -1 0 5590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3370_
timestamp 0
transform 1 0 2730 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3371_
timestamp 0
transform 1 0 2230 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3372_
timestamp 0
transform -1 0 2350 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3373_
timestamp 0
transform -1 0 4010 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3374_
timestamp 0
transform -1 0 2330 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3375_
timestamp 0
transform 1 0 2330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3376_
timestamp 0
transform -1 0 2990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3377_
timestamp 0
transform 1 0 2450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3378_
timestamp 0
transform -1 0 2310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3379_
timestamp 0
transform -1 0 1470 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3380_
timestamp 0
transform 1 0 1250 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3381_
timestamp 0
transform -1 0 1510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3382_
timestamp 0
transform -1 0 1970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3383_
timestamp 0
transform -1 0 1530 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3384_
timestamp 0
transform 1 0 1790 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3385_
timestamp 0
transform 1 0 1490 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3386_
timestamp 0
transform -1 0 2070 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3387_
timestamp 0
transform 1 0 2330 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3388_
timestamp 0
transform -1 0 670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3389_
timestamp 0
transform 1 0 2530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3390_
timestamp 0
transform 1 0 3350 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3391_
timestamp 0
transform 1 0 3070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3392_
timestamp 0
transform -1 0 2910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3393_
timestamp 0
transform 1 0 2310 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3394_
timestamp 0
transform 1 0 710 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3395_
timestamp 0
transform -1 0 670 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3396_
timestamp 0
transform -1 0 410 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3397_
timestamp 0
transform -1 0 430 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3398_
timestamp 0
transform -1 0 130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3399_
timestamp 0
transform 1 0 110 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3400_
timestamp 0
transform -1 0 910 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3401_
timestamp 0
transform -1 0 1490 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3402_
timestamp 0
transform 1 0 1470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3403_
timestamp 0
transform 1 0 1190 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3404_
timestamp 0
transform -1 0 130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3405_
timestamp 0
transform -1 0 390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3406_
timestamp 0
transform -1 0 130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3407_
timestamp 0
transform -1 0 410 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3408_
timestamp 0
transform -1 0 130 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3409_
timestamp 0
transform -1 0 130 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3410_
timestamp 0
transform 1 0 1450 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3411_
timestamp 0
transform 1 0 1170 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3412_
timestamp 0
transform -1 0 650 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3413_
timestamp 0
transform 1 0 390 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3414_
timestamp 0
transform 1 0 650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5__3415_
timestamp 0
transform -1 0 970 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3416_
timestamp 0
transform 1 0 650 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3417_
timestamp 0
transform -1 0 690 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3418_
timestamp 0
transform -1 0 390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3419_
timestamp 0
transform -1 0 1210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3420_
timestamp 0
transform 1 0 910 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3421_
timestamp 0
transform 1 0 1210 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3422_
timestamp 0
transform 1 0 930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3423_
timestamp 0
transform 1 0 1230 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3424_
timestamp 0
transform -1 0 1250 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3425_
timestamp 0
transform -1 0 970 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3426_
timestamp 0
transform 1 0 950 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5__3427_
timestamp 0
transform -1 0 1470 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3428_
timestamp 0
transform 1 0 1150 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3429_
timestamp 0
transform -1 0 930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3430_
timestamp 0
transform 1 0 1450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3431_
timestamp 0
transform 1 0 1170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3432_
timestamp 0
transform -1 0 970 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3433_
timestamp 0
transform -1 0 130 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3434_
timestamp 0
transform -1 0 710 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3435_
timestamp 0
transform -1 0 990 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3436_
timestamp 0
transform -1 0 930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3437_
timestamp 0
transform 1 0 1750 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3438_
timestamp 0
transform 1 0 1210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3439_
timestamp 0
transform -1 0 1490 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3440_
timestamp 0
transform 1 0 1210 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3441_
timestamp 0
transform -1 0 650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3442_
timestamp 0
transform 1 0 1230 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3443_
timestamp 0
transform 1 0 1150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3444_
timestamp 0
transform -1 0 2050 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3445_
timestamp 0
transform 1 0 1730 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3446_
timestamp 0
transform 1 0 2090 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3447_
timestamp 0
transform 1 0 1990 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3448_
timestamp 0
transform -1 0 1790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3449_
timestamp 0
transform 1 0 1470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3450_
timestamp 0
transform -1 0 930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3451_
timestamp 0
transform 1 0 1190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3452_
timestamp 0
transform 1 0 890 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3453_
timestamp 0
transform -1 0 2210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3454_
timestamp 0
transform 1 0 3130 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3455_
timestamp 0
transform -1 0 2070 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3456_
timestamp 0
transform -1 0 1730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3457_
timestamp 0
transform -1 0 2910 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3458_
timestamp 0
transform -1 0 1770 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3459_
timestamp 0
transform -1 0 1710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3460_
timestamp 0
transform 1 0 1750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3461_
timestamp 0
transform -1 0 1970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3462_
timestamp 0
transform -1 0 1730 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3463_
timestamp 0
transform -1 0 1490 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3464_
timestamp 0
transform 1 0 1210 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3465_
timestamp 0
transform -1 0 1470 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3466_
timestamp 0
transform 1 0 2010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3467_
timestamp 0
transform 1 0 2010 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3468_
timestamp 0
transform 1 0 2770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3469_
timestamp 0
transform 1 0 2630 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3470_
timestamp 0
transform -1 0 2530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3471_
timestamp 0
transform 1 0 2350 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3472_
timestamp 0
transform -1 0 2250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3473_
timestamp 0
transform 1 0 1490 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3474_
timestamp 0
transform -1 0 1750 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3475_
timestamp 0
transform 1 0 1230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3476_
timestamp 0
transform -1 0 970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3477_
timestamp 0
transform 1 0 390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3478_
timestamp 0
transform -1 0 370 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3479_
timestamp 0
transform -1 0 130 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3480_
timestamp 0
transform -1 0 130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3481_
timestamp 0
transform -1 0 130 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3482_
timestamp 0
transform 1 0 650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3483_
timestamp 0
transform -1 0 370 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3484_
timestamp 0
transform 1 0 1990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3485_
timestamp 0
transform -1 0 2050 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3486_
timestamp 0
transform -1 0 1430 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3487_
timestamp 0
transform -1 0 1750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3488_
timestamp 0
transform -1 0 1550 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3489_
timestamp 0
transform 1 0 1490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3490_
timestamp 0
transform 1 0 1170 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3491_
timestamp 0
transform -1 0 1250 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3492_
timestamp 0
transform 1 0 1150 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3493_
timestamp 0
transform -1 0 970 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3494_
timestamp 0
transform 1 0 890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3495_
timestamp 0
transform -1 0 650 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3496_
timestamp 0
transform 1 0 410 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3497_
timestamp 0
transform -1 0 370 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3498_
timestamp 0
transform 1 0 670 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3499_
timestamp 0
transform -1 0 730 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3500_
timestamp 0
transform 1 0 670 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3501_
timestamp 0
transform 1 0 910 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3502_
timestamp 0
transform -1 0 430 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3503_
timestamp 0
transform -1 0 410 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3504_
timestamp 0
transform -1 0 650 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3505_
timestamp 0
transform -1 0 410 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3506_
timestamp 0
transform -1 0 130 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3507_
timestamp 0
transform -1 0 130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3508_
timestamp 0
transform 1 0 650 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3509_
timestamp 0
transform -1 0 910 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3510_
timestamp 0
transform -1 0 410 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3511_
timestamp 0
transform -1 0 130 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3512_
timestamp 0
transform 1 0 610 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3513_
timestamp 0
transform -1 0 430 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3514_
timestamp 0
transform -1 0 370 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3515_
timestamp 0
transform -1 0 130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3516_
timestamp 0
transform -1 0 130 0 1 10150
box -6 -8 26 268
use FILL  FILL_5__3517_
timestamp 0
transform 1 0 670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3518_
timestamp 0
transform 1 0 890 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3519_
timestamp 0
transform 1 0 2590 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3520_
timestamp 0
transform 1 0 2870 0 1 9110
box -6 -8 26 268
use FILL  FILL_5__3521_
timestamp 0
transform 1 0 3350 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3522_
timestamp 0
transform 1 0 3050 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3523_
timestamp 0
transform 1 0 2610 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3524_
timestamp 0
transform -1 0 990 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3525_
timestamp 0
transform -1 0 130 0 1 10670
box -6 -8 26 268
use FILL  FILL_5__3526_
timestamp 0
transform -1 0 130 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3527_
timestamp 0
transform -1 0 630 0 1 11190
box -6 -8 26 268
use FILL  FILL_5__3528_
timestamp 0
transform -1 0 650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_5__3529_
timestamp 0
transform -1 0 130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5__3530_
timestamp 0
transform -1 0 130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3531_
timestamp 0
transform 1 0 110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3532_
timestamp 0
transform 1 0 350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3533_
timestamp 0
transform -1 0 130 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3534_
timestamp 0
transform -1 0 650 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3535_
timestamp 0
transform -1 0 410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5__3536_
timestamp 0
transform -1 0 390 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3537_
timestamp 0
transform -1 0 1750 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3538_
timestamp 0
transform 1 0 2510 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3539_
timestamp 0
transform -1 0 2610 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3540_
timestamp 0
transform -1 0 2350 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3541_
timestamp 0
transform -1 0 2070 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3542_
timestamp 0
transform -1 0 2250 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3543_
timestamp 0
transform 1 0 1650 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3544_
timestamp 0
transform 1 0 2010 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3545_
timestamp 0
transform 1 0 1810 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3546_
timestamp 0
transform 1 0 1930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5__3547_
timestamp 0
transform -1 0 2590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3548_
timestamp 0
transform 1 0 2290 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5__3549_
timestamp 0
transform -1 0 2390 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3550_
timestamp 0
transform 1 0 2090 0 1 11710
box -6 -8 26 268
use FILL  FILL_5__3551_
timestamp 0
transform -1 0 2570 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3552_
timestamp 0
transform 1 0 2270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5__3553_
timestamp 0
transform -1 0 1810 0 1 8070
box -6 -8 26 268
use FILL  FILL_5__3554_
timestamp 0
transform 1 0 950 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3555_
timestamp 0
transform 1 0 350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3556_
timestamp 0
transform 1 0 1210 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5__3557_
timestamp 0
transform -1 0 3110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3558_
timestamp 0
transform 1 0 2810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5__3559_
timestamp 0
transform -1 0 2570 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3560_
timestamp 0
transform 1 0 2270 0 1 9630
box -6 -8 26 268
use FILL  FILL_5__3561_
timestamp 0
transform -1 0 1990 0 1 7550
box -6 -8 26 268
use FILL  FILL_5__3562_
timestamp 0
transform -1 0 2810 0 1 8590
box -6 -8 26 268
use FILL  FILL_5__3563_
timestamp 0
transform 1 0 2210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5__3564_
timestamp 0
transform 1 0 2490 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3565_
timestamp 0
transform -1 0 1490 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3566_
timestamp 0
transform -1 0 1750 0 1 7030
box -6 -8 26 268
use FILL  FILL_5__3579_
timestamp 0
transform -1 0 5090 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3580_
timestamp 0
transform -1 0 130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5__3581_
timestamp 0
transform -1 0 3510 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3582_
timestamp 0
transform -1 0 3250 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3583_
timestamp 0
transform -1 0 5370 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__3584_
timestamp 0
transform 1 0 4550 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3585_
timestamp 0
transform 1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3586_
timestamp 0
transform -1 0 5890 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__3587_
timestamp 0
transform 1 0 110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3588_
timestamp 0
transform -1 0 130 0 1 3910
box -6 -8 26 268
use FILL  FILL_5__3589_
timestamp 0
transform -1 0 130 0 1 4950
box -6 -8 26 268
use FILL  FILL_5__3590_
timestamp 0
transform -1 0 130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5__3591_
timestamp 0
transform -1 0 410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3592_
timestamp 0
transform -1 0 130 0 1 4430
box -6 -8 26 268
use FILL  FILL_5__3593_
timestamp 0
transform -1 0 4830 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3594_
timestamp 0
transform 1 0 5870 0 -1 270
box -6 -8 26 268
use FILL  FILL_5__3595_
timestamp 0
transform 1 0 5610 0 -1 790
box -6 -8 26 268
use FILL  FILL_5__3596_
timestamp 0
transform -1 0 910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3597_
timestamp 0
transform -1 0 130 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__3598_
timestamp 0
transform -1 0 390 0 1 5990
box -6 -8 26 268
use FILL  FILL_5__3599_
timestamp 0
transform -1 0 130 0 1 6510
box -6 -8 26 268
use FILL  FILL_5__3600_
timestamp 0
transform -1 0 130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5__3601_
timestamp 0
transform -1 0 130 0 1 5470
box -6 -8 26 268
use FILL  FILL_5__3602_
timestamp 0
transform -1 0 1750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5__3603_
timestamp 0
transform 1 0 6910 0 -1 270
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert0
timestamp 0
transform 1 0 7930 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert1
timestamp 0
transform 1 0 9430 0 1 1830
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert2
timestamp 0
transform 1 0 8190 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert3
timestamp 0
transform 1 0 11050 0 1 1830
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert4
timestamp 0
transform 1 0 650 0 1 1830
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert5
timestamp 0
transform -1 0 12130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert6
timestamp 0
transform -1 0 9630 0 1 5470
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert7
timestamp 0
transform 1 0 7090 0 1 2350
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert8
timestamp 0
transform -1 0 910 0 1 5470
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert9
timestamp 0
transform 1 0 10170 0 1 3910
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert10
timestamp 0
transform -1 0 950 0 1 5990
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert11
timestamp 0
transform -1 0 6030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert12
timestamp 0
transform 1 0 11590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert13
timestamp 0
transform -1 0 6210 0 1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert14
timestamp 0
transform 1 0 6830 0 1 2350
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert15
timestamp 0
transform -1 0 3370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert16
timestamp 0
transform -1 0 3990 0 1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert17
timestamp 0
transform 1 0 7230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert18
timestamp 0
transform -1 0 7050 0 1 11190
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert19
timestamp 0
transform 1 0 5370 0 1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert20
timestamp 0
transform 1 0 8610 0 1 11190
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert21
timestamp 0
transform -1 0 8530 0 -1 7550
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert22
timestamp 0
transform -1 0 1490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert23
timestamp 0
transform 1 0 3470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert24
timestamp 0
transform -1 0 4370 0 1 5470
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert25
timestamp 0
transform 1 0 8210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert26
timestamp 0
transform 1 0 5150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert27
timestamp 0
transform -1 0 1290 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert39
timestamp 0
transform 1 0 6370 0 1 4950
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert40
timestamp 0
transform 1 0 7730 0 1 3910
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert41
timestamp 0
transform -1 0 8870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert42
timestamp 0
transform -1 0 7010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert43
timestamp 0
transform -1 0 8910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert44
timestamp 0
transform -1 0 9030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert45
timestamp 0
transform 1 0 11090 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert46
timestamp 0
transform 1 0 9530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert47
timestamp 0
transform 1 0 9250 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert48
timestamp 0
transform 1 0 6990 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert49
timestamp 0
transform 1 0 7250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert50
timestamp 0
transform -1 0 7630 0 1 9110
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert51
timestamp 0
transform 1 0 7590 0 1 10150
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert52
timestamp 0
transform 1 0 8990 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert53
timestamp 0
transform 1 0 10030 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert54
timestamp 0
transform 1 0 8870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert55
timestamp 0
transform 1 0 8730 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert56
timestamp 0
transform -1 0 2270 0 1 8590
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert57
timestamp 0
transform 1 0 2570 0 1 11190
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert58
timestamp 0
transform 1 0 2710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert59
timestamp 0
transform -1 0 2270 0 1 10670
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert60
timestamp 0
transform -1 0 10530 0 1 7550
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert61
timestamp 0
transform 1 0 10590 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert62
timestamp 0
transform 1 0 10550 0 1 8070
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert63
timestamp 0
transform -1 0 9210 0 1 7550
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert64
timestamp 0
transform -1 0 8650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert65
timestamp 0
transform 1 0 5250 0 1 270
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert66
timestamp 0
transform 1 0 5770 0 1 790
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert67
timestamp 0
transform -1 0 3070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert68
timestamp 0
transform 1 0 3190 0 1 270
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert69
timestamp 0
transform -1 0 6690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert70
timestamp 0
transform 1 0 8630 0 1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert71
timestamp 0
transform -1 0 9290 0 1 2870
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert72
timestamp 0
transform -1 0 6810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert73
timestamp 0
transform 1 0 8970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert74
timestamp 0
transform 1 0 10830 0 1 7030
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert75
timestamp 0
transform 1 0 2610 0 1 1310
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert76
timestamp 0
transform -1 0 3110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert77
timestamp 0
transform 1 0 10490 0 1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert78
timestamp 0
transform 1 0 9350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert79
timestamp 0
transform -1 0 8390 0 1 7550
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert80
timestamp 0
transform 1 0 7190 0 1 5470
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert81
timestamp 0
transform 1 0 7650 0 -1 790
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert82
timestamp 0
transform -1 0 7630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert83
timestamp 0
transform -1 0 7410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert84
timestamp 0
transform 1 0 9470 0 1 8590
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert85
timestamp 0
transform -1 0 8950 0 1 8590
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert86
timestamp 0
transform -1 0 9550 0 1 2870
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert87
timestamp 0
transform 1 0 9450 0 1 4430
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert88
timestamp 0
transform -1 0 10790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert89
timestamp 0
transform 1 0 9430 0 1 3390
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert90
timestamp 0
transform 1 0 5410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert91
timestamp 0
transform -1 0 4950 0 1 10670
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert92
timestamp 0
transform -1 0 4790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert93
timestamp 0
transform 1 0 5210 0 1 10150
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert94
timestamp 0
transform -1 0 11370 0 1 9630
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert95
timestamp 0
transform -1 0 11410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert96
timestamp 0
transform -1 0 10130 0 1 11710
box -6 -8 26 268
use FILL  FILL_5_BUFX2_insert97
timestamp 0
transform 1 0 11490 0 1 11710
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert28
timestamp 0
transform -1 0 6070 0 -1 11710
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert29
timestamp 0
transform -1 0 2250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert30
timestamp 0
transform 1 0 4590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert31
timestamp 0
transform -1 0 3290 0 1 2870
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert32
timestamp 0
transform 1 0 7190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert33
timestamp 0
transform 1 0 5770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert34
timestamp 0
transform -1 0 2530 0 1 10670
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert35
timestamp 0
transform -1 0 5290 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert36
timestamp 0
transform -1 0 2410 0 1 3910
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert37
timestamp 0
transform 1 0 7430 0 -1 12230
box -6 -8 26 268
use FILL  FILL_5_CLKBUF1_insert38
timestamp 0
transform -1 0 4410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__1688_
timestamp 0
transform -1 0 950 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1689_
timestamp 0
transform -1 0 410 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1690_
timestamp 0
transform -1 0 670 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1691_
timestamp 0
transform 1 0 130 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1692_
timestamp 0
transform -1 0 390 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1693_
timestamp 0
transform 1 0 630 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1694_
timestamp 0
transform -1 0 5630 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__1695_
timestamp 0
transform -1 0 410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1696_
timestamp 0
transform -1 0 410 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1697_
timestamp 0
transform -1 0 1530 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__1698_
timestamp 0
transform -1 0 3470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1699_
timestamp 0
transform 1 0 2910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1700_
timestamp 0
transform -1 0 3950 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__1701_
timestamp 0
transform -1 0 650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1702_
timestamp 0
transform -1 0 650 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1703_
timestamp 0
transform 1 0 3290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1704_
timestamp 0
transform -1 0 430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1705_
timestamp 0
transform 1 0 130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1706_
timestamp 0
transform -1 0 3910 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1707_
timestamp 0
transform -1 0 670 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1708_
timestamp 0
transform 1 0 670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1709_
timestamp 0
transform 1 0 4190 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1710_
timestamp 0
transform -1 0 5670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1711_
timestamp 0
transform 1 0 5210 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1712_
timestamp 0
transform 1 0 7350 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1713_
timestamp 0
transform -1 0 9730 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1714_
timestamp 0
transform -1 0 9930 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1715_
timestamp 0
transform -1 0 8610 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1716_
timestamp 0
transform 1 0 11370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1717_
timestamp 0
transform 1 0 11170 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1718_
timestamp 0
transform 1 0 11990 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1719_
timestamp 0
transform -1 0 8870 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1720_
timestamp 0
transform -1 0 10190 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1721_
timestamp 0
transform -1 0 10210 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1722_
timestamp 0
transform -1 0 9970 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1723_
timestamp 0
transform 1 0 10070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1724_
timestamp 0
transform 1 0 9290 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1725_
timestamp 0
transform 1 0 9130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1726_
timestamp 0
transform 1 0 10230 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1727_
timestamp 0
transform -1 0 8850 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1728_
timestamp 0
transform 1 0 11630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1729_
timestamp 0
transform 1 0 10230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1730_
timestamp 0
transform 1 0 8410 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1731_
timestamp 0
transform 1 0 8650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1732_
timestamp 0
transform -1 0 7850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1733_
timestamp 0
transform 1 0 9790 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1734_
timestamp 0
transform 1 0 7490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1735_
timestamp 0
transform 1 0 10930 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1736_
timestamp 0
transform -1 0 10730 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1737_
timestamp 0
transform -1 0 10990 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1738_
timestamp 0
transform -1 0 10370 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1739_
timestamp 0
transform -1 0 10370 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1740_
timestamp 0
transform 1 0 10590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1741_
timestamp 0
transform -1 0 8490 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1742_
timestamp 0
transform -1 0 8390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1743_
timestamp 0
transform -1 0 9950 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1744_
timestamp 0
transform 1 0 9830 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1745_
timestamp 0
transform -1 0 9530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1746_
timestamp 0
transform 1 0 11390 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1747_
timestamp 0
transform 1 0 10870 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1748_
timestamp 0
transform 1 0 7590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1749_
timestamp 0
transform 1 0 8010 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__1750_
timestamp 0
transform -1 0 8130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1751_
timestamp 0
transform 1 0 7530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1752_
timestamp 0
transform -1 0 8950 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1753_
timestamp 0
transform 1 0 9810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1754_
timestamp 0
transform -1 0 8350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1755_
timestamp 0
transform -1 0 8930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__1756_
timestamp 0
transform -1 0 11270 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1757_
timestamp 0
transform 1 0 11130 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1758_
timestamp 0
transform -1 0 9190 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1759_
timestamp 0
transform -1 0 7430 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__1760_
timestamp 0
transform 1 0 8930 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__1761_
timestamp 0
transform -1 0 9650 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1762_
timestamp 0
transform 1 0 10670 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1763_
timestamp 0
transform -1 0 9110 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1764_
timestamp 0
transform 1 0 11370 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1765_
timestamp 0
transform 1 0 8190 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1766_
timestamp 0
transform 1 0 8570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1767_
timestamp 0
transform 1 0 9270 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__1768_
timestamp 0
transform 1 0 8130 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__1769_
timestamp 0
transform 1 0 8650 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__1770_
timestamp 0
transform 1 0 9090 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__1771_
timestamp 0
transform 1 0 9050 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__1772_
timestamp 0
transform 1 0 8770 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__1773_
timestamp 0
transform 1 0 10850 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1774_
timestamp 0
transform 1 0 10850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1775_
timestamp 0
transform 1 0 10090 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1776_
timestamp 0
transform -1 0 8090 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1777_
timestamp 0
transform 1 0 8130 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1778_
timestamp 0
transform -1 0 7610 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1779_
timestamp 0
transform 1 0 5750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1780_
timestamp 0
transform -1 0 4150 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1781_
timestamp 0
transform -1 0 10870 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1782_
timestamp 0
transform 1 0 8350 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1783_
timestamp 0
transform 1 0 10590 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1784_
timestamp 0
transform -1 0 10070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1785_
timestamp 0
transform -1 0 9830 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1786_
timestamp 0
transform 1 0 10250 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1787_
timestamp 0
transform -1 0 9190 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1788_
timestamp 0
transform -1 0 8610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1789_
timestamp 0
transform 1 0 10050 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1790_
timestamp 0
transform -1 0 10110 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1791_
timestamp 0
transform -1 0 10190 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1792_
timestamp 0
transform -1 0 9730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1793_
timestamp 0
transform -1 0 9470 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1794_
timestamp 0
transform 1 0 9190 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1795_
timestamp 0
transform -1 0 8390 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1796_
timestamp 0
transform -1 0 8330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1797_
timestamp 0
transform 1 0 7170 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1798_
timestamp 0
transform 1 0 7430 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1799_
timestamp 0
transform -1 0 9450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1800_
timestamp 0
transform 1 0 11330 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1801_
timestamp 0
transform 1 0 9350 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1802_
timestamp 0
transform -1 0 9010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1803_
timestamp 0
transform 1 0 10610 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1804_
timestamp 0
transform -1 0 8630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1805_
timestamp 0
transform -1 0 8730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1806_
timestamp 0
transform 1 0 7670 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1807_
timestamp 0
transform -1 0 8130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1808_
timestamp 0
transform -1 0 8450 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1809_
timestamp 0
transform 1 0 8670 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1810_
timestamp 0
transform 1 0 8070 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1811_
timestamp 0
transform -1 0 7810 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1812_
timestamp 0
transform -1 0 8450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1813_
timestamp 0
transform -1 0 8170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1814_
timestamp 0
transform -1 0 7910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1815_
timestamp 0
transform 1 0 7930 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1816_
timestamp 0
transform -1 0 3930 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1817_
timestamp 0
transform 1 0 1410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1818_
timestamp 0
transform -1 0 6230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1819_
timestamp 0
transform -1 0 990 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1820_
timestamp 0
transform 1 0 430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1821_
timestamp 0
transform 1 0 950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1822_
timestamp 0
transform -1 0 410 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1823_
timestamp 0
transform 1 0 1770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1824_
timestamp 0
transform 1 0 1350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__1825_
timestamp 0
transform -1 0 1190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1826_
timestamp 0
transform -1 0 450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1827_
timestamp 0
transform 1 0 950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1828_
timestamp 0
transform -1 0 1550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1829_
timestamp 0
transform -1 0 690 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1830_
timestamp 0
transform -1 0 1490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1831_
timestamp 0
transform 1 0 2070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1832_
timestamp 0
transform -1 0 8070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1833_
timestamp 0
transform 1 0 9710 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1834_
timestamp 0
transform 1 0 9290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1835_
timestamp 0
transform -1 0 7810 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1836_
timestamp 0
transform -1 0 6470 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1837_
timestamp 0
transform -1 0 7810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1838_
timestamp 0
transform -1 0 7250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1839_
timestamp 0
transform -1 0 6230 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1840_
timestamp 0
transform 1 0 8610 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1841_
timestamp 0
transform -1 0 8230 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1842_
timestamp 0
transform -1 0 6990 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1843_
timestamp 0
transform -1 0 6710 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1844_
timestamp 0
transform 1 0 9130 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1845_
timestamp 0
transform 1 0 9670 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1846_
timestamp 0
transform -1 0 9270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1847_
timestamp 0
transform -1 0 8430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1848_
timestamp 0
transform 1 0 11270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1849_
timestamp 0
transform -1 0 11590 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1850_
timestamp 0
transform -1 0 11050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1851_
timestamp 0
transform 1 0 10410 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1852_
timestamp 0
transform -1 0 10470 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1853_
timestamp 0
transform -1 0 10490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__1854_
timestamp 0
transform -1 0 7470 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1855_
timestamp 0
transform 1 0 7450 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1856_
timestamp 0
transform 1 0 7730 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1857_
timestamp 0
transform -1 0 8870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__1858_
timestamp 0
transform -1 0 9410 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1859_
timestamp 0
transform -1 0 8870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1860_
timestamp 0
transform 1 0 9130 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1861_
timestamp 0
transform 1 0 6870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1862_
timestamp 0
transform -1 0 8370 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__1863_
timestamp 0
transform 1 0 7730 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1864_
timestamp 0
transform -1 0 6370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1865_
timestamp 0
transform -1 0 7810 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__1866_
timestamp 0
transform -1 0 7270 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1867_
timestamp 0
transform -1 0 8050 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1868_
timestamp 0
transform 1 0 7770 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1869_
timestamp 0
transform -1 0 6070 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__1870_
timestamp 0
transform 1 0 9410 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1871_
timestamp 0
transform 1 0 8890 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1872_
timestamp 0
transform -1 0 8630 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1873_
timestamp 0
transform -1 0 7830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1874_
timestamp 0
transform -1 0 7550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1875_
timestamp 0
transform -1 0 8350 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1876_
timestamp 0
transform -1 0 6990 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1877_
timestamp 0
transform -1 0 5830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__1878_
timestamp 0
transform 1 0 6710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1879_
timestamp 0
transform -1 0 7510 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1880_
timestamp 0
transform 1 0 6030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__1881_
timestamp 0
transform 1 0 6030 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__1882_
timestamp 0
transform -1 0 4990 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__1883_
timestamp 0
transform -1 0 7890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1884_
timestamp 0
transform -1 0 8130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1885_
timestamp 0
transform -1 0 8690 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__1886_
timestamp 0
transform 1 0 8530 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1887_
timestamp 0
transform -1 0 8510 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1888_
timestamp 0
transform 1 0 11650 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1889_
timestamp 0
transform -1 0 8510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1890_
timestamp 0
transform 1 0 9770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1891_
timestamp 0
transform 1 0 8930 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1892_
timestamp 0
transform -1 0 8650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1893_
timestamp 0
transform 1 0 12170 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1894_
timestamp 0
transform 1 0 12150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1895_
timestamp 0
transform 1 0 12170 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1896_
timestamp 0
transform -1 0 10790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1897_
timestamp 0
transform -1 0 9190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1898_
timestamp 0
transform 1 0 9070 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1899_
timestamp 0
transform 1 0 7510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1900_
timestamp 0
transform 1 0 9710 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1901_
timestamp 0
transform 1 0 8050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1902_
timestamp 0
transform -1 0 8270 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1903_
timestamp 0
transform 1 0 7990 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1904_
timestamp 0
transform 1 0 11910 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1905_
timestamp 0
transform 1 0 11670 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1906_
timestamp 0
transform -1 0 6550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1907_
timestamp 0
transform -1 0 7090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1908_
timestamp 0
transform -1 0 7010 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1909_
timestamp 0
transform -1 0 6770 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__1910_
timestamp 0
transform -1 0 6270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1911_
timestamp 0
transform 1 0 6850 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1912_
timestamp 0
transform 1 0 6310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__1913_
timestamp 0
transform 1 0 6250 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1914_
timestamp 0
transform 1 0 5750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1915_
timestamp 0
transform 1 0 5270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1916_
timestamp 0
transform 1 0 5270 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__1917_
timestamp 0
transform -1 0 3770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__1918_
timestamp 0
transform 1 0 3650 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__1919_
timestamp 0
transform -1 0 3930 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__1920_
timestamp 0
transform -1 0 3650 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__1921_
timestamp 0
transform -1 0 1770 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__1922_
timestamp 0
transform 1 0 7570 0 1 270
box -6 -8 26 268
use FILL  FILL_6__1923_
timestamp 0
transform 1 0 7830 0 1 790
box -6 -8 26 268
use FILL  FILL_6__1924_
timestamp 0
transform -1 0 6430 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__1925_
timestamp 0
transform -1 0 4670 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1926_
timestamp 0
transform -1 0 4030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1927_
timestamp 0
transform 1 0 2070 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__1928_
timestamp 0
transform -1 0 3230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__1929_
timestamp 0
transform 1 0 4610 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__1930_
timestamp 0
transform 1 0 3170 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__1931_
timestamp 0
transform -1 0 2950 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__1932_
timestamp 0
transform -1 0 1550 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1933_
timestamp 0
transform -1 0 8510 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1934_
timestamp 0
transform 1 0 3910 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__1935_
timestamp 0
transform -1 0 3930 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1936_
timestamp 0
transform -1 0 2610 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1937_
timestamp 0
transform -1 0 1270 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1938_
timestamp 0
transform -1 0 3630 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1939_
timestamp 0
transform -1 0 4190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1940_
timestamp 0
transform -1 0 3410 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1941_
timestamp 0
transform -1 0 3350 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1942_
timestamp 0
transform -1 0 1850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__1943_
timestamp 0
transform -1 0 3650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__1944_
timestamp 0
transform -1 0 3750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1945_
timestamp 0
transform -1 0 3010 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__1946_
timestamp 0
transform -1 0 1570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__1947_
timestamp 0
transform -1 0 4990 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__1948_
timestamp 0
transform 1 0 5190 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__1949_
timestamp 0
transform 1 0 5250 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__1950_
timestamp 0
transform -1 0 4990 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__1951_
timestamp 0
transform -1 0 2030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1952_
timestamp 0
transform 1 0 4150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__1953_
timestamp 0
transform 1 0 4090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__1954_
timestamp 0
transform 1 0 4230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1955_
timestamp 0
transform -1 0 1750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1956_
timestamp 0
transform -1 0 4370 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__1957_
timestamp 0
transform 1 0 4950 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__1958_
timestamp 0
transform -1 0 5230 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__1959_
timestamp 0
transform -1 0 4210 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__1960_
timestamp 0
transform -1 0 2370 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1961_
timestamp 0
transform 1 0 4190 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1962_
timestamp 0
transform 1 0 3950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1963_
timestamp 0
transform 1 0 3730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1964_
timestamp 0
transform 1 0 2070 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1965_
timestamp 0
transform 1 0 6450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__1966_
timestamp 0
transform 1 0 6390 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1967_
timestamp 0
transform 1 0 7230 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1968_
timestamp 0
transform 1 0 6690 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1969_
timestamp 0
transform -1 0 3350 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__1970_
timestamp 0
transform 1 0 2890 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1971_
timestamp 0
transform -1 0 4770 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1972_
timestamp 0
transform 1 0 3630 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1973_
timestamp 0
transform -1 0 3650 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__1974_
timestamp 0
transform -1 0 3150 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__1975_
timestamp 0
transform 1 0 3050 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__1976_
timestamp 0
transform -1 0 3150 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__1977_
timestamp 0
transform 1 0 4430 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__1978_
timestamp 0
transform 1 0 3130 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__1979_
timestamp 0
transform -1 0 2870 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__1980_
timestamp 0
transform -1 0 2390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1981_
timestamp 0
transform 1 0 6010 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__1982_
timestamp 0
transform 1 0 6130 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__1983_
timestamp 0
transform 1 0 6330 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__1984_
timestamp 0
transform 1 0 5330 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__1985_
timestamp 0
transform -1 0 4830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1986_
timestamp 0
transform 1 0 2610 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__1987_
timestamp 0
transform -1 0 7330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__1988_
timestamp 0
transform 1 0 7630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__1989_
timestamp 0
transform 1 0 7690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__1990_
timestamp 0
transform -1 0 7490 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1991_
timestamp 0
transform -1 0 7770 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__1992_
timestamp 0
transform 1 0 10510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__1993_
timestamp 0
transform 1 0 9630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__1994_
timestamp 0
transform -1 0 6310 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__1995_
timestamp 0
transform 1 0 6690 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__1996_
timestamp 0
transform -1 0 6830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1997_
timestamp 0
transform 1 0 6530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__1998_
timestamp 0
transform 1 0 6530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__1999_
timestamp 0
transform 1 0 7590 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2000_
timestamp 0
transform 1 0 6510 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2001_
timestamp 0
transform 1 0 6750 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2002_
timestamp 0
transform 1 0 6710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2003_
timestamp 0
transform 1 0 9590 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2004_
timestamp 0
transform 1 0 7530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2005_
timestamp 0
transform -1 0 7330 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2006_
timestamp 0
transform 1 0 6810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2007_
timestamp 0
transform 1 0 6650 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2008_
timestamp 0
transform -1 0 6290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2009_
timestamp 0
transform 1 0 6890 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2010_
timestamp 0
transform -1 0 7110 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2011_
timestamp 0
transform 1 0 7350 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2012_
timestamp 0
transform -1 0 9490 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2013_
timestamp 0
transform 1 0 10630 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2014_
timestamp 0
transform -1 0 10890 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2015_
timestamp 0
transform -1 0 6330 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2016_
timestamp 0
transform -1 0 7370 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2017_
timestamp 0
transform -1 0 7150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2018_
timestamp 0
transform 1 0 7390 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2019_
timestamp 0
transform 1 0 9470 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2020_
timestamp 0
transform -1 0 10370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2021_
timestamp 0
transform -1 0 7410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2022_
timestamp 0
transform 1 0 7650 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2023_
timestamp 0
transform -1 0 7950 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2024_
timestamp 0
transform 1 0 6170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2025_
timestamp 0
transform -1 0 6050 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2026_
timestamp 0
transform 1 0 9750 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2027_
timestamp 0
transform 1 0 10290 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2028_
timestamp 0
transform -1 0 10290 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2029_
timestamp 0
transform -1 0 11170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2030_
timestamp 0
transform 1 0 10790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2031_
timestamp 0
transform -1 0 11090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2032_
timestamp 0
transform 1 0 9010 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2033_
timestamp 0
transform 1 0 8470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2034_
timestamp 0
transform 1 0 8710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2035_
timestamp 0
transform 1 0 8670 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2036_
timestamp 0
transform 1 0 11630 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2037_
timestamp 0
transform 1 0 11830 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2038_
timestamp 0
transform -1 0 7670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2039_
timestamp 0
transform -1 0 6750 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2040_
timestamp 0
transform 1 0 11010 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2041_
timestamp 0
transform 1 0 11090 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2042_
timestamp 0
transform -1 0 10170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2043_
timestamp 0
transform -1 0 10550 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2044_
timestamp 0
transform -1 0 11070 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2045_
timestamp 0
transform -1 0 11410 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2046_
timestamp 0
transform 1 0 8890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2047_
timestamp 0
transform -1 0 9450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2048_
timestamp 0
transform 1 0 9250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2049_
timestamp 0
transform 1 0 9390 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2050_
timestamp 0
transform 1 0 9150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2051_
timestamp 0
transform 1 0 8850 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2052_
timestamp 0
transform 1 0 9130 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2053_
timestamp 0
transform -1 0 9690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2054_
timestamp 0
transform 1 0 9910 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2055_
timestamp 0
transform -1 0 6550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2056_
timestamp 0
transform -1 0 6130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2057_
timestamp 0
transform 1 0 10330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2058_
timestamp 0
transform -1 0 10070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2059_
timestamp 0
transform -1 0 10210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2060_
timestamp 0
transform -1 0 9970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2061_
timestamp 0
transform 1 0 10150 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2062_
timestamp 0
transform -1 0 9230 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2063_
timestamp 0
transform 1 0 8310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2064_
timestamp 0
transform -1 0 7990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2065_
timestamp 0
transform -1 0 8810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2066_
timestamp 0
transform 1 0 8790 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2067_
timestamp 0
transform -1 0 8050 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2068_
timestamp 0
transform -1 0 8330 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2069_
timestamp 0
transform 1 0 8050 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2070_
timestamp 0
transform -1 0 8350 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2071_
timestamp 0
transform -1 0 8630 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2072_
timestamp 0
transform 1 0 8850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2073_
timestamp 0
transform 1 0 9110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2074_
timestamp 0
transform 1 0 9330 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2075_
timestamp 0
transform -1 0 9630 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2076_
timestamp 0
transform 1 0 11290 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2077_
timestamp 0
transform -1 0 11350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2078_
timestamp 0
transform -1 0 11150 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2079_
timestamp 0
transform 1 0 11290 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2080_
timestamp 0
transform -1 0 11130 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2081_
timestamp 0
transform 1 0 11130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2082_
timestamp 0
transform 1 0 10390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2083_
timestamp 0
transform 1 0 9650 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2084_
timestamp 0
transform 1 0 11670 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2085_
timestamp 0
transform 1 0 11090 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2086_
timestamp 0
transform 1 0 11590 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2087_
timestamp 0
transform 1 0 11610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2088_
timestamp 0
transform -1 0 12170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2089_
timestamp 0
transform 1 0 11890 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2090_
timestamp 0
transform 1 0 12070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2091_
timestamp 0
transform 1 0 9970 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2092_
timestamp 0
transform 1 0 10590 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2093_
timestamp 0
transform -1 0 11150 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2094_
timestamp 0
transform 1 0 11390 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2095_
timestamp 0
transform -1 0 11050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2096_
timestamp 0
transform 1 0 11570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2097_
timestamp 0
transform -1 0 11910 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2098_
timestamp 0
transform -1 0 12090 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2099_
timestamp 0
transform -1 0 11390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2100_
timestamp 0
transform 1 0 11350 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2101_
timestamp 0
transform -1 0 11310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2102_
timestamp 0
transform -1 0 11690 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2103_
timestamp 0
transform 1 0 12170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2104_
timestamp 0
transform 1 0 12170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2105_
timestamp 0
transform -1 0 11630 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2106_
timestamp 0
transform -1 0 11610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2107_
timestamp 0
transform -1 0 12170 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2108_
timestamp 0
transform 1 0 8910 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2109_
timestamp 0
transform 1 0 12170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2110_
timestamp 0
transform -1 0 12190 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2111_
timestamp 0
transform -1 0 12190 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2112_
timestamp 0
transform -1 0 12090 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2113_
timestamp 0
transform 1 0 11850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2114_
timestamp 0
transform 1 0 10630 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2115_
timestamp 0
transform -1 0 9370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2116_
timestamp 0
transform -1 0 10250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2117_
timestamp 0
transform -1 0 10850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2118_
timestamp 0
transform -1 0 10810 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2119_
timestamp 0
transform 1 0 10710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2120_
timestamp 0
transform 1 0 10750 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2121_
timestamp 0
transform -1 0 10490 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2122_
timestamp 0
transform 1 0 10690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2123_
timestamp 0
transform -1 0 8190 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2124_
timestamp 0
transform -1 0 7890 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2125_
timestamp 0
transform -1 0 10250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2126_
timestamp 0
transform 1 0 10650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2127_
timestamp 0
transform -1 0 7070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2128_
timestamp 0
transform -1 0 9210 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2129_
timestamp 0
transform 1 0 7330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2130_
timestamp 0
transform -1 0 10950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2131_
timestamp 0
transform -1 0 7990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2132_
timestamp 0
transform 1 0 6770 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2133_
timestamp 0
transform -1 0 7070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2134_
timestamp 0
transform -1 0 7330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2135_
timestamp 0
transform -1 0 11210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2136_
timestamp 0
transform -1 0 11370 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2137_
timestamp 0
transform 1 0 11350 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2138_
timestamp 0
transform 1 0 11430 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2139_
timestamp 0
transform -1 0 11350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2140_
timestamp 0
transform -1 0 11070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2141_
timestamp 0
transform 1 0 9990 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2142_
timestamp 0
transform 1 0 10790 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2143_
timestamp 0
transform -1 0 10530 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2144_
timestamp 0
transform -1 0 11090 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2145_
timestamp 0
transform -1 0 5090 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2146_
timestamp 0
transform 1 0 9810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2147_
timestamp 0
transform 1 0 10370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2148_
timestamp 0
transform -1 0 6310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2149_
timestamp 0
transform 1 0 10090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2150_
timestamp 0
transform 1 0 8870 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2151_
timestamp 0
transform 1 0 7490 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2152_
timestamp 0
transform 1 0 8570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2153_
timestamp 0
transform 1 0 8830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2154_
timestamp 0
transform 1 0 9110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2155_
timestamp 0
transform -1 0 10190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2156_
timestamp 0
transform -1 0 10970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2157_
timestamp 0
transform 1 0 11210 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2158_
timestamp 0
transform -1 0 11790 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2159_
timestamp 0
transform -1 0 11910 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2160_
timestamp 0
transform -1 0 11450 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2161_
timestamp 0
transform 1 0 8190 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2162_
timestamp 0
transform 1 0 8950 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2163_
timestamp 0
transform -1 0 10050 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2164_
timestamp 0
transform 1 0 9810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2165_
timestamp 0
transform 1 0 11050 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2166_
timestamp 0
transform 1 0 10870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2167_
timestamp 0
transform 1 0 9250 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2168_
timestamp 0
transform 1 0 10070 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2169_
timestamp 0
transform -1 0 8810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2170_
timestamp 0
transform -1 0 9230 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2171_
timestamp 0
transform 1 0 10370 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2172_
timestamp 0
transform 1 0 9790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2173_
timestamp 0
transform 1 0 9910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2174_
timestamp 0
transform -1 0 9550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2175_
timestamp 0
transform 1 0 9630 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2176_
timestamp 0
transform -1 0 9750 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2177_
timestamp 0
transform -1 0 9450 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2178_
timestamp 0
transform -1 0 11050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2179_
timestamp 0
transform 1 0 9530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2180_
timestamp 0
transform 1 0 11890 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2181_
timestamp 0
transform 1 0 11870 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2182_
timestamp 0
transform 1 0 11950 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2183_
timestamp 0
transform -1 0 11330 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2184_
timestamp 0
transform 1 0 11070 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2185_
timestamp 0
transform -1 0 10310 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2186_
timestamp 0
transform 1 0 10250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2187_
timestamp 0
transform -1 0 10650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2188_
timestamp 0
transform 1 0 11610 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2189_
timestamp 0
transform 1 0 9990 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2190_
timestamp 0
transform 1 0 10550 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2191_
timestamp 0
transform 1 0 11170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2192_
timestamp 0
transform 1 0 11110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2193_
timestamp 0
transform -1 0 11050 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2194_
timestamp 0
transform -1 0 10610 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2195_
timestamp 0
transform -1 0 9490 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2196_
timestamp 0
transform -1 0 11130 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2197_
timestamp 0
transform 1 0 11390 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2198_
timestamp 0
transform -1 0 9930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2199_
timestamp 0
transform -1 0 9990 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2200_
timestamp 0
transform -1 0 5850 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2201_
timestamp 0
transform 1 0 6370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2202_
timestamp 0
transform 1 0 6110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2203_
timestamp 0
transform 1 0 6110 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2204_
timestamp 0
transform 1 0 6850 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2205_
timestamp 0
transform 1 0 7150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2206_
timestamp 0
transform 1 0 9490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2207_
timestamp 0
transform -1 0 9990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2208_
timestamp 0
transform -1 0 9410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2209_
timestamp 0
transform 1 0 10450 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2210_
timestamp 0
transform 1 0 10450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2211_
timestamp 0
transform 1 0 11290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2212_
timestamp 0
transform -1 0 11650 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2213_
timestamp 0
transform -1 0 11690 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2214_
timestamp 0
transform 1 0 11650 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2215_
timestamp 0
transform 1 0 11750 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2216_
timestamp 0
transform 1 0 12130 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2217_
timestamp 0
transform 1 0 11410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2218_
timestamp 0
transform 1 0 9690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2219_
timestamp 0
transform -1 0 9930 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2220_
timestamp 0
transform -1 0 9970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2221_
timestamp 0
transform -1 0 11910 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2222_
timestamp 0
transform 1 0 11850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2223_
timestamp 0
transform -1 0 11890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2224_
timestamp 0
transform 1 0 11870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2225_
timestamp 0
transform 1 0 10970 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2226_
timestamp 0
transform 1 0 11930 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2227_
timestamp 0
transform 1 0 11650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2228_
timestamp 0
transform -1 0 11510 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2229_
timestamp 0
transform -1 0 10590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2230_
timestamp 0
transform -1 0 10310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2231_
timestamp 0
transform -1 0 8510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2232_
timestamp 0
transform 1 0 8750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2233_
timestamp 0
transform 1 0 9530 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2234_
timestamp 0
transform -1 0 9790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2235_
timestamp 0
transform -1 0 9910 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2236_
timestamp 0
transform 1 0 7210 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2237_
timestamp 0
transform -1 0 6690 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2238_
timestamp 0
transform -1 0 6970 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2239_
timestamp 0
transform -1 0 8990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2240_
timestamp 0
transform -1 0 8710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2241_
timestamp 0
transform -1 0 8350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2242_
timestamp 0
transform -1 0 7530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2243_
timestamp 0
transform 1 0 7790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2244_
timestamp 0
transform 1 0 8070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2245_
timestamp 0
transform -1 0 7770 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2246_
timestamp 0
transform 1 0 9150 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2247_
timestamp 0
transform -1 0 12150 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2248_
timestamp 0
transform 1 0 11350 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2249_
timestamp 0
transform -1 0 9510 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2250_
timestamp 0
transform 1 0 11030 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2251_
timestamp 0
transform 1 0 10590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2252_
timestamp 0
transform 1 0 11330 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2253_
timestamp 0
transform -1 0 11930 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2254_
timestamp 0
transform 1 0 12170 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2255_
timestamp 0
transform -1 0 10530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2256_
timestamp 0
transform -1 0 10810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2257_
timestamp 0
transform 1 0 11050 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2258_
timestamp 0
transform 1 0 12210 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2259_
timestamp 0
transform -1 0 11890 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2260_
timestamp 0
transform 1 0 10070 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2261_
timestamp 0
transform 1 0 10330 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2262_
timestamp 0
transform -1 0 10850 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2263_
timestamp 0
transform 1 0 11330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2264_
timestamp 0
transform 1 0 12150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2265_
timestamp 0
transform -1 0 11410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2266_
timestamp 0
transform -1 0 10770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2267_
timestamp 0
transform 1 0 11990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2268_
timestamp 0
transform 1 0 12150 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2269_
timestamp 0
transform -1 0 11930 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2270_
timestamp 0
transform 1 0 11350 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2271_
timestamp 0
transform -1 0 11650 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2272_
timestamp 0
transform 1 0 11910 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2273_
timestamp 0
transform -1 0 12170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2274_
timestamp 0
transform 1 0 10090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2275_
timestamp 0
transform -1 0 8250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2276_
timestamp 0
transform 1 0 8910 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2277_
timestamp 0
transform 1 0 9190 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2278_
timestamp 0
transform -1 0 9270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2279_
timestamp 0
transform 1 0 9070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2280_
timestamp 0
transform 1 0 10230 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2281_
timestamp 0
transform 1 0 12110 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2282_
timestamp 0
transform 1 0 12170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2283_
timestamp 0
transform -1 0 11050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2284_
timestamp 0
transform 1 0 12130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2285_
timestamp 0
transform 1 0 12130 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2286_
timestamp 0
transform -1 0 11910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2287_
timestamp 0
transform 1 0 11850 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2288_
timestamp 0
transform -1 0 11010 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2289_
timestamp 0
transform -1 0 10790 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2290_
timestamp 0
transform -1 0 10970 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2291_
timestamp 0
transform 1 0 11330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2292_
timestamp 0
transform 1 0 10470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2293_
timestamp 0
transform 1 0 10750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2294_
timestamp 0
transform 1 0 11070 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2295_
timestamp 0
transform 1 0 10950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2296_
timestamp 0
transform 1 0 11210 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2297_
timestamp 0
transform 1 0 11870 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2298_
timestamp 0
transform -1 0 11970 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2299_
timestamp 0
transform -1 0 10530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2300_
timestamp 0
transform 1 0 10230 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2301_
timestamp 0
transform 1 0 11850 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2302_
timestamp 0
transform 1 0 11790 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2303_
timestamp 0
transform -1 0 11770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2304_
timestamp 0
transform 1 0 11910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2305_
timestamp 0
transform 1 0 10790 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2306_
timestamp 0
transform -1 0 11650 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2307_
timestamp 0
transform 1 0 11350 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2308_
timestamp 0
transform 1 0 12130 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2309_
timestamp 0
transform -1 0 11690 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2310_
timestamp 0
transform -1 0 11630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2311_
timestamp 0
transform 1 0 11610 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2312_
timestamp 0
transform 1 0 11670 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2313_
timestamp 0
transform 1 0 11950 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2314_
timestamp 0
transform -1 0 11270 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2315_
timestamp 0
transform 1 0 12130 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2316_
timestamp 0
transform 1 0 11530 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2317_
timestamp 0
transform -1 0 12030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2318_
timestamp 0
transform 1 0 11570 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2319_
timestamp 0
transform 1 0 11210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2320_
timestamp 0
transform 1 0 11630 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2321_
timestamp 0
transform 1 0 11490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2322_
timestamp 0
transform -1 0 11350 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2323_
timestamp 0
transform -1 0 11590 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2324_
timestamp 0
transform 1 0 11830 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2325_
timestamp 0
transform -1 0 12210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2326_
timestamp 0
transform 1 0 12130 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2327_
timestamp 0
transform 1 0 11490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2328_
timestamp 0
transform 1 0 11070 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2329_
timestamp 0
transform 1 0 8590 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2330_
timestamp 0
transform -1 0 10270 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2331_
timestamp 0
transform -1 0 9710 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2332_
timestamp 0
transform -1 0 11930 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2333_
timestamp 0
transform -1 0 10810 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2334_
timestamp 0
transform 1 0 10530 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2335_
timestamp 0
transform 1 0 10510 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2336_
timestamp 0
transform 1 0 10690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2337_
timestamp 0
transform -1 0 10810 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2338_
timestamp 0
transform -1 0 10730 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2339_
timestamp 0
transform -1 0 9650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2340_
timestamp 0
transform -1 0 9930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2341_
timestamp 0
transform 1 0 9630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2342_
timestamp 0
transform -1 0 10510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2343_
timestamp 0
transform -1 0 10450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2344_
timestamp 0
transform -1 0 10690 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2345_
timestamp 0
transform 1 0 11810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2346_
timestamp 0
transform 1 0 11550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2347_
timestamp 0
transform -1 0 8890 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2348_
timestamp 0
transform -1 0 9990 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2349_
timestamp 0
transform -1 0 11650 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2350_
timestamp 0
transform -1 0 11370 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2351_
timestamp 0
transform -1 0 10430 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2352_
timestamp 0
transform -1 0 10190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2353_
timestamp 0
transform -1 0 9490 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2354_
timestamp 0
transform 1 0 7890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2355_
timestamp 0
transform -1 0 6970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2356_
timestamp 0
transform -1 0 6910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2357_
timestamp 0
transform -1 0 7570 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2358_
timestamp 0
transform -1 0 7150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2359_
timestamp 0
transform 1 0 7370 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2360_
timestamp 0
transform -1 0 8050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2361_
timestamp 0
transform -1 0 7110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2362_
timestamp 0
transform 1 0 8830 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2363_
timestamp 0
transform -1 0 7510 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2364_
timestamp 0
transform 1 0 7250 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2365_
timestamp 0
transform 1 0 6970 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2366_
timestamp 0
transform 1 0 6450 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2367_
timestamp 0
transform -1 0 7290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2368_
timestamp 0
transform 1 0 6690 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2369_
timestamp 0
transform 1 0 7070 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2370_
timestamp 0
transform -1 0 7330 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2371_
timestamp 0
transform 1 0 7270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2372_
timestamp 0
transform -1 0 6850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2373_
timestamp 0
transform 1 0 6790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2374_
timestamp 0
transform 1 0 8290 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2375_
timestamp 0
transform 1 0 8350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2376_
timestamp 0
transform -1 0 6790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2377_
timestamp 0
transform 1 0 5490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2378_
timestamp 0
transform -1 0 3810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2379_
timestamp 0
transform -1 0 8070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2380_
timestamp 0
transform -1 0 5710 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2381_
timestamp 0
transform -1 0 5990 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2382_
timestamp 0
transform -1 0 5850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2383_
timestamp 0
transform 1 0 4770 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2384_
timestamp 0
transform 1 0 4690 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2385_
timestamp 0
transform 1 0 4930 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2386_
timestamp 0
transform 1 0 5210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2387_
timestamp 0
transform 1 0 1730 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2388_
timestamp 0
transform 1 0 1670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2389_
timestamp 0
transform 1 0 5250 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2390_
timestamp 0
transform 1 0 2530 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2391_
timestamp 0
transform -1 0 2330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2392_
timestamp 0
transform -1 0 2050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2393_
timestamp 0
transform -1 0 2610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2394_
timestamp 0
transform -1 0 3030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2395_
timestamp 0
transform 1 0 4430 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2396_
timestamp 0
transform 1 0 3070 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2397_
timestamp 0
transform -1 0 3150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2398_
timestamp 0
transform -1 0 2870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2399_
timestamp 0
transform 1 0 1970 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2400_
timestamp 0
transform -1 0 1410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2401_
timestamp 0
transform -1 0 2890 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2402_
timestamp 0
transform 1 0 2630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2403_
timestamp 0
transform -1 0 2270 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2404_
timestamp 0
transform -1 0 1710 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2405_
timestamp 0
transform -1 0 1570 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2406_
timestamp 0
transform 1 0 5950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2407_
timestamp 0
transform -1 0 4310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2408_
timestamp 0
transform -1 0 5670 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2409_
timestamp 0
transform -1 0 6490 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2410_
timestamp 0
transform -1 0 4270 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2411_
timestamp 0
transform -1 0 4030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2412_
timestamp 0
transform -1 0 1290 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2413_
timestamp 0
transform -1 0 4570 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2414_
timestamp 0
transform 1 0 3090 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2415_
timestamp 0
transform -1 0 2830 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2416_
timestamp 0
transform 1 0 1790 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2417_
timestamp 0
transform -1 0 2290 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2418_
timestamp 0
transform -1 0 2170 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2419_
timestamp 0
transform -1 0 3490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2420_
timestamp 0
transform 1 0 2910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2421_
timestamp 0
transform -1 0 2830 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2422_
timestamp 0
transform -1 0 2010 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2423_
timestamp 0
transform -1 0 3710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2424_
timestamp 0
transform -1 0 3550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2425_
timestamp 0
transform -1 0 3430 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2426_
timestamp 0
transform 1 0 3190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2427_
timestamp 0
transform 1 0 3350 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2428_
timestamp 0
transform -1 0 3430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2429_
timestamp 0
transform -1 0 5150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2430_
timestamp 0
transform -1 0 7850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2431_
timestamp 0
transform -1 0 5410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2432_
timestamp 0
transform -1 0 9530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2433_
timestamp 0
transform 1 0 11630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2434_
timestamp 0
transform 1 0 10810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2435_
timestamp 0
transform -1 0 7290 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2436_
timestamp 0
transform -1 0 6970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2437_
timestamp 0
transform -1 0 9650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2438_
timestamp 0
transform -1 0 9390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2439_
timestamp 0
transform -1 0 6170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2440_
timestamp 0
transform 1 0 7790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2441_
timestamp 0
transform -1 0 7630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2442_
timestamp 0
transform 1 0 10330 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2443_
timestamp 0
transform -1 0 7230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2444_
timestamp 0
transform -1 0 7230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2445_
timestamp 0
transform 1 0 5330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2446_
timestamp 0
transform 1 0 6450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2447_
timestamp 0
transform -1 0 4830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2448_
timestamp 0
transform -1 0 6430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2449_
timestamp 0
transform -1 0 7050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2450_
timestamp 0
transform 1 0 4190 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2451_
timestamp 0
transform -1 0 4070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2452_
timestamp 0
transform 1 0 4710 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2453_
timestamp 0
transform 1 0 8570 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2454_
timestamp 0
transform 1 0 4450 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2455_
timestamp 0
transform 1 0 4450 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2456_
timestamp 0
transform -1 0 4310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2457_
timestamp 0
transform -1 0 4570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2458_
timestamp 0
transform -1 0 4930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2459_
timestamp 0
transform 1 0 5070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2460_
timestamp 0
transform 1 0 4950 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2461_
timestamp 0
transform 1 0 5230 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2462_
timestamp 0
transform 1 0 5370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2463_
timestamp 0
transform 1 0 6310 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2464_
timestamp 0
transform -1 0 3250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2465_
timestamp 0
transform -1 0 2970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2466_
timestamp 0
transform -1 0 2970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2467_
timestamp 0
transform 1 0 2110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2468_
timestamp 0
transform -1 0 1670 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2469_
timestamp 0
transform 1 0 630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2470_
timestamp 0
transform -1 0 2730 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2471_
timestamp 0
transform -1 0 2750 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2472_
timestamp 0
transform -1 0 2450 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2473_
timestamp 0
transform 1 0 1950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2474_
timestamp 0
transform -1 0 1470 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2475_
timestamp 0
transform -1 0 410 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2476_
timestamp 0
transform -1 0 3830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2477_
timestamp 0
transform -1 0 5070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2478_
timestamp 0
transform 1 0 3930 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2479_
timestamp 0
transform -1 0 3570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2480_
timestamp 0
transform 1 0 1810 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2481_
timestamp 0
transform -1 0 3370 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2482_
timestamp 0
transform 1 0 3650 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2483_
timestamp 0
transform 1 0 3070 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2484_
timestamp 0
transform 1 0 2790 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2485_
timestamp 0
transform -1 0 410 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2486_
timestamp 0
transform -1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2487_
timestamp 0
transform 1 0 2410 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2488_
timestamp 0
transform -1 0 2410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2489_
timestamp 0
transform -1 0 1850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2490_
timestamp 0
transform -1 0 1410 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2491_
timestamp 0
transform -1 0 410 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2492_
timestamp 0
transform 1 0 4630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2493_
timestamp 0
transform 1 0 3630 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2494_
timestamp 0
transform 1 0 6210 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2495_
timestamp 0
transform 1 0 3870 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2496_
timestamp 0
transform 1 0 4170 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2497_
timestamp 0
transform -1 0 4090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2498_
timestamp 0
transform 1 0 3550 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2499_
timestamp 0
transform 1 0 3810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2500_
timestamp 0
transform -1 0 410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2501_
timestamp 0
transform -1 0 3410 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2502_
timestamp 0
transform -1 0 3050 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2503_
timestamp 0
transform -1 0 3530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__2504_
timestamp 0
transform -1 0 3290 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__2505_
timestamp 0
transform 1 0 2730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2506_
timestamp 0
transform -1 0 2550 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__2507_
timestamp 0
transform 1 0 670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2508_
timestamp 0
transform 1 0 3170 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2509_
timestamp 0
transform 1 0 2710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2510_
timestamp 0
transform -1 0 3270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2511_
timestamp 0
transform 1 0 3350 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__2512_
timestamp 0
transform 1 0 3190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2513_
timestamp 0
transform -1 0 2450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2514_
timestamp 0
transform 1 0 2150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2515_
timestamp 0
transform -1 0 2170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2516_
timestamp 0
transform -1 0 410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__2517_
timestamp 0
transform -1 0 2250 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2518_
timestamp 0
transform 1 0 5350 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2519_
timestamp 0
transform -1 0 5890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2520_
timestamp 0
transform -1 0 5990 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2521_
timestamp 0
transform 1 0 5690 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2522_
timestamp 0
transform -1 0 5690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2523_
timestamp 0
transform -1 0 5610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2524_
timestamp 0
transform -1 0 5550 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2525_
timestamp 0
transform -1 0 2770 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2526_
timestamp 0
transform 1 0 6170 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2527_
timestamp 0
transform 1 0 6570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2528_
timestamp 0
transform 1 0 6550 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2529_
timestamp 0
transform 1 0 6150 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2530_
timestamp 0
transform 1 0 5610 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2531_
timestamp 0
transform 1 0 2970 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2532_
timestamp 0
transform 1 0 4250 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2533_
timestamp 0
transform 1 0 5190 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2534_
timestamp 0
transform 1 0 4910 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2535_
timestamp 0
transform -1 0 4650 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2536_
timestamp 0
transform 1 0 3490 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2537_
timestamp 0
transform 1 0 2130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2538_
timestamp 0
transform 1 0 4530 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2539_
timestamp 0
transform 1 0 3910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2540_
timestamp 0
transform 1 0 4250 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2541_
timestamp 0
transform -1 0 4230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2542_
timestamp 0
transform -1 0 3750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2543_
timestamp 0
transform 1 0 3510 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2544_
timestamp 0
transform 1 0 4230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2545_
timestamp 0
transform 1 0 4490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2546_
timestamp 0
transform 1 0 4850 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2547_
timestamp 0
transform -1 0 4790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2548_
timestamp 0
transform -1 0 4510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2549_
timestamp 0
transform 1 0 4730 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2550_
timestamp 0
transform 1 0 4730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2551_
timestamp 0
transform 1 0 5250 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2552_
timestamp 0
transform 1 0 5490 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2553_
timestamp 0
transform 1 0 2390 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2554_
timestamp 0
transform 1 0 4530 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2555_
timestamp 0
transform -1 0 4710 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2556_
timestamp 0
transform -1 0 4950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2557_
timestamp 0
transform 1 0 4650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2558_
timestamp 0
transform 1 0 4730 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2559_
timestamp 0
transform 1 0 4450 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2560_
timestamp 0
transform 1 0 3950 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2561_
timestamp 0
transform 1 0 3650 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2562_
timestamp 0
transform 1 0 2270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2563_
timestamp 0
transform -1 0 4490 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2564_
timestamp 0
transform 1 0 4410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2565_
timestamp 0
transform -1 0 3890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2566_
timestamp 0
transform 1 0 2490 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2567_
timestamp 0
transform 1 0 3970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2568_
timestamp 0
transform -1 0 5770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2569_
timestamp 0
transform -1 0 5910 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2570_
timestamp 0
transform 1 0 5990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2571_
timestamp 0
transform 1 0 5990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2572_
timestamp 0
transform 1 0 5850 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2573_
timestamp 0
transform 1 0 5770 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2574_
timestamp 0
transform 1 0 5750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2575_
timestamp 0
transform -1 0 4790 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2576_
timestamp 0
transform -1 0 4270 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2577_
timestamp 0
transform -1 0 4530 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2578_
timestamp 0
transform 1 0 7030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2579_
timestamp 0
transform 1 0 7050 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2580_
timestamp 0
transform 1 0 8050 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2581_
timestamp 0
transform -1 0 8910 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2582_
timestamp 0
transform 1 0 6950 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2583_
timestamp 0
transform -1 0 6950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2584_
timestamp 0
transform 1 0 7370 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2585_
timestamp 0
transform 1 0 7410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2586_
timestamp 0
transform -1 0 8490 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2587_
timestamp 0
transform -1 0 6830 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2588_
timestamp 0
transform -1 0 5870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2589_
timestamp 0
transform 1 0 7490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2590_
timestamp 0
transform -1 0 6270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2591_
timestamp 0
transform 1 0 6510 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2592_
timestamp 0
transform -1 0 4490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2593_
timestamp 0
transform 1 0 5010 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2594_
timestamp 0
transform -1 0 8590 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2595_
timestamp 0
transform -1 0 5310 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2596_
timestamp 0
transform 1 0 5310 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2597_
timestamp 0
transform 1 0 5490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2598_
timestamp 0
transform -1 0 5230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2599_
timestamp 0
transform -1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2600_
timestamp 0
transform -1 0 5030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2601_
timestamp 0
transform -1 0 5290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2602_
timestamp 0
transform -1 0 8230 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2603_
timestamp 0
transform -1 0 6670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2604_
timestamp 0
transform -1 0 6430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2605_
timestamp 0
transform 1 0 6110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2606_
timestamp 0
transform -1 0 5610 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2607_
timestamp 0
transform 1 0 5770 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2608_
timestamp 0
transform 1 0 5590 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2609_
timestamp 0
transform -1 0 5570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2610_
timestamp 0
transform 1 0 4950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2611_
timestamp 0
transform -1 0 5210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2612_
timestamp 0
transform -1 0 5470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2613_
timestamp 0
transform -1 0 1290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2614_
timestamp 0
transform 1 0 2270 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2615_
timestamp 0
transform -1 0 2550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2616_
timestamp 0
transform -1 0 2530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2617_
timestamp 0
transform 1 0 1510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2618_
timestamp 0
transform 1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2619_
timestamp 0
transform -1 0 430 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2620_
timestamp 0
transform -1 0 670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2621_
timestamp 0
transform 1 0 990 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2622_
timestamp 0
transform 1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2623_
timestamp 0
transform 1 0 2810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2624_
timestamp 0
transform 1 0 2010 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2625_
timestamp 0
transform -1 0 2270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2626_
timestamp 0
transform -1 0 1990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2627_
timestamp 0
transform 1 0 130 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2628_
timestamp 0
transform 1 0 130 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2629_
timestamp 0
transform -1 0 390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2630_
timestamp 0
transform 1 0 130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2631_
timestamp 0
transform 1 0 5070 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2632_
timestamp 0
transform 1 0 2310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2633_
timestamp 0
transform -1 0 2610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2634_
timestamp 0
transform -1 0 150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2635_
timestamp 0
transform 1 0 130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2636_
timestamp 0
transform 1 0 670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2637_
timestamp 0
transform 1 0 1010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2638_
timestamp 0
transform 1 0 430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2639_
timestamp 0
transform -1 0 750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2640_
timestamp 0
transform -1 0 150 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2641_
timestamp 0
transform -1 0 150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2642_
timestamp 0
transform 1 0 1390 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2643_
timestamp 0
transform -1 0 1930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2644_
timestamp 0
transform 1 0 2330 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2645_
timestamp 0
transform -1 0 2070 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2646_
timestamp 0
transform -1 0 1270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2647_
timestamp 0
transform 1 0 130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2648_
timestamp 0
transform 1 0 630 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__2649_
timestamp 0
transform 1 0 130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2650_
timestamp 0
transform -1 0 3730 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2651_
timestamp 0
transform -1 0 3450 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2652_
timestamp 0
transform 1 0 670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2653_
timestamp 0
transform 1 0 390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2654_
timestamp 0
transform 1 0 1270 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2655_
timestamp 0
transform 1 0 710 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2656_
timestamp 0
transform -1 0 990 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2657_
timestamp 0
transform 1 0 130 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2658_
timestamp 0
transform 1 0 130 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2659_
timestamp 0
transform -1 0 430 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2660_
timestamp 0
transform 1 0 370 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2661_
timestamp 0
transform -1 0 2690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__2662_
timestamp 0
transform -1 0 2630 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2663_
timestamp 0
transform -1 0 2050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2664_
timestamp 0
transform 1 0 950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2665_
timestamp 0
transform -1 0 910 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2666_
timestamp 0
transform -1 0 430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2667_
timestamp 0
transform -1 0 650 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2668_
timestamp 0
transform 1 0 1150 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2669_
timestamp 0
transform -1 0 2910 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2670_
timestamp 0
transform -1 0 3030 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2671_
timestamp 0
transform 1 0 1190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2672_
timestamp 0
transform -1 0 690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2673_
timestamp 0
transform -1 0 650 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2674_
timestamp 0
transform 1 0 910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2675_
timestamp 0
transform 1 0 890 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2676_
timestamp 0
transform -1 0 1190 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2677_
timestamp 0
transform 1 0 6530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__2678_
timestamp 0
transform -1 0 6450 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2679_
timestamp 0
transform 1 0 7070 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2680_
timestamp 0
transform -1 0 6870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2681_
timestamp 0
transform 1 0 7130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2682_
timestamp 0
transform -1 0 6850 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2683_
timestamp 0
transform -1 0 1970 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2684_
timestamp 0
transform -1 0 1790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__2685_
timestamp 0
transform 1 0 1710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2686_
timestamp 0
transform 1 0 1710 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2687_
timestamp 0
transform 1 0 1450 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2688_
timestamp 0
transform -1 0 890 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2689_
timestamp 0
transform -1 0 870 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2690_
timestamp 0
transform 1 0 7370 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2691_
timestamp 0
transform -1 0 7210 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2692_
timestamp 0
transform -1 0 5150 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2693_
timestamp 0
transform -1 0 3110 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2694_
timestamp 0
transform -1 0 1410 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2695_
timestamp 0
transform -1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2696_
timestamp 0
transform -1 0 1410 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2697_
timestamp 0
transform 1 0 1990 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2698_
timestamp 0
transform -1 0 630 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2699_
timestamp 0
transform 1 0 6390 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2700_
timestamp 0
transform -1 0 7110 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2701_
timestamp 0
transform 1 0 7690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2702_
timestamp 0
transform 1 0 7390 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2703_
timestamp 0
transform 1 0 7550 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2704_
timestamp 0
transform -1 0 6750 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2705_
timestamp 0
transform 1 0 1670 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2706_
timestamp 0
transform 1 0 1110 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2707_
timestamp 0
transform 1 0 2810 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2708_
timestamp 0
transform 1 0 2490 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2709_
timestamp 0
transform -1 0 1170 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2710_
timestamp 0
transform -1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2711_
timestamp 0
transform -1 0 1230 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2712_
timestamp 0
transform 1 0 2970 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2713_
timestamp 0
transform -1 0 4370 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2714_
timestamp 0
transform -1 0 4790 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2715_
timestamp 0
transform 1 0 3630 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2716_
timestamp 0
transform -1 0 4390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2717_
timestamp 0
transform -1 0 5950 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__2718_
timestamp 0
transform -1 0 4190 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2719_
timestamp 0
transform 1 0 3790 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2720_
timestamp 0
transform -1 0 4090 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2721_
timestamp 0
transform -1 0 2250 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2722_
timestamp 0
transform 1 0 2370 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2723_
timestamp 0
transform 1 0 2670 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2724_
timestamp 0
transform -1 0 910 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2725_
timestamp 0
transform -1 0 5510 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2726_
timestamp 0
transform -1 0 6690 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2727_
timestamp 0
transform 1 0 3950 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2728_
timestamp 0
transform 1 0 3670 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2729_
timestamp 0
transform -1 0 3630 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2730_
timestamp 0
transform 1 0 3230 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2731_
timestamp 0
transform 1 0 2090 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2732_
timestamp 0
transform -1 0 1970 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2733_
timestamp 0
transform 1 0 1510 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2734_
timestamp 0
transform -1 0 1810 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2735_
timestamp 0
transform -1 0 3970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2736_
timestamp 0
transform -1 0 4110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2737_
timestamp 0
transform -1 0 4190 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2738_
timestamp 0
transform -1 0 3890 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2739_
timestamp 0
transform -1 0 3330 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2740_
timestamp 0
transform -1 0 3410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2741_
timestamp 0
transform -1 0 1170 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2742_
timestamp 0
transform 1 0 1470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2743_
timestamp 0
transform 1 0 1410 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2744_
timestamp 0
transform 1 0 1950 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2745_
timestamp 0
transform 1 0 610 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2746_
timestamp 0
transform 1 0 3670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2747_
timestamp 0
transform 1 0 4790 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__2748_
timestamp 0
transform 1 0 4450 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2749_
timestamp 0
transform -1 0 3610 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2750_
timestamp 0
transform -1 0 3050 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2751_
timestamp 0
transform 1 0 2890 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2752_
timestamp 0
transform 1 0 1190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2753_
timestamp 0
transform 1 0 690 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2754_
timestamp 0
transform -1 0 630 0 1 790
box -6 -8 26 268
use FILL  FILL_6__2755_
timestamp 0
transform -1 0 3150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2756_
timestamp 0
transform -1 0 2590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2757_
timestamp 0
transform 1 0 2830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2758_
timestamp 0
transform 1 0 2310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2759_
timestamp 0
transform -1 0 4390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2760_
timestamp 0
transform 1 0 3830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2761_
timestamp 0
transform 1 0 4170 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2762_
timestamp 0
transform -1 0 3910 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2763_
timestamp 0
transform -1 0 2150 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2764_
timestamp 0
transform -1 0 1870 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2765_
timestamp 0
transform -1 0 1790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2766_
timestamp 0
transform -1 0 2050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__2767_
timestamp 0
transform -1 0 1570 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__2768_
timestamp 0
transform 1 0 2230 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2769_
timestamp 0
transform 1 0 1670 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__2770_
timestamp 0
transform 1 0 6030 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2771_
timestamp 0
transform 1 0 6570 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2772_
timestamp 0
transform 1 0 5010 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__2773_
timestamp 0
transform 1 0 4210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2774_
timestamp 0
transform 1 0 2370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2775_
timestamp 0
transform 1 0 2610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2776_
timestamp 0
transform 1 0 3430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2777_
timestamp 0
transform -1 0 2910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2778_
timestamp 0
transform -1 0 3170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__2779_
timestamp 0
transform -1 0 7210 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2780_
timestamp 0
transform -1 0 7450 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__2781_
timestamp 0
transform 1 0 7930 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__2782_
timestamp 0
transform 1 0 7810 0 1 270
box -6 -8 26 268
use FILL  FILL_6__2783_
timestamp 0
transform 1 0 9750 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2784_
timestamp 0
transform 1 0 10890 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2785_
timestamp 0
transform 1 0 10270 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2786_
timestamp 0
transform 1 0 9990 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2787_
timestamp 0
transform 1 0 8450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2788_
timestamp 0
transform 1 0 8710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2789_
timestamp 0
transform 1 0 8230 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2790_
timestamp 0
transform -1 0 7970 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2791_
timestamp 0
transform 1 0 6230 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2792_
timestamp 0
transform 1 0 9850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2793_
timestamp 0
transform 1 0 10050 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2794_
timestamp 0
transform -1 0 10310 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2795_
timestamp 0
transform 1 0 8490 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2796_
timestamp 0
transform 1 0 8470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2797_
timestamp 0
transform 1 0 10870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2798_
timestamp 0
transform -1 0 10010 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2799_
timestamp 0
transform -1 0 8390 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2800_
timestamp 0
transform -1 0 7790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2801_
timestamp 0
transform 1 0 9730 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2802_
timestamp 0
transform -1 0 10050 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2803_
timestamp 0
transform 1 0 8490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2804_
timestamp 0
transform -1 0 8390 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2805_
timestamp 0
transform -1 0 10130 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2806_
timestamp 0
transform 1 0 9810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2807_
timestamp 0
transform -1 0 8430 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2808_
timestamp 0
transform -1 0 6670 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2809_
timestamp 0
transform 1 0 8190 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2810_
timestamp 0
transform -1 0 7610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2811_
timestamp 0
transform 1 0 10090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2812_
timestamp 0
transform 1 0 9730 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2813_
timestamp 0
transform 1 0 8310 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2814_
timestamp 0
transform -1 0 8190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2815_
timestamp 0
transform -1 0 8270 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2816_
timestamp 0
transform 1 0 9530 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2817_
timestamp 0
transform -1 0 10390 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2818_
timestamp 0
transform 1 0 11210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2819_
timestamp 0
transform 1 0 10190 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2820_
timestamp 0
transform -1 0 9970 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2821_
timestamp 0
transform -1 0 9830 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2822_
timestamp 0
transform -1 0 7550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2823_
timestamp 0
transform -1 0 9550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2824_
timestamp 0
transform -1 0 9290 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2825_
timestamp 0
transform 1 0 8750 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2826_
timestamp 0
transform 1 0 8790 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2827_
timestamp 0
transform 1 0 9210 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2828_
timestamp 0
transform 1 0 10330 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2829_
timestamp 0
transform -1 0 9270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2830_
timestamp 0
transform 1 0 9890 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2831_
timestamp 0
transform 1 0 9070 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2832_
timestamp 0
transform -1 0 8990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2833_
timestamp 0
transform -1 0 8750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2834_
timestamp 0
transform -1 0 8330 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2835_
timestamp 0
transform -1 0 9350 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2836_
timestamp 0
transform -1 0 8050 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2837_
timestamp 0
transform 1 0 8130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2838_
timestamp 0
transform 1 0 9370 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2839_
timestamp 0
transform 1 0 9630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2840_
timestamp 0
transform -1 0 9370 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2841_
timestamp 0
transform 1 0 8270 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2842_
timestamp 0
transform 1 0 11590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2843_
timestamp 0
transform -1 0 11090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2844_
timestamp 0
transform 1 0 10810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2845_
timestamp 0
transform 1 0 10550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2846_
timestamp 0
transform -1 0 10190 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2847_
timestamp 0
transform 1 0 10390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2848_
timestamp 0
transform -1 0 9670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2849_
timestamp 0
transform 1 0 10970 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__2850_
timestamp 0
transform 1 0 11130 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2851_
timestamp 0
transform 1 0 11370 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2852_
timestamp 0
transform 1 0 12070 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2853_
timestamp 0
transform 1 0 12130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2854_
timestamp 0
transform 1 0 11810 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2855_
timestamp 0
transform 1 0 12090 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2856_
timestamp 0
transform -1 0 9130 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2857_
timestamp 0
transform 1 0 9630 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2858_
timestamp 0
transform -1 0 9930 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2859_
timestamp 0
transform 1 0 10870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2860_
timestamp 0
transform 1 0 7750 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2861_
timestamp 0
transform 1 0 8430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2862_
timestamp 0
transform -1 0 7810 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2863_
timestamp 0
transform 1 0 7510 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2864_
timestamp 0
transform 1 0 9750 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2865_
timestamp 0
transform 1 0 8910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2866_
timestamp 0
transform -1 0 7010 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2867_
timestamp 0
transform -1 0 8850 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2868_
timestamp 0
transform -1 0 8570 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2869_
timestamp 0
transform -1 0 9010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2870_
timestamp 0
transform 1 0 8650 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2871_
timestamp 0
transform 1 0 8610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2872_
timestamp 0
transform 1 0 5550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2873_
timestamp 0
transform -1 0 5570 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2874_
timestamp 0
transform 1 0 5490 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2875_
timestamp 0
transform -1 0 5850 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2876_
timestamp 0
transform 1 0 5530 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2877_
timestamp 0
transform 1 0 6110 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2878_
timestamp 0
transform -1 0 5850 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2879_
timestamp 0
transform -1 0 8990 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2880_
timestamp 0
transform -1 0 11990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2881_
timestamp 0
transform 1 0 11670 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2882_
timestamp 0
transform -1 0 9270 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2883_
timestamp 0
transform 1 0 9070 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2884_
timestamp 0
transform -1 0 9390 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2885_
timestamp 0
transform -1 0 10570 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2886_
timestamp 0
transform 1 0 10530 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2887_
timestamp 0
transform -1 0 8950 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2888_
timestamp 0
transform -1 0 9230 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2889_
timestamp 0
transform 1 0 9510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2890_
timestamp 0
transform -1 0 9870 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__2891_
timestamp 0
transform -1 0 9810 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2892_
timestamp 0
transform 1 0 9190 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2893_
timestamp 0
transform -1 0 9350 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2894_
timestamp 0
transform -1 0 11170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2895_
timestamp 0
transform 1 0 10850 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2896_
timestamp 0
transform -1 0 11130 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2897_
timestamp 0
transform -1 0 10850 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2898_
timestamp 0
transform 1 0 9470 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2899_
timestamp 0
transform -1 0 9770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2900_
timestamp 0
transform 1 0 10450 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2901_
timestamp 0
transform -1 0 10470 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2902_
timestamp 0
transform 1 0 10650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2903_
timestamp 0
transform -1 0 10770 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2904_
timestamp 0
transform -1 0 9930 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2905_
timestamp 0
transform -1 0 9430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2906_
timestamp 0
transform -1 0 8590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2907_
timestamp 0
transform -1 0 9150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2908_
timestamp 0
transform -1 0 10490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2909_
timestamp 0
transform 1 0 11850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2910_
timestamp 0
transform 1 0 10930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2911_
timestamp 0
transform 1 0 11790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2912_
timestamp 0
transform 1 0 12070 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__2913_
timestamp 0
transform 1 0 10670 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__2914_
timestamp 0
transform -1 0 7850 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2915_
timestamp 0
transform 1 0 10990 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2916_
timestamp 0
transform 1 0 11230 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__2917_
timestamp 0
transform 1 0 10730 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2918_
timestamp 0
transform -1 0 10890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2919_
timestamp 0
transform 1 0 8570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2920_
timestamp 0
transform 1 0 11270 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2921_
timestamp 0
transform 1 0 11790 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__2922_
timestamp 0
transform -1 0 11910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2923_
timestamp 0
transform 1 0 11370 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2924_
timestamp 0
transform 1 0 10290 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2925_
timestamp 0
transform 1 0 10050 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2926_
timestamp 0
transform 1 0 10190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2927_
timestamp 0
transform -1 0 10030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2928_
timestamp 0
transform -1 0 10290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__2929_
timestamp 0
transform -1 0 10410 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__2930_
timestamp 0
transform -1 0 11290 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2931_
timestamp 0
transform -1 0 11550 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__2932_
timestamp 0
transform 1 0 11510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__2933_
timestamp 0
transform 1 0 11470 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__2934_
timestamp 0
transform 1 0 11550 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__2935_
timestamp 0
transform 1 0 11630 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2936_
timestamp 0
transform 1 0 10570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__2937_
timestamp 0
transform -1 0 3570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__2938_
timestamp 0
transform -1 0 7790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2939_
timestamp 0
transform 1 0 6550 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2940_
timestamp 0
transform -1 0 6330 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2941_
timestamp 0
transform -1 0 6250 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2942_
timestamp 0
transform 1 0 5150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2943_
timestamp 0
transform -1 0 7050 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__2944_
timestamp 0
transform 1 0 5430 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2945_
timestamp 0
transform -1 0 6830 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2946_
timestamp 0
transform 1 0 6430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__2947_
timestamp 0
transform 1 0 7910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2948_
timestamp 0
transform 1 0 7650 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2949_
timestamp 0
transform 1 0 5750 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__2950_
timestamp 0
transform -1 0 6090 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2951_
timestamp 0
transform 1 0 6850 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2952_
timestamp 0
transform 1 0 6570 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2953_
timestamp 0
transform 1 0 5730 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2954_
timestamp 0
transform -1 0 6030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__2955_
timestamp 0
transform 1 0 7110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2956_
timestamp 0
transform 1 0 6590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__2957_
timestamp 0
transform -1 0 8210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__2958_
timestamp 0
transform 1 0 6590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__2959_
timestamp 0
transform 1 0 6330 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2960_
timestamp 0
transform -1 0 7210 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2961_
timestamp 0
transform 1 0 6590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2962_
timestamp 0
transform -1 0 6370 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__2963_
timestamp 0
transform -1 0 6670 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2964_
timestamp 0
transform 1 0 4730 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2965_
timestamp 0
transform 1 0 5790 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2966_
timestamp 0
transform -1 0 6690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__2967_
timestamp 0
transform -1 0 5110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2968_
timestamp 0
transform -1 0 5370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2969_
timestamp 0
transform 1 0 4450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2970_
timestamp 0
transform 1 0 4810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2971_
timestamp 0
transform 1 0 4690 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2972_
timestamp 0
transform -1 0 6130 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2973_
timestamp 0
transform -1 0 6390 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2974_
timestamp 0
transform -1 0 6390 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2975_
timestamp 0
transform 1 0 5850 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2976_
timestamp 0
transform -1 0 4770 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2977_
timestamp 0
transform -1 0 5030 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2978_
timestamp 0
transform 1 0 5290 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__2979_
timestamp 0
transform 1 0 5570 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__2980_
timestamp 0
transform -1 0 7450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2981_
timestamp 0
transform -1 0 6410 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2982_
timestamp 0
transform -1 0 6690 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__2983_
timestamp 0
transform 1 0 7210 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2984_
timestamp 0
transform 1 0 6610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__2985_
timestamp 0
transform -1 0 6950 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2986_
timestamp 0
transform 1 0 6650 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2987_
timestamp 0
transform 1 0 6090 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2988_
timestamp 0
transform -1 0 6370 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__2989_
timestamp 0
transform -1 0 7950 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2990_
timestamp 0
transform 1 0 7070 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__2991_
timestamp 0
transform -1 0 6930 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2992_
timestamp 0
transform -1 0 5230 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__2993_
timestamp 0
transform -1 0 6090 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2994_
timestamp 0
transform 1 0 5550 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2995_
timestamp 0
transform 1 0 6630 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2996_
timestamp 0
transform 1 0 6350 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__2997_
timestamp 0
transform 1 0 6070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2998_
timestamp 0
transform -1 0 5810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__2999_
timestamp 0
transform 1 0 6470 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3000_
timestamp 0
transform -1 0 5810 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__3001_
timestamp 0
transform 1 0 5030 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3002_
timestamp 0
transform -1 0 5530 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__3003_
timestamp 0
transform -1 0 5890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3004_
timestamp 0
transform -1 0 5310 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3005_
timestamp 0
transform -1 0 5570 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3006_
timestamp 0
transform -1 0 7470 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3007_
timestamp 0
transform 1 0 6890 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3008_
timestamp 0
transform 1 0 8690 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3009_
timestamp 0
transform 1 0 8150 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3010_
timestamp 0
transform 1 0 7170 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3011_
timestamp 0
transform -1 0 7270 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3012_
timestamp 0
transform -1 0 7150 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3013_
timestamp 0
transform -1 0 7890 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3014_
timestamp 0
transform 1 0 7090 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3015_
timestamp 0
transform -1 0 7370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3016_
timestamp 0
transform -1 0 6130 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3017_
timestamp 0
transform -1 0 6930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3018_
timestamp 0
transform -1 0 6610 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3019_
timestamp 0
transform -1 0 6870 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3020_
timestamp 0
transform 1 0 5510 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__3021_
timestamp 0
transform 1 0 5950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3022_
timestamp 0
transform 1 0 5750 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__3023_
timestamp 0
transform -1 0 6830 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3024_
timestamp 0
transform -1 0 6750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3025_
timestamp 0
transform 1 0 6030 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__3026_
timestamp 0
transform 1 0 5450 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__3027_
timestamp 0
transform -1 0 5550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3028_
timestamp 0
transform 1 0 6030 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3029_
timestamp 0
transform 1 0 6790 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3030_
timestamp 0
transform 1 0 4930 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__3031_
timestamp 0
transform 1 0 4470 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3032_
timestamp 0
transform -1 0 5250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3033_
timestamp 0
transform 1 0 5510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3034_
timestamp 0
transform -1 0 3450 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3035_
timestamp 0
transform -1 0 4010 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3036_
timestamp 0
transform -1 0 3510 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3037_
timestamp 0
transform -1 0 3390 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3038_
timestamp 0
transform 1 0 3610 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3039_
timestamp 0
transform -1 0 3110 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3040_
timestamp 0
transform 1 0 2990 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3041_
timestamp 0
transform 1 0 3230 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3042_
timestamp 0
transform -1 0 3790 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3043_
timestamp 0
transform -1 0 3890 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3044_
timestamp 0
transform -1 0 3650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3045_
timestamp 0
transform 1 0 4450 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3046_
timestamp 0
transform 1 0 4170 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3047_
timestamp 0
transform -1 0 3130 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3048_
timestamp 0
transform 1 0 3170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3049_
timestamp 0
transform -1 0 2870 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3050_
timestamp 0
transform 1 0 2910 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3051_
timestamp 0
transform 1 0 2650 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3052_
timestamp 0
transform 1 0 2550 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3053_
timestamp 0
transform 1 0 3310 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3054_
timestamp 0
transform -1 0 3590 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3055_
timestamp 0
transform 1 0 3410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3056_
timestamp 0
transform -1 0 3670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3057_
timestamp 0
transform 1 0 3870 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3058_
timestamp 0
transform 1 0 4050 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3059_
timestamp 0
transform 1 0 4330 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3060_
timestamp 0
transform 1 0 4170 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3061_
timestamp 0
transform 1 0 3650 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3062_
timestamp 0
transform -1 0 3890 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3063_
timestamp 0
transform -1 0 5130 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__3064_
timestamp 0
transform 1 0 4990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__3065_
timestamp 0
transform -1 0 4730 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3066_
timestamp 0
transform 1 0 4630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3067_
timestamp 0
transform -1 0 3730 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3068_
timestamp 0
transform -1 0 3470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3069_
timestamp 0
transform 1 0 3670 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3070_
timestamp 0
transform -1 0 4570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__3071_
timestamp 0
transform 1 0 4290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__3072_
timestamp 0
transform -1 0 4230 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3073_
timestamp 0
transform -1 0 4490 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3074_
timestamp 0
transform 1 0 5770 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3075_
timestamp 0
transform 1 0 5490 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3076_
timestamp 0
transform 1 0 3730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3077_
timestamp 0
transform 1 0 4050 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3078_
timestamp 0
transform 1 0 4110 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3079_
timestamp 0
transform -1 0 4190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3080_
timestamp 0
transform 1 0 6330 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3081_
timestamp 0
transform -1 0 6990 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3082_
timestamp 0
transform 1 0 6690 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3083_
timestamp 0
transform -1 0 3870 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3084_
timestamp 0
transform 1 0 3570 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3085_
timestamp 0
transform 1 0 3190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3086_
timestamp 0
transform -1 0 2910 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3087_
timestamp 0
transform 1 0 4390 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3088_
timestamp 0
transform -1 0 4990 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3089_
timestamp 0
transform 1 0 3470 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3090_
timestamp 0
transform -1 0 3750 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3091_
timestamp 0
transform -1 0 6290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3092_
timestamp 0
transform 1 0 5510 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3093_
timestamp 0
transform 1 0 5770 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3094_
timestamp 0
transform 1 0 5490 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3095_
timestamp 0
transform -1 0 4690 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3096_
timestamp 0
transform 1 0 4390 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3097_
timestamp 0
transform -1 0 4150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3098_
timestamp 0
transform 1 0 3850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3099_
timestamp 0
transform -1 0 3910 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3100_
timestamp 0
transform -1 0 3730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3101_
timestamp 0
transform 1 0 4950 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3102_
timestamp 0
transform -1 0 5250 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3103_
timestamp 0
transform -1 0 4630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3104_
timestamp 0
transform -1 0 4910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3105_
timestamp 0
transform 1 0 5690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3106_
timestamp 0
transform -1 0 5990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3107_
timestamp 0
transform -1 0 4090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3108_
timestamp 0
transform 1 0 3790 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3109_
timestamp 0
transform 1 0 6270 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3110_
timestamp 0
transform 1 0 3950 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3111_
timestamp 0
transform 1 0 5810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3112_
timestamp 0
transform -1 0 5230 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3113_
timestamp 0
transform -1 0 4690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3114_
timestamp 0
transform 1 0 4390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3115_
timestamp 0
transform 1 0 4910 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3116_
timestamp 0
transform 1 0 3850 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3117_
timestamp 0
transform 1 0 4470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3118_
timestamp 0
transform -1 0 4770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3119_
timestamp 0
transform 1 0 4950 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3120_
timestamp 0
transform 1 0 4650 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3121_
timestamp 0
transform 1 0 5250 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3122_
timestamp 0
transform 1 0 5530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3123_
timestamp 0
transform 1 0 5510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3124_
timestamp 0
transform -1 0 5810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3125_
timestamp 0
transform -1 0 4170 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3126_
timestamp 0
transform 1 0 3870 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3127_
timestamp 0
transform 1 0 6530 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3128_
timestamp 0
transform 1 0 6090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3129_
timestamp 0
transform 1 0 5490 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3130_
timestamp 0
transform -1 0 3410 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3131_
timestamp 0
transform -1 0 3650 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3132_
timestamp 0
transform 1 0 4750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3133_
timestamp 0
transform 1 0 3990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3134_
timestamp 0
transform 1 0 5170 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3135_
timestamp 0
transform 1 0 4870 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3136_
timestamp 0
transform 1 0 5770 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3137_
timestamp 0
transform 1 0 5490 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3138_
timestamp 0
transform 1 0 5770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3139_
timestamp 0
transform 1 0 5490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3140_
timestamp 0
transform -1 0 5690 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3141_
timestamp 0
transform -1 0 5950 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3142_
timestamp 0
transform -1 0 4290 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3143_
timestamp 0
transform -1 0 4550 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3144_
timestamp 0
transform 1 0 11630 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__3145_
timestamp 0
transform 1 0 11870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__3146_
timestamp 0
transform -1 0 11930 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__3147_
timestamp 0
transform 1 0 9550 0 1 790
box -6 -8 26 268
use FILL  FILL_6__3148_
timestamp 0
transform -1 0 11930 0 1 790
box -6 -8 26 268
use FILL  FILL_6__3149_
timestamp 0
transform -1 0 11550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3150_
timestamp 0
transform -1 0 11830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3151_
timestamp 0
transform -1 0 10770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3152_
timestamp 0
transform 1 0 9410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3153_
timestamp 0
transform -1 0 9710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3154_
timestamp 0
transform -1 0 10230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3155_
timestamp 0
transform -1 0 10350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3156_
timestamp 0
transform -1 0 8990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__3157_
timestamp 0
transform -1 0 9030 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__3158_
timestamp 0
transform -1 0 8750 0 1 2870
box -6 -8 26 268
use FILL  FILL_6__3159_
timestamp 0
transform -1 0 8730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__3160_
timestamp 0
transform 1 0 10570 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3161_
timestamp 0
transform 1 0 10290 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3162_
timestamp 0
transform -1 0 9830 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3163_
timestamp 0
transform 1 0 9550 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3164_
timestamp 0
transform -1 0 9030 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3165_
timestamp 0
transform -1 0 7250 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3166_
timestamp 0
transform 1 0 7650 0 1 1310
box -6 -8 26 268
use FILL  FILL_6__3167_
timestamp 0
transform 1 0 7510 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3168_
timestamp 0
transform 1 0 7670 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3169_
timestamp 0
transform -1 0 8750 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3170_
timestamp 0
transform -1 0 8470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3171_
timestamp 0
transform -1 0 9190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3172_
timestamp 0
transform -1 0 8190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3173_
timestamp 0
transform 1 0 8450 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3174_
timestamp 0
transform 1 0 7930 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3175_
timestamp 0
transform -1 0 7910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3176_
timestamp 0
transform -1 0 7630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3177_
timestamp 0
transform -1 0 11910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__3178_
timestamp 0
transform -1 0 11850 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3179_
timestamp 0
transform 1 0 12110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3180_
timestamp 0
transform 1 0 12170 0 1 790
box -6 -8 26 268
use FILL  FILL_6__3181_
timestamp 0
transform 1 0 12150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__3182_
timestamp 0
transform -1 0 11370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3183_
timestamp 0
transform 1 0 11630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3184_
timestamp 0
transform 1 0 11910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3185_
timestamp 0
transform 1 0 11930 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3186_
timestamp 0
transform 1 0 12110 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3187_
timestamp 0
transform 1 0 9970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6__3188_
timestamp 0
transform 1 0 10850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3189_
timestamp 0
transform -1 0 11110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_6__3190_
timestamp 0
transform 1 0 11150 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3191_
timestamp 0
transform 1 0 11090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3192_
timestamp 0
transform -1 0 10810 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3193_
timestamp 0
transform 1 0 10230 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3194_
timestamp 0
transform 1 0 10850 0 1 2350
box -6 -8 26 268
use FILL  FILL_6__3195_
timestamp 0
transform -1 0 10590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3196_
timestamp 0
transform 1 0 10490 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3197_
timestamp 0
transform -1 0 7350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3198_
timestamp 0
transform -1 0 4710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3199_
timestamp 0
transform 1 0 2870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6__3200_
timestamp 0
transform 1 0 4850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__3201_
timestamp 0
transform 1 0 4570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__3202_
timestamp 0
transform 1 0 1630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6__3203_
timestamp 0
transform 1 0 1590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3204_
timestamp 0
transform 1 0 1550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__3205_
timestamp 0
transform 1 0 1110 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__3206_
timestamp 0
transform 1 0 1530 0 1 3390
box -6 -8 26 268
use FILL  FILL_6__3207_
timestamp 0
transform -1 0 1670 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__3208_
timestamp 0
transform -1 0 1010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__3209_
timestamp 0
transform -1 0 710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__3210_
timestamp 0
transform -1 0 4370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__3211_
timestamp 0
transform 1 0 4310 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__3212_
timestamp 0
transform 1 0 1270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6__3213_
timestamp 0
transform 1 0 1170 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__3214_
timestamp 0
transform -1 0 2450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3215_
timestamp 0
transform 1 0 1870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3216_
timestamp 0
transform 1 0 5810 0 1 270
box -6 -8 26 268
use FILL  FILL_6__3217_
timestamp 0
transform -1 0 6110 0 1 270
box -6 -8 26 268
use FILL  FILL_6__3218_
timestamp 0
transform 1 0 6150 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3219_
timestamp 0
transform -1 0 6430 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3220_
timestamp 0
transform 1 0 3770 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3221_
timestamp 0
transform -1 0 4050 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3222_
timestamp 0
transform -1 0 3650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3223_
timestamp 0
transform 1 0 3370 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__3224_
timestamp 0
transform -1 0 3350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3225_
timestamp 0
transform 1 0 5490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__3226_
timestamp 0
transform 1 0 5210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__3227_
timestamp 0
transform -1 0 4330 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3228_
timestamp 0
transform -1 0 4530 0 1 270
box -6 -8 26 268
use FILL  FILL_6__3229_
timestamp 0
transform 1 0 2770 0 1 1830
box -6 -8 26 268
use FILL  FILL_6__3230_
timestamp 0
transform -1 0 2810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6__3231_
timestamp 0
transform 1 0 6050 0 1 790
box -6 -8 26 268
use FILL  FILL_6__3232_
timestamp 0
transform 1 0 6030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6__3364_
timestamp 0
transform 1 0 5310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3365_
timestamp 0
transform 1 0 4510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3366_
timestamp 0
transform 1 0 4990 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__3367_
timestamp 0
transform -1 0 4790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3368_
timestamp 0
transform -1 0 5050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3369_
timestamp 0
transform -1 0 5610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3370_
timestamp 0
transform 1 0 2750 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3371_
timestamp 0
transform 1 0 2250 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3372_
timestamp 0
transform -1 0 2370 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3373_
timestamp 0
transform -1 0 4030 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3374_
timestamp 0
transform -1 0 2350 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3375_
timestamp 0
transform 1 0 2350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3376_
timestamp 0
transform -1 0 3010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3377_
timestamp 0
transform 1 0 2470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3378_
timestamp 0
transform -1 0 2330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3379_
timestamp 0
transform -1 0 1490 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3380_
timestamp 0
transform 1 0 1270 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3381_
timestamp 0
transform -1 0 1530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3382_
timestamp 0
transform -1 0 1990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3383_
timestamp 0
transform -1 0 1550 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3384_
timestamp 0
transform 1 0 1810 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3385_
timestamp 0
transform 1 0 1510 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3386_
timestamp 0
transform -1 0 2090 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3387_
timestamp 0
transform 1 0 2350 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3388_
timestamp 0
transform -1 0 690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3389_
timestamp 0
transform 1 0 2550 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3390_
timestamp 0
transform 1 0 3370 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3391_
timestamp 0
transform 1 0 3090 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3392_
timestamp 0
transform -1 0 2930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3393_
timestamp 0
transform 1 0 2330 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3394_
timestamp 0
transform 1 0 730 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3395_
timestamp 0
transform -1 0 690 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3396_
timestamp 0
transform -1 0 430 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3397_
timestamp 0
transform -1 0 450 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3398_
timestamp 0
transform -1 0 150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3399_
timestamp 0
transform 1 0 130 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3400_
timestamp 0
transform -1 0 930 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3401_
timestamp 0
transform -1 0 1510 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3402_
timestamp 0
transform 1 0 1490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3403_
timestamp 0
transform 1 0 1210 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3404_
timestamp 0
transform -1 0 150 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3405_
timestamp 0
transform -1 0 410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3406_
timestamp 0
transform -1 0 150 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3407_
timestamp 0
transform -1 0 430 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3408_
timestamp 0
transform -1 0 150 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3409_
timestamp 0
transform -1 0 150 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3410_
timestamp 0
transform 1 0 1470 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3411_
timestamp 0
transform 1 0 1190 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3412_
timestamp 0
transform -1 0 670 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3413_
timestamp 0
transform 1 0 410 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3414_
timestamp 0
transform 1 0 670 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6__3415_
timestamp 0
transform -1 0 990 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3416_
timestamp 0
transform 1 0 670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3417_
timestamp 0
transform -1 0 710 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3418_
timestamp 0
transform -1 0 410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3419_
timestamp 0
transform -1 0 1230 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3420_
timestamp 0
transform 1 0 930 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3421_
timestamp 0
transform 1 0 1230 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3422_
timestamp 0
transform 1 0 950 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3423_
timestamp 0
transform 1 0 1250 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3424_
timestamp 0
transform -1 0 1270 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3425_
timestamp 0
transform -1 0 990 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3426_
timestamp 0
transform 1 0 970 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6__3427_
timestamp 0
transform -1 0 1490 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3428_
timestamp 0
transform 1 0 1170 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3429_
timestamp 0
transform -1 0 950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3430_
timestamp 0
transform 1 0 1470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3431_
timestamp 0
transform 1 0 1190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3432_
timestamp 0
transform -1 0 990 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3433_
timestamp 0
transform -1 0 150 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3434_
timestamp 0
transform -1 0 730 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3435_
timestamp 0
transform -1 0 1010 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3436_
timestamp 0
transform -1 0 950 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3437_
timestamp 0
transform 1 0 1770 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3438_
timestamp 0
transform 1 0 1230 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3439_
timestamp 0
transform -1 0 1510 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3440_
timestamp 0
transform 1 0 1230 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3441_
timestamp 0
transform -1 0 670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3442_
timestamp 0
transform 1 0 1250 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3443_
timestamp 0
transform 1 0 1170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3444_
timestamp 0
transform -1 0 2070 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3445_
timestamp 0
transform 1 0 1750 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3446_
timestamp 0
transform 1 0 2110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3447_
timestamp 0
transform 1 0 2010 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3448_
timestamp 0
transform -1 0 1810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3449_
timestamp 0
transform 1 0 1490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3450_
timestamp 0
transform -1 0 950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3451_
timestamp 0
transform 1 0 1210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3452_
timestamp 0
transform 1 0 910 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3453_
timestamp 0
transform -1 0 2230 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3454_
timestamp 0
transform 1 0 3150 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3455_
timestamp 0
transform -1 0 2090 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3456_
timestamp 0
transform -1 0 1750 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3457_
timestamp 0
transform -1 0 2930 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3458_
timestamp 0
transform -1 0 1790 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3459_
timestamp 0
transform -1 0 1730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3460_
timestamp 0
transform 1 0 1770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3461_
timestamp 0
transform -1 0 1990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3462_
timestamp 0
transform -1 0 1750 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3463_
timestamp 0
transform -1 0 1510 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3464_
timestamp 0
transform 1 0 1230 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3465_
timestamp 0
transform -1 0 1490 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3466_
timestamp 0
transform 1 0 2030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3467_
timestamp 0
transform 1 0 2030 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3468_
timestamp 0
transform 1 0 2790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3469_
timestamp 0
transform 1 0 2650 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3470_
timestamp 0
transform -1 0 2550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3471_
timestamp 0
transform 1 0 2370 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3472_
timestamp 0
transform -1 0 2270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3473_
timestamp 0
transform 1 0 1510 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3474_
timestamp 0
transform -1 0 1770 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3475_
timestamp 0
transform 1 0 1250 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3476_
timestamp 0
transform -1 0 990 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3477_
timestamp 0
transform 1 0 410 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3478_
timestamp 0
transform -1 0 390 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3479_
timestamp 0
transform -1 0 150 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3480_
timestamp 0
transform -1 0 150 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3481_
timestamp 0
transform -1 0 150 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3482_
timestamp 0
transform 1 0 670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3483_
timestamp 0
transform -1 0 390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3484_
timestamp 0
transform 1 0 2010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3485_
timestamp 0
transform -1 0 2070 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3486_
timestamp 0
transform -1 0 1450 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3487_
timestamp 0
transform -1 0 1770 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3488_
timestamp 0
transform -1 0 1570 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3489_
timestamp 0
transform 1 0 1510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3490_
timestamp 0
transform 1 0 1190 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3491_
timestamp 0
transform -1 0 1270 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3492_
timestamp 0
transform 1 0 1170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3493_
timestamp 0
transform -1 0 990 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3494_
timestamp 0
transform 1 0 910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3495_
timestamp 0
transform -1 0 670 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3496_
timestamp 0
transform 1 0 430 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3497_
timestamp 0
transform -1 0 390 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3498_
timestamp 0
transform 1 0 690 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3499_
timestamp 0
transform -1 0 750 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3500_
timestamp 0
transform 1 0 690 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3501_
timestamp 0
transform 1 0 930 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3502_
timestamp 0
transform -1 0 450 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3503_
timestamp 0
transform -1 0 430 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3504_
timestamp 0
transform -1 0 670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3505_
timestamp 0
transform -1 0 430 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3506_
timestamp 0
transform -1 0 150 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3507_
timestamp 0
transform -1 0 150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3508_
timestamp 0
transform 1 0 670 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3509_
timestamp 0
transform -1 0 930 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3510_
timestamp 0
transform -1 0 430 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3511_
timestamp 0
transform -1 0 150 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3512_
timestamp 0
transform 1 0 630 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3513_
timestamp 0
transform -1 0 450 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3514_
timestamp 0
transform -1 0 390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3515_
timestamp 0
transform -1 0 150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3516_
timestamp 0
transform -1 0 150 0 1 10150
box -6 -8 26 268
use FILL  FILL_6__3517_
timestamp 0
transform 1 0 690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3518_
timestamp 0
transform 1 0 910 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3519_
timestamp 0
transform 1 0 2610 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3520_
timestamp 0
transform 1 0 2890 0 1 9110
box -6 -8 26 268
use FILL  FILL_6__3521_
timestamp 0
transform 1 0 3370 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3522_
timestamp 0
transform 1 0 3070 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3523_
timestamp 0
transform 1 0 2630 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3524_
timestamp 0
transform -1 0 1010 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3525_
timestamp 0
transform -1 0 150 0 1 10670
box -6 -8 26 268
use FILL  FILL_6__3526_
timestamp 0
transform -1 0 150 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3527_
timestamp 0
transform -1 0 650 0 1 11190
box -6 -8 26 268
use FILL  FILL_6__3528_
timestamp 0
transform -1 0 670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_6__3529_
timestamp 0
transform -1 0 150 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6__3530_
timestamp 0
transform -1 0 150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3531_
timestamp 0
transform 1 0 130 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3532_
timestamp 0
transform 1 0 370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3533_
timestamp 0
transform -1 0 150 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3534_
timestamp 0
transform -1 0 670 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3535_
timestamp 0
transform -1 0 430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6__3536_
timestamp 0
transform -1 0 410 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3537_
timestamp 0
transform -1 0 1770 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3538_
timestamp 0
transform 1 0 2530 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3539_
timestamp 0
transform -1 0 2630 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3540_
timestamp 0
transform -1 0 2370 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3541_
timestamp 0
transform -1 0 2090 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3542_
timestamp 0
transform -1 0 2270 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3543_
timestamp 0
transform 1 0 1670 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3544_
timestamp 0
transform 1 0 2030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3545_
timestamp 0
transform 1 0 1830 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3546_
timestamp 0
transform 1 0 1950 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6__3547_
timestamp 0
transform -1 0 2610 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3548_
timestamp 0
transform 1 0 2310 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6__3549_
timestamp 0
transform -1 0 2410 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3550_
timestamp 0
transform 1 0 2110 0 1 11710
box -6 -8 26 268
use FILL  FILL_6__3551_
timestamp 0
transform -1 0 2590 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3552_
timestamp 0
transform 1 0 2290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6__3553_
timestamp 0
transform -1 0 1830 0 1 8070
box -6 -8 26 268
use FILL  FILL_6__3554_
timestamp 0
transform 1 0 970 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3555_
timestamp 0
transform 1 0 370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3556_
timestamp 0
transform 1 0 1230 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6__3557_
timestamp 0
transform -1 0 3130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3558_
timestamp 0
transform 1 0 2830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6__3559_
timestamp 0
transform -1 0 2590 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3560_
timestamp 0
transform 1 0 2290 0 1 9630
box -6 -8 26 268
use FILL  FILL_6__3561_
timestamp 0
transform -1 0 2010 0 1 7550
box -6 -8 26 268
use FILL  FILL_6__3562_
timestamp 0
transform -1 0 2830 0 1 8590
box -6 -8 26 268
use FILL  FILL_6__3563_
timestamp 0
transform 1 0 2230 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6__3564_
timestamp 0
transform 1 0 2510 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3565_
timestamp 0
transform -1 0 1510 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3566_
timestamp 0
transform -1 0 1770 0 1 7030
box -6 -8 26 268
use FILL  FILL_6__3579_
timestamp 0
transform -1 0 5110 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3580_
timestamp 0
transform -1 0 150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6__3581_
timestamp 0
transform -1 0 3530 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3582_
timestamp 0
transform -1 0 3270 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3583_
timestamp 0
transform -1 0 5390 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__3584_
timestamp 0
transform 1 0 4570 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3585_
timestamp 0
transform 1 0 2990 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3586_
timestamp 0
transform -1 0 5910 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__3587_
timestamp 0
transform 1 0 130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3588_
timestamp 0
transform -1 0 150 0 1 3910
box -6 -8 26 268
use FILL  FILL_6__3589_
timestamp 0
transform -1 0 150 0 1 4950
box -6 -8 26 268
use FILL  FILL_6__3590_
timestamp 0
transform -1 0 150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6__3591_
timestamp 0
transform -1 0 430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3592_
timestamp 0
transform -1 0 150 0 1 4430
box -6 -8 26 268
use FILL  FILL_6__3593_
timestamp 0
transform -1 0 4850 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3594_
timestamp 0
transform 1 0 5890 0 -1 270
box -6 -8 26 268
use FILL  FILL_6__3595_
timestamp 0
transform 1 0 5630 0 -1 790
box -6 -8 26 268
use FILL  FILL_6__3596_
timestamp 0
transform -1 0 930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3597_
timestamp 0
transform -1 0 150 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__3598_
timestamp 0
transform -1 0 410 0 1 5990
box -6 -8 26 268
use FILL  FILL_6__3599_
timestamp 0
transform -1 0 150 0 1 6510
box -6 -8 26 268
use FILL  FILL_6__3600_
timestamp 0
transform -1 0 150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6__3601_
timestamp 0
transform -1 0 150 0 1 5470
box -6 -8 26 268
use FILL  FILL_6__3602_
timestamp 0
transform -1 0 1770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6__3603_
timestamp 0
transform 1 0 6930 0 -1 270
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert0
timestamp 0
transform 1 0 7950 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert1
timestamp 0
transform 1 0 9450 0 1 1830
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert2
timestamp 0
transform 1 0 8210 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert3
timestamp 0
transform 1 0 11070 0 1 1830
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert4
timestamp 0
transform 1 0 670 0 1 1830
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert5
timestamp 0
transform -1 0 12150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert6
timestamp 0
transform -1 0 9650 0 1 5470
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert7
timestamp 0
transform 1 0 7110 0 1 2350
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert8
timestamp 0
transform -1 0 930 0 1 5470
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert9
timestamp 0
transform 1 0 10190 0 1 3910
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert10
timestamp 0
transform -1 0 970 0 1 5990
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert11
timestamp 0
transform -1 0 6050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert12
timestamp 0
transform 1 0 11610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert13
timestamp 0
transform -1 0 6230 0 1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert14
timestamp 0
transform 1 0 6850 0 1 2350
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert15
timestamp 0
transform -1 0 3390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert16
timestamp 0
transform -1 0 4010 0 1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert17
timestamp 0
transform 1 0 7250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert18
timestamp 0
transform -1 0 7070 0 1 11190
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert19
timestamp 0
transform 1 0 5390 0 1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert20
timestamp 0
transform 1 0 8630 0 1 11190
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert21
timestamp 0
transform -1 0 8550 0 -1 7550
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert22
timestamp 0
transform -1 0 1510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert23
timestamp 0
transform 1 0 3490 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert24
timestamp 0
transform -1 0 4390 0 1 5470
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert25
timestamp 0
transform 1 0 8230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert26
timestamp 0
transform 1 0 5170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert27
timestamp 0
transform -1 0 1310 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert39
timestamp 0
transform 1 0 6390 0 1 4950
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert40
timestamp 0
transform 1 0 7750 0 1 3910
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert41
timestamp 0
transform -1 0 8890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert42
timestamp 0
transform -1 0 7030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert43
timestamp 0
transform -1 0 8930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert44
timestamp 0
transform -1 0 9050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert45
timestamp 0
transform 1 0 11110 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert46
timestamp 0
transform 1 0 9550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert47
timestamp 0
transform 1 0 9270 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert48
timestamp 0
transform 1 0 7010 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert49
timestamp 0
transform 1 0 7270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert50
timestamp 0
transform -1 0 7650 0 1 9110
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert51
timestamp 0
transform 1 0 7610 0 1 10150
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert52
timestamp 0
transform 1 0 9010 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert53
timestamp 0
transform 1 0 10050 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert54
timestamp 0
transform 1 0 8890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert55
timestamp 0
transform 1 0 8750 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert56
timestamp 0
transform -1 0 2290 0 1 8590
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert57
timestamp 0
transform 1 0 2590 0 1 11190
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert58
timestamp 0
transform 1 0 2730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert59
timestamp 0
transform -1 0 2290 0 1 10670
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert60
timestamp 0
transform -1 0 10550 0 1 7550
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert61
timestamp 0
transform 1 0 10610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert62
timestamp 0
transform 1 0 10570 0 1 8070
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert63
timestamp 0
transform -1 0 9230 0 1 7550
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert64
timestamp 0
transform -1 0 8670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert65
timestamp 0
transform 1 0 5270 0 1 270
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert66
timestamp 0
transform 1 0 5790 0 1 790
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert67
timestamp 0
transform -1 0 3090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert68
timestamp 0
transform 1 0 3210 0 1 270
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert69
timestamp 0
transform -1 0 6710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert70
timestamp 0
transform 1 0 8650 0 1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert71
timestamp 0
transform -1 0 9310 0 1 2870
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert72
timestamp 0
transform -1 0 6830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert73
timestamp 0
transform 1 0 8990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert74
timestamp 0
transform 1 0 10850 0 1 7030
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert75
timestamp 0
transform 1 0 2630 0 1 1310
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert76
timestamp 0
transform -1 0 3130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert77
timestamp 0
transform 1 0 10510 0 1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert78
timestamp 0
transform 1 0 9370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert79
timestamp 0
transform -1 0 8410 0 1 7550
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert80
timestamp 0
transform 1 0 7210 0 1 5470
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert81
timestamp 0
transform 1 0 7670 0 -1 790
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert82
timestamp 0
transform -1 0 7650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert83
timestamp 0
transform -1 0 7430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert84
timestamp 0
transform 1 0 9490 0 1 8590
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert85
timestamp 0
transform -1 0 8970 0 1 8590
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert86
timestamp 0
transform -1 0 9570 0 1 2870
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert87
timestamp 0
transform 1 0 9470 0 1 4430
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert88
timestamp 0
transform -1 0 10810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert89
timestamp 0
transform 1 0 9450 0 1 3390
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert90
timestamp 0
transform 1 0 5430 0 -1 11190
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert91
timestamp 0
transform -1 0 4970 0 1 10670
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert92
timestamp 0
transform -1 0 4810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert93
timestamp 0
transform 1 0 5230 0 1 10150
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert94
timestamp 0
transform -1 0 11390 0 1 9630
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert95
timestamp 0
transform -1 0 11430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert96
timestamp 0
transform -1 0 10150 0 1 11710
box -6 -8 26 268
use FILL  FILL_6_BUFX2_insert97
timestamp 0
transform 1 0 11510 0 1 11710
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert28
timestamp 0
transform -1 0 6090 0 -1 11710
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert29
timestamp 0
transform -1 0 2270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert30
timestamp 0
transform 1 0 4610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert31
timestamp 0
transform -1 0 3310 0 1 2870
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert32
timestamp 0
transform 1 0 7210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert33
timestamp 0
transform 1 0 5790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert34
timestamp 0
transform -1 0 2550 0 1 10670
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert35
timestamp 0
transform -1 0 5310 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert36
timestamp 0
transform -1 0 2430 0 1 3910
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert37
timestamp 0
transform 1 0 7450 0 -1 12230
box -6 -8 26 268
use FILL  FILL_6_CLKBUF1_insert38
timestamp 0
transform -1 0 4430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__1688_
timestamp 0
transform -1 0 970 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1689_
timestamp 0
transform -1 0 430 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1690_
timestamp 0
transform -1 0 690 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1691_
timestamp 0
transform 1 0 150 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1692_
timestamp 0
transform -1 0 410 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1693_
timestamp 0
transform 1 0 650 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1694_
timestamp 0
transform -1 0 5650 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__1695_
timestamp 0
transform -1 0 430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1696_
timestamp 0
transform -1 0 430 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1697_
timestamp 0
transform -1 0 1550 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__1698_
timestamp 0
transform -1 0 3490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1699_
timestamp 0
transform 1 0 2930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1700_
timestamp 0
transform -1 0 3970 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__1701_
timestamp 0
transform -1 0 670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1702_
timestamp 0
transform -1 0 670 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1703_
timestamp 0
transform 1 0 3310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1704_
timestamp 0
transform -1 0 450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1705_
timestamp 0
transform 1 0 150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1706_
timestamp 0
transform -1 0 3930 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1707_
timestamp 0
transform -1 0 690 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1708_
timestamp 0
transform 1 0 690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1709_
timestamp 0
transform 1 0 4210 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1710_
timestamp 0
transform -1 0 5690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1711_
timestamp 0
transform 1 0 5230 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1712_
timestamp 0
transform 1 0 7370 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1713_
timestamp 0
transform -1 0 9750 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1714_
timestamp 0
transform -1 0 9950 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1715_
timestamp 0
transform -1 0 8630 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1716_
timestamp 0
transform 1 0 11390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1717_
timestamp 0
transform 1 0 11190 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1718_
timestamp 0
transform 1 0 12010 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1719_
timestamp 0
transform -1 0 8890 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1720_
timestamp 0
transform -1 0 10210 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1721_
timestamp 0
transform -1 0 10230 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1722_
timestamp 0
transform -1 0 9990 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1723_
timestamp 0
transform 1 0 10090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1724_
timestamp 0
transform 1 0 9310 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1725_
timestamp 0
transform 1 0 9150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1726_
timestamp 0
transform 1 0 10250 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1727_
timestamp 0
transform -1 0 8870 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1728_
timestamp 0
transform 1 0 11650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1729_
timestamp 0
transform 1 0 10250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1730_
timestamp 0
transform 1 0 8430 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1731_
timestamp 0
transform 1 0 8670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1732_
timestamp 0
transform -1 0 7870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1733_
timestamp 0
transform 1 0 9810 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1734_
timestamp 0
transform 1 0 7510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1735_
timestamp 0
transform 1 0 10950 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1736_
timestamp 0
transform -1 0 10750 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1737_
timestamp 0
transform -1 0 11010 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1738_
timestamp 0
transform -1 0 10390 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1739_
timestamp 0
transform -1 0 10390 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1740_
timestamp 0
transform 1 0 10610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1741_
timestamp 0
transform -1 0 8510 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1742_
timestamp 0
transform -1 0 8410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1743_
timestamp 0
transform -1 0 9970 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1744_
timestamp 0
transform 1 0 9850 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1745_
timestamp 0
transform -1 0 9550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1746_
timestamp 0
transform 1 0 11410 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1747_
timestamp 0
transform 1 0 10890 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1748_
timestamp 0
transform 1 0 7610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1749_
timestamp 0
transform 1 0 8030 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__1750_
timestamp 0
transform -1 0 8150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1751_
timestamp 0
transform 1 0 7550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1752_
timestamp 0
transform -1 0 8970 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1753_
timestamp 0
transform 1 0 9830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1754_
timestamp 0
transform -1 0 8370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1755_
timestamp 0
transform -1 0 8950 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__1756_
timestamp 0
transform -1 0 11290 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1757_
timestamp 0
transform 1 0 11150 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1758_
timestamp 0
transform -1 0 9210 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1759_
timestamp 0
transform -1 0 7450 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__1760_
timestamp 0
transform 1 0 8950 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__1761_
timestamp 0
transform -1 0 9670 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1762_
timestamp 0
transform 1 0 10690 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1763_
timestamp 0
transform -1 0 9130 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1764_
timestamp 0
transform 1 0 11390 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1765_
timestamp 0
transform 1 0 8210 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1766_
timestamp 0
transform 1 0 8590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1767_
timestamp 0
transform 1 0 9290 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__1768_
timestamp 0
transform 1 0 8150 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__1769_
timestamp 0
transform 1 0 8670 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__1770_
timestamp 0
transform 1 0 9110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__1771_
timestamp 0
transform 1 0 9070 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__1772_
timestamp 0
transform 1 0 8790 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__1773_
timestamp 0
transform 1 0 10870 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1774_
timestamp 0
transform 1 0 10870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1775_
timestamp 0
transform 1 0 10110 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1776_
timestamp 0
transform -1 0 8110 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1777_
timestamp 0
transform 1 0 8150 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1778_
timestamp 0
transform -1 0 7630 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1779_
timestamp 0
transform 1 0 5770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1780_
timestamp 0
transform -1 0 4170 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1781_
timestamp 0
transform -1 0 10890 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1782_
timestamp 0
transform 1 0 8370 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1783_
timestamp 0
transform 1 0 10610 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1784_
timestamp 0
transform -1 0 10090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1785_
timestamp 0
transform -1 0 9850 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1786_
timestamp 0
transform 1 0 10270 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1787_
timestamp 0
transform -1 0 9210 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1788_
timestamp 0
transform -1 0 8630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1789_
timestamp 0
transform 1 0 10070 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1790_
timestamp 0
transform -1 0 10130 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1791_
timestamp 0
transform -1 0 10210 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1792_
timestamp 0
transform -1 0 9750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1793_
timestamp 0
transform -1 0 9490 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1794_
timestamp 0
transform 1 0 9210 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1795_
timestamp 0
transform -1 0 8410 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1796_
timestamp 0
transform -1 0 8350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1797_
timestamp 0
transform 1 0 7190 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1798_
timestamp 0
transform 1 0 7450 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1799_
timestamp 0
transform -1 0 9470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1800_
timestamp 0
transform 1 0 11350 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1801_
timestamp 0
transform 1 0 9370 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1802_
timestamp 0
transform -1 0 9030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1803_
timestamp 0
transform 1 0 10630 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1804_
timestamp 0
transform -1 0 8650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1805_
timestamp 0
transform -1 0 8750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1806_
timestamp 0
transform 1 0 7690 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1807_
timestamp 0
transform -1 0 8150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1808_
timestamp 0
transform -1 0 8470 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1809_
timestamp 0
transform 1 0 8690 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1810_
timestamp 0
transform 1 0 8090 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1811_
timestamp 0
transform -1 0 7830 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1812_
timestamp 0
transform -1 0 8470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1813_
timestamp 0
transform -1 0 8190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1814_
timestamp 0
transform -1 0 7930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1815_
timestamp 0
transform 1 0 7950 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1816_
timestamp 0
transform -1 0 3950 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1817_
timestamp 0
transform 1 0 1430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1818_
timestamp 0
transform -1 0 6250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1819_
timestamp 0
transform -1 0 1010 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1820_
timestamp 0
transform 1 0 450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1821_
timestamp 0
transform 1 0 970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1822_
timestamp 0
transform -1 0 430 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1823_
timestamp 0
transform 1 0 1790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1824_
timestamp 0
transform 1 0 1370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__1825_
timestamp 0
transform -1 0 1210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1826_
timestamp 0
transform -1 0 470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1827_
timestamp 0
transform 1 0 970 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1828_
timestamp 0
transform -1 0 1570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1829_
timestamp 0
transform -1 0 710 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1830_
timestamp 0
transform -1 0 1510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1831_
timestamp 0
transform 1 0 2090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1832_
timestamp 0
transform -1 0 8090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1833_
timestamp 0
transform 1 0 9730 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1834_
timestamp 0
transform 1 0 9310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1835_
timestamp 0
transform -1 0 7830 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1836_
timestamp 0
transform -1 0 6490 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1837_
timestamp 0
transform -1 0 7830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1838_
timestamp 0
transform -1 0 7270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1839_
timestamp 0
transform -1 0 6250 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1840_
timestamp 0
transform 1 0 8630 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1841_
timestamp 0
transform -1 0 8250 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1842_
timestamp 0
transform -1 0 7010 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1843_
timestamp 0
transform -1 0 6730 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1844_
timestamp 0
transform 1 0 9150 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1845_
timestamp 0
transform 1 0 9690 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1846_
timestamp 0
transform -1 0 9290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1847_
timestamp 0
transform -1 0 8450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1848_
timestamp 0
transform 1 0 11290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1849_
timestamp 0
transform -1 0 11610 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1850_
timestamp 0
transform -1 0 11070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1851_
timestamp 0
transform 1 0 10430 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1852_
timestamp 0
transform -1 0 10490 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1853_
timestamp 0
transform -1 0 10510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__1854_
timestamp 0
transform -1 0 7490 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1855_
timestamp 0
transform 1 0 7470 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1856_
timestamp 0
transform 1 0 7750 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1857_
timestamp 0
transform -1 0 8890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__1858_
timestamp 0
transform -1 0 9430 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1859_
timestamp 0
transform -1 0 8890 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1860_
timestamp 0
transform 1 0 9150 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1861_
timestamp 0
transform 1 0 6890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1862_
timestamp 0
transform -1 0 8390 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__1863_
timestamp 0
transform 1 0 7750 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1864_
timestamp 0
transform -1 0 6390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1865_
timestamp 0
transform -1 0 7830 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__1866_
timestamp 0
transform -1 0 7290 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1867_
timestamp 0
transform -1 0 8070 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1868_
timestamp 0
transform 1 0 7790 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1869_
timestamp 0
transform -1 0 6090 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__1870_
timestamp 0
transform 1 0 9430 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1871_
timestamp 0
transform 1 0 8910 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1872_
timestamp 0
transform -1 0 8650 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1873_
timestamp 0
transform -1 0 7850 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1874_
timestamp 0
transform -1 0 7570 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1875_
timestamp 0
transform -1 0 8370 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1876_
timestamp 0
transform -1 0 7010 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1877_
timestamp 0
transform -1 0 5850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__1878_
timestamp 0
transform 1 0 6730 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1879_
timestamp 0
transform -1 0 7530 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1880_
timestamp 0
transform 1 0 6050 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__1881_
timestamp 0
transform 1 0 6050 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__1882_
timestamp 0
transform -1 0 5010 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__1883_
timestamp 0
transform -1 0 7910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1884_
timestamp 0
transform -1 0 8150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1885_
timestamp 0
transform -1 0 8710 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__1886_
timestamp 0
transform 1 0 8550 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1887_
timestamp 0
transform -1 0 8530 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1888_
timestamp 0
transform 1 0 11670 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1889_
timestamp 0
transform -1 0 8530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1890_
timestamp 0
transform 1 0 9790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1891_
timestamp 0
transform 1 0 8950 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1892_
timestamp 0
transform -1 0 8670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1893_
timestamp 0
transform 1 0 12190 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1894_
timestamp 0
transform 1 0 12170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1895_
timestamp 0
transform 1 0 12190 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1896_
timestamp 0
transform -1 0 10810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1897_
timestamp 0
transform -1 0 9210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1898_
timestamp 0
transform 1 0 9090 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1899_
timestamp 0
transform 1 0 7530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1900_
timestamp 0
transform 1 0 9730 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1901_
timestamp 0
transform 1 0 8070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1902_
timestamp 0
transform -1 0 8290 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1903_
timestamp 0
transform 1 0 8010 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1904_
timestamp 0
transform 1 0 11930 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1905_
timestamp 0
transform 1 0 11690 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1906_
timestamp 0
transform -1 0 6570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1907_
timestamp 0
transform -1 0 7110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1908_
timestamp 0
transform -1 0 7030 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1909_
timestamp 0
transform -1 0 6790 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__1910_
timestamp 0
transform -1 0 6290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1911_
timestamp 0
transform 1 0 6870 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1912_
timestamp 0
transform 1 0 6330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__1913_
timestamp 0
transform 1 0 6270 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1914_
timestamp 0
transform 1 0 5770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1915_
timestamp 0
transform 1 0 5290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1916_
timestamp 0
transform 1 0 5290 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__1917_
timestamp 0
transform -1 0 3790 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__1918_
timestamp 0
transform 1 0 3670 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__1919_
timestamp 0
transform -1 0 3950 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__1920_
timestamp 0
transform -1 0 3670 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__1921_
timestamp 0
transform -1 0 1790 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__1922_
timestamp 0
transform 1 0 7590 0 1 270
box -6 -8 26 268
use FILL  FILL_7__1923_
timestamp 0
transform 1 0 7850 0 1 790
box -6 -8 26 268
use FILL  FILL_7__1924_
timestamp 0
transform -1 0 6450 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__1925_
timestamp 0
transform -1 0 4690 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1926_
timestamp 0
transform -1 0 4050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1927_
timestamp 0
transform 1 0 2090 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__1928_
timestamp 0
transform -1 0 3250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__1929_
timestamp 0
transform 1 0 4630 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__1930_
timestamp 0
transform 1 0 3190 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__1931_
timestamp 0
transform -1 0 2970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__1932_
timestamp 0
transform -1 0 1570 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1933_
timestamp 0
transform -1 0 8530 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1934_
timestamp 0
transform 1 0 3930 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__1935_
timestamp 0
transform -1 0 3950 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1936_
timestamp 0
transform -1 0 2630 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1937_
timestamp 0
transform -1 0 1290 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1938_
timestamp 0
transform -1 0 3650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1939_
timestamp 0
transform -1 0 4210 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1940_
timestamp 0
transform -1 0 3430 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1941_
timestamp 0
transform -1 0 3370 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1942_
timestamp 0
transform -1 0 1870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__1943_
timestamp 0
transform -1 0 3670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__1944_
timestamp 0
transform -1 0 3770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1945_
timestamp 0
transform -1 0 3030 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__1946_
timestamp 0
transform -1 0 1590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__1947_
timestamp 0
transform -1 0 5010 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__1948_
timestamp 0
transform 1 0 5210 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__1949_
timestamp 0
transform 1 0 5270 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__1950_
timestamp 0
transform -1 0 5010 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__1951_
timestamp 0
transform -1 0 2050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1952_
timestamp 0
transform 1 0 4170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__1953_
timestamp 0
transform 1 0 4110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__1954_
timestamp 0
transform 1 0 4250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1955_
timestamp 0
transform -1 0 1770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1956_
timestamp 0
transform -1 0 4390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__1957_
timestamp 0
transform 1 0 4970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__1958_
timestamp 0
transform -1 0 5250 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__1959_
timestamp 0
transform -1 0 4230 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__1960_
timestamp 0
transform -1 0 2390 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1961_
timestamp 0
transform 1 0 4210 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1962_
timestamp 0
transform 1 0 3970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1963_
timestamp 0
transform 1 0 3750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1964_
timestamp 0
transform 1 0 2090 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1965_
timestamp 0
transform 1 0 6470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__1966_
timestamp 0
transform 1 0 6410 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1967_
timestamp 0
transform 1 0 7250 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1968_
timestamp 0
transform 1 0 6710 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1969_
timestamp 0
transform -1 0 3370 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__1970_
timestamp 0
transform 1 0 2910 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1971_
timestamp 0
transform -1 0 4790 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1972_
timestamp 0
transform 1 0 3650 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1973_
timestamp 0
transform -1 0 3670 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__1974_
timestamp 0
transform -1 0 3170 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__1975_
timestamp 0
transform 1 0 3070 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__1976_
timestamp 0
transform -1 0 3170 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__1977_
timestamp 0
transform 1 0 4450 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__1978_
timestamp 0
transform 1 0 3150 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__1979_
timestamp 0
transform -1 0 2890 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__1980_
timestamp 0
transform -1 0 2410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1981_
timestamp 0
transform 1 0 6030 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__1982_
timestamp 0
transform 1 0 6150 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__1983_
timestamp 0
transform 1 0 6350 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__1984_
timestamp 0
transform 1 0 5350 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__1985_
timestamp 0
transform -1 0 4850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1986_
timestamp 0
transform 1 0 2630 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__1987_
timestamp 0
transform -1 0 7350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__1988_
timestamp 0
transform 1 0 7650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__1989_
timestamp 0
transform 1 0 7710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__1990_
timestamp 0
transform -1 0 7510 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1991_
timestamp 0
transform -1 0 7790 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__1992_
timestamp 0
transform 1 0 10530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__1993_
timestamp 0
transform 1 0 9650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__1994_
timestamp 0
transform -1 0 6330 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__1995_
timestamp 0
transform 1 0 6710 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__1996_
timestamp 0
transform -1 0 6850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1997_
timestamp 0
transform 1 0 6550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__1998_
timestamp 0
transform 1 0 6550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__1999_
timestamp 0
transform 1 0 7610 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2000_
timestamp 0
transform 1 0 6530 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2001_
timestamp 0
transform 1 0 6770 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2002_
timestamp 0
transform 1 0 6730 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2003_
timestamp 0
transform 1 0 9610 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2004_
timestamp 0
transform 1 0 7550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2005_
timestamp 0
transform -1 0 7350 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2006_
timestamp 0
transform 1 0 6830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2007_
timestamp 0
transform 1 0 6670 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2008_
timestamp 0
transform -1 0 6310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2009_
timestamp 0
transform 1 0 6910 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2010_
timestamp 0
transform -1 0 7130 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2011_
timestamp 0
transform 1 0 7370 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2012_
timestamp 0
transform -1 0 9510 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2013_
timestamp 0
transform 1 0 10650 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2014_
timestamp 0
transform -1 0 10910 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2015_
timestamp 0
transform -1 0 6350 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2016_
timestamp 0
transform -1 0 7390 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2017_
timestamp 0
transform -1 0 7170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2018_
timestamp 0
transform 1 0 7410 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2019_
timestamp 0
transform 1 0 9490 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2020_
timestamp 0
transform -1 0 10390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2021_
timestamp 0
transform -1 0 7430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2022_
timestamp 0
transform 1 0 7670 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2023_
timestamp 0
transform -1 0 7970 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2024_
timestamp 0
transform 1 0 6190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2025_
timestamp 0
transform -1 0 6070 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2026_
timestamp 0
transform 1 0 9770 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2027_
timestamp 0
transform 1 0 10310 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2028_
timestamp 0
transform -1 0 10310 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2029_
timestamp 0
transform -1 0 11190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2030_
timestamp 0
transform 1 0 10810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2031_
timestamp 0
transform -1 0 11110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2032_
timestamp 0
transform 1 0 9030 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2033_
timestamp 0
transform 1 0 8490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2034_
timestamp 0
transform 1 0 8730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2035_
timestamp 0
transform 1 0 8690 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2036_
timestamp 0
transform 1 0 11650 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2037_
timestamp 0
transform 1 0 11850 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2038_
timestamp 0
transform -1 0 7690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2039_
timestamp 0
transform -1 0 6770 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2040_
timestamp 0
transform 1 0 11030 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2041_
timestamp 0
transform 1 0 11110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2042_
timestamp 0
transform -1 0 10190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2043_
timestamp 0
transform -1 0 10570 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2044_
timestamp 0
transform -1 0 11090 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2045_
timestamp 0
transform -1 0 11430 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2046_
timestamp 0
transform 1 0 8910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2047_
timestamp 0
transform -1 0 9470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2048_
timestamp 0
transform 1 0 9270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2049_
timestamp 0
transform 1 0 9410 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2050_
timestamp 0
transform 1 0 9170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2051_
timestamp 0
transform 1 0 8870 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2052_
timestamp 0
transform 1 0 9150 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2053_
timestamp 0
transform -1 0 9710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2054_
timestamp 0
transform 1 0 9930 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2055_
timestamp 0
transform -1 0 6570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2056_
timestamp 0
transform -1 0 6150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2057_
timestamp 0
transform 1 0 10350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2058_
timestamp 0
transform -1 0 10090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2059_
timestamp 0
transform -1 0 10230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2060_
timestamp 0
transform -1 0 9990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2061_
timestamp 0
transform 1 0 10170 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2062_
timestamp 0
transform -1 0 9250 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2063_
timestamp 0
transform 1 0 8330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2064_
timestamp 0
transform -1 0 8010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2065_
timestamp 0
transform -1 0 8830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2066_
timestamp 0
transform 1 0 8810 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2067_
timestamp 0
transform -1 0 8070 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2068_
timestamp 0
transform -1 0 8350 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2069_
timestamp 0
transform 1 0 8070 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2070_
timestamp 0
transform -1 0 8370 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2071_
timestamp 0
transform -1 0 8650 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2072_
timestamp 0
transform 1 0 8870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2073_
timestamp 0
transform 1 0 9130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2074_
timestamp 0
transform 1 0 9350 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2075_
timestamp 0
transform -1 0 9650 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2076_
timestamp 0
transform 1 0 11310 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2077_
timestamp 0
transform -1 0 11370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2078_
timestamp 0
transform -1 0 11170 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2079_
timestamp 0
transform 1 0 11310 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2080_
timestamp 0
transform -1 0 11150 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2081_
timestamp 0
transform 1 0 11150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2082_
timestamp 0
transform 1 0 10410 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2083_
timestamp 0
transform 1 0 9670 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2084_
timestamp 0
transform 1 0 11690 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2085_
timestamp 0
transform 1 0 11110 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2086_
timestamp 0
transform 1 0 11610 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2087_
timestamp 0
transform 1 0 11630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2088_
timestamp 0
transform -1 0 12190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2089_
timestamp 0
transform 1 0 11910 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2090_
timestamp 0
transform 1 0 12090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2091_
timestamp 0
transform 1 0 9990 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2092_
timestamp 0
transform 1 0 10610 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2093_
timestamp 0
transform -1 0 11170 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2094_
timestamp 0
transform 1 0 11410 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2095_
timestamp 0
transform -1 0 11070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2096_
timestamp 0
transform 1 0 11590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2097_
timestamp 0
transform -1 0 11930 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2098_
timestamp 0
transform -1 0 12110 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2099_
timestamp 0
transform -1 0 11410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2100_
timestamp 0
transform 1 0 11370 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2101_
timestamp 0
transform -1 0 11330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2102_
timestamp 0
transform -1 0 11710 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2103_
timestamp 0
transform 1 0 12190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2104_
timestamp 0
transform 1 0 12190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2105_
timestamp 0
transform -1 0 11650 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2106_
timestamp 0
transform -1 0 11630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2107_
timestamp 0
transform -1 0 12190 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2108_
timestamp 0
transform 1 0 8930 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2109_
timestamp 0
transform 1 0 12190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2110_
timestamp 0
transform -1 0 12210 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2111_
timestamp 0
transform -1 0 12210 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2112_
timestamp 0
transform -1 0 12110 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2113_
timestamp 0
transform 1 0 11870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2114_
timestamp 0
transform 1 0 10650 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2115_
timestamp 0
transform -1 0 9390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2116_
timestamp 0
transform -1 0 10270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2117_
timestamp 0
transform -1 0 10870 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2118_
timestamp 0
transform -1 0 10830 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2119_
timestamp 0
transform 1 0 10730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2120_
timestamp 0
transform 1 0 10770 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2121_
timestamp 0
transform -1 0 10510 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2122_
timestamp 0
transform 1 0 10710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2123_
timestamp 0
transform -1 0 8210 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2124_
timestamp 0
transform -1 0 7910 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2125_
timestamp 0
transform -1 0 10270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2126_
timestamp 0
transform 1 0 10670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2127_
timestamp 0
transform -1 0 7090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2128_
timestamp 0
transform -1 0 9230 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2129_
timestamp 0
transform 1 0 7350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2130_
timestamp 0
transform -1 0 10970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2131_
timestamp 0
transform -1 0 8010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2132_
timestamp 0
transform 1 0 6790 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2133_
timestamp 0
transform -1 0 7090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2134_
timestamp 0
transform -1 0 7350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2135_
timestamp 0
transform -1 0 11230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2136_
timestamp 0
transform -1 0 11390 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2137_
timestamp 0
transform 1 0 11370 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2138_
timestamp 0
transform 1 0 11450 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2139_
timestamp 0
transform -1 0 11370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2140_
timestamp 0
transform -1 0 11090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2141_
timestamp 0
transform 1 0 10010 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2142_
timestamp 0
transform 1 0 10810 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2143_
timestamp 0
transform -1 0 10550 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2144_
timestamp 0
transform -1 0 11110 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2145_
timestamp 0
transform -1 0 5110 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2146_
timestamp 0
transform 1 0 9830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2147_
timestamp 0
transform 1 0 10390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2148_
timestamp 0
transform -1 0 6330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2149_
timestamp 0
transform 1 0 10110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2150_
timestamp 0
transform 1 0 8890 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2151_
timestamp 0
transform 1 0 7510 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2152_
timestamp 0
transform 1 0 8590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2153_
timestamp 0
transform 1 0 8850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2154_
timestamp 0
transform 1 0 9130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2155_
timestamp 0
transform -1 0 10210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2156_
timestamp 0
transform -1 0 10990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2157_
timestamp 0
transform 1 0 11230 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2158_
timestamp 0
transform -1 0 11810 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2159_
timestamp 0
transform -1 0 11930 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2160_
timestamp 0
transform -1 0 11470 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2161_
timestamp 0
transform 1 0 8210 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2162_
timestamp 0
transform 1 0 8970 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2163_
timestamp 0
transform -1 0 10070 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2164_
timestamp 0
transform 1 0 9830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2165_
timestamp 0
transform 1 0 11070 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2166_
timestamp 0
transform 1 0 10890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2167_
timestamp 0
transform 1 0 9270 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2168_
timestamp 0
transform 1 0 10090 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2169_
timestamp 0
transform -1 0 8830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2170_
timestamp 0
transform -1 0 9250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2171_
timestamp 0
transform 1 0 10390 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2172_
timestamp 0
transform 1 0 9810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2173_
timestamp 0
transform 1 0 9930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2174_
timestamp 0
transform -1 0 9570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2175_
timestamp 0
transform 1 0 9650 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2176_
timestamp 0
transform -1 0 9770 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2177_
timestamp 0
transform -1 0 9470 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2178_
timestamp 0
transform -1 0 11070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2179_
timestamp 0
transform 1 0 9550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2180_
timestamp 0
transform 1 0 11910 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2181_
timestamp 0
transform 1 0 11890 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2182_
timestamp 0
transform 1 0 11970 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2183_
timestamp 0
transform -1 0 11350 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2184_
timestamp 0
transform 1 0 11090 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2185_
timestamp 0
transform -1 0 10330 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2186_
timestamp 0
transform 1 0 10270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2187_
timestamp 0
transform -1 0 10670 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2188_
timestamp 0
transform 1 0 11630 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2189_
timestamp 0
transform 1 0 10010 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2190_
timestamp 0
transform 1 0 10570 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2191_
timestamp 0
transform 1 0 11190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2192_
timestamp 0
transform 1 0 11130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2193_
timestamp 0
transform -1 0 11070 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2194_
timestamp 0
transform -1 0 10630 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2195_
timestamp 0
transform -1 0 9510 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2196_
timestamp 0
transform -1 0 11150 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2197_
timestamp 0
transform 1 0 11410 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2198_
timestamp 0
transform -1 0 9950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2199_
timestamp 0
transform -1 0 10010 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2200_
timestamp 0
transform -1 0 5870 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2201_
timestamp 0
transform 1 0 6390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2202_
timestamp 0
transform 1 0 6130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2203_
timestamp 0
transform 1 0 6130 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2204_
timestamp 0
transform 1 0 6870 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2205_
timestamp 0
transform 1 0 7170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2206_
timestamp 0
transform 1 0 9510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2207_
timestamp 0
transform -1 0 10010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2208_
timestamp 0
transform -1 0 9430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2209_
timestamp 0
transform 1 0 10470 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2210_
timestamp 0
transform 1 0 10470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2211_
timestamp 0
transform 1 0 11310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2212_
timestamp 0
transform -1 0 11670 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2213_
timestamp 0
transform -1 0 11710 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2214_
timestamp 0
transform 1 0 11670 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2215_
timestamp 0
transform 1 0 11770 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2216_
timestamp 0
transform 1 0 12150 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2217_
timestamp 0
transform 1 0 11430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2218_
timestamp 0
transform 1 0 9710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2219_
timestamp 0
transform -1 0 9950 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2220_
timestamp 0
transform -1 0 9990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2221_
timestamp 0
transform -1 0 11930 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2222_
timestamp 0
transform 1 0 11870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2223_
timestamp 0
transform -1 0 11910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2224_
timestamp 0
transform 1 0 11890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2225_
timestamp 0
transform 1 0 10990 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2226_
timestamp 0
transform 1 0 11950 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2227_
timestamp 0
transform 1 0 11670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2228_
timestamp 0
transform -1 0 11530 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2229_
timestamp 0
transform -1 0 10610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2230_
timestamp 0
transform -1 0 10330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2231_
timestamp 0
transform -1 0 8530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2232_
timestamp 0
transform 1 0 8770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2233_
timestamp 0
transform 1 0 9550 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2234_
timestamp 0
transform -1 0 9810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2235_
timestamp 0
transform -1 0 9930 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2236_
timestamp 0
transform 1 0 7230 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2237_
timestamp 0
transform -1 0 6710 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2238_
timestamp 0
transform -1 0 6990 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2239_
timestamp 0
transform -1 0 9010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2240_
timestamp 0
transform -1 0 8730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2241_
timestamp 0
transform -1 0 8370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2242_
timestamp 0
transform -1 0 7550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2243_
timestamp 0
transform 1 0 7810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2244_
timestamp 0
transform 1 0 8090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2245_
timestamp 0
transform -1 0 7790 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2246_
timestamp 0
transform 1 0 9170 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2247_
timestamp 0
transform -1 0 12170 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2248_
timestamp 0
transform 1 0 11370 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2249_
timestamp 0
transform -1 0 9530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2250_
timestamp 0
transform 1 0 11050 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2251_
timestamp 0
transform 1 0 10610 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2252_
timestamp 0
transform 1 0 11350 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2253_
timestamp 0
transform -1 0 11950 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2254_
timestamp 0
transform 1 0 12190 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2255_
timestamp 0
transform -1 0 10550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2256_
timestamp 0
transform -1 0 10830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2257_
timestamp 0
transform 1 0 11070 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2258_
timestamp 0
transform 1 0 12230 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2259_
timestamp 0
transform -1 0 11910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2260_
timestamp 0
transform 1 0 10090 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2261_
timestamp 0
transform 1 0 10350 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2262_
timestamp 0
transform -1 0 10870 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2263_
timestamp 0
transform 1 0 11350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2264_
timestamp 0
transform 1 0 12170 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2265_
timestamp 0
transform -1 0 11430 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2266_
timestamp 0
transform -1 0 10790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2267_
timestamp 0
transform 1 0 12010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2268_
timestamp 0
transform 1 0 12170 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2269_
timestamp 0
transform -1 0 11950 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2270_
timestamp 0
transform 1 0 11370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2271_
timestamp 0
transform -1 0 11670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2272_
timestamp 0
transform 1 0 11930 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2273_
timestamp 0
transform -1 0 12190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2274_
timestamp 0
transform 1 0 10110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2275_
timestamp 0
transform -1 0 8270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2276_
timestamp 0
transform 1 0 8930 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2277_
timestamp 0
transform 1 0 9210 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2278_
timestamp 0
transform -1 0 9290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2279_
timestamp 0
transform 1 0 9090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2280_
timestamp 0
transform 1 0 10250 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2281_
timestamp 0
transform 1 0 12130 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2282_
timestamp 0
transform 1 0 12190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2283_
timestamp 0
transform -1 0 11070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2284_
timestamp 0
transform 1 0 12150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2285_
timestamp 0
transform 1 0 12150 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2286_
timestamp 0
transform -1 0 11930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2287_
timestamp 0
transform 1 0 11870 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2288_
timestamp 0
transform -1 0 11030 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2289_
timestamp 0
transform -1 0 10810 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2290_
timestamp 0
transform -1 0 10990 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2291_
timestamp 0
transform 1 0 11350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2292_
timestamp 0
transform 1 0 10490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2293_
timestamp 0
transform 1 0 10770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2294_
timestamp 0
transform 1 0 11090 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2295_
timestamp 0
transform 1 0 10970 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2296_
timestamp 0
transform 1 0 11230 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2297_
timestamp 0
transform 1 0 11890 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2298_
timestamp 0
transform -1 0 11990 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2299_
timestamp 0
transform -1 0 10550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2300_
timestamp 0
transform 1 0 10250 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2301_
timestamp 0
transform 1 0 11870 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2302_
timestamp 0
transform 1 0 11810 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2303_
timestamp 0
transform -1 0 11790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2304_
timestamp 0
transform 1 0 11930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2305_
timestamp 0
transform 1 0 10810 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2306_
timestamp 0
transform -1 0 11670 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2307_
timestamp 0
transform 1 0 11370 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2308_
timestamp 0
transform 1 0 12150 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2309_
timestamp 0
transform -1 0 11710 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2310_
timestamp 0
transform -1 0 11650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2311_
timestamp 0
transform 1 0 11630 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2312_
timestamp 0
transform 1 0 11690 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2313_
timestamp 0
transform 1 0 11970 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2314_
timestamp 0
transform -1 0 11290 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2315_
timestamp 0
transform 1 0 12150 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2316_
timestamp 0
transform 1 0 11550 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2317_
timestamp 0
transform -1 0 12050 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2318_
timestamp 0
transform 1 0 11590 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2319_
timestamp 0
transform 1 0 11230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2320_
timestamp 0
transform 1 0 11650 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2321_
timestamp 0
transform 1 0 11510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2322_
timestamp 0
transform -1 0 11370 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2323_
timestamp 0
transform -1 0 11610 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2324_
timestamp 0
transform 1 0 11850 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2325_
timestamp 0
transform -1 0 12230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2326_
timestamp 0
transform 1 0 12150 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2327_
timestamp 0
transform 1 0 11510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2328_
timestamp 0
transform 1 0 11090 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2329_
timestamp 0
transform 1 0 8610 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2330_
timestamp 0
transform -1 0 10290 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2331_
timestamp 0
transform -1 0 9730 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2332_
timestamp 0
transform -1 0 11950 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2333_
timestamp 0
transform -1 0 10830 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2334_
timestamp 0
transform 1 0 10550 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2335_
timestamp 0
transform 1 0 10530 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2336_
timestamp 0
transform 1 0 10710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2337_
timestamp 0
transform -1 0 10830 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2338_
timestamp 0
transform -1 0 10750 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2339_
timestamp 0
transform -1 0 9670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2340_
timestamp 0
transform -1 0 9950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2341_
timestamp 0
transform 1 0 9650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2342_
timestamp 0
transform -1 0 10530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2343_
timestamp 0
transform -1 0 10470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2344_
timestamp 0
transform -1 0 10710 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2345_
timestamp 0
transform 1 0 11830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2346_
timestamp 0
transform 1 0 11570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2347_
timestamp 0
transform -1 0 8910 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2348_
timestamp 0
transform -1 0 10010 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2349_
timestamp 0
transform -1 0 11670 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2350_
timestamp 0
transform -1 0 11390 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2351_
timestamp 0
transform -1 0 10450 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2352_
timestamp 0
transform -1 0 10210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2353_
timestamp 0
transform -1 0 9510 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2354_
timestamp 0
transform 1 0 7910 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2355_
timestamp 0
transform -1 0 6990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2356_
timestamp 0
transform -1 0 6930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2357_
timestamp 0
transform -1 0 7590 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2358_
timestamp 0
transform -1 0 7170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2359_
timestamp 0
transform 1 0 7390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2360_
timestamp 0
transform -1 0 8070 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2361_
timestamp 0
transform -1 0 7130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2362_
timestamp 0
transform 1 0 8850 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2363_
timestamp 0
transform -1 0 7530 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2364_
timestamp 0
transform 1 0 7270 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2365_
timestamp 0
transform 1 0 6990 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2366_
timestamp 0
transform 1 0 6470 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2367_
timestamp 0
transform -1 0 7310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2368_
timestamp 0
transform 1 0 6710 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2369_
timestamp 0
transform 1 0 7090 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2370_
timestamp 0
transform -1 0 7350 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2371_
timestamp 0
transform 1 0 7290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2372_
timestamp 0
transform -1 0 6870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2373_
timestamp 0
transform 1 0 6810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2374_
timestamp 0
transform 1 0 8310 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2375_
timestamp 0
transform 1 0 8370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2376_
timestamp 0
transform -1 0 6810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2377_
timestamp 0
transform 1 0 5510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2378_
timestamp 0
transform -1 0 3830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2379_
timestamp 0
transform -1 0 8090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2380_
timestamp 0
transform -1 0 5730 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2381_
timestamp 0
transform -1 0 6010 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2382_
timestamp 0
transform -1 0 5870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2383_
timestamp 0
transform 1 0 4790 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2384_
timestamp 0
transform 1 0 4710 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2385_
timestamp 0
transform 1 0 4950 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2386_
timestamp 0
transform 1 0 5230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2387_
timestamp 0
transform 1 0 1750 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2388_
timestamp 0
transform 1 0 1690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2389_
timestamp 0
transform 1 0 5270 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2390_
timestamp 0
transform 1 0 2550 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2391_
timestamp 0
transform -1 0 2350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2392_
timestamp 0
transform -1 0 2070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2393_
timestamp 0
transform -1 0 2630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2394_
timestamp 0
transform -1 0 3050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2395_
timestamp 0
transform 1 0 4450 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2396_
timestamp 0
transform 1 0 3090 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2397_
timestamp 0
transform -1 0 3170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2398_
timestamp 0
transform -1 0 2890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2399_
timestamp 0
transform 1 0 1990 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2400_
timestamp 0
transform -1 0 1430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2401_
timestamp 0
transform -1 0 2910 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2402_
timestamp 0
transform 1 0 2650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2403_
timestamp 0
transform -1 0 2290 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2404_
timestamp 0
transform -1 0 1730 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2405_
timestamp 0
transform -1 0 1590 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2406_
timestamp 0
transform 1 0 5970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2407_
timestamp 0
transform -1 0 4330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2408_
timestamp 0
transform -1 0 5690 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2409_
timestamp 0
transform -1 0 6510 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2410_
timestamp 0
transform -1 0 4290 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2411_
timestamp 0
transform -1 0 4050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2412_
timestamp 0
transform -1 0 1310 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2413_
timestamp 0
transform -1 0 4590 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2414_
timestamp 0
transform 1 0 3110 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2415_
timestamp 0
transform -1 0 2850 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2416_
timestamp 0
transform 1 0 1810 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2417_
timestamp 0
transform -1 0 2310 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2418_
timestamp 0
transform -1 0 2190 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2419_
timestamp 0
transform -1 0 3510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2420_
timestamp 0
transform 1 0 2930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2421_
timestamp 0
transform -1 0 2850 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2422_
timestamp 0
transform -1 0 2030 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2423_
timestamp 0
transform -1 0 3730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2424_
timestamp 0
transform -1 0 3570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2425_
timestamp 0
transform -1 0 3450 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2426_
timestamp 0
transform 1 0 3210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2427_
timestamp 0
transform 1 0 3370 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2428_
timestamp 0
transform -1 0 3450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2429_
timestamp 0
transform -1 0 5170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2430_
timestamp 0
transform -1 0 7870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2431_
timestamp 0
transform -1 0 5430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2432_
timestamp 0
transform -1 0 9550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2433_
timestamp 0
transform 1 0 11650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2434_
timestamp 0
transform 1 0 10830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2435_
timestamp 0
transform -1 0 7310 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2436_
timestamp 0
transform -1 0 6990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2437_
timestamp 0
transform -1 0 9670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2438_
timestamp 0
transform -1 0 9410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2439_
timestamp 0
transform -1 0 6190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2440_
timestamp 0
transform 1 0 7810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2441_
timestamp 0
transform -1 0 7650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2442_
timestamp 0
transform 1 0 10350 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2443_
timestamp 0
transform -1 0 7250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2444_
timestamp 0
transform -1 0 7250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2445_
timestamp 0
transform 1 0 5350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2446_
timestamp 0
transform 1 0 6470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2447_
timestamp 0
transform -1 0 4850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2448_
timestamp 0
transform -1 0 6450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2449_
timestamp 0
transform -1 0 7070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2450_
timestamp 0
transform 1 0 4210 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2451_
timestamp 0
transform -1 0 4090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2452_
timestamp 0
transform 1 0 4730 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2453_
timestamp 0
transform 1 0 8590 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2454_
timestamp 0
transform 1 0 4470 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2455_
timestamp 0
transform 1 0 4470 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2456_
timestamp 0
transform -1 0 4330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2457_
timestamp 0
transform -1 0 4590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2458_
timestamp 0
transform -1 0 4950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2459_
timestamp 0
transform 1 0 5090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2460_
timestamp 0
transform 1 0 4970 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2461_
timestamp 0
transform 1 0 5250 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2462_
timestamp 0
transform 1 0 5390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2463_
timestamp 0
transform 1 0 6330 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2464_
timestamp 0
transform -1 0 3270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2465_
timestamp 0
transform -1 0 2990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2466_
timestamp 0
transform -1 0 2990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2467_
timestamp 0
transform 1 0 2130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2468_
timestamp 0
transform -1 0 1690 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2469_
timestamp 0
transform 1 0 650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2470_
timestamp 0
transform -1 0 2750 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2471_
timestamp 0
transform -1 0 2770 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2472_
timestamp 0
transform -1 0 2470 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2473_
timestamp 0
transform 1 0 1970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2474_
timestamp 0
transform -1 0 1490 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2475_
timestamp 0
transform -1 0 430 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2476_
timestamp 0
transform -1 0 3850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2477_
timestamp 0
transform -1 0 5090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2478_
timestamp 0
transform 1 0 3950 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2479_
timestamp 0
transform -1 0 3590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2480_
timestamp 0
transform 1 0 1830 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2481_
timestamp 0
transform -1 0 3390 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2482_
timestamp 0
transform 1 0 3670 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2483_
timestamp 0
transform 1 0 3090 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2484_
timestamp 0
transform 1 0 2810 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2485_
timestamp 0
transform -1 0 430 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2486_
timestamp 0
transform -1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2487_
timestamp 0
transform 1 0 2430 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2488_
timestamp 0
transform -1 0 2430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2489_
timestamp 0
transform -1 0 1870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2490_
timestamp 0
transform -1 0 1430 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2491_
timestamp 0
transform -1 0 430 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2492_
timestamp 0
transform 1 0 4650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2493_
timestamp 0
transform 1 0 3650 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2494_
timestamp 0
transform 1 0 6230 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2495_
timestamp 0
transform 1 0 3890 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2496_
timestamp 0
transform 1 0 4190 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2497_
timestamp 0
transform -1 0 4110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2498_
timestamp 0
transform 1 0 3570 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2499_
timestamp 0
transform 1 0 3830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2500_
timestamp 0
transform -1 0 430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2501_
timestamp 0
transform -1 0 3430 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2502_
timestamp 0
transform -1 0 3070 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2503_
timestamp 0
transform -1 0 3550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__2504_
timestamp 0
transform -1 0 3310 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__2505_
timestamp 0
transform 1 0 2750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2506_
timestamp 0
transform -1 0 2570 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__2507_
timestamp 0
transform 1 0 690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2508_
timestamp 0
transform 1 0 3190 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2509_
timestamp 0
transform 1 0 2730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2510_
timestamp 0
transform -1 0 3290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2511_
timestamp 0
transform 1 0 3370 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__2512_
timestamp 0
transform 1 0 3210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2513_
timestamp 0
transform -1 0 2470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2514_
timestamp 0
transform 1 0 2170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2515_
timestamp 0
transform -1 0 2190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2516_
timestamp 0
transform -1 0 430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__2517_
timestamp 0
transform -1 0 2270 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2518_
timestamp 0
transform 1 0 5370 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2519_
timestamp 0
transform -1 0 5910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2520_
timestamp 0
transform -1 0 6010 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2521_
timestamp 0
transform 1 0 5710 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2522_
timestamp 0
transform -1 0 5710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2523_
timestamp 0
transform -1 0 5630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2524_
timestamp 0
transform -1 0 5570 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2525_
timestamp 0
transform -1 0 2790 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2526_
timestamp 0
transform 1 0 6190 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2527_
timestamp 0
transform 1 0 6590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2528_
timestamp 0
transform 1 0 6570 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2529_
timestamp 0
transform 1 0 6170 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2530_
timestamp 0
transform 1 0 5630 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2531_
timestamp 0
transform 1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2532_
timestamp 0
transform 1 0 4270 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2533_
timestamp 0
transform 1 0 5210 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2534_
timestamp 0
transform 1 0 4930 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2535_
timestamp 0
transform -1 0 4670 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2536_
timestamp 0
transform 1 0 3510 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2537_
timestamp 0
transform 1 0 2150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2538_
timestamp 0
transform 1 0 4550 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2539_
timestamp 0
transform 1 0 3930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2540_
timestamp 0
transform 1 0 4270 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2541_
timestamp 0
transform -1 0 4250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2542_
timestamp 0
transform -1 0 3770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2543_
timestamp 0
transform 1 0 3530 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2544_
timestamp 0
transform 1 0 4250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2545_
timestamp 0
transform 1 0 4510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2546_
timestamp 0
transform 1 0 4870 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2547_
timestamp 0
transform -1 0 4810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2548_
timestamp 0
transform -1 0 4530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2549_
timestamp 0
transform 1 0 4750 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2550_
timestamp 0
transform 1 0 4750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2551_
timestamp 0
transform 1 0 5270 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2552_
timestamp 0
transform 1 0 5510 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2553_
timestamp 0
transform 1 0 2410 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2554_
timestamp 0
transform 1 0 4550 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2555_
timestamp 0
transform -1 0 4730 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2556_
timestamp 0
transform -1 0 4970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2557_
timestamp 0
transform 1 0 4670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2558_
timestamp 0
transform 1 0 4750 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2559_
timestamp 0
transform 1 0 4470 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2560_
timestamp 0
transform 1 0 3970 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2561_
timestamp 0
transform 1 0 3670 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2562_
timestamp 0
transform 1 0 2290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2563_
timestamp 0
transform -1 0 4510 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2564_
timestamp 0
transform 1 0 4430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2565_
timestamp 0
transform -1 0 3910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2566_
timestamp 0
transform 1 0 2510 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2567_
timestamp 0
transform 1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2568_
timestamp 0
transform -1 0 5790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2569_
timestamp 0
transform -1 0 5930 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2570_
timestamp 0
transform 1 0 6010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2571_
timestamp 0
transform 1 0 6010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2572_
timestamp 0
transform 1 0 5870 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2573_
timestamp 0
transform 1 0 5790 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2574_
timestamp 0
transform 1 0 5770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2575_
timestamp 0
transform -1 0 4810 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2576_
timestamp 0
transform -1 0 4290 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2577_
timestamp 0
transform -1 0 4550 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2578_
timestamp 0
transform 1 0 7050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2579_
timestamp 0
transform 1 0 7070 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2580_
timestamp 0
transform 1 0 8070 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2581_
timestamp 0
transform -1 0 8930 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2582_
timestamp 0
transform 1 0 6970 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2583_
timestamp 0
transform -1 0 6970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2584_
timestamp 0
transform 1 0 7390 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2585_
timestamp 0
transform 1 0 7430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2586_
timestamp 0
transform -1 0 8510 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2587_
timestamp 0
transform -1 0 6850 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2588_
timestamp 0
transform -1 0 5890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2589_
timestamp 0
transform 1 0 7510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2590_
timestamp 0
transform -1 0 6290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2591_
timestamp 0
transform 1 0 6530 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2592_
timestamp 0
transform -1 0 4510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2593_
timestamp 0
transform 1 0 5030 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2594_
timestamp 0
transform -1 0 8610 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2595_
timestamp 0
transform -1 0 5330 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2596_
timestamp 0
transform 1 0 5330 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2597_
timestamp 0
transform 1 0 5510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2598_
timestamp 0
transform -1 0 5250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2599_
timestamp 0
transform -1 0 5050 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2600_
timestamp 0
transform -1 0 5050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2601_
timestamp 0
transform -1 0 5310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2602_
timestamp 0
transform -1 0 8250 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2603_
timestamp 0
transform -1 0 6690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2604_
timestamp 0
transform -1 0 6450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2605_
timestamp 0
transform 1 0 6130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2606_
timestamp 0
transform -1 0 5630 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2607_
timestamp 0
transform 1 0 5790 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2608_
timestamp 0
transform 1 0 5610 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2609_
timestamp 0
transform -1 0 5590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2610_
timestamp 0
transform 1 0 4970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2611_
timestamp 0
transform -1 0 5230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2612_
timestamp 0
transform -1 0 5490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2613_
timestamp 0
transform -1 0 1310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2614_
timestamp 0
transform 1 0 2290 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2615_
timestamp 0
transform -1 0 2570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2616_
timestamp 0
transform -1 0 2550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2617_
timestamp 0
transform 1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2618_
timestamp 0
transform 1 0 950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2619_
timestamp 0
transform -1 0 450 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2620_
timestamp 0
transform -1 0 690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2621_
timestamp 0
transform 1 0 1010 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2622_
timestamp 0
transform 1 0 450 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2623_
timestamp 0
transform 1 0 2830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2624_
timestamp 0
transform 1 0 2030 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2625_
timestamp 0
transform -1 0 2290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2626_
timestamp 0
transform -1 0 2010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2627_
timestamp 0
transform 1 0 150 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2628_
timestamp 0
transform 1 0 150 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2629_
timestamp 0
transform -1 0 410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2630_
timestamp 0
transform 1 0 150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2631_
timestamp 0
transform 1 0 5090 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2632_
timestamp 0
transform 1 0 2330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2633_
timestamp 0
transform -1 0 2630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2634_
timestamp 0
transform -1 0 170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2635_
timestamp 0
transform 1 0 150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2636_
timestamp 0
transform 1 0 690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2637_
timestamp 0
transform 1 0 1030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2638_
timestamp 0
transform 1 0 450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2639_
timestamp 0
transform -1 0 770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2640_
timestamp 0
transform -1 0 170 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2641_
timestamp 0
transform -1 0 170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2642_
timestamp 0
transform 1 0 1410 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2643_
timestamp 0
transform -1 0 1950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2644_
timestamp 0
transform 1 0 2350 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2645_
timestamp 0
transform -1 0 2090 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2646_
timestamp 0
transform -1 0 1290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2647_
timestamp 0
transform 1 0 150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2648_
timestamp 0
transform 1 0 650 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__2649_
timestamp 0
transform 1 0 150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2650_
timestamp 0
transform -1 0 3750 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2651_
timestamp 0
transform -1 0 3470 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2652_
timestamp 0
transform 1 0 690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2653_
timestamp 0
transform 1 0 410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2654_
timestamp 0
transform 1 0 1290 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2655_
timestamp 0
transform 1 0 730 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2656_
timestamp 0
transform -1 0 1010 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2657_
timestamp 0
transform 1 0 150 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2658_
timestamp 0
transform 1 0 150 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2659_
timestamp 0
transform -1 0 450 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2660_
timestamp 0
transform 1 0 390 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2661_
timestamp 0
transform -1 0 2710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__2662_
timestamp 0
transform -1 0 2650 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2663_
timestamp 0
transform -1 0 2070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2664_
timestamp 0
transform 1 0 970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2665_
timestamp 0
transform -1 0 930 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2666_
timestamp 0
transform -1 0 450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2667_
timestamp 0
transform -1 0 670 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2668_
timestamp 0
transform 1 0 1170 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2669_
timestamp 0
transform -1 0 2930 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2670_
timestamp 0
transform -1 0 3050 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2671_
timestamp 0
transform 1 0 1210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2672_
timestamp 0
transform -1 0 710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2673_
timestamp 0
transform -1 0 670 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2674_
timestamp 0
transform 1 0 930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2675_
timestamp 0
transform 1 0 910 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2676_
timestamp 0
transform -1 0 1210 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2677_
timestamp 0
transform 1 0 6550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__2678_
timestamp 0
transform -1 0 6470 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2679_
timestamp 0
transform 1 0 7090 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2680_
timestamp 0
transform -1 0 6890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2681_
timestamp 0
transform 1 0 7150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2682_
timestamp 0
transform -1 0 6870 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2683_
timestamp 0
transform -1 0 1990 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2684_
timestamp 0
transform -1 0 1810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__2685_
timestamp 0
transform 1 0 1730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2686_
timestamp 0
transform 1 0 1730 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2687_
timestamp 0
transform 1 0 1470 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2688_
timestamp 0
transform -1 0 910 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2689_
timestamp 0
transform -1 0 890 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2690_
timestamp 0
transform 1 0 7390 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2691_
timestamp 0
transform -1 0 7230 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2692_
timestamp 0
transform -1 0 5170 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2693_
timestamp 0
transform -1 0 3130 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2694_
timestamp 0
transform -1 0 1430 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2695_
timestamp 0
transform -1 0 1710 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2696_
timestamp 0
transform -1 0 1430 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2697_
timestamp 0
transform 1 0 2010 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2698_
timestamp 0
transform -1 0 650 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2699_
timestamp 0
transform 1 0 6410 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2700_
timestamp 0
transform -1 0 7130 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2701_
timestamp 0
transform 1 0 7710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2702_
timestamp 0
transform 1 0 7410 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2703_
timestamp 0
transform 1 0 7570 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2704_
timestamp 0
transform -1 0 6770 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2705_
timestamp 0
transform 1 0 1690 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2706_
timestamp 0
transform 1 0 1130 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2707_
timestamp 0
transform 1 0 2830 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2708_
timestamp 0
transform 1 0 2510 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2709_
timestamp 0
transform -1 0 1190 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2710_
timestamp 0
transform -1 0 970 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2711_
timestamp 0
transform -1 0 1250 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2712_
timestamp 0
transform 1 0 2990 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2713_
timestamp 0
transform -1 0 4390 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2714_
timestamp 0
transform -1 0 4810 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2715_
timestamp 0
transform 1 0 3650 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2716_
timestamp 0
transform -1 0 4410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2717_
timestamp 0
transform -1 0 5970 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__2718_
timestamp 0
transform -1 0 4210 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2719_
timestamp 0
transform 1 0 3810 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2720_
timestamp 0
transform -1 0 4110 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2721_
timestamp 0
transform -1 0 2270 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2722_
timestamp 0
transform 1 0 2390 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2723_
timestamp 0
transform 1 0 2690 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2724_
timestamp 0
transform -1 0 930 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2725_
timestamp 0
transform -1 0 5530 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2726_
timestamp 0
transform -1 0 6710 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2727_
timestamp 0
transform 1 0 3970 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2728_
timestamp 0
transform 1 0 3690 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2729_
timestamp 0
transform -1 0 3650 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2730_
timestamp 0
transform 1 0 3250 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2731_
timestamp 0
transform 1 0 2110 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2732_
timestamp 0
transform -1 0 1990 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2733_
timestamp 0
transform 1 0 1530 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2734_
timestamp 0
transform -1 0 1830 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2735_
timestamp 0
transform -1 0 3990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2736_
timestamp 0
transform -1 0 4130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2737_
timestamp 0
transform -1 0 4210 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2738_
timestamp 0
transform -1 0 3910 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2739_
timestamp 0
transform -1 0 3350 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2740_
timestamp 0
transform -1 0 3430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2741_
timestamp 0
transform -1 0 1190 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2742_
timestamp 0
transform 1 0 1490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2743_
timestamp 0
transform 1 0 1430 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2744_
timestamp 0
transform 1 0 1970 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2745_
timestamp 0
transform 1 0 630 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2746_
timestamp 0
transform 1 0 3690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2747_
timestamp 0
transform 1 0 4810 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__2748_
timestamp 0
transform 1 0 4470 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2749_
timestamp 0
transform -1 0 3630 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2750_
timestamp 0
transform -1 0 3070 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2751_
timestamp 0
transform 1 0 2910 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2752_
timestamp 0
transform 1 0 1210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2753_
timestamp 0
transform 1 0 710 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2754_
timestamp 0
transform -1 0 650 0 1 790
box -6 -8 26 268
use FILL  FILL_7__2755_
timestamp 0
transform -1 0 3170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2756_
timestamp 0
transform -1 0 2610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2757_
timestamp 0
transform 1 0 2850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2758_
timestamp 0
transform 1 0 2330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2759_
timestamp 0
transform -1 0 4410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2760_
timestamp 0
transform 1 0 3850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2761_
timestamp 0
transform 1 0 4190 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2762_
timestamp 0
transform -1 0 3930 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2763_
timestamp 0
transform -1 0 2170 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2764_
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2765_
timestamp 0
transform -1 0 1810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2766_
timestamp 0
transform -1 0 2070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__2767_
timestamp 0
transform -1 0 1590 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__2768_
timestamp 0
transform 1 0 2250 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2769_
timestamp 0
transform 1 0 1690 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__2770_
timestamp 0
transform 1 0 6050 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2771_
timestamp 0
transform 1 0 6590 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2772_
timestamp 0
transform 1 0 5030 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__2773_
timestamp 0
transform 1 0 4230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2774_
timestamp 0
transform 1 0 2390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2775_
timestamp 0
transform 1 0 2630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2776_
timestamp 0
transform 1 0 3450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2777_
timestamp 0
transform -1 0 2930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2778_
timestamp 0
transform -1 0 3190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__2779_
timestamp 0
transform -1 0 7230 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2780_
timestamp 0
transform -1 0 7470 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__2781_
timestamp 0
transform 1 0 7950 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__2782_
timestamp 0
transform 1 0 7830 0 1 270
box -6 -8 26 268
use FILL  FILL_7__2783_
timestamp 0
transform 1 0 9770 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2784_
timestamp 0
transform 1 0 10910 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2785_
timestamp 0
transform 1 0 10290 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2786_
timestamp 0
transform 1 0 10010 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2787_
timestamp 0
transform 1 0 8470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2788_
timestamp 0
transform 1 0 8730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2789_
timestamp 0
transform 1 0 8250 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2790_
timestamp 0
transform -1 0 7990 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2791_
timestamp 0
transform 1 0 6250 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2792_
timestamp 0
transform 1 0 9870 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2793_
timestamp 0
transform 1 0 10070 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2794_
timestamp 0
transform -1 0 10330 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2795_
timestamp 0
transform 1 0 8510 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2796_
timestamp 0
transform 1 0 8490 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2797_
timestamp 0
transform 1 0 10890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2798_
timestamp 0
transform -1 0 10030 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2799_
timestamp 0
transform -1 0 8410 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2800_
timestamp 0
transform -1 0 7810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2801_
timestamp 0
transform 1 0 9750 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2802_
timestamp 0
transform -1 0 10070 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2803_
timestamp 0
transform 1 0 8510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2804_
timestamp 0
transform -1 0 8410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2805_
timestamp 0
transform -1 0 10150 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2806_
timestamp 0
transform 1 0 9830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2807_
timestamp 0
transform -1 0 8450 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2808_
timestamp 0
transform -1 0 6690 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2809_
timestamp 0
transform 1 0 8210 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2810_
timestamp 0
transform -1 0 7630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2811_
timestamp 0
transform 1 0 10110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2812_
timestamp 0
transform 1 0 9750 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2813_
timestamp 0
transform 1 0 8330 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2814_
timestamp 0
transform -1 0 8210 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2815_
timestamp 0
transform -1 0 8290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2816_
timestamp 0
transform 1 0 9550 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2817_
timestamp 0
transform -1 0 10410 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2818_
timestamp 0
transform 1 0 11230 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2819_
timestamp 0
transform 1 0 10210 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2820_
timestamp 0
transform -1 0 9990 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2821_
timestamp 0
transform -1 0 9850 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2822_
timestamp 0
transform -1 0 7570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2823_
timestamp 0
transform -1 0 9570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2824_
timestamp 0
transform -1 0 9310 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2825_
timestamp 0
transform 1 0 8770 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2826_
timestamp 0
transform 1 0 8810 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2827_
timestamp 0
transform 1 0 9230 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2828_
timestamp 0
transform 1 0 10350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2829_
timestamp 0
transform -1 0 9290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2830_
timestamp 0
transform 1 0 9910 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2831_
timestamp 0
transform 1 0 9090 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2832_
timestamp 0
transform -1 0 9010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2833_
timestamp 0
transform -1 0 8770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2834_
timestamp 0
transform -1 0 8350 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2835_
timestamp 0
transform -1 0 9370 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2836_
timestamp 0
transform -1 0 8070 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2837_
timestamp 0
transform 1 0 8150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2838_
timestamp 0
transform 1 0 9390 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2839_
timestamp 0
transform 1 0 9650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2840_
timestamp 0
transform -1 0 9390 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2841_
timestamp 0
transform 1 0 8290 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2842_
timestamp 0
transform 1 0 11610 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2843_
timestamp 0
transform -1 0 11110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2844_
timestamp 0
transform 1 0 10830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2845_
timestamp 0
transform 1 0 10570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2846_
timestamp 0
transform -1 0 10210 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2847_
timestamp 0
transform 1 0 10410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2848_
timestamp 0
transform -1 0 9690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2849_
timestamp 0
transform 1 0 10990 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__2850_
timestamp 0
transform 1 0 11150 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2851_
timestamp 0
transform 1 0 11390 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2852_
timestamp 0
transform 1 0 12090 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2853_
timestamp 0
transform 1 0 12150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2854_
timestamp 0
transform 1 0 11830 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2855_
timestamp 0
transform 1 0 12110 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2856_
timestamp 0
transform -1 0 9150 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2857_
timestamp 0
transform 1 0 9650 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2858_
timestamp 0
transform -1 0 9950 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2859_
timestamp 0
transform 1 0 10890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2860_
timestamp 0
transform 1 0 7770 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2861_
timestamp 0
transform 1 0 8450 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2862_
timestamp 0
transform -1 0 7830 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2863_
timestamp 0
transform 1 0 7530 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2864_
timestamp 0
transform 1 0 9770 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2865_
timestamp 0
transform 1 0 8930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2866_
timestamp 0
transform -1 0 7030 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2867_
timestamp 0
transform -1 0 8870 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2868_
timestamp 0
transform -1 0 8590 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2869_
timestamp 0
transform -1 0 9030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2870_
timestamp 0
transform 1 0 8670 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2871_
timestamp 0
transform 1 0 8630 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2872_
timestamp 0
transform 1 0 5570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2873_
timestamp 0
transform -1 0 5590 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2874_
timestamp 0
transform 1 0 5510 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2875_
timestamp 0
transform -1 0 5870 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2876_
timestamp 0
transform 1 0 5550 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2877_
timestamp 0
transform 1 0 6130 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2878_
timestamp 0
transform -1 0 5870 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2879_
timestamp 0
transform -1 0 9010 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2880_
timestamp 0
transform -1 0 12010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2881_
timestamp 0
transform 1 0 11690 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2882_
timestamp 0
transform -1 0 9290 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2883_
timestamp 0
transform 1 0 9090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2884_
timestamp 0
transform -1 0 9410 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2885_
timestamp 0
transform -1 0 10590 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2886_
timestamp 0
transform 1 0 10550 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2887_
timestamp 0
transform -1 0 8970 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2888_
timestamp 0
transform -1 0 9250 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2889_
timestamp 0
transform 1 0 9530 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2890_
timestamp 0
transform -1 0 9890 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__2891_
timestamp 0
transform -1 0 9830 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2892_
timestamp 0
transform 1 0 9210 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2893_
timestamp 0
transform -1 0 9370 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2894_
timestamp 0
transform -1 0 11190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2895_
timestamp 0
transform 1 0 10870 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2896_
timestamp 0
transform -1 0 11150 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2897_
timestamp 0
transform -1 0 10870 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2898_
timestamp 0
transform 1 0 9490 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2899_
timestamp 0
transform -1 0 9790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2900_
timestamp 0
transform 1 0 10470 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2901_
timestamp 0
transform -1 0 10490 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2902_
timestamp 0
transform 1 0 10670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2903_
timestamp 0
transform -1 0 10790 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2904_
timestamp 0
transform -1 0 9950 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2905_
timestamp 0
transform -1 0 9450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2906_
timestamp 0
transform -1 0 8610 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2907_
timestamp 0
transform -1 0 9170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2908_
timestamp 0
transform -1 0 10510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2909_
timestamp 0
transform 1 0 11870 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2910_
timestamp 0
transform 1 0 10950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2911_
timestamp 0
transform 1 0 11810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2912_
timestamp 0
transform 1 0 12090 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__2913_
timestamp 0
transform 1 0 10690 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__2914_
timestamp 0
transform -1 0 7870 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2915_
timestamp 0
transform 1 0 11010 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2916_
timestamp 0
transform 1 0 11250 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__2917_
timestamp 0
transform 1 0 10750 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2918_
timestamp 0
transform -1 0 10910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2919_
timestamp 0
transform 1 0 8590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2920_
timestamp 0
transform 1 0 11290 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2921_
timestamp 0
transform 1 0 11810 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__2922_
timestamp 0
transform -1 0 11930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2923_
timestamp 0
transform 1 0 11390 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2924_
timestamp 0
transform 1 0 10310 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2925_
timestamp 0
transform 1 0 10070 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2926_
timestamp 0
transform 1 0 10210 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2927_
timestamp 0
transform -1 0 10050 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2928_
timestamp 0
transform -1 0 10310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__2929_
timestamp 0
transform -1 0 10430 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__2930_
timestamp 0
transform -1 0 11310 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2931_
timestamp 0
transform -1 0 11570 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__2932_
timestamp 0
transform 1 0 11530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__2933_
timestamp 0
transform 1 0 11490 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__2934_
timestamp 0
transform 1 0 11570 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__2935_
timestamp 0
transform 1 0 11650 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2936_
timestamp 0
transform 1 0 10590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__2937_
timestamp 0
transform -1 0 3590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__2938_
timestamp 0
transform -1 0 7810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2939_
timestamp 0
transform 1 0 6570 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2940_
timestamp 0
transform -1 0 6350 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2941_
timestamp 0
transform -1 0 6270 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2942_
timestamp 0
transform 1 0 5170 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2943_
timestamp 0
transform -1 0 7070 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__2944_
timestamp 0
transform 1 0 5450 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2945_
timestamp 0
transform -1 0 6850 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2946_
timestamp 0
transform 1 0 6450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__2947_
timestamp 0
transform 1 0 7930 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2948_
timestamp 0
transform 1 0 7670 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2949_
timestamp 0
transform 1 0 5770 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__2950_
timestamp 0
transform -1 0 6110 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2951_
timestamp 0
transform 1 0 6870 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2952_
timestamp 0
transform 1 0 6590 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2953_
timestamp 0
transform 1 0 5750 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2954_
timestamp 0
transform -1 0 6050 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__2955_
timestamp 0
transform 1 0 7130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2956_
timestamp 0
transform 1 0 6610 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__2957_
timestamp 0
transform -1 0 8230 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__2958_
timestamp 0
transform 1 0 6610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__2959_
timestamp 0
transform 1 0 6350 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2960_
timestamp 0
transform -1 0 7230 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2961_
timestamp 0
transform 1 0 6610 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2962_
timestamp 0
transform -1 0 6390 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__2963_
timestamp 0
transform -1 0 6690 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2964_
timestamp 0
transform 1 0 4750 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2965_
timestamp 0
transform 1 0 5810 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2966_
timestamp 0
transform -1 0 6710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__2967_
timestamp 0
transform -1 0 5130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2968_
timestamp 0
transform -1 0 5390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2969_
timestamp 0
transform 1 0 4470 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2970_
timestamp 0
transform 1 0 4830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2971_
timestamp 0
transform 1 0 4710 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2972_
timestamp 0
transform -1 0 6150 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2973_
timestamp 0
transform -1 0 6410 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2974_
timestamp 0
transform -1 0 6410 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2975_
timestamp 0
transform 1 0 5870 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2976_
timestamp 0
transform -1 0 4790 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2977_
timestamp 0
transform -1 0 5050 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2978_
timestamp 0
transform 1 0 5310 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__2979_
timestamp 0
transform 1 0 5590 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__2980_
timestamp 0
transform -1 0 7470 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2981_
timestamp 0
transform -1 0 6430 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2982_
timestamp 0
transform -1 0 6710 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__2983_
timestamp 0
transform 1 0 7230 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2984_
timestamp 0
transform 1 0 6630 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__2985_
timestamp 0
transform -1 0 6970 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2986_
timestamp 0
transform 1 0 6670 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2987_
timestamp 0
transform 1 0 6110 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2988_
timestamp 0
transform -1 0 6390 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__2989_
timestamp 0
transform -1 0 7970 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2990_
timestamp 0
transform 1 0 7090 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__2991_
timestamp 0
transform -1 0 6950 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2992_
timestamp 0
transform -1 0 5250 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__2993_
timestamp 0
transform -1 0 6110 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2994_
timestamp 0
transform 1 0 5570 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2995_
timestamp 0
transform 1 0 6650 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2996_
timestamp 0
transform 1 0 6370 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__2997_
timestamp 0
transform 1 0 6090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2998_
timestamp 0
transform -1 0 5830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__2999_
timestamp 0
transform 1 0 6490 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3000_
timestamp 0
transform -1 0 5830 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__3001_
timestamp 0
transform 1 0 5050 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3002_
timestamp 0
transform -1 0 5550 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__3003_
timestamp 0
transform -1 0 5910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3004_
timestamp 0
transform -1 0 5330 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3005_
timestamp 0
transform -1 0 5590 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3006_
timestamp 0
transform -1 0 7490 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3007_
timestamp 0
transform 1 0 6910 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3008_
timestamp 0
transform 1 0 8710 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3009_
timestamp 0
transform 1 0 8170 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3010_
timestamp 0
transform 1 0 7190 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3011_
timestamp 0
transform -1 0 7290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3012_
timestamp 0
transform -1 0 7170 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3013_
timestamp 0
transform -1 0 7910 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3014_
timestamp 0
transform 1 0 7110 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3015_
timestamp 0
transform -1 0 7390 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3016_
timestamp 0
transform -1 0 6150 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3017_
timestamp 0
transform -1 0 6950 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3018_
timestamp 0
transform -1 0 6630 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3019_
timestamp 0
transform -1 0 6890 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3020_
timestamp 0
transform 1 0 5530 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__3021_
timestamp 0
transform 1 0 5970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3022_
timestamp 0
transform 1 0 5770 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__3023_
timestamp 0
transform -1 0 6850 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3024_
timestamp 0
transform -1 0 6770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3025_
timestamp 0
transform 1 0 6050 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__3026_
timestamp 0
transform 1 0 5470 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__3027_
timestamp 0
transform -1 0 5570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3028_
timestamp 0
transform 1 0 6050 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3029_
timestamp 0
transform 1 0 6810 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3030_
timestamp 0
transform 1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__3031_
timestamp 0
transform 1 0 4490 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3032_
timestamp 0
transform -1 0 5270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3033_
timestamp 0
transform 1 0 5530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3034_
timestamp 0
transform -1 0 3470 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3035_
timestamp 0
transform -1 0 4030 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3036_
timestamp 0
transform -1 0 3530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3037_
timestamp 0
transform -1 0 3410 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3038_
timestamp 0
transform 1 0 3630 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3039_
timestamp 0
transform -1 0 3130 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3040_
timestamp 0
transform 1 0 3010 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3041_
timestamp 0
transform 1 0 3250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3042_
timestamp 0
transform -1 0 3810 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3043_
timestamp 0
transform -1 0 3910 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3044_
timestamp 0
transform -1 0 3670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3045_
timestamp 0
transform 1 0 4470 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3046_
timestamp 0
transform 1 0 4190 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3047_
timestamp 0
transform -1 0 3150 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3048_
timestamp 0
transform 1 0 3190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3049_
timestamp 0
transform -1 0 2890 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3050_
timestamp 0
transform 1 0 2930 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3051_
timestamp 0
transform 1 0 2670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3052_
timestamp 0
transform 1 0 2570 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3053_
timestamp 0
transform 1 0 3330 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3054_
timestamp 0
transform -1 0 3610 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3055_
timestamp 0
transform 1 0 3430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3056_
timestamp 0
transform -1 0 3690 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3057_
timestamp 0
transform 1 0 3890 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3058_
timestamp 0
transform 1 0 4070 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3059_
timestamp 0
transform 1 0 4350 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3060_
timestamp 0
transform 1 0 4190 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3061_
timestamp 0
transform 1 0 3670 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3062_
timestamp 0
transform -1 0 3910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3063_
timestamp 0
transform -1 0 5150 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__3064_
timestamp 0
transform 1 0 5010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__3065_
timestamp 0
transform -1 0 4750 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3066_
timestamp 0
transform 1 0 4650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3067_
timestamp 0
transform -1 0 3750 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3068_
timestamp 0
transform -1 0 3490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3069_
timestamp 0
transform 1 0 3690 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3070_
timestamp 0
transform -1 0 4590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__3071_
timestamp 0
transform 1 0 4310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__3072_
timestamp 0
transform -1 0 4250 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3073_
timestamp 0
transform -1 0 4510 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3074_
timestamp 0
transform 1 0 5790 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3075_
timestamp 0
transform 1 0 5510 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3076_
timestamp 0
transform 1 0 3750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3077_
timestamp 0
transform 1 0 4070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3078_
timestamp 0
transform 1 0 4130 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3079_
timestamp 0
transform -1 0 4210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3080_
timestamp 0
transform 1 0 6350 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3081_
timestamp 0
transform -1 0 7010 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3082_
timestamp 0
transform 1 0 6710 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3083_
timestamp 0
transform -1 0 3890 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3084_
timestamp 0
transform 1 0 3590 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3085_
timestamp 0
transform 1 0 3210 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3086_
timestamp 0
transform -1 0 2930 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3087_
timestamp 0
transform 1 0 4410 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3088_
timestamp 0
transform -1 0 5010 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3089_
timestamp 0
transform 1 0 3490 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3090_
timestamp 0
transform -1 0 3770 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3091_
timestamp 0
transform -1 0 6310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3092_
timestamp 0
transform 1 0 5530 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3093_
timestamp 0
transform 1 0 5790 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3094_
timestamp 0
transform 1 0 5510 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3095_
timestamp 0
transform -1 0 4710 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3096_
timestamp 0
transform 1 0 4410 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3097_
timestamp 0
transform -1 0 4170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3098_
timestamp 0
transform 1 0 3870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3099_
timestamp 0
transform -1 0 3930 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3100_
timestamp 0
transform -1 0 3750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3101_
timestamp 0
transform 1 0 4970 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3102_
timestamp 0
transform -1 0 5270 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3103_
timestamp 0
transform -1 0 4650 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3104_
timestamp 0
transform -1 0 4930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3105_
timestamp 0
transform 1 0 5710 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3106_
timestamp 0
transform -1 0 6010 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3107_
timestamp 0
transform -1 0 4110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3108_
timestamp 0
transform 1 0 3810 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3109_
timestamp 0
transform 1 0 6290 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3110_
timestamp 0
transform 1 0 3970 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3111_
timestamp 0
transform 1 0 5830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3112_
timestamp 0
transform -1 0 5250 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3113_
timestamp 0
transform -1 0 4710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3114_
timestamp 0
transform 1 0 4410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3115_
timestamp 0
transform 1 0 4930 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3116_
timestamp 0
transform 1 0 3870 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3117_
timestamp 0
transform 1 0 4490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3118_
timestamp 0
transform -1 0 4790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3119_
timestamp 0
transform 1 0 4970 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3120_
timestamp 0
transform 1 0 4670 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3121_
timestamp 0
transform 1 0 5270 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3122_
timestamp 0
transform 1 0 5550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3123_
timestamp 0
transform 1 0 5530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3124_
timestamp 0
transform -1 0 5830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3125_
timestamp 0
transform -1 0 4190 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3126_
timestamp 0
transform 1 0 3890 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3127_
timestamp 0
transform 1 0 6550 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3128_
timestamp 0
transform 1 0 6110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3129_
timestamp 0
transform 1 0 5510 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3130_
timestamp 0
transform -1 0 3430 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3131_
timestamp 0
transform -1 0 3670 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3132_
timestamp 0
transform 1 0 4770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3133_
timestamp 0
transform 1 0 4010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3134_
timestamp 0
transform 1 0 5190 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3135_
timestamp 0
transform 1 0 4890 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3136_
timestamp 0
transform 1 0 5790 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3137_
timestamp 0
transform 1 0 5510 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3138_
timestamp 0
transform 1 0 5790 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3139_
timestamp 0
transform 1 0 5510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3140_
timestamp 0
transform -1 0 5710 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3141_
timestamp 0
transform -1 0 5970 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3142_
timestamp 0
transform -1 0 4310 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3143_
timestamp 0
transform -1 0 4570 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3144_
timestamp 0
transform 1 0 11650 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__3145_
timestamp 0
transform 1 0 11890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__3146_
timestamp 0
transform -1 0 11950 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__3147_
timestamp 0
transform 1 0 9570 0 1 790
box -6 -8 26 268
use FILL  FILL_7__3148_
timestamp 0
transform -1 0 11950 0 1 790
box -6 -8 26 268
use FILL  FILL_7__3149_
timestamp 0
transform -1 0 11570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3150_
timestamp 0
transform -1 0 11850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3151_
timestamp 0
transform -1 0 10790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3152_
timestamp 0
transform 1 0 9430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3153_
timestamp 0
transform -1 0 9730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3154_
timestamp 0
transform -1 0 10250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3155_
timestamp 0
transform -1 0 10370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3156_
timestamp 0
transform -1 0 9010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__3157_
timestamp 0
transform -1 0 9050 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__3158_
timestamp 0
transform -1 0 8770 0 1 2870
box -6 -8 26 268
use FILL  FILL_7__3159_
timestamp 0
transform -1 0 8750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__3160_
timestamp 0
transform 1 0 10590 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3161_
timestamp 0
transform 1 0 10310 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3162_
timestamp 0
transform -1 0 9850 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3163_
timestamp 0
transform 1 0 9570 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3164_
timestamp 0
transform -1 0 9050 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3165_
timestamp 0
transform -1 0 7270 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3166_
timestamp 0
transform 1 0 7670 0 1 1310
box -6 -8 26 268
use FILL  FILL_7__3167_
timestamp 0
transform 1 0 7530 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3168_
timestamp 0
transform 1 0 7690 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3169_
timestamp 0
transform -1 0 8770 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3170_
timestamp 0
transform -1 0 8490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3171_
timestamp 0
transform -1 0 9210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3172_
timestamp 0
transform -1 0 8210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3173_
timestamp 0
transform 1 0 8470 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3174_
timestamp 0
transform 1 0 7950 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3175_
timestamp 0
transform -1 0 7930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3176_
timestamp 0
transform -1 0 7650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3177_
timestamp 0
transform -1 0 11930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__3178_
timestamp 0
transform -1 0 11870 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3179_
timestamp 0
transform 1 0 12130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3180_
timestamp 0
transform 1 0 12190 0 1 790
box -6 -8 26 268
use FILL  FILL_7__3181_
timestamp 0
transform 1 0 12170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__3182_
timestamp 0
transform -1 0 11390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3183_
timestamp 0
transform 1 0 11650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3184_
timestamp 0
transform 1 0 11930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3185_
timestamp 0
transform 1 0 11950 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3186_
timestamp 0
transform 1 0 12130 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3187_
timestamp 0
transform 1 0 9990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7__3188_
timestamp 0
transform 1 0 10870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3189_
timestamp 0
transform -1 0 11130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_7__3190_
timestamp 0
transform 1 0 11170 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3191_
timestamp 0
transform 1 0 11110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3192_
timestamp 0
transform -1 0 10830 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3193_
timestamp 0
transform 1 0 10250 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3194_
timestamp 0
transform 1 0 10870 0 1 2350
box -6 -8 26 268
use FILL  FILL_7__3195_
timestamp 0
transform -1 0 10610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3196_
timestamp 0
transform 1 0 10510 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3197_
timestamp 0
transform -1 0 7370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3198_
timestamp 0
transform -1 0 4730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3199_
timestamp 0
transform 1 0 2890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7__3200_
timestamp 0
transform 1 0 4870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__3201_
timestamp 0
transform 1 0 4590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__3202_
timestamp 0
transform 1 0 1650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7__3203_
timestamp 0
transform 1 0 1610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3204_
timestamp 0
transform 1 0 1570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__3205_
timestamp 0
transform 1 0 1130 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__3206_
timestamp 0
transform 1 0 1550 0 1 3390
box -6 -8 26 268
use FILL  FILL_7__3207_
timestamp 0
transform -1 0 1690 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__3208_
timestamp 0
transform -1 0 1030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__3209_
timestamp 0
transform -1 0 730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__3210_
timestamp 0
transform -1 0 4390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__3211_
timestamp 0
transform 1 0 4330 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__3212_
timestamp 0
transform 1 0 1290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7__3213_
timestamp 0
transform 1 0 1190 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__3214_
timestamp 0
transform -1 0 2470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3215_
timestamp 0
transform 1 0 1890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3216_
timestamp 0
transform 1 0 5830 0 1 270
box -6 -8 26 268
use FILL  FILL_7__3217_
timestamp 0
transform -1 0 6130 0 1 270
box -6 -8 26 268
use FILL  FILL_7__3218_
timestamp 0
transform 1 0 6170 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3219_
timestamp 0
transform -1 0 6450 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3220_
timestamp 0
transform 1 0 3790 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3221_
timestamp 0
transform -1 0 4070 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3222_
timestamp 0
transform -1 0 3670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3223_
timestamp 0
transform 1 0 3390 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__3224_
timestamp 0
transform -1 0 3370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3225_
timestamp 0
transform 1 0 5510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__3226_
timestamp 0
transform 1 0 5230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__3227_
timestamp 0
transform -1 0 4350 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3228_
timestamp 0
transform -1 0 4550 0 1 270
box -6 -8 26 268
use FILL  FILL_7__3229_
timestamp 0
transform 1 0 2790 0 1 1830
box -6 -8 26 268
use FILL  FILL_7__3230_
timestamp 0
transform -1 0 2830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7__3231_
timestamp 0
transform 1 0 6070 0 1 790
box -6 -8 26 268
use FILL  FILL_7__3232_
timestamp 0
transform 1 0 6050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7__3364_
timestamp 0
transform 1 0 5330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3365_
timestamp 0
transform 1 0 4530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3366_
timestamp 0
transform 1 0 5010 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__3367_
timestamp 0
transform -1 0 4810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3368_
timestamp 0
transform -1 0 5070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3369_
timestamp 0
transform -1 0 5630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3370_
timestamp 0
transform 1 0 2770 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3371_
timestamp 0
transform 1 0 2270 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3372_
timestamp 0
transform -1 0 2390 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3373_
timestamp 0
transform -1 0 4050 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3374_
timestamp 0
transform -1 0 2370 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3375_
timestamp 0
transform 1 0 2370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3376_
timestamp 0
transform -1 0 3030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3377_
timestamp 0
transform 1 0 2490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3378_
timestamp 0
transform -1 0 2350 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3379_
timestamp 0
transform -1 0 1510 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3380_
timestamp 0
transform 1 0 1290 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3381_
timestamp 0
transform -1 0 1550 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3382_
timestamp 0
transform -1 0 2010 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3383_
timestamp 0
transform -1 0 1570 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3384_
timestamp 0
transform 1 0 1830 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3385_
timestamp 0
transform 1 0 1530 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3386_
timestamp 0
transform -1 0 2110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3387_
timestamp 0
transform 1 0 2370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3388_
timestamp 0
transform -1 0 710 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3389_
timestamp 0
transform 1 0 2570 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3390_
timestamp 0
transform 1 0 3390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3391_
timestamp 0
transform 1 0 3110 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3392_
timestamp 0
transform -1 0 2950 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3393_
timestamp 0
transform 1 0 2350 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3394_
timestamp 0
transform 1 0 750 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3395_
timestamp 0
transform -1 0 710 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3396_
timestamp 0
transform -1 0 450 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3397_
timestamp 0
transform -1 0 470 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3398_
timestamp 0
transform -1 0 170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3399_
timestamp 0
transform 1 0 150 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3400_
timestamp 0
transform -1 0 950 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3401_
timestamp 0
transform -1 0 1530 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3402_
timestamp 0
transform 1 0 1510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3403_
timestamp 0
transform 1 0 1230 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3404_
timestamp 0
transform -1 0 170 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3405_
timestamp 0
transform -1 0 430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3406_
timestamp 0
transform -1 0 170 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3407_
timestamp 0
transform -1 0 450 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3408_
timestamp 0
transform -1 0 170 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3409_
timestamp 0
transform -1 0 170 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3410_
timestamp 0
transform 1 0 1490 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3411_
timestamp 0
transform 1 0 1210 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3412_
timestamp 0
transform -1 0 690 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3413_
timestamp 0
transform 1 0 430 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3414_
timestamp 0
transform 1 0 690 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7__3415_
timestamp 0
transform -1 0 1010 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3416_
timestamp 0
transform 1 0 690 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3417_
timestamp 0
transform -1 0 730 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3418_
timestamp 0
transform -1 0 430 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3419_
timestamp 0
transform -1 0 1250 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3420_
timestamp 0
transform 1 0 950 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3421_
timestamp 0
transform 1 0 1250 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3422_
timestamp 0
transform 1 0 970 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3423_
timestamp 0
transform 1 0 1270 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3424_
timestamp 0
transform -1 0 1290 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3425_
timestamp 0
transform -1 0 1010 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3426_
timestamp 0
transform 1 0 990 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7__3427_
timestamp 0
transform -1 0 1510 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3428_
timestamp 0
transform 1 0 1190 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3429_
timestamp 0
transform -1 0 970 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3430_
timestamp 0
transform 1 0 1490 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3431_
timestamp 0
transform 1 0 1210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3432_
timestamp 0
transform -1 0 1010 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3433_
timestamp 0
transform -1 0 170 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3434_
timestamp 0
transform -1 0 750 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3435_
timestamp 0
transform -1 0 1030 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3436_
timestamp 0
transform -1 0 970 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3437_
timestamp 0
transform 1 0 1790 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3438_
timestamp 0
transform 1 0 1250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3439_
timestamp 0
transform -1 0 1530 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3440_
timestamp 0
transform 1 0 1250 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3441_
timestamp 0
transform -1 0 690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3442_
timestamp 0
transform 1 0 1270 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3443_
timestamp 0
transform 1 0 1190 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3444_
timestamp 0
transform -1 0 2090 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3445_
timestamp 0
transform 1 0 1770 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3446_
timestamp 0
transform 1 0 2130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3447_
timestamp 0
transform 1 0 2030 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3448_
timestamp 0
transform -1 0 1830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3449_
timestamp 0
transform 1 0 1510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3450_
timestamp 0
transform -1 0 970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3451_
timestamp 0
transform 1 0 1230 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3452_
timestamp 0
transform 1 0 930 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3453_
timestamp 0
transform -1 0 2250 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3454_
timestamp 0
transform 1 0 3170 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3455_
timestamp 0
transform -1 0 2110 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3456_
timestamp 0
transform -1 0 1770 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3457_
timestamp 0
transform -1 0 2950 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3458_
timestamp 0
transform -1 0 1810 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3459_
timestamp 0
transform -1 0 1750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3460_
timestamp 0
transform 1 0 1790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3461_
timestamp 0
transform -1 0 2010 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3462_
timestamp 0
transform -1 0 1770 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3463_
timestamp 0
transform -1 0 1530 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3464_
timestamp 0
transform 1 0 1250 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3465_
timestamp 0
transform -1 0 1510 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3466_
timestamp 0
transform 1 0 2050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3467_
timestamp 0
transform 1 0 2050 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3468_
timestamp 0
transform 1 0 2810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3469_
timestamp 0
transform 1 0 2670 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3470_
timestamp 0
transform -1 0 2570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3471_
timestamp 0
transform 1 0 2390 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3472_
timestamp 0
transform -1 0 2290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3473_
timestamp 0
transform 1 0 1530 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3474_
timestamp 0
transform -1 0 1790 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3475_
timestamp 0
transform 1 0 1270 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3476_
timestamp 0
transform -1 0 1010 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3477_
timestamp 0
transform 1 0 430 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3478_
timestamp 0
transform -1 0 410 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3479_
timestamp 0
transform -1 0 170 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3480_
timestamp 0
transform -1 0 170 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3481_
timestamp 0
transform -1 0 170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3482_
timestamp 0
transform 1 0 690 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3483_
timestamp 0
transform -1 0 410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3484_
timestamp 0
transform 1 0 2030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3485_
timestamp 0
transform -1 0 2090 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3486_
timestamp 0
transform -1 0 1470 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3487_
timestamp 0
transform -1 0 1790 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3488_
timestamp 0
transform -1 0 1590 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3489_
timestamp 0
transform 1 0 1530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3490_
timestamp 0
transform 1 0 1210 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3491_
timestamp 0
transform -1 0 1290 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3492_
timestamp 0
transform 1 0 1190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3493_
timestamp 0
transform -1 0 1010 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3494_
timestamp 0
transform 1 0 930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3495_
timestamp 0
transform -1 0 690 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3496_
timestamp 0
transform 1 0 450 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3497_
timestamp 0
transform -1 0 410 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3498_
timestamp 0
transform 1 0 710 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3499_
timestamp 0
transform -1 0 770 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3500_
timestamp 0
transform 1 0 710 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3501_
timestamp 0
transform 1 0 950 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3502_
timestamp 0
transform -1 0 470 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3503_
timestamp 0
transform -1 0 450 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3504_
timestamp 0
transform -1 0 690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3505_
timestamp 0
transform -1 0 450 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3506_
timestamp 0
transform -1 0 170 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3507_
timestamp 0
transform -1 0 170 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3508_
timestamp 0
transform 1 0 690 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3509_
timestamp 0
transform -1 0 950 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3510_
timestamp 0
transform -1 0 450 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3511_
timestamp 0
transform -1 0 170 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3512_
timestamp 0
transform 1 0 650 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3513_
timestamp 0
transform -1 0 470 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3514_
timestamp 0
transform -1 0 410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3515_
timestamp 0
transform -1 0 170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3516_
timestamp 0
transform -1 0 170 0 1 10150
box -6 -8 26 268
use FILL  FILL_7__3517_
timestamp 0
transform 1 0 710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3518_
timestamp 0
transform 1 0 930 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3519_
timestamp 0
transform 1 0 2630 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3520_
timestamp 0
transform 1 0 2910 0 1 9110
box -6 -8 26 268
use FILL  FILL_7__3521_
timestamp 0
transform 1 0 3390 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3522_
timestamp 0
transform 1 0 3090 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3523_
timestamp 0
transform 1 0 2650 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3524_
timestamp 0
transform -1 0 1030 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3525_
timestamp 0
transform -1 0 170 0 1 10670
box -6 -8 26 268
use FILL  FILL_7__3526_
timestamp 0
transform -1 0 170 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3527_
timestamp 0
transform -1 0 670 0 1 11190
box -6 -8 26 268
use FILL  FILL_7__3528_
timestamp 0
transform -1 0 690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_7__3529_
timestamp 0
transform -1 0 170 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7__3530_
timestamp 0
transform -1 0 170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3531_
timestamp 0
transform 1 0 150 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3532_
timestamp 0
transform 1 0 390 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3533_
timestamp 0
transform -1 0 170 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3534_
timestamp 0
transform -1 0 690 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3535_
timestamp 0
transform -1 0 450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7__3536_
timestamp 0
transform -1 0 430 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3537_
timestamp 0
transform -1 0 1790 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3538_
timestamp 0
transform 1 0 2550 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3539_
timestamp 0
transform -1 0 2650 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3540_
timestamp 0
transform -1 0 2390 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3541_
timestamp 0
transform -1 0 2110 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3542_
timestamp 0
transform -1 0 2290 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3543_
timestamp 0
transform 1 0 1690 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3544_
timestamp 0
transform 1 0 2050 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3545_
timestamp 0
transform 1 0 1850 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3546_
timestamp 0
transform 1 0 1970 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7__3547_
timestamp 0
transform -1 0 2630 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3548_
timestamp 0
transform 1 0 2330 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7__3549_
timestamp 0
transform -1 0 2430 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3550_
timestamp 0
transform 1 0 2130 0 1 11710
box -6 -8 26 268
use FILL  FILL_7__3551_
timestamp 0
transform -1 0 2610 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3552_
timestamp 0
transform 1 0 2310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7__3553_
timestamp 0
transform -1 0 1850 0 1 8070
box -6 -8 26 268
use FILL  FILL_7__3554_
timestamp 0
transform 1 0 990 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3555_
timestamp 0
transform 1 0 390 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3556_
timestamp 0
transform 1 0 1250 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7__3557_
timestamp 0
transform -1 0 3150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3558_
timestamp 0
transform 1 0 2850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7__3559_
timestamp 0
transform -1 0 2610 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3560_
timestamp 0
transform 1 0 2310 0 1 9630
box -6 -8 26 268
use FILL  FILL_7__3561_
timestamp 0
transform -1 0 2030 0 1 7550
box -6 -8 26 268
use FILL  FILL_7__3562_
timestamp 0
transform -1 0 2850 0 1 8590
box -6 -8 26 268
use FILL  FILL_7__3563_
timestamp 0
transform 1 0 2250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7__3564_
timestamp 0
transform 1 0 2530 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3565_
timestamp 0
transform -1 0 1530 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3566_
timestamp 0
transform -1 0 1790 0 1 7030
box -6 -8 26 268
use FILL  FILL_7__3579_
timestamp 0
transform -1 0 5130 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3580_
timestamp 0
transform -1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7__3581_
timestamp 0
transform -1 0 3550 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3582_
timestamp 0
transform -1 0 3290 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3583_
timestamp 0
transform -1 0 5410 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__3584_
timestamp 0
transform 1 0 4590 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3585_
timestamp 0
transform 1 0 3010 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3586_
timestamp 0
transform -1 0 5930 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__3587_
timestamp 0
transform 1 0 150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3588_
timestamp 0
transform -1 0 170 0 1 3910
box -6 -8 26 268
use FILL  FILL_7__3589_
timestamp 0
transform -1 0 170 0 1 4950
box -6 -8 26 268
use FILL  FILL_7__3590_
timestamp 0
transform -1 0 170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7__3591_
timestamp 0
transform -1 0 450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3592_
timestamp 0
transform -1 0 170 0 1 4430
box -6 -8 26 268
use FILL  FILL_7__3593_
timestamp 0
transform -1 0 4870 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3594_
timestamp 0
transform 1 0 5910 0 -1 270
box -6 -8 26 268
use FILL  FILL_7__3595_
timestamp 0
transform 1 0 5650 0 -1 790
box -6 -8 26 268
use FILL  FILL_7__3596_
timestamp 0
transform -1 0 950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3597_
timestamp 0
transform -1 0 170 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__3598_
timestamp 0
transform -1 0 430 0 1 5990
box -6 -8 26 268
use FILL  FILL_7__3599_
timestamp 0
transform -1 0 170 0 1 6510
box -6 -8 26 268
use FILL  FILL_7__3600_
timestamp 0
transform -1 0 170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7__3601_
timestamp 0
transform -1 0 170 0 1 5470
box -6 -8 26 268
use FILL  FILL_7__3602_
timestamp 0
transform -1 0 1790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7__3603_
timestamp 0
transform 1 0 6950 0 -1 270
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert0
timestamp 0
transform 1 0 7970 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert1
timestamp 0
transform 1 0 9470 0 1 1830
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert2
timestamp 0
transform 1 0 8230 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert3
timestamp 0
transform 1 0 11090 0 1 1830
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert4
timestamp 0
transform 1 0 690 0 1 1830
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert5
timestamp 0
transform -1 0 12170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert6
timestamp 0
transform -1 0 9670 0 1 5470
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert7
timestamp 0
transform 1 0 7130 0 1 2350
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert8
timestamp 0
transform -1 0 950 0 1 5470
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert9
timestamp 0
transform 1 0 10210 0 1 3910
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert10
timestamp 0
transform -1 0 990 0 1 5990
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert11
timestamp 0
transform -1 0 6070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert12
timestamp 0
transform 1 0 11630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert13
timestamp 0
transform -1 0 6250 0 1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert14
timestamp 0
transform 1 0 6870 0 1 2350
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert15
timestamp 0
transform -1 0 3410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert16
timestamp 0
transform -1 0 4030 0 1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert17
timestamp 0
transform 1 0 7270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert18
timestamp 0
transform -1 0 7090 0 1 11190
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert19
timestamp 0
transform 1 0 5410 0 1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert20
timestamp 0
transform 1 0 8650 0 1 11190
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert21
timestamp 0
transform -1 0 8570 0 -1 7550
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert22
timestamp 0
transform -1 0 1530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert23
timestamp 0
transform 1 0 3510 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert24
timestamp 0
transform -1 0 4410 0 1 5470
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert25
timestamp 0
transform 1 0 8250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert26
timestamp 0
transform 1 0 5190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert27
timestamp 0
transform -1 0 1330 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert39
timestamp 0
transform 1 0 6410 0 1 4950
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert40
timestamp 0
transform 1 0 7770 0 1 3910
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert41
timestamp 0
transform -1 0 8910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert42
timestamp 0
transform -1 0 7050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert43
timestamp 0
transform -1 0 8950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert44
timestamp 0
transform -1 0 9070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert45
timestamp 0
transform 1 0 11130 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert46
timestamp 0
transform 1 0 9570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert47
timestamp 0
transform 1 0 9290 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert48
timestamp 0
transform 1 0 7030 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert49
timestamp 0
transform 1 0 7290 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert50
timestamp 0
transform -1 0 7670 0 1 9110
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert51
timestamp 0
transform 1 0 7630 0 1 10150
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert52
timestamp 0
transform 1 0 9030 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert53
timestamp 0
transform 1 0 10070 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert54
timestamp 0
transform 1 0 8910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert55
timestamp 0
transform 1 0 8770 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert56
timestamp 0
transform -1 0 2310 0 1 8590
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert57
timestamp 0
transform 1 0 2610 0 1 11190
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert58
timestamp 0
transform 1 0 2750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert59
timestamp 0
transform -1 0 2310 0 1 10670
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert60
timestamp 0
transform -1 0 10570 0 1 7550
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert61
timestamp 0
transform 1 0 10630 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert62
timestamp 0
transform 1 0 10590 0 1 8070
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert63
timestamp 0
transform -1 0 9250 0 1 7550
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert64
timestamp 0
transform -1 0 8690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert65
timestamp 0
transform 1 0 5290 0 1 270
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert66
timestamp 0
transform 1 0 5810 0 1 790
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert67
timestamp 0
transform -1 0 3110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert68
timestamp 0
transform 1 0 3230 0 1 270
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert69
timestamp 0
transform -1 0 6730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert70
timestamp 0
transform 1 0 8670 0 1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert71
timestamp 0
transform -1 0 9330 0 1 2870
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert72
timestamp 0
transform -1 0 6850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert73
timestamp 0
transform 1 0 9010 0 -1 7030
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert74
timestamp 0
transform 1 0 10870 0 1 7030
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert75
timestamp 0
transform 1 0 2650 0 1 1310
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert76
timestamp 0
transform -1 0 3150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert77
timestamp 0
transform 1 0 10530 0 1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert78
timestamp 0
transform 1 0 9390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert79
timestamp 0
transform -1 0 8430 0 1 7550
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert80
timestamp 0
transform 1 0 7230 0 1 5470
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert81
timestamp 0
transform 1 0 7690 0 -1 790
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert82
timestamp 0
transform -1 0 7670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert83
timestamp 0
transform -1 0 7450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert84
timestamp 0
transform 1 0 9510 0 1 8590
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert85
timestamp 0
transform -1 0 8990 0 1 8590
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert86
timestamp 0
transform -1 0 9590 0 1 2870
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert87
timestamp 0
transform 1 0 9490 0 1 4430
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert88
timestamp 0
transform -1 0 10830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert89
timestamp 0
transform 1 0 9470 0 1 3390
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert90
timestamp 0
transform 1 0 5450 0 -1 11190
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert91
timestamp 0
transform -1 0 4990 0 1 10670
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert92
timestamp 0
transform -1 0 4830 0 -1 9630
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert93
timestamp 0
transform 1 0 5250 0 1 10150
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert94
timestamp 0
transform -1 0 11410 0 1 9630
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert95
timestamp 0
transform -1 0 11450 0 -1 10150
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert96
timestamp 0
transform -1 0 10170 0 1 11710
box -6 -8 26 268
use FILL  FILL_7_BUFX2_insert97
timestamp 0
transform 1 0 11530 0 1 11710
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert28
timestamp 0
transform -1 0 6110 0 -1 11710
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert29
timestamp 0
transform -1 0 2290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert30
timestamp 0
transform 1 0 4630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert31
timestamp 0
transform -1 0 3330 0 1 2870
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert32
timestamp 0
transform 1 0 7230 0 -1 8070
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert33
timestamp 0
transform 1 0 5810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert34
timestamp 0
transform -1 0 2570 0 1 10670
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert35
timestamp 0
transform -1 0 5330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert36
timestamp 0
transform -1 0 2450 0 1 3910
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert37
timestamp 0
transform 1 0 7470 0 -1 12230
box -6 -8 26 268
use FILL  FILL_7_CLKBUF1_insert38
timestamp 0
transform -1 0 4450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__1688_
timestamp 0
transform -1 0 990 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1689_
timestamp 0
transform -1 0 450 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1690_
timestamp 0
transform -1 0 710 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1691_
timestamp 0
transform 1 0 170 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1692_
timestamp 0
transform -1 0 430 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1693_
timestamp 0
transform 1 0 670 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1694_
timestamp 0
transform -1 0 5670 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__1695_
timestamp 0
transform -1 0 450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1696_
timestamp 0
transform -1 0 450 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1697_
timestamp 0
transform -1 0 1570 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__1698_
timestamp 0
transform -1 0 3510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1699_
timestamp 0
transform 1 0 2950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1700_
timestamp 0
transform -1 0 3990 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__1701_
timestamp 0
transform -1 0 690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1702_
timestamp 0
transform -1 0 690 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1703_
timestamp 0
transform 1 0 3330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1704_
timestamp 0
transform -1 0 470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1705_
timestamp 0
transform 1 0 170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1706_
timestamp 0
transform -1 0 3950 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1707_
timestamp 0
transform -1 0 710 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1708_
timestamp 0
transform 1 0 710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1709_
timestamp 0
transform 1 0 4230 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1710_
timestamp 0
transform -1 0 5710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1711_
timestamp 0
transform 1 0 5250 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1712_
timestamp 0
transform 1 0 7390 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1713_
timestamp 0
transform -1 0 9770 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1714_
timestamp 0
transform -1 0 9970 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1715_
timestamp 0
transform -1 0 8650 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1716_
timestamp 0
transform 1 0 11410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1717_
timestamp 0
transform 1 0 11210 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1718_
timestamp 0
transform 1 0 12030 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1719_
timestamp 0
transform -1 0 8910 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1720_
timestamp 0
transform -1 0 10230 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1721_
timestamp 0
transform -1 0 10250 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1722_
timestamp 0
transform -1 0 10010 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1723_
timestamp 0
transform 1 0 10110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1724_
timestamp 0
transform 1 0 9330 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1725_
timestamp 0
transform 1 0 9170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1726_
timestamp 0
transform 1 0 10270 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1727_
timestamp 0
transform -1 0 8890 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1728_
timestamp 0
transform 1 0 11670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1729_
timestamp 0
transform 1 0 10270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1730_
timestamp 0
transform 1 0 8450 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1731_
timestamp 0
transform 1 0 8690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1732_
timestamp 0
transform -1 0 7890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1733_
timestamp 0
transform 1 0 9830 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1734_
timestamp 0
transform 1 0 7530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1735_
timestamp 0
transform 1 0 10970 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1736_
timestamp 0
transform -1 0 10770 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1737_
timestamp 0
transform -1 0 11030 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1738_
timestamp 0
transform -1 0 10410 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1739_
timestamp 0
transform -1 0 10410 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1740_
timestamp 0
transform 1 0 10630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1741_
timestamp 0
transform -1 0 8530 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1742_
timestamp 0
transform -1 0 8430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1743_
timestamp 0
transform -1 0 9990 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1744_
timestamp 0
transform 1 0 9870 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1745_
timestamp 0
transform -1 0 9570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1746_
timestamp 0
transform 1 0 11430 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1747_
timestamp 0
transform 1 0 10910 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1748_
timestamp 0
transform 1 0 7630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1749_
timestamp 0
transform 1 0 8050 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__1750_
timestamp 0
transform -1 0 8170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1751_
timestamp 0
transform 1 0 7570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1752_
timestamp 0
transform -1 0 8990 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1753_
timestamp 0
transform 1 0 9850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1754_
timestamp 0
transform -1 0 8390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1755_
timestamp 0
transform -1 0 8970 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__1756_
timestamp 0
transform -1 0 11310 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1757_
timestamp 0
transform 1 0 11170 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1758_
timestamp 0
transform -1 0 9230 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1759_
timestamp 0
transform -1 0 7470 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__1760_
timestamp 0
transform 1 0 8970 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__1761_
timestamp 0
transform -1 0 9690 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1762_
timestamp 0
transform 1 0 10710 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1763_
timestamp 0
transform -1 0 9150 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1764_
timestamp 0
transform 1 0 11410 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1765_
timestamp 0
transform 1 0 8230 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1766_
timestamp 0
transform 1 0 8610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1767_
timestamp 0
transform 1 0 9310 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__1768_
timestamp 0
transform 1 0 8170 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__1769_
timestamp 0
transform 1 0 8690 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__1770_
timestamp 0
transform 1 0 9130 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__1771_
timestamp 0
transform 1 0 9090 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__1772_
timestamp 0
transform 1 0 8810 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__1773_
timestamp 0
transform 1 0 10890 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1774_
timestamp 0
transform 1 0 10890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1775_
timestamp 0
transform 1 0 10130 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1776_
timestamp 0
transform -1 0 8130 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1777_
timestamp 0
transform 1 0 8170 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1778_
timestamp 0
transform -1 0 7650 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1779_
timestamp 0
transform 1 0 5790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1780_
timestamp 0
transform -1 0 4190 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1781_
timestamp 0
transform -1 0 10910 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1782_
timestamp 0
transform 1 0 8390 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1783_
timestamp 0
transform 1 0 10630 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1784_
timestamp 0
transform -1 0 10110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1785_
timestamp 0
transform -1 0 9870 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1786_
timestamp 0
transform 1 0 10290 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1787_
timestamp 0
transform -1 0 9230 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1788_
timestamp 0
transform -1 0 8650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1789_
timestamp 0
transform 1 0 10090 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1790_
timestamp 0
transform -1 0 10150 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1791_
timestamp 0
transform -1 0 10230 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1792_
timestamp 0
transform -1 0 9770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1793_
timestamp 0
transform -1 0 9510 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1794_
timestamp 0
transform 1 0 9230 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1795_
timestamp 0
transform -1 0 8430 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1796_
timestamp 0
transform -1 0 8370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1797_
timestamp 0
transform 1 0 7210 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1798_
timestamp 0
transform 1 0 7470 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1799_
timestamp 0
transform -1 0 9490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1800_
timestamp 0
transform 1 0 11370 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1801_
timestamp 0
transform 1 0 9390 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1802_
timestamp 0
transform -1 0 9050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1803_
timestamp 0
transform 1 0 10650 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1804_
timestamp 0
transform -1 0 8670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1805_
timestamp 0
transform -1 0 8770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1806_
timestamp 0
transform 1 0 7710 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1807_
timestamp 0
transform -1 0 8170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1808_
timestamp 0
transform -1 0 8490 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1809_
timestamp 0
transform 1 0 8710 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1810_
timestamp 0
transform 1 0 8110 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1811_
timestamp 0
transform -1 0 7850 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1812_
timestamp 0
transform -1 0 8490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1813_
timestamp 0
transform -1 0 8210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1814_
timestamp 0
transform -1 0 7950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1815_
timestamp 0
transform 1 0 7970 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1816_
timestamp 0
transform -1 0 3970 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1817_
timestamp 0
transform 1 0 1450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1818_
timestamp 0
transform -1 0 6270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1819_
timestamp 0
transform -1 0 1030 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1820_
timestamp 0
transform 1 0 470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1821_
timestamp 0
transform 1 0 990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1822_
timestamp 0
transform -1 0 450 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1823_
timestamp 0
transform 1 0 1810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1824_
timestamp 0
transform 1 0 1390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__1825_
timestamp 0
transform -1 0 1230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1826_
timestamp 0
transform -1 0 490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1827_
timestamp 0
transform 1 0 990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1828_
timestamp 0
transform -1 0 1590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1829_
timestamp 0
transform -1 0 730 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1830_
timestamp 0
transform -1 0 1530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1831_
timestamp 0
transform 1 0 2110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1832_
timestamp 0
transform -1 0 8110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1833_
timestamp 0
transform 1 0 9750 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1834_
timestamp 0
transform 1 0 9330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1835_
timestamp 0
transform -1 0 7850 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1836_
timestamp 0
transform -1 0 6510 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1837_
timestamp 0
transform -1 0 7850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1838_
timestamp 0
transform -1 0 7290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1839_
timestamp 0
transform -1 0 6270 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1840_
timestamp 0
transform 1 0 8650 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1841_
timestamp 0
transform -1 0 8270 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1842_
timestamp 0
transform -1 0 7030 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1843_
timestamp 0
transform -1 0 6750 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1844_
timestamp 0
transform 1 0 9170 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1845_
timestamp 0
transform 1 0 9710 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1846_
timestamp 0
transform -1 0 9310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1847_
timestamp 0
transform -1 0 8470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1848_
timestamp 0
transform 1 0 11310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1849_
timestamp 0
transform -1 0 11630 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1850_
timestamp 0
transform -1 0 11090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1851_
timestamp 0
transform 1 0 10450 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1852_
timestamp 0
transform -1 0 10510 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1853_
timestamp 0
transform -1 0 10530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__1854_
timestamp 0
transform -1 0 7510 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1855_
timestamp 0
transform 1 0 7490 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1856_
timestamp 0
transform 1 0 7770 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1857_
timestamp 0
transform -1 0 8910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__1858_
timestamp 0
transform -1 0 9450 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1859_
timestamp 0
transform -1 0 8910 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1860_
timestamp 0
transform 1 0 9170 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1861_
timestamp 0
transform 1 0 6910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1862_
timestamp 0
transform -1 0 8410 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__1863_
timestamp 0
transform 1 0 7770 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1864_
timestamp 0
transform -1 0 6410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1865_
timestamp 0
transform -1 0 7850 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__1866_
timestamp 0
transform -1 0 7310 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1867_
timestamp 0
transform -1 0 8090 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1868_
timestamp 0
transform 1 0 7810 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1869_
timestamp 0
transform -1 0 6110 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__1870_
timestamp 0
transform 1 0 9450 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1871_
timestamp 0
transform 1 0 8930 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1872_
timestamp 0
transform -1 0 8670 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1873_
timestamp 0
transform -1 0 7870 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1874_
timestamp 0
transform -1 0 7590 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1875_
timestamp 0
transform -1 0 8390 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1876_
timestamp 0
transform -1 0 7030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1877_
timestamp 0
transform -1 0 5870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__1878_
timestamp 0
transform 1 0 6750 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1879_
timestamp 0
transform -1 0 7550 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1880_
timestamp 0
transform 1 0 6070 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__1881_
timestamp 0
transform 1 0 6070 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__1882_
timestamp 0
transform -1 0 5030 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__1883_
timestamp 0
transform -1 0 7930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1884_
timestamp 0
transform -1 0 8170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1885_
timestamp 0
transform -1 0 8730 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__1886_
timestamp 0
transform 1 0 8570 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1887_
timestamp 0
transform -1 0 8550 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1888_
timestamp 0
transform 1 0 11690 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1889_
timestamp 0
transform -1 0 8550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1890_
timestamp 0
transform 1 0 9810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1891_
timestamp 0
transform 1 0 8970 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1892_
timestamp 0
transform -1 0 8690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1893_
timestamp 0
transform 1 0 12210 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1894_
timestamp 0
transform 1 0 12190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1895_
timestamp 0
transform 1 0 12210 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1896_
timestamp 0
transform -1 0 10830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1897_
timestamp 0
transform -1 0 9230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1898_
timestamp 0
transform 1 0 9110 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1899_
timestamp 0
transform 1 0 7550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1900_
timestamp 0
transform 1 0 9750 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1901_
timestamp 0
transform 1 0 8090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1902_
timestamp 0
transform -1 0 8310 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1903_
timestamp 0
transform 1 0 8030 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1904_
timestamp 0
transform 1 0 11950 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1905_
timestamp 0
transform 1 0 11710 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1906_
timestamp 0
transform -1 0 6590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1907_
timestamp 0
transform -1 0 7130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1908_
timestamp 0
transform -1 0 7050 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1909_
timestamp 0
transform -1 0 6810 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__1910_
timestamp 0
transform -1 0 6310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1911_
timestamp 0
transform 1 0 6890 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1912_
timestamp 0
transform 1 0 6350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__1913_
timestamp 0
transform 1 0 6290 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1914_
timestamp 0
transform 1 0 5790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1915_
timestamp 0
transform 1 0 5310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1916_
timestamp 0
transform 1 0 5310 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__1917_
timestamp 0
transform -1 0 3810 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__1918_
timestamp 0
transform 1 0 3690 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__1919_
timestamp 0
transform -1 0 3970 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__1920_
timestamp 0
transform -1 0 3690 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__1921_
timestamp 0
transform -1 0 1810 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__1922_
timestamp 0
transform 1 0 7610 0 1 270
box -6 -8 26 268
use FILL  FILL_8__1923_
timestamp 0
transform 1 0 7870 0 1 790
box -6 -8 26 268
use FILL  FILL_8__1924_
timestamp 0
transform -1 0 6470 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__1925_
timestamp 0
transform -1 0 4710 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1926_
timestamp 0
transform -1 0 4070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1927_
timestamp 0
transform 1 0 2110 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__1928_
timestamp 0
transform -1 0 3270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__1929_
timestamp 0
transform 1 0 4650 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__1930_
timestamp 0
transform 1 0 3210 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__1931_
timestamp 0
transform -1 0 2990 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__1932_
timestamp 0
transform -1 0 1590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1933_
timestamp 0
transform -1 0 8550 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1934_
timestamp 0
transform 1 0 3950 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__1935_
timestamp 0
transform -1 0 3970 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1936_
timestamp 0
transform -1 0 2650 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1937_
timestamp 0
transform -1 0 1310 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1938_
timestamp 0
transform -1 0 3670 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1939_
timestamp 0
transform -1 0 4230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1940_
timestamp 0
transform -1 0 3450 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1941_
timestamp 0
transform -1 0 3390 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1942_
timestamp 0
transform -1 0 1890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__1943_
timestamp 0
transform -1 0 3690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__1944_
timestamp 0
transform -1 0 3790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1945_
timestamp 0
transform -1 0 3050 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__1946_
timestamp 0
transform -1 0 1610 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__1947_
timestamp 0
transform -1 0 5030 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__1948_
timestamp 0
transform 1 0 5230 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__1949_
timestamp 0
transform 1 0 5290 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__1950_
timestamp 0
transform -1 0 5030 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__1951_
timestamp 0
transform -1 0 2070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1952_
timestamp 0
transform 1 0 4190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__1953_
timestamp 0
transform 1 0 4130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__1954_
timestamp 0
transform 1 0 4270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1955_
timestamp 0
transform -1 0 1790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1956_
timestamp 0
transform -1 0 4410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__1957_
timestamp 0
transform 1 0 4990 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__1958_
timestamp 0
transform -1 0 5270 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__1959_
timestamp 0
transform -1 0 4250 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__1960_
timestamp 0
transform -1 0 2410 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1961_
timestamp 0
transform 1 0 4230 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1962_
timestamp 0
transform 1 0 3990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1963_
timestamp 0
transform 1 0 3770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1964_
timestamp 0
transform 1 0 2110 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1965_
timestamp 0
transform 1 0 6490 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__1966_
timestamp 0
transform 1 0 6430 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1967_
timestamp 0
transform 1 0 7270 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1968_
timestamp 0
transform 1 0 6730 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1969_
timestamp 0
transform -1 0 3390 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__1970_
timestamp 0
transform 1 0 2930 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1971_
timestamp 0
transform -1 0 4810 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1972_
timestamp 0
transform 1 0 3670 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1973_
timestamp 0
transform -1 0 3690 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__1974_
timestamp 0
transform -1 0 3190 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__1975_
timestamp 0
transform 1 0 3090 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__1976_
timestamp 0
transform -1 0 3190 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__1977_
timestamp 0
transform 1 0 4470 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__1978_
timestamp 0
transform 1 0 3170 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__1979_
timestamp 0
transform -1 0 2910 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__1980_
timestamp 0
transform -1 0 2430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1981_
timestamp 0
transform 1 0 6050 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__1982_
timestamp 0
transform 1 0 6170 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__1983_
timestamp 0
transform 1 0 6370 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__1984_
timestamp 0
transform 1 0 5370 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__1985_
timestamp 0
transform -1 0 4870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1986_
timestamp 0
transform 1 0 2650 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__1987_
timestamp 0
transform -1 0 7370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__1988_
timestamp 0
transform 1 0 7670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__1989_
timestamp 0
transform 1 0 7730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__1990_
timestamp 0
transform -1 0 7530 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1991_
timestamp 0
transform -1 0 7810 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__1992_
timestamp 0
transform 1 0 10550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__1993_
timestamp 0
transform 1 0 9670 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__1994_
timestamp 0
transform -1 0 6350 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__1995_
timestamp 0
transform 1 0 6730 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__1996_
timestamp 0
transform -1 0 6870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1997_
timestamp 0
transform 1 0 6570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__1998_
timestamp 0
transform 1 0 6570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__1999_
timestamp 0
transform 1 0 7630 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2000_
timestamp 0
transform 1 0 6550 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2001_
timestamp 0
transform 1 0 6790 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2002_
timestamp 0
transform 1 0 6750 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2003_
timestamp 0
transform 1 0 9630 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2004_
timestamp 0
transform 1 0 7570 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2005_
timestamp 0
transform -1 0 7370 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2006_
timestamp 0
transform 1 0 6850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2007_
timestamp 0
transform 1 0 6690 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2008_
timestamp 0
transform -1 0 6330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2009_
timestamp 0
transform 1 0 6930 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2010_
timestamp 0
transform -1 0 7150 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2011_
timestamp 0
transform 1 0 7390 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2012_
timestamp 0
transform -1 0 9530 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2013_
timestamp 0
transform 1 0 10670 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2014_
timestamp 0
transform -1 0 10930 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2015_
timestamp 0
transform -1 0 6370 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2016_
timestamp 0
transform -1 0 7410 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2017_
timestamp 0
transform -1 0 7190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2018_
timestamp 0
transform 1 0 7430 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2019_
timestamp 0
transform 1 0 9510 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2020_
timestamp 0
transform -1 0 10410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2021_
timestamp 0
transform -1 0 7450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2022_
timestamp 0
transform 1 0 7690 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2023_
timestamp 0
transform -1 0 7990 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2024_
timestamp 0
transform 1 0 6210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2025_
timestamp 0
transform -1 0 6090 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2026_
timestamp 0
transform 1 0 9790 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2027_
timestamp 0
transform 1 0 10330 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2028_
timestamp 0
transform -1 0 10330 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2029_
timestamp 0
transform -1 0 11210 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2030_
timestamp 0
transform 1 0 10830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2031_
timestamp 0
transform -1 0 11130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2032_
timestamp 0
transform 1 0 9050 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2033_
timestamp 0
transform 1 0 8510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2034_
timestamp 0
transform 1 0 8750 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2035_
timestamp 0
transform 1 0 8710 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2036_
timestamp 0
transform 1 0 11670 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2037_
timestamp 0
transform 1 0 11870 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2038_
timestamp 0
transform -1 0 7710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2039_
timestamp 0
transform -1 0 6790 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2040_
timestamp 0
transform 1 0 11050 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2041_
timestamp 0
transform 1 0 11130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2042_
timestamp 0
transform -1 0 10210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2043_
timestamp 0
transform -1 0 10590 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2044_
timestamp 0
transform -1 0 11110 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2045_
timestamp 0
transform -1 0 11450 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2046_
timestamp 0
transform 1 0 8930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2047_
timestamp 0
transform -1 0 9490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2048_
timestamp 0
transform 1 0 9290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2049_
timestamp 0
transform 1 0 9430 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2050_
timestamp 0
transform 1 0 9190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2051_
timestamp 0
transform 1 0 8890 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2052_
timestamp 0
transform 1 0 9170 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2053_
timestamp 0
transform -1 0 9730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2054_
timestamp 0
transform 1 0 9950 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2055_
timestamp 0
transform -1 0 6590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2056_
timestamp 0
transform -1 0 6170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2057_
timestamp 0
transform 1 0 10370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2058_
timestamp 0
transform -1 0 10110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2059_
timestamp 0
transform -1 0 10250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2060_
timestamp 0
transform -1 0 10010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2061_
timestamp 0
transform 1 0 10190 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2062_
timestamp 0
transform -1 0 9270 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2063_
timestamp 0
transform 1 0 8350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2064_
timestamp 0
transform -1 0 8030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2065_
timestamp 0
transform -1 0 8850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2066_
timestamp 0
transform 1 0 8830 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2067_
timestamp 0
transform -1 0 8090 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2068_
timestamp 0
transform -1 0 8370 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2069_
timestamp 0
transform 1 0 8090 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2070_
timestamp 0
transform -1 0 8390 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2071_
timestamp 0
transform -1 0 8670 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2072_
timestamp 0
transform 1 0 8890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2073_
timestamp 0
transform 1 0 9150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2074_
timestamp 0
transform 1 0 9370 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2075_
timestamp 0
transform -1 0 9670 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2076_
timestamp 0
transform 1 0 11330 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2077_
timestamp 0
transform -1 0 11390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2078_
timestamp 0
transform -1 0 11190 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2079_
timestamp 0
transform 1 0 11330 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2080_
timestamp 0
transform -1 0 11170 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2081_
timestamp 0
transform 1 0 11170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2082_
timestamp 0
transform 1 0 10430 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2083_
timestamp 0
transform 1 0 9690 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2084_
timestamp 0
transform 1 0 11710 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2085_
timestamp 0
transform 1 0 11130 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2086_
timestamp 0
transform 1 0 11630 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2087_
timestamp 0
transform 1 0 11650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2088_
timestamp 0
transform -1 0 12210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2089_
timestamp 0
transform 1 0 11930 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2090_
timestamp 0
transform 1 0 12110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2091_
timestamp 0
transform 1 0 10010 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2092_
timestamp 0
transform 1 0 10630 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2093_
timestamp 0
transform -1 0 11190 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2094_
timestamp 0
transform 1 0 11430 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2095_
timestamp 0
transform -1 0 11090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2096_
timestamp 0
transform 1 0 11610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2097_
timestamp 0
transform -1 0 11950 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2098_
timestamp 0
transform -1 0 12130 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2099_
timestamp 0
transform -1 0 11430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2100_
timestamp 0
transform 1 0 11390 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2101_
timestamp 0
transform -1 0 11350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2102_
timestamp 0
transform -1 0 11730 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2103_
timestamp 0
transform 1 0 12210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2104_
timestamp 0
transform 1 0 12210 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2105_
timestamp 0
transform -1 0 11670 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2106_
timestamp 0
transform -1 0 11650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2107_
timestamp 0
transform -1 0 12210 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2108_
timestamp 0
transform 1 0 8950 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2109_
timestamp 0
transform 1 0 12210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2110_
timestamp 0
transform -1 0 12230 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2111_
timestamp 0
transform -1 0 12230 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2112_
timestamp 0
transform -1 0 12130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2113_
timestamp 0
transform 1 0 11890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2114_
timestamp 0
transform 1 0 10670 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2115_
timestamp 0
transform -1 0 9410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2116_
timestamp 0
transform -1 0 10290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2117_
timestamp 0
transform -1 0 10890 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2118_
timestamp 0
transform -1 0 10850 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2119_
timestamp 0
transform 1 0 10750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2120_
timestamp 0
transform 1 0 10790 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2121_
timestamp 0
transform -1 0 10530 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2122_
timestamp 0
transform 1 0 10730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2123_
timestamp 0
transform -1 0 8230 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2124_
timestamp 0
transform -1 0 7930 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2125_
timestamp 0
transform -1 0 10290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2126_
timestamp 0
transform 1 0 10690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2127_
timestamp 0
transform -1 0 7110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2128_
timestamp 0
transform -1 0 9250 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2129_
timestamp 0
transform 1 0 7370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2130_
timestamp 0
transform -1 0 10990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2131_
timestamp 0
transform -1 0 8030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2132_
timestamp 0
transform 1 0 6810 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2133_
timestamp 0
transform -1 0 7110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2134_
timestamp 0
transform -1 0 7370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2135_
timestamp 0
transform -1 0 11250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2136_
timestamp 0
transform -1 0 11410 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2137_
timestamp 0
transform 1 0 11390 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2138_
timestamp 0
transform 1 0 11470 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2139_
timestamp 0
transform -1 0 11390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2140_
timestamp 0
transform -1 0 11110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2141_
timestamp 0
transform 1 0 10030 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2142_
timestamp 0
transform 1 0 10830 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2143_
timestamp 0
transform -1 0 10570 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2144_
timestamp 0
transform -1 0 11130 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2145_
timestamp 0
transform -1 0 5130 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2146_
timestamp 0
transform 1 0 9850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2147_
timestamp 0
transform 1 0 10410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2148_
timestamp 0
transform -1 0 6350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2149_
timestamp 0
transform 1 0 10130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2150_
timestamp 0
transform 1 0 8910 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2151_
timestamp 0
transform 1 0 7530 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2152_
timestamp 0
transform 1 0 8610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2153_
timestamp 0
transform 1 0 8870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2154_
timestamp 0
transform 1 0 9150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2155_
timestamp 0
transform -1 0 10230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2156_
timestamp 0
transform -1 0 11010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2157_
timestamp 0
transform 1 0 11250 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2158_
timestamp 0
transform -1 0 11830 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2159_
timestamp 0
transform -1 0 11950 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2160_
timestamp 0
transform -1 0 11490 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2161_
timestamp 0
transform 1 0 8230 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2162_
timestamp 0
transform 1 0 8990 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2163_
timestamp 0
transform -1 0 10090 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2164_
timestamp 0
transform 1 0 9850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2165_
timestamp 0
transform 1 0 11090 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2166_
timestamp 0
transform 1 0 10910 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2167_
timestamp 0
transform 1 0 9290 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2168_
timestamp 0
transform 1 0 10110 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2169_
timestamp 0
transform -1 0 8850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2170_
timestamp 0
transform -1 0 9270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2171_
timestamp 0
transform 1 0 10410 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2172_
timestamp 0
transform 1 0 9830 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2173_
timestamp 0
transform 1 0 9950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2174_
timestamp 0
transform -1 0 9590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2175_
timestamp 0
transform 1 0 9670 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2176_
timestamp 0
transform -1 0 9790 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2177_
timestamp 0
transform -1 0 9490 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2178_
timestamp 0
transform -1 0 11090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2179_
timestamp 0
transform 1 0 9570 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2180_
timestamp 0
transform 1 0 11930 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2181_
timestamp 0
transform 1 0 11910 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2182_
timestamp 0
transform 1 0 11990 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2183_
timestamp 0
transform -1 0 11370 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2184_
timestamp 0
transform 1 0 11110 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2185_
timestamp 0
transform -1 0 10350 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2186_
timestamp 0
transform 1 0 10290 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2187_
timestamp 0
transform -1 0 10690 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2188_
timestamp 0
transform 1 0 11650 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2189_
timestamp 0
transform 1 0 10030 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2190_
timestamp 0
transform 1 0 10590 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2191_
timestamp 0
transform 1 0 11210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2192_
timestamp 0
transform 1 0 11150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2193_
timestamp 0
transform -1 0 11090 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2194_
timestamp 0
transform -1 0 10650 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2195_
timestamp 0
transform -1 0 9530 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2196_
timestamp 0
transform -1 0 11170 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2197_
timestamp 0
transform 1 0 11430 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2198_
timestamp 0
transform -1 0 9970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2199_
timestamp 0
transform -1 0 10030 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2200_
timestamp 0
transform -1 0 5890 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2201_
timestamp 0
transform 1 0 6410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2202_
timestamp 0
transform 1 0 6150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2203_
timestamp 0
transform 1 0 6150 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2204_
timestamp 0
transform 1 0 6890 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2205_
timestamp 0
transform 1 0 7190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2206_
timestamp 0
transform 1 0 9530 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2207_
timestamp 0
transform -1 0 10030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2208_
timestamp 0
transform -1 0 9450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2209_
timestamp 0
transform 1 0 10490 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2210_
timestamp 0
transform 1 0 10490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2211_
timestamp 0
transform 1 0 11330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2212_
timestamp 0
transform -1 0 11690 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2213_
timestamp 0
transform -1 0 11730 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2214_
timestamp 0
transform 1 0 11690 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2215_
timestamp 0
transform 1 0 11790 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2216_
timestamp 0
transform 1 0 12170 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2217_
timestamp 0
transform 1 0 11450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2218_
timestamp 0
transform 1 0 9730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2219_
timestamp 0
transform -1 0 9970 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2220_
timestamp 0
transform -1 0 10010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2221_
timestamp 0
transform -1 0 11950 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2222_
timestamp 0
transform 1 0 11890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2223_
timestamp 0
transform -1 0 11930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2224_
timestamp 0
transform 1 0 11910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2225_
timestamp 0
transform 1 0 11010 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2226_
timestamp 0
transform 1 0 11970 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2227_
timestamp 0
transform 1 0 11690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2228_
timestamp 0
transform -1 0 11550 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2229_
timestamp 0
transform -1 0 10630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2230_
timestamp 0
transform -1 0 10350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2231_
timestamp 0
transform -1 0 8550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2232_
timestamp 0
transform 1 0 8790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2233_
timestamp 0
transform 1 0 9570 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2234_
timestamp 0
transform -1 0 9830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2235_
timestamp 0
transform -1 0 9950 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2236_
timestamp 0
transform 1 0 7250 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2237_
timestamp 0
transform -1 0 6730 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2238_
timestamp 0
transform -1 0 7010 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2239_
timestamp 0
transform -1 0 9030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2240_
timestamp 0
transform -1 0 8750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2241_
timestamp 0
transform -1 0 8390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2242_
timestamp 0
transform -1 0 7570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2243_
timestamp 0
transform 1 0 7830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2244_
timestamp 0
transform 1 0 8110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2245_
timestamp 0
transform -1 0 7810 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2246_
timestamp 0
transform 1 0 9190 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2247_
timestamp 0
transform -1 0 12190 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2248_
timestamp 0
transform 1 0 11390 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2249_
timestamp 0
transform -1 0 9550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2250_
timestamp 0
transform 1 0 11070 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2251_
timestamp 0
transform 1 0 10630 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2252_
timestamp 0
transform 1 0 11370 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2253_
timestamp 0
transform -1 0 11970 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2254_
timestamp 0
transform 1 0 12210 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2255_
timestamp 0
transform -1 0 10570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2256_
timestamp 0
transform -1 0 10850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2257_
timestamp 0
transform 1 0 11090 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2258_
timestamp 0
transform 1 0 12250 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2259_
timestamp 0
transform -1 0 11930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2260_
timestamp 0
transform 1 0 10110 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2261_
timestamp 0
transform 1 0 10370 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2262_
timestamp 0
transform -1 0 10890 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2263_
timestamp 0
transform 1 0 11370 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2264_
timestamp 0
transform 1 0 12190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2265_
timestamp 0
transform -1 0 11450 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2266_
timestamp 0
transform -1 0 10810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2267_
timestamp 0
transform 1 0 12030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2268_
timestamp 0
transform 1 0 12190 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2269_
timestamp 0
transform -1 0 11970 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2270_
timestamp 0
transform 1 0 11390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2271_
timestamp 0
transform -1 0 11690 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2272_
timestamp 0
transform 1 0 11950 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2273_
timestamp 0
transform -1 0 12210 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2274_
timestamp 0
transform 1 0 10130 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2275_
timestamp 0
transform -1 0 8290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2276_
timestamp 0
transform 1 0 8950 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2277_
timestamp 0
transform 1 0 9230 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2278_
timestamp 0
transform -1 0 9310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2279_
timestamp 0
transform 1 0 9110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2280_
timestamp 0
transform 1 0 10270 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2281_
timestamp 0
transform 1 0 12150 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2282_
timestamp 0
transform 1 0 12210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2283_
timestamp 0
transform -1 0 11090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2284_
timestamp 0
transform 1 0 12170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2285_
timestamp 0
transform 1 0 12170 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2286_
timestamp 0
transform -1 0 11950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2287_
timestamp 0
transform 1 0 11890 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2288_
timestamp 0
transform -1 0 11050 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2289_
timestamp 0
transform -1 0 10830 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2290_
timestamp 0
transform -1 0 11010 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2291_
timestamp 0
transform 1 0 11370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2292_
timestamp 0
transform 1 0 10510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2293_
timestamp 0
transform 1 0 10790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2294_
timestamp 0
transform 1 0 11110 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2295_
timestamp 0
transform 1 0 10990 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2296_
timestamp 0
transform 1 0 11250 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2297_
timestamp 0
transform 1 0 11910 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2298_
timestamp 0
transform -1 0 12010 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2299_
timestamp 0
transform -1 0 10570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2300_
timestamp 0
transform 1 0 10270 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2301_
timestamp 0
transform 1 0 11890 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2302_
timestamp 0
transform 1 0 11830 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2303_
timestamp 0
transform -1 0 11810 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2304_
timestamp 0
transform 1 0 11950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2305_
timestamp 0
transform 1 0 10830 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2306_
timestamp 0
transform -1 0 11690 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2307_
timestamp 0
transform 1 0 11390 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2308_
timestamp 0
transform 1 0 12170 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2309_
timestamp 0
transform -1 0 11730 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2310_
timestamp 0
transform -1 0 11670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2311_
timestamp 0
transform 1 0 11650 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2312_
timestamp 0
transform 1 0 11710 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2313_
timestamp 0
transform 1 0 11990 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2314_
timestamp 0
transform -1 0 11310 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2315_
timestamp 0
transform 1 0 12170 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2316_
timestamp 0
transform 1 0 11570 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2317_
timestamp 0
transform -1 0 12070 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2318_
timestamp 0
transform 1 0 11610 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2319_
timestamp 0
transform 1 0 11250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2320_
timestamp 0
transform 1 0 11670 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2321_
timestamp 0
transform 1 0 11530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2322_
timestamp 0
transform -1 0 11390 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2323_
timestamp 0
transform -1 0 11630 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2324_
timestamp 0
transform 1 0 11870 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2325_
timestamp 0
transform -1 0 12250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2326_
timestamp 0
transform 1 0 12170 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2327_
timestamp 0
transform 1 0 11530 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2328_
timestamp 0
transform 1 0 11110 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2329_
timestamp 0
transform 1 0 8630 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2330_
timestamp 0
transform -1 0 10310 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2331_
timestamp 0
transform -1 0 9750 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2332_
timestamp 0
transform -1 0 11970 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2333_
timestamp 0
transform -1 0 10850 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2334_
timestamp 0
transform 1 0 10570 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2335_
timestamp 0
transform 1 0 10550 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2336_
timestamp 0
transform 1 0 10730 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2337_
timestamp 0
transform -1 0 10850 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2338_
timestamp 0
transform -1 0 10770 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2339_
timestamp 0
transform -1 0 9690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2340_
timestamp 0
transform -1 0 9970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2341_
timestamp 0
transform 1 0 9670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2342_
timestamp 0
transform -1 0 10550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2343_
timestamp 0
transform -1 0 10490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2344_
timestamp 0
transform -1 0 10730 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2345_
timestamp 0
transform 1 0 11850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2346_
timestamp 0
transform 1 0 11590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2347_
timestamp 0
transform -1 0 8930 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2348_
timestamp 0
transform -1 0 10030 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2349_
timestamp 0
transform -1 0 11690 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2350_
timestamp 0
transform -1 0 11410 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2351_
timestamp 0
transform -1 0 10470 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2352_
timestamp 0
transform -1 0 10230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2353_
timestamp 0
transform -1 0 9530 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2354_
timestamp 0
transform 1 0 7930 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2355_
timestamp 0
transform -1 0 7010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2356_
timestamp 0
transform -1 0 6950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2357_
timestamp 0
transform -1 0 7610 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2358_
timestamp 0
transform -1 0 7190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2359_
timestamp 0
transform 1 0 7410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2360_
timestamp 0
transform -1 0 8090 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2361_
timestamp 0
transform -1 0 7150 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2362_
timestamp 0
transform 1 0 8870 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2363_
timestamp 0
transform -1 0 7550 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2364_
timestamp 0
transform 1 0 7290 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2365_
timestamp 0
transform 1 0 7010 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2366_
timestamp 0
transform 1 0 6490 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2367_
timestamp 0
transform -1 0 7330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2368_
timestamp 0
transform 1 0 6730 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2369_
timestamp 0
transform 1 0 7110 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2370_
timestamp 0
transform -1 0 7370 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2371_
timestamp 0
transform 1 0 7310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2372_
timestamp 0
transform -1 0 6890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2373_
timestamp 0
transform 1 0 6830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2374_
timestamp 0
transform 1 0 8330 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2375_
timestamp 0
transform 1 0 8390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2376_
timestamp 0
transform -1 0 6830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2377_
timestamp 0
transform 1 0 5530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2378_
timestamp 0
transform -1 0 3850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2379_
timestamp 0
transform -1 0 8110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2380_
timestamp 0
transform -1 0 5750 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2381_
timestamp 0
transform -1 0 6030 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2382_
timestamp 0
transform -1 0 5890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2383_
timestamp 0
transform 1 0 4810 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2384_
timestamp 0
transform 1 0 4730 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2385_
timestamp 0
transform 1 0 4970 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2386_
timestamp 0
transform 1 0 5250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2387_
timestamp 0
transform 1 0 1770 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2388_
timestamp 0
transform 1 0 1710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2389_
timestamp 0
transform 1 0 5290 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2390_
timestamp 0
transform 1 0 2570 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2391_
timestamp 0
transform -1 0 2370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2392_
timestamp 0
transform -1 0 2090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2393_
timestamp 0
transform -1 0 2650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2394_
timestamp 0
transform -1 0 3070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2395_
timestamp 0
transform 1 0 4470 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2396_
timestamp 0
transform 1 0 3110 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2397_
timestamp 0
transform -1 0 3190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2398_
timestamp 0
transform -1 0 2910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2399_
timestamp 0
transform 1 0 2010 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2400_
timestamp 0
transform -1 0 1450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2401_
timestamp 0
transform -1 0 2930 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2402_
timestamp 0
transform 1 0 2670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2403_
timestamp 0
transform -1 0 2310 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2404_
timestamp 0
transform -1 0 1750 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2405_
timestamp 0
transform -1 0 1610 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2406_
timestamp 0
transform 1 0 5990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2407_
timestamp 0
transform -1 0 4350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2408_
timestamp 0
transform -1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2409_
timestamp 0
transform -1 0 6530 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2410_
timestamp 0
transform -1 0 4310 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2411_
timestamp 0
transform -1 0 4070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2412_
timestamp 0
transform -1 0 1330 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2413_
timestamp 0
transform -1 0 4610 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2414_
timestamp 0
transform 1 0 3130 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2415_
timestamp 0
transform -1 0 2870 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2416_
timestamp 0
transform 1 0 1830 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2417_
timestamp 0
transform -1 0 2330 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2418_
timestamp 0
transform -1 0 2210 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2419_
timestamp 0
transform -1 0 3530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2420_
timestamp 0
transform 1 0 2950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2421_
timestamp 0
transform -1 0 2870 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2422_
timestamp 0
transform -1 0 2050 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2423_
timestamp 0
transform -1 0 3750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2424_
timestamp 0
transform -1 0 3590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2425_
timestamp 0
transform -1 0 3470 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2426_
timestamp 0
transform 1 0 3230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2427_
timestamp 0
transform 1 0 3390 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2428_
timestamp 0
transform -1 0 3470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2429_
timestamp 0
transform -1 0 5190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2430_
timestamp 0
transform -1 0 7890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2431_
timestamp 0
transform -1 0 5450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2432_
timestamp 0
transform -1 0 9570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2433_
timestamp 0
transform 1 0 11670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2434_
timestamp 0
transform 1 0 10850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2435_
timestamp 0
transform -1 0 7330 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2436_
timestamp 0
transform -1 0 7010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2437_
timestamp 0
transform -1 0 9690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2438_
timestamp 0
transform -1 0 9430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2439_
timestamp 0
transform -1 0 6210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2440_
timestamp 0
transform 1 0 7830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2441_
timestamp 0
transform -1 0 7670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2442_
timestamp 0
transform 1 0 10370 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2443_
timestamp 0
transform -1 0 7270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2444_
timestamp 0
transform -1 0 7270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2445_
timestamp 0
transform 1 0 5370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2446_
timestamp 0
transform 1 0 6490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2447_
timestamp 0
transform -1 0 4870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2448_
timestamp 0
transform -1 0 6470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2449_
timestamp 0
transform -1 0 7090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2450_
timestamp 0
transform 1 0 4230 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2451_
timestamp 0
transform -1 0 4110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2452_
timestamp 0
transform 1 0 4750 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2453_
timestamp 0
transform 1 0 8610 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2454_
timestamp 0
transform 1 0 4490 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2455_
timestamp 0
transform 1 0 4490 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2456_
timestamp 0
transform -1 0 4350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2457_
timestamp 0
transform -1 0 4610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2458_
timestamp 0
transform -1 0 4970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2459_
timestamp 0
transform 1 0 5110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2460_
timestamp 0
transform 1 0 4990 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2461_
timestamp 0
transform 1 0 5270 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2462_
timestamp 0
transform 1 0 5410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2463_
timestamp 0
transform 1 0 6350 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2464_
timestamp 0
transform -1 0 3290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2465_
timestamp 0
transform -1 0 3010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2466_
timestamp 0
transform -1 0 3010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2467_
timestamp 0
transform 1 0 2150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2468_
timestamp 0
transform -1 0 1710 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2469_
timestamp 0
transform 1 0 670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2470_
timestamp 0
transform -1 0 2770 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2471_
timestamp 0
transform -1 0 2790 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2472_
timestamp 0
transform -1 0 2490 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2473_
timestamp 0
transform 1 0 1990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2474_
timestamp 0
transform -1 0 1510 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2475_
timestamp 0
transform -1 0 450 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2476_
timestamp 0
transform -1 0 3870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2477_
timestamp 0
transform -1 0 5110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2478_
timestamp 0
transform 1 0 3970 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2479_
timestamp 0
transform -1 0 3610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2480_
timestamp 0
transform 1 0 1850 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2481_
timestamp 0
transform -1 0 3410 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2482_
timestamp 0
transform 1 0 3690 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2483_
timestamp 0
transform 1 0 3110 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2484_
timestamp 0
transform 1 0 2830 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2485_
timestamp 0
transform -1 0 450 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2486_
timestamp 0
transform -1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2487_
timestamp 0
transform 1 0 2450 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2488_
timestamp 0
transform -1 0 2450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2489_
timestamp 0
transform -1 0 1890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2490_
timestamp 0
transform -1 0 1450 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2491_
timestamp 0
transform -1 0 450 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2492_
timestamp 0
transform 1 0 4670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2493_
timestamp 0
transform 1 0 3670 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2494_
timestamp 0
transform 1 0 6250 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2495_
timestamp 0
transform 1 0 3910 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2496_
timestamp 0
transform 1 0 4210 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2497_
timestamp 0
transform -1 0 4130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2498_
timestamp 0
transform 1 0 3590 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2499_
timestamp 0
transform 1 0 3850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2500_
timestamp 0
transform -1 0 450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2501_
timestamp 0
transform -1 0 3450 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2502_
timestamp 0
transform -1 0 3090 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2503_
timestamp 0
transform -1 0 3570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__2504_
timestamp 0
transform -1 0 3330 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__2505_
timestamp 0
transform 1 0 2770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2506_
timestamp 0
transform -1 0 2590 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__2507_
timestamp 0
transform 1 0 710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2508_
timestamp 0
transform 1 0 3210 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2509_
timestamp 0
transform 1 0 2750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2510_
timestamp 0
transform -1 0 3310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2511_
timestamp 0
transform 1 0 3390 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__2512_
timestamp 0
transform 1 0 3230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2513_
timestamp 0
transform -1 0 2490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2514_
timestamp 0
transform 1 0 2190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2515_
timestamp 0
transform -1 0 2210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2516_
timestamp 0
transform -1 0 450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__2517_
timestamp 0
transform -1 0 2290 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2518_
timestamp 0
transform 1 0 5390 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2519_
timestamp 0
transform -1 0 5930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2520_
timestamp 0
transform -1 0 6030 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2521_
timestamp 0
transform 1 0 5730 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2522_
timestamp 0
transform -1 0 5730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2523_
timestamp 0
transform -1 0 5650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2524_
timestamp 0
transform -1 0 5590 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2525_
timestamp 0
transform -1 0 2810 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2526_
timestamp 0
transform 1 0 6210 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2527_
timestamp 0
transform 1 0 6610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2528_
timestamp 0
transform 1 0 6590 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2529_
timestamp 0
transform 1 0 6190 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2530_
timestamp 0
transform 1 0 5650 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2531_
timestamp 0
transform 1 0 3010 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2532_
timestamp 0
transform 1 0 4290 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2533_
timestamp 0
transform 1 0 5230 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2534_
timestamp 0
transform 1 0 4950 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2535_
timestamp 0
transform -1 0 4690 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2536_
timestamp 0
transform 1 0 3530 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2537_
timestamp 0
transform 1 0 2170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2538_
timestamp 0
transform 1 0 4570 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2539_
timestamp 0
transform 1 0 3950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2540_
timestamp 0
transform 1 0 4290 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2541_
timestamp 0
transform -1 0 4270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2542_
timestamp 0
transform -1 0 3790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2543_
timestamp 0
transform 1 0 3550 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2544_
timestamp 0
transform 1 0 4270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2545_
timestamp 0
transform 1 0 4530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2546_
timestamp 0
transform 1 0 4890 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2547_
timestamp 0
transform -1 0 4830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2548_
timestamp 0
transform -1 0 4550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2549_
timestamp 0
transform 1 0 4770 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2550_
timestamp 0
transform 1 0 4770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2551_
timestamp 0
transform 1 0 5290 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2552_
timestamp 0
transform 1 0 5530 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2553_
timestamp 0
transform 1 0 2430 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2554_
timestamp 0
transform 1 0 4570 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2555_
timestamp 0
transform -1 0 4750 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2556_
timestamp 0
transform -1 0 4990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2557_
timestamp 0
transform 1 0 4690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2558_
timestamp 0
transform 1 0 4770 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2559_
timestamp 0
transform 1 0 4490 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2560_
timestamp 0
transform 1 0 3990 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2561_
timestamp 0
transform 1 0 3690 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2562_
timestamp 0
transform 1 0 2310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2563_
timestamp 0
transform -1 0 4530 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2564_
timestamp 0
transform 1 0 4450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2565_
timestamp 0
transform -1 0 3930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2566_
timestamp 0
transform 1 0 2530 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2567_
timestamp 0
transform 1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2568_
timestamp 0
transform -1 0 5810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2569_
timestamp 0
transform -1 0 5950 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2570_
timestamp 0
transform 1 0 6030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2571_
timestamp 0
transform 1 0 6030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2572_
timestamp 0
transform 1 0 5890 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2573_
timestamp 0
transform 1 0 5810 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2574_
timestamp 0
transform 1 0 5790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2575_
timestamp 0
transform -1 0 4830 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2576_
timestamp 0
transform -1 0 4310 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2577_
timestamp 0
transform -1 0 4570 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2578_
timestamp 0
transform 1 0 7070 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2579_
timestamp 0
transform 1 0 7090 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2580_
timestamp 0
transform 1 0 8090 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2581_
timestamp 0
transform -1 0 8950 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2582_
timestamp 0
transform 1 0 6990 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2583_
timestamp 0
transform -1 0 6990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2584_
timestamp 0
transform 1 0 7410 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2585_
timestamp 0
transform 1 0 7450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2586_
timestamp 0
transform -1 0 8530 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2587_
timestamp 0
transform -1 0 6870 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2588_
timestamp 0
transform -1 0 5910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2589_
timestamp 0
transform 1 0 7530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2590_
timestamp 0
transform -1 0 6310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2591_
timestamp 0
transform 1 0 6550 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2592_
timestamp 0
transform -1 0 4530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2593_
timestamp 0
transform 1 0 5050 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2594_
timestamp 0
transform -1 0 8630 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2595_
timestamp 0
transform -1 0 5350 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2596_
timestamp 0
transform 1 0 5350 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2597_
timestamp 0
transform 1 0 5530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2598_
timestamp 0
transform -1 0 5270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2599_
timestamp 0
transform -1 0 5070 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2600_
timestamp 0
transform -1 0 5070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2601_
timestamp 0
transform -1 0 5330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2602_
timestamp 0
transform -1 0 8270 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2603_
timestamp 0
transform -1 0 6710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2604_
timestamp 0
transform -1 0 6470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2605_
timestamp 0
transform 1 0 6150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2606_
timestamp 0
transform -1 0 5650 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2607_
timestamp 0
transform 1 0 5810 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2608_
timestamp 0
transform 1 0 5630 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2609_
timestamp 0
transform -1 0 5610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2610_
timestamp 0
transform 1 0 4990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2611_
timestamp 0
transform -1 0 5250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2612_
timestamp 0
transform -1 0 5510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2613_
timestamp 0
transform -1 0 1330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2614_
timestamp 0
transform 1 0 2310 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2615_
timestamp 0
transform -1 0 2590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2616_
timestamp 0
transform -1 0 2570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2617_
timestamp 0
transform 1 0 1550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2618_
timestamp 0
transform 1 0 970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2619_
timestamp 0
transform -1 0 470 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2620_
timestamp 0
transform -1 0 710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2621_
timestamp 0
transform 1 0 1030 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2622_
timestamp 0
transform 1 0 470 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2623_
timestamp 0
transform 1 0 2850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2624_
timestamp 0
transform 1 0 2050 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2625_
timestamp 0
transform -1 0 2310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2626_
timestamp 0
transform -1 0 2030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2627_
timestamp 0
transform 1 0 170 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2628_
timestamp 0
transform 1 0 170 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2629_
timestamp 0
transform -1 0 430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2630_
timestamp 0
transform 1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2631_
timestamp 0
transform 1 0 5110 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2632_
timestamp 0
transform 1 0 2350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2633_
timestamp 0
transform -1 0 2650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2634_
timestamp 0
transform -1 0 190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2635_
timestamp 0
transform 1 0 170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2636_
timestamp 0
transform 1 0 710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2637_
timestamp 0
transform 1 0 1050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2638_
timestamp 0
transform 1 0 470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2639_
timestamp 0
transform -1 0 790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2640_
timestamp 0
transform -1 0 190 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2641_
timestamp 0
transform -1 0 190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2642_
timestamp 0
transform 1 0 1430 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2643_
timestamp 0
transform -1 0 1970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2644_
timestamp 0
transform 1 0 2370 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2645_
timestamp 0
transform -1 0 2110 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2646_
timestamp 0
transform -1 0 1310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2647_
timestamp 0
transform 1 0 170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2648_
timestamp 0
transform 1 0 670 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__2649_
timestamp 0
transform 1 0 170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2650_
timestamp 0
transform -1 0 3770 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2651_
timestamp 0
transform -1 0 3490 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2652_
timestamp 0
transform 1 0 710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2653_
timestamp 0
transform 1 0 430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2654_
timestamp 0
transform 1 0 1310 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2655_
timestamp 0
transform 1 0 750 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2656_
timestamp 0
transform -1 0 1030 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2657_
timestamp 0
transform 1 0 170 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2658_
timestamp 0
transform 1 0 170 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2659_
timestamp 0
transform -1 0 470 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2660_
timestamp 0
transform 1 0 410 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2661_
timestamp 0
transform -1 0 2730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__2662_
timestamp 0
transform -1 0 2670 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2663_
timestamp 0
transform -1 0 2090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2664_
timestamp 0
transform 1 0 990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2665_
timestamp 0
transform -1 0 950 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2666_
timestamp 0
transform -1 0 470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2667_
timestamp 0
transform -1 0 690 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2668_
timestamp 0
transform 1 0 1190 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2669_
timestamp 0
transform -1 0 2950 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2670_
timestamp 0
transform -1 0 3070 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2671_
timestamp 0
transform 1 0 1230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2672_
timestamp 0
transform -1 0 730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2673_
timestamp 0
transform -1 0 690 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2674_
timestamp 0
transform 1 0 950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2675_
timestamp 0
transform 1 0 930 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2676_
timestamp 0
transform -1 0 1230 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2677_
timestamp 0
transform 1 0 6570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__2678_
timestamp 0
transform -1 0 6490 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2679_
timestamp 0
transform 1 0 7110 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2680_
timestamp 0
transform -1 0 6910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2681_
timestamp 0
transform 1 0 7170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2682_
timestamp 0
transform -1 0 6890 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2683_
timestamp 0
transform -1 0 2010 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2684_
timestamp 0
transform -1 0 1830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__2685_
timestamp 0
transform 1 0 1750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2686_
timestamp 0
transform 1 0 1750 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2687_
timestamp 0
transform 1 0 1490 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2688_
timestamp 0
transform -1 0 930 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2689_
timestamp 0
transform -1 0 910 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2690_
timestamp 0
transform 1 0 7410 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2691_
timestamp 0
transform -1 0 7250 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2692_
timestamp 0
transform -1 0 5190 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2693_
timestamp 0
transform -1 0 3150 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2694_
timestamp 0
transform -1 0 1450 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2695_
timestamp 0
transform -1 0 1730 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2696_
timestamp 0
transform -1 0 1450 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2697_
timestamp 0
transform 1 0 2030 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2698_
timestamp 0
transform -1 0 670 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2699_
timestamp 0
transform 1 0 6430 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2700_
timestamp 0
transform -1 0 7150 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2701_
timestamp 0
transform 1 0 7730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2702_
timestamp 0
transform 1 0 7430 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2703_
timestamp 0
transform 1 0 7590 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2704_
timestamp 0
transform -1 0 6790 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2705_
timestamp 0
transform 1 0 1710 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2706_
timestamp 0
transform 1 0 1150 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2707_
timestamp 0
transform 1 0 2850 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2708_
timestamp 0
transform 1 0 2530 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2709_
timestamp 0
transform -1 0 1210 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2710_
timestamp 0
transform -1 0 990 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2711_
timestamp 0
transform -1 0 1270 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2712_
timestamp 0
transform 1 0 3010 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2713_
timestamp 0
transform -1 0 4410 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2714_
timestamp 0
transform -1 0 4830 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2715_
timestamp 0
transform 1 0 3670 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2716_
timestamp 0
transform -1 0 4430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2717_
timestamp 0
transform -1 0 5990 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__2718_
timestamp 0
transform -1 0 4230 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2719_
timestamp 0
transform 1 0 3830 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2720_
timestamp 0
transform -1 0 4130 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2721_
timestamp 0
transform -1 0 2290 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2722_
timestamp 0
transform 1 0 2410 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2723_
timestamp 0
transform 1 0 2710 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2724_
timestamp 0
transform -1 0 950 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2725_
timestamp 0
transform -1 0 5550 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2726_
timestamp 0
transform -1 0 6730 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2727_
timestamp 0
transform 1 0 3990 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2728_
timestamp 0
transform 1 0 3710 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2729_
timestamp 0
transform -1 0 3670 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2730_
timestamp 0
transform 1 0 3270 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2731_
timestamp 0
transform 1 0 2130 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2732_
timestamp 0
transform -1 0 2010 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2733_
timestamp 0
transform 1 0 1550 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2734_
timestamp 0
transform -1 0 1850 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2735_
timestamp 0
transform -1 0 4010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2736_
timestamp 0
transform -1 0 4150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2737_
timestamp 0
transform -1 0 4230 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2738_
timestamp 0
transform -1 0 3930 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2739_
timestamp 0
transform -1 0 3370 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2740_
timestamp 0
transform -1 0 3450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2741_
timestamp 0
transform -1 0 1210 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2742_
timestamp 0
transform 1 0 1510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2743_
timestamp 0
transform 1 0 1450 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2744_
timestamp 0
transform 1 0 1990 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2745_
timestamp 0
transform 1 0 650 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2746_
timestamp 0
transform 1 0 3710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2747_
timestamp 0
transform 1 0 4830 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__2748_
timestamp 0
transform 1 0 4490 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2749_
timestamp 0
transform -1 0 3650 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2750_
timestamp 0
transform -1 0 3090 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2751_
timestamp 0
transform 1 0 2930 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2752_
timestamp 0
transform 1 0 1230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2753_
timestamp 0
transform 1 0 730 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2754_
timestamp 0
transform -1 0 670 0 1 790
box -6 -8 26 268
use FILL  FILL_8__2755_
timestamp 0
transform -1 0 3190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2756_
timestamp 0
transform -1 0 2630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2757_
timestamp 0
transform 1 0 2870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2758_
timestamp 0
transform 1 0 2350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2759_
timestamp 0
transform -1 0 4430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2760_
timestamp 0
transform 1 0 3870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2761_
timestamp 0
transform 1 0 4210 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2762_
timestamp 0
transform -1 0 3950 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2763_
timestamp 0
transform -1 0 2190 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2764_
timestamp 0
transform -1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2765_
timestamp 0
transform -1 0 1830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2766_
timestamp 0
transform -1 0 2090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__2767_
timestamp 0
transform -1 0 1610 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__2768_
timestamp 0
transform 1 0 2270 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2769_
timestamp 0
transform 1 0 1710 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__2770_
timestamp 0
transform 1 0 6070 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2771_
timestamp 0
transform 1 0 6610 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2772_
timestamp 0
transform 1 0 5050 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__2773_
timestamp 0
transform 1 0 4250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2774_
timestamp 0
transform 1 0 2410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2775_
timestamp 0
transform 1 0 2650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2776_
timestamp 0
transform 1 0 3470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2777_
timestamp 0
transform -1 0 2950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2778_
timestamp 0
transform -1 0 3210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__2779_
timestamp 0
transform -1 0 7250 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2780_
timestamp 0
transform -1 0 7490 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__2781_
timestamp 0
transform 1 0 7970 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__2782_
timestamp 0
transform 1 0 7850 0 1 270
box -6 -8 26 268
use FILL  FILL_8__2783_
timestamp 0
transform 1 0 9790 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2784_
timestamp 0
transform 1 0 10930 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2785_
timestamp 0
transform 1 0 10310 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2786_
timestamp 0
transform 1 0 10030 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2787_
timestamp 0
transform 1 0 8490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2788_
timestamp 0
transform 1 0 8750 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2789_
timestamp 0
transform 1 0 8270 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2790_
timestamp 0
transform -1 0 8010 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2791_
timestamp 0
transform 1 0 6270 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2792_
timestamp 0
transform 1 0 9890 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2793_
timestamp 0
transform 1 0 10090 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2794_
timestamp 0
transform -1 0 10350 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2795_
timestamp 0
transform 1 0 8530 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2796_
timestamp 0
transform 1 0 8510 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2797_
timestamp 0
transform 1 0 10910 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2798_
timestamp 0
transform -1 0 10050 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2799_
timestamp 0
transform -1 0 8430 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2800_
timestamp 0
transform -1 0 7830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2801_
timestamp 0
transform 1 0 9770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2802_
timestamp 0
transform -1 0 10090 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2803_
timestamp 0
transform 1 0 8530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2804_
timestamp 0
transform -1 0 8430 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2805_
timestamp 0
transform -1 0 10170 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2806_
timestamp 0
transform 1 0 9850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2807_
timestamp 0
transform -1 0 8470 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2808_
timestamp 0
transform -1 0 6710 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2809_
timestamp 0
transform 1 0 8230 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2810_
timestamp 0
transform -1 0 7650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2811_
timestamp 0
transform 1 0 10130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2812_
timestamp 0
transform 1 0 9770 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2813_
timestamp 0
transform 1 0 8350 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2814_
timestamp 0
transform -1 0 8230 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2815_
timestamp 0
transform -1 0 8310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2816_
timestamp 0
transform 1 0 9570 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2817_
timestamp 0
transform -1 0 10430 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2818_
timestamp 0
transform 1 0 11250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2819_
timestamp 0
transform 1 0 10230 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2820_
timestamp 0
transform -1 0 10010 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2821_
timestamp 0
transform -1 0 9870 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2822_
timestamp 0
transform -1 0 7590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2823_
timestamp 0
transform -1 0 9590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2824_
timestamp 0
transform -1 0 9330 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2825_
timestamp 0
transform 1 0 8790 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2826_
timestamp 0
transform 1 0 8830 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2827_
timestamp 0
transform 1 0 9250 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2828_
timestamp 0
transform 1 0 10370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2829_
timestamp 0
transform -1 0 9310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2830_
timestamp 0
transform 1 0 9930 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2831_
timestamp 0
transform 1 0 9110 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2832_
timestamp 0
transform -1 0 9030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2833_
timestamp 0
transform -1 0 8790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2834_
timestamp 0
transform -1 0 8370 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2835_
timestamp 0
transform -1 0 9390 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2836_
timestamp 0
transform -1 0 8090 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2837_
timestamp 0
transform 1 0 8170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2838_
timestamp 0
transform 1 0 9410 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2839_
timestamp 0
transform 1 0 9670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2840_
timestamp 0
transform -1 0 9410 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2841_
timestamp 0
transform 1 0 8310 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2842_
timestamp 0
transform 1 0 11630 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2843_
timestamp 0
transform -1 0 11130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2844_
timestamp 0
transform 1 0 10850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2845_
timestamp 0
transform 1 0 10590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2846_
timestamp 0
transform -1 0 10230 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2847_
timestamp 0
transform 1 0 10430 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2848_
timestamp 0
transform -1 0 9710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2849_
timestamp 0
transform 1 0 11010 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__2850_
timestamp 0
transform 1 0 11170 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2851_
timestamp 0
transform 1 0 11410 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2852_
timestamp 0
transform 1 0 12110 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2853_
timestamp 0
transform 1 0 12170 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2854_
timestamp 0
transform 1 0 11850 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2855_
timestamp 0
transform 1 0 12130 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2856_
timestamp 0
transform -1 0 9170 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2857_
timestamp 0
transform 1 0 9670 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2858_
timestamp 0
transform -1 0 9970 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2859_
timestamp 0
transform 1 0 10910 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2860_
timestamp 0
transform 1 0 7790 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2861_
timestamp 0
transform 1 0 8470 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2862_
timestamp 0
transform -1 0 7850 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2863_
timestamp 0
transform 1 0 7550 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2864_
timestamp 0
transform 1 0 9790 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2865_
timestamp 0
transform 1 0 8950 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2866_
timestamp 0
transform -1 0 7050 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2867_
timestamp 0
transform -1 0 8890 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2868_
timestamp 0
transform -1 0 8610 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2869_
timestamp 0
transform -1 0 9050 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2870_
timestamp 0
transform 1 0 8690 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2871_
timestamp 0
transform 1 0 8650 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2872_
timestamp 0
transform 1 0 5590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2873_
timestamp 0
transform -1 0 5610 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2874_
timestamp 0
transform 1 0 5530 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2875_
timestamp 0
transform -1 0 5890 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2876_
timestamp 0
transform 1 0 5570 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2877_
timestamp 0
transform 1 0 6150 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2878_
timestamp 0
transform -1 0 5890 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2879_
timestamp 0
transform -1 0 9030 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2880_
timestamp 0
transform -1 0 12030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2881_
timestamp 0
transform 1 0 11710 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2882_
timestamp 0
transform -1 0 9310 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2883_
timestamp 0
transform 1 0 9110 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2884_
timestamp 0
transform -1 0 9430 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2885_
timestamp 0
transform -1 0 10610 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2886_
timestamp 0
transform 1 0 10570 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2887_
timestamp 0
transform -1 0 8990 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2888_
timestamp 0
transform -1 0 9270 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2889_
timestamp 0
transform 1 0 9550 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2890_
timestamp 0
transform -1 0 9910 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__2891_
timestamp 0
transform -1 0 9850 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2892_
timestamp 0
transform 1 0 9230 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2893_
timestamp 0
transform -1 0 9390 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2894_
timestamp 0
transform -1 0 11210 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2895_
timestamp 0
transform 1 0 10890 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2896_
timestamp 0
transform -1 0 11170 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2897_
timestamp 0
transform -1 0 10890 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2898_
timestamp 0
transform 1 0 9510 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2899_
timestamp 0
transform -1 0 9810 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2900_
timestamp 0
transform 1 0 10490 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2901_
timestamp 0
transform -1 0 10510 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2902_
timestamp 0
transform 1 0 10690 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2903_
timestamp 0
transform -1 0 10810 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2904_
timestamp 0
transform -1 0 9970 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2905_
timestamp 0
transform -1 0 9470 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2906_
timestamp 0
transform -1 0 8630 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2907_
timestamp 0
transform -1 0 9190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2908_
timestamp 0
transform -1 0 10530 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2909_
timestamp 0
transform 1 0 11890 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2910_
timestamp 0
transform 1 0 10970 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2911_
timestamp 0
transform 1 0 11830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2912_
timestamp 0
transform 1 0 12110 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__2913_
timestamp 0
transform 1 0 10710 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__2914_
timestamp 0
transform -1 0 7890 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2915_
timestamp 0
transform 1 0 11030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2916_
timestamp 0
transform 1 0 11270 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__2917_
timestamp 0
transform 1 0 10770 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2918_
timestamp 0
transform -1 0 10930 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2919_
timestamp 0
transform 1 0 8610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2920_
timestamp 0
transform 1 0 11310 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2921_
timestamp 0
transform 1 0 11830 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__2922_
timestamp 0
transform -1 0 11950 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2923_
timestamp 0
transform 1 0 11410 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2924_
timestamp 0
transform 1 0 10330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2925_
timestamp 0
transform 1 0 10090 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2926_
timestamp 0
transform 1 0 10230 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2927_
timestamp 0
transform -1 0 10070 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2928_
timestamp 0
transform -1 0 10330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__2929_
timestamp 0
transform -1 0 10450 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__2930_
timestamp 0
transform -1 0 11330 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2931_
timestamp 0
transform -1 0 11590 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__2932_
timestamp 0
transform 1 0 11550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__2933_
timestamp 0
transform 1 0 11510 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__2934_
timestamp 0
transform 1 0 11590 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__2935_
timestamp 0
transform 1 0 11670 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2936_
timestamp 0
transform 1 0 10610 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__2937_
timestamp 0
transform -1 0 3610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__2938_
timestamp 0
transform -1 0 7830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2939_
timestamp 0
transform 1 0 6590 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2940_
timestamp 0
transform -1 0 6370 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2941_
timestamp 0
transform -1 0 6290 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2942_
timestamp 0
transform 1 0 5190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2943_
timestamp 0
transform -1 0 7090 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__2944_
timestamp 0
transform 1 0 5470 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2945_
timestamp 0
transform -1 0 6870 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2946_
timestamp 0
transform 1 0 6470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__2947_
timestamp 0
transform 1 0 7950 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2948_
timestamp 0
transform 1 0 7690 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2949_
timestamp 0
transform 1 0 5790 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__2950_
timestamp 0
transform -1 0 6130 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2951_
timestamp 0
transform 1 0 6890 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2952_
timestamp 0
transform 1 0 6610 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2953_
timestamp 0
transform 1 0 5770 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2954_
timestamp 0
transform -1 0 6070 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__2955_
timestamp 0
transform 1 0 7150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2956_
timestamp 0
transform 1 0 6630 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__2957_
timestamp 0
transform -1 0 8250 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__2958_
timestamp 0
transform 1 0 6630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__2959_
timestamp 0
transform 1 0 6370 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2960_
timestamp 0
transform -1 0 7250 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2961_
timestamp 0
transform 1 0 6630 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2962_
timestamp 0
transform -1 0 6410 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__2963_
timestamp 0
transform -1 0 6710 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2964_
timestamp 0
transform 1 0 4770 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2965_
timestamp 0
transform 1 0 5830 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2966_
timestamp 0
transform -1 0 6730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__2967_
timestamp 0
transform -1 0 5150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2968_
timestamp 0
transform -1 0 5410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2969_
timestamp 0
transform 1 0 4490 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2970_
timestamp 0
transform 1 0 4850 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2971_
timestamp 0
transform 1 0 4730 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2972_
timestamp 0
transform -1 0 6170 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2973_
timestamp 0
transform -1 0 6430 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2974_
timestamp 0
transform -1 0 6430 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2975_
timestamp 0
transform 1 0 5890 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2976_
timestamp 0
transform -1 0 4810 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2977_
timestamp 0
transform -1 0 5070 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2978_
timestamp 0
transform 1 0 5330 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__2979_
timestamp 0
transform 1 0 5610 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__2980_
timestamp 0
transform -1 0 7490 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2981_
timestamp 0
transform -1 0 6450 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2982_
timestamp 0
transform -1 0 6730 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__2983_
timestamp 0
transform 1 0 7250 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2984_
timestamp 0
transform 1 0 6650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__2985_
timestamp 0
transform -1 0 6990 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2986_
timestamp 0
transform 1 0 6690 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2987_
timestamp 0
transform 1 0 6130 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2988_
timestamp 0
transform -1 0 6410 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__2989_
timestamp 0
transform -1 0 7990 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2990_
timestamp 0
transform 1 0 7110 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__2991_
timestamp 0
transform -1 0 6970 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2992_
timestamp 0
transform -1 0 5270 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__2993_
timestamp 0
transform -1 0 6130 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2994_
timestamp 0
transform 1 0 5590 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2995_
timestamp 0
transform 1 0 6670 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2996_
timestamp 0
transform 1 0 6390 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__2997_
timestamp 0
transform 1 0 6110 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2998_
timestamp 0
transform -1 0 5850 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__2999_
timestamp 0
transform 1 0 6510 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3000_
timestamp 0
transform -1 0 5850 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__3001_
timestamp 0
transform 1 0 5070 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3002_
timestamp 0
transform -1 0 5570 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__3003_
timestamp 0
transform -1 0 5930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3004_
timestamp 0
transform -1 0 5350 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3005_
timestamp 0
transform -1 0 5610 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3006_
timestamp 0
transform -1 0 7510 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3007_
timestamp 0
transform 1 0 6930 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3008_
timestamp 0
transform 1 0 8730 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3009_
timestamp 0
transform 1 0 8190 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3010_
timestamp 0
transform 1 0 7210 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3011_
timestamp 0
transform -1 0 7310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3012_
timestamp 0
transform -1 0 7190 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3013_
timestamp 0
transform -1 0 7930 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3014_
timestamp 0
transform 1 0 7130 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3015_
timestamp 0
transform -1 0 7410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3016_
timestamp 0
transform -1 0 6170 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3017_
timestamp 0
transform -1 0 6970 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3018_
timestamp 0
transform -1 0 6650 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3019_
timestamp 0
transform -1 0 6910 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3020_
timestamp 0
transform 1 0 5550 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__3021_
timestamp 0
transform 1 0 5990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3022_
timestamp 0
transform 1 0 5790 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__3023_
timestamp 0
transform -1 0 6870 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3024_
timestamp 0
transform -1 0 6790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3025_
timestamp 0
transform 1 0 6070 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__3026_
timestamp 0
transform 1 0 5490 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__3027_
timestamp 0
transform -1 0 5590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3028_
timestamp 0
transform 1 0 6070 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3029_
timestamp 0
transform 1 0 6830 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3030_
timestamp 0
transform 1 0 4970 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__3031_
timestamp 0
transform 1 0 4510 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3032_
timestamp 0
transform -1 0 5290 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3033_
timestamp 0
transform 1 0 5550 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3034_
timestamp 0
transform -1 0 3490 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3035_
timestamp 0
transform -1 0 4050 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3036_
timestamp 0
transform -1 0 3550 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3037_
timestamp 0
transform -1 0 3430 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3038_
timestamp 0
transform 1 0 3650 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3039_
timestamp 0
transform -1 0 3150 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3040_
timestamp 0
transform 1 0 3030 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3041_
timestamp 0
transform 1 0 3270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3042_
timestamp 0
transform -1 0 3830 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3043_
timestamp 0
transform -1 0 3930 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3044_
timestamp 0
transform -1 0 3690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3045_
timestamp 0
transform 1 0 4490 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3046_
timestamp 0
transform 1 0 4210 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3047_
timestamp 0
transform -1 0 3170 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3048_
timestamp 0
transform 1 0 3210 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3049_
timestamp 0
transform -1 0 2910 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3050_
timestamp 0
transform 1 0 2950 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3051_
timestamp 0
transform 1 0 2690 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3052_
timestamp 0
transform 1 0 2590 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3053_
timestamp 0
transform 1 0 3350 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3054_
timestamp 0
transform -1 0 3630 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3055_
timestamp 0
transform 1 0 3450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3056_
timestamp 0
transform -1 0 3710 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3057_
timestamp 0
transform 1 0 3910 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3058_
timestamp 0
transform 1 0 4090 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3059_
timestamp 0
transform 1 0 4370 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3060_
timestamp 0
transform 1 0 4210 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3061_
timestamp 0
transform 1 0 3690 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3062_
timestamp 0
transform -1 0 3930 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3063_
timestamp 0
transform -1 0 5170 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__3064_
timestamp 0
transform 1 0 5030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__3065_
timestamp 0
transform -1 0 4770 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3066_
timestamp 0
transform 1 0 4670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3067_
timestamp 0
transform -1 0 3770 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3068_
timestamp 0
transform -1 0 3510 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3069_
timestamp 0
transform 1 0 3710 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3070_
timestamp 0
transform -1 0 4610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__3071_
timestamp 0
transform 1 0 4330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__3072_
timestamp 0
transform -1 0 4270 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3073_
timestamp 0
transform -1 0 4530 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3074_
timestamp 0
transform 1 0 5810 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3075_
timestamp 0
transform 1 0 5530 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3076_
timestamp 0
transform 1 0 3770 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3077_
timestamp 0
transform 1 0 4090 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3078_
timestamp 0
transform 1 0 4150 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3079_
timestamp 0
transform -1 0 4230 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3080_
timestamp 0
transform 1 0 6370 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3081_
timestamp 0
transform -1 0 7030 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3082_
timestamp 0
transform 1 0 6730 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3083_
timestamp 0
transform -1 0 3910 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3084_
timestamp 0
transform 1 0 3610 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3085_
timestamp 0
transform 1 0 3230 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3086_
timestamp 0
transform -1 0 2950 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3087_
timestamp 0
transform 1 0 4430 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3088_
timestamp 0
transform -1 0 5030 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3089_
timestamp 0
transform 1 0 3510 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3090_
timestamp 0
transform -1 0 3790 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3091_
timestamp 0
transform -1 0 6330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3092_
timestamp 0
transform 1 0 5550 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3093_
timestamp 0
transform 1 0 5810 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3094_
timestamp 0
transform 1 0 5530 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3095_
timestamp 0
transform -1 0 4730 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3096_
timestamp 0
transform 1 0 4430 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3097_
timestamp 0
transform -1 0 4190 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3098_
timestamp 0
transform 1 0 3890 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3099_
timestamp 0
transform -1 0 3950 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3100_
timestamp 0
transform -1 0 3770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3101_
timestamp 0
transform 1 0 4990 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3102_
timestamp 0
transform -1 0 5290 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3103_
timestamp 0
transform -1 0 4670 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3104_
timestamp 0
transform -1 0 4950 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3105_
timestamp 0
transform 1 0 5730 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3106_
timestamp 0
transform -1 0 6030 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3107_
timestamp 0
transform -1 0 4130 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3108_
timestamp 0
transform 1 0 3830 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3109_
timestamp 0
transform 1 0 6310 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3110_
timestamp 0
transform 1 0 3990 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3111_
timestamp 0
transform 1 0 5850 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3112_
timestamp 0
transform -1 0 5270 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3113_
timestamp 0
transform -1 0 4730 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3114_
timestamp 0
transform 1 0 4430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3115_
timestamp 0
transform 1 0 4950 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3116_
timestamp 0
transform 1 0 3890 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3117_
timestamp 0
transform 1 0 4510 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3118_
timestamp 0
transform -1 0 4810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3119_
timestamp 0
transform 1 0 4990 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3120_
timestamp 0
transform 1 0 4690 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3121_
timestamp 0
transform 1 0 5290 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3122_
timestamp 0
transform 1 0 5570 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3123_
timestamp 0
transform 1 0 5550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3124_
timestamp 0
transform -1 0 5850 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3125_
timestamp 0
transform -1 0 4210 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3126_
timestamp 0
transform 1 0 3910 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3127_
timestamp 0
transform 1 0 6570 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3128_
timestamp 0
transform 1 0 6130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3129_
timestamp 0
transform 1 0 5530 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3130_
timestamp 0
transform -1 0 3450 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3131_
timestamp 0
transform -1 0 3690 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3132_
timestamp 0
transform 1 0 4790 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3133_
timestamp 0
transform 1 0 4030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3134_
timestamp 0
transform 1 0 5210 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3135_
timestamp 0
transform 1 0 4910 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3136_
timestamp 0
transform 1 0 5810 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3137_
timestamp 0
transform 1 0 5530 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3138_
timestamp 0
transform 1 0 5810 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3139_
timestamp 0
transform 1 0 5530 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3140_
timestamp 0
transform -1 0 5730 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3141_
timestamp 0
transform -1 0 5990 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3142_
timestamp 0
transform -1 0 4330 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3143_
timestamp 0
transform -1 0 4590 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3144_
timestamp 0
transform 1 0 11670 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__3145_
timestamp 0
transform 1 0 11910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__3146_
timestamp 0
transform -1 0 11970 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__3147_
timestamp 0
transform 1 0 9590 0 1 790
box -6 -8 26 268
use FILL  FILL_8__3148_
timestamp 0
transform -1 0 11970 0 1 790
box -6 -8 26 268
use FILL  FILL_8__3149_
timestamp 0
transform -1 0 11590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3150_
timestamp 0
transform -1 0 11870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3151_
timestamp 0
transform -1 0 10810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3152_
timestamp 0
transform 1 0 9450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3153_
timestamp 0
transform -1 0 9750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3154_
timestamp 0
transform -1 0 10270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3155_
timestamp 0
transform -1 0 10390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3156_
timestamp 0
transform -1 0 9030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__3157_
timestamp 0
transform -1 0 9070 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__3158_
timestamp 0
transform -1 0 8790 0 1 2870
box -6 -8 26 268
use FILL  FILL_8__3159_
timestamp 0
transform -1 0 8770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__3160_
timestamp 0
transform 1 0 10610 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3161_
timestamp 0
transform 1 0 10330 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3162_
timestamp 0
transform -1 0 9870 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3163_
timestamp 0
transform 1 0 9590 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3164_
timestamp 0
transform -1 0 9070 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3165_
timestamp 0
transform -1 0 7290 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3166_
timestamp 0
transform 1 0 7690 0 1 1310
box -6 -8 26 268
use FILL  FILL_8__3167_
timestamp 0
transform 1 0 7550 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3168_
timestamp 0
transform 1 0 7710 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3169_
timestamp 0
transform -1 0 8790 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3170_
timestamp 0
transform -1 0 8510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3171_
timestamp 0
transform -1 0 9230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3172_
timestamp 0
transform -1 0 8230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3173_
timestamp 0
transform 1 0 8490 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3174_
timestamp 0
transform 1 0 7970 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3175_
timestamp 0
transform -1 0 7950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3176_
timestamp 0
transform -1 0 7670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3177_
timestamp 0
transform -1 0 11950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__3178_
timestamp 0
transform -1 0 11890 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3179_
timestamp 0
transform 1 0 12150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3180_
timestamp 0
transform 1 0 12210 0 1 790
box -6 -8 26 268
use FILL  FILL_8__3181_
timestamp 0
transform 1 0 12190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__3182_
timestamp 0
transform -1 0 11410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3183_
timestamp 0
transform 1 0 11670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3184_
timestamp 0
transform 1 0 11950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3185_
timestamp 0
transform 1 0 11970 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3186_
timestamp 0
transform 1 0 12150 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3187_
timestamp 0
transform 1 0 10010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8__3188_
timestamp 0
transform 1 0 10890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3189_
timestamp 0
transform -1 0 11150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_8__3190_
timestamp 0
transform 1 0 11190 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3191_
timestamp 0
transform 1 0 11130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3192_
timestamp 0
transform -1 0 10850 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3193_
timestamp 0
transform 1 0 10270 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3194_
timestamp 0
transform 1 0 10890 0 1 2350
box -6 -8 26 268
use FILL  FILL_8__3195_
timestamp 0
transform -1 0 10630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3196_
timestamp 0
transform 1 0 10530 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3197_
timestamp 0
transform -1 0 7390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3198_
timestamp 0
transform -1 0 4750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3199_
timestamp 0
transform 1 0 2910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8__3200_
timestamp 0
transform 1 0 4890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__3201_
timestamp 0
transform 1 0 4610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__3202_
timestamp 0
transform 1 0 1670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8__3203_
timestamp 0
transform 1 0 1630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3204_
timestamp 0
transform 1 0 1590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__3205_
timestamp 0
transform 1 0 1150 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__3206_
timestamp 0
transform 1 0 1570 0 1 3390
box -6 -8 26 268
use FILL  FILL_8__3207_
timestamp 0
transform -1 0 1710 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__3208_
timestamp 0
transform -1 0 1050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__3209_
timestamp 0
transform -1 0 750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__3210_
timestamp 0
transform -1 0 4410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__3211_
timestamp 0
transform 1 0 4350 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__3212_
timestamp 0
transform 1 0 1310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8__3213_
timestamp 0
transform 1 0 1210 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__3214_
timestamp 0
transform -1 0 2490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3215_
timestamp 0
transform 1 0 1910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3216_
timestamp 0
transform 1 0 5850 0 1 270
box -6 -8 26 268
use FILL  FILL_8__3217_
timestamp 0
transform -1 0 6150 0 1 270
box -6 -8 26 268
use FILL  FILL_8__3218_
timestamp 0
transform 1 0 6190 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3219_
timestamp 0
transform -1 0 6470 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3220_
timestamp 0
transform 1 0 3810 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3221_
timestamp 0
transform -1 0 4090 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3222_
timestamp 0
transform -1 0 3690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3223_
timestamp 0
transform 1 0 3410 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__3224_
timestamp 0
transform -1 0 3390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3225_
timestamp 0
transform 1 0 5530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__3226_
timestamp 0
transform 1 0 5250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__3227_
timestamp 0
transform -1 0 4370 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3228_
timestamp 0
transform -1 0 4570 0 1 270
box -6 -8 26 268
use FILL  FILL_8__3229_
timestamp 0
transform 1 0 2810 0 1 1830
box -6 -8 26 268
use FILL  FILL_8__3230_
timestamp 0
transform -1 0 2850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8__3231_
timestamp 0
transform 1 0 6090 0 1 790
box -6 -8 26 268
use FILL  FILL_8__3232_
timestamp 0
transform 1 0 6070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8__3364_
timestamp 0
transform 1 0 5350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3365_
timestamp 0
transform 1 0 4550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3366_
timestamp 0
transform 1 0 5030 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__3367_
timestamp 0
transform -1 0 4830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3368_
timestamp 0
transform -1 0 5090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3369_
timestamp 0
transform -1 0 5650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3370_
timestamp 0
transform 1 0 2790 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3371_
timestamp 0
transform 1 0 2290 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3372_
timestamp 0
transform -1 0 2410 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3373_
timestamp 0
transform -1 0 4070 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3374_
timestamp 0
transform -1 0 2390 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3375_
timestamp 0
transform 1 0 2390 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3376_
timestamp 0
transform -1 0 3050 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3377_
timestamp 0
transform 1 0 2510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3378_
timestamp 0
transform -1 0 2370 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3379_
timestamp 0
transform -1 0 1530 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3380_
timestamp 0
transform 1 0 1310 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3381_
timestamp 0
transform -1 0 1570 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3382_
timestamp 0
transform -1 0 2030 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3383_
timestamp 0
transform -1 0 1590 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3384_
timestamp 0
transform 1 0 1850 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3385_
timestamp 0
transform 1 0 1550 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3386_
timestamp 0
transform -1 0 2130 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3387_
timestamp 0
transform 1 0 2390 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3388_
timestamp 0
transform -1 0 730 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3389_
timestamp 0
transform 1 0 2590 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3390_
timestamp 0
transform 1 0 3410 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3391_
timestamp 0
transform 1 0 3130 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3392_
timestamp 0
transform -1 0 2970 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3393_
timestamp 0
transform 1 0 2370 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3394_
timestamp 0
transform 1 0 770 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3395_
timestamp 0
transform -1 0 730 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3396_
timestamp 0
transform -1 0 470 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3397_
timestamp 0
transform -1 0 490 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3398_
timestamp 0
transform -1 0 190 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3399_
timestamp 0
transform 1 0 170 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3400_
timestamp 0
transform -1 0 970 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3401_
timestamp 0
transform -1 0 1550 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3402_
timestamp 0
transform 1 0 1530 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3403_
timestamp 0
transform 1 0 1250 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3404_
timestamp 0
transform -1 0 190 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3405_
timestamp 0
transform -1 0 450 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3406_
timestamp 0
transform -1 0 190 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3407_
timestamp 0
transform -1 0 470 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3408_
timestamp 0
transform -1 0 190 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3409_
timestamp 0
transform -1 0 190 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3410_
timestamp 0
transform 1 0 1510 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3411_
timestamp 0
transform 1 0 1230 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3412_
timestamp 0
transform -1 0 710 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3413_
timestamp 0
transform 1 0 450 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3414_
timestamp 0
transform 1 0 710 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8__3415_
timestamp 0
transform -1 0 1030 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3416_
timestamp 0
transform 1 0 710 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3417_
timestamp 0
transform -1 0 750 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3418_
timestamp 0
transform -1 0 450 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3419_
timestamp 0
transform -1 0 1270 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3420_
timestamp 0
transform 1 0 970 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3421_
timestamp 0
transform 1 0 1270 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3422_
timestamp 0
transform 1 0 990 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3423_
timestamp 0
transform 1 0 1290 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3424_
timestamp 0
transform -1 0 1310 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3425_
timestamp 0
transform -1 0 1030 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3426_
timestamp 0
transform 1 0 1010 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8__3427_
timestamp 0
transform -1 0 1530 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3428_
timestamp 0
transform 1 0 1210 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3429_
timestamp 0
transform -1 0 990 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3430_
timestamp 0
transform 1 0 1510 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3431_
timestamp 0
transform 1 0 1230 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3432_
timestamp 0
transform -1 0 1030 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3433_
timestamp 0
transform -1 0 190 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3434_
timestamp 0
transform -1 0 770 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3435_
timestamp 0
transform -1 0 1050 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3436_
timestamp 0
transform -1 0 990 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3437_
timestamp 0
transform 1 0 1810 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3438_
timestamp 0
transform 1 0 1270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3439_
timestamp 0
transform -1 0 1550 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3440_
timestamp 0
transform 1 0 1270 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3441_
timestamp 0
transform -1 0 710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3442_
timestamp 0
transform 1 0 1290 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3443_
timestamp 0
transform 1 0 1210 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3444_
timestamp 0
transform -1 0 2110 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3445_
timestamp 0
transform 1 0 1790 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3446_
timestamp 0
transform 1 0 2150 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3447_
timestamp 0
transform 1 0 2050 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3448_
timestamp 0
transform -1 0 1850 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3449_
timestamp 0
transform 1 0 1530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3450_
timestamp 0
transform -1 0 990 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3451_
timestamp 0
transform 1 0 1250 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3452_
timestamp 0
transform 1 0 950 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3453_
timestamp 0
transform -1 0 2270 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3454_
timestamp 0
transform 1 0 3190 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3455_
timestamp 0
transform -1 0 2130 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3456_
timestamp 0
transform -1 0 1790 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3457_
timestamp 0
transform -1 0 2970 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3458_
timestamp 0
transform -1 0 1830 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3459_
timestamp 0
transform -1 0 1770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3460_
timestamp 0
transform 1 0 1810 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3461_
timestamp 0
transform -1 0 2030 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3462_
timestamp 0
transform -1 0 1790 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3463_
timestamp 0
transform -1 0 1550 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3464_
timestamp 0
transform 1 0 1270 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3465_
timestamp 0
transform -1 0 1530 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3466_
timestamp 0
transform 1 0 2070 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3467_
timestamp 0
transform 1 0 2070 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3468_
timestamp 0
transform 1 0 2830 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3469_
timestamp 0
transform 1 0 2690 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3470_
timestamp 0
transform -1 0 2590 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3471_
timestamp 0
transform 1 0 2410 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3472_
timestamp 0
transform -1 0 2310 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3473_
timestamp 0
transform 1 0 1550 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3474_
timestamp 0
transform -1 0 1810 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3475_
timestamp 0
transform 1 0 1290 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3476_
timestamp 0
transform -1 0 1030 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3477_
timestamp 0
transform 1 0 450 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3478_
timestamp 0
transform -1 0 430 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3479_
timestamp 0
transform -1 0 190 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3480_
timestamp 0
transform -1 0 190 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3481_
timestamp 0
transform -1 0 190 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3482_
timestamp 0
transform 1 0 710 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3483_
timestamp 0
transform -1 0 430 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3484_
timestamp 0
transform 1 0 2050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3485_
timestamp 0
transform -1 0 2110 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3486_
timestamp 0
transform -1 0 1490 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3487_
timestamp 0
transform -1 0 1810 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3488_
timestamp 0
transform -1 0 1610 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3489_
timestamp 0
transform 1 0 1550 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3490_
timestamp 0
transform 1 0 1230 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3491_
timestamp 0
transform -1 0 1310 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3492_
timestamp 0
transform 1 0 1210 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3493_
timestamp 0
transform -1 0 1030 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3494_
timestamp 0
transform 1 0 950 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3495_
timestamp 0
transform -1 0 710 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3496_
timestamp 0
transform 1 0 470 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3497_
timestamp 0
transform -1 0 430 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3498_
timestamp 0
transform 1 0 730 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3499_
timestamp 0
transform -1 0 790 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3500_
timestamp 0
transform 1 0 730 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3501_
timestamp 0
transform 1 0 970 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3502_
timestamp 0
transform -1 0 490 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3503_
timestamp 0
transform -1 0 470 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3504_
timestamp 0
transform -1 0 710 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3505_
timestamp 0
transform -1 0 470 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3506_
timestamp 0
transform -1 0 190 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3507_
timestamp 0
transform -1 0 190 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3508_
timestamp 0
transform 1 0 710 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3509_
timestamp 0
transform -1 0 970 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3510_
timestamp 0
transform -1 0 470 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3511_
timestamp 0
transform -1 0 190 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3512_
timestamp 0
transform 1 0 670 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3513_
timestamp 0
transform -1 0 490 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3514_
timestamp 0
transform -1 0 430 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3515_
timestamp 0
transform -1 0 190 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3516_
timestamp 0
transform -1 0 190 0 1 10150
box -6 -8 26 268
use FILL  FILL_8__3517_
timestamp 0
transform 1 0 730 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3518_
timestamp 0
transform 1 0 950 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3519_
timestamp 0
transform 1 0 2650 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3520_
timestamp 0
transform 1 0 2930 0 1 9110
box -6 -8 26 268
use FILL  FILL_8__3521_
timestamp 0
transform 1 0 3410 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3522_
timestamp 0
transform 1 0 3110 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3523_
timestamp 0
transform 1 0 2670 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3524_
timestamp 0
transform -1 0 1050 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3525_
timestamp 0
transform -1 0 190 0 1 10670
box -6 -8 26 268
use FILL  FILL_8__3526_
timestamp 0
transform -1 0 190 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3527_
timestamp 0
transform -1 0 690 0 1 11190
box -6 -8 26 268
use FILL  FILL_8__3528_
timestamp 0
transform -1 0 710 0 -1 10670
box -6 -8 26 268
use FILL  FILL_8__3529_
timestamp 0
transform -1 0 190 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8__3530_
timestamp 0
transform -1 0 190 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3531_
timestamp 0
transform 1 0 170 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3532_
timestamp 0
transform 1 0 410 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3533_
timestamp 0
transform -1 0 190 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3534_
timestamp 0
transform -1 0 710 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3535_
timestamp 0
transform -1 0 470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8__3536_
timestamp 0
transform -1 0 450 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3537_
timestamp 0
transform -1 0 1810 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3538_
timestamp 0
transform 1 0 2570 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3539_
timestamp 0
transform -1 0 2670 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3540_
timestamp 0
transform -1 0 2410 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3541_
timestamp 0
transform -1 0 2130 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3542_
timestamp 0
transform -1 0 2310 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3543_
timestamp 0
transform 1 0 1710 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3544_
timestamp 0
transform 1 0 2070 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3545_
timestamp 0
transform 1 0 1870 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3546_
timestamp 0
transform 1 0 1990 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8__3547_
timestamp 0
transform -1 0 2650 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3548_
timestamp 0
transform 1 0 2350 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8__3549_
timestamp 0
transform -1 0 2450 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3550_
timestamp 0
transform 1 0 2150 0 1 11710
box -6 -8 26 268
use FILL  FILL_8__3551_
timestamp 0
transform -1 0 2630 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3552_
timestamp 0
transform 1 0 2330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8__3553_
timestamp 0
transform -1 0 1870 0 1 8070
box -6 -8 26 268
use FILL  FILL_8__3554_
timestamp 0
transform 1 0 1010 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3555_
timestamp 0
transform 1 0 410 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3556_
timestamp 0
transform 1 0 1270 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8__3557_
timestamp 0
transform -1 0 3170 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3558_
timestamp 0
transform 1 0 2870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8__3559_
timestamp 0
transform -1 0 2630 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3560_
timestamp 0
transform 1 0 2330 0 1 9630
box -6 -8 26 268
use FILL  FILL_8__3561_
timestamp 0
transform -1 0 2050 0 1 7550
box -6 -8 26 268
use FILL  FILL_8__3562_
timestamp 0
transform -1 0 2870 0 1 8590
box -6 -8 26 268
use FILL  FILL_8__3563_
timestamp 0
transform 1 0 2270 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8__3564_
timestamp 0
transform 1 0 2550 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3565_
timestamp 0
transform -1 0 1550 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3566_
timestamp 0
transform -1 0 1810 0 1 7030
box -6 -8 26 268
use FILL  FILL_8__3579_
timestamp 0
transform -1 0 5150 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3580_
timestamp 0
transform -1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8__3581_
timestamp 0
transform -1 0 3570 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3582_
timestamp 0
transform -1 0 3310 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3583_
timestamp 0
transform -1 0 5430 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__3584_
timestamp 0
transform 1 0 4610 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3585_
timestamp 0
transform 1 0 3030 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3586_
timestamp 0
transform -1 0 5950 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__3587_
timestamp 0
transform 1 0 170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3588_
timestamp 0
transform -1 0 190 0 1 3910
box -6 -8 26 268
use FILL  FILL_8__3589_
timestamp 0
transform -1 0 190 0 1 4950
box -6 -8 26 268
use FILL  FILL_8__3590_
timestamp 0
transform -1 0 190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8__3591_
timestamp 0
transform -1 0 470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3592_
timestamp 0
transform -1 0 190 0 1 4430
box -6 -8 26 268
use FILL  FILL_8__3593_
timestamp 0
transform -1 0 4890 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3594_
timestamp 0
transform 1 0 5930 0 -1 270
box -6 -8 26 268
use FILL  FILL_8__3595_
timestamp 0
transform 1 0 5670 0 -1 790
box -6 -8 26 268
use FILL  FILL_8__3596_
timestamp 0
transform -1 0 970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3597_
timestamp 0
transform -1 0 190 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__3598_
timestamp 0
transform -1 0 450 0 1 5990
box -6 -8 26 268
use FILL  FILL_8__3599_
timestamp 0
transform -1 0 190 0 1 6510
box -6 -8 26 268
use FILL  FILL_8__3600_
timestamp 0
transform -1 0 190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8__3601_
timestamp 0
transform -1 0 190 0 1 5470
box -6 -8 26 268
use FILL  FILL_8__3602_
timestamp 0
transform -1 0 1810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8__3603_
timestamp 0
transform 1 0 6970 0 -1 270
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert0
timestamp 0
transform 1 0 7990 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert1
timestamp 0
transform 1 0 9490 0 1 1830
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert2
timestamp 0
transform 1 0 8250 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert3
timestamp 0
transform 1 0 11110 0 1 1830
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert4
timestamp 0
transform 1 0 710 0 1 1830
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert5
timestamp 0
transform -1 0 12190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert6
timestamp 0
transform -1 0 9690 0 1 5470
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert7
timestamp 0
transform 1 0 7150 0 1 2350
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert8
timestamp 0
transform -1 0 970 0 1 5470
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert9
timestamp 0
transform 1 0 10230 0 1 3910
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert10
timestamp 0
transform -1 0 1010 0 1 5990
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert11
timestamp 0
transform -1 0 6090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert12
timestamp 0
transform 1 0 11650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert13
timestamp 0
transform -1 0 6270 0 1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert14
timestamp 0
transform 1 0 6890 0 1 2350
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert15
timestamp 0
transform -1 0 3430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert16
timestamp 0
transform -1 0 4050 0 1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert17
timestamp 0
transform 1 0 7290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert18
timestamp 0
transform -1 0 7110 0 1 11190
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert19
timestamp 0
transform 1 0 5430 0 1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert20
timestamp 0
transform 1 0 8670 0 1 11190
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert21
timestamp 0
transform -1 0 8590 0 -1 7550
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert22
timestamp 0
transform -1 0 1550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert23
timestamp 0
transform 1 0 3530 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert24
timestamp 0
transform -1 0 4430 0 1 5470
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert25
timestamp 0
transform 1 0 8270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert26
timestamp 0
transform 1 0 5210 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert27
timestamp 0
transform -1 0 1350 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert39
timestamp 0
transform 1 0 6430 0 1 4950
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert40
timestamp 0
transform 1 0 7790 0 1 3910
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert41
timestamp 0
transform -1 0 8930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert42
timestamp 0
transform -1 0 7070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert43
timestamp 0
transform -1 0 8970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert44
timestamp 0
transform -1 0 9090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert45
timestamp 0
transform 1 0 11150 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert46
timestamp 0
transform 1 0 9590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert47
timestamp 0
transform 1 0 9310 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert48
timestamp 0
transform 1 0 7050 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert49
timestamp 0
transform 1 0 7310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert50
timestamp 0
transform -1 0 7690 0 1 9110
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert51
timestamp 0
transform 1 0 7650 0 1 10150
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert52
timestamp 0
transform 1 0 9050 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert53
timestamp 0
transform 1 0 10090 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert54
timestamp 0
transform 1 0 8930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert55
timestamp 0
transform 1 0 8790 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert56
timestamp 0
transform -1 0 2330 0 1 8590
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert57
timestamp 0
transform 1 0 2630 0 1 11190
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert58
timestamp 0
transform 1 0 2770 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert59
timestamp 0
transform -1 0 2330 0 1 10670
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert60
timestamp 0
transform -1 0 10590 0 1 7550
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert61
timestamp 0
transform 1 0 10650 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert62
timestamp 0
transform 1 0 10610 0 1 8070
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert63
timestamp 0
transform -1 0 9270 0 1 7550
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert64
timestamp 0
transform -1 0 8710 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert65
timestamp 0
transform 1 0 5310 0 1 270
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert66
timestamp 0
transform 1 0 5830 0 1 790
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert67
timestamp 0
transform -1 0 3130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert68
timestamp 0
transform 1 0 3250 0 1 270
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert69
timestamp 0
transform -1 0 6750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert70
timestamp 0
transform 1 0 8690 0 1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert71
timestamp 0
transform -1 0 9350 0 1 2870
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert72
timestamp 0
transform -1 0 6870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert73
timestamp 0
transform 1 0 9030 0 -1 7030
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert74
timestamp 0
transform 1 0 10890 0 1 7030
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert75
timestamp 0
transform 1 0 2670 0 1 1310
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert76
timestamp 0
transform -1 0 3170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert77
timestamp 0
transform 1 0 10550 0 1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert78
timestamp 0
transform 1 0 9410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert79
timestamp 0
transform -1 0 8450 0 1 7550
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert80
timestamp 0
transform 1 0 7250 0 1 5470
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert81
timestamp 0
transform 1 0 7710 0 -1 790
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert82
timestamp 0
transform -1 0 7690 0 -1 8590
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert83
timestamp 0
transform -1 0 7470 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert84
timestamp 0
transform 1 0 9530 0 1 8590
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert85
timestamp 0
transform -1 0 9010 0 1 8590
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert86
timestamp 0
transform -1 0 9610 0 1 2870
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert87
timestamp 0
transform 1 0 9510 0 1 4430
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert88
timestamp 0
transform -1 0 10850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert89
timestamp 0
transform 1 0 9490 0 1 3390
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert90
timestamp 0
transform 1 0 5470 0 -1 11190
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert91
timestamp 0
transform -1 0 5010 0 1 10670
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert92
timestamp 0
transform -1 0 4850 0 -1 9630
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert93
timestamp 0
transform 1 0 5270 0 1 10150
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert94
timestamp 0
transform -1 0 11430 0 1 9630
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert95
timestamp 0
transform -1 0 11470 0 -1 10150
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert96
timestamp 0
transform -1 0 10190 0 1 11710
box -6 -8 26 268
use FILL  FILL_8_BUFX2_insert97
timestamp 0
transform 1 0 11550 0 1 11710
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert28
timestamp 0
transform -1 0 6130 0 -1 11710
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert29
timestamp 0
transform -1 0 2310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert30
timestamp 0
transform 1 0 4650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert31
timestamp 0
transform -1 0 3350 0 1 2870
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert32
timestamp 0
transform 1 0 7250 0 -1 8070
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert33
timestamp 0
transform 1 0 5830 0 -1 9110
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert34
timestamp 0
transform -1 0 2590 0 1 10670
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert35
timestamp 0
transform -1 0 5350 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert36
timestamp 0
transform -1 0 2470 0 1 3910
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert37
timestamp 0
transform 1 0 7490 0 -1 12230
box -6 -8 26 268
use FILL  FILL_8_CLKBUF1_insert38
timestamp 0
transform -1 0 4470 0 -1 9630
box -6 -8 26 268
use FILL  FILL_9__1693_
timestamp 0
transform 1 0 690 0 -1 270
box -6 -8 26 268
use FILL  FILL_9__1707_
timestamp 0
transform -1 0 730 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__1722_
timestamp 0
transform -1 0 10030 0 -1 270
box -6 -8 26 268
use FILL  FILL_9__1737_
timestamp 0
transform -1 0 11050 0 -1 790
box -6 -8 26 268
use FILL  FILL_9__1751_
timestamp 0
transform 1 0 7590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_9__1766_
timestamp 0
transform 1 0 8630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__1781_
timestamp 0
transform -1 0 10930 0 1 2870
box -6 -8 26 268
use FILL  FILL_9__1796_
timestamp 0
transform -1 0 8390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_9__1810_
timestamp 0
transform 1 0 8130 0 1 3390
box -6 -8 26 268
use FILL  FILL_9__1825_
timestamp 0
transform -1 0 1250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__1840_
timestamp 0
transform 1 0 8670 0 1 1830
box -6 -8 26 268
use FILL  FILL_9__1854_
timestamp 0
transform -1 0 7530 0 1 6510
box -6 -8 26 268
use FILL  FILL_9__1869_
timestamp 0
transform -1 0 6130 0 1 10150
box -6 -8 26 268
use FILL  FILL_9__1884_
timestamp 0
transform -1 0 8190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_9__1899_
timestamp 0
transform 1 0 7570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__1913_
timestamp 0
transform 1 0 6310 0 1 1310
box -6 -8 26 268
use FILL  FILL_9__1928_
timestamp 0
transform -1 0 3290 0 -1 9110
box -6 -8 26 268
use FILL  FILL_9__1943_
timestamp 0
transform -1 0 3710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_9__1958_
timestamp 0
transform -1 0 5290 0 1 11190
box -6 -8 26 268
use FILL  FILL_9__1972_
timestamp 0
transform 1 0 3690 0 1 5470
box -6 -8 26 268
use FILL  FILL_9__1987_
timestamp 0
transform -1 0 7390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_9__2002_
timestamp 0
transform 1 0 6770 0 -1 9110
box -6 -8 26 268
use FILL  FILL_9__2016_
timestamp 0
transform -1 0 7430 0 1 9630
box -6 -8 26 268
use FILL  FILL_9__2031_
timestamp 0
transform -1 0 11150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__2046_
timestamp 0
transform 1 0 8950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_9__2061_
timestamp 0
transform 1 0 10210 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__2075_
timestamp 0
transform -1 0 9690 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__2090_
timestamp 0
transform 1 0 12130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_9__2105_
timestamp 0
transform -1 0 11690 0 1 3390
box -6 -8 26 268
use FILL  FILL_9__2119_
timestamp 0
transform 1 0 10770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_9__2134_
timestamp 0
transform -1 0 7390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_9__2149_
timestamp 0
transform 1 0 10150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_9__2164_
timestamp 0
transform 1 0 9870 0 -1 9630
box -6 -8 26 268
use FILL  FILL_9__2178_
timestamp 0
transform -1 0 11110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_9__2193_
timestamp 0
transform -1 0 11110 0 1 3910
box -6 -8 26 268
use FILL  FILL_9__2208_
timestamp 0
transform -1 0 9470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__2223_
timestamp 0
transform -1 0 11950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_9__2237_
timestamp 0
transform -1 0 6750 0 1 4950
box -6 -8 26 268
use FILL  FILL_9__2252_
timestamp 0
transform 1 0 11390 0 1 9110
box -6 -8 26 268
use FILL  FILL_9__2267_
timestamp 0
transform 1 0 12050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_9__2281_
timestamp 0
transform 1 0 12170 0 1 6510
box -6 -8 26 268
use FILL  FILL_9__2296_
timestamp 0
transform 1 0 11270 0 -1 7030
box -6 -8 26 268
use FILL  FILL_9__2311_
timestamp 0
transform 1 0 11670 0 1 8070
box -6 -8 26 268
use FILL  FILL_9__2326_
timestamp 0
transform 1 0 12190 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__2340_
timestamp 0
transform -1 0 9990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_9__2355_
timestamp 0
transform -1 0 7030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__2370_
timestamp 0
transform -1 0 7390 0 1 10150
box -6 -8 26 268
use FILL  FILL_9__2384_
timestamp 0
transform 1 0 4750 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__2399_
timestamp 0
transform 1 0 2030 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__2414_
timestamp 0
transform 1 0 3150 0 1 5470
box -6 -8 26 268
use FILL  FILL_9__2429_
timestamp 0
transform -1 0 5210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_9__2443_
timestamp 0
transform -1 0 7290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_9__2458_
timestamp 0
transform -1 0 4990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_9__2473_
timestamp 0
transform 1 0 2010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_9__2487_
timestamp 0
transform 1 0 2470 0 1 4430
box -6 -8 26 268
use FILL  FILL_9__2502_
timestamp 0
transform -1 0 3110 0 1 4430
box -6 -8 26 268
use FILL  FILL_9__2517_
timestamp 0
transform -1 0 2310 0 1 270
box -6 -8 26 268
use FILL  FILL_9__2532_
timestamp 0
transform 1 0 4310 0 1 270
box -6 -8 26 268
use FILL  FILL_9__2546_
timestamp 0
transform 1 0 4910 0 1 3390
box -6 -8 26 268
use FILL  FILL_9__2561_
timestamp 0
transform 1 0 3710 0 1 1310
box -6 -8 26 268
use FILL  FILL_9__2576_
timestamp 0
transform -1 0 4330 0 1 7550
box -6 -8 26 268
use FILL  FILL_9__2591_
timestamp 0
transform 1 0 6570 0 1 1310
box -6 -8 26 268
use FILL  FILL_9__2605_
timestamp 0
transform 1 0 6170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_9__2620_
timestamp 0
transform -1 0 730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_9__2635_
timestamp 0
transform 1 0 190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_9__2649_
timestamp 0
transform 1 0 190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_9__2664_
timestamp 0
transform 1 0 1010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_9__2679_
timestamp 0
transform 1 0 7130 0 1 1310
box -6 -8 26 268
use FILL  FILL_9__2694_
timestamp 0
transform -1 0 1470 0 -1 790
box -6 -8 26 268
use FILL  FILL_9__2708_
timestamp 0
transform 1 0 2550 0 -1 790
box -6 -8 26 268
use FILL  FILL_9__2723_
timestamp 0
transform 1 0 2730 0 1 790
box -6 -8 26 268
use FILL  FILL_9__2738_
timestamp 0
transform -1 0 3950 0 1 1830
box -6 -8 26 268
use FILL  FILL_9__2752_
timestamp 0
transform 1 0 1250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_9__2767_
timestamp 0
transform -1 0 1630 0 1 1310
box -6 -8 26 268
use FILL  FILL_9__2782_
timestamp 0
transform 1 0 7870 0 1 270
box -6 -8 26 268
use FILL  FILL_9__2797_
timestamp 0
transform 1 0 10930 0 -1 8070
box -6 -8 26 268
use FILL  FILL_9__2811_
timestamp 0
transform 1 0 10150 0 -1 9630
box -6 -8 26 268
use FILL  FILL_9__2826_
timestamp 0
transform 1 0 8850 0 -1 7550
box -6 -8 26 268
use FILL  FILL_9__2841_
timestamp 0
transform 1 0 8330 0 -1 11190
box -6 -8 26 268
use FILL  FILL_9__2856_
timestamp 0
transform -1 0 9190 0 1 10670
box -6 -8 26 268
use FILL  FILL_9__2870_
timestamp 0
transform 1 0 8710 0 1 9110
box -6 -8 26 268
use FILL  FILL_9__2885_
timestamp 0
transform -1 0 10630 0 1 9630
box -6 -8 26 268
use FILL  FILL_9__2900_
timestamp 0
transform 1 0 10510 0 1 11190
box -6 -8 26 268
use FILL  FILL_9__2914_
timestamp 0
transform -1 0 7910 0 -1 12230
box -6 -8 26 268
use FILL  FILL_9__2929_
timestamp 0
transform -1 0 10470 0 1 11710
box -6 -8 26 268
use FILL  FILL_9__2944_
timestamp 0
transform 1 0 5490 0 -1 8590
box -6 -8 26 268
use FILL  FILL_9__2959_
timestamp 0
transform 1 0 6390 0 -1 7030
box -6 -8 26 268
use FILL  FILL_9__2973_
timestamp 0
transform -1 0 6450 0 1 8070
box -6 -8 26 268
use FILL  FILL_9__2988_
timestamp 0
transform -1 0 6430 0 1 5990
box -6 -8 26 268
use FILL  FILL_9__3003_
timestamp 0
transform -1 0 5950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__3017_
timestamp 0
transform -1 0 6990 0 -1 8070
box -6 -8 26 268
use FILL  FILL_9__3032_
timestamp 0
transform -1 0 5310 0 -1 9110
box -6 -8 26 268
use FILL  FILL_9__3047_
timestamp 0
transform -1 0 3190 0 1 7550
box -6 -8 26 268
use FILL  FILL_9__3062_
timestamp 0
transform -1 0 3950 0 -1 11710
box -6 -8 26 268
use FILL  FILL_9__3076_
timestamp 0
transform 1 0 3790 0 -1 7030
box -6 -8 26 268
use FILL  FILL_9__3091_
timestamp 0
transform -1 0 6350 0 -1 11190
box -6 -8 26 268
use FILL  FILL_9__3106_
timestamp 0
transform -1 0 6050 0 -1 11190
box -6 -8 26 268
use FILL  FILL_9__3120_
timestamp 0
transform 1 0 4710 0 1 10150
box -6 -8 26 268
use FILL  FILL_9__3135_
timestamp 0
transform 1 0 4930 0 1 11710
box -6 -8 26 268
use FILL  FILL_9__3150_
timestamp 0
transform -1 0 11890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_9__3165_
timestamp 0
transform -1 0 7310 0 1 1830
box -6 -8 26 268
use FILL  FILL_9__3179_
timestamp 0
transform 1 0 12170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_9__3194_
timestamp 0
transform 1 0 10910 0 1 2350
box -6 -8 26 268
use FILL  FILL_9__3209_
timestamp 0
transform -1 0 770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_9__3224_
timestamp 0
transform -1 0 3410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_9__3369_
timestamp 0
transform -1 0 5670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__3384_
timestamp 0
transform 1 0 1870 0 -1 8590
box -6 -8 26 268
use FILL  FILL_9__3399_
timestamp 0
transform 1 0 190 0 1 8070
box -6 -8 26 268
use FILL  FILL_9__3413_
timestamp 0
transform 1 0 470 0 1 7030
box -6 -8 26 268
use FILL  FILL_9__3428_
timestamp 0
transform 1 0 1230 0 1 9630
box -6 -8 26 268
use FILL  FILL_9__3443_
timestamp 0
transform 1 0 1230 0 -1 10670
box -6 -8 26 268
use FILL  FILL_9__3458_
timestamp 0
transform -1 0 1850 0 1 10150
box -6 -8 26 268
use FILL  FILL_9__3472_
timestamp 0
transform -1 0 2330 0 -1 10670
box -6 -8 26 268
use FILL  FILL_9__3487_
timestamp 0
transform -1 0 1830 0 -1 11710
box -6 -8 26 268
use FILL  FILL_9__3502_
timestamp 0
transform -1 0 510 0 1 10670
box -6 -8 26 268
use FILL  FILL_9__3516_
timestamp 0
transform -1 0 210 0 1 10150
box -6 -8 26 268
use FILL  FILL_9__3531_
timestamp 0
transform 1 0 190 0 -1 10150
box -6 -8 26 268
use FILL  FILL_9__3546_
timestamp 0
transform 1 0 2010 0 -1 12230
box -6 -8 26 268
use FILL  FILL_9__3561_
timestamp 0
transform -1 0 2070 0 1 7550
box -6 -8 26 268
use FILL  FILL_9__3587_
timestamp 0
transform 1 0 190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9__3602_
timestamp 0
transform -1 0 1830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert9
timestamp 0
transform 1 0 10250 0 1 3910
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert24
timestamp 0
transform -1 0 4450 0 1 5470
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert39
timestamp 0
transform 1 0 6450 0 1 4950
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert53
timestamp 0
transform 1 0 10110 0 1 1310
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert68
timestamp 0
transform 1 0 3270 0 1 270
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert83
timestamp 0
transform -1 0 7490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_9_BUFX2_insert97
timestamp 0
transform 1 0 11570 0 1 11710
box -6 -8 26 268
<< labels >>
flabel metal1 s 12343 2 12403 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 5917 -23 5923 -17 7 FreeSans 16 270 0 0 AB[15]
port 2 nsew
flabel metal2 s 3077 -23 3083 -17 7 FreeSans 16 270 0 0 AB[14]
port 3 nsew
flabel metal2 s 4657 -23 4663 -17 7 FreeSans 16 270 0 0 AB[13]
port 4 nsew
flabel metal2 s 5457 -23 5463 -17 7 FreeSans 16 270 0 0 AB[12]
port 5 nsew
flabel metal2 s 3337 -23 3343 -17 7 FreeSans 16 270 0 0 AB[11]
port 6 nsew
flabel metal2 s 3597 -23 3603 -17 7 FreeSans 16 270 0 0 AB[10]
port 7 nsew
flabel metal2 s 5977 -23 5983 -17 7 FreeSans 16 270 0 0 AB[9]
port 8 nsew
flabel metal2 s 4917 -23 4923 -17 7 FreeSans 16 270 0 0 AB[8]
port 9 nsew
flabel metal3 s -24 4556 -16 4564 7 FreeSans 16 0 0 0 AB[7]
port 10 nsew
flabel metal3 s -24 5896 -16 5904 7 FreeSans 16 0 0 0 AB[6]
port 11 nsew
flabel metal3 s -24 5336 -16 5344 7 FreeSans 16 0 0 0 AB[5]
port 12 nsew
flabel metal3 s -24 5076 -16 5084 7 FreeSans 16 0 0 0 AB[4]
port 13 nsew
flabel metal3 s -24 4036 -16 4044 7 FreeSans 16 0 0 0 AB[3]
port 14 nsew
flabel metal3 s -24 6156 -16 6164 7 FreeSans 16 0 0 0 AB[2]
port 15 nsew
flabel metal3 s -24 4296 -16 4304 7 FreeSans 16 0 0 0 AB[1]
port 16 nsew
flabel metal2 s 5177 -23 5183 -17 7 FreeSans 16 270 0 0 AB[0]
port 17 nsew
flabel metal2 s 6037 -23 6043 -17 7 FreeSans 16 270 0 0 DI[7]
port 18 nsew
flabel metal3 s -24 6416 -16 6424 7 FreeSans 16 0 0 0 DI[6]
port 19 nsew
flabel metal3 s -24 4816 -16 4824 7 FreeSans 16 0 0 0 DI[5]
port 20 nsew
flabel metal3 s -24 5596 -16 5604 7 FreeSans 16 0 0 0 DI[4]
port 21 nsew
flabel metal3 s -24 3776 -16 3784 7 FreeSans 16 0 0 0 DI[3]
port 22 nsew
flabel metal3 s -24 6676 -16 6684 7 FreeSans 16 0 0 0 DI[2]
port 23 nsew
flabel metal2 s 457 -23 463 -17 7 FreeSans 16 270 0 0 DI[1]
port 24 nsew
flabel metal3 s -24 4596 -16 4604 7 FreeSans 16 0 0 0 DI[0]
port 25 nsew
flabel metal3 s -24 5856 -16 5864 7 FreeSans 16 0 0 0 DO[7]
port 26 nsew
flabel metal3 s -24 5636 -16 5644 7 FreeSans 16 0 0 0 DO[6]
port 27 nsew
flabel metal3 s -24 6376 -16 6384 7 FreeSans 16 0 0 0 DO[5]
port 28 nsew
flabel metal3 s -24 6636 -16 6644 7 FreeSans 16 0 0 0 DO[4]
port 29 nsew
flabel metal3 s -24 6116 -16 6124 7 FreeSans 16 0 0 0 DO[3]
port 30 nsew
flabel metal3 s -24 6196 -16 6204 7 FreeSans 16 0 0 0 DO[2]
port 31 nsew
flabel metal3 s -24 5936 -16 5944 7 FreeSans 16 0 0 0 DO[1]
port 32 nsew
flabel metal2 s 5717 -23 5723 -17 7 FreeSans 16 270 0 0 DO[0]
port 33 nsew
flabel metal2 s 6777 -23 6783 -17 7 FreeSans 16 270 0 0 IRQ
port 34 nsew
flabel metal2 s 7517 -23 7523 -17 7 FreeSans 16 270 0 0 NMI
port 35 nsew
flabel metal3 s 12376 3816 12384 3824 3 FreeSans 16 0 0 0 RDY
port 36 nsew
flabel metal2 s 7017 -23 7023 -17 7 FreeSans 16 270 0 0 WE
port 37 nsew
flabel metal2 s 5437 12277 5443 12283 3 FreeSans 16 90 0 0 clk
port 38 nsew
flabel metal2 s 4097 12277 4103 12283 3 FreeSans 16 90 0 0 reset
port 39 nsew
<< properties >>
string FIXED_BBOX -40 -40 12380 12280
<< end >>
