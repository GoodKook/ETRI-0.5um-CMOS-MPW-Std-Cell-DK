magic
tech scmos
magscale 1 2
timestamp 1702316108
<< nwell >>
rect -13 154 235 272
rect 8 152 47 154
<< ntransistor >>
rect 16 14 20 54
rect 36 14 40 34
rect 48 14 52 34
rect 68 14 72 34
rect 78 14 82 34
rect 100 14 104 34
rect 140 14 144 34
rect 150 14 154 34
rect 170 14 174 34
rect 180 14 184 34
rect 200 14 204 54
<< ptransistor >>
rect 16 166 20 246
rect 36 206 40 246
rect 48 206 52 246
rect 68 206 72 246
rect 80 206 84 246
rect 100 206 104 246
rect 140 206 144 246
rect 150 206 154 246
rect 170 226 174 246
rect 180 226 184 246
rect 200 166 204 246
<< ndiffusion >>
rect 14 14 16 54
rect 20 14 22 54
rect 34 14 36 34
rect 40 14 48 34
rect 52 14 54 34
rect 66 14 68 34
rect 72 14 78 34
rect 82 14 84 34
rect 96 14 100 34
rect 104 14 106 34
rect 138 14 140 34
rect 144 14 150 34
rect 154 14 156 34
rect 168 14 170 34
rect 174 14 180 34
rect 184 14 186 34
rect 198 14 200 54
rect 204 14 206 54
<< pdiffusion >>
rect 14 166 16 246
rect 20 169 22 246
rect 34 206 36 246
rect 40 206 48 246
rect 52 206 54 246
rect 66 206 68 246
rect 72 206 80 246
rect 84 206 86 246
rect 98 206 100 246
rect 104 206 106 246
rect 138 206 140 246
rect 144 206 150 246
rect 154 206 156 246
rect 168 226 170 246
rect 174 226 180 246
rect 184 226 186 246
rect 20 166 34 169
rect 198 166 200 246
rect 204 166 206 246
<< ndcontact >>
rect 2 14 14 54
rect 22 14 34 54
rect 54 14 66 34
rect 84 14 96 34
rect 106 14 118 34
rect 126 14 138 34
rect 156 14 168 34
rect 186 14 198 54
rect 206 14 218 54
<< pdcontact >>
rect 2 166 14 246
rect 22 169 34 246
rect 54 206 66 246
rect 86 206 98 246
rect 106 206 118 246
rect 126 206 138 246
rect 156 206 168 246
rect 186 166 198 246
rect 206 166 218 246
<< psubstratepcontact >>
rect -6 -6 226 6
<< nsubstratencontact >>
rect -6 254 226 266
<< polysilicon >>
rect 16 246 20 250
rect 36 246 40 250
rect 48 246 52 250
rect 68 246 72 250
rect 80 246 84 250
rect 100 246 104 250
rect 140 246 144 250
rect 150 246 154 250
rect 170 246 174 250
rect 180 246 184 250
rect 200 246 204 250
rect 16 80 20 166
rect 36 131 40 206
rect 48 162 52 206
rect 68 200 72 206
rect 80 200 84 206
rect 60 150 72 154
rect 36 119 43 131
rect 16 54 20 68
rect 36 34 40 119
rect 48 34 52 56
rect 68 34 72 150
rect 80 54 84 188
rect 100 100 104 206
rect 140 204 144 206
rect 78 52 84 54
rect 78 40 80 52
rect 78 34 82 40
rect 100 34 104 88
rect 112 200 144 204
rect 150 197 154 206
rect 148 192 154 197
rect 112 40 116 188
rect 126 50 130 168
rect 148 76 152 192
rect 170 184 174 226
rect 172 172 174 184
rect 180 152 184 226
rect 200 96 204 166
rect 196 84 204 96
rect 150 68 152 76
rect 150 64 164 68
rect 160 50 164 64
rect 126 46 154 50
rect 160 46 174 50
rect 112 36 144 40
rect 140 34 144 36
rect 150 34 154 46
rect 170 34 174 46
rect 180 34 184 63
rect 200 54 204 84
rect 16 10 20 14
rect 36 10 40 14
rect 48 10 52 14
rect 68 10 72 14
rect 78 10 82 14
rect 100 10 104 14
rect 140 10 144 14
rect 150 10 154 14
rect 170 10 174 14
rect 180 10 184 14
rect 200 10 204 14
<< polycontact >>
rect 60 188 72 200
rect 80 188 92 200
rect 48 150 60 162
rect 43 119 55 131
rect 14 68 26 80
rect 48 56 60 68
rect 92 88 104 100
rect 80 40 92 52
rect 112 188 124 200
rect 126 168 138 180
rect 160 172 172 184
rect 176 140 188 152
rect 184 84 196 96
rect 138 64 150 76
rect 176 63 188 75
<< metal1 >>
rect -6 266 226 268
rect -6 252 226 254
rect 22 246 34 252
rect 86 246 98 252
rect 126 246 138 252
rect 186 246 198 252
rect 40 206 54 214
rect 106 200 112 206
rect 92 194 112 200
rect 60 182 72 188
rect 138 172 160 180
rect 2 162 14 166
rect 126 162 132 168
rect 2 156 48 162
rect 2 54 8 156
rect 60 154 132 162
rect 206 152 214 166
rect 188 140 214 152
rect 203 137 214 140
rect 18 123 37 137
rect 18 80 26 123
rect 83 128 97 137
rect 55 119 97 128
rect 203 123 217 137
rect 53 94 92 100
rect 26 74 58 76
rect 168 84 184 96
rect 72 74 138 76
rect 26 68 138 74
rect 206 71 214 123
rect 188 63 214 71
rect 206 54 214 63
rect 92 40 112 46
rect 106 34 112 40
rect 42 27 54 34
rect 154 28 156 34
rect 22 8 34 14
rect 84 8 96 14
rect 126 8 138 14
rect 186 8 198 14
rect -6 6 226 8
rect -6 -8 226 -6
<< m2contact >>
rect 40 192 54 206
rect 154 192 168 206
rect 60 168 74 182
rect 39 92 53 106
rect 58 74 72 88
rect 154 84 168 98
rect 42 34 56 48
rect 154 34 168 48
<< metal2 >>
rect 43 106 50 192
rect 154 180 162 192
rect 154 172 160 180
rect 43 48 50 92
rect 63 88 72 168
rect 154 98 162 172
rect 154 48 162 84
<< m1p >>
rect -6 252 226 268
rect 23 123 37 137
rect 83 123 97 137
rect 203 123 217 137
rect -6 -8 226 8
<< labels >>
rlabel nsubstratencontact 110 260 110 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 110 0 110 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 30 131 30 131 0 CLK
port 2 nsew clock input
rlabel metal1 90 130 90 130 0 D
port 1 nsew signal input
rlabel metal1 210 131 210 131 0 Q
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 220 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
