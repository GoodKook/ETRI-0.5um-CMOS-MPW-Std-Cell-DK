/* Verilog module written by vlog2Verilog (qflow) */

module fir8(
    input [7:0] Xin,
    output [7:0] Xout,
    input [15:0] Yin,
    output [15:0] Yout,
    input clk
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire [15:5] _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire [15:0] \u_fir_pe2.mul  ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _2712_ ;
wire _5184_ ;
wire \X[1]_5_bF$buf0  ;
wire _3917_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire [15:0] \u_fir_pe4.mul  ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire [2:2] _4778_ ;
wire _4358_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6313_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6122_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6351_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6160_ ;
wire [15:0] \u_fir_pe6.mul  ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6254_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6063_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire [15:0] \Y[4]  ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire [15:1] _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6251_ ;
wire _2591_ ;
wire _2171_ ;
wire _3796_ ;
wire _3376_ ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire \X[6]_5_bF$buf1  ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire [15:0] \u_fir_pe4.rYin  ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6060_ ;
wire [3:3] _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6057_ ;
wire _1192_ ;
wire [7:0] \X[2]  ;
wire _2397_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _197_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6210_ ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire [15:5] _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire \X[5]_5_bF$buf3  ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire [0:0] _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6113_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _5783_ ;
wire _5363_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire [15:0] _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire [2:2] _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire [15:0] \u_fir_pe2.rYin  ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire \X[5]_5_bF$buf0  ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire [15:1] _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _5704_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6242_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire Xin_5_bF$buf0 ;
wire Xin_5_bF$buf1 ;
wire Xin_5_bF$buf2 ;
wire Xin_5_bF$buf3 ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire [4:4] _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _5683_ ;
wire _5263_ ;
wire _6048_ ;
wire _1183_ ;
wire [3:3] _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire \X[4]_5_bF$buf2  ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire [15:0] \u_fir_pe7.rYin  ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6201_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire [1:1] _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6045_ ;
wire _1180_ ;
wire [0:0] _2385_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6274_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire [15:5] _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire [15:0] \Y[6]  ;
wire _5583_ ;
wire _5163_ ;
wire [0:0] _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire _5601_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6233_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6271_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire [2:2] _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire \X[3]_5_bF$buf1  ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6365_ ;
wire _1080_ ;
wire [15:0] \u_fir_pe5.rYin  ;
wire _2285_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _5674_ ;
wire _5254_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire _5483_ ;
wire _5063_ ;
wire _6268_ ;
wire _2188_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6077_ ;
wire [7:0] \X[4]  ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire [4:4] _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6230_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6324_ ;
wire [15:1] _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire \X[2]_5_bF$buf3  ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _5633_ ;
wire _5213_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6036_ ;
wire [3:3] _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6265_ ;
wire _2185_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _5994_ ;
wire [1:1] _5574_ ;
wire _5154_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire _5383_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire _2088_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire [0:0] _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6321_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire \X[2]_5_bF$buf0  ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6224_ ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _5724_ ;
wire _5304_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6262_ ;
wire _2182_ ;
wire [15:0] \Y[1]  ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire [0:0] _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _4707_ ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6068_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire \X[1]_5_bF$buf2  ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6221_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _6353_ ;
wire _2693_ ;
wire _2273_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6162_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _4704_ ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire \X[7]_5_bF$buf1  ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire [4:4] _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire [1:1] _4777_ ;
wire _4357_ ;
wire _56_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6312_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6121_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6350_ ;
wire [15:0] \u_fir_pe5.mul  ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6253_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire \X[6]_5_bF$buf3  ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6062_ ;
wire [15:0] \u_fir_pe7.mul  ;
wire [15:5] _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6059_ ;
wire _1194_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire [0:0] _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire [7:0] \X[6]  ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _199_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6250_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire \X[6]_5_bF$buf0  ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire [2:2] _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire [15:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _196_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _1094_ ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire [4:4] _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire \X[5]_5_bF$buf2  ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire [15:1] _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _5803_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6244_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire [15:0] \Y[3]  ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire [7:0] _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire _1185_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6279_ ;
wire _2199_ ;
wire [1:1] _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire [0:0] _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _5703_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6241_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6050_ ;
wire [15:5] _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire [3:3] _6373_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _5644_ ;
wire _5224_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire [15:0] \u_fir_pe0.rYin  ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6047_ ;
wire _1182_ ;
wire [7:0] \X[1]  ;
wire [2:2] _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire \X[4]_5_bF$buf1  ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire _2731_ ;
wire _2311_ ;
wire [15:0] Yout ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6200_ ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire [0:0] _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6044_ ;
wire [15:1] _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6273_ ;
wire _2193_ ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire [4:4] _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire \X[3]_5_bF$buf3  ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4624_ ;
wire _4204_ ;
wire _5829_ ;
wire _5409_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6079_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _2631_ ;
wire _2211_ ;
wire [7:0] Xout ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6232_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6041_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6270_ ;
wire _2190_ ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire [1:1] _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire \X[3]_5_bF$buf0  ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _4621_ ;
wire _4201_ ;
wire _5826_ ;
wire _5406_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _5673_ ;
wire _5253_ ;
wire _6038_ ;
wire [15:5] _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire _6267_ ;
wire _2187_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire [0:0] _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire [3:3] _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire [15:0] \u_fir_pe3.rYin  ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire \X[2]_5_bF$buf2  ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _3677_ ;
wire _3257_ ;
wire _5823_ ;
wire _5403_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6035_ ;
wire [2:2] _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6264_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire [15:0] \Y[5]  ;
wire _5993_ ;
wire [0:0] _5573_ ;
wire _5153_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6167_ ;
wire _2087_ ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _4709_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire [15:1] _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6320_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6223_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _5723_ ;
wire _5303_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6261_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _4706_ ;
wire _3098_ ;
wire _5664_ ;
wire _5244_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire [15:0] \u_fir_pe1.mul  ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire \X[7]_5_bF$buf3  ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6067_ ;
wire [7:0] \X[3]  ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _1678_ ;
wire _1258_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire [15:0] \u_fir_pe3.mul  ;
wire \X[1]_5_bF$buf1  ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6220_ ;
wire _1199_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire [3:3] _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6123_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6352_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6161_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire \X[7]_5_bF$buf0  ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire [15:0] \u_fir_pe6.rYin  ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire [0:0] _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6311_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6120_ ;
wire _1099_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6252_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire \X[6]_5_bF$buf2  ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6061_ ;
wire [4:4] _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _198_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6211_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _3794_ ;
wire _3374_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire [1:1] _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _5708_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _5784_ ;
wire _5364_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire [15:0] \Y[7]  ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire [3:3] _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire \X[5]_5_bF$buf1  ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire [0:0] _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6111_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6014_ ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire [0:0] _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5705_ ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6243_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire [15:5] _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire _6049_ ;
wire _1184_ ;
wire [4:4] _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire [7:0] \X[5]  ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire \X[4]_5_bF$buf3  ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6240_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _5605_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _1754_ ;
wire _1334_ ;
wire [7:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire [2:2] _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _5643_ ;
wire _5223_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6046_ ;
wire _1181_ ;
wire [1:1] _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire \X[4]_5_bF$buf0  ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _5584_ ;
wire _5164_ ;
wire [15:1] _6369_ ;
wire _1084_ ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6178_ ;
wire _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _1598_ ;
wire _1178_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire _5602_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _3494_ ;
wire _3074_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6234_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6043_ ;
wire [0:0] _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6272_ ;
wire _2192_ ;
wire [15:0] \Y[2]  ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire [3:3] _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire \X[3]_5_bF$buf2  ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _4623_ ;
wire _4203_ ;
wire _5828_ ;
wire _5408_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _5484_ ;
wire _5064_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire [15:5] _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire _4238_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6231_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6040_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire [0:0] _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6363_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6037_ ;
wire [4:4] _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6266_ ;
wire _2186_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6075_ ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire [2:2] _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire [1:1] _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6322_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire \X[2]_5_bF$buf1  ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6360_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6034_ ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6263_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6072_ ;
wire _4805_ ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire [15:1] _5572_ ;
wire _5152_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6166_ ;
wire _2086_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _4708_ ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire [0:0] _1586_ ;
wire _1166_ ;
wire [15:0] \u_fir_pe1.rYin  ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6069_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire [7:0] \X[7]  ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire \X[1]_5_bF$buf3  ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6222_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6031_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _5722_ ;
wire _5302_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6260_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6354_ ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6163_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire [15:0] \u_fir_pe0.mul  ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire \X[7]_5_bF$buf2  ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire [7:1] \X  ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6066_ ;

INVX1 _11689_ (
    .A(_4810_),
    .Y(_4811_)
);

OAI21X1 _11269_ (
    .A(_4059_),
    .B(_4304_),
    .C(_4458_),
    .Y(_4465_)
);

FILL FILL_2__7905_ (
);

FILL FILL_0__12765_ (
);

NAND3X1 _12630_ (
    .A(vdd),
    .B(\X[6] [3]),
    .C(_5662_),
    .Y(_5671_)
);

FILL FILL_0__12345_ (
);

INVX1 _12210_ (
    .A(_5297_),
    .Y(_5325_)
);

DFFPOSX1 _9837_ (
    .D(_3181_[7]),
    .CLK(clk_bF$buf53),
    .Q(\Y[4] [7])
);

OAI21X1 _9417_ (
    .A(_2695_),
    .B(_2699_),
    .C(_2704_),
    .Y(_2774_)
);

FILL FILL_1__8794_ (
);

FILL FILL_1__8374_ (
);

FILL FILL_3__9661_ (
);

BUFX2 _13415_ (
    .A(_6377_[7]),
    .Y(Yout[7])
);

FILL FILL_1__9999_ (
);

FILL FILL_1__9579_ (
);

FILL FILL_1__9159_ (
);

FILL FILL_2__11484_ (
);

FILL FILL_2__11064_ (
);

FILL FILL_1__10897_ (
);

FILL FILL_1__10477_ (
);

FILL FILL_1__10057_ (
);

FILL FILL_0__7484_ (
);

NAND3X1 _9590_ (
    .A(_2902_),
    .B(_2944_),
    .C(_2903_),
    .Y(_2945_)
);

FILL FILL_0__7064_ (
);

NAND2X1 _9170_ (
    .A(\X[3] [1]),
    .B(vdd),
    .Y(_2530_)
);

FILL FILL_3__10804_ (
);

FILL FILL_2__8863_ (
);

FILL FILL_2__8443_ (
);

FILL FILL_0__10831_ (
);

FILL FILL_3__13276_ (
);

FILL FILL_0__10411_ (
);

FILL FILL_2__8023_ (
);

FILL FILL_2__12689_ (
);

FILL FILL_2__12269_ (
);

AND2X2 _7903_ (
    .A(_1393_),
    .B(_1392_),
    .Y(_1415_)
);

FILL FILL_1__6860_ (
);

FILL FILL_1__6440_ (
);

FILL FILL_0__8689_ (
);

FILL FILL_2__13210_ (
);

FILL FILL_3__6786_ (
);

FILL FILL_0__8269_ (
);

FILL FILL_1__12623_ (
);

FILL FILL_1__12203_ (
);

FILL FILL_0__9630_ (
);

FILL FILL_2__9648_ (
);

FILL FILL_0__9210_ (
);

FILL FILL_2__9228_ (
);

NAND2X1 _11901_ (
    .A(_5014_),
    .B(_5019_),
    .Y(_5020_)
);

FILL FILL_1__7645_ (
);

FILL FILL_1__13408_ (
);

FILL FILL_3__8932_ (
);

OAI21X1 _10293_ (
    .A(_3489_),
    .B(_3569_),
    .C(_3552_),
    .Y(_3570_)
);

FILL FILL_3__11762_ (
);

FILL FILL_3__11342_ (
);

FILL FILL_2__10335_ (
);

FILL FILL_3__9717_ (
);

FILL FILL_0__6755_ (
);

INVX1 _8861_ (
    .A(\u_fir_pe2.rYin [8]),
    .Y(_2284_)
);

NAND3X1 _8441_ (
    .A(_1875_),
    .B(_1876_),
    .C(_1877_),
    .Y(_1880_)
);

NOR2X1 _8021_ (
    .A(_1524_),
    .B(_1523_),
    .Y(_1525_)
);

NAND2X1 _11498_ (
    .A(_4660_),
    .B(_4672_),
    .Y(_4681_)
);

AOI21X1 _11078_ (
    .A(_4272_),
    .B(_4271_),
    .C(_4173_),
    .Y(_4277_)
);

FILL FILL_2__7714_ (
);

FILL FILL_3__12547_ (
);

FILL FILL_3__12127_ (
);

FILL FILL_1__13161_ (
);

FILL FILL_0__12994_ (
);

FILL FILL_0__12574_ (
);

FILL FILL_0__12154_ (
);

FILL FILL_2__12901_ (
);

NAND2X1 _9646_ (
    .A(_2997_),
    .B(_2998_),
    .Y(_2999_)
);

AOI21X1 _9226_ (
    .A(_2509_),
    .B(_2508_),
    .C(_2445_),
    .Y(_2586_)
);

FILL FILL_1__8183_ (
);

FILL FILL_0__8901_ (
);

FILL FILL_2__8919_ (
);

FILL FILL_3__9050_ (
);

NAND2X1 _13224_ (
    .A(_6248_),
    .B(_6243_),
    .Y(_6249_)
);

FILL FILL_1__6916_ (
);

FILL FILL_1__9388_ (
);

FILL FILL_2__11293_ (
);

FILL FILL_1__10286_ (
);

FILL FILL_0__7293_ (
);

FILL FILL_3__10613_ (
);

FILL FILL_2__8672_ (
);

FILL FILL_2__8252_ (
);

FILL FILL_0__10640_ (
);

FILL FILL_0__10220_ (
);

FILL FILL_2__12078_ (
);

INVX1 _7712_ (
    .A(_1151_),
    .Y(_1229_)
);

FILL FILL_0__8498_ (
);

AOI22X1 _10769_ (
    .A(\X[5] [0]),
    .B(gnd),
    .C(\X[5] [1]),
    .D(gnd),
    .Y(_4735_)
);

INVX1 _10349_ (
    .A(_3571_),
    .Y(_3626_)
);

FILL FILL_1__12852_ (
);

FILL FILL_1__12432_ (
);

FILL FILL_1__12012_ (
);

FILL FILL_2__9457_ (
);

FILL FILL_0__11845_ (
);

FILL FILL_2__9037_ (
);

NAND2X1 _11710_ (
    .A(_4814_),
    .B(_4829_),
    .Y(_4832_)
);

FILL FILL_0__11425_ (
);

FILL FILL_0__11005_ (
);

NAND2X1 _8917_ (
    .A(_2340_),
    .B(_2335_),
    .Y(_2341_)
);

FILL FILL_1__7874_ (
);

FILL FILL_1__7454_ (
);

FILL FILL_1__7034_ (
);

FILL FILL_1__13217_ (
);

NAND2X1 _12915_ (
    .A(_5952_),
    .B(_5876_),
    .Y(_5953_)
);

FILL FILL_3__8321_ (
);

FILL FILL_3__11991_ (
);

FILL FILL_1__8659_ (
);

FILL FILL_1__8239_ (
);

FILL FILL_3__11571_ (
);

FILL FILL_3__11151_ (
);

FILL FILL_2__10984_ (
);

FILL FILL_2__10564_ (
);

FILL FILL_2__10144_ (
);

FILL FILL_1__9600_ (
);

FILL FILL_3__9946_ (
);

FILL FILL_3__9526_ (
);

FILL FILL_3__9106_ (
);

FILL FILL_0__6984_ (
);

FILL FILL_0__6564_ (
);

NAND3X1 _8670_ (
    .A(_2089_),
    .B(_2095_),
    .C(_2053_),
    .Y(_2105_)
);

INVX1 _8250_ (
    .A(_1678_),
    .Y(_1691_)
);

FILL FILL_2__7943_ (
);

FILL FILL_3__12776_ (
);

FILL FILL_2__7523_ (
);

FILL FILL_3__12356_ (
);

FILL FILL_2__7103_ (
);

FILL FILL_2__11769_ (
);

FILL FILL_2__11349_ (
);

FILL FILL_0__12383_ (
);

FILL FILL_2__12710_ (
);

FILL FILL_0__7769_ (
);

DFFPOSX1 _9875_ (
    .D(_3187_[5]),
    .CLK(clk_bF$buf14),
    .Q(\u_fir_pe3.mul [5])
);

FILL FILL_0__7349_ (
);

NAND2X1 _9455_ (
    .A(_2797_),
    .B(_2800_),
    .Y(_2812_)
);

NOR2X1 _9035_ (
    .A(_3122_),
    .B(_2393_),
    .Y(_2398_)
);

FILL FILL_1__11703_ (
);

FILL FILL_0__8710_ (
);

FILL FILL_2__8728_ (
);

FILL FILL_2__8308_ (
);

FILL FILL_0__13168_ (
);

NAND3X1 _13033_ (
    .A(_5986_),
    .B(_6062_),
    .C(_5994_),
    .Y(_6069_)
);

FILL FILL_1__6725_ (
);

FILL FILL_1__9197_ (
);

FILL FILL_1__12908_ (
);

FILL FILL_0__9915_ (
);

FILL FILL_1__10095_ (
);

FILL FILL_3__10842_ (
);

FILL FILL_3__10002_ (
);

FILL FILL_2__8481_ (
);

FILL FILL_2__8061_ (
);

NOR2X1 _7941_ (
    .A(\u_fir_pe1.rYin [3]),
    .B(\u_fir_pe1.mul [3]),
    .Y(_1448_)
);

NAND2X1 _7521_ (
    .A(_1038_),
    .B(_1039_),
    .Y(_1040_)
);

NOR2X1 _7101_ (
    .A(\u_fir_pe0.rYin [7]),
    .B(\u_fir_pe0.mul [7]),
    .Y(_684_)
);

NAND2X1 _10998_ (
    .A(\X[5] [1]),
    .B(gnd),
    .Y(_4197_)
);

INVX1 _10578_ (
    .A(\u_fir_pe4.mul [4]),
    .Y(_3844_)
);

INVX1 _10158_ (
    .A(_3436_),
    .Y(_3437_)
);

FILL FILL_1__12661_ (
);

FILL FILL_1__12241_ (
);

FILL FILL_2__9686_ (
);

FILL FILL_2__9266_ (
);

FILL FILL_0__11654_ (
);

FILL FILL_0__11234_ (
);

NOR2X1 _8726_ (
    .A(_2067_),
    .B(_2120_),
    .Y(_2160_)
);

AND2X2 _8306_ (
    .A(_1741_),
    .B(_1745_),
    .Y(_1746_)
);

FILL FILL_1__7683_ (
);

FILL FILL_1__7263_ (
);

FILL FILL_1__13026_ (
);

FILL FILL_0__12859_ (
);

FILL FILL_3__8550_ (
);

OAI21X1 _12724_ (
    .A(_5759_),
    .B(_5760_),
    .C(_5717_),
    .Y(_5764_)
);

FILL FILL_0__12439_ (
);

FILL FILL_0__12019_ (
);

AND2X2 _12304_ (
    .A(\u_fir_pe6.rYin [0]),
    .B(\u_fir_pe6.mul [0]),
    .Y(_5413_)
);

FILL FILL_1__8888_ (
);

FILL FILL_1__8468_ (
);

FILL FILL_1__8048_ (
);

FILL FILL_2__10793_ (
);

FILL FILL_2__10373_ (
);

FILL FILL_3__9755_ (
);

FILL FILL_3__9335_ (
);

FILL FILL_0__6793_ (
);

FILL FILL_2__7752_ (
);

FILL FILL_2__7332_ (
);

FILL FILL_2__11998_ (
);

FILL FILL_2__11578_ (
);

FILL FILL_2__11158_ (
);

FILL FILL_0__12192_ (
);

FILL FILL_0__7998_ (
);

FILL FILL_0__7578_ (
);

AND2X2 _9684_ (
    .A(\u_fir_pe3.rYin [2]),
    .B(\u_fir_pe3.mul [2]),
    .Y(_3032_)
);

FILL FILL_0__7158_ (
);

NAND3X1 _9264_ (
    .A(_2617_),
    .B(_2622_),
    .C(_2620_),
    .Y(_2623_)
);

FILL FILL_1__11932_ (
);

FILL FILL_1__11512_ (
);

FILL FILL_2__8537_ (
);

FILL FILL_0__10925_ (
);

FILL FILL_0__10505_ (
);

FILL FILL_0__13397_ (
);

NAND2X1 _13262_ (
    .A(_6284_),
    .B(_6285_),
    .Y(_6286_)
);

FILL FILL_1__6954_ (
);

FILL FILL_1__6534_ (
);

FILL FILL_2__13304_ (
);

FILL FILL_1__12717_ (
);

FILL FILL_0__9724_ (
);

FILL FILL_0__9304_ (
);

FILL FILL_3__7401_ (
);

FILL FILL_1__7739_ (
);

FILL FILL_1__7319_ (
);

FILL FILL_3__10231_ (
);

FILL FILL_2__8290_ (
);

NAND2X1 _6389_ (
    .A(_780_),
    .B(_760_),
    .Y(_781_)
);

NAND3X1 _7750_ (
    .A(_1264_),
    .B(_1261_),
    .C(_1265_),
    .Y(_1266_)
);

NAND2X1 _7330_ (
    .A(_806_),
    .B(_811_),
    .Y(_852_)
);

AND2X2 _10387_ (
    .A(_3661_),
    .B(_3604_),
    .Y(_3663_)
);

FILL FILL_3__11856_ (
);

FILL FILL_2__6603_ (
);

FILL FILL_1__12890_ (
);

FILL FILL_3__11016_ (
);

FILL FILL_1__12050_ (
);

FILL FILL_2__10849_ (
);

FILL FILL_2__9495_ (
);

FILL FILL_0__11883_ (
);

FILL FILL_2__10429_ (
);

FILL FILL_2__9075_ (
);

FILL FILL_0__11463_ (
);

FILL FILL_2__10009_ (
);

FILL FILL_0__11043_ (
);

FILL FILL_0__6849_ (
);

DFFPOSX1 _8955_ (
    .D(_2384_[2]),
    .CLK(clk_bF$buf36),
    .Q(\Y[3] [2])
);

FILL FILL_0__6429_ (
);

NAND2X1 _8535_ (
    .A(_1968_),
    .B(_1972_),
    .Y(_2390_[8])
);

DFFPOSX1 _8115_ (
    .D(\Y[1] [15]),
    .CLK(clk_bF$buf25),
    .Q(\u_fir_pe1.rYin [15])
);

FILL FILL_1__7492_ (
);

FILL FILL_1__7072_ (
);

FILL FILL_2__7808_ (
);

FILL FILL_1__13255_ (
);

NAND2X1 _12953_ (
    .A(_5980_),
    .B(_5989_),
    .Y(_5990_)
);

FILL FILL_0__12668_ (
);

FILL FILL_0__12248_ (
);

INVX1 _12533_ (
    .A(_6364_),
    .Y(_6365_)
);

AOI21X1 _12113_ (
    .A(_5218_),
    .B(_5213_),
    .C(_5165_),
    .Y(_5230_)
);

FILL FILL_1__8697_ (
);

FILL FILL_1__8277_ (
);

FILL FILL_2__10182_ (
);

FILL FILL254250x72150 (
);

NOR2X1 _13318_ (
    .A(\u_fir_pe7.rYin [14]),
    .B(\u_fir_pe7.mul [14]),
    .Y(_6342_)
);

FILL FILL_1_CLKBUF1_insert60 (
);

FILL FILL_1_CLKBUF1_insert61 (
);

FILL FILL_1_CLKBUF1_insert62 (
);

FILL FILL_1_CLKBUF1_insert63 (
);

FILL FILL_1_CLKBUF1_insert64 (
);

FILL FILL_2__7981_ (
);

FILL FILL_1_CLKBUF1_insert65 (
);

FILL FILL_2__7561_ (
);

FILL FILL_1_CLKBUF1_insert66 (
);

FILL FILL_2__7141_ (
);

FILL FILL_1_CLKBUF1_insert67 (
);

FILL FILL_1_CLKBUF1_insert68 (
);

FILL FILL_1_CLKBUF1_insert69 (
);

FILL FILL_2__11387_ (
);

OAI21X1 _6601_ (
    .A(_199_),
    .B(_200_),
    .C(_198_),
    .Y(_201_)
);

FILL FILL_0__7387_ (
);

INVX1 _9493_ (
    .A(_2848_),
    .Y(_2849_)
);

NAND3X1 _9073_ (
    .A(_2424_),
    .B(_2432_),
    .C(_2434_),
    .Y(_2435_)
);

FILL FILL_1__11741_ (
);

FILL FILL_1__11321_ (
);

FILL FILL_2__8766_ (
);

FILL FILL_2__8346_ (
);

FILL FILL_0__10314_ (
);

OAI22X1 _13071_ (
    .A(_5812_),
    .B(_5814_),
    .C(_5898_),
    .D(_5723_),
    .Y(_6106_)
);

NAND2X1 _7806_ (
    .A(_1316_),
    .B(_1320_),
    .Y(_1321_)
);

FILL FILL_1__6763_ (
);

FILL FILL_2__13113_ (
);

FILL FILL_1__12946_ (
);

FILL FILL_1__12526_ (
);

FILL FILL_1__12106_ (
);

FILL FILL_0__9953_ (
);

FILL FILL_0__9533_ (
);

FILL FILL_0__11939_ (
);

FILL FILL_3__7630_ (
);

FILL FILL_0__9113_ (
);

AND2X2 _11804_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_4924_)
);

FILL FILL_0__11519_ (
);

FILL FILL_1__7968_ (
);

FILL FILL_1__7548_ (
);

FILL FILL_3__10460_ (
);

FILL FILL_1__7128_ (
);

FILL FILL_3__8415_ (
);

NAND3X1 _10196_ (
    .A(_3323_),
    .B(_3462_),
    .C(_3467_),
    .Y(_3475_)
);

FILL FILL_2__6832_ (
);

FILL FILL_2__6412_ (
);

FILL FILL_3__11245_ (
);

FILL FILL_2__10658_ (
);

FILL FILL_0__11692_ (
);

FILL FILL_2__10238_ (
);

FILL FILL_0__11272_ (
);

FILL FILL_0__6658_ (
);

OR2X2 _8764_ (
    .A(_2195_),
    .B(_2188_),
    .Y(_2197_)
);

OAI21X1 _8344_ (
    .A(_1706_),
    .B(_1783_),
    .C(_1700_),
    .Y(_1784_)
);

FILL FILL_2__7617_ (
);

FILL FILL_1__13064_ (
);

FILL FILL_0__12897_ (
);

NAND2X1 _12762_ (
    .A(_5797_),
    .B(_5800_),
    .Y(_5801_)
);

FILL FILL_0__12057_ (
);

INVX1 _12342_ (
    .A(\u_fir_pe6.rYin [5]),
    .Y(_5447_)
);

FILL FILL_2__12804_ (
);

AOI21X1 _9969_ (
    .A(_3228_),
    .B(_3232_),
    .C(_3220_),
    .Y(_3251_)
);

NOR2X1 _9549_ (
    .A(_2884_),
    .B(_2889_),
    .Y(_2904_)
);

AOI22X1 _9129_ (
    .A(vdd),
    .B(\X[3] [4]),
    .C(_2479_),
    .D(_2481_),
    .Y(_2490_)
);

FILL FILL_0__8804_ (
);

FILL FILL_3__6901_ (
);

FILL FILL_3__9373_ (
);

OAI21X1 _13127_ (
    .A(_6158_),
    .B(_6160_),
    .C(_6139_),
    .Y(_6161_)
);

FILL FILL_1__6819_ (
);

FILL FILL_2__7790_ (
);

FILL FILL_2__7370_ (
);

FILL FILL_2__11196_ (
);

NAND2X1 _6830_ (
    .A(_391_),
    .B(_394_),
    .Y(_427_)
);

NAND3X1 _6410_ (
    .A(_10_),
    .B(_12_),
    .C(_11_),
    .Y(_13_)
);

FILL FILL_1__10189_ (
);

FILL FILL_0__7196_ (
);

FILL FILL_3__10936_ (
);

FILL FILL_1__11970_ (
);

FILL FILL_1__11550_ (
);

FILL FILL_1__11130_ (
);

FILL FILL_2__8575_ (
);

FILL FILL_0__10963_ (
);

FILL FILL_2__8155_ (
);

FILL FILL_0__10543_ (
);

FILL FILL_0__10123_ (
);

OAI21X1 _7615_ (
    .A(_1132_),
    .B(_1126_),
    .C(_1120_),
    .Y(_1133_)
);

FILL FILL_1__6992_ (
);

FILL FILL_1__6572_ (
);

FILL FILL_3__6498_ (
);

FILL FILL_1__12755_ (
);

FILL FILL_1__12335_ (
);

FILL FILL_0__9762_ (
);

FILL FILL_0__9342_ (
);

FILL FILL_0__11748_ (
);

DFFPOSX1 _11613_ (
    .D(\Y[5] [5]),
    .CLK(clk_bF$buf57),
    .Q(\u_fir_pe5.rYin [5])
);

FILL FILL_0__11328_ (
);

FILL FILL_1__7777_ (
);

FILL FILL_1__7357_ (
);

FILL FILL_3__8644_ (
);

NAND3X1 _12818_ (
    .A(_5801_),
    .B(_5842_),
    .C(_5847_),
    .Y(_5857_)
);

FILL FILL_2__6641_ (
);

FILL FILL_2__10887_ (
);

FILL FILL_2__10467_ (
);

FILL FILL_2__10047_ (
);

FILL FILL_0__11081_ (
);

FILL FILL_1__9923_ (
);

FILL FILL_1__9503_ (
);

FILL FILL_3__9429_ (
);

FILL FILL_0__6887_ (
);

DFFPOSX1 _8993_ (
    .D(_2385_[0]),
    .CLK(clk_bF$buf36),
    .Q(\u_fir_pe2.mul [0])
);

FILL FILL_0__6467_ (
);

NAND2X1 _8573_ (
    .A(\X[2]_5_bF$buf2 ),
    .B(gnd),
    .Y(_2010_)
);

NAND2X1 _8153_ (
    .A(vdd),
    .B(\X[2] [0]),
    .Y(_1596_)
);

FILL FILL_1__10821_ (
);

FILL FILL_1__10401_ (
);

FILL FILL_2__7846_ (
);

FILL FILL_2__7426_ (
);

FILL FILL_2__7006_ (
);

FILL FILL_1__13293_ (
);

OAI21X1 _12991_ (
    .A(_6026_),
    .B(_6027_),
    .C(_6023_),
    .Y(_6028_)
);

FILL FILL_0__12286_ (
);

INVX1 _12571_ (
    .A(_5612_),
    .Y(_5613_)
);

NAND2X1 _12151_ (
    .A(_5264_),
    .B(_5258_),
    .Y(_5267_)
);

FILL FILL_3__13200_ (
);

FILL FILL_2__12613_ (
);

AND2X2 _9778_ (
    .A(_3120_),
    .B(_3121_),
    .Y(_3181_[10])
);

NAND2X1 _9358_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .Y(_2716_)
);

FILL FILL_0__8613_ (
);

DFFPOSX1 _13356_ (
    .D(\X[6] [2]),
    .CLK(clk_bF$buf2),
    .Q(\X[7] [2])
);

FILL FILL_1__6628_ (
);

FILL FILL_0__9818_ (
);

FILL FILL_3__10325_ (
);

FILL FILL_2__8384_ (
);

FILL FILL_0__10772_ (
);

FILL FILL_0__10352_ (
);

OAI21X1 _7844_ (
    .A(_1102_),
    .B(_1276_),
    .C(_1320_),
    .Y(_1358_)
);

NAND3X1 _7424_ (
    .A(_943_),
    .B(_937_),
    .C(_940_),
    .Y(_944_)
);

OAI22X1 _7004_ (
    .A(_144_),
    .B(_462_),
    .C(_305_),
    .D(_235_),
    .Y(_597_)
);

FILL FILL_1__6381_ (
);

FILL FILL_2__13151_ (
);

FILL FILL_1__12984_ (
);

FILL FILL_1__12564_ (
);

FILL FILL_1__12144_ (
);

FILL FILL_0__9991_ (
);

FILL FILL_0__11977_ (
);

FILL FILL_2__9589_ (
);

FILL FILL_0__9571_ (
);

FILL FILL_2__9169_ (
);

FILL FILL_0__9151_ (
);

AOI21X1 _11842_ (
    .A(_4956_),
    .B(_4957_),
    .C(_4955_),
    .Y(_4962_)
);

FILL FILL_0__11557_ (
);

NAND2X1 _11422_ (
    .A(_4613_),
    .B(_4607_),
    .Y(_4781_[14])
);

FILL FILL_0__11137_ (
);

NAND2X1 _11002_ (
    .A(_4198_),
    .B(_4200_),
    .Y(_4201_)
);

NOR2X1 _8629_ (
    .A(_2000_),
    .B(_1997_),
    .Y(_2065_)
);

OR2X2 _8209_ (
    .A(_1650_),
    .B(_1649_),
    .Y(_1651_)
);

FILL FILL_1__7586_ (
);

FILL FILL_1__7166_ (
);

FILL FILL_3__8873_ (
);

INVX1 _12627_ (
    .A(vdd),
    .Y(_5668_)
);

NAND2X1 _12207_ (
    .A(_5314_),
    .B(_5317_),
    .Y(_5322_)
);

FILL FILL_2__6870_ (
);

FILL FILL_2__6450_ (
);

FILL FILL_3__11283_ (
);

FILL FILL_2__10696_ (
);

FILL FILL_2__10276_ (
);

FILL FILL_1__9732_ (
);

FILL FILL_1__9312_ (
);

FILL FILL_0__6696_ (
);

AND2X2 _8382_ (
    .A(\X[2] [3]),
    .B(vdd),
    .Y(_1821_)
);

FILL FILL_1__10630_ (
);

FILL FILL_1__10210_ (
);

FILL FILL_2__7655_ (
);

FILL FILL_3__12068_ (
);

FILL FILL_0__12095_ (
);

NAND3X1 _12380_ (
    .A(_5483_),
    .B(_5480_),
    .C(_5443_),
    .Y(_5484_)
);

FILL FILL_2__12842_ (
);

FILL FILL_2__12422_ (
);

FILL FILL_2__12002_ (
);

NAND3X1 _9587_ (
    .A(_2933_),
    .B(_2937_),
    .C(_2941_),
    .Y(_2942_)
);

NAND2X1 _9167_ (
    .A(_2526_),
    .B(_2525_),
    .Y(_2527_)
);

FILL FILL_1__11835_ (
);

FILL FILL_1__11415_ (
);

FILL FILL_0__8842_ (
);

FILL FILL_0__8422_ (
);

FILL FILL_0__10828_ (
);

FILL FILL_0__10408_ (
);

FILL FILL_0__8002_ (
);

AND2X2 _13165_ (
    .A(_6175_),
    .B(_6174_),
    .Y(_6197_)
);

FILL FILL_2__9801_ (
);

FILL FILL_1__6857_ (
);

FILL FILL_1__6437_ (
);

FILL FILL_2__13207_ (
);

FILL FILL_0__9627_ (
);

FILL FILL_3__7724_ (
);

FILL FILL_0__9207_ (
);

FILL FILL_3__7304_ (
);

FILL FILL_3__10554_ (
);

FILL FILL_2__8193_ (
);

FILL FILL_0__10581_ (
);

FILL FILL_0__10161_ (
);

FILL FILL_3__8509_ (
);

NAND2X1 _7653_ (
    .A(_1170_),
    .B(_1094_),
    .Y(_1171_)
);

DFFPOSX1 _7233_ (
    .D(Yin[10]),
    .CLK(clk_bF$buf1),
    .Q(\u_fir_pe0.rYin [10])
);

FILL FILL_2__6926_ (
);

FILL FILL_2__6506_ (
);

FILL FILL_1__12793_ (
);

FILL FILL_3__11339_ (
);

FILL FILL_1__12373_ (
);

FILL FILL_0__9380_ (
);

FILL FILL_2__9398_ (
);

FILL FILL_0__11786_ (
);

NAND2X1 _11651_ (
    .A(_5562_),
    .B(_5542_),
    .Y(_5563_)
);

FILL FILL_0__11366_ (
);

INVX1 _11231_ (
    .A(_4349_),
    .Y(_4428_)
);

FILL FILL_3__12700_ (
);

NOR2X1 _8858_ (
    .A(_2278_),
    .B(_2277_),
    .Y(_2281_)
);

OAI21X1 _8438_ (
    .A(_1863_),
    .B(_1867_),
    .C(_1870_),
    .Y(_1877_)
);

INVX1 _8018_ (
    .A(\u_fir_pe1.mul [10]),
    .Y(_1522_)
);

FILL FILL_1__7395_ (
);

FILL FILL_1__13158_ (
);

NAND2X1 _12856_ (
    .A(_5889_),
    .B(_5893_),
    .Y(_5894_)
);

FILL FILL_3__8262_ (
);

AND2X2 _12436_ (
    .A(_5539_),
    .B(_5538_),
    .Y(_5572_[13])
);

AOI21X1 _12016_ (
    .A(_5133_),
    .B(_5128_),
    .C(_5097_),
    .Y(_5134_)
);

FILL FILL_2__10085_ (
);

FILL FILL_1__9961_ (
);

FILL FILL_1__9541_ (
);

FILL FILL_1__9121_ (
);

FILL FILL_3__9887_ (
);

FILL FILL_3__9467_ (
);

FILL FILL_3__9047_ (
);

INVX1 _8191_ (
    .A(_1632_),
    .Y(_1633_)
);

FILL FILL_2__7884_ (
);

FILL FILL_2__7464_ (
);

FILL FILL_3__12297_ (
);

FILL FILL_2__7044_ (
);

OAI22X1 _6924_ (
    .A(_417_),
    .B(_462_),
    .C(_518_),
    .D(_517_),
    .Y(_519_)
);

NAND3X1 _6504_ (
    .A(_102_),
    .B(_104_),
    .C(_103_),
    .Y(_105_)
);

FILL FILL_2__12651_ (
);

FILL FILL_2__12231_ (
);

AOI21X1 _9396_ (
    .A(_2748_),
    .B(_2753_),
    .C(_2692_),
    .Y(_2754_)
);

FILL FILL_1__11644_ (
);

FILL FILL_1__11224_ (
);

FILL FILL_0__8651_ (
);

FILL FILL_2__8669_ (
);

FILL FILL_0__8231_ (
);

FILL FILL_2__8249_ (
);

FILL FILL_0__10637_ (
);

AOI21X1 _10922_ (
    .A(_4076_),
    .B(_4080_),
    .C(_4069_),
    .Y(_4122_)
);

OAI21X1 _10502_ (
    .A(_3564_),
    .B(_3775_),
    .C(_3747_),
    .Y(_3776_)
);

FILL FILL_0__10217_ (
);

BUFX2 _13394_ (
    .A(_6376_[0]),
    .Y(Xout[0])
);

FILL FILL_2__9610_ (
);

AOI21X1 _7709_ (
    .A(_1212_),
    .B(_1219_),
    .C(_1194_),
    .Y(_1226_)
);

FILL FILL_1__6666_ (
);

FILL FILL_2__13016_ (
);

FILL FILL_1__12849_ (
);

FILL FILL_1__12429_ (
);

FILL FILL_1__12009_ (
);

FILL FILL_3__7953_ (
);

FILL FILL_0__9436_ (
);

FILL FILL_0__9016_ (
);

NAND2X1 _11707_ (
    .A(_4826_),
    .B(_4822_),
    .Y(_4829_)
);

FILL FILL_3__7113_ (
);

FILL FILL_3__10783_ (
);

FILL FILL_0__10390_ (
);

FILL FILL_1__8812_ (
);

FILL FILL_3__8738_ (
);

NAND2X1 _7882_ (
    .A(_1394_),
    .B(_1393_),
    .Y(_1395_)
);

OAI21X1 _7462_ (
    .A(_977_),
    .B(_978_),
    .C(_935_),
    .Y(_982_)
);

AND2X2 _7042_ (
    .A(\u_fir_pe0.rYin [0]),
    .B(\u_fir_pe0.mul [0]),
    .Y(_631_)
);

NAND3X1 _10099_ (
    .A(_3372_),
    .B(_3365_),
    .C(_3370_),
    .Y(_3379_)
);

FILL FILL_2__6735_ (
);

FILL FILL_3__11568_ (
);

FILL FILL_1__12182_ (
);

NAND3X1 _11880_ (
    .A(_4925_),
    .B(_4994_),
    .C(_4929_),
    .Y(_4999_)
);

OAI21X1 _11460_ (
    .A(_4636_),
    .B(_4632_),
    .C(_4645_),
    .Y(_4646_)
);

FILL FILL_0__11175_ (
);

NAND2X1 _11040_ (
    .A(gnd),
    .B(\X[5]_5_bF$buf0 ),
    .Y(_4239_)
);

FILL FILL_2__11922_ (
);

FILL FILL_2__11502_ (
);

OAI21X1 _8667_ (
    .A(_2102_),
    .B(_1970_),
    .C(_2052_),
    .Y(_2103_)
);

NAND3X1 _8247_ (
    .A(vdd),
    .B(\X[2] [2]),
    .C(_1687_),
    .Y(_1688_)
);

FILL FILL_1__10915_ (
);

FILL FILL_0__7922_ (
);

FILL FILL_0__7502_ (
);

FILL FILL_3__8491_ (
);

INVX1 _12665_ (
    .A(_5646_),
    .Y(_5706_)
);

FILL FILL_3__8071_ (
);

NAND2X1 _12245_ (
    .A(_5345_),
    .B(_5358_),
    .Y(_5359_)
);

FILL FILL_2__12707_ (
);

FILL FILL_0__13321_ (
);

FILL FILL_0__8707_ (
);

FILL FILL_1__9770_ (
);

FILL FILL_1__9350_ (
);

FILL FILL_3__9696_ (
);

FILL FILL_3__9276_ (
);

FILL FILL_2__7693_ (
);

FILL FILL_2__7273_ (
);

FILL FILL_2__11099_ (
);

AND2X2 _6733_ (
    .A(vdd),
    .B(Xin[6]),
    .Y(_331_)
);

FILL FILL_2__12880_ (
);

FILL FILL_2__12460_ (
);

FILL FILL_2__12040_ (
);

FILL FILL_0__7099_ (
);

FILL FILL_3__10839_ (
);

FILL FILL_1__11873_ (
);

FILL FILL_3__10419_ (
);

FILL FILL_1__11453_ (
);

FILL FILL_1__11033_ (
);

FILL FILL_0__8880_ (
);

FILL FILL_2__8898_ (
);

FILL FILL_2__8478_ (
);

FILL FILL_0__8460_ (
);

FILL FILL_0__10866_ (
);

DFFPOSX1 _10731_ (
    .D(\Y[4] [0]),
    .CLK(clk_bF$buf26),
    .Q(\u_fir_pe4.rYin [0])
);

FILL FILL_0__10446_ (
);

FILL FILL_2__8058_ (
);

FILL FILL_0__8040_ (
);

NOR2X1 _10311_ (
    .A(_3586_),
    .B(_3587_),
    .Y(_3588_)
);

FILL FILL_0__10026_ (
);

INVX1 _7938_ (
    .A(\u_fir_pe1.rYin [3]),
    .Y(_1445_)
);

NAND2X1 _7518_ (
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_1037_)
);

FILL FILL_1__6895_ (
);

FILL FILL_1__6475_ (
);

FILL FILL_2__13245_ (
);

FILL FILL_3_CLKBUF1_insert12 (
);

FILL FILL_3_CLKBUF1_insert13 (
);

FILL FILL_1__12658_ (
);

FILL FILL_3_CLKBUF1_insert15 (
);

FILL FILL_1__12238_ (
);

FILL FILL_3_CLKBUF1_insert17 (
);

FILL FILL_3_CLKBUF1_insert19 (
);

FILL FILL_0__9665_ (
);

FILL FILL_0__9245_ (
);

AOI21X1 _11936_ (
    .A(_5054_),
    .B(_5053_),
    .C(_5052_),
    .Y(_5055_)
);

FILL FILL_3__7342_ (
);

INVX1 _11516_ (
    .A(_4699_),
    .Y(_4700_)
);

FILL FILL_3__10172_ (
);

FILL FILL_1__8621_ (
);

FILL FILL_1__8201_ (
);

NAND2X1 _7691_ (
    .A(_1198_),
    .B(_1207_),
    .Y(_1208_)
);

INVX1 _7271_ (
    .A(_1582_),
    .Y(_1583_)
);

FILL FILL_2__6964_ (
);

FILL FILL_3__11797_ (
);

FILL FILL_2__6544_ (
);

FILL FILL_3__11377_ (
);

FILL FILL_1__9826_ (
);

FILL FILL_1__9406_ (
);

FILL FILL_2__11731_ (
);

FILL FILL_2__11311_ (
);

NOR2X1 _8896_ (
    .A(_2318_),
    .B(_2319_),
    .Y(_2320_)
);

OAI21X1 _8476_ (
    .A(_1609_),
    .B(_1913_),
    .C(_1619_),
    .Y(_1914_)
);

NOR2X1 _8056_ (
    .A(\u_fir_pe1.rYin [14]),
    .B(\u_fir_pe1.mul [14]),
    .Y(_1560_)
);

FILL FILL_1__10304_ (
);

FILL FILL_0__7731_ (
);

FILL FILL_2__7749_ (
);

FILL FILL_2__7329_ (
);

FILL FILL_0__7311_ (
);

FILL FILL_1__13196_ (
);

AND2X2 _12894_ (
    .A(_5893_),
    .B(_5889_),
    .Y(_5932_)
);

FILL FILL_0__12189_ (
);

DFFPOSX1 _12474_ (
    .D(_5572_[13]),
    .CLK(clk_bF$buf8),
    .Q(_6377_[13])
);

INVX1 _12054_ (
    .A(_5170_),
    .Y(_5171_)
);

FILL FILL_2__12936_ (
);

FILL FILL_0__13130_ (
);

FILL FILL_1__11929_ (
);

FILL FILL_1__11509_ (
);

FILL FILL_0__8936_ (
);

FILL FILL_0__8516_ (
);

FILL FILL_3__6613_ (
);

FILL FILL_3__9085_ (
);

OAI21X1 _13259_ (
    .A(_6271_),
    .B(_6272_),
    .C(_6282_),
    .Y(_6283_)
);

FILL FILL_2__7082_ (
);

FILL FILL_3__7818_ (
);

NOR3X1 _6962_ (
    .A(_502_),
    .B(_504_),
    .C(_552_),
    .Y(_556_)
);

AND2X2 _6542_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_142_)
);

FILL FILL_3__10648_ (
);

FILL FILL_1__11682_ (
);

FILL FILL_1__11262_ (
);

FILL FILL_2__8287_ (
);

FILL FILL_0__10675_ (
);

NAND3X1 _10960_ (
    .A(_4147_),
    .B(_4151_),
    .C(_4153_),
    .Y(_4160_)
);

NOR3X1 _10540_ (
    .A(_3811_),
    .B(_3779_),
    .C(_3797_),
    .Y(_3812_)
);

FILL FILL_0__10255_ (
);

INVX1 _10120_ (
    .A(_3398_),
    .Y(_3399_)
);

OAI22X1 _7747_ (
    .A(_812_),
    .B(_1259_),
    .C(_1260_),
    .D(_1262_),
    .Y(_1263_)
);

NAND3X1 _7327_ (
    .A(_825_),
    .B(_848_),
    .C(_847_),
    .Y(_849_)
);

FILL FILL_2__13054_ (
);

FILL FILL_1__12887_ (
);

FILL FILL_1__12047_ (
);

FILL FILL_0__9894_ (
);

FILL FILL_0__9474_ (
);

FILL FILL_3__7571_ (
);

FILL FILL_0__9054_ (
);

OAI22X1 _11745_ (
    .A(_5513_),
    .B(_4865_),
    .C(_4815_),
    .D(_4820_),
    .Y(_4866_)
);

NAND3X1 _11325_ (
    .A(_4514_),
    .B(_4519_),
    .C(_4518_),
    .Y(_4520_)
);

FILL FILL_0__12821_ (
);

FILL FILL_0__12401_ (
);

FILL FILL_1__7489_ (
);

FILL FILL_1__7069_ (
);

FILL FILL_1__8850_ (
);

FILL FILL_1__8430_ (
);

FILL FILL_1__8010_ (
);

FILL FILL_3__8356_ (
);

INVX1 _7080_ (
    .A(\u_fir_pe0.rYin [5]),
    .Y(_665_)
);

FILL FILL_2__6773_ (
);

FILL FILL_3__11186_ (
);

FILL FILL_2__10599_ (
);

FILL FILL_2__10179_ (
);

FILL FILL_1__9635_ (
);

FILL FILL_1__9215_ (
);

FILL FILL_2__11960_ (
);

FILL FILL_2__11540_ (
);

FILL FILL_2__11120_ (
);

FILL FILL_0__6599_ (
);

AND2X2 _8285_ (
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1725_)
);

FILL FILL_1__10953_ (
);

FILL FILL_1__10533_ (
);

FILL FILL_1__10113_ (
);

FILL FILL_0__7960_ (
);

FILL FILL_2__7978_ (
);

FILL FILL_2__7558_ (
);

FILL FILL_0__7540_ (
);

FILL FILL_2__7138_ (
);

FILL FILL_0__7120_ (
);

NAND2X1 _12283_ (
    .A(_5395_),
    .B(_5392_),
    .Y(_5578_[13])
);

FILL FILL_2__12745_ (
);

FILL FILL_2__12325_ (
);

FILL FILL_1__11738_ (
);

FILL FILL_1__11318_ (
);

FILL FILL_0__8745_ (
);

FILL FILL_3__6842_ (
);

FILL FILL_0__8325_ (
);

NAND2X1 _13068_ (
    .A(_6098_),
    .B(_6102_),
    .Y(_6103_)
);

FILL FILL_2__9704_ (
);

FILL FILL_1__7701_ (
);

OAI21X1 _6771_ (
    .A(_135_),
    .B(_368_),
    .C(_282_),
    .Y(_369_)
);

FILL FILL_3__10877_ (
);

FILL FILL_1__11491_ (
);

FILL FILL_3__10037_ (
);

FILL FILL_1__11071_ (
);

FILL FILL_0__10484_ (
);

FILL FILL_0__10064_ (
);

FILL FILL_1__8906_ (
);

FILL FILL_2__10811_ (
);

INVX1 _7976_ (
    .A(\u_fir_pe1.mul [7]),
    .Y(_1479_)
);

NAND3X1 _7556_ (
    .A(_1019_),
    .B(_1060_),
    .C(_1065_),
    .Y(_1075_)
);

AOI21X1 _7136_ (
    .A(_714_),
    .B(_692_),
    .C(_712_),
    .Y(_719_)
);

FILL FILL_2__13283_ (
);

FILL FILL_0__6811_ (
);

FILL FILL_2__6829_ (
);

FILL FILL_2__6409_ (
);

FILL FILL_1__12696_ (
);

FILL FILL_1__12276_ (
);

FILL FILL_0__9283_ (
);

OAI21X1 _11974_ (
    .A(_5090_),
    .B(_5091_),
    .C(_5086_),
    .Y(_5092_)
);

FILL FILL_0__11689_ (
);

NOR2X1 _11554_ (
    .A(_4736_),
    .B(_4737_),
    .Y(_4738_)
);

FILL FILL_0__11269_ (
);

INVX1 _11134_ (
    .A(_4245_),
    .Y(_4332_)
);

FILL FILL_0__12630_ (
);

FILL FILL_0__12210_ (
);

FILL FILL_1__7298_ (
);

NOR2X1 _9702_ (
    .A(_3046_),
    .B(_3047_),
    .Y(_3048_)
);

FILL FILL_3__8585_ (
);

AOI21X1 _12759_ (
    .A(_5726_),
    .B(_5722_),
    .C(_5791_),
    .Y(_5798_)
);

OR2X2 _12339_ (
    .A(_5443_),
    .B(_5441_),
    .Y(_5445_)
);

FILL FILL_0__13415_ (
);

FILL FILL_2__6582_ (
);

FILL FILL_1__9444_ (
);

FILL FILL_1__9024_ (
);

DFFPOSX1 _8094_ (
    .D(\X[1] [2]),
    .CLK(clk_bF$buf54),
    .Q(\X[2] [2])
);

FILL FILL_1__10342_ (
);

FILL FILL_2__7787_ (
);

FILL FILL_2__7367_ (
);

NAND2X1 _12092_ (
    .A(_5173_),
    .B(_5176_),
    .Y(_5209_)
);

FILL FILL_3__13141_ (
);

NAND2X1 _6827_ (
    .A(_415_),
    .B(_422_),
    .Y(_424_)
);

INVX1 _6407_ (
    .A(_740_),
    .Y(_10_)
);

FILL FILL_2__12974_ (
);

FILL FILL_2__12554_ (
);

FILL FILL_2__12134_ (
);

NAND3X1 _9299_ (
    .A(_2629_),
    .B(_2648_),
    .C(_2642_),
    .Y(_2658_)
);

FILL FILL_1__11967_ (
);

FILL FILL_1__11547_ (
);

FILL FILL_1__11127_ (
);

FILL FILL_0__8554_ (
);

FILL FILL_0__8134_ (
);

NAND2X1 _10825_ (
    .A(gnd),
    .B(\X[5] [2]),
    .Y(_4027_)
);

NAND2X1 _10405_ (
    .A(_3679_),
    .B(_3675_),
    .Y(_3681_)
);

INVX1 _13297_ (
    .A(\u_fir_pe7.rYin [12]),
    .Y(_6321_)
);

FILL FILL_2__9933_ (
);

FILL FILL_0__11901_ (
);

FILL FILL_2__9513_ (
);

FILL FILL_1__6989_ (
);

FILL FILL_1__6569_ (
);

FILL FILL_1__7930_ (
);

FILL FILL_1__7510_ (
);

FILL FILL_0__9759_ (
);

FILL FILL_0__9339_ (
);

FILL FILL_3__7436_ (
);

AOI21X1 _6580_ (
    .A(_174_),
    .B(_175_),
    .C(_173_),
    .Y(_180_)
);

FILL FILL_3__10266_ (
);

FILL FILL_0__10293_ (
);

FILL FILL_1__8715_ (
);

FILL FILL_2__10620_ (
);

FILL FILL_2__10200_ (
);

AOI21X1 _7785_ (
    .A(_1228_),
    .B(_1234_),
    .C(_1300_),
    .Y(_1301_)
);

INVX1 _7365_ (
    .A(vdd),
    .Y(_886_)
);

FILL FILL_2__13092_ (
);

FILL FILL_2__6638_ (
);

FILL FILL_0__6620_ (
);

FILL FILL_1__12085_ (
);

FILL FILL_0__9092_ (
);

NAND3X1 _11783_ (
    .A(_4903_),
    .B(_4836_),
    .C(_4839_),
    .Y(_4904_)
);

FILL FILL_0__11498_ (
);

FILL FILL_0__11078_ (
);

NAND3X1 _11363_ (
    .A(_4549_),
    .B(_4556_),
    .C(_4555_),
    .Y(_4557_)
);

FILL FILL_2__11825_ (
);

FILL FILL_2__11405_ (
);

FILL FILL_1__10818_ (
);

FILL FILL_0__7825_ (
);

NAND2X1 _9931_ (
    .A(\X[4] [4]),
    .B(gnd),
    .Y(_3213_)
);

FILL FILL_0__7405_ (
);

OAI22X1 _9511_ (
    .A(_2722_),
    .B(_2803_),
    .C(_2865_),
    .D(_2866_),
    .Y(_2867_)
);

NAND3X1 _12988_ (
    .A(_6005_),
    .B(_6009_),
    .C(_6012_),
    .Y(_6025_)
);

NAND2X1 _12568_ (
    .A(vdd),
    .B(\X[6] [1]),
    .Y(_5610_)
);

NAND3X1 _12148_ (
    .A(_5262_),
    .B(_5263_),
    .C(_5261_),
    .Y(_5264_)
);

FILL FILL_0__13224_ (
);

FILL FILL_2__6391_ (
);

FILL FILL_3__6707_ (
);

FILL FILL_1__9673_ (
);

FILL FILL_1__9253_ (
);

FILL FILL253950x244950 (
);

FILL FILL_1__10991_ (
);

FILL FILL_1__10571_ (
);

FILL FILL_1__10151_ (
);

FILL FILL_2__7596_ (
);

FILL FILL_2__7176_ (
);

INVX1 _6636_ (
    .A(Xin[7]),
    .Y(_235_)
);

FILL FILL_2__12783_ (
);

FILL FILL_2__12363_ (
);

FILL FILL_1__11776_ (
);

FILL FILL_1__11356_ (
);

FILL FILL_0__8783_ (
);

FILL FILL_3__6880_ (
);

FILL FILL_0__8363_ (
);

FILL FILL_0__10769_ (
);

FILL FILL_3__6460_ (
);

FILL FILL_0__10349_ (
);

INVX1 _10634_ (
    .A(_3893_),
    .Y(_3897_)
);

NAND2X1 _10214_ (
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3492_)
);

FILL FILL_2__9742_ (
);

FILL FILL_2__9322_ (
);

FILL FILL_0__11710_ (
);

FILL FILL_1__6798_ (
);

FILL FILL_1__6378_ (
);

FILL FILL_2__13148_ (
);

FILL FILL_0__9988_ (
);

FILL FILL_0__9568_ (
);

FILL FILL_3__7665_ (
);

FILL FILL_0__9148_ (
);

NAND3X1 _11839_ (
    .A(_4954_),
    .B(_4920_),
    .C(_4958_),
    .Y(_4959_)
);

INVX1 _11419_ (
    .A(_4601_),
    .Y(_4611_)
);

FILL FILL_0__12915_ (
);

FILL FILL_3__10495_ (
);

FILL FILL_1__8944_ (
);

FILL FILL_1__8524_ (
);

NAND2X1 _7594_ (
    .A(_1107_),
    .B(_1111_),
    .Y(_1112_)
);

AND2X2 _7174_ (
    .A(_757_),
    .B(_756_),
    .Y(_790_[13])
);

FILL FILL_3__9811_ (
);

FILL FILL_2__6867_ (
);

FILL FILL_2__6447_ (
);

DFFPOSX1 _11592_ (
    .D(_4775_[8]),
    .CLK(clk_bF$buf5),
    .Q(\Y[6] [8])
);

AOI21X1 _11172_ (
    .A(_4334_),
    .B(_4335_),
    .C(_4302_),
    .Y(_4369_)
);

FILL FILL_1__9729_ (
);

FILL FILL_1__9309_ (
);

FILL FILL_3__12641_ (
);

FILL FILL_3__12221_ (
);

FILL FILL_2__11214_ (
);

FILL FILL254250x154950 (
);

NOR2X1 _8799_ (
    .A(_2226_),
    .B(_2227_),
    .Y(_2228_)
);

OAI21X1 _8379_ (
    .A(_1767_),
    .B(_1817_),
    .C(_1761_),
    .Y(_1818_)
);

FILL FILL_1__10627_ (
);

FILL FILL_1__10207_ (
);

FILL FILL_0__7634_ (
);

NOR2X1 _9740_ (
    .A(_3081_),
    .B(_3082_),
    .Y(_3083_)
);

NAND3X1 _9320_ (
    .A(_2579_),
    .B(_2677_),
    .C(_2678_),
    .Y(_2679_)
);

FILL FILL_1__13099_ (
);

NAND3X1 _12797_ (
    .A(_5832_),
    .B(_5831_),
    .C(_5835_),
    .Y(_5836_)
);

AND2X2 _12377_ (
    .A(_5459_),
    .B(_5469_),
    .Y(_5480_)
);

FILL FILL_3__13006_ (
);

FILL FILL_2__12839_ (
);

FILL FILL253950x93750 (
);

FILL FILL_2__12419_ (
);

FILL FILL_0__13033_ (
);

FILL FILL_0__8839_ (
);

FILL FILL_3__6936_ (
);

FILL FILL_0__8419_ (
);

FILL FILL_1__9482_ (
);

FILL FILL_1__9062_ (
);

FILL FILL_1__10380_ (
);

OAI21X1 _6865_ (
    .A(_427_),
    .B(_429_),
    .C(_423_),
    .Y(_461_)
);

NAND2X1 _6445_ (
    .A(_44_),
    .B(_40_),
    .Y(_47_)
);

FILL FILL_2__12592_ (
);

FILL FILL_2__12172_ (
);

FILL FILL_1__11165_ (
);

FILL FILL_0__8592_ (
);

FILL FILL_0__10998_ (
);

FILL FILL_0__8172_ (
);

FILL FILL_0__10578_ (
);

NAND2X1 _10863_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf2 ),
    .Y(_4064_)
);

INVX1 _10443_ (
    .A(_3717_),
    .Y(_3718_)
);

FILL FILL_0__10158_ (
);

NAND3X1 _10023_ (
    .A(_3241_),
    .B(_3299_),
    .C(_3303_),
    .Y(_3304_)
);

FILL FILL_2__10905_ (
);

FILL FILL_2__9971_ (
);

FILL FILL_2__9551_ (
);

FILL FILL_2__9131_ (
);

FILL FILL_0__6905_ (
);

FILL FILL_0__9797_ (
);

FILL FILL_3__7894_ (
);

FILL FILL_0__9377_ (
);

INVX1 _11648_ (
    .A(\X[7] [2]),
    .Y(_5552_)
);

FILL FILL_3__7054_ (
);

AOI21X1 _11228_ (
    .A(_4415_),
    .B(_4411_),
    .C(_4370_),
    .Y(_4425_)
);

FILL FILL_1__13311_ (
);

FILL FILL_0__12724_ (
);

FILL FILL_0__12304_ (
);

FILL FILL_1__8753_ (
);

FILL FILL_1__8333_ (
);

FILL FILL_3__8679_ (
);

FILL FILL_3__9200_ (
);

FILL FILL_2__6676_ (
);

FILL FILL_1__9958_ (
);

FILL FILL_3__12870_ (
);

FILL FILL_1__9538_ (
);

FILL FILL_1__9118_ (
);

FILL FILL_3__12450_ (
);

FILL FILL_3__12030_ (
);

FILL FILL_2__11863_ (
);

FILL FILL_2__11443_ (
);

FILL FILL_2__11023_ (
);

AND2X2 _8188_ (
    .A(vdd),
    .B(\X[2] [2]),
    .Y(_1630_)
);

FILL FILL_1__10856_ (
);

FILL FILL_1__10436_ (
);

FILL FILL_1__10016_ (
);

FILL FILL_0__7863_ (
);

FILL FILL_0__7443_ (
);

FILL FILL_0__7023_ (
);

OAI22X1 _12186_ (
    .A(_5199_),
    .B(_5244_),
    .C(_5300_),
    .D(_5299_),
    .Y(_5301_)
);

FILL FILL_2__8822_ (
);

FILL FILL_2__8402_ (
);

FILL FILL_3__13235_ (
);

FILL FILL_2__12648_ (
);

FILL FILL_2__12228_ (
);

FILL FILL_0__13262_ (
);

FILL FILL_0__8648_ (
);

FILL FILL_0__8228_ (
);

OR2X2 _10919_ (
    .A(_4118_),
    .B(_4116_),
    .Y(_4119_)
);

FILL FILL_1__9291_ (
);

FILL FILL_2_CLKBUF1_insert20 (
);

FILL FILL_2_CLKBUF1_insert21 (
);

FILL FILL_2__9607_ (
);

FILL FILL_2_CLKBUF1_insert22 (
);

FILL FILL_2_CLKBUF1_insert23 (
);

FILL FILL_2_CLKBUF1_insert24 (
);

FILL FILL_2_CLKBUF1_insert25 (
);

FILL FILL_2_CLKBUF1_insert26 (
);

FILL FILL_2_CLKBUF1_insert27 (
);

FILL FILL_2_CLKBUF1_insert28 (
);

FILL FILL_2_CLKBUF1_insert29 (
);

FILL FILL_1__7604_ (
);

AOI21X1 _6674_ (
    .A(_272_),
    .B(_271_),
    .C(_270_),
    .Y(_273_)
);

FILL FILL_1__11394_ (
);

FILL FILL_0__10387_ (
);

OR2X2 _10672_ (
    .A(_3929_),
    .B(_3934_),
    .Y(_3936_)
);

FILL FILL253650x230550 (
);

INVX1 _10252_ (
    .A(_3510_),
    .Y(_3530_)
);

FILL FILL_1__8809_ (
);

FILL FILL_3__11721_ (
);

FILL FILL_2__9780_ (
);

FILL FILL_2__9360_ (
);

NOR2X1 _7879_ (
    .A(_1032_),
    .B(_1259_),
    .Y(_1392_)
);

OAI21X1 _7459_ (
    .A(_977_),
    .B(_978_),
    .C(_976_),
    .Y(_979_)
);

OAI21X1 _7039_ (
    .A(_567_),
    .B(_617_),
    .C(_595_),
    .Y(_630_)
);

FILL FILL_2__13186_ (
);

FILL FILL_0__6714_ (
);

NAND2X1 _8820_ (
    .A(_2246_),
    .B(_2241_),
    .Y(_2247_)
);

FILL FILL_1__12599_ (
);

AOI21X1 _8400_ (
    .A(_1838_),
    .B(_1837_),
    .C(_1834_),
    .Y(_1839_)
);

FILL FILL_1__12179_ (
);

FILL FILL_0__9186_ (
);

AND2X2 _11877_ (
    .A(_4927_),
    .B(_4931_),
    .Y(_4996_)
);

FILL FILL_3__7283_ (
);

NOR2X1 _11457_ (
    .A(\u_fir_pe5.rYin [4]),
    .B(\u_fir_pe5.mul [4]),
    .Y(_4643_)
);

OAI21X1 _11037_ (
    .A(_4235_),
    .B(_4230_),
    .C(_4224_),
    .Y(_4236_)
);

FILL FILL_1__13120_ (
);

FILL FILL_2__11919_ (
);

FILL FILL_0__12953_ (
);

FILL FILL_0__12533_ (
);

FILL FILL_0__12113_ (
);

FILL FILL_0__7919_ (
);

NOR2X1 _9605_ (
    .A(_2958_),
    .B(_2957_),
    .Y(_2959_)
);

FILL FILL_1__8562_ (
);

FILL FILL_1__8142_ (
);

FILL FILL_0__13318_ (
);

FILL FILL_2__6485_ (
);

FILL FILL_1__9767_ (
);

FILL FILL_1__9347_ (
);

FILL FILL_2__11672_ (
);

FILL FILL_2__11252_ (
);

FILL FILL_1__10665_ (
);

FILL FILL_1__10245_ (
);

FILL FILL_0__7672_ (
);

FILL FILL_2__8631_ (
);

FILL FILL_2__8211_ (
);

FILL FILL_2__12877_ (
);

FILL FILL_2__12457_ (
);

FILL FILL_2__12037_ (
);

FILL FILL_0__13071_ (
);

FILL FILL_0__8877_ (
);

FILL FILL_3__6974_ (
);

FILL FILL_0__8457_ (
);

FILL FILL_3__6554_ (
);

DFFPOSX1 _10728_ (
    .D(\X[4]_5_bF$buf1 ),
    .CLK(clk_bF$buf21),
    .Q(\X[5] [5])
);

FILL FILL_0__8037_ (
);

OAI21X1 _10308_ (
    .A(_3510_),
    .B(_3584_),
    .C(_3531_),
    .Y(_3585_)
);

FILL FILL_1__12811_ (
);

FILL FILL_2__9416_ (
);

FILL FILL_0__11804_ (
);

FILL FILL_1__7833_ (
);

FILL FILL_1__7413_ (
);

FILL FILL_3__7759_ (
);

FILL FILL_3__7339_ (
);

OAI22X1 _6483_ (
    .A(_731_),
    .B(_83_),
    .C(_33_),
    .D(_38_),
    .Y(_84_)
);

FILL FILL_3__10589_ (
);

FILL FILL254550x133350 (
);

NOR2X1 _10481_ (
    .A(_3332_),
    .B(_3493_),
    .Y(_3755_)
);

FILL FILL_0__10196_ (
);

NAND2X1 _10061_ (
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3341_)
);

FILL FILL_1__8618_ (
);

FILL FILL_3__11950_ (
);

FILL FILL_3__11110_ (
);

FILL FILL_2__10943_ (
);

FILL FILL_2__10523_ (
);

FILL FILL_2__10103_ (
);

AND2X2 _7688_ (
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1205_)
);

NOR2X1 _7268_ (
    .A(_1577_),
    .B(_1557_),
    .Y(_1580_)
);

FILL FILL_3__9905_ (
);

FILL FILL_0__6943_ (
);

FILL FILL_0__6523_ (
);

NOR2X1 _11686_ (
    .A(_4806_),
    .B(_4807_),
    .Y(_4808_)
);

AND2X2 _11266_ (
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4462_)
);

FILL FILL_2__7902_ (
);

FILL FILL_3__12735_ (
);

FILL FILL_2__11728_ (
);

FILL FILL_0__12762_ (
);

FILL FILL_2__11308_ (
);

FILL FILL_0__12342_ (
);

FILL FILL_0__7728_ (
);

DFFPOSX1 _9834_ (
    .D(_3181_[4]),
    .CLK(clk_bF$buf38),
    .Q(\Y[4] [4])
);

FILL FILL_0__7308_ (
);

AOI21X1 _9414_ (
    .A(_2688_),
    .B(_2758_),
    .C(_2770_),
    .Y(_2771_)
);

FILL FILL_1__8791_ (
);

FILL FILL_1__8371_ (
);

FILL FILL_3__8297_ (
);

BUFX2 _13412_ (
    .A(_6377_[4]),
    .Y(Yout[4])
);

FILL FILL_0__13127_ (
);

FILL FILL_1__9996_ (
);

FILL FILL_1__9576_ (
);

FILL FILL_1__9156_ (
);

FILL FILL_2__11481_ (
);

FILL FILL_2__11061_ (
);

FILL FILL_1__10894_ (
);

FILL FILL_1__10474_ (
);

FILL FILL_1__10054_ (
);

FILL FILL_0__7481_ (
);

FILL FILL_2__7499_ (
);

FILL FILL_0__7061_ (
);

FILL FILL_2__7079_ (
);

FILL FILL_2__8860_ (
);

FILL FILL_2__8440_ (
);

FILL FILL_2__8020_ (
);

NAND3X1 _6959_ (
    .A(_511_),
    .B(_553_),
    .C(_512_),
    .Y(_554_)
);

NAND2X1 _6539_ (
    .A(Xin[1]),
    .B(gnd),
    .Y(_139_)
);

FILL FILL_2__12686_ (
);

FILL FILL_2__12266_ (
);

AOI21X1 _7900_ (
    .A(_1354_),
    .B(_1356_),
    .C(_1411_),
    .Y(_1412_)
);

FILL FILL_1__11679_ (
);

FILL FILL_1__11259_ (
);

FILL FILL_0__8686_ (
);

FILL FILL_3__6783_ (
);

FILL FILL_0__8266_ (
);

NAND3X1 _10957_ (
    .A(_4152_),
    .B(_4137_),
    .C(_4156_),
    .Y(_4157_)
);

NAND2X1 _10537_ (
    .A(_3808_),
    .B(_3807_),
    .Y(_3809_)
);

AOI21X1 _10117_ (
    .A(_3360_),
    .B(_3364_),
    .C(_3326_),
    .Y(_3396_)
);

FILL FILL_1__12620_ (
);

FILL FILL_1__12200_ (
);

FILL FILL_2__9645_ (
);

FILL FILL_2__9225_ (
);

FILL FILL_1__7642_ (
);

FILL FILL_3__7988_ (
);

FILL FILL_3__7148_ (
);

FILL FILL_1__13405_ (
);

FILL FILL_0__12818_ (
);

INVX1 _10290_ (
    .A(_3560_),
    .Y(_3567_)
);

FILL FILL_1__8847_ (
);

FILL FILL_1__8427_ (
);

FILL FILL_1__8007_ (
);

FILL FILL_2__10332_ (
);

AOI21X1 _7497_ (
    .A(_944_),
    .B(_940_),
    .C(_1009_),
    .Y(_1016_)
);

OR2X2 _7077_ (
    .A(_661_),
    .B(_659_),
    .Y(_663_)
);

FILL FILL_0__6752_ (
);

NOR2X1 _11495_ (
    .A(\u_fir_pe5.rYin [8]),
    .B(\u_fir_pe5.mul [8]),
    .Y(_4678_)
);

AND2X2 _11075_ (
    .A(_4270_),
    .B(_4273_),
    .Y(_4274_)
);

FILL FILL_3__12964_ (
);

FILL FILL_2__7711_ (
);

FILL FILL_3__12124_ (
);

FILL FILL_2__11957_ (
);

FILL FILL_0__12991_ (
);

FILL FILL_2__11537_ (
);

FILL FILL_0__12571_ (
);

FILL FILL_2__11117_ (
);

FILL FILL_0__12151_ (
);

FILL FILL_0__7957_ (
);

FILL FILL_0__7537_ (
);

NAND3X1 _9643_ (
    .A(_2969_),
    .B(_2971_),
    .C(_2995_),
    .Y(_2996_)
);

FILL FILL_0__7117_ (
);

NAND3X1 _9223_ (
    .A(_2527_),
    .B(_2576_),
    .C(_2577_),
    .Y(_2583_)
);

FILL FILL_1__8180_ (
);

FILL FILL_2__8916_ (
);

FILL FILL_3__13329_ (
);

NOR2X1 _13221_ (
    .A(_6244_),
    .B(_6245_),
    .Y(_6246_)
);

FILL FILL_1__6913_ (
);

FILL FILL_3__6419_ (
);

FILL FILL_1__9385_ (
);

FILL FILL_2__11290_ (
);

FILL FILL_1__10283_ (
);

FILL FILL_0__7290_ (
);

FILL FILL_3__13082_ (
);

AOI21X1 _6768_ (
    .A(_365_),
    .B(_364_),
    .C(_300_),
    .Y(_366_)
);

FILL FILL_2__12075_ (
);

FILL FILL_1__11488_ (
);

FILL FILL_1__11068_ (
);

FILL FILL_0__8495_ (
);

FILL FILL_3__6592_ (
);

NOR2X1 _10766_ (
    .A(_4674_),
    .B(_4695_),
    .Y(_4705_)
);

FILL FILL_0__8075_ (
);

AOI21X1 _10346_ (
    .A(_3613_),
    .B(_3611_),
    .C(_3583_),
    .Y(_3623_)
);

FILL FILL_3__11815_ (
);

FILL FILL_2__10808_ (
);

FILL FILL_2__9454_ (
);

FILL FILL_0__11842_ (
);

FILL FILL_2__9034_ (
);

FILL FILL_0__11422_ (
);

FILL FILL_0__11002_ (
);

FILL FILL_0__6808_ (
);

NOR2X1 _8914_ (
    .A(_2336_),
    .B(_2337_),
    .Y(_2338_)
);

FILL FILL_1__7871_ (
);

FILL FILL_1__7451_ (
);

FILL FILL_1__7031_ (
);

FILL FILL_3__7377_ (
);

FILL FILL_1__13214_ (
);

NAND3X1 _12912_ (
    .A(_5880_),
    .B(_5941_),
    .C(_5936_),
    .Y(_5950_)
);

FILL FILL_0__12627_ (
);

FILL FILL_0__12207_ (
);

FILL FILL_1__8656_ (
);

FILL FILL_1__8236_ (
);

FILL FILL_2__10981_ (
);

FILL FILL_2__10561_ (
);

FILL FILL_2__10141_ (
);

FILL FILL_3__9523_ (
);

FILL FILL_0__6981_ (
);

FILL FILL_2__6999_ (
);

FILL FILL_0__6561_ (
);

FILL FILL_2__6579_ (
);

FILL FILL_2__7940_ (
);

FILL FILL_2__7520_ (
);

FILL FILL_2__7100_ (
);

FILL FILL_2__11766_ (
);

FILL FILL_2__11346_ (
);

FILL FILL_0__12380_ (
);

FILL FILL_1__10339_ (
);

FILL FILL_0__7766_ (
);

DFFPOSX1 _9872_ (
    .D(_3184_[2]),
    .CLK(clk_bF$buf42),
    .Q(\u_fir_pe3.mul [2])
);

FILL FILL_0__7346_ (
);

OAI21X1 _9452_ (
    .A(_2808_),
    .B(_2710_),
    .C(_2523_),
    .Y(_2809_)
);

AOI22X1 _9032_ (
    .A(gnd),
    .B(\X[3] [0]),
    .C(gnd),
    .D(\X[3] [1]),
    .Y(_2395_)
);

FILL FILL_1__11700_ (
);

NAND2X1 _12089_ (
    .A(_5197_),
    .B(_5204_),
    .Y(_5206_)
);

FILL FILL_2__8725_ (
);

FILL FILL_2__8305_ (
);

FILL FILL_0__13165_ (
);

NAND3X1 _13030_ (
    .A(_6049_),
    .B(_6065_),
    .C(_6063_),
    .Y(_6066_)
);

FILL FILL_1__6722_ (
);

FILL FILL_3__6648_ (
);

FILL FILL_1__9194_ (
);

FILL FILL_1__12905_ (
);

FILL FILL_0__9912_ (
);

FILL FILL253950x25350 (
);

FILL FILL_1__10092_ (
);

FILL FILL_1__7927_ (
);

FILL FILL_1__7507_ (
);

NOR2X1 _6997_ (
    .A(_586_),
    .B(_590_),
    .Y(_796_[12])
);

NAND3X1 _6577_ (
    .A(_172_),
    .B(_138_),
    .C(_176_),
    .Y(_177_)
);

FILL FILL_1__11297_ (
);

OAI21X1 _10995_ (
    .A(_4121_),
    .B(_4193_),
    .C(_4162_),
    .Y(_4194_)
);

OR2X2 _10575_ (
    .A(_3835_),
    .B(_3840_),
    .Y(_3842_)
);

INVX1 _10155_ (
    .A(_3428_),
    .Y(_3434_)
);

FILL FILL_3__11204_ (
);

FILL FILL_2__9683_ (
);

FILL FILL_2__10617_ (
);

FILL FILL_2__9263_ (
);

FILL FILL_0__11651_ (
);

FILL FILL_0__11231_ (
);

FILL FILL_2__13089_ (
);

FILL FILL_0__6617_ (
);

INVX1 _8723_ (
    .A(_2156_),
    .Y(_2157_)
);

NAND2X1 _8303_ (
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_1743_)
);

FILL FILL_1__7680_ (
);

FILL FILL_1__7260_ (
);

FILL FILL_0__9089_ (
);

FILL FILL_3__12829_ (
);

FILL FILL_1__13023_ (
);

FILL FILL_0__12856_ (
);

OAI21X1 _12721_ (
    .A(_5759_),
    .B(_5760_),
    .C(_5758_),
    .Y(_5761_)
);

FILL FILL_0__12436_ (
);

FILL FILL_0__12016_ (
);

OAI21X1 _12301_ (
    .A(_5349_),
    .B(_5399_),
    .C(_5377_),
    .Y(_5412_)
);

AOI21X1 _9928_ (
    .A(_3207_),
    .B(_3208_),
    .C(_3974_),
    .Y(_3211_)
);

NAND2X1 _9508_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2864_)
);

FILL FILL_1__8885_ (
);

FILL FILL_1__8465_ (
);

FILL FILL_1__8045_ (
);

FILL FILL_2__10790_ (
);

FILL FILL_2__10370_ (
);

FILL FILL_3__9752_ (
);

FILL FILL_0__6790_ (
);

FILL FILL_2__6388_ (
);

FILL FILL_3__12582_ (
);

FILL FILL_3__12162_ (
);

FILL FILL_2__11995_ (
);

FILL FILL_2__11575_ (
);

FILL FILL_2__11155_ (
);

FILL FILL_1__10988_ (
);

FILL FILL_1__10568_ (
);

FILL FILL_1__10148_ (
);

FILL FILL_0__7995_ (
);

FILL FILL_0__7575_ (
);

NOR2X1 _9681_ (
    .A(_3022_),
    .B(_3027_),
    .Y(_3030_)
);

FILL FILL_0__7155_ (
);

NAND2X1 _9261_ (
    .A(_2618_),
    .B(_2619_),
    .Y(_2620_)
);

FILL FILL_2__8534_ (
);

FILL FILL_0__10922_ (
);

FILL FILL_0__10502_ (
);

FILL FILL_0__13394_ (
);

FILL FILL_1__6951_ (
);

FILL FILL_1__6531_ (
);

FILL FILL_2__13301_ (
);

FILL FILL_3__6877_ (
);

FILL FILL_1__12714_ (
);

FILL FILL_0__9721_ (
);

FILL FILL_2__9739_ (
);

FILL FILL_0__9301_ (
);

FILL FILL_2__9319_ (
);

FILL FILL_0__11707_ (
);

FILL FILL_1__7736_ (
);

FILL FILL_1__7316_ (
);

INVX1 _6386_ (
    .A(Xin[2]),
    .Y(_770_)
);

FILL FILL_3__8603_ (
);

OAI21X1 _10384_ (
    .A(_3607_),
    .B(_3659_),
    .C(_3595_),
    .Y(_3660_)
);

FILL FILL_0__10099_ (
);

FILL FILL_2__6600_ (
);

FILL FILL_3__11433_ (
);

FILL FILL_2__10846_ (
);

FILL FILL_2__9492_ (
);

FILL FILL_0__11880_ (
);

FILL FILL_2__10426_ (
);

FILL FILL_2__9072_ (
);

FILL FILL_0__11460_ (
);

FILL FILL_2__10006_ (
);

FILL FILL_0__11040_ (
);

FILL FILL_0__6846_ (
);

NOR2X1 _8952_ (
    .A(_2373_),
    .B(_2380_),
    .Y(_2387_[2])
);

FILL FILL_0__6426_ (
);

AOI21X1 _8532_ (
    .A(_1883_),
    .B(_1798_),
    .C(_1969_),
    .Y(_1970_)
);

DFFPOSX1 _8112_ (
    .D(\Y[1] [12]),
    .CLK(clk_bF$buf25),
    .Q(\u_fir_pe1.rYin [12])
);

DFFPOSX1 _11589_ (
    .D(_4775_[5]),
    .CLK(clk_bF$buf39),
    .Q(\Y[6] [5])
);

AOI21X1 _11169_ (
    .A(_4346_),
    .B(_4345_),
    .C(_4288_),
    .Y(_4366_)
);

FILL FILL_2__7805_ (
);

FILL FILL_3__12218_ (
);

FILL FILL_1__13252_ (
);

AND2X2 _12950_ (
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5987_)
);

FILL FILL_0__12665_ (
);

FILL FILL_0__12245_ (
);

NOR2X1 _12530_ (
    .A(_6359_),
    .B(_6339_),
    .Y(_6362_)
);

OAI21X1 _12110_ (
    .A(_5217_),
    .B(_5216_),
    .C(_5167_),
    .Y(_5227_)
);

NAND2X1 _9737_ (
    .A(_3076_),
    .B(_3079_),
    .Y(_3181_[7])
);

OAI21X1 _9317_ (
    .A(_2675_),
    .B(_2671_),
    .C(_2587_),
    .Y(_2676_)
);

FILL FILL_1__8694_ (
);

FILL FILL_1__8274_ (
);

FILL FILL_3__9981_ (
);

FILL FILL_3__9141_ (
);

INVX1 _13315_ (
    .A(\u_fir_pe7.rYin [14]),
    .Y(_6338_)
);

FILL FILL_1_CLKBUF1_insert30 (
);

FILL FILL_1_CLKBUF1_insert31 (
);

FILL FILL_1_CLKBUF1_insert32 (
);

FILL FILL_1_CLKBUF1_insert33 (
);

FILL FILL_1_CLKBUF1_insert34 (
);

FILL FILL_1__9899_ (
);

FILL FILL_1__9479_ (
);

FILL FILL_1_CLKBUF1_insert35 (
);

FILL FILL_1__9059_ (
);

FILL FILL_3__12391_ (
);

FILL FILL_1_CLKBUF1_insert36 (
);

FILL FILL_1_CLKBUF1_insert37 (
);

FILL FILL_1_CLKBUF1_insert38 (
);

FILL FILL_1_CLKBUF1_insert39 (
);

FILL FILL_2__11384_ (
);

FILL FILL_1__10797_ (
);

FILL FILL_1__10377_ (
);

FILL FILL_0__7384_ (
);

NAND2X1 _9490_ (
    .A(_2845_),
    .B(_2688_),
    .Y(_2846_)
);

NAND3X1 _9070_ (
    .A(gnd),
    .B(\X[3] [2]),
    .C(_2422_),
    .Y(_2432_)
);

FILL FILL_2__8763_ (
);

FILL FILL_2__8343_ (
);

FILL FILL_3__13176_ (
);

FILL FILL_0__10311_ (
);

FILL FILL_2__12589_ (
);

FILL FILL_2__12169_ (
);

NAND2X1 _7803_ (
    .A(gnd),
    .B(_1271_),
    .Y(_1318_)
);

FILL FILL_1__6760_ (
);

FILL FILL_2__13110_ (
);

FILL FILL_0__8589_ (
);

FILL FILL_0__8169_ (
);

FILL FILL_1__12943_ (
);

FILL FILL_1__12523_ (
);

FILL FILL_1__12103_ (
);

FILL FILL_2__9968_ (
);

FILL FILL_0__9950_ (
);

FILL FILL_0__9530_ (
);

FILL FILL_2__9548_ (
);

FILL FILL_0__11936_ (
);

FILL FILL_2__9128_ (
);

FILL FILL_0__9110_ (
);

NAND2X1 _11801_ (
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_4921_)
);

FILL FILL_0__11516_ (
);

FILL FILL_1__7965_ (
);

FILL FILL_1__7545_ (
);

FILL FILL_1__7125_ (
);

FILL FILL_1__13308_ (
);

FILL FILL_3__8832_ (
);

FILL FILL254250x93750 (
);

AOI21X1 _10193_ (
    .A(_3471_),
    .B(_3470_),
    .C(_3469_),
    .Y(_3472_)
);

FILL FILL_3__11662_ (
);

FILL FILL_2__10655_ (
);

FILL FILL_2__10235_ (
);

FILL FILL_3__9617_ (
);

FILL FILL_0__6655_ (
);

OR2X2 _8761_ (
    .A(_2166_),
    .B(_2192_),
    .Y(_2194_)
);

NAND3X1 _8341_ (
    .A(_1778_),
    .B(_1779_),
    .C(_1780_),
    .Y(_1781_)
);

FILL FILL253950x144150 (
);

OAI21X1 _11398_ (
    .A(_4548_),
    .B(_4561_),
    .C(_4565_),
    .Y(_4591_)
);

FILL FILL_2__7614_ (
);

FILL FILL_3__12447_ (
);

FILL FILL_1__13061_ (
);

FILL FILL_0__12894_ (
);

FILL FILL_0__12054_ (
);

FILL FILL_2__12801_ (
);

OR2X2 _9966_ (
    .A(_3247_),
    .B(_3246_),
    .Y(_3248_)
);

NOR2X1 _9546_ (
    .A(_2898_),
    .B(_2901_),
    .Y(_3187_[10])
);

NAND3X1 _9126_ (
    .A(_2475_),
    .B(_2486_),
    .C(_2482_),
    .Y(_2487_)
);

FILL FILL_0__8801_ (
);

FILL FILL_2__8819_ (
);

FILL FILL_3__9790_ (
);

FILL FILL_3__9370_ (
);

FILL FILL_0__13259_ (
);

AOI21X1 _13124_ (
    .A(_6156_),
    .B(_6157_),
    .C(_6140_),
    .Y(_6158_)
);

FILL FILL_1__6816_ (
);

FILL FILL_1__9288_ (
);

FILL FILL_2__11193_ (
);

FILL FILL_1__10186_ (
);

FILL FILL_0__7193_ (
);

FILL FILL_3__10933_ (
);

FILL FILL_3__10513_ (
);

FILL FILL_2__8572_ (
);

FILL FILL_0__10960_ (
);

FILL FILL_2__8152_ (
);

FILL FILL_0__10540_ (
);

FILL FILL_0__10120_ (
);

FILL FILL_2__12398_ (
);

NAND2X1 _7612_ (
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1130_)
);

FILL FILL_0__8398_ (
);

FILL FILL_3__6495_ (
);

NOR2X1 _10669_ (
    .A(\u_fir_pe4.rYin [12]),
    .B(\u_fir_pe4.mul [12]),
    .Y(_3933_)
);

NAND3X1 _10249_ (
    .A(_3512_),
    .B(_3514_),
    .C(_3516_),
    .Y(_3527_)
);

FILL FILL_3__11718_ (
);

FILL FILL_1__12752_ (
);

FILL FILL_1__12332_ (
);

FILL FILL_2__9777_ (
);

FILL FILL_2__9357_ (
);

FILL FILL_0__11745_ (
);

DFFPOSX1 _11610_ (
    .D(\Y[5] [2]),
    .CLK(clk_bF$buf5),
    .Q(\u_fir_pe5.rYin [2])
);

FILL FILL_0__11325_ (
);

NOR2X1 _8817_ (
    .A(_2242_),
    .B(_2243_),
    .Y(_2244_)
);

FILL FILL_1__7774_ (
);

FILL FILL_1__7354_ (
);

FILL FILL_1__13117_ (
);

INVX1 _12815_ (
    .A(_5756_),
    .Y(_5854_)
);

FILL FILL_3__8221_ (
);

FILL FILL_3__11891_ (
);

FILL FILL_1__8559_ (
);

FILL FILL_1__8139_ (
);

FILL FILL_3__11051_ (
);

FILL FILL_2__10884_ (
);

FILL FILL_2__10464_ (
);

FILL FILL_2__10044_ (
);

FILL FILL_1__9920_ (
);

FILL FILL_1__9500_ (
);

FILL FILL_0__6884_ (
);

DFFPOSX1 _8990_ (
    .D(\Y[2] [13]),
    .CLK(clk_bF$buf3),
    .Q(\u_fir_pe2.rYin [13])
);

FILL FILL_0__6464_ (
);

OAI21X1 _8570_ (
    .A(_1927_),
    .B(_2006_),
    .C(_2005_),
    .Y(_2007_)
);

INVX1 _8150_ (
    .A(_2381_),
    .Y(_2382_)
);

FILL FILL_2__7843_ (
);

FILL FILL_3__12676_ (
);

FILL FILL_2__7423_ (
);

FILL FILL_3__12256_ (
);

FILL FILL_2__7003_ (
);

FILL FILL_1__13290_ (
);

FILL FILL_2__11669_ (
);

FILL FILL_2__11249_ (
);

FILL FILL_0__12283_ (
);

FILL FILL_2__12610_ (
);

FILL FILL_0__7669_ (
);

NOR2X1 _9775_ (
    .A(_3118_),
    .B(_3117_),
    .Y(_3119_)
);

OAI21X1 _9355_ (
    .A(_2709_),
    .B(_2712_),
    .C(_2711_),
    .Y(_2713_)
);

FILL FILL_2__8628_ (
);

FILL FILL_0__8610_ (
);

FILL FILL_2__8208_ (
);

FILL FILL_0__13068_ (
);

DFFPOSX1 _13353_ (
    .D(_6369_[15]),
    .CLK(clk_bF$buf9),
    .Q(\Y[7] [15])
);

FILL FILL_1__6625_ (
);

FILL FILL_1__9097_ (
);

FILL FILL_1__12808_ (
);

FILL FILL_0__9815_ (
);

FILL FILL_3__7912_ (
);

FILL FILL_2__8381_ (
);

OAI21X1 _7841_ (
    .A(_1308_),
    .B(_1349_),
    .C(_1348_),
    .Y(_1355_)
);

INVX2 _7421_ (
    .A(\X[1] [6]),
    .Y(_941_)
);

INVX1 _7001_ (
    .A(_593_),
    .Y(_594_)
);

NAND3X1 _10898_ (
    .A(_4086_),
    .B(_4090_),
    .C(_4092_),
    .Y(_4099_)
);

INVX1 _10478_ (
    .A(_3714_),
    .Y(_3752_)
);

NAND2X1 _10058_ (
    .A(_3337_),
    .B(_3329_),
    .Y(_3338_)
);

FILL FILL_1__12981_ (
);

FILL FILL_3__11527_ (
);

FILL FILL_1__12561_ (
);

FILL FILL_1__12141_ (
);

FILL FILL_0__11974_ (
);

FILL FILL_2__9586_ (
);

FILL FILL_2__9166_ (
);

FILL FILL_0__11554_ (
);

FILL FILL_0__11134_ (
);

NAND2X1 _8626_ (
    .A(gnd),
    .B(_1992_),
    .Y(_2062_)
);

INVX1 _8206_ (
    .A(_1647_),
    .Y(_1648_)
);

FILL FILL_1__7583_ (
);

FILL FILL_1__7163_ (
);

FILL FILL_3__7089_ (
);

FILL FILL_0__12759_ (
);

FILL FILL_3__8450_ (
);

INVX1 _12624_ (
    .A(_5664_),
    .Y(_5665_)
);

FILL FILL_0__12339_ (
);

NAND2X1 _12204_ (
    .A(_5318_),
    .B(_5298_),
    .Y(_5319_)
);

FILL FILL_1__8788_ (
);

FILL FILL_1__8368_ (
);

FILL FILL_3__11280_ (
);

FILL FILL_2__10693_ (
);

FILL FILL_2__10273_ (
);

FILL FILL_3__9235_ (
);

BUFX2 _13409_ (
    .A(_6377_[15]),
    .Y(Yout[15])
);

FILL FILL_0__6693_ (
);

FILL FILL_2__7652_ (
);

FILL FILL_3__12065_ (
);

FILL FILL_2__11898_ (
);

FILL FILL_2__11478_ (
);

FILL FILL_2__11058_ (
);

FILL FILL_0__12092_ (
);

FILL FILL_0__7898_ (
);

FILL FILL_0__7478_ (
);

NAND2X1 _9584_ (
    .A(_2938_),
    .B(_2905_),
    .Y(_2939_)
);

FILL FILL_0__7058_ (
);

OAI21X1 _9164_ (
    .A(_3101_),
    .B(_2523_),
    .C(_2468_),
    .Y(_2524_)
);

FILL FILL_1__11832_ (
);

FILL FILL_1__11412_ (
);

FILL FILL_2__8857_ (
);

FILL FILL_2__8437_ (
);

FILL FILL_0__10825_ (
);

FILL FILL_0__10405_ (
);

FILL FILL_2__8017_ (
);

FILL FILL_0__13297_ (
);

AOI21X1 _13162_ (
    .A(_6136_),
    .B(_6138_),
    .C(_6193_),
    .Y(_6194_)
);

FILL FILL_1__6854_ (
);

FILL FILL_1__6434_ (
);

FILL FILL_2__13204_ (
);

FILL FILL_1__12617_ (
);

FILL FILL_0__9624_ (
);

FILL FILL_3__7721_ (
);

FILL FILL_0__9204_ (
);

FILL FILL_1__7639_ (
);

FILL FILL_3__10131_ (
);

FILL FILL_2__8190_ (
);

FILL FILL_3__8926_ (
);

NAND3X1 _7650_ (
    .A(_1098_),
    .B(_1159_),
    .C(_1154_),
    .Y(_1168_)
);

DFFPOSX1 _7230_ (
    .D(Yin[7]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.rYin [7])
);

AND2X2 _10287_ (
    .A(_3555_),
    .B(_3560_),
    .Y(_3565_)
);

FILL FILL_2__6923_ (
);

FILL FILL_3__11756_ (
);

FILL FILL_2__6503_ (
);

FILL FILL_1__12790_ (
);

FILL FILL_1__12370_ (
);

FILL FILL_2__9395_ (
);

FILL FILL_0__11783_ (
);

FILL FILL_2__10329_ (
);

FILL FILL_0__11363_ (
);

FILL FILL_0__6749_ (
);

NOR2X1 _8855_ (
    .A(\u_fir_pe2.rYin [7]),
    .B(\u_fir_pe2.mul [7]),
    .Y(_2278_)
);

AOI21X1 _8435_ (
    .A(_1873_),
    .B(_1868_),
    .C(_1729_),
    .Y(_1874_)
);

AOI21X1 _8015_ (
    .A(_1500_),
    .B(_1515_),
    .C(_1518_),
    .Y(_1519_)
);

FILL FILL_1__7392_ (
);

FILL FILL_2__7708_ (
);

FILL FILL_1__13155_ (
);

FILL FILL_0__12988_ (
);

OR2X2 _12853_ (
    .A(_5886_),
    .B(_5885_),
    .Y(_5891_)
);

FILL FILL_0__12568_ (
);

FILL FILL_0__12148_ (
);

NOR2X1 _12433_ (
    .A(_5536_),
    .B(_5535_),
    .Y(_5537_)
);

NAND3X1 _12013_ (
    .A(_5124_),
    .B(_5125_),
    .C(_5126_),
    .Y(_5131_)
);

FILL FILL_1__8597_ (
);

FILL FILL_1__8177_ (
);

FILL FILL_2__10082_ (
);

FILL FILL_3__9464_ (
);

OAI21X1 _13218_ (
    .A(_6234_),
    .B(_6235_),
    .C(_6241_),
    .Y(_6243_)
);

FILL FILL_2__7881_ (
);

FILL FILL_2__7461_ (
);

FILL FILL_2__7041_ (
);

FILL FILL_2__11287_ (
);

NAND2X1 _6921_ (
    .A(_484_),
    .B(_487_),
    .Y(_516_)
);

NAND2X1 _6501_ (
    .A(_81_),
    .B(_77_),
    .Y(_102_)
);

FILL FILL_0__7287_ (
);

NAND3X1 _9393_ (
    .A(_2744_),
    .B(_2745_),
    .C(_2746_),
    .Y(_2751_)
);

FILL FILL_3__10607_ (
);

FILL FILL_1__11641_ (
);

FILL FILL_1__11221_ (
);

FILL FILL_2__8666_ (
);

FILL FILL_2__8246_ (
);

FILL FILL_0__10634_ (
);

FILL FILL_0__10214_ (
);

DFFPOSX1 _13391_ (
    .D(_6375_[13]),
    .CLK(clk_bF$buf26),
    .Q(\u_fir_pe7.mul [13])
);

NAND3X1 _7706_ (
    .A(_1192_),
    .B(_1220_),
    .C(_1222_),
    .Y(_1223_)
);

FILL FILL_1__6663_ (
);

FILL FILL_2__13013_ (
);

FILL FILL_3__6589_ (
);

FILL FILL_1__12846_ (
);

FILL FILL_1__12426_ (
);

FILL FILL_1__12006_ (
);

FILL FILL_0__9433_ (
);

FILL FILL_0__11839_ (
);

FILL FILL_3__7530_ (
);

FILL FILL_0__9013_ (
);

NAND3X1 _11704_ (
    .A(_4815_),
    .B(_4823_),
    .C(_4825_),
    .Y(_4826_)
);

FILL FILL_0__11419_ (
);

FILL FILL_1__7868_ (
);

FILL FILL_3__10780_ (
);

FILL FILL_1__7448_ (
);

FILL FILL_3__10360_ (
);

FILL FILL_1__7028_ (
);

AOI21X1 _12909_ (
    .A(_5857_),
    .B(_5856_),
    .C(_5788_),
    .Y(_5947_)
);

FILL FILL_3__8315_ (
);

AOI22X1 _10096_ (
    .A(_3299_),
    .B(_3294_),
    .C(_3371_),
    .D(_3375_),
    .Y(_3376_)
);

FILL FILL_3__11985_ (
);

FILL FILL_2__6732_ (
);

FILL FILL_3__11145_ (
);

FILL FILL_2__10978_ (
);

FILL FILL_2__10558_ (
);

FILL FILL_2__10138_ (
);

FILL FILL_0__11172_ (
);

FILL FILL_0__6978_ (
);

FILL FILL_0__6558_ (
);

INVX1 _8664_ (
    .A(_2099_),
    .Y(_2100_)
);

NAND3X1 _8244_ (
    .A(_1680_),
    .B(_1684_),
    .C(_1682_),
    .Y(_1685_)
);

FILL FILL_1__10912_ (
);

FILL FILL_2__7937_ (
);

FILL FILL_2__7517_ (
);

FILL FILL_0__12797_ (
);

NAND3X1 _12662_ (
    .A(_5632_),
    .B(_5696_),
    .C(_5697_),
    .Y(_5703_)
);

FILL FILL_0__12377_ (
);

INVX1 _12242_ (
    .A(_5353_),
    .Y(_5356_)
);

FILL FILL_2__12704_ (
);

DFFPOSX1 _9869_ (
    .D(\Y[3] [15]),
    .CLK(clk_bF$buf4),
    .Q(\u_fir_pe3.rYin [15])
);

NAND3X1 _9449_ (
    .A(_2791_),
    .B(_2798_),
    .C(_2805_),
    .Y(_2806_)
);

INVX1 _9029_ (
    .A(_2391_),
    .Y(_2392_)
);

FILL FILL_0__8704_ (
);

FILL FILL_3__6801_ (
);

FILL FILL_3__9693_ (
);

NAND2X1 _13027_ (
    .A(_6062_),
    .B(_6051_),
    .Y(_6063_)
);

FILL FILL_1__6719_ (
);

FILL FILL_2__7690_ (
);

FILL FILL_2__7270_ (
);

FILL FILL_0__9909_ (
);

FILL FILL_2__11096_ (
);

OAI21X1 _6730_ (
    .A(_89_),
    .B(_144_),
    .C(_327_),
    .Y(_328_)
);

FILL FILL_1__10089_ (
);

FILL FILL_0__7096_ (
);

FILL FILL_1__11870_ (
);

FILL FILL_1__11450_ (
);

FILL FILL_1__11030_ (
);

FILL FILL_2__8895_ (
);

FILL FILL_2__8475_ (
);

FILL FILL_0__10863_ (
);

FILL FILL_0__10443_ (
);

FILL FILL_2__8055_ (
);

FILL FILL_0__10023_ (
);

NAND2X1 _7935_ (
    .A(_1442_),
    .B(_1441_),
    .Y(_1443_)
);

NAND3X1 _7515_ (
    .A(_1022_),
    .B(_1031_),
    .C(_1033_),
    .Y(_1034_)
);

FILL FILL_1__6892_ (
);

FILL FILL_1__6472_ (
);

FILL FILL_2__13242_ (
);

FILL FILL_1__12655_ (
);

FILL FILL_1__12235_ (
);

FILL FILL_0__9662_ (
);

FILL FILL_0__9242_ (
);

FILL FILL_0__11648_ (
);

AND2X2 _11933_ (
    .A(_5003_),
    .B(_5000_),
    .Y(_5052_)
);

AND2X2 _11513_ (
    .A(\u_fir_pe5.rYin [9]),
    .B(\u_fir_pe5.mul [9]),
    .Y(_4697_)
);

FILL FILL_0__11228_ (
);

FILL FILL_1__7677_ (
);

FILL FILL_1__7257_ (
);

FILL FILL254550x18150 (
);

FILL FILL_3__8544_ (
);

AOI21X1 _12718_ (
    .A(_5661_),
    .B(_5679_),
    .C(_5757_),
    .Y(_5758_)
);

FILL FILL_2__6961_ (
);

FILL FILL_2__6541_ (
);

FILL FILL_3__11374_ (
);

FILL FILL_2__10787_ (
);

FILL FILL_2__10367_ (
);

FILL FILL_1__9823_ (
);

FILL FILL_1__9403_ (
);

FILL FILL_0_CLKBUF1_insert40 (
);

FILL FILL254250x25350 (
);

FILL FILL_3__9329_ (
);

FILL FILL_0_CLKBUF1_insert41 (
);

FILL FILL_0_CLKBUF1_insert42 (
);

FILL FILL_0_CLKBUF1_insert43 (
);

FILL FILL_0_CLKBUF1_insert44 (
);

FILL FILL_0__6787_ (
);

FILL FILL_0_CLKBUF1_insert45 (
);

INVX1 _8893_ (
    .A(_2316_),
    .Y(_2317_)
);

OAI21X1 _8473_ (
    .A(_1832_),
    .B(_1910_),
    .C(_1854_),
    .Y(_1911_)
);

FILL FILL_0_CLKBUF1_insert46 (
);

FILL FILL_0_CLKBUF1_insert47 (
);

INVX1 _8053_ (
    .A(\u_fir_pe1.rYin [14]),
    .Y(_1556_)
);

FILL FILL_0_CLKBUF1_insert48 (
);

FILL FILL_0_CLKBUF1_insert49 (
);

FILL FILL_1__10301_ (
);

FILL FILL_3__12999_ (
);

FILL FILL_2__7746_ (
);

FILL FILL_2__7326_ (
);

FILL FILL_3__12159_ (
);

FILL FILL_1__13193_ (
);

NAND3X1 _12891_ (
    .A(_5901_),
    .B(_5919_),
    .C(_5915_),
    .Y(_5929_)
);

FILL FILL_0__12186_ (
);

DFFPOSX1 _12471_ (
    .D(_5572_[10]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[10])
);

NAND2X1 _12051_ (
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_5168_)
);

FILL FILL_3__13100_ (
);

FILL FILL_2__12933_ (
);

NOR2X1 _9678_ (
    .A(_3026_),
    .B(_3025_),
    .Y(_3027_)
);

INVX1 _9258_ (
    .A(_2616_),
    .Y(_2617_)
);

FILL FILL_1__11926_ (
);

FILL FILL_1__11506_ (
);

FILL FILL_0__8933_ (
);

FILL FILL_0__8513_ (
);

FILL FILL_0__10919_ (
);

FILL FILL_3__9082_ (
);

AND2X2 _13256_ (
    .A(_6238_),
    .B(_6248_),
    .Y(_6280_)
);

FILL FILL_1__6948_ (
);

FILL FILL_1__6528_ (
);

FILL FILL_0__9718_ (
);

FILL FILL_3__7815_ (
);

FILL FILL_3__10225_ (
);

FILL FILL_2__8284_ (
);

FILL FILL_0__10672_ (
);

FILL FILL_0__10252_ (
);

NOR3X1 _7744_ (
    .A(_1102_),
    .B(_929_),
    .C(_1118_),
    .Y(_1260_)
);

NAND3X1 _7324_ (
    .A(_826_),
    .B(_842_),
    .C(_845_),
    .Y(_846_)
);

FILL FILL_2__13051_ (
);

FILL FILL_1__12884_ (
);

FILL FILL_1__12044_ (
);

FILL FILL_0__9891_ (
);

FILL FILL_0__9471_ (
);

FILL FILL_2__9489_ (
);

FILL FILL_0__11877_ (
);

FILL FILL_2__9069_ (
);

FILL FILL_0__9051_ (
);

NAND3X1 _11742_ (
    .A(_4852_),
    .B(_4860_),
    .C(_4862_),
    .Y(_4863_)
);

FILL FILL_0__11457_ (
);

FILL FILL_0__11037_ (
);

OAI21X1 _11322_ (
    .A(_4516_),
    .B(_4515_),
    .C(_4509_),
    .Y(_4517_)
);

AOI21X1 _8949_ (
    .A(\X[2] [0]),
    .B(gnd),
    .C(_2294_),
    .Y(_2371_)
);

NAND2X1 _8529_ (
    .A(_1966_),
    .B(_1961_),
    .Y(_1967_)
);

DFFPOSX1 _8109_ (
    .D(\Y[1] [9]),
    .CLK(clk_bF$buf25),
    .Q(\u_fir_pe1.rYin [9])
);

FILL FILL_1__7486_ (
);

FILL FILL_1__7066_ (
);

FILL FILL_1__13249_ (
);

FILL FILL_3__8773_ (
);

AND2X2 _12947_ (
    .A(vdd),
    .B(\X[6] [7]),
    .Y(_5984_)
);

NOR2X1 _12527_ (
    .A(_6349_),
    .B(_6357_),
    .Y(_6359_)
);

NAND3X1 _12107_ (
    .A(_5164_),
    .B(_5219_),
    .C(_5223_),
    .Y(_5224_)
);

FILL FILL_2__6770_ (
);

FILL FILL_2__10596_ (
);

FILL FILL_2__10176_ (
);

FILL FILL_1__9632_ (
);

FILL FILL_1__9212_ (
);

FILL FILL_3__9558_ (
);

FILL FILL_0__6596_ (
);

INVX1 _8282_ (
    .A(_1719_),
    .Y(_1723_)
);

FILL FILL_1__10950_ (
);

FILL FILL_1__10530_ (
);

FILL FILL_1__10110_ (
);

FILL FILL_2__7975_ (
);

FILL FILL_2__7555_ (
);

FILL FILL_2__7135_ (
);

NAND2X1 _12280_ (
    .A(_5371_),
    .B(_5370_),
    .Y(_5393_)
);

FILL FILL_2__12742_ (
);

FILL FILL_2__12322_ (
);

NAND2X1 _9487_ (
    .A(_2843_),
    .B(_2842_),
    .Y(_3187_[9])
);

AOI22X1 _9067_ (
    .A(gnd),
    .B(\X[3] [1]),
    .C(gnd),
    .D(\X[3] [2]),
    .Y(_2429_)
);

FILL FILL_1__11735_ (
);

FILL FILL_1__11315_ (
);

FILL FILL_0__8742_ (
);

FILL FILL_0__8322_ (
);

FILL FILL_0__10308_ (
);

NAND2X1 _13065_ (
    .A(gnd),
    .B(_6053_),
    .Y(_6100_)
);

FILL FILL_2__9701_ (
);

FILL FILL_1__6757_ (
);

FILL FILL_2__13107_ (
);

FILL FILL_0__9947_ (
);

FILL FILL_0__9527_ (
);

FILL FILL_0__9107_ (
);

FILL FILL_3__10874_ (
);

FILL FILL_3__10454_ (
);

FILL FILL_3__10034_ (
);

FILL FILL_0__10481_ (
);

FILL FILL_0__10061_ (
);

FILL FILL_1__8903_ (
);

FILL FILL_3__8409_ (
);

AND2X2 _7973_ (
    .A(_1476_),
    .B(_1475_),
    .Y(_1587_[6])
);

INVX1 _7553_ (
    .A(_974_),
    .Y(_1072_)
);

OAI21X1 _7133_ (
    .A(_712_),
    .B(_713_),
    .C(_711_),
    .Y(_717_)
);

FILL FILL_2__13280_ (
);

FILL FILL_2__6826_ (
);

FILL FILL_3__11659_ (
);

FILL FILL_2__6406_ (
);

FILL FILL_1__12693_ (
);

FILL FILL_3__11239_ (
);

FILL FILL_1__12273_ (
);

FILL FILL_0__9280_ (
);

FILL FILL_2__9298_ (
);

OAI21X1 _11971_ (
    .A(_5007_),
    .B(_5012_),
    .C(_5011_),
    .Y(_5089_)
);

FILL FILL_0__11686_ (
);

OAI21X1 _11551_ (
    .A(_4727_),
    .B(_4728_),
    .C(_4732_),
    .Y(_4734_)
);

FILL FILL_0__11266_ (
);

OAI21X1 _11131_ (
    .A(_4320_),
    .B(_4314_),
    .C(_4322_),
    .Y(_4329_)
);

FILL FILL_3__12600_ (
);

OAI22X1 _8758_ (
    .A(_1738_),
    .B(_2056_),
    .C(_1899_),
    .D(_1829_),
    .Y(_2191_)
);

AND2X2 _8338_ (
    .A(_1728_),
    .B(_1729_),
    .Y(_1778_)
);

FILL FILL_1__7295_ (
);

FILL FILL_1__13058_ (
);

NAND2X1 _12756_ (
    .A(_5792_),
    .B(_5794_),
    .Y(_5795_)
);

FILL FILL_3__8162_ (
);

INVX1 _12336_ (
    .A(_5432_),
    .Y(_5442_)
);

FILL FILL_0__13412_ (
);

FILL FILL_1__9441_ (
);

FILL FILL_1__9021_ (
);

FILL FILL_3__9787_ (
);

DFFPOSX1 _8091_ (
    .D(_1587_[15]),
    .CLK(clk_bF$buf3),
    .Q(\Y[2] [15])
);

FILL FILL_2__7784_ (
);

FILL FILL_2__7364_ (
);

FILL FILL_3__12197_ (
);

NAND2X1 _6824_ (
    .A(_406_),
    .B(_409_),
    .Y(_421_)
);

NOR2X1 _6404_ (
    .A(_731_),
    .B(_2_),
    .Y(_7_)
);

FILL FILL_2__12971_ (
);

FILL FILL_2__12551_ (
);

FILL FILL_2__12131_ (
);

INVX1 _9296_ (
    .A(_2558_),
    .Y(_2655_)
);

FILL FILL_1__11964_ (
);

FILL FILL_1__11544_ (
);

FILL FILL_1__11124_ (
);

FILL FILL_0__8551_ (
);

FILL FILL_2__8569_ (
);

FILL FILL_0__10957_ (
);

FILL FILL_2__8149_ (
);

FILL FILL_0__10537_ (
);

INVX1 _10822_ (
    .A(_4023_),
    .Y(_4024_)
);

NAND3X1 _10402_ (
    .A(_3595_),
    .B(_3671_),
    .C(_3603_),
    .Y(_3678_)
);

FILL FILL_0__10117_ (
);

AOI21X1 _13294_ (
    .A(_6314_),
    .B(_6305_),
    .C(_6312_),
    .Y(_6317_)
);

FILL FILL_2__9930_ (
);

FILL FILL_2__9510_ (
);

INVX1 _7609_ (
    .A(_1121_),
    .Y(_1127_)
);

FILL FILL_1__6986_ (
);

FILL FILL_1__6566_ (
);

FILL FILL_2__13336_ (
);

FILL FILL_1__12749_ (
);

FILL FILL_1__12329_ (
);

FILL FILL_0__9756_ (
);

FILL FILL_3__7853_ (
);

FILL FILL_0__9336_ (
);

FILL FILL_3__7433_ (
);

DFFPOSX1 _11607_ (
    .D(\X[5] [7]),
    .CLK(clk_bF$buf45),
    .Q(\X[6] [7])
);

FILL FILL_3__7013_ (
);

FILL FILL_3__10683_ (
);

FILL FILL_0__10290_ (
);

FILL FILL_1__8712_ (
);

FILL FILL_3__8638_ (
);

FILL FILL_3__8218_ (
);

NAND3X1 _7782_ (
    .A(_1293_),
    .B(_1294_),
    .C(_1297_),
    .Y(_1298_)
);

INVX1 _7362_ (
    .A(_882_),
    .Y(_883_)
);

FILL FILL_2__6635_ (
);

FILL FILL_3__11468_ (
);

FILL FILL_1__12082_ (
);

NAND3X1 _11780_ (
    .A(_4836_),
    .B(_4899_),
    .C(_4900_),
    .Y(_4901_)
);

FILL FILL_0__11495_ (
);

FILL FILL_0__11075_ (
);

AOI21X1 _11360_ (
    .A(gnd),
    .B(_4551_),
    .C(_4553_),
    .Y(_4554_)
);

FILL FILL_1__9917_ (
);

FILL FILL_2__11822_ (
);

FILL FILL_2__11402_ (
);

DFFPOSX1 _8987_ (
    .D(\Y[2] [10]),
    .CLK(clk_bF$buf10),
    .Q(\u_fir_pe2.rYin [10])
);

NAND2X1 _8567_ (
    .A(gnd),
    .B(\X[2] [7]),
    .Y(_2004_)
);

NAND2X1 _8147_ (
    .A(_2314_),
    .B(_2378_),
    .Y(_2379_)
);

FILL FILL_1__10815_ (
);

FILL FILL_0__7822_ (
);

FILL FILL_0__7402_ (
);

FILL FILL_1__13287_ (
);

INVX1 _12985_ (
    .A(_5943_),
    .Y(_6022_)
);

FILL FILL_3__8391_ (
);

NOR2X1 _12565_ (
    .A(_5606_),
    .B(_5605_),
    .Y(_5607_)
);

NAND2X1 _12145_ (
    .A(_5259_),
    .B(_5260_),
    .Y(_5261_)
);

FILL FILL_2__12607_ (
);

FILL FILL_0__13221_ (
);

FILL FILL_0__8607_ (
);

FILL FILL_1__9670_ (
);

FILL FILL_1__9250_ (
);

FILL FILL_3__9176_ (
);

FILL FILL_2__7593_ (
);

FILL FILL_2__7173_ (
);

FILL FILL_3__7909_ (
);

NAND3X1 _6633_ (
    .A(_226_),
    .B(_231_),
    .C(_229_),
    .Y(_232_)
);

FILL FILL_2__12780_ (
);

FILL FILL_2__12360_ (
);

FILL FILL_1__11773_ (
);

FILL FILL_1__11353_ (
);

FILL FILL_0__8780_ (
);

FILL FILL_2__8798_ (
);

FILL FILL_2__8378_ (
);

FILL FILL_0__8360_ (
);

FILL FILL_0__10766_ (
);

FILL FILL_0__10346_ (
);

NAND2X1 _10631_ (
    .A(_3893_),
    .B(_3894_),
    .Y(_3895_)
);

INVX1 _10211_ (
    .A(_3488_),
    .Y(_3489_)
);

NAND2X1 _7838_ (
    .A(_1351_),
    .B(_1352_),
    .Y(_1593_[11])
);

AND2X2 _7418_ (
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_938_)
);

FILL FILL_1__6795_ (
);

FILL FILL_2__13145_ (
);

FILL FILL_1__12978_ (
);

FILL FILL_1__12558_ (
);

FILL FILL_1__12138_ (
);

FILL FILL_0__9985_ (
);

FILL FILL_0__9565_ (
);

FILL FILL_0__9145_ (
);

OAI21X1 _11836_ (
    .A(_4951_),
    .B(_4952_),
    .C(_4937_),
    .Y(_4956_)
);

INVX1 _11416_ (
    .A(_4567_),
    .Y(_4608_)
);

FILL FILL_0__12912_ (
);

FILL FILL_3__10072_ (
);

FILL FILL_1__8941_ (
);

FILL FILL_1__8521_ (
);

FILL FILL_3__8867_ (
);

FILL FILL_3__8027_ (
);

OR2X2 _7591_ (
    .A(_1104_),
    .B(_1103_),
    .Y(_1109_)
);

NOR2X1 _7171_ (
    .A(_754_),
    .B(_753_),
    .Y(_755_)
);

FILL FILL_2__6864_ (
);

FILL FILL_3__11697_ (
);

FILL FILL_2__6444_ (
);

FILL FILL_1__9726_ (
);

FILL FILL_1__9306_ (
);

FILL FILL_2__11211_ (
);

AND2X2 _8796_ (
    .A(\u_fir_pe2.rYin [0]),
    .B(\u_fir_pe2.mul [0]),
    .Y(_2225_)
);

OAI21X1 _8376_ (
    .A(_1813_),
    .B(_1814_),
    .C(_1804_),
    .Y(_1815_)
);

FILL FILL_1__10624_ (
);

FILL FILL_1__10204_ (
);

FILL FILL_0__7631_ (
);

FILL FILL_2__7649_ (
);

FILL FILL_1__13096_ (
);

NAND2X1 _12794_ (
    .A(vdd),
    .B(\X[6]_5_bF$buf0 ),
    .Y(_5833_)
);

FILL FILL_0__12089_ (
);

OAI21X1 _12374_ (
    .A(_5447_),
    .B(_5448_),
    .C(_5476_),
    .Y(_5477_)
);

FILL FILL_3__13003_ (
);

FILL FILL_2__12836_ (
);

FILL FILL_2__12416_ (
);

FILL FILL_0__13030_ (
);

FILL FILL_1__11829_ (
);

FILL FILL_1__11409_ (
);

FILL FILL_0__8836_ (
);

FILL FILL_0__8416_ (
);

FILL FILL_3__6513_ (
);

NAND3X1 _13159_ (
    .A(_6163_),
    .B(_6191_),
    .C(_6190_),
    .Y(_6192_)
);

INVX1 _6862_ (
    .A(_457_),
    .Y(_458_)
);

NAND3X1 _6442_ (
    .A(_33_),
    .B(_41_),
    .C(_43_),
    .Y(_44_)
);

FILL FILL_3__10968_ (
);

FILL FILL_3__10548_ (
);

FILL FILL_1__11582_ (
);

FILL FILL_3__10128_ (
);

FILL FILL_1__11162_ (
);

FILL FILL_0__10995_ (
);

FILL FILL_2__8187_ (
);

FILL FILL_0__10575_ (
);

OAI21X1 _10860_ (
    .A(_4763_),
    .B(_4059_),
    .C(_4060_),
    .Y(_4061_)
);

OAI22X1 _10440_ (
    .A(_3421_),
    .B(_3423_),
    .C(_3507_),
    .D(_3332_),
    .Y(_3715_)
);

FILL FILL_0__10155_ (
);

OAI21X1 _10020_ (
    .A(_3296_),
    .B(_3297_),
    .C(_3257_),
    .Y(_3301_)
);

FILL FILL_2__10902_ (
);

AOI21X1 _7647_ (
    .A(_1075_),
    .B(_1074_),
    .C(_1006_),
    .Y(_1165_)
);

DFFPOSX1 _7227_ (
    .D(Yin[4]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [4])
);

FILL FILL_0__6902_ (
);

FILL FILL_1__12787_ (
);

FILL FILL_1__12367_ (
);

FILL FILL_0__9794_ (
);

FILL FILL_0__9374_ (
);

FILL FILL_3__7471_ (
);

NOR2X1 _11645_ (
    .A(_5471_),
    .B(_5513_),
    .Y(_5522_)
);

NAND3X1 _11225_ (
    .A(_4368_),
    .B(_4416_),
    .C(_4421_),
    .Y(_4422_)
);

FILL FILL_0__12721_ (
);

FILL FILL_0__12301_ (
);

FILL FILL_1__7389_ (
);

FILL FILL_1__8750_ (
);

FILL FILL_1__8330_ (
);

FILL FILL_3__8256_ (
);

FILL FILL_2__6673_ (
);

FILL FILL_3__11086_ (
);

FILL FILL_2__10499_ (
);

FILL FILL_2__10079_ (
);

FILL FILL_1__9955_ (
);

FILL FILL_1__9535_ (
);

FILL FILL_1__9115_ (
);

FILL FILL_2__11860_ (
);

FILL FILL_2__11440_ (
);

FILL FILL_2__11020_ (
);

FILL FILL_0__6499_ (
);

NAND2X1 _8185_ (
    .A(gnd),
    .B(\X[2] [3]),
    .Y(_1627_)
);

FILL FILL_1__10853_ (
);

FILL FILL_1__10433_ (
);

FILL FILL_1__10013_ (
);

FILL FILL_2__7878_ (
);

FILL FILL_0__7860_ (
);

FILL FILL_2__7458_ (
);

FILL FILL_0__7440_ (
);

FILL FILL_0__7020_ (
);

FILL FILL_2__7038_ (
);

NAND2X1 _12183_ (
    .A(_5266_),
    .B(_5269_),
    .Y(_5298_)
);

NOR2X1 _6918_ (
    .A(_493_),
    .B(_498_),
    .Y(_513_)
);

FILL FILL_2__12645_ (
);

FILL FILL_2__12225_ (
);

FILL FILL_1__11218_ (
);

FILL FILL_0__8645_ (
);

FILL FILL_3__6742_ (
);

FILL FILL_0__8225_ (
);

AND2X2 _10916_ (
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4116_)
);

DFFPOSX1 _13388_ (
    .D(_6375_[10]),
    .CLK(clk_bF$buf24),
    .Q(\u_fir_pe7.mul [10])
);

FILL FILL_2__9604_ (
);

FILL FILL_1__7601_ (
);

FILL FILL_3__7527_ (
);

FILL FILL_3__7107_ (
);

AND2X2 _6671_ (
    .A(_221_),
    .B(_218_),
    .Y(_270_)
);

FILL FILL_1__11391_ (
);

FILL FILL_0__10384_ (
);

FILL FILL_1__8806_ (
);

INVX1 _7876_ (
    .A(_1363_),
    .Y(_1389_)
);

AOI21X1 _7456_ (
    .A(_879_),
    .B(_897_),
    .C(_975_),
    .Y(_976_)
);

NAND3X1 _7036_ (
    .A(_626_),
    .B(_627_),
    .C(_625_),
    .Y(_628_)
);

FILL FILL_2__13183_ (
);

FILL FILL_2__6729_ (
);

FILL FILL_0__6711_ (
);

FILL FILL_1__12596_ (
);

FILL FILL_1__12176_ (
);

FILL FILL_0__9183_ (
);

INVX1 _11874_ (
    .A(_4992_),
    .Y(_4993_)
);

FILL FILL_3__7280_ (
);

INVX1 _11454_ (
    .A(\u_fir_pe5.rYin [4]),
    .Y(_4640_)
);

FILL FILL_0__11169_ (
);

AOI22X1 _11034_ (
    .A(vdd),
    .B(\X[5] [4]),
    .C(gnd),
    .D(\X[5]_5_bF$buf3 ),
    .Y(_4233_)
);

FILL FILL_3__12923_ (
);

FILL FILL_2__11916_ (
);

FILL FILL_0__12950_ (
);

FILL FILL_0__12530_ (
);

FILL FILL_0__12110_ (
);

FILL FILL_1__7198_ (
);

FILL FILL_1__10909_ (
);

FILL FILL_0__7916_ (
);

NOR2X1 _9602_ (
    .A(_2465_),
    .B(_2853_),
    .Y(_2956_)
);

FILL FILL_3__8485_ (
);

INVX1 _12659_ (
    .A(_5599_),
    .Y(_5700_)
);

NAND2X1 _12239_ (
    .A(_5347_),
    .B(_5351_),
    .Y(_5353_)
);

FILL FILL_0__13315_ (
);

FILL FILL_2__6482_ (
);

FILL FILL_1__9764_ (
);

FILL FILL_1__9344_ (
);

FILL FILL_1__10662_ (
);

FILL FILL_1__10242_ (
);

FILL FILL_2__7687_ (
);

FILL FILL_2__7267_ (
);

FILL FILL_3__13041_ (
);

NAND2X1 _6727_ (
    .A(gnd),
    .B(Xin_5_bF$buf0),
    .Y(_325_)
);

FILL FILL_2__12874_ (
);

FILL FILL_2__12454_ (
);

FILL FILL_2__12034_ (
);

INVX1 _9199_ (
    .A(_2546_),
    .Y(_2559_)
);

FILL FILL_1__11867_ (
);

FILL FILL_1__11447_ (
);

FILL FILL_1__11027_ (
);

FILL FILL_0__8874_ (
);

FILL FILL_3__6971_ (
);

FILL FILL_0__8454_ (
);

DFFPOSX1 _10725_ (
    .D(\X[4] [2]),
    .CLK(clk_bF$buf13),
    .Q(\X[5] [2])
);

FILL FILL_0__8034_ (
);

NAND3X1 _10305_ (
    .A(_3580_),
    .B(_3576_),
    .C(_3581_),
    .Y(_3582_)
);

NAND2X1 _13197_ (
    .A(_6224_),
    .B(_6223_),
    .Y(_6225_)
);

FILL FILL_0__11801_ (
);

FILL FILL_2__9413_ (
);

FILL FILL_1__6889_ (
);

FILL FILL_1__6469_ (
);

FILL FILL_2__13239_ (
);

FILL FILL_1__7830_ (
);

FILL FILL_1__7410_ (
);

FILL FILL_0__9659_ (
);

FILL FILL_3__7756_ (
);

FILL FILL_0__9239_ (
);

NAND3X1 _6480_ (
    .A(_70_),
    .B(_78_),
    .C(_80_),
    .Y(_81_)
);

FILL FILL_3__10166_ (
);

FILL FILL_0__10193_ (
);

FILL FILL_1__8615_ (
);

FILL FILL_2__10940_ (
);

FILL FILL_2__10520_ (
);

FILL FILL_2__10100_ (
);

AND2X2 _7685_ (
    .A(vdd),
    .B(\X[1] [7]),
    .Y(_1202_)
);

NOR2X1 _7265_ (
    .A(_1567_),
    .B(_1575_),
    .Y(_1577_)
);

FILL FILL_3__9902_ (
);

FILL FILL_0__6940_ (
);

FILL FILL_2__6958_ (
);

FILL FILL_2__6538_ (
);

FILL FILL_0__6520_ (
);

NOR2X1 _11683_ (
    .A(_4805_),
    .B(_4804_),
    .Y(_5576_[3])
);

FILL FILL_0__11398_ (
);

NOR2X1 _11263_ (
    .A(_4458_),
    .B(_4401_),
    .Y(_4459_)
);

FILL FILL_3__12312_ (
);

FILL FILL_2__11725_ (
);

FILL FILL_2__11305_ (
);

FILL FILL_0__7725_ (
);

DFFPOSX1 _9831_ (
    .D(_3181_[1]),
    .CLK(clk_bF$buf56),
    .Q(\Y[4] [1])
);

FILL FILL_0__7305_ (
);

NAND2X1 _9411_ (
    .A(_2768_),
    .B(_2767_),
    .Y(_2769_)
);

INVX1 _12888_ (
    .A(_5839_),
    .Y(_5926_)
);

DFFPOSX1 _12468_ (
    .D(_5572_[7]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[7])
);

OAI21X1 _12048_ (
    .A(_5086_),
    .B(_5090_),
    .C(_5095_),
    .Y(_5165_)
);

FILL FILL_0__13124_ (
);

FILL FILL_3__6607_ (
);

FILL FILL_1__9993_ (
);

FILL FILL_1__9573_ (
);

FILL FILL_1__9153_ (
);

FILL FILL_3__9499_ (
);

FILL FILL_1__10891_ (
);

FILL FILL_1__10471_ (
);

FILL FILL_1__10051_ (
);

FILL FILL_2__7496_ (
);

FILL FILL_2__7076_ (
);

FILL FILL254550x154950 (
);

FILL FILL_3__13270_ (
);

NAND3X1 _6956_ (
    .A(_542_),
    .B(_546_),
    .C(_550_),
    .Y(_551_)
);

NAND2X1 _6536_ (
    .A(_135_),
    .B(_134_),
    .Y(_136_)
);

FILL FILL_2__12683_ (
);

FILL FILL_2__12263_ (
);

FILL FILL_1__11676_ (
);

FILL FILL_1__11256_ (
);

FILL FILL_0__8683_ (
);

FILL FILL_0__8263_ (
);

FILL FILL_0__10669_ (
);

AOI21X1 _10954_ (
    .A(_4148_),
    .B(_4150_),
    .C(_4141_),
    .Y(_4154_)
);

AND2X2 _10534_ (
    .A(_3784_),
    .B(_3783_),
    .Y(_3806_)
);

FILL FILL_0__10249_ (
);

AOI21X1 _10114_ (
    .A(_3382_),
    .B(_3390_),
    .C(_3393_),
    .Y(_3394_)
);

FILL FILL_2__9642_ (
);

FILL FILL_2__9222_ (
);

FILL FILL_1__6698_ (
);

FILL FILL_2__13048_ (
);

FILL FILL_0__9888_ (
);

FILL FILL_0__9468_ (
);

FILL FILL_0__9048_ (
);

NAND3X1 _11739_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf1 ),
    .C(_4857_),
    .Y(_4860_)
);

NAND3X1 _11319_ (
    .A(_4510_),
    .B(_4513_),
    .C(_4467_),
    .Y(_4514_)
);

FILL FILL_1__13402_ (
);

FILL FILL_0__12815_ (
);

FILL FILL_3__10395_ (
);

FILL FILL_1__8844_ (
);

FILL FILL_1__8424_ (
);

FILL FILL_1__8004_ (
);

NAND2X1 _7494_ (
    .A(_1010_),
    .B(_1012_),
    .Y(_1013_)
);

INVX1 _7074_ (
    .A(_650_),
    .Y(_660_)
);

FILL FILL_3__9711_ (
);

FILL FILL_2__6767_ (
);

INVX1 _11492_ (
    .A(\u_fir_pe5.rYin [8]),
    .Y(_4675_)
);

NAND3X1 _11072_ (
    .A(_4266_),
    .B(_4267_),
    .C(_4268_),
    .Y(_4271_)
);

FILL FILL_1__9629_ (
);

FILL FILL_1__9209_ (
);

FILL FILL_3__12541_ (
);

FILL FILL_2__11954_ (
);

FILL FILL_2__11534_ (
);

FILL FILL_2__11114_ (
);

NAND2X1 _8699_ (
    .A(_2126_),
    .B(_2129_),
    .Y(_2134_)
);

NAND3X1 _8279_ (
    .A(_1714_),
    .B(_1719_),
    .C(_1661_),
    .Y(_1720_)
);

FILL FILL_1__10947_ (
);

FILL FILL_1__10527_ (
);

FILL FILL_1__10107_ (
);

FILL FILL_0__7954_ (
);

FILL FILL_0__7534_ (
);

NAND2X1 _9640_ (
    .A(_2985_),
    .B(_2992_),
    .Y(_2993_)
);

FILL FILL_0__7114_ (
);

AOI21X1 _9220_ (
    .A(_2492_),
    .B(_2496_),
    .C(_2460_),
    .Y(_2580_)
);

AND2X2 _12697_ (
    .A(vdd),
    .B(\X[6] [4]),
    .Y(_5737_)
);

NAND2X1 _12277_ (
    .A(_5388_),
    .B(_5389_),
    .Y(_5390_)
);

FILL FILL_2__8913_ (
);

FILL FILL_3__13326_ (
);

FILL FILL_2__12739_ (
);

FILL FILL_2__12319_ (
);

FILL FILL_1__6910_ (
);

FILL FILL_0__8739_ (
);

FILL FILL_3__6836_ (
);

FILL FILL_0__8319_ (
);

FILL FILL_1__9382_ (
);

FILL FILL_1__10280_ (
);

AOI21X1 _6765_ (
    .A(_357_),
    .B(_362_),
    .C(_301_),
    .Y(_363_)
);

FILL FILL_2__12072_ (
);

FILL FILL_1__11485_ (
);

FILL FILL_1__11065_ (
);

FILL FILL_0__8492_ (
);

FILL FILL_0__10898_ (
);

FILL FILL_0__10478_ (
);

NAND2X1 _10763_ (
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4674_)
);

FILL FILL_0__8072_ (
);

INVX1 _10343_ (
    .A(_3542_),
    .Y(_3620_)
);

FILL FILL_0__10058_ (
);

FILL FILL_3__11812_ (
);

FILL FILL_2__10805_ (
);

FILL FILL_2__9451_ (
);

FILL FILL_2__9031_ (
);

FILL FILL_2__13277_ (
);

FILL FILL_0__6805_ (
);

OAI21X1 _8911_ (
    .A(_2333_),
    .B(_2316_),
    .C(_2332_),
    .Y(_2335_)
);

FILL FILL_0__9697_ (
);

FILL FILL_3__7794_ (
);

FILL FILL_0__9277_ (
);

NAND2X1 _11968_ (
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_5086_)
);

FILL FILL_3__7374_ (
);

NAND2X1 _11548_ (
    .A(_4731_),
    .B(_4726_),
    .Y(_4732_)
);

AOI21X1 _11128_ (
    .A(_4321_),
    .B(_4325_),
    .C(_4307_),
    .Y(_4326_)
);

FILL FILL_1__13211_ (
);

FILL FILL_0__12624_ (
);

FILL FILL_0__12204_ (
);

FILL FILL_1__8653_ (
);

FILL FILL_1__8233_ (
);

FILL FILL_3__8579_ (
);

FILL FILL_3__8159_ (
);

FILL FILL253950x230550 (
);

FILL FILL_3__9940_ (
);

FILL FILL_3__9100_ (
);

FILL FILL_0__13409_ (
);

FILL FILL_2__6996_ (
);

FILL FILL_2__6576_ (
);

FILL FILL_1__9438_ (
);

FILL FILL_3__12770_ (
);

FILL FILL_1__9018_ (
);

FILL FILL_2__11763_ (
);

FILL FILL_2__11343_ (
);

DFFPOSX1 _8088_ (
    .D(_1587_[12]),
    .CLK(clk_bF$buf10),
    .Q(\Y[2] [12])
);

FILL FILL_1__10336_ (
);

FILL FILL_0__7763_ (
);

FILL FILL_0__7343_ (
);

NAND2X1 _12086_ (
    .A(_5188_),
    .B(_5191_),
    .Y(_5203_)
);

FILL FILL_2__8722_ (
);

FILL FILL_2__8302_ (
);

FILL FILL_3__13135_ (
);

FILL FILL_2__12968_ (
);

FILL FILL_2__12548_ (
);

FILL FILL_2__12128_ (
);

FILL FILL_0__13162_ (
);

FILL FILL_0__8548_ (
);

AND2X2 _10819_ (
    .A(vdd),
    .B(\X[5] [2]),
    .Y(_4021_)
);

FILL FILL_1__9191_ (
);

FILL FILL_1__12902_ (
);

FILL FILL_2__9927_ (
);

FILL FILL_2__9507_ (
);

FILL FILL_1__7924_ (
);

FILL FILL_1__7504_ (
);

OAI21X1 _6994_ (
    .A(_376_),
    .B(_587_),
    .C(_559_),
    .Y(_588_)
);

OAI21X1 _6574_ (
    .A(_169_),
    .B(_170_),
    .C(_155_),
    .Y(_174_)
);

FILL FILL_1__11294_ (
);

NOR2X1 _10992_ (
    .A(_4189_),
    .B(_4191_),
    .Y(_4781_[6])
);

NOR2X1 _10572_ (
    .A(\u_fir_pe4.rYin [3]),
    .B(\u_fir_pe4.mul [3]),
    .Y(_3839_)
);

FILL FILL_0__10287_ (
);

NAND2X1 _10152_ (
    .A(_3429_),
    .B(_3430_),
    .Y(_3431_)
);

FILL FILL_1__8709_ (
);

FILL FILL_2__9680_ (
);

FILL FILL_2__10614_ (
);

FILL FILL_2__9260_ (
);

AOI21X1 _7779_ (
    .A(_1192_),
    .B(_1222_),
    .C(_1225_),
    .Y(_1295_)
);

FILL FILL254250x140550 (
);

NAND2X1 _7359_ (
    .A(vdd),
    .B(\X[1] [2]),
    .Y(_880_)
);

FILL FILL_2__13086_ (
);

FILL FILL_0__6614_ (
);

AND2X2 _8720_ (
    .A(_2136_),
    .B(_2131_),
    .Y(_2154_)
);

OAI21X1 _8300_ (
    .A(_2372_),
    .B(_1738_),
    .C(_1739_),
    .Y(_1740_)
);

FILL FILL_1__12079_ (
);

FILL FILL_0__9086_ (
);

NAND3X1 _11777_ (
    .A(_4835_),
    .B(_4893_),
    .C(_4897_),
    .Y(_4898_)
);

FILL FILL_3__7183_ (
);

NOR2X1 _11357_ (
    .A(_4458_),
    .B(_4511_),
    .Y(_4551_)
);

FILL FILL_3__12406_ (
);

FILL FILL_1__13020_ (
);

FILL FILL_2__11819_ (
);

FILL FILL_0__12853_ (
);

FILL FILL_0__12433_ (
);

FILL FILL_0__12013_ (
);

FILL FILL_0__7819_ (
);

NAND3X1 _9925_ (
    .A(_3970_),
    .B(_3202_),
    .C(_3205_),
    .Y(_3208_)
);

AND2X2 _9505_ (
    .A(_2857_),
    .B(_2860_),
    .Y(_2861_)
);

FILL FILL_1__8882_ (
);

FILL FILL_1__8462_ (
);

FILL FILL_1__8042_ (
);

FILL FILL_0__13218_ (
);

FILL FILL_2__6385_ (
);

FILL FILL_1__9667_ (
);

FILL FILL_1__9247_ (
);

FILL FILL_2__11992_ (
);

FILL FILL_2__11572_ (
);

FILL FILL_2__11152_ (
);

FILL FILL_1__10985_ (
);

FILL FILL_1__10565_ (
);

FILL FILL_1__10145_ (
);

FILL FILL_0__7992_ (
);

FILL FILL_0__7572_ (
);

FILL FILL_0__7152_ (
);

FILL FILL_2__8951_ (
);

FILL FILL_2__8531_ (
);

FILL FILL_2__12777_ (
);

FILL FILL_2__12357_ (
);

FILL FILL_0__8777_ (
);

FILL FILL_0__8357_ (
);

FILL FILL_3__6454_ (
);

OAI21X1 _10628_ (
    .A(_3880_),
    .B(_3881_),
    .C(_3891_),
    .Y(_3892_)
);

INVX1 _10208_ (
    .A(_3470_),
    .Y(_3486_)
);

FILL FILL_1__12711_ (
);

FILL FILL_2__9736_ (
);

FILL FILL_2__9316_ (
);

FILL FILL_0__11704_ (
);

FILL FILL_1__7733_ (
);

FILL FILL_1__7313_ (
);

NOR2X1 _6383_ (
    .A(_689_),
    .B(_731_),
    .Y(_740_)
);

FILL FILL_0__12909_ (
);

FILL FILL_3__8600_ (
);

FILL FILL_3__10489_ (
);

FILL FILL_3__10069_ (
);

NAND3X1 _10381_ (
    .A(_3655_),
    .B(_3652_),
    .C(_3656_),
    .Y(_3657_)
);

FILL FILL_0__10096_ (
);

FILL FILL_1__8938_ (
);

FILL FILL_1__8518_ (
);

FILL FILL_3__11010_ (
);

FILL FILL_2__10843_ (
);

FILL FILL_2__10423_ (
);

FILL FILL_2__10003_ (
);

AND2X2 _7588_ (
    .A(_1104_),
    .B(_1103_),
    .Y(_1106_)
);

INVX1 _7168_ (
    .A(\u_fir_pe0.mul [13]),
    .Y(_752_)
);

FILL FILL_3__9805_ (
);

FILL FILL_0__6843_ (
);

FILL FILL_0__6423_ (
);

DFFPOSX1 _11586_ (
    .D(_4775_[2]),
    .CLK(clk_bF$buf5),
    .Q(\Y[6] [2])
);

NAND2X1 _11166_ (
    .A(_4359_),
    .B(_4363_),
    .Y(_4781_[8])
);

FILL FILL_2__7802_ (
);

FILL FILL_3__12635_ (
);

FILL FILL_0__12662_ (
);

FILL FILL_2__11208_ (
);

FILL FILL_0__12242_ (
);

FILL FILL_0__7628_ (
);

INVX1 _9734_ (
    .A(_3071_),
    .Y(_3077_)
);

NAND3X1 _9314_ (
    .A(_2600_),
    .B(_2668_),
    .C(_2669_),
    .Y(_2673_)
);

FILL FILL_1__8691_ (
);

FILL FILL_1__8271_ (
);

FILL FILL_3__8197_ (
);

FILL FILL_0__13027_ (
);

OR2X2 _13312_ (
    .A(_6328_),
    .B(_6334_),
    .Y(_6336_)
);

FILL FILL_1__9896_ (
);

FILL FILL_1__9476_ (
);

FILL FILL_1__9056_ (
);

FILL FILL_2__11381_ (
);

FILL FILL_1__10794_ (
);

FILL FILL_1__10374_ (
);

FILL FILL_2__7399_ (
);

FILL FILL_0__7381_ (
);

FILL FILL_3__10701_ (
);

FILL FILL_2__8760_ (
);

FILL FILL_2__8340_ (
);

NAND2X1 _6859_ (
    .A(_454_),
    .B(_297_),
    .Y(_455_)
);

NAND3X1 _6439_ (
    .A(vdd),
    .B(Xin[2]),
    .C(_31_),
    .Y(_41_)
);

FILL FILL_2__12586_ (
);

FILL FILL_2__12166_ (
);

FILL FILL_1__11999_ (
);

AOI22X1 _7800_ (
    .A(\X[1]_5_bF$buf0 ),
    .B(gnd),
    .C(_1274_),
    .D(_1275_),
    .Y(_1315_)
);

FILL FILL_1__11579_ (
);

FILL FILL_1__11159_ (
);

FILL FILL_0__8586_ (
);

FILL FILL_3__6683_ (
);

FILL FILL_0__8166_ (
);

NAND2X1 _10857_ (
    .A(_4685_),
    .B(_4057_),
    .Y(_4058_)
);

NAND2X1 _10437_ (
    .A(_3707_),
    .B(_3711_),
    .Y(_3712_)
);

OAI21X1 _10017_ (
    .A(_3296_),
    .B(_3297_),
    .C(_3295_),
    .Y(_3298_)
);

FILL FILL_3__11906_ (
);

FILL FILL_1__12940_ (
);

FILL FILL_1__12520_ (
);

FILL FILL_1__12100_ (
);

FILL FILL_2__9965_ (
);

FILL FILL_2__9545_ (
);

FILL FILL_0__11933_ (
);

FILL FILL_2__9125_ (
);

FILL FILL_0__11513_ (
);

FILL FILL_1__7962_ (
);

FILL FILL_1__7542_ (
);

FILL FILL_1__7122_ (
);

FILL FILL_3__7888_ (
);

FILL FILL_3__7468_ (
);

FILL FILL_3__7048_ (
);

FILL FILL_1__13305_ (
);

FILL FILL_0__12718_ (
);

INVX1 _10190_ (
    .A(_3323_),
    .Y(_3469_)
);

FILL FILL_1__8747_ (
);

FILL FILL_1__8327_ (
);

FILL FILL_2__10652_ (
);

FILL FILL_2__10232_ (
);

INVX1 _7397_ (
    .A(_817_),
    .Y(_918_)
);

FILL FILL_0__6652_ (
);

OR2X2 _11395_ (
    .A(_4586_),
    .B(_4579_),
    .Y(_4588_)
);

FILL FILL_3__12864_ (
);

FILL FILL_2__7611_ (
);

FILL FILL_3__12024_ (
);

FILL FILL_2__11857_ (
);

FILL FILL_0__12891_ (
);

FILL FILL_2__11437_ (
);

FILL FILL_2__11017_ (
);

FILL FILL_0__12051_ (
);

FILL FILL_0__7857_ (
);

OR2X2 _9963_ (
    .A(_3244_),
    .B(_3243_),
    .Y(_3245_)
);

FILL FILL_0__7437_ (
);

NAND2X1 _9543_ (
    .A(_2768_),
    .B(_2841_),
    .Y(_2899_)
);

FILL FILL_0__7017_ (
);

NAND2X1 _9123_ (
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_2484_)
);

FILL FILL_2__8816_ (
);

FILL FILL_0__13256_ (
);

NAND2X1 _13121_ (
    .A(_6151_),
    .B(_6154_),
    .Y(_6155_)
);

FILL FILL_1__6813_ (
);

FILL FILL_1__9285_ (
);

FILL FILL_2__11190_ (
);

FILL FILL_1__10183_ (
);

FILL FILL_0__7190_ (
);

FILL FILL_3__10510_ (
);

NAND3X1 _6668_ (
    .A(_238_),
    .B(_257_),
    .C(_251_),
    .Y(_267_)
);

FILL FILL_2__12395_ (
);

FILL FILL_1__11388_ (
);

FILL FILL_0__8395_ (
);

INVX1 _10666_ (
    .A(\u_fir_pe4.rYin [12]),
    .Y(_3930_)
);

OAI21X1 _10246_ (
    .A(_3523_),
    .B(_3517_),
    .C(_3511_),
    .Y(_3524_)
);

FILL FILL253950x165750 (
);

FILL FILL_2__9774_ (
);

FILL FILL_2__9354_ (
);

FILL FILL_0__11742_ (
);

FILL FILL_0__11322_ (
);

FILL FILL_0__6708_ (
);

AOI21X1 _8814_ (
    .A(_2234_),
    .B(_2239_),
    .C(_2235_),
    .Y(_2241_)
);

FILL FILL_1__7771_ (
);

FILL FILL_1__7351_ (
);

FILL FILL_3__7697_ (
);

FILL FILL_1__13114_ (
);

FILL FILL_0__12947_ (
);

OAI21X1 _12812_ (
    .A(_5837_),
    .B(_5841_),
    .C(_5844_),
    .Y(_5851_)
);

FILL FILL_0__12527_ (
);

FILL FILL_0__12107_ (
);

FILL FILL_1__8556_ (
);

FILL FILL_1__8136_ (
);

FILL FILL_2__10881_ (
);

FILL FILL_2__10461_ (
);

FILL FILL_2__10041_ (
);

FILL FILL_3__9423_ (
);

FILL FILL_0__6881_ (
);

FILL FILL_2__6899_ (
);

FILL FILL_2__6479_ (
);

FILL FILL_0__6461_ (
);

FILL FILL_2__7840_ (
);

FILL FILL_2__7420_ (
);

FILL FILL_3__12253_ (
);

FILL FILL_2__7000_ (
);

FILL FILL_2__11666_ (
);

FILL FILL_2__11246_ (
);

FILL FILL_0__12280_ (
);

FILL FILL_1__10659_ (
);

FILL FILL_1__10239_ (
);

FILL FILL_0__7666_ (
);

INVX1 _9772_ (
    .A(\u_fir_pe3.mul [10]),
    .Y(_3116_)
);

INVX1 _9352_ (
    .A(vdd),
    .Y(_2710_)
);

FILL FILL_2__8625_ (
);

FILL FILL_2__8205_ (
);

FILL FILL_3__13038_ (
);

FILL FILL_0__13065_ (
);

DFFPOSX1 _13350_ (
    .D(_6369_[12]),
    .CLK(clk_bF$buf5),
    .Q(\Y[7] [12])
);

FILL FILL_1__6622_ (
);

FILL FILL_3__6548_ (
);

FILL FILL_1__9094_ (
);

FILL FILL_1__12805_ (
);

FILL FILL_0__9812_ (
);

FILL FILL_1__7827_ (
);

FILL FILL_1__7407_ (
);

NAND2X1 _6897_ (
    .A(_491_),
    .B(_487_),
    .Y(_493_)
);

NAND3X1 _6477_ (
    .A(gnd),
    .B(Xin_5_bF$buf1),
    .C(_75_),
    .Y(_78_)
);

FILL FILL_1__11197_ (
);

NAND3X1 _10895_ (
    .A(_4011_),
    .B(_4091_),
    .C(_4095_),
    .Y(_4096_)
);

OAI21X1 _10475_ (
    .A(_3493_),
    .B(_3667_),
    .C(_3711_),
    .Y(_3749_)
);

NAND3X1 _10055_ (
    .A(_3334_),
    .B(_3328_),
    .C(_3331_),
    .Y(_3335_)
);

FILL FILL_3__11104_ (
);

FILL FILL_2__10937_ (
);

FILL FILL_2__9583_ (
);

FILL FILL_0__11971_ (
);

FILL FILL_2__10517_ (
);

FILL FILL_2__9163_ (
);

FILL FILL_0__11551_ (
);

FILL FILL_0__11131_ (
);

FILL FILL_0__6937_ (
);

FILL FILL_0__6517_ (
);

INVX1 _8623_ (
    .A(_2058_),
    .Y(_2059_)
);

NAND3X1 _8203_ (
    .A(_1634_),
    .B(_1638_),
    .C(_1640_),
    .Y(_1645_)
);

FILL FILL_1__7580_ (
);

FILL FILL_1__7160_ (
);

FILL FILL_3__12729_ (
);

FILL FILL_0__12756_ (
);

NAND2X1 _12621_ (
    .A(vdd),
    .B(\X[6] [2]),
    .Y(_5662_)
);

FILL FILL_0__12336_ (
);

INVX1 _12201_ (
    .A(_5313_),
    .Y(_5316_)
);

NOR2X1 _9828_ (
    .A(_3111_),
    .B(_3175_),
    .Y(_3170_)
);

OAI21X1 _9408_ (
    .A(_2593_),
    .B(_2683_),
    .C(_2679_),
    .Y(_2766_)
);

FILL FILL_1__8785_ (
);

FILL FILL_1__8365_ (
);

FILL FILL_2__10690_ (
);

FILL FILL_2__10270_ (
);

FILL FILL_3__9652_ (
);

BUFX2 _13406_ (
    .A(_6377_[12]),
    .Y(Yout[12])
);

FILL FILL_0__6690_ (
);

FILL FILL_2__11895_ (
);

FILL FILL_2__11475_ (
);

FILL FILL_2__11055_ (
);

FILL FILL_1__10888_ (
);

FILL FILL_1__10468_ (
);

FILL FILL_1__10048_ (
);

FILL FILL_0__7895_ (
);

FILL FILL_0__7475_ (
);

NAND2X1 _9581_ (
    .A(_2930_),
    .B(_2927_),
    .Y(_2936_)
);

FILL FILL_0__7055_ (
);

AND2X2 _9161_ (
    .A(_2521_),
    .B(_2517_),
    .Y(_3187_[5])
);

FILL FILL_2__8854_ (
);

FILL FILL_2__8434_ (
);

FILL FILL_0__10822_ (
);

FILL FILL_0__10402_ (
);

FILL FILL_2__8014_ (
);

FILL FILL_0__13294_ (
);

FILL FILL_1__6851_ (
);

FILL FILL_1__6431_ (
);

FILL FILL_2__13201_ (
);

FILL FILL_3__6777_ (
);

FILL FILL_1__12614_ (
);

FILL FILL_0__9621_ (
);

FILL FILL_2__9639_ (
);

FILL FILL_0__9201_ (
);

FILL FILL_2__9219_ (
);

FILL FILL_1__7636_ (
);

NAND2X1 _10284_ (
    .A(_3561_),
    .B(_3485_),
    .Y(_3562_)
);

FILL FILL_2__6920_ (
);

FILL FILL_3__11753_ (
);

FILL FILL_2__6500_ (
);

FILL FILL_3__11333_ (
);

FILL FILL_2__9392_ (
);

FILL FILL_0__11780_ (
);

FILL FILL_2__10326_ (
);

FILL FILL_0__11360_ (
);

FILL FILL_0__6746_ (
);

INVX1 _8852_ (
    .A(\u_fir_pe2.rYin [7]),
    .Y(_2275_)
);

NAND3X1 _8432_ (
    .A(_1865_),
    .B(_1864_),
    .C(_1866_),
    .Y(_1871_)
);

NOR2X1 _8012_ (
    .A(_1512_),
    .B(_1506_),
    .Y(_1515_)
);

NOR2X1 _11489_ (
    .A(_4669_),
    .B(_4668_),
    .Y(_4672_)
);

OAI21X1 _11069_ (
    .A(_4254_),
    .B(_4258_),
    .C(_4261_),
    .Y(_4268_)
);

FILL FILL_3__12958_ (
);

FILL FILL_2__7705_ (
);

FILL FILL_3__12538_ (
);

FILL FILL_3__12118_ (
);

FILL FILL_1__13152_ (
);

FILL FILL_0__12985_ (
);

AND2X2 _12850_ (
    .A(_5886_),
    .B(_5885_),
    .Y(_5888_)
);

FILL FILL_0__12565_ (
);

FILL FILL_0__12145_ (
);

INVX1 _12430_ (
    .A(\u_fir_pe6.mul [13]),
    .Y(_5534_)
);

OAI21X1 _12010_ (
    .A(_5123_),
    .B(_5127_),
    .C(_5099_),
    .Y(_5128_)
);

NAND2X1 _9637_ (
    .A(_2989_),
    .B(_2963_),
    .Y(_2990_)
);

NAND3X1 _9217_ (
    .A(_2563_),
    .B(_2567_),
    .C(_2570_),
    .Y(_2577_)
);

FILL FILL_1__8594_ (
);

FILL FILL_1__8174_ (
);

FILL FILL_3__9041_ (
);

NAND2X1 _13215_ (
    .A(_6238_),
    .B(_6240_),
    .Y(_6241_)
);

FILL FILL_1__6907_ (
);

FILL FILL_1__9799_ (
);

FILL FILL_1__9379_ (
);

FILL FILL_2__11284_ (
);

FILL FILL_1__10697_ (
);

FILL FILL_1__10277_ (
);

FILL FILL_0__7284_ (
);

OAI21X1 _9390_ (
    .A(_2747_),
    .B(_2743_),
    .C(_2694_),
    .Y(_2748_)
);

FILL FILL_3__10604_ (
);

FILL FILL_2__8663_ (
);

FILL FILL_2__8243_ (
);

FILL FILL_0__10631_ (
);

FILL FILL_3__13076_ (
);

FILL FILL_0__10211_ (
);

FILL FILL_2__12069_ (
);

NAND3X1 _7703_ (
    .A(_1212_),
    .B(_1219_),
    .C(_1194_),
    .Y(_1220_)
);

FILL FILL_1__6660_ (
);

FILL FILL_2__13010_ (
);

FILL FILL_0__8489_ (
);

FILL FILL_0__8069_ (
);

FILL FILL_1__12843_ (
);

FILL FILL_1__12423_ (
);

FILL FILL_1__12003_ (
);

FILL FILL_0__9430_ (
);

FILL FILL_2__9448_ (
);

FILL FILL_0__11836_ (
);

FILL FILL_2__9028_ (
);

FILL FILL_0__9010_ (
);

NAND3X1 _11701_ (
    .A(vdd),
    .B(\X[7] [2]),
    .C(_4813_),
    .Y(_4823_)
);

FILL FILL_0__11416_ (
);

NOR2X1 _8908_ (
    .A(_2330_),
    .B(_2331_),
    .Y(_2384_[11])
);

FILL FILL_1__7865_ (
);

FILL FILL_1__7445_ (
);

FILL FILL_1__7025_ (
);

FILL FILL_1__13208_ (
);

FILL FILL_3__8732_ (
);

OAI21X1 _12906_ (
    .A(_5935_),
    .B(_5931_),
    .C(_5938_),
    .Y(_5944_)
);

FILL FILL_3__8312_ (
);

OAI21X1 _10093_ (
    .A(_3368_),
    .B(_3369_),
    .C(_3326_),
    .Y(_3373_)
);

FILL FILL_3__11982_ (
);

FILL FILL_3__11562_ (
);

FILL FILL_2__10975_ (
);

FILL FILL_2__10555_ (
);

FILL FILL_2__10135_ (
);

FILL FILL_3__9937_ (
);

FILL FILL_3__9517_ (
);

FILL FILL_0__6975_ (
);

FILL FILL_0__6555_ (
);

NAND2X1 _8661_ (
    .A(_2089_),
    .B(_2095_),
    .Y(_2097_)
);

NAND2X1 _8241_ (
    .A(_1630_),
    .B(_1681_),
    .Y(_1682_)
);

OAI21X1 _11298_ (
    .A(_4493_),
    .B(_4361_),
    .C(_4443_),
    .Y(_4494_)
);

FILL FILL_2__7934_ (
);

FILL FILL_2__7514_ (
);

FILL FILL_3__12347_ (
);

FILL FILL_0__12794_ (
);

FILL FILL_0__12374_ (
);

FILL FILL_2__12701_ (
);

DFFPOSX1 _9866_ (
    .D(\Y[3] [12]),
    .CLK(clk_bF$buf17),
    .Q(\u_fir_pe3.rYin [12])
);

NAND2X1 _9446_ (
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2803_)
);

NAND2X1 _9026_ (
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_3178_)
);

FILL FILL_0__8701_ (
);

FILL FILL_2__8719_ (
);

FILL FILL_3__9270_ (
);

FILL FILL_0__13159_ (
);

AOI21X1 _13024_ (
    .A(vdd),
    .B(\X[6] [6]),
    .C(_5991_),
    .Y(_6060_)
);

FILL FILL_1__6716_ (
);

FILL FILL_1__9188_ (
);

FILL FILL_0__9906_ (
);

FILL FILL_2__11093_ (
);

FILL FILL_1__10086_ (
);

FILL FILL_0__7093_ (
);

FILL FILL_3__10833_ (
);

FILL FILL_2__8892_ (
);

FILL FILL_2__8472_ (
);

FILL FILL_0__10860_ (
);

FILL FILL_0__10440_ (
);

FILL FILL_2__8052_ (
);

FILL FILL_0__10020_ (
);

FILL FILL_2__12298_ (
);

OAI21X1 _7932_ (
    .A(_1438_),
    .B(_1439_),
    .C(_1437_),
    .Y(_1440_)
);

OAI21X1 _7512_ (
    .A(_812_),
    .B(_1030_),
    .C(_1025_),
    .Y(_1031_)
);

FILL FILL_0__8298_ (
);

AOI21X1 _10989_ (
    .A(_4105_),
    .B(_4111_),
    .C(_4188_),
    .Y(_4189_)
);

FILL FILL_3__6395_ (
);

INVX1 _10569_ (
    .A(\u_fir_pe4.rYin [3]),
    .Y(_3836_)
);

NAND2X1 _10149_ (
    .A(vdd),
    .B(\X[4] [6]),
    .Y(_3428_)
);

FILL FILL_1__12652_ (
);

FILL FILL_1__12232_ (
);

FILL FILL_2__9677_ (
);

FILL FILL_2__9257_ (
);

NAND3X1 _11930_ (
    .A(_5020_),
    .B(_5039_),
    .C(_5033_),
    .Y(_5049_)
);

FILL FILL_0__11645_ (
);

INVX1 _11510_ (
    .A(_4677_),
    .Y(_4693_)
);

FILL FILL_0__11225_ (
);

NAND3X1 _8717_ (
    .A(_2048_),
    .B(_2150_),
    .C(_1891_),
    .Y(_2151_)
);

FILL FILL_1__7674_ (
);

FILL FILL_1__13017_ (
);

NAND3X1 _12715_ (
    .A(_5752_),
    .B(_5754_),
    .C(_5753_),
    .Y(_5755_)
);

FILL FILL_1__8879_ (
);

FILL FILL_3__11791_ (
);

FILL FILL_1__8459_ (
);

FILL FILL_1__8039_ (
);

FILL FILL_2__10784_ (
);

FILL FILL_2__10364_ (
);

FILL FILL_1__9820_ (
);

FILL FILL_1__9400_ (
);

FILL FILL_3__9746_ (
);

FILL FILL_0_CLKBUF1_insert12 (
);

FILL FILL_0_CLKBUF1_insert13 (
);

FILL FILL_0_CLKBUF1_insert14 (
);

FILL FILL_0__6784_ (
);

AOI21X1 _8890_ (
    .A(_2308_),
    .B(_2286_),
    .C(_2306_),
    .Y(_2313_)
);

FILL FILL_0_CLKBUF1_insert15 (
);

NAND3X1 _8470_ (
    .A(_1905_),
    .B(_1907_),
    .C(_1906_),
    .Y(_1908_)
);

FILL FILL_0_CLKBUF1_insert16 (
);

OR2X2 _8050_ (
    .A(_1546_),
    .B(_1552_),
    .Y(_1554_)
);

FILL FILL_0_CLKBUF1_insert17 (
);

FILL FILL_0_CLKBUF1_insert18 (
);

FILL FILL_0_CLKBUF1_insert19 (
);

FILL FILL_2__7743_ (
);

FILL FILL_3__12576_ (
);

FILL FILL_2__7323_ (
);

FILL FILL_1__13190_ (
);

FILL FILL_2__11989_ (
);

FILL FILL_2__11569_ (
);

FILL FILL_2__11149_ (
);

FILL FILL_0__12183_ (
);

FILL FILL_2__12930_ (
);

FILL FILL_0__7989_ (
);

FILL FILL_0__7569_ (
);

INVX1 _9675_ (
    .A(\u_fir_pe3.mul [1]),
    .Y(_3024_)
);

FILL FILL_0__7149_ (
);

AOI21X1 _9255_ (
    .A(_2553_),
    .B(_2557_),
    .C(_2546_),
    .Y(_2614_)
);

FILL FILL_1__11923_ (
);

FILL FILL_1__11503_ (
);

FILL FILL_0__8930_ (
);

FILL FILL_2__8948_ (
);

FILL FILL_0__8510_ (
);

FILL FILL_2__8528_ (
);

FILL FILL_0__10916_ (
);

OAI21X1 _13253_ (
    .A(_6260_),
    .B(_6261_),
    .C(_6275_),
    .Y(_6276_)
);

FILL FILL_1__6945_ (
);

FILL FILL_1__6525_ (
);

FILL FILL_1__12708_ (
);

FILL FILL254550x39750 (
);

FILL FILL_0__9715_ (
);

FILL FILL_3__10642_ (
);

FILL FILL_3__10222_ (
);

FILL FILL_2__8281_ (
);

OAI21X1 _7741_ (
    .A(_1183_),
    .B(_1187_),
    .C(_1185_),
    .Y(_1257_)
);

INVX1 _7321_ (
    .A(_829_),
    .Y(_843_)
);

FILL FILL254250x46950 (
);

NAND2X1 _10798_ (
    .A(_3998_),
    .B(_3994_),
    .Y(_4001_)
);

OAI22X1 _10378_ (
    .A(_3203_),
    .B(_3650_),
    .C(_3651_),
    .D(_3653_),
    .Y(_3654_)
);

FILL FILL_3__11847_ (
);

FILL FILL_1__12881_ (
);

FILL FILL_3__11427_ (
);

FILL FILL_3__11007_ (
);

FILL FILL_1__12041_ (
);

FILL FILL_2__9486_ (
);

FILL FILL_0__11874_ (
);

FILL FILL_2__9066_ (
);

FILL FILL_0__11454_ (
);

FILL FILL_0__11034_ (
);

NAND2X1 _8946_ (
    .A(_2368_),
    .B(_2369_),
    .Y(_2384_[15])
);

NAND3X1 _8526_ (
    .A(_1894_),
    .B(_1958_),
    .C(_1959_),
    .Y(_1964_)
);

DFFPOSX1 _8106_ (
    .D(\Y[1] [6]),
    .CLK(clk_bF$buf16),
    .Q(\u_fir_pe1.rYin [6])
);

FILL FILL_1__7483_ (
);

FILL FILL_1__7063_ (
);

FILL FILL_1__13246_ (
);

AOI22X1 _12944_ (
    .A(vdd),
    .B(\X[6]_5_bF$buf0 ),
    .C(vdd),
    .D(\X[6] [6]),
    .Y(_5981_)
);

FILL FILL_0__12659_ (
);

FILL FILL_3__8350_ (
);

FILL FILL_0__12239_ (
);

NOR2X1 _12524_ (
    .A(_6329_),
    .B(_6319_),
    .Y(_6339_)
);

INVX1 _12104_ (
    .A(_5213_),
    .Y(_5221_)
);

FILL FILL_1__8688_ (
);

FILL FILL_1__8268_ (
);

FILL FILL_3__11180_ (
);

FILL FILL_2__10593_ (
);

FILL FILL_2__10173_ (
);

FILL FILL_3__9135_ (
);

NOR2X1 _13309_ (
    .A(\u_fir_pe7.rYin [13]),
    .B(\u_fir_pe7.mul [13]),
    .Y(_6333_)
);

FILL FILL_0__6593_ (
);

FILL FILL_2__7972_ (
);

FILL FILL_2__7552_ (
);

FILL FILL253050x61350 (
);

FILL FILL_2__7132_ (
);

FILL FILL_2__11798_ (
);

FILL FILL_2__11378_ (
);

FILL FILL_0__7798_ (
);

FILL FILL_0__7378_ (
);

AND2X2 _9484_ (
    .A(_2840_),
    .B(_2833_),
    .Y(_2841_)
);

AND2X2 _9064_ (
    .A(gnd),
    .B(\X[3] [1]),
    .Y(_2426_)
);

FILL FILL_1__11732_ (
);

FILL FILL_1__11312_ (
);

FILL FILL_2__8757_ (
);

FILL FILL_2__8337_ (
);

FILL FILL_0__10305_ (
);

FILL FILL_0__13197_ (
);

AOI22X1 _13062_ (
    .A(\X[6]_5_bF$buf2 ),
    .B(gnd),
    .C(_6056_),
    .D(_6057_),
    .Y(_6097_)
);

FILL FILL_1__6754_ (
);

FILL FILL_2__13104_ (
);

FILL FILL_1__12937_ (
);

FILL FILL_1__12517_ (
);

FILL FILL_0__9944_ (
);

FILL FILL_0__9524_ (
);

FILL FILL_3__7621_ (
);

FILL FILL_0__9104_ (
);

FILL FILL_1__7959_ (
);

FILL FILL_1__7539_ (
);

FILL FILL_3__10451_ (
);

FILL FILL_1__7119_ (
);

FILL FILL_1__8900_ (
);

FILL FILL_3__8826_ (
);

FILL FILL_3__8406_ (
);

NOR2X1 _7970_ (
    .A(_1473_),
    .B(_1472_),
    .Y(_1474_)
);

OAI21X1 _7550_ (
    .A(_1055_),
    .B(_1059_),
    .C(_1062_),
    .Y(_1069_)
);

NOR2X1 _7130_ (
    .A(_713_),
    .B(_712_),
    .Y(_714_)
);

NAND3X1 _10187_ (
    .A(_3410_),
    .B(_3451_),
    .C(_3456_),
    .Y(_3466_)
);

FILL FILL_2__6823_ (
);

FILL FILL_2__6403_ (
);

FILL FILL_1__12690_ (
);

FILL FILL_1__12270_ (
);

FILL FILL_2__10649_ (
);

FILL FILL_2__9295_ (
);

FILL FILL_0__11683_ (
);

FILL FILL_2__10229_ (
);

FILL FILL_0__11263_ (
);

FILL FILL_0__6649_ (
);

INVX1 _8755_ (
    .A(_2187_),
    .Y(_2188_)
);

AOI21X1 _8335_ (
    .A(_1765_),
    .B(_1761_),
    .C(_1746_),
    .Y(_1775_)
);

FILL FILL_1__7292_ (
);

FILL FILL_2__7608_ (
);

FILL FILL_1__13055_ (
);

FILL FILL_0__12888_ (
);

INVX1 _12753_ (
    .A(_5791_),
    .Y(_5792_)
);

FILL FILL_0__12048_ (
);

NOR2X1 _12333_ (
    .A(_5437_),
    .B(_5438_),
    .Y(_5439_)
);

FILL FILL_1__8497_ (
);

FILL FILL_3__9364_ (
);

NOR2X1 _13118_ (
    .A(_6144_),
    .B(_6148_),
    .Y(_6152_)
);

FILL FILL_2__7781_ (
);

FILL FILL_2__7361_ (
);

FILL FILL_3__12194_ (
);

FILL FILL_2__11187_ (
);

OAI21X1 _6821_ (
    .A(_417_),
    .B(_319_),
    .C(_132_),
    .Y(_418_)
);

AOI22X1 _6401_ (
    .A(gnd),
    .B(Xin[0]),
    .C(vdd),
    .D(Xin[1]),
    .Y(_4_)
);

FILL FILL_2_BUFX2_insert80 (
);

FILL FILL_0__7187_ (
);

OAI21X1 _9293_ (
    .A(_2641_),
    .B(_2636_),
    .C(_2643_),
    .Y(_2652_)
);

FILL FILL_2_BUFX2_insert81 (
);

FILL FILL_2_BUFX2_insert82 (
);

FILL FILL_3__10927_ (
);

FILL FILL_2_BUFX2_insert83 (
);

FILL FILL_1__11961_ (
);

FILL FILL_2_BUFX2_insert84 (
);

FILL FILL_1__11541_ (
);

FILL FILL_2_BUFX2_insert85 (
);

FILL FILL_2_BUFX2_insert86 (
);

FILL FILL_1__11121_ (
);

FILL FILL_2_BUFX2_insert87 (
);

FILL FILL_2_BUFX2_insert88 (
);

FILL FILL_2_BUFX2_insert89 (
);

FILL FILL_2__8566_ (
);

FILL FILL_0__10954_ (
);

FILL FILL_2__8146_ (
);

FILL FILL_0__10534_ (
);

FILL FILL_0__10114_ (
);

NOR2X1 _13291_ (
    .A(_6314_),
    .B(_6311_),
    .Y(_6315_)
);

AND2X2 _7606_ (
    .A(vdd),
    .B(\X[1]_5_bF$buf2 ),
    .Y(_1124_)
);

FILL FILL_1__6983_ (
);

FILL FILL_1__6563_ (
);

FILL FILL_2__13333_ (
);

FILL FILL_3__6489_ (
);

FILL FILL_1__12746_ (
);

FILL FILL_1__12326_ (
);

FILL FILL_0__9753_ (
);

FILL FILL_3__7850_ (
);

FILL FILL_0__9333_ (
);

FILL FILL_0__11739_ (
);

DFFPOSX1 _11604_ (
    .D(\X[5] [4]),
    .CLK(clk_bF$buf24),
    .Q(\X[6] [4])
);

FILL FILL_0__11319_ (
);

FILL FILL_1__7768_ (
);

FILL FILL_1__7348_ (
);

FILL FILL_3__10260_ (
);

FILL FILL_3__8635_ (
);

AOI21X1 _12809_ (
    .A(_5847_),
    .B(_5842_),
    .C(_5801_),
    .Y(_5848_)
);

FILL FILL_2__6632_ (
);

FILL FILL_3__11045_ (
);

FILL FILL_2__10878_ (
);

FILL FILL_2__10458_ (
);

FILL FILL_0__11492_ (
);

FILL FILL_2__10038_ (
);

FILL FILL_0__11072_ (
);

FILL FILL_1__9914_ (
);

FILL FILL_0__6878_ (
);

DFFPOSX1 _8984_ (
    .D(\Y[2] [7]),
    .CLK(clk_bF$buf38),
    .Q(\u_fir_pe2.rYin [7])
);

FILL FILL_0__6458_ (
);

NAND2X1 _8564_ (
    .A(_2000_),
    .B(_1997_),
    .Y(_2001_)
);

INVX1 _8144_ (
    .A(_2375_),
    .Y(_2376_)
);

FILL FILL_1__10812_ (
);

FILL FILL_2__7837_ (
);

FILL FILL_2__7417_ (
);

FILL FILL_1__13284_ (
);

AOI21X1 _12982_ (
    .A(_6009_),
    .B(_6005_),
    .C(_5964_),
    .Y(_6019_)
);

FILL FILL_0__12697_ (
);

FILL FILL_0__12277_ (
);

NAND2X1 _12562_ (
    .A(\X[6] [4]),
    .B(gnd),
    .Y(_5604_)
);

OAI22X1 _12142_ (
    .A(_5113_),
    .B(_5194_),
    .C(_5256_),
    .D(_5257_),
    .Y(_5258_)
);

FILL FILL_2__12604_ (
);

AOI21X1 _9769_ (
    .A(_3094_),
    .B(_3109_),
    .C(_3112_),
    .Y(_3113_)
);

AOI21X1 _9349_ (
    .A(_2647_),
    .B(_2644_),
    .C(_2630_),
    .Y(_2707_)
);

FILL FILL_0__8604_ (
);

FILL FILL_3__6701_ (
);

FILL FILL_3__9593_ (
);

DFFPOSX1 _13347_ (
    .D(_6369_[9]),
    .CLK(clk_bF$buf39),
    .Q(\Y[7] [9])
);

FILL FILL_1__6619_ (
);

FILL FILL_2__7590_ (
);

FILL FILL_2__7170_ (
);

FILL FILL_0__9809_ (
);

NAND2X1 _6630_ (
    .A(_227_),
    .B(_228_),
    .Y(_229_)
);

FILL FILL_1__11770_ (
);

FILL FILL_3__10316_ (
);

FILL FILL_1__11350_ (
);

FILL FILL_2__8795_ (
);

FILL FILL_2__8375_ (
);

FILL FILL_0__10763_ (
);

FILL FILL_0__10343_ (
);

INVX1 _7835_ (
    .A(_1349_),
    .Y(_1350_)
);

OAI21X1 _7415_ (
    .A(_899_),
    .B(_934_),
    .C(_893_),
    .Y(_935_)
);

FILL FILL_1__6792_ (
);

FILL FILL_2__13142_ (
);

FILL FILL_1__12975_ (
);

FILL FILL_1__12555_ (
);

FILL FILL_1__12135_ (
);

FILL FILL_0__9982_ (
);

FILL FILL_0__11968_ (
);

FILL FILL_0__9562_ (
);

FILL FILL_0__9142_ (
);

OAI21X1 _11833_ (
    .A(_4951_),
    .B(_4952_),
    .C(_4950_),
    .Y(_4953_)
);

FILL FILL_0__11548_ (
);

NAND2X1 _11413_ (
    .A(_4603_),
    .B(_4602_),
    .Y(_4605_)
);

FILL FILL_0__11128_ (
);

FILL FILL_1__7997_ (
);

FILL FILL_1__7577_ (
);

FILL FILL_1__7157_ (
);

NAND3X1 _12618_ (
    .A(\X[6] [1]),
    .B(gnd),
    .C(_5658_),
    .Y(_5659_)
);

FILL FILL_2__6861_ (
);

FILL FILL_3__11694_ (
);

FILL FILL_2__6441_ (
);

FILL FILL_3__11274_ (
);

FILL FILL_2__10687_ (
);

FILL FILL_2__10267_ (
);

FILL FILL_1__9723_ (
);

FILL FILL_1__9303_ (
);

FILL FILL_3__9229_ (
);

FILL FILL_0__6687_ (
);

OAI21X1 _8793_ (
    .A(_2161_),
    .B(_2211_),
    .C(_2189_),
    .Y(_2224_)
);

NAND3X1 _8373_ (
    .A(_1805_),
    .B(_1811_),
    .C(_1810_),
    .Y(_1812_)
);

FILL FILL_1__10621_ (
);

FILL FILL_1__10201_ (
);

FILL FILL_3__12899_ (
);

FILL FILL_2__7646_ (
);

FILL FILL_3__12059_ (
);

FILL FILL_1__13093_ (
);

OAI21X1 _12791_ (
    .A(_5829_),
    .B(_5824_),
    .C(_5818_),
    .Y(_5830_)
);

FILL FILL_0__12086_ (
);

NOR2X1 _12371_ (
    .A(_5472_),
    .B(_5473_),
    .Y(_5474_)
);

FILL FILL_2__12833_ (
);

FILL FILL_2__12413_ (
);

NAND3X1 _9998_ (
    .A(_3274_),
    .B(_3278_),
    .C(_3276_),
    .Y(_3279_)
);

NAND3X1 _9578_ (
    .A(_2906_),
    .B(_2932_),
    .C(_2928_),
    .Y(_2933_)
);

INVX1 _9158_ (
    .A(_2511_),
    .Y(_2519_)
);

FILL FILL_1__11826_ (
);

FILL FILL_1__11406_ (
);

FILL FILL_0__8833_ (
);

FILL FILL_3__6930_ (
);

FILL FILL_0__8413_ (
);

FILL FILL_0__10819_ (
);

OAI21X1 _13156_ (
    .A(_6170_),
    .B(_6165_),
    .C(_6188_),
    .Y(_6189_)
);

FILL FILL_1__6848_ (
);

FILL FILL_1__6428_ (
);

FILL FILL_0__9618_ (
);

FILL FILL_3__7715_ (
);

FILL FILL_3__10545_ (
);

FILL FILL_0__10992_ (
);

FILL FILL_2__8184_ (
);

FILL FILL_0__10572_ (
);

FILL FILL_0__10152_ (
);

OAI21X1 _7644_ (
    .A(_1153_),
    .B(_1149_),
    .C(_1156_),
    .Y(_1162_)
);

DFFPOSX1 _7224_ (
    .D(Yin[1]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [1])
);

FILL FILL_2__6917_ (
);

FILL FILL_1__12784_ (
);

FILL FILL_1__12364_ (
);

FILL FILL_0__9791_ (
);

FILL FILL_0__9371_ (
);

FILL FILL_2__9389_ (
);

FILL FILL_0__11777_ (
);

INVX1 _11642_ (
    .A(_5482_),
    .Y(_5492_)
);

FILL FILL_0__11357_ (
);

INVX1 _11222_ (
    .A(_4411_),
    .Y(_4419_)
);

OR2X2 _8849_ (
    .A(_2266_),
    .B(_2271_),
    .Y(_2273_)
);

OAI21X1 _8429_ (
    .A(_1867_),
    .B(_1863_),
    .C(_1803_),
    .Y(_1868_)
);

OR2X2 _8009_ (
    .A(_1508_),
    .B(_1512_),
    .Y(_1513_)
);

FILL FILL_1__7386_ (
);

FILL FILL_1__13149_ (
);

FILL FILL_3__8673_ (
);

NOR2X1 _12847_ (
    .A(_6349_),
    .B(_5884_),
    .Y(_5885_)
);

FILL FILL_3__8253_ (
);

AND2X2 _12427_ (
    .A(_5530_),
    .B(_5529_),
    .Y(_5572_[12])
);

NAND3X1 _12007_ (
    .A(_5105_),
    .B(_5120_),
    .C(_5121_),
    .Y(_5125_)
);

FILL FILL_2__6670_ (
);

FILL FILL_2__10496_ (
);

FILL FILL_2__10076_ (
);

FILL FILL_1__9952_ (
);

FILL FILL_1__9532_ (
);

FILL FILL_1__9112_ (
);

FILL FILL_3__9458_ (
);

FILL FILL_0__6496_ (
);

NAND2X1 _8182_ (
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1624_)
);

FILL FILL_1__10850_ (
);

FILL FILL_1__10430_ (
);

FILL FILL_1__10010_ (
);

FILL FILL_2__7875_ (
);

FILL FILL_2__7455_ (
);

FILL FILL_3__12288_ (
);

FILL FILL_2__7035_ (
);

NOR2X1 _12180_ (
    .A(_5275_),
    .B(_5280_),
    .Y(_5295_)
);

NOR2X1 _6915_ (
    .A(_507_),
    .B(_510_),
    .Y(_796_[10])
);

FILL FILL_2__12642_ (
);

FILL FILL_2__12222_ (
);

NAND3X1 _9387_ (
    .A(_2740_),
    .B(_2741_),
    .C(_2708_),
    .Y(_2745_)
);

FILL FILL_1__11215_ (
);

FILL FILL_0__8642_ (
);

FILL FILL_0__8222_ (
);

FILL FILL_0__10628_ (
);

INVX1 _10913_ (
    .A(_4110_),
    .Y(_4114_)
);

FILL FILL_0__10208_ (
);

DFFPOSX1 _13385_ (
    .D(_6375_[7]),
    .CLK(clk_bF$buf2),
    .Q(\u_fir_pe7.mul [7])
);

FILL FILL_2__9601_ (
);

FILL FILL_1__6657_ (
);

FILL FILL_2__13007_ (
);

FILL FILL_3__7944_ (
);

FILL FILL_0__9427_ (
);

FILL FILL_3__7104_ (
);

FILL FILL_3__10774_ (
);

FILL FILL_0__10381_ (
);

FILL FILL_1__8803_ (
);

FILL FILL_3__8729_ (
);

NOR2X1 _7873_ (
    .A(_1386_),
    .B(_1385_),
    .Y(_1387_)
);

NAND3X1 _7453_ (
    .A(_970_),
    .B(_972_),
    .C(_971_),
    .Y(_973_)
);

NAND2X1 _7033_ (
    .A(_624_),
    .B(_588_),
    .Y(_625_)
);

FILL FILL_2__13180_ (
);

FILL FILL_2__6726_ (
);

FILL FILL_1__12593_ (
);

FILL FILL_3__11139_ (
);

FILL FILL_1__12173_ (
);

FILL FILL_2__9198_ (
);

FILL FILL_0__9180_ (
);

AOI21X1 _11871_ (
    .A(_4954_),
    .B(_4958_),
    .C(_4920_),
    .Y(_4990_)
);

NAND2X1 _11451_ (
    .A(_4637_),
    .B(_4632_),
    .Y(_4638_)
);

FILL FILL_0__11166_ (
);

AOI21X1 _11031_ (
    .A(_4229_),
    .B(_4228_),
    .C(_4225_),
    .Y(_4230_)
);

FILL FILL_3__12920_ (
);

FILL FILL_2__11913_ (
);

NAND2X1 _8658_ (
    .A(_2092_),
    .B(_2093_),
    .Y(_2094_)
);

NAND2X1 _8238_ (
    .A(gnd),
    .B(\X[2] [4]),
    .Y(_1679_)
);

FILL FILL_1__7195_ (
);

FILL FILL_1__10906_ (
);

FILL FILL_0__7913_ (
);

NAND3X1 _12656_ (
    .A(_5605_),
    .B(_5692_),
    .C(_5693_),
    .Y(_5697_)
);

FILL FILL_3__8062_ (
);

NOR2X1 _12236_ (
    .A(_5349_),
    .B(_5348_),
    .Y(_5350_)
);

FILL FILL_0__13312_ (
);

FILL FILL_1__9761_ (
);

FILL FILL_1__9341_ (
);

FILL FILL_3__9687_ (
);

FILL FILL_2__7684_ (
);

FILL FILL_2__7264_ (
);

OAI21X1 _6724_ (
    .A(_318_),
    .B(_321_),
    .C(_320_),
    .Y(_322_)
);

FILL FILL_2__12871_ (
);

FILL FILL_2__12451_ (
);

FILL FILL_2__12031_ (
);

NAND3X1 _9196_ (
    .A(gnd),
    .B(\X[3] [3]),
    .C(_2555_),
    .Y(_2556_)
);

FILL FILL_1__11864_ (
);

FILL FILL_1__11444_ (
);

FILL FILL_1__11024_ (
);

FILL FILL_0__8871_ (
);

FILL FILL_2__8889_ (
);

FILL FILL_2__8469_ (
);

FILL FILL_0__8451_ (
);

FILL FILL_0__10857_ (
);

FILL FILL_0__10437_ (
);

DFFPOSX1 _10722_ (
    .D(_3978_[15]),
    .CLK(clk_bF$buf6),
    .Q(\Y[5] [15])
);

FILL FILL_2__8049_ (
);

FILL FILL_0__8031_ (
);

OAI21X1 _10302_ (
    .A(_3578_),
    .B(_3577_),
    .C(_3574_),
    .Y(_3579_)
);

FILL FILL_0__10017_ (
);

OAI21X1 _13194_ (
    .A(_6220_),
    .B(_6221_),
    .C(_6219_),
    .Y(_6222_)
);

FILL FILL_2__9410_ (
);

OAI21X1 _7929_ (
    .A(_1429_),
    .B(_1430_),
    .C(_1434_),
    .Y(_1437_)
);

INVX1 _7509_ (
    .A(_1027_),
    .Y(_1028_)
);

FILL FILL_1__6886_ (
);

FILL FILL_1__6466_ (
);

FILL FILL_2__13236_ (
);

FILL FILL_1__12649_ (
);

FILL FILL_1__12229_ (
);

FILL FILL_0__9656_ (
);

FILL FILL_0__9236_ (
);

INVX1 _11927_ (
    .A(_4949_),
    .Y(_5046_)
);

FILL FILL_3__7333_ (
);

INVX1 _11507_ (
    .A(_4688_),
    .Y(_4691_)
);

FILL FILL_3__10583_ (
);

FILL FILL_3__10163_ (
);

FILL FILL_0__10190_ (
);

FILL FILL_1__8612_ (
);

AOI22X1 _7682_ (
    .A(vdd),
    .B(\X[1]_5_bF$buf2 ),
    .C(vdd),
    .D(\X[1] [6]),
    .Y(_1199_)
);

NOR2X1 _7262_ (
    .A(_1547_),
    .B(_1537_),
    .Y(_1557_)
);

FILL FILL_2__6955_ (
);

FILL FILL_3__11788_ (
);

FILL FILL_2__6535_ (
);

FILL FILL_3__11368_ (
);

NAND3X1 _11680_ (
    .A(_4802_),
    .B(_5568_),
    .C(_4801_),
    .Y(_4803_)
);

FILL FILL_0__11395_ (
);

NOR2X1 _11260_ (
    .A(_4391_),
    .B(_4388_),
    .Y(_4456_)
);

FILL FILL_1__9817_ (
);

FILL FILL_2__11722_ (
);

FILL FILL_2__11302_ (
);

OAI21X1 _8887_ (
    .A(_2306_),
    .B(_2307_),
    .C(_2305_),
    .Y(_2311_)
);

INVX1 _8467_ (
    .A(_1898_),
    .Y(_1905_)
);

NOR2X1 _8047_ (
    .A(\u_fir_pe1.rYin [13]),
    .B(\u_fir_pe1.mul [13]),
    .Y(_1551_)
);

FILL FILL_0__7722_ (
);

FILL FILL_0__7302_ (
);

FILL FILL_1__13187_ (
);

OAI21X1 _12885_ (
    .A(_5914_),
    .B(_5908_),
    .C(_5916_),
    .Y(_5923_)
);

FILL FILL_3__8291_ (
);

DFFPOSX1 _12465_ (
    .D(_5572_[4]),
    .CLK(clk_bF$buf22),
    .Q(_6377_[4])
);

AOI21X1 _12045_ (
    .A(_5079_),
    .B(_5149_),
    .C(_5161_),
    .Y(_5162_)
);

FILL FILL_2__12927_ (
);

FILL FILL_0__13121_ (
);

FILL FILL_1_BUFX2_insert0 (
);

FILL FILL_1_BUFX2_insert1 (
);

FILL FILL_1_BUFX2_insert2 (
);

FILL FILL_1_BUFX2_insert3 (
);

FILL FILL_1_BUFX2_insert4 (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_0__8927_ (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_0__8507_ (
);

FILL FILL_3__6604_ (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

FILL FILL_1__9990_ (
);

FILL FILL_1__9570_ (
);

FILL FILL_1__9150_ (
);

FILL FILL_3__9076_ (
);

FILL FILL_2__7493_ (
);

FILL FILL_2__7073_ (
);

FILL FILL_3__7809_ (
);

NAND2X1 _6953_ (
    .A(_547_),
    .B(_514_),
    .Y(_548_)
);

OAI21X1 _6533_ (
    .A(_710_),
    .B(_132_),
    .C(_77_),
    .Y(_133_)
);

FILL FILL_2__12680_ (
);

FILL FILL_2__12260_ (
);

FILL FILL_3__10639_ (
);

FILL FILL_1__11673_ (
);

FILL FILL_1__11253_ (
);

FILL FILL_2__8698_ (
);

FILL FILL_0__8680_ (
);

FILL FILL_0__8260_ (
);

FILL FILL_2__8278_ (
);

FILL FILL_0__10666_ (
);

NAND3X1 _10951_ (
    .A(_4141_),
    .B(_4148_),
    .C(_4150_),
    .Y(_4151_)
);

AOI21X1 _10531_ (
    .A(_3745_),
    .B(_3747_),
    .C(_3802_),
    .Y(_3803_)
);

FILL FILL_0__10246_ (
);

NAND2X1 _10111_ (
    .A(_3390_),
    .B(_3382_),
    .Y(_3391_)
);

AOI21X1 _7738_ (
    .A(_1169_),
    .B(_1239_),
    .C(_1253_),
    .Y(_1254_)
);

NAND3X1 _7318_ (
    .A(vdd),
    .B(\X[1] [1]),
    .C(_839_),
    .Y(_840_)
);

FILL FILL_1__6695_ (
);

FILL FILL_2__13045_ (
);

FILL FILL_1__12878_ (
);

FILL FILL_1__12458_ (
);

FILL FILL_1__12038_ (
);

FILL FILL_0__9465_ (
);

FILL FILL_3__7562_ (
);

FILL FILL_0__9045_ (
);

NAND2X1 _11736_ (
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_4857_)
);

FILL FILL_3__7142_ (
);

NAND2X1 _11316_ (
    .A(gnd),
    .B(\X[5] [7]),
    .Y(_4511_)
);

FILL FILL_0__12812_ (
);

FILL FILL_1__8841_ (
);

FILL FILL_1__8421_ (
);

FILL FILL_1__8001_ (
);

FILL FILL_3__8767_ (
);

FILL FILL_3__8347_ (
);

INVX1 _7491_ (
    .A(_1009_),
    .Y(_1010_)
);

NOR2X1 _7071_ (
    .A(_655_),
    .B(_656_),
    .Y(_657_)
);

FILL FILL_2__6764_ (
);

FILL FILL_1__9626_ (
);

FILL FILL_1__9206_ (
);

FILL FILL_2__11951_ (
);

FILL FILL_2__11531_ (
);

FILL FILL_2__11111_ (
);

NAND2X1 _8696_ (
    .A(_2130_),
    .B(_2110_),
    .Y(_2131_)
);

NAND3X1 _8276_ (
    .A(_1648_),
    .B(_1705_),
    .C(_1709_),
    .Y(_1717_)
);

FILL FILL_1__10944_ (
);

FILL FILL_1__10524_ (
);

FILL FILL_1__10104_ (
);

FILL FILL_0__7951_ (
);

FILL FILL_2__7969_ (
);

FILL FILL_0__7531_ (
);

FILL FILL_2__7549_ (
);

FILL FILL_2__7129_ (
);

FILL FILL_0__7111_ (
);

OAI22X1 _12694_ (
    .A(_5621_),
    .B(_5732_),
    .C(_5664_),
    .D(_5733_),
    .Y(_5734_)
);

NAND3X1 _12274_ (
    .A(_5360_),
    .B(_5362_),
    .C(_5386_),
    .Y(_5387_)
);

FILL FILL_2__8910_ (
);

FILL FILL_2__12736_ (
);

FILL FILL_2__12316_ (
);

FILL FILL_1__11729_ (
);

FILL FILL_1__11309_ (
);

FILL FILL_0__8736_ (
);

FILL FILL_0__8316_ (
);

FILL FILL_3__6413_ (
);

NAND2X1 _13059_ (
    .A(_6047_),
    .B(_6048_),
    .Y(_6094_)
);

NAND3X1 _6762_ (
    .A(_353_),
    .B(_354_),
    .C(_355_),
    .Y(_360_)
);

FILL FILL_3__10868_ (
);

FILL FILL_1__11482_ (
);

FILL FILL_3__10028_ (
);

FILL FILL_1__11062_ (
);

FILL FILL_0__10895_ (
);

FILL FILL_0__10475_ (
);

DFFPOSX1 _10760_ (
    .D(_3984_[13]),
    .CLK(clk_bF$buf44),
    .Q(\u_fir_pe4.mul [13])
);

AOI21X1 _10340_ (
    .A(_3603_),
    .B(_3610_),
    .C(_3585_),
    .Y(_3617_)
);

FILL FILL_0__10055_ (
);

FILL FILL_2__10802_ (
);

INVX1 _7967_ (
    .A(\u_fir_pe1.mul [6]),
    .Y(_1471_)
);

AOI21X1 _7547_ (
    .A(_1065_),
    .B(_1060_),
    .C(_1019_),
    .Y(_1066_)
);

OAI21X1 _7127_ (
    .A(_709_),
    .B(_706_),
    .C(_708_),
    .Y(_711_)
);

FILL FILL_2__13274_ (
);

FILL FILL_0__6802_ (
);

FILL FILL_1__12687_ (
);

FILL FILL_1__12267_ (
);

FILL FILL_0__9694_ (
);

FILL FILL_3__7791_ (
);

FILL FILL_0__9274_ (
);

INVX1 _11965_ (
    .A(_5082_),
    .Y(_5083_)
);

NOR2X1 _11545_ (
    .A(_4727_),
    .B(_4728_),
    .Y(_4729_)
);

NAND3X1 _11125_ (
    .A(_4315_),
    .B(_4319_),
    .C(_4317_),
    .Y(_4323_)
);

FILL FILL_0__12621_ (
);

FILL FILL_0__12201_ (
);

FILL FILL_1__7289_ (
);

FILL FILL_1__8650_ (
);

FILL FILL_1__8230_ (
);

FILL FILL_3__8576_ (
);

FILL FILL_0__13406_ (
);

FILL FILL_2__6993_ (
);

FILL FILL_2__6573_ (
);

FILL FILL_2__10399_ (
);

FILL FILL_1__9435_ (
);

FILL FILL_1__9015_ (
);

FILL FILL_2__11760_ (
);

FILL FILL_2__11340_ (
);

FILL FILL_0__6399_ (
);

DFFPOSX1 _8085_ (
    .D(_1587_[9]),
    .CLK(clk_bF$buf13),
    .Q(\Y[2] [9])
);

FILL FILL_1__10333_ (
);

FILL FILL_0__7760_ (
);

FILL FILL_2__7778_ (
);

FILL FILL_0__7340_ (
);

FILL FILL_2__7358_ (
);

OAI21X1 _12083_ (
    .A(_5199_),
    .B(_5101_),
    .C(_4914_),
    .Y(_5200_)
);

FILL FILL_3__13132_ (
);

NAND3X1 _6818_ (
    .A(_400_),
    .B(_407_),
    .C(_414_),
    .Y(_415_)
);

FILL FILL_2__12965_ (
);

FILL FILL_2__12545_ (
);

FILL FILL_2__12125_ (
);

FILL FILL_1__11958_ (
);

FILL FILL_1__11538_ (
);

FILL FILL_1__11118_ (
);

FILL FILL_0__8545_ (
);

FILL FILL_3__6642_ (
);

NAND2X1 _10816_ (
    .A(gnd),
    .B(\X[5] [3]),
    .Y(_4018_)
);

AND2X2 _13288_ (
    .A(\u_fir_pe7.rYin [11]),
    .B(\u_fir_pe7.mul [11]),
    .Y(_6312_)
);

FILL FILL_2__9924_ (
);

FILL FILL_2__9504_ (
);

FILL FILL_1__7921_ (
);

FILL FILL_1__7501_ (
);

FILL FILL_3__7427_ (
);

NAND2X1 _6991_ (
    .A(_582_),
    .B(_584_),
    .Y(_585_)
);

OAI21X1 _6571_ (
    .A(_169_),
    .B(_170_),
    .C(_168_),
    .Y(_171_)
);

FILL FILL_3__10257_ (
);

FILL FILL_1__11291_ (
);

FILL FILL_0__10284_ (
);

FILL FILL_1__8706_ (
);

FILL FILL_2__10611_ (
);

NAND3X1 _7776_ (
    .A(_1257_),
    .B(_1291_),
    .C(_1289_),
    .Y(_1292_)
);

NAND3X1 _7356_ (
    .A(\X[1] [1]),
    .B(gnd),
    .C(_876_),
    .Y(_877_)
);

FILL FILL_2__13083_ (
);

FILL FILL_2__6629_ (
);

FILL FILL_0__6611_ (
);

FILL FILL_1__12076_ (
);

FILL FILL_0__9083_ (
);

OAI21X1 _11774_ (
    .A(_4890_),
    .B(_4891_),
    .C(_4851_),
    .Y(_4895_)
);

FILL FILL_0__11489_ (
);

FILL FILL_0__11069_ (
);

INVX1 _11354_ (
    .A(_4547_),
    .Y(_4548_)
);

FILL FILL_2__11816_ (
);

FILL FILL_0__12850_ (
);

FILL FILL_0__12430_ (
);

FILL FILL_0__12010_ (
);

FILL FILL_1__7098_ (
);

FILL FILL_1__10809_ (
);

FILL FILL_0__7816_ (
);

OAI21X1 _9922_ (
    .A(_3966_),
    .B(_3203_),
    .C(_3204_),
    .Y(_3205_)
);

NOR2X1 _9502_ (
    .A(_2406_),
    .B(_2853_),
    .Y(_2858_)
);

NAND3X1 _12979_ (
    .A(_5962_),
    .B(_6010_),
    .C(_6015_),
    .Y(_6016_)
);

FILL FILL_3__8385_ (
);

AOI21X1 _12559_ (
    .A(_5598_),
    .B(_5599_),
    .C(_6365_),
    .Y(_5602_)
);

NAND2X1 _12139_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5255_)
);

FILL FILL_0__13215_ (
);

FILL FILL_2__6382_ (
);

FILL FILL_1__9664_ (
);

FILL FILL_1__9244_ (
);

FILL FILL_1__10982_ (
);

FILL FILL_1__10562_ (
);

FILL FILL_1__10142_ (
);

FILL FILL_2__7587_ (
);

FILL FILL_2__7167_ (
);

INVX1 _6627_ (
    .A(_225_),
    .Y(_226_)
);

FILL FILL_2__12774_ (
);

FILL FILL_2__12354_ (
);

OAI21X1 _9099_ (
    .A(_2420_),
    .B(_2454_),
    .C(_2436_),
    .Y(_2460_)
);

FILL FILL_1__11767_ (
);

FILL FILL_1__11347_ (
);

FILL FILL_0__8774_ (
);

FILL FILL_3__6871_ (
);

FILL FILL_0__8354_ (
);

AND2X2 _10625_ (
    .A(_3847_),
    .B(_3857_),
    .Y(_3889_)
);

NAND3X1 _10205_ (
    .A(_3473_),
    .B(_3476_),
    .C(_3392_),
    .Y(_3483_)
);

INVX1 _13097_ (
    .A(_6131_),
    .Y(_6132_)
);

FILL FILL_2__9733_ (
);

FILL FILL_2__9313_ (
);

FILL FILL_0__11701_ (
);

FILL FILL_1__6789_ (
);

FILL FILL_2__13139_ (
);

FILL FILL_1__7730_ (
);

FILL FILL_1__7310_ (
);

FILL FILL_0__9979_ (
);

FILL FILL_0__9559_ (
);

FILL FILL_3__7656_ (
);

FILL FILL_0__9139_ (
);

INVX1 _6380_ (
    .A(_700_),
    .Y(_710_)
);

FILL FILL_0__12906_ (
);

FILL FILL_3__10486_ (
);

FILL FILL_0__10093_ (
);

FILL FILL_1__8935_ (
);

FILL FILL_1__8515_ (
);

FILL FILL_2__10840_ (
);

FILL FILL_2__10420_ (
);

FILL FILL_2__10000_ (
);

NOR2X1 _7585_ (
    .A(_1567_),
    .B(_1102_),
    .Y(_1103_)
);

AND2X2 _7165_ (
    .A(_748_),
    .B(_747_),
    .Y(_790_[12])
);

FILL FILL_2__6858_ (
);

FILL FILL_0__6840_ (
);

FILL FILL_0__6420_ (
);

FILL FILL_2__6438_ (
);

NOR2X1 _11583_ (
    .A(_4764_),
    .B(_4771_),
    .Y(_4778_[2])
);

FILL FILL_0__11298_ (
);

AOI21X1 _11163_ (
    .A(_4274_),
    .B(_4189_),
    .C(_4360_),
    .Y(_4361_)
);

FILL FILL_3__12632_ (
);

FILL FILL_3__12212_ (
);

FILL FILL_2__11205_ (
);

FILL FILL_1__10618_ (
);

FILL FILL_0__7625_ (
);

NOR2X1 _9731_ (
    .A(_3072_),
    .B(_3073_),
    .Y(_3074_)
);

NAND3X1 _9311_ (
    .A(_2668_),
    .B(_2669_),
    .C(_2667_),
    .Y(_2670_)
);

AOI22X1 _12788_ (
    .A(vdd),
    .B(\X[6] [4]),
    .C(vdd),
    .D(\X[6]_5_bF$buf1 ),
    .Y(_5827_)
);

FILL FILL_3__8194_ (
);

NAND2X1 _12368_ (
    .A(_5467_),
    .B(_5470_),
    .Y(_5572_[7])
);

FILL FILL_3__13417_ (
);

FILL FILL_0__13024_ (
);

FILL FILL_1__9893_ (
);

FILL FILL_1__9473_ (
);

FILL FILL_1__9053_ (
);

FILL FILL_3__9399_ (
);

FILL FILL_1__10791_ (
);

FILL FILL_3_BUFX2_insert1 (
);

FILL FILL_1__10371_ (
);

FILL FILL_3_BUFX2_insert2 (
);

FILL FILL_3_BUFX2_insert4 (
);

FILL FILL_3_BUFX2_insert6 (
);

FILL FILL_2__7396_ (
);

FILL FILL_3_BUFX2_insert8 (
);

NAND2X1 _6856_ (
    .A(_452_),
    .B(_451_),
    .Y(_796_[9])
);

AOI22X1 _6436_ (
    .A(gnd),
    .B(Xin[1]),
    .C(vdd),
    .D(Xin[2]),
    .Y(_38_)
);

FILL FILL_2__12583_ (
);

FILL FILL_2__12163_ (
);

FILL FILL_1__11996_ (
);

FILL FILL_1__11576_ (
);

FILL FILL_1__11156_ (
);

FILL FILL_0__8583_ (
);

FILL FILL_0__10989_ (
);

FILL FILL_0__8163_ (
);

FILL FILL_0__10569_ (
);

NAND2X1 _10854_ (
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4055_)
);

NAND2X1 _10434_ (
    .A(gnd),
    .B(_3662_),
    .Y(_3709_)
);

FILL FILL_0__10149_ (
);

AOI21X1 _10014_ (
    .A(_3216_),
    .B(_3236_),
    .C(_3250_),
    .Y(_3295_)
);

FILL FILL_2__9962_ (
);

FILL FILL_0__11930_ (
);

FILL FILL_2__9542_ (
);

FILL FILL_2__9122_ (
);

FILL FILL_0__11510_ (
);

FILL FILL_1__6598_ (
);

FILL FILL_0__9788_ (
);

FILL FILL_3__7885_ (
);

FILL FILL_0__9368_ (
);

DFFPOSX1 _11639_ (
    .D(_4781_[15]),
    .CLK(clk_bF$buf35),
    .Q(\u_fir_pe5.mul [15])
);

FILL FILL_3__7045_ (
);

NAND3X1 _11219_ (
    .A(_4411_),
    .B(_4415_),
    .C(_4370_),
    .Y(_4416_)
);

FILL FILL_1__13302_ (
);

FILL FILL_0__12715_ (
);

FILL FILL_1__8744_ (
);

FILL FILL_1__8324_ (
);

NAND3X1 _7394_ (
    .A(_823_),
    .B(_910_),
    .C(_911_),
    .Y(_915_)
);

FILL FILL_3__9611_ (
);

FILL FILL_2__6667_ (
);

OR2X2 _11392_ (
    .A(_4557_),
    .B(_4583_),
    .Y(_4585_)
);

FILL FILL_1__9949_ (
);

FILL FILL_1__9529_ (
);

FILL FILL_3__12861_ (
);

FILL FILL_1__9109_ (
);

FILL FILL_3__12441_ (
);

FILL FILL_2__11854_ (
);

FILL FILL_2__11434_ (
);

FILL FILL_2__11014_ (
);

NAND3X1 _8599_ (
    .A(_1976_),
    .B(_2031_),
    .C(_2035_),
    .Y(_2036_)
);

AOI22X1 _8179_ (
    .A(\X[2] [0]),
    .B(vdd),
    .C(vdd),
    .D(\X[2] [4]),
    .Y(_1621_)
);

FILL FILL_1__10847_ (
);

FILL FILL_1__10427_ (
);

FILL FILL_1__10007_ (
);

FILL FILL_0__7854_ (
);

INVX1 _9960_ (
    .A(_3241_),
    .Y(_3242_)
);

FILL FILL_0__7434_ (
);

NOR2X1 _9540_ (
    .A(_2893_),
    .B(_2895_),
    .Y(_2896_)
);

FILL FILL_0__7014_ (
);

OAI21X1 _9120_ (
    .A(_2480_),
    .B(_2406_),
    .C(_2474_),
    .Y(_2481_)
);

OR2X2 _12597_ (
    .A(_5638_),
    .B(_5637_),
    .Y(_5639_)
);

NOR2X1 _12177_ (
    .A(_5289_),
    .B(_5292_),
    .Y(_5578_[10])
);

FILL FILL_2__8813_ (
);

FILL FILL_3__13226_ (
);

FILL FILL_2__12639_ (
);

FILL FILL_2__12219_ (
);

FILL FILL_0__13253_ (
);

FILL FILL_1__6810_ (
);

FILL FILL_0__8639_ (
);

FILL FILL_3__6736_ (
);

FILL FILL_0__8219_ (
);

FILL FILL_1__9282_ (
);

FILL FILL_1__10180_ (
);

INVX1 _6665_ (
    .A(_167_),
    .Y(_264_)
);

FILL FILL_2__12392_ (
);

FILL FILL_1__11385_ (
);

FILL FILL_0__8392_ (
);

FILL FILL_0__10798_ (
);

FILL FILL_0__10378_ (
);

AOI21X1 _10663_ (
    .A(_3923_),
    .B(_3914_),
    .C(_3921_),
    .Y(_3926_)
);

NAND2X1 _10243_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3521_)
);

FILL FILL_3__11712_ (
);

FILL FILL_2__9771_ (
);

FILL FILL_2__10705_ (
);

FILL FILL_2__9351_ (
);

FILL FILL_2__13177_ (
);

FILL FILL_0__6705_ (
);

NOR2X1 _8811_ (
    .A(_2236_),
    .B(_2235_),
    .Y(_2239_)
);

FILL FILL_0__9597_ (
);

FILL FILL_0__9177_ (
);

AOI21X1 _11868_ (
    .A(_4976_),
    .B(_4984_),
    .C(_4987_),
    .Y(_4988_)
);

FILL FILL_3__7274_ (
);

NOR2X1 _11448_ (
    .A(_4633_),
    .B(_4634_),
    .Y(_4635_)
);

AND2X2 _11028_ (
    .A(gnd),
    .B(\X[5]_5_bF$buf3 ),
    .Y(_4227_)
);

FILL FILL_1__13111_ (
);

FILL FILL_0__12944_ (
);

FILL FILL_0__12524_ (
);

FILL FILL_0__12104_ (
);

FILL FILL_1__8553_ (
);

FILL FILL_1__8133_ (
);

FILL FILL_0__13309_ (
);

FILL FILL_2__6896_ (
);

FILL FILL_2__6476_ (
);

FILL FILL254550x140550 (
);

FILL FILL_1__9758_ (
);

FILL FILL_3__12670_ (
);

FILL FILL_1__9338_ (
);

FILL FILL_2__11663_ (
);

FILL FILL_2__11243_ (
);

FILL FILL_1__10656_ (
);

FILL FILL_1__10236_ (
);

FILL FILL_0__7663_ (
);

FILL FILL_2__8622_ (
);

FILL FILL_2__8202_ (
);

FILL FILL_2__12868_ (
);

FILL FILL_2__12448_ (
);

FILL FILL_2__12028_ (
);

FILL FILL_0__13062_ (
);

FILL FILL_0__8868_ (
);

FILL FILL_3__6965_ (
);

FILL FILL_0__8448_ (
);

DFFPOSX1 _10719_ (
    .D(_3978_[12]),
    .CLK(clk_bF$buf18),
    .Q(\Y[5] [12])
);

FILL FILL_0__8028_ (
);

FILL FILL_1__9091_ (
);

FILL FILL_1__12802_ (
);

FILL FILL_2__9827_ (
);

FILL FILL_2__9407_ (
);

FILL FILL_1__7824_ (
);

FILL FILL_1__7404_ (
);

NAND3X1 _6894_ (
    .A(_407_),
    .B(_483_),
    .C(_415_),
    .Y(_490_)
);

NAND2X1 _6474_ (
    .A(Xin[1]),
    .B(gnd),
    .Y(_75_)
);

FILL FILL_1__11194_ (
);

AOI21X1 _10892_ (
    .A(_4088_),
    .B(_4089_),
    .C(_4087_),
    .Y(_4093_)
);

OAI21X1 _10472_ (
    .A(_3699_),
    .B(_3740_),
    .C(_3739_),
    .Y(_3746_)
);

FILL FILL_0__10187_ (
);

INVX2 _10052_ (
    .A(\X[4] [6]),
    .Y(_3332_)
);

FILL FILL_3__11941_ (
);

FILL FILL_1__8609_ (
);

FILL FILL_3__11521_ (
);

FILL FILL_3__11101_ (
);

FILL FILL_2__10934_ (
);

FILL FILL_2__9580_ (
);

FILL FILL_2__10514_ (
);

FILL FILL_2__9160_ (
);

AND2X2 _7679_ (
    .A(_929_),
    .B(_1118_),
    .Y(_1196_)
);

NAND2X1 _7259_ (
    .A(vdd),
    .B(\X[1] [1]),
    .Y(_1528_)
);

FILL FILL_0__6934_ (
);

FILL FILL_0__6514_ (
);

INVX2 _8620_ (
    .A(gnd),
    .Y(_2056_)
);

NAND2X1 _8200_ (
    .A(_1640_),
    .B(_1641_),
    .Y(_1642_)
);

FILL FILL_1__12399_ (
);

NAND2X1 _11677_ (
    .A(_4796_),
    .B(_4799_),
    .Y(_4800_)
);

FILL FILL_3__7083_ (
);

NAND2X1 _11257_ (
    .A(gnd),
    .B(_4383_),
    .Y(_4453_)
);

FILL FILL_3__12726_ (
);

FILL FILL_3__12306_ (
);

FILL FILL_2__11719_ (
);

FILL FILL_0__12753_ (
);

FILL FILL_0__12333_ (
);

FILL FILL_0__7719_ (
);

NOR2X1 _9825_ (
    .A(_3167_),
    .B(_3022_),
    .Y(_3180_[0])
);

NAND3X1 _9405_ (
    .A(_2760_),
    .B(_2761_),
    .C(_2762_),
    .Y(_2763_)
);

FILL FILL_1__8782_ (
);

FILL FILL_1__8362_ (
);

FILL FILL_3__8288_ (
);

FILL FILL_0__13118_ (
);

BUFX2 _13403_ (
    .A(_6377_[1]),
    .Y(Yout[1])
);

FILL FILL_1__9987_ (
);

FILL FILL_1__9567_ (
);

FILL FILL_1__9147_ (
);

FILL FILL_2__11892_ (
);

FILL FILL_2__11472_ (
);

FILL FILL_2__11052_ (
);

FILL FILL_1__10885_ (
);

FILL FILL_1__10465_ (
);

FILL FILL_1__10045_ (
);

FILL FILL_0__7892_ (
);

FILL FILL_0__7472_ (
);

FILL FILL_0__7052_ (
);

FILL FILL_2__8851_ (
);

FILL FILL_2__8431_ (
);

FILL FILL_2__8011_ (
);

FILL FILL_2__12677_ (
);

FILL FILL_2__12257_ (
);

FILL FILL_0__13291_ (
);

FILL FILL_0__8677_ (
);

FILL FILL_0__8257_ (
);

NAND3X1 _10948_ (
    .A(gnd),
    .B(\X[5] [4]),
    .C(_4138_),
    .Y(_4148_)
);

NAND3X1 _10528_ (
    .A(_3772_),
    .B(_3800_),
    .C(_3799_),
    .Y(_3801_)
);

AOI21X1 _10108_ (
    .A(_3370_),
    .B(_3365_),
    .C(_3372_),
    .Y(_3388_)
);

FILL FILL_1__12611_ (
);

FILL FILL_2__9636_ (
);

FILL FILL_2__9216_ (
);

FILL FILL_1__7633_ (
);

FILL FILL_3__7979_ (
);

FILL FILL_3__7139_ (
);

FILL FILL_0__12809_ (
);

FILL FILL_3__8500_ (
);

NAND3X1 _10281_ (
    .A(_3489_),
    .B(_3550_),
    .C(_3545_),
    .Y(_3559_)
);

FILL FILL_1__8838_ (
);

FILL FILL_1__8418_ (
);

FILL FILL_3__11330_ (
);

FILL FILL_2__10323_ (
);

NAND2X1 _7488_ (
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_1007_)
);

NAND2X1 _7068_ (
    .A(_653_),
    .B(_654_),
    .Y(_790_[3])
);

FILL FILL_3__9705_ (
);

FILL FILL_0__6743_ (
);

NOR2X1 _11486_ (
    .A(\u_fir_pe5.rYin [7]),
    .B(\u_fir_pe5.mul [7]),
    .Y(_4669_)
);

AOI21X1 _11066_ (
    .A(_4264_),
    .B(_4259_),
    .C(_4120_),
    .Y(_4265_)
);

FILL FILL_3__12955_ (
);

FILL FILL_2__7702_ (
);

FILL FILL_2__11948_ (
);

FILL FILL_0__12982_ (
);

FILL FILL_2__11528_ (
);

FILL FILL_0__12562_ (
);

FILL FILL_2__11108_ (
);

FILL FILL_0__12142_ (
);

FILL FILL_0__7948_ (
);

FILL FILL_0__7528_ (
);

NAND2X1 _9634_ (
    .A(_2958_),
    .B(_2986_),
    .Y(_2987_)
);

FILL FILL_0__7108_ (
);

NAND3X1 _9214_ (
    .A(_2527_),
    .B(_2568_),
    .C(_2573_),
    .Y(_2574_)
);

FILL FILL_1__8591_ (
);

FILL FILL_1__8171_ (
);

FILL FILL_2__8907_ (
);

NOR2X1 _13212_ (
    .A(_6237_),
    .B(_6236_),
    .Y(_6238_)
);

FILL FILL_1__6904_ (
);

FILL FILL_1__9796_ (
);

FILL FILL_1__9376_ (
);

FILL FILL_2__11281_ (
);

FILL FILL_1__10694_ (
);

FILL FILL_1__10274_ (
);

FILL FILL_2__7299_ (
);

FILL FILL_0__7281_ (
);

FILL FILL_2__8660_ (
);

FILL FILL_2__8240_ (
);

FILL FILL_3__13073_ (
);

OAI21X1 _6759_ (
    .A(_356_),
    .B(_352_),
    .C(_303_),
    .Y(_357_)
);

FILL FILL_2__12066_ (
);

FILL FILL_1__11899_ (
);

NAND2X1 _7700_ (
    .A(_1200_),
    .B(_1210_),
    .Y(_1217_)
);

FILL FILL_1__11479_ (
);

FILL FILL_1__11059_ (
);

FILL FILL_0__8486_ (
);

FILL FILL_3__6583_ (
);

DFFPOSX1 _10757_ (
    .D(_3984_[10]),
    .CLK(clk_bF$buf3),
    .Q(\u_fir_pe4.mul [10])
);

FILL FILL_0__8066_ (
);

NAND3X1 _10337_ (
    .A(_3583_),
    .B(_3611_),
    .C(_3613_),
    .Y(_3614_)
);

FILL FILL_3__11806_ (
);

FILL FILL_1__12840_ (
);

FILL FILL_1__12420_ (
);

FILL FILL_1__12000_ (
);

FILL FILL_2__9445_ (
);

FILL FILL_0__11833_ (
);

FILL FILL_2__9025_ (
);

FILL FILL_0__11413_ (
);

FILL FILL253650x172950 (
);

NOR2X1 _8905_ (
    .A(_2328_),
    .B(_2327_),
    .Y(_2329_)
);

FILL FILL_1__7862_ (
);

FILL FILL_1__7442_ (
);

FILL FILL_1__7022_ (
);

FILL FILL_3__7368_ (
);

FILL FILL_1__13205_ (
);

NAND3X1 _12903_ (
    .A(_5939_),
    .B(_5940_),
    .C(_5938_),
    .Y(_5941_)
);

FILL FILL_0__12618_ (
);

FILL FILL253950x32550 (
);

FILL FILL_3__10198_ (
);

OAI21X1 _10090_ (
    .A(_3368_),
    .B(_3369_),
    .C(_3367_),
    .Y(_3370_)
);

FILL FILL_1__8647_ (
);

FILL FILL_1__8227_ (
);

FILL FILL_2__10972_ (
);

FILL FILL_2__10552_ (
);

FILL FILL_2__10132_ (
);

AOI21X1 _7297_ (
    .A(_816_),
    .B(_817_),
    .C(_1583_),
    .Y(_820_)
);

FILL FILL_3__9514_ (
);

FILL FILL_0__6972_ (
);

FILL FILL_0__6552_ (
);

INVX1 _11295_ (
    .A(_4490_),
    .Y(_4491_)
);

FILL FILL_2__7931_ (
);

FILL FILL_2__7511_ (
);

FILL FILL_2__11757_ (
);

FILL FILL_0__12791_ (
);

FILL FILL_2__11337_ (
);

FILL FILL_0__12371_ (
);

FILL FILL_0__7757_ (
);

DFFPOSX1 _9863_ (
    .D(\Y[3] [9]),
    .CLK(clk_bF$buf17),
    .Q(\u_fir_pe3.rYin [9])
);

FILL FILL_0__7337_ (
);

AOI22X1 _9443_ (
    .A(_2633_),
    .B(_2799_),
    .C(_2725_),
    .D(_2721_),
    .Y(_2800_)
);

NOR2X1 _9023_ (
    .A(_3174_),
    .B(_3173_),
    .Y(_3175_)
);

FILL FILL_2__8716_ (
);

FILL FILL_0__13156_ (
);

AND2X2 _13021_ (
    .A(\X[6]_5_bF$buf2 ),
    .B(gnd),
    .Y(_6057_)
);

FILL FILL_1__6713_ (
);

FILL FILL_3__6639_ (
);

FILL FILL_1__9185_ (
);

FILL FILL_0__9903_ (
);

FILL FILL_2__11090_ (
);

FILL FILL_1__10083_ (
);

FILL FILL_0__7090_ (
);

FILL FILL_1__7918_ (
);

FILL FILL_3__10410_ (
);

OAI21X1 _6988_ (
    .A(_579_),
    .B(_581_),
    .C(_560_),
    .Y(_582_)
);

INVX1 _6568_ (
    .A(_155_),
    .Y(_168_)
);

FILL FILL_2__12295_ (
);

FILL FILL_1__11288_ (
);

FILL FILL_0__8295_ (
);

OAI21X1 _10986_ (
    .A(_4184_),
    .B(_4185_),
    .C(_4183_),
    .Y(_4186_)
);

NAND2X1 _10566_ (
    .A(_3833_),
    .B(_3832_),
    .Y(_3834_)
);

NAND3X1 _10146_ (
    .A(_3413_),
    .B(_3422_),
    .C(_3424_),
    .Y(_3425_)
);

FILL FILL_2__9674_ (
);

FILL FILL_2__10608_ (
);

FILL FILL_2__9254_ (
);

FILL FILL_0__11642_ (
);

FILL FILL_0__11222_ (
);

FILL FILL_0__6608_ (
);

OAI21X1 _8714_ (
    .A(_2098_),
    .B(_2101_),
    .C(_2146_),
    .Y(_2149_)
);

FILL FILL_1__7671_ (
);

FILL FILL_3__7597_ (
);

FILL FILL_3__7177_ (
);

FILL FILL_1__13014_ (
);

FILL FILL_0__12847_ (
);

NAND2X1 _12712_ (
    .A(_5730_),
    .B(_5726_),
    .Y(_5752_)
);

FILL FILL_0__12427_ (
);

FILL FILL_0__12007_ (
);

NAND3X1 _9919_ (
    .A(_3976_),
    .B(_3201_),
    .C(_3197_),
    .Y(_3202_)
);

FILL FILL_1__8876_ (
);

FILL FILL_1__8456_ (
);

FILL FILL_1__8036_ (
);

FILL FILL_2__10781_ (
);

FILL FILL_2__10361_ (
);

FILL FILL_3__9323_ (
);

FILL FILL_0__6781_ (
);

FILL FILL_2__6799_ (
);

FILL FILL_2__6379_ (
);

FILL FILL_3__12993_ (
);

FILL FILL_2__7740_ (
);

FILL FILL_3__12573_ (
);

FILL FILL_2__7320_ (
);

FILL FILL_3__12153_ (
);

FILL FILL_2__11986_ (
);

FILL FILL_2__11566_ (
);

FILL FILL_2__11146_ (
);

FILL FILL_0__12180_ (
);

FILL FILL_1__10979_ (
);

FILL FILL_1__10559_ (
);

FILL FILL_1__10139_ (
);

FILL FILL_0__7986_ (
);

FILL FILL_0__7566_ (
);

INVX1 _9672_ (
    .A(_2415_),
    .Y(_3182_[0])
);

FILL FILL_0__7146_ (
);

NOR2X1 _9252_ (
    .A(_2604_),
    .B(_2606_),
    .Y(_2611_)
);

FILL FILL_1__11920_ (
);

FILL FILL_1__11500_ (
);

FILL FILL_2__8945_ (
);

FILL FILL_2__8525_ (
);

FILL FILL_0__10913_ (
);

NAND2X1 _13250_ (
    .A(_6236_),
    .B(_6248_),
    .Y(_6273_)
);

FILL FILL_1__6942_ (
);

FILL FILL_1__6522_ (
);

FILL FILL_1__12705_ (
);

FILL FILL_0__9712_ (
);

FILL FILL_1__7727_ (
);

FILL FILL_1__7307_ (
);

NAND3X1 _6797_ (
    .A(_392_),
    .B(_388_),
    .C(_393_),
    .Y(_394_)
);

FILL FILL_1__11097_ (
);

NAND3X1 _10795_ (
    .A(_3995_),
    .B(_3997_),
    .C(_3996_),
    .Y(_3998_)
);

NOR3X1 _10375_ (
    .A(_3493_),
    .B(_3320_),
    .C(_3509_),
    .Y(_3651_)
);

FILL FILL_3__11424_ (
);

FILL FILL_2__10837_ (
);

FILL FILL_2__9483_ (
);

FILL FILL_0__11871_ (
);

FILL FILL_2__10417_ (
);

FILL FILL_2__9063_ (
);

FILL FILL_0__11451_ (
);

FILL FILL_0__11031_ (
);

FILL FILL_0__6837_ (
);

INVX1 _8943_ (
    .A(_2366_),
    .Y(_2367_)
);

FILL FILL_0__6417_ (
);

OAI21X1 _8523_ (
    .A(_1960_),
    .B(_1957_),
    .C(_1893_),
    .Y(_1961_)
);

DFFPOSX1 _8103_ (
    .D(\Y[1] [3]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.rYin [3])
);

FILL FILL_1__7480_ (
);

FILL FILL_1__7060_ (
);

FILL FILL_1__13243_ (
);

AND2X2 _12941_ (
    .A(_5711_),
    .B(_5900_),
    .Y(_5978_)
);

FILL FILL_0__12656_ (
);

FILL FILL_0__12236_ (
);

NAND2X1 _12521_ (
    .A(vdd),
    .B(\X[6] [1]),
    .Y(_6310_)
);

OAI21X1 _12101_ (
    .A(_5217_),
    .B(_5216_),
    .C(_5215_),
    .Y(_5218_)
);

OAI21X1 _9728_ (
    .A(_3064_),
    .B(_3065_),
    .C(_3069_),
    .Y(_3071_)
);

AOI21X1 _9308_ (
    .A(_2575_),
    .B(_2573_),
    .C(_2666_),
    .Y(_2667_)
);

FILL FILL_1__8685_ (
);

FILL FILL_1__8265_ (
);

FILL FILL_2__10590_ (
);

FILL FILL_2__10170_ (
);

FILL FILL_3__9972_ (
);

FILL FILL_3__9552_ (
);

FILL FILL_3__9132_ (
);

INVX1 _13306_ (
    .A(\u_fir_pe7.rYin [13]),
    .Y(_6330_)
);

FILL FILL_0__6590_ (
);

FILL FILL_3__12382_ (
);

FILL FILL_2__11795_ (
);

FILL FILL_2__11375_ (
);

FILL FILL_1__10788_ (
);

FILL FILL_1__10368_ (
);

FILL FILL_0__7795_ (
);

FILL FILL_0__7375_ (
);

AOI21X1 _9481_ (
    .A(_2837_),
    .B(_2836_),
    .C(_2829_),
    .Y(_2838_)
);

OAI22X1 _9061_ (
    .A(_2421_),
    .B(_2422_),
    .C(_2391_),
    .D(_2395_),
    .Y(_2423_)
);

FILL FILL_2__8754_ (
);

FILL FILL_2__8334_ (
);

FILL FILL_3__13167_ (
);

FILL FILL_0__10302_ (
);

FILL FILL_0__13194_ (
);

FILL FILL_1__6751_ (
);

FILL FILL_2__13101_ (
);

FILL FILL_3__6677_ (
);

FILL FILL_1__12934_ (
);

FILL FILL_2__9959_ (
);

FILL FILL_0__9941_ (
);

FILL FILL_2__9539_ (
);

FILL FILL_0__9521_ (
);

FILL FILL_0__11927_ (
);

FILL FILL_2__9119_ (
);

FILL FILL_0__9101_ (
);

FILL FILL_0__11507_ (
);

FILL FILL_1__7956_ (
);

FILL FILL_1__7536_ (
);

FILL FILL_1__7116_ (
);

FILL FILL_3__8823_ (
);

INVX1 _10184_ (
    .A(_3365_),
    .Y(_3463_)
);

FILL FILL_2__6820_ (
);

FILL FILL_3__11653_ (
);

FILL FILL_2__6400_ (
);

FILL FILL_2__10646_ (
);

FILL FILL_2__9292_ (
);

FILL FILL_0__11680_ (
);

FILL FILL_2__10226_ (
);

FILL FILL_0__11260_ (
);

FILL FILL_3__9608_ (
);

FILL FILL_0__6646_ (
);

NOR2X1 _8752_ (
    .A(_2154_),
    .B(_2177_),
    .Y(_2185_)
);

INVX1 _8332_ (
    .A(_1690_),
    .Y(_1772_)
);

OAI22X1 _11389_ (
    .A(_4129_),
    .B(_4447_),
    .C(_4290_),
    .D(_4220_),
    .Y(_4582_)
);

FILL FILL_2__7605_ (
);

FILL FILL_3__12018_ (
);

FILL FILL_1__13052_ (
);

FILL FILL_0__12885_ (
);

NAND2X1 _12750_ (
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5789_)
);

FILL FILL_0__12045_ (
);

NAND2X1 _12330_ (
    .A(_5435_),
    .B(_5436_),
    .Y(_5572_[3])
);

NAND3X1 _9957_ (
    .A(_3228_),
    .B(_3232_),
    .C(_3234_),
    .Y(_3239_)
);

AOI21X1 _9537_ (
    .A(_2886_),
    .B(_2892_),
    .C(_2850_),
    .Y(_2893_)
);

AND2X2 _9117_ (
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_2478_)
);

FILL FILL_1__8494_ (
);

FILL FILL_1__8074_ (
);

FILL FILL_3__9781_ (
);

OR2X2 _13115_ (
    .A(_6148_),
    .B(_6144_),
    .Y(_6149_)
);

FILL FILL_1__6807_ (
);

FILL FILL_1__9699_ (
);

FILL FILL_1__9279_ (
);

FILL FILL_2__11184_ (
);

FILL FILL_1__10597_ (
);

FILL FILL_1__10177_ (
);

FILL FILL_0__7184_ (
);

AOI21X1 _9290_ (
    .A(_2642_),
    .B(_2648_),
    .C(_2629_),
    .Y(_2649_)
);

FILL FILL_3__10924_ (
);

FILL FILL_3__10504_ (
);

FILL FILL_2__8563_ (
);

FILL FILL_0__10951_ (
);

FILL FILL_3__13396_ (
);

FILL FILL_2__8143_ (
);

FILL FILL_0__10531_ (
);

FILL FILL_0__10111_ (
);

FILL FILL_2__12389_ (
);

NAND2X1 _7603_ (
    .A(gnd),
    .B(\X[1] [7]),
    .Y(_1121_)
);

FILL FILL_1__6980_ (
);

FILL FILL_1__6560_ (
);

FILL FILL_2__13330_ (
);

FILL FILL_0__8389_ (
);

FILL FILL_1__12743_ (
);

FILL FILL_1__12323_ (
);

FILL FILL_0__9750_ (
);

FILL FILL_2__9768_ (
);

FILL FILL_2__9348_ (
);

FILL FILL_0__9330_ (
);

FILL FILL_0__11736_ (
);

DFFPOSX1 _11601_ (
    .D(\X[5] [1]),
    .CLK(clk_bF$buf24),
    .Q(\X[6] [1])
);

FILL FILL_0__11316_ (
);

NOR2X1 _8808_ (
    .A(\u_fir_pe2.rYin [2]),
    .B(\u_fir_pe2.mul [2]),
    .Y(_2236_)
);

FILL FILL_1__7765_ (
);

FILL FILL_1__7345_ (
);

FILL FILL_1__13108_ (
);

NAND3X1 _12806_ (
    .A(_5839_),
    .B(_5838_),
    .C(_5840_),
    .Y(_5845_)
);

FILL FILL_3__8212_ (
);

FILL FILL_3__11882_ (
);

FILL FILL_3__11462_ (
);

FILL FILL_3__11042_ (
);

FILL FILL_2__10875_ (
);

FILL FILL_2__10455_ (
);

FILL FILL_2__10035_ (
);

FILL FILL_1__9911_ (
);

FILL FILL_0__6875_ (
);

DFFPOSX1 _8981_ (
    .D(\Y[2] [4]),
    .CLK(clk_bF$buf44),
    .Q(\u_fir_pe2.rYin [4])
);

FILL FILL_0__6455_ (
);

AOI22X1 _8561_ (
    .A(vdd),
    .B(\X[2] [6]),
    .C(gnd),
    .D(\X[2] [7]),
    .Y(_1998_)
);

INVX2 _8141_ (
    .A(vdd),
    .Y(_2372_)
);

NAND2X1 _11198_ (
    .A(gnd),
    .B(\X[5] [7]),
    .Y(_4395_)
);

FILL FILL_2__7834_ (
);

FILL FILL_3__12667_ (
);

FILL FILL_2__7414_ (
);

FILL FILL_3__12247_ (
);

FILL FILL_1__13281_ (
);

FILL FILL_0__12694_ (
);

FILL FILL_0__12274_ (
);

FILL FILL_2__12601_ (
);

NOR2X1 _9766_ (
    .A(_3106_),
    .B(_3100_),
    .Y(_3109_)
);

NAND2X1 _9346_ (
    .A(_2697_),
    .B(_2698_),
    .Y(_2704_)
);

FILL FILL_2__8619_ (
);

FILL FILL_0__8601_ (
);

FILL FILL_3__9170_ (
);

FILL FILL_0__13059_ (
);

DFFPOSX1 _13344_ (
    .D(_6369_[6]),
    .CLK(clk_bF$buf46),
    .Q(\Y[7] [6])
);

FILL FILL_1__6616_ (
);

FILL FILL_1__9088_ (
);

FILL FILL_0__9806_ (
);

FILL FILL_3__7903_ (
);

FILL FILL_2__8792_ (
);

FILL FILL_2__8372_ (
);

FILL FILL_0__10340_ (
);

FILL FILL_2__12198_ (
);

OAI21X1 _7832_ (
    .A(_1293_),
    .B(_1346_),
    .C(_1289_),
    .Y(_1347_)
);

NAND2X1 _7412_ (
    .A(_928_),
    .B(_930_),
    .Y(_932_)
);

FILL FILL_0__8198_ (
);

NAND3X1 _10889_ (
    .A(_4087_),
    .B(_4089_),
    .C(_4088_),
    .Y(_4090_)
);

NAND2X1 _10469_ (
    .A(_3742_),
    .B(_3743_),
    .Y(_3984_[11])
);

AND2X2 _10049_ (
    .A(\X[4] [2]),
    .B(gnd),
    .Y(_3329_)
);

FILL FILL_1__12972_ (
);

FILL FILL_3__11518_ (
);

FILL FILL_1__12552_ (
);

FILL FILL_1__12132_ (
);

FILL FILL_2__9997_ (
);

FILL FILL_0__11965_ (
);

FILL FILL_2__9577_ (
);

FILL FILL_2__9157_ (
);

INVX1 _11830_ (
    .A(_4937_),
    .Y(_4950_)
);

FILL FILL_0__11545_ (
);

OAI21X1 _11410_ (
    .A(_4579_),
    .B(_4586_),
    .C(_4585_),
    .Y(_4602_)
);

FILL FILL_0__11125_ (
);

OAI21X1 _8617_ (
    .A(_2032_),
    .B(_2034_),
    .C(_2025_),
    .Y(_2053_)
);

FILL FILL_1__7994_ (
);

FILL FILL_1__7574_ (
);

FILL FILL_1__7154_ (
);

FILL FILL_1__13337_ (
);

FILL FILL_3__8441_ (
);

NAND3X1 _12615_ (
    .A(_5655_),
    .B(_5650_),
    .C(_5652_),
    .Y(_5656_)
);

FILL FILL_3__8021_ (
);

FILL FILL_1__8779_ (
);

FILL FILL_1__8359_ (
);

FILL FILL_2__10684_ (
);

FILL FILL_2__10264_ (
);

FILL FILL_1__9720_ (
);

FILL FILL_1__9300_ (
);

FILL FILL_3__9646_ (
);

FILL FILL_3__9226_ (
);

FILL FILL_0__6684_ (
);

NAND3X1 _8790_ (
    .A(_2220_),
    .B(_2221_),
    .C(_2219_),
    .Y(_2222_)
);

OAI21X1 _8370_ (
    .A(_1733_),
    .B(_1808_),
    .C(_1737_),
    .Y(_1809_)
);

FILL FILL_3__12896_ (
);

FILL FILL_2__7643_ (
);

FILL FILL_1__13090_ (
);

FILL FILL_2__11889_ (
);

FILL FILL_2__11469_ (
);

FILL FILL_2__11049_ (
);

FILL FILL_0__12083_ (
);

FILL FILL_2__12830_ (
);

FILL FILL_2__12410_ (
);

FILL FILL_0__7889_ (
);

NAND2X1 _9995_ (
    .A(_3224_),
    .B(_3275_),
    .Y(_3276_)
);

FILL FILL_0__7469_ (
);

AOI21X1 _9575_ (
    .A(_2861_),
    .B(_2877_),
    .C(_2929_),
    .Y(_2930_)
);

FILL FILL_0__7049_ (
);

NAND3X1 _9155_ (
    .A(_2514_),
    .B(_2515_),
    .C(_2513_),
    .Y(_2516_)
);

FILL FILL_1__11823_ (
);

FILL FILL_1__11403_ (
);

FILL FILL_2__8848_ (
);

FILL FILL_0__8830_ (
);

FILL FILL_0__8410_ (
);

FILL FILL_2__8428_ (
);

FILL FILL_0__10816_ (
);

FILL FILL_2__8008_ (
);

FILL FILL_0__13288_ (
);

AND2X2 _13153_ (
    .A(_6182_),
    .B(_6181_),
    .Y(_6186_)
);

FILL FILL_1__6845_ (
);

FILL FILL_1__6425_ (
);

FILL FILL_1__12608_ (
);

FILL FILL_0__9615_ (
);

FILL FILL_3__10962_ (
);

FILL FILL_3__10122_ (
);

FILL FILL_2__8181_ (
);

FILL FILL_3__8917_ (
);

NAND3X1 _7641_ (
    .A(_1157_),
    .B(_1158_),
    .C(_1156_),
    .Y(_1159_)
);

DFFPOSX1 _7221_ (
    .D(Xin[6]),
    .CLK(clk_bF$buf1),
    .Q(\X[1] [6])
);

NAND3X1 _10698_ (
    .A(_3955_),
    .B(_3961_),
    .C(_3956_),
    .Y(_3962_)
);

AOI21X1 _10278_ (
    .A(_3466_),
    .B(_3465_),
    .C(_3397_),
    .Y(_3556_)
);

FILL FILL_2__6914_ (
);

FILL FILL_3__11747_ (
);

FILL FILL_1__12781_ (
);

FILL FILL_1__12361_ (
);

FILL FILL_2__9386_ (
);

FILL FILL_0__11774_ (
);

FILL FILL_0__11354_ (
);

NOR2X1 _8846_ (
    .A(\u_fir_pe2.rYin [6]),
    .B(\u_fir_pe2.mul [6]),
    .Y(_2270_)
);

NAND3X1 _8426_ (
    .A(_1818_),
    .B(_1860_),
    .C(_1861_),
    .Y(_1865_)
);

NOR2X1 _8006_ (
    .A(\u_fir_pe1.rYin [9]),
    .B(\u_fir_pe1.mul [9]),
    .Y(_1510_)
);

FILL FILL_1__7383_ (
);

FILL FILL_1__13146_ (
);

FILL FILL_0__12979_ (
);

FILL FILL_3__8670_ (
);

OAI21X1 _12844_ (
    .A(_5801_),
    .B(_5881_),
    .C(_5850_),
    .Y(_5882_)
);

FILL FILL_0__12559_ (
);

FILL FILL_0__12139_ (
);

NOR2X1 _12424_ (
    .A(_5527_),
    .B(_5526_),
    .Y(_5528_)
);

NAND3X1 _12004_ (
    .A(_5120_),
    .B(_5121_),
    .C(_5119_),
    .Y(_5122_)
);

FILL FILL_1__8588_ (
);

FILL FILL_1__8168_ (
);

FILL FILL_3__11080_ (
);

FILL FILL_2__10493_ (
);

FILL FILL_2__10073_ (
);

FILL FILL_3__9455_ (
);

INVX1 _13209_ (
    .A(\u_fir_pe7.mul [4]),
    .Y(_6235_)
);

FILL FILL_0__6493_ (
);

FILL FILL_2__7872_ (
);

FILL FILL_2__7452_ (
);

FILL FILL_2__7032_ (
);

FILL FILL_2__11698_ (
);

FILL FILL_2__11278_ (
);

NAND2X1 _6912_ (
    .A(_377_),
    .B(_450_),
    .Y(_508_)
);

FILL FILL_0__7698_ (
);

FILL FILL_0__7278_ (
);

NAND3X1 _9384_ (
    .A(_2740_),
    .B(_2741_),
    .C(_2739_),
    .Y(_2742_)
);

FILL FILL_1__11212_ (
);

FILL FILL_2__8657_ (
);

FILL FILL_2__8237_ (
);

FILL FILL_0__10625_ (
);

NAND3X1 _10910_ (
    .A(_4105_),
    .B(_4110_),
    .C(_4052_),
    .Y(_4111_)
);

FILL FILL_0__10205_ (
);

FILL FILL_0__13097_ (
);

DFFPOSX1 _13382_ (
    .D(_6374_[4]),
    .CLK(clk_bF$buf27),
    .Q(\u_fir_pe7.mul [4])
);

FILL FILL_1__6654_ (
);

FILL FILL_2__13004_ (
);

FILL FILL_1__12837_ (
);

FILL FILL_1__12417_ (
);

FILL FILL_0__9424_ (
);

FILL FILL_3__7521_ (
);

FILL FILL_1__7859_ (
);

FILL FILL_1__7439_ (
);

FILL FILL_3__10351_ (
);

FILL FILL_1__7019_ (
);

FILL FILL_1__8800_ (
);

FILL FILL_3__8306_ (
);

NAND3X1 _7870_ (
    .A(_1174_),
    .B(_1247_),
    .C(_1353_),
    .Y(_1384_)
);

NAND2X1 _7450_ (
    .A(_948_),
    .B(_944_),
    .Y(_970_)
);

OAI21X1 _7030_ (
    .A(_616_),
    .B(_615_),
    .C(_621_),
    .Y(_622_)
);

AOI21X1 _10087_ (
    .A(_3270_),
    .B(_3288_),
    .C(_3366_),
    .Y(_3367_)
);

FILL FILL_3__11976_ (
);

FILL FILL_2__6723_ (
);

FILL FILL_3__11556_ (
);

FILL FILL_1__12590_ (
);

FILL FILL_3__11136_ (
);

FILL FILL_1__12170_ (
);

FILL FILL_2__10969_ (
);

FILL FILL_2__10549_ (
);

FILL FILL_2__9195_ (
);

FILL FILL_0__11583_ (
);

FILL FILL_2__10129_ (
);

FILL FILL_0__11163_ (
);

FILL FILL_2__11910_ (
);

FILL FILL_0__6969_ (
);

FILL FILL_0__6549_ (
);

NAND2X1 _8655_ (
    .A(_2087_),
    .B(_2055_),
    .Y(_2091_)
);

AND2X2 _8235_ (
    .A(_1671_),
    .B(_1675_),
    .Y(_1676_)
);

FILL FILL_1__7192_ (
);

FILL FILL_1__10903_ (
);

FILL FILL_2__7928_ (
);

FILL FILL_0__7910_ (
);

FILL FILL_2__7508_ (
);

FILL FILL_0__12788_ (
);

NAND3X1 _12653_ (
    .A(_5691_),
    .B(_5692_),
    .C(_5693_),
    .Y(_5694_)
);

FILL FILL_0__12368_ (
);

NOR2X1 _12233_ (
    .A(_4856_),
    .B(_5244_),
    .Y(_5347_)
);

FILL FILL_1__8397_ (
);

FILL FILL254550x25350 (
);

FILL FILL_3__9264_ (
);

AND2X2 _13018_ (
    .A(_6052_),
    .B(_5995_),
    .Y(_6054_)
);

FILL FILL_2__7681_ (
);

FILL FILL_2__7261_ (
);

FILL FILL_3__12094_ (
);

FILL FILL_2__11087_ (
);

INVX1 _6721_ (
    .A(gnd),
    .Y(_319_)
);

FILL FILL254250x32550 (
);

FILL FILL_0__7087_ (
);

NAND3X1 _9193_ (
    .A(_2548_),
    .B(_2552_),
    .C(_2550_),
    .Y(_2553_)
);

FILL FILL_1__11861_ (
);

FILL FILL_1__11441_ (
);

FILL FILL_1__11021_ (
);

FILL FILL_2__8886_ (
);

FILL FILL_2__8466_ (
);

FILL FILL_0__10854_ (
);

FILL FILL_0__10434_ (
);

FILL FILL_2__8046_ (
);

FILL FILL_0__10014_ (
);

OAI21X1 _13191_ (
    .A(_6211_),
    .B(_6212_),
    .C(_6216_),
    .Y(_6219_)
);

INVX1 _7926_ (
    .A(_1434_),
    .Y(_1435_)
);

AND2X2 _7506_ (
    .A(gnd),
    .B(\X[1] [7]),
    .Y(_1025_)
);

FILL FILL_1__6883_ (
);

FILL FILL_1__6463_ (
);

FILL FILL_2__13233_ (
);

FILL FILL_3__6389_ (
);

FILL FILL_1__12646_ (
);

FILL FILL_1__12226_ (
);

FILL FILL_0__9653_ (
);

FILL FILL_3__7750_ (
);

FILL FILL_0__9233_ (
);

OAI21X1 _11924_ (
    .A(_5032_),
    .B(_5027_),
    .C(_5034_),
    .Y(_5043_)
);

NAND2X1 _11504_ (
    .A(_4684_),
    .B(_4687_),
    .Y(_4688_)
);

FILL FILL_0__11219_ (
);

FILL FILL_1__7668_ (
);

FILL FILL_3__10580_ (
);

FILL FILL_3__8535_ (
);

AOI22X1 _12709_ (
    .A(gnd),
    .B(\X[6]_5_bF$buf3 ),
    .C(_5738_),
    .D(_5740_),
    .Y(_5749_)
);

FILL FILL_2__6952_ (
);

FILL FILL_2__6532_ (
);

FILL FILL_3__11365_ (
);

FILL FILL_2__10778_ (
);

FILL FILL_2__10358_ (
);

FILL FILL_0__11392_ (
);

FILL FILL_1__9814_ (
);

FILL FILL_0__6778_ (
);

NOR2X1 _8884_ (
    .A(_2307_),
    .B(_2306_),
    .Y(_2308_)
);

NOR2X1 _8464_ (
    .A(_1900_),
    .B(_1901_),
    .Y(_1902_)
);

INVX1 _8044_ (
    .A(\u_fir_pe1.rYin [13]),
    .Y(_1548_)
);

FILL FILL_2__7737_ (
);

FILL FILL_2__7317_ (
);

FILL FILL_1__13184_ (
);

AOI21X1 _12882_ (
    .A(_5915_),
    .B(_5919_),
    .C(_5901_),
    .Y(_5920_)
);

FILL FILL_0__12597_ (
);

FILL FILL_0__12177_ (
);

DFFPOSX1 _12462_ (
    .D(_5572_[1]),
    .CLK(clk_bF$buf29),
    .Q(_6377_[1])
);

NAND2X1 _12042_ (
    .A(_5159_),
    .B(_5158_),
    .Y(_5160_)
);

FILL FILL_2__12924_ (
);

OAI21X1 _9669_ (
    .A(_3007_),
    .B(_3006_),
    .C(_3018_),
    .Y(_3020_)
);

NAND3X1 _9249_ (
    .A(_2534_),
    .B(_2603_),
    .C(_2538_),
    .Y(_2608_)
);

FILL FILL_1__11917_ (
);

FILL FILL_0__8924_ (
);

FILL FILL_0__8504_ (
);

FILL FILL_3__9493_ (
);

FILL FILL_3__9073_ (
);

INVX1 _13247_ (
    .A(\u_fir_pe7.mul [8]),
    .Y(_6270_)
);

FILL FILL_1__6939_ (
);

FILL FILL_1__6519_ (
);

FILL FILL_2__7490_ (
);

FILL FILL_2__7070_ (
);

FILL FILL_0__9709_ (
);

NAND2X1 _6950_ (
    .A(_539_),
    .B(_536_),
    .Y(_545_)
);

AND2X2 _6530_ (
    .A(_130_),
    .B(_126_),
    .Y(_796_[5])
);

FILL FILL_1__11670_ (
);

FILL FILL_3__10216_ (
);

FILL FILL_1__11250_ (
);

FILL FILL_2__8695_ (
);

FILL FILL_2__8275_ (
);

FILL FILL_0__10663_ (
);

FILL FILL_0__10243_ (
);

NOR2X1 _7735_ (
    .A(_1170_),
    .B(_1250_),
    .Y(_1251_)
);

NAND3X1 _7315_ (
    .A(_831_),
    .B(_836_),
    .C(_834_),
    .Y(_837_)
);

FILL FILL_1__6692_ (
);

FILL FILL_2__13042_ (
);

FILL FILL_1__12875_ (
);

FILL FILL_1__12455_ (
);

FILL FILL_1__12035_ (
);

FILL FILL_0__9462_ (
);

FILL FILL_0__11868_ (
);

FILL FILL_0__9042_ (
);

AND2X2 _11733_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf2 ),
    .Y(_4854_)
);

FILL FILL_0__11448_ (
);

FILL FILL_0__11028_ (
);

NAND3X1 _11313_ (
    .A(_4505_),
    .B(_4506_),
    .C(_4507_),
    .Y(_4508_)
);

FILL FILL_1__7897_ (
);

FILL FILL_1__7477_ (
);

FILL FILL_1__7057_ (
);

FILL FILL_3__8764_ (
);

AOI21X1 _12938_ (
    .A(_5918_),
    .B(_5917_),
    .C(_5902_),
    .Y(_5975_)
);

AND2X2 _12518_ (
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_6279_)
);

FILL FILL_2__6761_ (
);

FILL FILL_2__10587_ (
);

FILL FILL_2__10167_ (
);

FILL FILL_1__9623_ (
);

FILL FILL_1__9203_ (
);

FILL FILL_3__9549_ (
);

FILL FILL_0__6587_ (
);

INVX1 _8693_ (
    .A(_2125_),
    .Y(_2128_)
);

NAND3X1 _8273_ (
    .A(_1710_),
    .B(_1713_),
    .C(_1662_),
    .Y(_1714_)
);

FILL FILL_1__10941_ (
);

FILL FILL_1__10521_ (
);

FILL FILL_1__10101_ (
);

FILL FILL_2__7966_ (
);

FILL FILL_2__7546_ (
);

FILL FILL_2__7126_ (
);

AND2X2 _12691_ (
    .A(_5726_),
    .B(_5730_),
    .Y(_5731_)
);

NAND2X1 _12271_ (
    .A(_5376_),
    .B(_5383_),
    .Y(_5384_)
);

FILL FILL_3__13320_ (
);

FILL FILL_2__12733_ (
);

FILL FILL_2__12313_ (
);

INVX1 _9898_ (
    .A(_3969_),
    .Y(_3970_)
);

AOI21X1 _9478_ (
    .A(_2691_),
    .B(_2756_),
    .C(_2834_),
    .Y(_2835_)
);

INVX1 _9058_ (
    .A(_2419_),
    .Y(_2420_)
);

FILL FILL_1__11726_ (
);

FILL FILL_1__11306_ (
);

FILL FILL_0__8733_ (
);

FILL FILL_3__6830_ (
);

FILL FILL_0__8313_ (
);

FILL FILL_3__6410_ (
);

NAND2X1 _13056_ (
    .A(_6084_),
    .B(_6088_),
    .Y(_6091_)
);

FILL FILL_1__6748_ (
);

FILL FILL_0__9938_ (
);

FILL FILL_0__9518_ (
);

FILL FILL_3__7615_ (
);

FILL FILL_3__10865_ (
);

FILL FILL_3__10445_ (
);

FILL FILL_0__10892_ (
);

FILL FILL_0__10472_ (
);

FILL FILL_0__10052_ (
);

AND2X2 _7964_ (
    .A(_1468_),
    .B(_1467_),
    .Y(_1587_[5])
);

NAND3X1 _7544_ (
    .A(_1057_),
    .B(_1056_),
    .C(_1058_),
    .Y(_1063_)
);

NAND2X1 _7124_ (
    .A(_704_),
    .B(_707_),
    .Y(_790_[8])
);

FILL FILL_2__13271_ (
);

FILL FILL_2__6817_ (
);

FILL FILL_1__12684_ (
);

FILL FILL_1__12264_ (
);

FILL FILL_0__9691_ (
);

FILL FILL_2__9289_ (
);

FILL FILL_0__9271_ (
);

INVX1 _11962_ (
    .A(_5064_),
    .Y(_5080_)
);

FILL FILL_0__11677_ (
);

OAI21X1 _11542_ (
    .A(_4724_),
    .B(_4707_),
    .C(_4723_),
    .Y(_4726_)
);

FILL FILL_0__11257_ (
);

AOI21X1 _11122_ (
    .A(_4317_),
    .B(_4319_),
    .C(_4315_),
    .Y(_4320_)
);

INVX1 _8749_ (
    .A(_2179_),
    .Y(_2183_)
);

NAND3X1 _8329_ (
    .A(_1756_),
    .B(_1760_),
    .C(_1762_),
    .Y(_1769_)
);

FILL FILL_1__7286_ (
);

FILL FILL_1__13049_ (
);

INVX1 _12747_ (
    .A(_5781_),
    .Y(_5786_)
);

FILL FILL_3__8153_ (
);

NOR2X1 _12327_ (
    .A(_5433_),
    .B(_5432_),
    .Y(_5434_)
);

FILL FILL254250x219750 (
);

FILL FILL_0__13403_ (
);

FILL FILL_2__6990_ (
);

FILL FILL_2__6570_ (
);

FILL FILL_2__10396_ (
);

FILL FILL_1__9432_ (
);

FILL FILL_1__9012_ (
);

FILL FILL_0__6396_ (
);

DFFPOSX1 _8082_ (
    .D(_1587_[6]),
    .CLK(clk_bF$buf54),
    .Q(\Y[2] [6])
);

FILL FILL_1__10330_ (
);

FILL FILL_2__7775_ (
);

FILL FILL_2__7355_ (
);

FILL FILL_3__12188_ (
);

NAND3X1 _12080_ (
    .A(_5182_),
    .B(_5189_),
    .C(_5196_),
    .Y(_5197_)
);

NAND2X1 _6815_ (
    .A(gnd),
    .B(Xin[7]),
    .Y(_412_)
);

FILL FILL_2__12962_ (
);

FILL FILL_2__12542_ (
);

FILL FILL_2__12122_ (
);

NOR2X1 _9287_ (
    .A(_2632_),
    .B(_2645_),
    .Y(_2646_)
);

FILL FILL_1__11955_ (
);

FILL FILL_1__11535_ (
);

FILL FILL_1__11115_ (
);

FILL FILL254550x75750 (
);

FILL FILL_0__8542_ (
);

FILL FILL_0__10948_ (
);

FILL FILL_0__10528_ (
);

NAND2X1 _10813_ (
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4015_)
);

FILL FILL_0__10108_ (
);

OAI21X1 _13285_ (
    .A(_6305_),
    .B(_6306_),
    .C(_6301_),
    .Y(_6309_)
);

FILL FILL_2__9921_ (
);

FILL FILL_2__9501_ (
);

FILL FILL_1__6977_ (
);

FILL FILL_1__6557_ (
);

FILL FILL_2__13327_ (
);

FILL FILL_0__9747_ (
);

FILL FILL_3__7844_ (
);

FILL FILL_0__9327_ (
);

FILL FILL_3__7004_ (
);

FILL FILL_3__10674_ (
);

FILL FILL_0__10281_ (
);

FILL FILL_1__8703_ (
);

FILL FILL_3__8629_ (
);

NAND3X1 _7773_ (
    .A(_1284_),
    .B(_1288_),
    .C(_1258_),
    .Y(_1289_)
);

NAND3X1 _7353_ (
    .A(_873_),
    .B(_868_),
    .C(_870_),
    .Y(_874_)
);

FILL FILL_2__13080_ (
);

FILL FILL_2__6626_ (
);

FILL FILL_3__11459_ (
);

FILL FILL_1__12073_ (
);

FILL FILL_0__9080_ (
);

FILL FILL_2__9098_ (
);

OAI21X1 _11771_ (
    .A(_4890_),
    .B(_4891_),
    .C(_4889_),
    .Y(_4892_)
);

FILL FILL_0__11486_ (
);

FILL FILL_0__11066_ (
);

AND2X2 _11351_ (
    .A(_4527_),
    .B(_4522_),
    .Y(_4545_)
);

FILL FILL_1__9908_ (
);

FILL FILL_3__12820_ (
);

FILL FILL_3__12400_ (
);

FILL FILL_2__11813_ (
);

DFFPOSX1 _8978_ (
    .D(\Y[2] [1]),
    .CLK(clk_bF$buf45),
    .Q(\u_fir_pe2.rYin [1])
);

NAND2X1 _8558_ (
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_1995_)
);

AOI22X1 _8138_ (
    .A(\X[2] [0]),
    .B(gnd),
    .C(\X[2] [1]),
    .D(gnd),
    .Y(_2344_)
);

FILL FILL_1__7095_ (
);

FILL FILL_1__10806_ (
);

FILL FILL_0__7813_ (
);

FILL FILL_1__13278_ (
);

INVX1 _12976_ (
    .A(_6005_),
    .Y(_6013_)
);

FILL FILL_3__8382_ (
);

NAND3X1 _12556_ (
    .A(_6361_),
    .B(_5593_),
    .C(_5596_),
    .Y(_5599_)
);

AND2X2 _12136_ (
    .A(_5248_),
    .B(_5251_),
    .Y(_5252_)
);

FILL FILL_0__13212_ (
);

FILL FILL_1__9661_ (
);

FILL FILL_1__9241_ (
);

FILL FILL_3__9587_ (
);

FILL FILL_3__9167_ (
);

FILL FILL_2__7584_ (
);

FILL FILL_2__7164_ (
);

AOI21X1 _6624_ (
    .A(_162_),
    .B(_166_),
    .C(_155_),
    .Y(_223_)
);

FILL FILL_2__12771_ (
);

FILL FILL_2__12351_ (
);

NAND2X1 _9096_ (
    .A(_2457_),
    .B(_2451_),
    .Y(_3186_[4])
);

FILL FILL_1__11764_ (
);

FILL FILL_1__11344_ (
);

FILL FILL_2__8789_ (
);

FILL FILL_0__8771_ (
);

FILL FILL_0__8351_ (
);

FILL FILL_2__8369_ (
);

FILL FILL_0__10337_ (
);

OAI21X1 _10622_ (
    .A(_3869_),
    .B(_3870_),
    .C(_3884_),
    .Y(_3885_)
);

INVX1 _10202_ (
    .A(_3476_),
    .Y(_3481_)
);

OAI21X1 _13094_ (
    .A(_6075_),
    .B(_6128_),
    .C(_6071_),
    .Y(_6129_)
);

FILL FILL_2__9730_ (
);

FILL FILL_2__9310_ (
);

NAND2X1 _7829_ (
    .A(_1339_),
    .B(_1343_),
    .Y(_1344_)
);

NAND2X1 _7409_ (
    .A(gnd),
    .B(\X[1]_5_bF$buf2 ),
    .Y(_929_)
);

FILL FILL_1__6786_ (
);

FILL FILL_2__13136_ (
);

FILL FILL_1__12969_ (
);

FILL FILL_1__12549_ (
);

FILL FILL_1__12129_ (
);

FILL FILL_0__9976_ (
);

FILL FILL_0__9556_ (
);

FILL FILL_0__9136_ (
);

NAND3X1 _11827_ (
    .A(gnd),
    .B(\X[7] [3]),
    .C(_4946_),
    .Y(_4947_)
);

NAND3X1 _11407_ (
    .A(_4567_),
    .B(_4569_),
    .C(_4597_),
    .Y(_4599_)
);

FILL FILL_0__12903_ (
);

FILL FILL_3__10063_ (
);

FILL FILL_0__10090_ (
);

FILL FILL_1__8932_ (
);

FILL FILL_1__8512_ (
);

FILL FILL_3__8858_ (
);

FILL FILL_3__8018_ (
);

OAI21X1 _7582_ (
    .A(_1019_),
    .B(_1099_),
    .C(_1068_),
    .Y(_1100_)
);

NOR2X1 _7162_ (
    .A(_745_),
    .B(_744_),
    .Y(_746_)
);

FILL FILL_2__6855_ (
);

FILL FILL_3__11688_ (
);

FILL FILL_2__6435_ (
);

AOI21X1 _11580_ (
    .A(\X[5] [0]),
    .B(gnd),
    .C(_4685_),
    .Y(_4762_)
);

FILL FILL_0__11295_ (
);

NAND2X1 _11160_ (
    .A(_4357_),
    .B(_4352_),
    .Y(_4358_)
);

FILL FILL_1__9717_ (
);

FILL FILL_2__11202_ (
);

NAND2X1 _8787_ (
    .A(_2218_),
    .B(_2182_),
    .Y(_2219_)
);

NAND2X1 _8367_ (
    .A(\X[2] [1]),
    .B(gnd),
    .Y(_1806_)
);

FILL FILL_1__10615_ (
);

FILL FILL_0__7622_ (
);

FILL FILL_1__13087_ (
);

AOI21X1 _12785_ (
    .A(_5823_),
    .B(_5822_),
    .C(_5819_),
    .Y(_5824_)
);

INVX1 _12365_ (
    .A(_5462_),
    .Y(_5468_)
);

FILL FILL_2__12827_ (
);

FILL FILL_2__12407_ (
);

FILL FILL_0__13021_ (
);

FILL FILL_0__8827_ (
);

FILL FILL_0__8407_ (
);

FILL FILL_3__6504_ (
);

FILL FILL_1__9890_ (
);

FILL FILL_1__9470_ (
);

FILL FILL_1__9050_ (
);

FILL FILL_2__7393_ (
);

FILL FILL_3__7709_ (
);

AND2X2 _6853_ (
    .A(_449_),
    .B(_442_),
    .Y(_450_)
);

AND2X2 _6433_ (
    .A(vdd),
    .B(Xin[1]),
    .Y(_35_)
);

FILL FILL_2__12580_ (
);

FILL FILL_2__12160_ (
);

FILL FILL_3__10959_ (
);

FILL FILL_1__11993_ (
);

FILL FILL_3__10539_ (
);

FILL FILL_1__11573_ (
);

FILL FILL_1__11153_ (
);

FILL FILL_0__8580_ (
);

FILL FILL_2__8598_ (
);

FILL FILL_0__10986_ (
);

FILL FILL_0__8160_ (
);

FILL FILL_2__8178_ (
);

FILL FILL_0__10566_ (
);

NOR2X1 _10851_ (
    .A(_4006_),
    .B(_4043_),
    .Y(_4052_)
);

AOI22X1 _10431_ (
    .A(\X[4]_5_bF$buf0 ),
    .B(gnd),
    .C(_3665_),
    .D(_3666_),
    .Y(_3706_)
);

FILL FILL_0__10146_ (
);

NAND3X1 _10011_ (
    .A(_3283_),
    .B(_3279_),
    .C(_3285_),
    .Y(_3292_)
);

FILL FILL_3__11900_ (
);

AOI21X1 _7638_ (
    .A(_1067_),
    .B(_1069_),
    .C(_1155_),
    .Y(_1156_)
);

DFFPOSX1 _7218_ (
    .D(Xin[3]),
    .CLK(clk_bF$buf41),
    .Q(\X[1] [3])
);

FILL FILL_1__6595_ (
);

FILL FILL_1__12778_ (
);

FILL FILL_1__12358_ (
);

FILL FILL_0__9785_ (
);

FILL FILL_0__9365_ (
);

FILL FILL_3__7462_ (
);

DFFPOSX1 _11636_ (
    .D(_4781_[12]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [12])
);

AOI21X1 _11216_ (
    .A(_4328_),
    .B(_4334_),
    .C(_4409_),
    .Y(_4413_)
);

FILL FILL_0__12712_ (
);

FILL FILL_3__10292_ (
);

FILL FILL_1__8741_ (
);

FILL FILL_1__8321_ (
);

FILL FILL_3__8247_ (
);

NAND3X1 _7391_ (
    .A(_909_),
    .B(_910_),
    .C(_911_),
    .Y(_912_)
);

FILL FILL_2__6664_ (
);

FILL FILL_3__11497_ (
);

FILL FILL_3__11077_ (
);

FILL FILL_1__9946_ (
);

FILL FILL_1__9526_ (
);

FILL FILL_1__9106_ (
);

FILL FILL_2__11851_ (
);

FILL FILL_2__11431_ (
);

FILL FILL_2__11011_ (
);

INVX1 _8596_ (
    .A(_2025_),
    .Y(_2033_)
);

NAND2X1 _8176_ (
    .A(\X[2] [0]),
    .B(vdd),
    .Y(_1618_)
);

FILL FILL_1__10844_ (
);

FILL FILL_1__10424_ (
);

FILL FILL_1__10004_ (
);

FILL FILL_2__7869_ (
);

FILL FILL_0__7851_ (
);

FILL FILL_2__7449_ (
);

FILL FILL_0__7431_ (
);

FILL FILL_0__7011_ (
);

FILL FILL_2__7029_ (
);

OR2X2 _12594_ (
    .A(_5635_),
    .B(_5634_),
    .Y(_5636_)
);

NAND2X1 _12174_ (
    .A(_5159_),
    .B(_5232_),
    .Y(_5290_)
);

FILL FILL_2__8810_ (
);

NOR2X1 _6909_ (
    .A(_502_),
    .B(_504_),
    .Y(_505_)
);

FILL FILL_2__12636_ (
);

FILL FILL_2__12216_ (
);

FILL FILL_0__13250_ (
);

FILL FILL_1__11209_ (
);

FILL FILL_0__8636_ (
);

FILL FILL_3__6733_ (
);

FILL FILL_0__8216_ (
);

NAND3X1 _10907_ (
    .A(_4039_),
    .B(_4096_),
    .C(_4100_),
    .Y(_4108_)
);

DFFPOSX1 _13379_ (
    .D(_6371_[1]),
    .CLK(clk_bF$buf24),
    .Q(\u_fir_pe7.mul [1])
);

FILL FILL_3__7938_ (
);

FILL FILL_3__7518_ (
);

OAI21X1 _6662_ (
    .A(_250_),
    .B(_245_),
    .C(_252_),
    .Y(_261_)
);

FILL FILL_1__11382_ (
);

FILL FILL_0__10795_ (
);

FILL FILL_0__10375_ (
);

NOR2X1 _10660_ (
    .A(_3923_),
    .B(_3920_),
    .Y(_3924_)
);

INVX1 _10240_ (
    .A(_3512_),
    .Y(_3518_)
);

FILL FILL_2__10702_ (
);

OR2X2 _7867_ (
    .A(_1380_),
    .B(_1357_),
    .Y(_1381_)
);

AOI22X1 _7447_ (
    .A(gnd),
    .B(\X[1]_5_bF$buf3 ),
    .C(_956_),
    .D(_958_),
    .Y(_967_)
);

OR2X2 _7027_ (
    .A(_617_),
    .B(_618_),
    .Y(_619_)
);

FILL FILL_2__13174_ (
);

FILL FILL_0__6702_ (
);

FILL FILL_1__12587_ (
);

FILL FILL_1__12167_ (
);

FILL FILL_0__9594_ (
);

FILL FILL_3__7691_ (
);

FILL FILL_0__9174_ (
);

NAND2X1 _11865_ (
    .A(_4984_),
    .B(_4976_),
    .Y(_4985_)
);

AOI21X1 _11445_ (
    .A(_4625_),
    .B(_4630_),
    .C(_4626_),
    .Y(_4632_)
);

OAI21X1 _11025_ (
    .A(_4141_),
    .B(_4145_),
    .C(_4144_),
    .Y(_4224_)
);

FILL FILL_3__12914_ (
);

FILL FILL_2__11907_ (
);

FILL FILL_0__12941_ (
);

FILL FILL_0__12521_ (
);

FILL FILL_0__12101_ (
);

FILL FILL_1__7189_ (
);

FILL FILL_0__7907_ (
);

FILL FILL_1__8550_ (
);

FILL FILL_3__8476_ (
);

FILL FILL_3__8056_ (
);

FILL FILL_0__13306_ (
);

FILL FILL_2__6893_ (
);

FILL FILL_2__6473_ (
);

FILL FILL_2__10299_ (
);

FILL FILL_1__9755_ (
);

FILL FILL_1__9335_ (
);

FILL FILL_2__11660_ (
);

FILL FILL_2__11240_ (
);

FILL FILL_1__10653_ (
);

FILL FILL_1__10233_ (
);

FILL FILL_0__7660_ (
);

FILL FILL_2__7678_ (
);

FILL FILL_2__7258_ (
);

FILL FILL_3__13032_ (
);

AOI21X1 _6718_ (
    .A(_256_),
    .B(_253_),
    .C(_239_),
    .Y(_316_)
);

FILL FILL_2__12865_ (
);

FILL FILL_2__12445_ (
);

FILL FILL_2__12025_ (
);

FILL FILL_1__11858_ (
);

FILL FILL_1__11438_ (
);

FILL FILL_1__11018_ (
);

FILL FILL_0__8865_ (
);

FILL FILL_3__6962_ (
);

FILL FILL_0__8445_ (
);

DFFPOSX1 _10716_ (
    .D(_3978_[9]),
    .CLK(clk_bF$buf57),
    .Q(\Y[5] [9])
);

FILL FILL_0__8025_ (
);

INVX1 _13188_ (
    .A(_6216_),
    .Y(_6217_)
);

FILL FILL_2__9824_ (
);

FILL FILL_2__9404_ (
);

FILL FILL253650x10950 (
);

FILL FILL_1__7821_ (
);

FILL FILL_1__7401_ (
);

NAND3X1 _6891_ (
    .A(_470_),
    .B(_486_),
    .C(_484_),
    .Y(_487_)
);

AND2X2 _6471_ (
    .A(gnd),
    .B(Xin_5_bF$buf1),
    .Y(_72_)
);

FILL FILL_3__10997_ (
);

FILL FILL_3__10157_ (
);

FILL FILL_1__11191_ (
);

FILL FILL_0__10184_ (
);

FILL FILL_1__8606_ (
);

FILL FILL_2__10931_ (
);

FILL FILL_2__10511_ (
);

AOI21X1 _7676_ (
    .A(_1136_),
    .B(_1135_),
    .C(_1120_),
    .Y(_1193_)
);

AND2X2 _7256_ (
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_1497_)
);

FILL FILL_2__6949_ (
);

FILL FILL_0__6931_ (
);

FILL FILL_2__6529_ (
);

FILL FILL_0__6511_ (
);

FILL FILL_1__12396_ (
);

INVX2 _11674_ (
    .A(\X[7] [3]),
    .Y(_4797_)
);

FILL FILL_0__11389_ (
);

FILL FILL_3__7080_ (
);

INVX1 _11254_ (
    .A(_4449_),
    .Y(_4450_)
);

FILL FILL_3__12303_ (
);

FILL FILL_2__11716_ (
);

FILL FILL_0__12750_ (
);

FILL FILL_0__12330_ (
);

FILL FILL_0__7716_ (
);

OAI21X1 _9822_ (
    .A(_3153_),
    .B(_3156_),
    .C(_3163_),
    .Y(_3166_)
);

OAI21X1 _9402_ (
    .A(_2526_),
    .B(_2759_),
    .C(_2673_),
    .Y(_2760_)
);

NAND3X1 _12879_ (
    .A(_5909_),
    .B(_5913_),
    .C(_5911_),
    .Y(_5917_)
);

NOR2X1 _12459_ (
    .A(_5502_),
    .B(_5566_),
    .Y(_5561_)
);

OAI21X1 _12039_ (
    .A(_4984_),
    .B(_5074_),
    .C(_5070_),
    .Y(_5157_)
);

BUFX2 _13400_ (
    .A(_6376_[6]),
    .Y(Xout[6])
);

FILL FILL_0__13115_ (
);

FILL FILL_1__9984_ (
);

FILL FILL_1__9564_ (
);

FILL FILL_1__9144_ (
);

FILL FILL_1__10882_ (
);

FILL FILL_1__10462_ (
);

FILL FILL_1__10042_ (
);

FILL FILL_2__7487_ (
);

FILL FILL_2__7067_ (
);

FILL FILL_3__13261_ (
);

NAND3X1 _6947_ (
    .A(_515_),
    .B(_541_),
    .C(_537_),
    .Y(_542_)
);

INVX1 _6527_ (
    .A(_120_),
    .Y(_128_)
);

FILL FILL_2__12674_ (
);

FILL FILL_2__12254_ (
);

FILL FILL_1__11667_ (
);

FILL FILL_1__11247_ (
);

FILL FILL_0__8674_ (
);

FILL FILL_3__6771_ (
);

FILL FILL_0__8254_ (
);

AOI22X1 _10945_ (
    .A(vdd),
    .B(\X[5] [3]),
    .C(gnd),
    .D(\X[5] [4]),
    .Y(_4145_)
);

OAI21X1 _10525_ (
    .A(_3779_),
    .B(_3774_),
    .C(_3797_),
    .Y(_3798_)
);

INVX1 _10105_ (
    .A(_3294_),
    .Y(_3385_)
);

FILL FILL_2__9633_ (
);

FILL FILL_2__9213_ (
);

FILL FILL_1__6689_ (
);

FILL FILL_2__13039_ (
);

FILL FILL_1__7630_ (
);

FILL FILL_0__9459_ (
);

FILL FILL_3__7556_ (
);

FILL FILL_0__9039_ (
);

FILL FILL_0__12806_ (
);

FILL FILL_3__10386_ (
);

FILL FILL_1__8835_ (
);

FILL FILL_1__8415_ (
);

FILL FILL_2__10320_ (
);

INVX1 _7485_ (
    .A(_999_),
    .Y(_1004_)
);

NOR2X1 _7065_ (
    .A(_651_),
    .B(_650_),
    .Y(_652_)
);

FILL FILL_3__9702_ (
);

FILL FILL_0__6740_ (
);

FILL FILL_2__6758_ (
);

INVX1 _11483_ (
    .A(\u_fir_pe5.rYin [7]),
    .Y(_4666_)
);

FILL FILL_0__11198_ (
);

NAND3X1 _11063_ (
    .A(_4256_),
    .B(_4255_),
    .C(_4257_),
    .Y(_4262_)
);

FILL FILL_3__12532_ (
);

FILL FILL_2__11945_ (
);

FILL FILL_2__11525_ (
);

FILL FILL_2__11105_ (
);

FILL FILL_1__10938_ (
);

FILL FILL_1__10518_ (
);

FILL FILL_0__7945_ (
);

FILL FILL_0__7525_ (
);

OAI21X1 _9631_ (
    .A(_2696_),
    .B(_2983_),
    .C(_2962_),
    .Y(_2984_)
);

FILL FILL_0__7105_ (
);

AOI21X1 _9211_ (
    .A(_2565_),
    .B(_2566_),
    .C(_2564_),
    .Y(_2571_)
);

NAND2X1 _12688_ (
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_5728_)
);

NAND2X1 _12268_ (
    .A(_5380_),
    .B(_5354_),
    .Y(_5381_)
);

FILL FILL_2__8904_ (
);

FILL FILL_1__6901_ (
);

FILL FILL_3__6827_ (
);

FILL FILL_1__9793_ (
);

FILL FILL_1__9373_ (
);

FILL FILL_1__10691_ (
);

FILL FILL_1__10271_ (
);

FILL FILL_2__7296_ (
);

NAND3X1 _6756_ (
    .A(_349_),
    .B(_350_),
    .C(_317_),
    .Y(_354_)
);

FILL FILL_2__12063_ (
);

FILL FILL_1__11896_ (
);

FILL FILL_1__11476_ (
);

FILL FILL_1__11056_ (
);

FILL FILL_0__8483_ (
);

FILL FILL_0__10889_ (
);

FILL FILL_3__6580_ (
);

FILL FILL_0__10469_ (
);

DFFPOSX1 _10754_ (
    .D(_3984_[7]),
    .CLK(clk_bF$buf21),
    .Q(\u_fir_pe4.mul [7])
);

FILL FILL_0__8063_ (
);

NAND3X1 _10334_ (
    .A(_3603_),
    .B(_3610_),
    .C(_3585_),
    .Y(_3611_)
);

FILL FILL_0__10049_ (
);

FILL FILL_3__11803_ (
);

FILL FILL_2__9442_ (
);

FILL FILL_0__11830_ (
);

FILL FILL_2__9022_ (
);

FILL FILL_0__11410_ (
);

FILL FILL_1__6498_ (
);

FILL FILL_2__13268_ (
);

OAI21X1 _8902_ (
    .A(_2318_),
    .B(_2319_),
    .C(_2323_),
    .Y(_2326_)
);

FILL FILL_0__9688_ (
);

FILL FILL_3__7785_ (
);

FILL FILL_0__9268_ (
);

NAND3X1 _11959_ (
    .A(_5067_),
    .B(_5070_),
    .C(_4986_),
    .Y(_5077_)
);

NOR2X1 _11539_ (
    .A(_4721_),
    .B(_4722_),
    .Y(_4775_[11])
);

NAND2X1 _11119_ (
    .A(_4312_),
    .B(_4316_),
    .Y(_4317_)
);

FILL FILL_1__13202_ (
);

AOI21X1 _12900_ (
    .A(_5849_),
    .B(_5851_),
    .C(_5937_),
    .Y(_5938_)
);

FILL FILL_0__12615_ (
);

FILL FILL_1__8644_ (
);

FILL FILL_1__8224_ (
);

NAND3X1 _7294_ (
    .A(_1579_),
    .B(_811_),
    .C(_814_),
    .Y(_817_)
);

FILL FILL_3__9931_ (
);

FILL FILL_2__6987_ (
);

FILL FILL_2__6567_ (
);

NAND2X1 _11292_ (
    .A(_4480_),
    .B(_4486_),
    .Y(_4488_)
);

FILL FILL_3__12761_ (
);

FILL FILL_1__9429_ (
);

FILL FILL_1__9009_ (
);

FILL FILL_3__12341_ (
);

FILL FILL_2__11754_ (
);

FILL FILL_2__11334_ (
);

NAND3X1 _8499_ (
    .A(_1917_),
    .B(_1932_),
    .C(_1933_),
    .Y(_1937_)
);

DFFPOSX1 _8079_ (
    .D(_1587_[3]),
    .CLK(clk_bF$buf43),
    .Q(\Y[2] [3])
);

FILL FILL_1__10327_ (
);

FILL FILL_0__7754_ (
);

DFFPOSX1 _9860_ (
    .D(\Y[3] [6]),
    .CLK(clk_bF$buf53),
    .Q(\u_fir_pe3.rYin [6])
);

FILL FILL_0__7334_ (
);

AOI21X1 _9440_ (
    .A(_2722_),
    .B(_2796_),
    .C(_2795_),
    .Y(_2797_)
);

NAND2X1 _9020_ (
    .A(_3171_),
    .B(_3151_),
    .Y(_3172_)
);

DFFPOSX1 _12497_ (
    .D(\Y[7] [12]),
    .CLK(clk_bF$buf39),
    .Q(\u_fir_pe6.rYin [12])
);

NAND2X1 _12077_ (
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5194_)
);

FILL FILL_2__8713_ (
);

FILL FILL_3__13126_ (
);

FILL FILL_2__12959_ (
);

FILL FILL_2__12539_ (
);

FILL FILL_2__12119_ (
);

FILL FILL_0__13153_ (
);

FILL FILL_1__6710_ (
);

FILL FILL_0__8539_ (
);

FILL FILL_1__9182_ (
);

FILL FILL_0__9900_ (
);

FILL FILL_2__9918_ (
);

FILL FILL_1__10080_ (
);

FILL FILL_1__7915_ (
);

AOI21X1 _6985_ (
    .A(_577_),
    .B(_578_),
    .C(_561_),
    .Y(_579_)
);

NAND3X1 _6565_ (
    .A(gnd),
    .B(Xin[3]),
    .C(_164_),
    .Y(_165_)
);

FILL FILL_2__12292_ (
);

FILL FILL_1__11285_ (
);

FILL FILL_0__8292_ (
);

FILL FILL_0__10698_ (
);

AOI21X1 _10983_ (
    .A(_4011_),
    .B(_4095_),
    .C(_4182_),
    .Y(_4183_)
);

OAI21X1 _10563_ (
    .A(_3829_),
    .B(_3830_),
    .C(_3828_),
    .Y(_3831_)
);

FILL FILL_0__10278_ (
);

OAI21X1 _10143_ (
    .A(_3203_),
    .B(_3421_),
    .C(_3416_),
    .Y(_3422_)
);

FILL FILL_2__9671_ (
);

FILL FILL_2__10605_ (
);

FILL FILL_2__9251_ (
);

FILL FILL_2__13077_ (
);

FILL FILL_0__6605_ (
);

NAND2X1 _8711_ (
    .A(_2142_),
    .B(_2145_),
    .Y(_2146_)
);

FILL FILL_0__9497_ (
);

FILL FILL_0__9077_ (
);

AOI21X1 _11768_ (
    .A(_4810_),
    .B(_4830_),
    .C(_4844_),
    .Y(_4889_)
);

FILL FILL_3__7174_ (
);

NAND3X1 _11348_ (
    .A(_4439_),
    .B(_4541_),
    .C(_4282_),
    .Y(_4542_)
);

FILL FILL_1__13011_ (
);

FILL FILL_0__12844_ (
);

FILL FILL_0__12424_ (
);

FILL FILL_0__12004_ (
);

NAND3X1 _9916_ (
    .A(_3188_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3199_)
);

FILL FILL_1__8873_ (
);

FILL FILL_1__8453_ (
);

FILL FILL_1__8033_ (
);

FILL FILL_3__8799_ (
);

FILL FILL_3__9320_ (
);

FILL FILL_0__13209_ (
);

FILL FILL_2__6796_ (
);

FILL FILL_3__12990_ (
);

FILL FILL_1__9658_ (
);

FILL FILL_1__9238_ (
);

FILL FILL_2__11983_ (
);

FILL FILL_2__11563_ (
);

FILL FILL_2__11143_ (
);

FILL FILL_1__10976_ (
);

FILL FILL_1__10556_ (
);

FILL FILL_1__10136_ (
);

FILL FILL_0__7983_ (
);

FILL FILL_0__7563_ (
);

FILL FILL_0__7143_ (
);

FILL FILL_2__8942_ (
);

FILL FILL_2__8522_ (
);

FILL FILL_0__10910_ (
);

FILL FILL_2__12768_ (
);

FILL FILL_2__12348_ (
);

FILL FILL_0__8768_ (
);

FILL FILL_0__8348_ (
);

FILL FILL_3__6445_ (
);

NAND2X1 _10619_ (
    .A(_3845_),
    .B(_3857_),
    .Y(_3882_)
);

FILL FILL_1__12702_ (
);

FILL FILL_2__9727_ (
);

FILL FILL_2__9307_ (
);

FILL FILL_1__7724_ (
);

FILL FILL_1__7304_ (
);

OAI21X1 _6794_ (
    .A(_390_),
    .B(_389_),
    .C(_386_),
    .Y(_391_)
);

FILL FILL_1__11094_ (
);

INVX1 _10792_ (
    .A(_4725_),
    .Y(_3995_)
);

OAI21X1 _10372_ (
    .A(_3574_),
    .B(_3578_),
    .C(_3576_),
    .Y(_3648_)
);

FILL FILL_0__10087_ (
);

FILL FILL_1__8929_ (
);

FILL FILL_3__11841_ (
);

FILL FILL_1__8509_ (
);

FILL FILL_3__11001_ (
);

FILL FILL_2__10834_ (
);

FILL FILL_2__9480_ (
);

FILL FILL_2__10414_ (
);

FILL FILL_2__9060_ (
);

INVX1 _7999_ (
    .A(_1500_),
    .Y(_1503_)
);

OAI21X1 _7579_ (
    .A(_1007_),
    .B(_1017_),
    .C(_1013_),
    .Y(_1097_)
);

INVX1 _7159_ (
    .A(\u_fir_pe0.mul [12]),
    .Y(_743_)
);

FILL FILL_0__6834_ (
);

NAND2X1 _8940_ (
    .A(\u_fir_pe2.rYin [15]),
    .B(\u_fir_pe2.mul [15]),
    .Y(_2363_)
);

FILL FILL_0__6414_ (
);

NAND3X1 _8520_ (
    .A(_1897_),
    .B(_1954_),
    .C(_1955_),
    .Y(_1958_)
);

FILL FILL_1__12299_ (
);

DFFPOSX1 _8100_ (
    .D(\Y[1] [0]),
    .CLK(clk_bF$buf43),
    .Q(\u_fir_pe1.rYin [0])
);

NAND2X1 _11997_ (
    .A(vdd),
    .B(\X[7] [6]),
    .Y(_5115_)
);

NAND2X1 _11577_ (
    .A(_4759_),
    .B(_4760_),
    .Y(_4775_[15])
);

NAND3X1 _11157_ (
    .A(_4285_),
    .B(_4349_),
    .C(_4350_),
    .Y(_4355_)
);

FILL FILL_3__12626_ (
);

FILL FILL_1__13240_ (
);

FILL FILL_0__12653_ (
);

FILL FILL_0__12233_ (
);

FILL FILL_0__7619_ (
);

NAND2X1 _9725_ (
    .A(_3068_),
    .B(_3063_),
    .Y(_3069_)
);

AOI21X1 _9305_ (
    .A(_2663_),
    .B(_2662_),
    .C(_2661_),
    .Y(_2664_)
);

FILL FILL_1__8682_ (
);

FILL FILL_1__8262_ (
);

FILL FILL_3__8188_ (
);

FILL FILL_0__13018_ (
);

OR2X2 _13303_ (
    .A(_6320_),
    .B(_6325_),
    .Y(_6327_)
);

FILL FILL_1__9887_ (
);

FILL FILL_1__9467_ (
);

FILL FILL_1__9047_ (
);

FILL FILL_2__11792_ (
);

FILL FILL_2__11372_ (
);

FILL FILL_1__10785_ (
);

FILL FILL_1__10365_ (
);

FILL FILL_0__7792_ (
);

FILL FILL_0__7372_ (
);

FILL FILL_2__8751_ (
);

FILL FILL_2__8331_ (
);

FILL FILL_2__12997_ (
);

FILL FILL_2__12577_ (
);

FILL FILL_2__12157_ (
);

FILL FILL_0__13191_ (
);

FILL FILL_0__8577_ (
);

FILL FILL_3__6674_ (
);

FILL FILL_0__8157_ (
);

AOI21X1 _10848_ (
    .A(_4046_),
    .B(_4049_),
    .C(_4040_),
    .Y(_4050_)
);

NAND2X1 _10428_ (
    .A(_3656_),
    .B(_3657_),
    .Y(_3703_)
);

NAND3X1 _10008_ (
    .A(_3284_),
    .B(_3270_),
    .C(_3288_),
    .Y(_3289_)
);

FILL FILL_1__12931_ (
);

FILL FILL_2__9956_ (
);

FILL FILL_2__9536_ (
);

FILL FILL_0__11924_ (
);

FILL FILL_2__9116_ (
);

FILL FILL_0__11504_ (
);

FILL FILL_1__7953_ (
);

FILL FILL_1__7533_ (
);

FILL FILL_1__7113_ (
);

FILL FILL_3__7879_ (
);

FILL FILL_3__7459_ (
);

FILL FILL_3__7039_ (
);

FILL FILL_0__12709_ (
);

FILL FILL_3__8400_ (
);

OAI21X1 _10181_ (
    .A(_3446_),
    .B(_3450_),
    .C(_3453_),
    .Y(_3460_)
);

FILL FILL_1__8738_ (
);

FILL FILL_1__8318_ (
);

FILL FILL_3__11230_ (
);

FILL FILL_2__10643_ (
);

FILL FILL_2__10223_ (
);

INVX1 _7388_ (
    .A(_823_),
    .Y(_909_)
);

FILL FILL_0__6643_ (
);

INVX1 _11386_ (
    .A(_4578_),
    .Y(_4579_)
);

FILL FILL253950x172950 (
);

FILL FILL_3__12855_ (
);

FILL FILL_2__7602_ (
);

FILL FILL_3__12435_ (
);

FILL FILL_3__12015_ (
);

FILL FILL_2__11848_ (
);

FILL FILL_0__12882_ (
);

FILL FILL_2__11428_ (
);

FILL FILL_2__11008_ (
);

FILL FILL_0__12042_ (
);

FILL FILL_0__7848_ (
);

NAND2X1 _9954_ (
    .A(_3234_),
    .B(_3235_),
    .Y(_3236_)
);

FILL FILL_0__7428_ (
);

AND2X2 _9534_ (
    .A(_2878_),
    .B(_2882_),
    .Y(_2890_)
);

FILL FILL_0__7008_ (
);

OAI22X1 _9114_ (
    .A(_3122_),
    .B(_2474_),
    .C(_2424_),
    .D(_2429_),
    .Y(_2475_)
);

FILL FILL_1__8491_ (
);

FILL FILL_1__8071_ (
);

FILL FILL_2__8807_ (
);

FILL FILL_0__13247_ (
);

NOR2X1 _13112_ (
    .A(_5723_),
    .B(_5884_),
    .Y(_6146_)
);

FILL FILL_1__6804_ (
);

FILL FILL_1__9696_ (
);

FILL FILL_1__9276_ (
);

FILL FILL_2__11181_ (
);

FILL FILL_1__10594_ (
);

FILL FILL_1__10174_ (
);

FILL FILL_0__7181_ (
);

FILL FILL_2__8560_ (
);

FILL FILL_2__8140_ (
);

AOI21X1 _6659_ (
    .A(_251_),
    .B(_257_),
    .C(_238_),
    .Y(_258_)
);

FILL FILL_2__12386_ (
);

FILL FILL_1__11799_ (
);

NAND2X1 _7600_ (
    .A(\X[1] [4]),
    .B(gnd),
    .Y(_1118_)
);

FILL FILL_1__11379_ (
);

FILL FILL_0__8386_ (
);

AND2X2 _10657_ (
    .A(\u_fir_pe4.rYin [11]),
    .B(\u_fir_pe4.mul [11]),
    .Y(_3921_)
);

AND2X2 _10237_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf2 ),
    .Y(_3515_)
);

FILL FILL_1__12740_ (
);

FILL FILL_1__12320_ (
);

FILL FILL_2__9765_ (
);

FILL FILL_2__9345_ (
);

FILL FILL_0__11733_ (
);

FILL FILL_0__11313_ (
);

NOR2X1 _8805_ (
    .A(_2233_),
    .B(_2232_),
    .Y(_2384_[1])
);

FILL FILL_1__7762_ (
);

FILL FILL_1__7342_ (
);

FILL FILL_3__7268_ (
);

FILL FILL_1__13105_ (
);

FILL FILL_0__12938_ (
);

OAI21X1 _12803_ (
    .A(_5837_),
    .B(_5841_),
    .C(_5803_),
    .Y(_5842_)
);

FILL FILL_0__12518_ (
);

FILL FILL_3__10098_ (
);

FILL FILL_1__8547_ (
);

FILL FILL_2__10872_ (
);

FILL FILL_2__10452_ (
);

FILL FILL_2__10032_ (
);

NOR2X1 _7197_ (
    .A(_720_),
    .B(_784_),
    .Y(_779_)
);

FILL FILL_3__9414_ (
);

FILL FILL_0__6872_ (
);

FILL FILL_0__6452_ (
);

NAND2X1 _11195_ (
    .A(_4391_),
    .B(_4388_),
    .Y(_4392_)
);

FILL FILL_2__7831_ (
);

FILL FILL_2__7411_ (
);

FILL FILL_3__12244_ (
);

FILL FILL_2__11657_ (
);

FILL FILL_0__12691_ (
);

FILL FILL_2__11237_ (
);

FILL FILL_0__12271_ (
);

FILL FILL_0__7657_ (
);

OR2X2 _9763_ (
    .A(_3102_),
    .B(_3106_),
    .Y(_3107_)
);

OAI21X1 _9343_ (
    .A(_2699_),
    .B(_2700_),
    .C(_2695_),
    .Y(_2701_)
);

FILL FILL_2__8616_ (
);

FILL FILL_0__13056_ (
);

DFFPOSX1 _13341_ (
    .D(_6369_[3]),
    .CLK(clk_bF$buf11),
    .Q(\Y[7] [3])
);

FILL FILL_1__6613_ (
);

FILL FILL_3__6539_ (
);

FILL FILL_1__9085_ (
);

FILL FILL_0__9803_ (
);

FILL FILL_3__7900_ (
);

FILL FILL_1__7818_ (
);

FILL FILL_3__10310_ (
);

NAND2X1 _6888_ (
    .A(_483_),
    .B(_472_),
    .Y(_484_)
);

OAI21X1 _6468_ (
    .A(_29_),
    .B(_63_),
    .C(_45_),
    .Y(_69_)
);

FILL FILL_2__12195_ (
);

FILL FILL_1__11188_ (
);

FILL FILL_0__8195_ (
);

NAND2X1 _10886_ (
    .A(_4066_),
    .B(_4062_),
    .Y(_4087_)
);

INVX1 _10466_ (
    .A(_3740_),
    .Y(_3741_)
);

OAI21X1 _10046_ (
    .A(_3290_),
    .B(_3325_),
    .C(_3284_),
    .Y(_3326_)
);

FILL FILL_3__11935_ (
);

FILL FILL_2__10928_ (
);

FILL FILL_2__9994_ (
);

FILL FILL_2__9574_ (
);

FILL FILL_0__11962_ (
);

FILL FILL_2__10508_ (
);

FILL FILL_2__9154_ (
);

FILL FILL_0__11542_ (
);

FILL FILL_0__11122_ (
);

FILL FILL_0__6928_ (
);

FILL FILL_0__6508_ (
);

AOI21X1 _8614_ (
    .A(_2035_),
    .B(_2031_),
    .C(_1976_),
    .Y(_2050_)
);

FILL FILL_1__7991_ (
);

FILL FILL_1__7571_ (
);

FILL FILL_1__7151_ (
);

FILL FILL_3__7497_ (
);

FILL FILL_1__13334_ (
);

FILL FILL_0__12747_ (
);

INVX2 _12612_ (
    .A(\X[6]_5_bF$buf1 ),
    .Y(_5653_)
);

FILL FILL_0__12327_ (
);

FILL FILL254250x169350 (
);

NAND2X1 _9819_ (
    .A(_3160_),
    .B(_3162_),
    .Y(_3163_)
);

FILL FILL_1__8776_ (
);

FILL FILL_1__8356_ (
);

FILL FILL_2__10681_ (
);

FILL FILL_2__10261_ (
);

FILL FILL_3__9643_ (
);

FILL FILL_2__6699_ (
);

FILL FILL_0__6681_ (
);

FILL FILL_2__7640_ (
);

FILL FILL_3__12053_ (
);

FILL FILL_2__11886_ (
);

FILL FILL_2__11466_ (
);

FILL FILL_2__11046_ (
);

FILL FILL_0__12080_ (
);

FILL FILL_1__10879_ (
);

FILL FILL_1__10459_ (
);

FILL FILL_1__10039_ (
);

FILL FILL_0__7886_ (
);

NAND2X1 _9992_ (
    .A(vdd),
    .B(\X[4] [4]),
    .Y(_3273_)
);

FILL FILL_0__7466_ (
);

AND2X2 _9572_ (
    .A(_2926_),
    .B(_2923_),
    .Y(_2927_)
);

FILL FILL_0__7046_ (
);

NAND3X1 _9152_ (
    .A(_2512_),
    .B(_2445_),
    .C(_2448_),
    .Y(_2513_)
);

FILL FILL_1__11820_ (
);

FILL FILL_1__11400_ (
);

FILL FILL_2__8845_ (
);

FILL FILL_2__8425_ (
);

FILL FILL_0__10813_ (
);

FILL FILL_2__8005_ (
);

FILL FILL_0__13285_ (
);

NAND2X1 _13150_ (
    .A(_6181_),
    .B(_6182_),
    .Y(_6183_)
);

FILL FILL_1__6842_ (
);

FILL FILL_1__6422_ (
);

FILL FILL_3__6768_ (
);

FILL FILL_1__12605_ (
);

FILL FILL_0__9612_ (
);

FILL FILL_1__7627_ (
);

NAND3X1 _6697_ (
    .A(_285_),
    .B(_288_),
    .C(_204_),
    .Y(_295_)
);

OR2X2 _10695_ (
    .A(\u_fir_pe4.rYin [15]),
    .B(\u_fir_pe4.mul [15]),
    .Y(_3959_)
);

OAI21X1 _10275_ (
    .A(_3544_),
    .B(_3540_),
    .C(_3547_),
    .Y(_3553_)
);

FILL FILL_2__6911_ (
);

FILL FILL_3__11324_ (
);

FILL FILL_2__9383_ (
);

FILL FILL_0__11771_ (
);

FILL FILL_2__10317_ (
);

FILL FILL_0__11351_ (
);

FILL FILL_0__6737_ (
);

INVX1 _8843_ (
    .A(\u_fir_pe2.rYin [6]),
    .Y(_2267_)
);

NAND3X1 _8423_ (
    .A(_1860_),
    .B(_1861_),
    .C(_1859_),
    .Y(_1862_)
);

INVX1 _8003_ (
    .A(_1502_),
    .Y(_1506_)
);

FILL FILL_1__7380_ (
);

FILL FILL_3__12949_ (
);

FILL FILL_3__12109_ (
);

FILL FILL_1__13143_ (
);

FILL FILL_0__12976_ (
);

OAI21X1 _12841_ (
    .A(_5789_),
    .B(_5799_),
    .C(_5795_),
    .Y(_5879_)
);

FILL FILL_0__12556_ (
);

FILL FILL_0__12136_ (
);

INVX1 _12421_ (
    .A(\u_fir_pe6.mul [12]),
    .Y(_5525_)
);

AOI21X1 _12001_ (
    .A(_5028_),
    .B(_5031_),
    .C(_5037_),
    .Y(_5119_)
);

NOR2X1 _9628_ (
    .A(_2977_),
    .B(_2981_),
    .Y(_3187_[12])
);

NAND3X1 _9208_ (
    .A(_2563_),
    .B(_2529_),
    .C(_2567_),
    .Y(_2568_)
);

FILL FILL_1__8585_ (
);

FILL FILL_1__8165_ (
);

FILL FILL_2__10490_ (
);

FILL FILL_2__10070_ (
);

FILL FILL_3__9032_ (
);

OR2X2 _13206_ (
    .A(_6226_),
    .B(_6231_),
    .Y(_6233_)
);

FILL FILL_0__6490_ (
);

FILL FILL_3__12282_ (
);

FILL FILL_2__11695_ (
);

FILL FILL_2__11275_ (
);

FILL FILL_1__10688_ (
);

FILL FILL_1__10268_ (
);

FILL FILL_0__7695_ (
);

FILL FILL_0__7275_ (
);

AOI21X1 _9381_ (
    .A(_2650_),
    .B(_2652_),
    .C(_2738_),
    .Y(_2739_)
);

FILL FILL_2__8654_ (
);

FILL FILL_2__8234_ (
);

FILL FILL_0__10622_ (
);

FILL FILL_3__13067_ (
);

FILL FILL_0__10202_ (
);

FILL FILL_0__13094_ (
);

FILL FILL_1__6651_ (
);

FILL FILL_3__6997_ (
);

FILL FILL_2__13001_ (
);

FILL FILL_1__12834_ (
);

FILL FILL_1__12414_ (
);

FILL FILL_0__9421_ (
);

FILL FILL_2__9439_ (
);

FILL FILL_0__11827_ (
);

FILL FILL_2__9019_ (
);

FILL FILL_0__11407_ (
);

FILL FILL_1__7856_ (
);

FILL FILL_1__7436_ (
);

FILL FILL_1__7016_ (
);

FILL FILL_3__8723_ (
);

NAND3X1 _10084_ (
    .A(_3361_),
    .B(_3363_),
    .C(_3362_),
    .Y(_3364_)
);

FILL FILL_2__6720_ (
);

FILL FILL_3__11553_ (
);

FILL FILL_2__10966_ (
);

FILL FILL_2__10546_ (
);

FILL FILL_2__9192_ (
);

FILL FILL_0__11580_ (
);

FILL FILL_2__10126_ (
);

FILL FILL_0__11160_ (
);

FILL FILL_3__9928_ (
);

FILL FILL_3__9508_ (
);

FILL FILL_0__6966_ (
);

FILL FILL_0__6546_ (
);

NAND3X1 _8652_ (
    .A(_2017_),
    .B(_2020_),
    .C(_2087_),
    .Y(_2088_)
);

NAND2X1 _8232_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf1 ),
    .Y(_1673_)
);

FILL FILL_1__10900_ (
);

NAND2X1 _11289_ (
    .A(_4483_),
    .B(_4484_),
    .Y(_4485_)
);

FILL FILL_2__7925_ (
);

FILL FILL_2__7505_ (
);

FILL FILL_3__12338_ (
);

FILL FILL_0__12785_ (
);

INVX1 _12650_ (
    .A(_5605_),
    .Y(_5691_)
);

FILL FILL_0__12365_ (
);

OAI21X1 _12230_ (
    .A(_5312_),
    .B(_5306_),
    .C(_5316_),
    .Y(_5344_)
);

DFFPOSX1 _9857_ (
    .D(\Y[3] [3]),
    .CLK(clk_bF$buf47),
    .Q(\u_fir_pe3.rYin [3])
);

OAI22X1 _9437_ (
    .A(_2645_),
    .B(_2792_),
    .C(_2715_),
    .D(_2793_),
    .Y(_2794_)
);

INVX1 _9017_ (
    .A(\X[3] [2]),
    .Y(_3161_)
);

FILL FILL_1__8394_ (
);

FILL FILL_3__9681_ (
);

FILL FILL_3__9261_ (
);

OAI21X1 _13015_ (
    .A(_5998_),
    .B(_6050_),
    .C(_5986_),
    .Y(_6051_)
);

FILL FILL_1__6707_ (
);

FILL FILL_1__9599_ (
);

FILL FILL_1__9179_ (
);

FILL FILL_2__11084_ (
);

FILL FILL_1__10497_ (
);

FILL FILL_1__10077_ (
);

FILL FILL_0__7084_ (
);

NAND2X1 _9190_ (
    .A(_2478_),
    .B(_2549_),
    .Y(_2550_)
);

FILL FILL_3__10824_ (
);

FILL FILL_3__10404_ (
);

FILL FILL_2__8883_ (
);

FILL FILL_2__8463_ (
);

FILL FILL_0__10851_ (
);

FILL FILL_0__10431_ (
);

FILL FILL_3__13296_ (
);

FILL FILL_2__8043_ (
);

FILL FILL_0__10011_ (
);

FILL FILL_2__12289_ (
);

NOR2X1 _7923_ (
    .A(\u_fir_pe1.rYin [1]),
    .B(\u_fir_pe1.mul [1]),
    .Y(_1432_)
);

NAND2X1 _7503_ (
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_1022_)
);

FILL FILL_1__6880_ (
);

FILL FILL_1__6460_ (
);

FILL FILL_2__13230_ (
);

FILL FILL_0__8289_ (
);

FILL FILL_3__6386_ (
);

FILL FILL_1__12643_ (
);

FILL FILL_1__12223_ (
);

FILL FILL_0__9650_ (
);

FILL FILL_2__9668_ (
);

FILL FILL_0__9230_ (
);

FILL FILL_2__9248_ (
);

AOI21X1 _11921_ (
    .A(_5033_),
    .B(_5039_),
    .C(_5020_),
    .Y(_5040_)
);

AOI21X1 _11501_ (
    .A(_4680_),
    .B(_4683_),
    .C(_4682_),
    .Y(_4684_)
);

FILL FILL_0__11216_ (
);

AOI21X1 _8708_ (
    .A(_2081_),
    .B(_2085_),
    .C(_2055_),
    .Y(_2143_)
);

FILL FILL_1__7665_ (
);

FILL FILL254550x46950 (
);

FILL FILL_1__13008_ (
);

FILL FILL_3__8952_ (
);

NAND3X1 _12706_ (
    .A(_5734_),
    .B(_5745_),
    .C(_5741_),
    .Y(_5746_)
);

FILL FILL_3__11782_ (
);

FILL FILL253350x111750 (
);

FILL FILL_2__10775_ (
);

FILL FILL_2__10355_ (
);

FILL FILL_1__9811_ (
);

FILL FILL_3__9737_ (
);

FILL FILL_0__6775_ (
);

OAI21X1 _8881_ (
    .A(_2303_),
    .B(_2300_),
    .C(_2302_),
    .Y(_2305_)
);

INVX2 _8461_ (
    .A(gnd),
    .Y(_1899_)
);

OR2X2 _8041_ (
    .A(_1538_),
    .B(_1543_),
    .Y(_1545_)
);

INVX1 _11098_ (
    .A(_4289_),
    .Y(_4296_)
);

FILL FILL_2__7734_ (
);

FILL FILL_3__12567_ (
);

FILL FILL_2__7314_ (
);

FILL FILL_1__13181_ (
);

FILL FILL_0__12594_ (
);

FILL FILL_0__12174_ (
);

FILL FILL_2__12921_ (
);

INVX1 _9666_ (
    .A(_3012_),
    .Y(_3018_)
);

AND2X2 _9246_ (
    .A(_2536_),
    .B(_2540_),
    .Y(_2605_)
);

FILL FILL_1__11914_ (
);

FILL FILL253950x104550 (
);

FILL FILL_2__8939_ (
);

FILL FILL_0__8921_ (
);

FILL FILL_0__8501_ (
);

FILL FILL_2__8519_ (
);

FILL FILL_0__10907_ (
);

FILL FILL_3__9490_ (
);

NAND2X1 _13244_ (
    .A(_6266_),
    .B(_6265_),
    .Y(_6267_)
);

FILL FILL_1__6936_ (
);

FILL FILL_1__6516_ (
);

FILL FILL_0__9706_ (
);

FILL FILL_3__10633_ (
);

FILL FILL_3__10213_ (
);

FILL FILL_2__8692_ (
);

FILL FILL_2__8272_ (
);

FILL FILL_0__10660_ (
);

FILL FILL_0__10240_ (
);

FILL FILL_2__12098_ (
);

NAND2X1 _7732_ (
    .A(_1247_),
    .B(_1177_),
    .Y(_1249_)
);

NAND2X1 _7312_ (
    .A(_832_),
    .B(_833_),
    .Y(_834_)
);

NOR2X1 _10789_ (
    .A(_4716_),
    .B(_3987_),
    .Y(_3992_)
);

AOI21X1 _10369_ (
    .A(_3560_),
    .B(_3630_),
    .C(_3644_),
    .Y(_3645_)
);

FILL FILL_3__11838_ (
);

FILL FILL_1__12872_ (
);

FILL FILL_3__11418_ (
);

FILL FILL_1__12452_ (
);

FILL FILL_1__12032_ (
);

FILL FILL_2__9897_ (
);

FILL FILL_2__9477_ (
);

FILL FILL_0__11865_ (
);

FILL FILL_2__9057_ (
);

OAI21X1 _11730_ (
    .A(_4811_),
    .B(_4845_),
    .C(_4827_),
    .Y(_4851_)
);

FILL FILL_0__11445_ (
);

FILL FILL_0__11025_ (
);

NOR2X1 _11310_ (
    .A(_4402_),
    .B(_4447_),
    .Y(_4505_)
);

NOR2X1 _8937_ (
    .A(_2360_),
    .B(_2359_),
    .Y(_2384_[14])
);

NAND3X1 _8517_ (
    .A(_1909_),
    .B(_1940_),
    .C(_1945_),
    .Y(_1955_)
);

FILL FILL_1__7894_ (
);

FILL FILL_1__7474_ (
);

FILL FILL_1__7054_ (
);

FILL FILL_1__13237_ (
);

INVX1 _12935_ (
    .A(_5969_),
    .Y(_5972_)
);

FILL FILL_3__8341_ (
);

DFFPOSX1 _12515_ (
    .D(_5578_[14]),
    .CLK(clk_bF$buf2),
    .Q(\u_fir_pe6.mul [14])
);

FILL FILL_1__8679_ (
);

FILL FILL_1__8259_ (
);

FILL FILL_3__11171_ (
);

FILL FILL_2__10584_ (
);

FILL FILL_2__10164_ (
);

FILL FILL_1__9620_ (
);

FILL FILL_1__9200_ (
);

FILL FILL_3__9966_ (
);

FILL FILL_3__9126_ (
);

FILL FILL_0__6584_ (
);

AOI21X1 _8690_ (
    .A(_2076_),
    .B(_2119_),
    .C(_2122_),
    .Y(_2125_)
);

NAND3X1 _8270_ (
    .A(_1706_),
    .B(_1700_),
    .C(_1704_),
    .Y(_1711_)
);

FILL FILL_2__7963_ (
);

FILL FILL_3__12796_ (
);

FILL FILL_2__7543_ (
);

FILL FILL_3__12376_ (
);

FILL FILL_2__7123_ (
);

FILL FILL_2__11789_ (
);

FILL FILL_2__11369_ (
);

FILL FILL_2__12730_ (
);

FILL FILL_2__12310_ (
);

FILL FILL_0__7789_ (
);

INVX2 _9895_ (
    .A(gnd),
    .Y(_3966_)
);

FILL FILL_0__7369_ (
);

OAI21X1 _9475_ (
    .A(_2831_),
    .B(_2830_),
    .C(_2829_),
    .Y(_2832_)
);

NOR2X1 _9055_ (
    .A(_2415_),
    .B(_2416_),
    .Y(_2417_)
);

FILL FILL_1__11723_ (
);

FILL FILL_1__11303_ (
);

FILL FILL_0__8730_ (
);

FILL FILL_2__8748_ (
);

FILL FILL_0__8310_ (
);

FILL FILL_2__8328_ (
);

FILL FILL_0__13188_ (
);

NOR2X1 _13053_ (
    .A(_6084_),
    .B(_6088_),
    .Y(_6089_)
);

FILL FILL_1__6745_ (
);

FILL FILL_1__12928_ (
);

FILL FILL_0__9935_ (
);

FILL FILL_0__9515_ (
);

FILL FILL_3__7612_ (
);

FILL FILL_3__10022_ (
);

FILL FILL_3__8817_ (
);

NOR2X1 _7961_ (
    .A(_1465_),
    .B(_1464_),
    .Y(_1466_)
);

OAI21X1 _7541_ (
    .A(_1055_),
    .B(_1059_),
    .C(_1021_),
    .Y(_1060_)
);

NOR2X1 _7121_ (
    .A(_693_),
    .B(_692_),
    .Y(_705_)
);

INVX1 _10598_ (
    .A(\u_fir_pe4.mul [6]),
    .Y(_3862_)
);

AOI21X1 _10178_ (
    .A(_3456_),
    .B(_3451_),
    .C(_3410_),
    .Y(_3457_)
);

FILL FILL_2__6814_ (
);

FILL FILL_1__12681_ (
);

FILL FILL_1__12261_ (
);

FILL FILL_2__9286_ (
);

FILL FILL_0__11674_ (
);

FILL FILL_0__11254_ (
);

AOI21X1 _8746_ (
    .A(_2151_),
    .B(_2153_),
    .C(_2179_),
    .Y(_2180_)
);

NAND3X1 _8326_ (
    .A(_1761_),
    .B(_1746_),
    .C(_1765_),
    .Y(_1766_)
);

FILL FILL_1__7283_ (
);

FILL FILL_1__13046_ (
);

FILL FILL_0__12879_ (
);

FILL FILL_3__8570_ (
);

OAI21X1 _12744_ (
    .A(_5708_),
    .B(_5706_),
    .C(_5699_),
    .Y(_5784_)
);

FILL FILL_0__12459_ (
);

FILL FILL_0__12039_ (
);

INVX1 _12324_ (
    .A(\u_fir_pe6.mul [3]),
    .Y(_5431_)
);

FILL FILL_0__13400_ (
);

FILL FILL_1__8488_ (
);

FILL FILL_1__8068_ (
);

FILL FILL_2__10393_ (
);

FILL FILL_3__9355_ (
);

INVX1 _13109_ (
    .A(_6105_),
    .Y(_6143_)
);

FILL FILL_0__6393_ (
);

FILL FILL_2__7772_ (
);

FILL FILL_2__7352_ (
);

FILL FILL_3__12185_ (
);

FILL FILL_2__11178_ (
);

AOI22X1 _6812_ (
    .A(_242_),
    .B(_408_),
    .C(_334_),
    .D(_330_),
    .Y(_409_)
);

FILL FILL_0__7598_ (
);

FILL FILL_0__7178_ (
);

AOI22X1 _9284_ (
    .A(_2478_),
    .B(_2549_),
    .C(_2552_),
    .D(_2548_),
    .Y(_2643_)
);

FILL FILL_3__10918_ (
);

FILL FILL_1__11952_ (
);

FILL FILL_1__11532_ (
);

FILL FILL_1__11112_ (
);

FILL FILL_2__8557_ (
);

FILL FILL_0__10945_ (
);

FILL FILL_2__8137_ (
);

FILL FILL_0__10525_ (
);

AOI22X1 _10810_ (
    .A(\X[5] [0]),
    .B(vdd),
    .C(vdd),
    .D(\X[5] [4]),
    .Y(_4012_)
);

FILL FILL_0__10105_ (
);

NOR2X1 _13282_ (
    .A(\u_fir_pe7.rYin [10]),
    .B(\u_fir_pe7.mul [10]),
    .Y(_6306_)
);

FILL FILL_1__6974_ (
);

FILL FILL_1__6554_ (
);

FILL FILL_2__13324_ (
);

FILL FILL_1__12737_ (
);

FILL FILL_1__12317_ (
);

FILL FILL_0__9744_ (
);

FILL FILL_0__9324_ (
);

FILL FILL_1__7759_ (
);

FILL FILL_1__7339_ (
);

FILL FILL_3__10251_ (
);

FILL FILL_1__8700_ (
);

FILL FILL_3__8206_ (
);

NAND2X1 _7770_ (
    .A(_1282_),
    .B(_1269_),
    .Y(_1286_)
);

INVX2 _7350_ (
    .A(\X[1]_5_bF$buf0 ),
    .Y(_871_)
);

FILL FILL_3__11876_ (
);

FILL FILL_2__6623_ (
);

FILL FILL_3__11036_ (
);

FILL FILL_1__12070_ (
);

FILL FILL_2__10869_ (
);

FILL FILL_2__10449_ (
);

FILL FILL_2__9095_ (
);

FILL FILL_0__11483_ (
);

FILL FILL_2__10029_ (
);

FILL FILL_0__11063_ (
);

FILL FILL_1__9905_ (
);

FILL FILL_2__11810_ (
);

FILL FILL_0__6869_ (
);

DFFPOSX1 _8975_ (
    .D(\X[2] [6]),
    .CLK(clk_bF$buf14),
    .Q(\X[3] [6])
);

FILL FILL_0__6449_ (
);

NOR2X1 _8555_ (
    .A(_1726_),
    .B(_1915_),
    .Y(_1992_)
);

NOR2X1 _8135_ (
    .A(_2283_),
    .B(_2304_),
    .Y(_2314_)
);

FILL FILL_1__7092_ (
);

FILL FILL_1__10803_ (
);

FILL FILL_2__7828_ (
);

FILL FILL_0__7810_ (
);

FILL FILL_2__7408_ (
);

FILL FILL_1__13275_ (
);

NAND3X1 _12973_ (
    .A(_6005_),
    .B(_6009_),
    .C(_5964_),
    .Y(_6010_)
);

FILL FILL_0__12688_ (
);

FILL FILL_0__12268_ (
);

OAI21X1 _12553_ (
    .A(_6357_),
    .B(_5594_),
    .C(_5595_),
    .Y(_5596_)
);

NOR2X1 _12133_ (
    .A(_4797_),
    .B(_5244_),
    .Y(_5249_)
);

FILL FILL_1__8297_ (
);

FILL FILL_3__9584_ (
);

DFFPOSX1 _13338_ (
    .D(_6368_[0]),
    .CLK(clk_bF$buf9),
    .Q(\Y[7] [0])
);

FILL FILL_2__7581_ (
);

FILL FILL_2__7161_ (
);

NOR2X1 _6621_ (
    .A(_213_),
    .B(_215_),
    .Y(_220_)
);

OAI21X1 _9093_ (
    .A(_2454_),
    .B(_2453_),
    .C(_2420_),
    .Y(_2455_)
);

FILL FILL_1__11761_ (
);

FILL FILL_3__10307_ (
);

FILL FILL_1__11341_ (
);

FILL FILL_2__8786_ (
);

FILL FILL_2__8366_ (
);

FILL FILL_0__10334_ (
);

NAND2X1 _13091_ (
    .A(_6121_),
    .B(_6125_),
    .Y(_6126_)
);

NAND2X1 _7826_ (
    .A(_1337_),
    .B(_1313_),
    .Y(_1341_)
);

OAI21X1 _7406_ (
    .A(_925_),
    .B(_926_),
    .C(_924_),
    .Y(_927_)
);

FILL FILL_1__6783_ (
);

FILL FILL_2__13133_ (
);

FILL FILL_1__12966_ (
);

FILL FILL_1__12546_ (
);

FILL FILL_1__12126_ (
);

FILL FILL_0__9973_ (
);

FILL FILL_0__9553_ (
);

FILL FILL_0__11959_ (
);

FILL FILL_3__7650_ (
);

FILL FILL_0__9133_ (
);

NAND3X1 _11824_ (
    .A(_4939_),
    .B(_4943_),
    .C(_4941_),
    .Y(_4944_)
);

FILL FILL_0__11539_ (
);

AND2X2 _11404_ (
    .A(_4593_),
    .B(_4590_),
    .Y(_4597_)
);

FILL FILL_0__11119_ (
);

FILL FILL_0__12900_ (
);

FILL FILL_1__7988_ (
);

FILL FILL_1__7568_ (
);

FILL FILL_3__10480_ (
);

FILL FILL_1__7148_ (
);

FILL FILL_3__8435_ (
);

INVX1 _12609_ (
    .A(_5649_),
    .Y(_5650_)
);

FILL FILL_2__6852_ (
);

FILL FILL_2__6432_ (
);

FILL FILL_3__11265_ (
);

FILL FILL_2__10678_ (
);

FILL FILL_2__10258_ (
);

FILL FILL_0__11292_ (
);

FILL FILL_1__9714_ (
);

FILL FILL_0__6678_ (
);

OAI21X1 _8784_ (
    .A(_2210_),
    .B(_2209_),
    .C(_2215_),
    .Y(_2216_)
);

OAI21X1 _8364_ (
    .A(_1730_),
    .B(_1802_),
    .C(_1771_),
    .Y(_1803_)
);

FILL FILL_1__10612_ (
);

FILL FILL_2__7637_ (
);

FILL FILL_1__13084_ (
);

AND2X2 _12782_ (
    .A(vdd),
    .B(\X[6]_5_bF$buf1 ),
    .Y(_5821_)
);

FILL FILL_0__12077_ (
);

NOR2X1 _12362_ (
    .A(_5463_),
    .B(_5464_),
    .Y(_5465_)
);

FILL FILL_3__13411_ (
);

FILL FILL_2__12824_ (
);

FILL FILL_2__12404_ (
);

AND2X2 _9989_ (
    .A(_3265_),
    .B(_3269_),
    .Y(_3270_)
);

AND2X2 _9569_ (
    .A(_2914_),
    .B(_2910_),
    .Y(_2924_)
);

NAND3X1 _9149_ (
    .A(_2445_),
    .B(_2508_),
    .C(_2509_),
    .Y(_2510_)
);

FILL FILL_1__11817_ (
);

FILL FILL_0__8824_ (
);

FILL FILL_3__6921_ (
);

FILL FILL_0__8404_ (
);

NAND2X1 _13147_ (
    .A(_6178_),
    .B(_6179_),
    .Y(_6180_)
);

FILL FILL_1__6839_ (
);

FILL FILL_1__6419_ (
);

FILL FILL_2__7390_ (
);

FILL FILL_0__9609_ (
);

FILL FILL_3__7706_ (
);

AOI21X1 _6850_ (
    .A(_446_),
    .B(_445_),
    .C(_438_),
    .Y(_447_)
);

OAI22X1 _6430_ (
    .A(_30_),
    .B(_31_),
    .C(_0_),
    .D(_4_),
    .Y(_32_)
);

FILL FILL_1__11990_ (
);

FILL FILL_1__11570_ (
);

FILL FILL_1__11150_ (
);

FILL FILL_2__8595_ (
);

FILL FILL_0__10983_ (
);

FILL FILL_2__8175_ (
);

FILL FILL_0__10563_ (
);

FILL FILL_0__10143_ (
);

AOI21X1 _7635_ (
    .A(_1152_),
    .B(_1151_),
    .C(_1150_),
    .Y(_1153_)
);

DFFPOSX1 _7215_ (
    .D(Xin[0]),
    .CLK(clk_bF$buf33),
    .Q(\X[1] [0])
);

FILL FILL_1__6592_ (
);

FILL FILL_2__6908_ (
);

FILL FILL_1__12775_ (
);

FILL FILL_1__12355_ (
);

FILL FILL_0__9782_ (
);

FILL FILL_0__9362_ (
);

FILL FILL_0__11768_ (
);

DFFPOSX1 _11633_ (
    .D(_4781_[9]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [9])
);

FILL FILL_0__11348_ (
);

NAND3X1 _11213_ (
    .A(_4328_),
    .B(_4334_),
    .C(_4409_),
    .Y(_4410_)
);

FILL FILL_1__7797_ (
);

FILL FILL_1__7377_ (
);

FILL FILL_3__8664_ (
);

NAND2X1 _12838_ (
    .A(_5875_),
    .B(_5874_),
    .Y(_5876_)
);

NAND2X1 _12418_ (
    .A(_5517_),
    .B(_5510_),
    .Y(_5521_)
);

FILL FILL_2__6661_ (
);

FILL FILL_3__11494_ (
);

FILL FILL_2__10487_ (
);

FILL FILL_2__10067_ (
);

FILL FILL_1__9943_ (
);

FILL FILL_1__9523_ (
);

FILL FILL_1__9103_ (
);

FILL FILL_3__9449_ (
);

FILL FILL_0__6487_ (
);

OAI21X1 _8593_ (
    .A(_2029_),
    .B(_2028_),
    .C(_2027_),
    .Y(_2030_)
);

INVX1 _8173_ (
    .A(_1615_),
    .Y(_1616_)
);

FILL FILL_1__10841_ (
);

FILL FILL_1__10421_ (
);

FILL FILL_1__10001_ (
);

FILL FILL_2__7866_ (
);

FILL FILL_2__7446_ (
);

FILL FILL_3__12279_ (
);

FILL FILL_2__7026_ (
);

INVX1 _12591_ (
    .A(_5632_),
    .Y(_5633_)
);

NOR2X1 _12171_ (
    .A(_5284_),
    .B(_5286_),
    .Y(_5287_)
);

FILL FILL_3__13220_ (
);

AOI21X1 _6906_ (
    .A(_495_),
    .B(_501_),
    .C(_459_),
    .Y(_502_)
);

FILL FILL_2__12633_ (
);

FILL FILL_2__12213_ (
);

INVX1 _9798_ (
    .A(\u_fir_pe3.rYin [13]),
    .Y(_3142_)
);

AOI21X1 _9378_ (
    .A(_2735_),
    .B(_2734_),
    .C(_2733_),
    .Y(_2736_)
);

FILL FILL_1__11206_ (
);

FILL FILL_0__8633_ (
);

FILL FILL_0__8213_ (
);

FILL FILL_0__10619_ (
);

NAND3X1 _10904_ (
    .A(_4101_),
    .B(_4104_),
    .C(_4053_),
    .Y(_4105_)
);

FILL FILL254550x219750 (
);

DFFPOSX1 _13376_ (
    .D(\Y[6] [14]),
    .CLK(clk_bF$buf40),
    .Q(\u_fir_pe7.rYin [14])
);

FILL FILL_1__6648_ (
);

FILL FILL_3__7935_ (
);

FILL FILL_0__9418_ (
);

FILL FILL_3__10765_ (
);

FILL FILL_3__10345_ (
);

FILL FILL_0__10792_ (
);

FILL FILL_0__10372_ (
);

INVX1 _7864_ (
    .A(_1377_),
    .Y(_1378_)
);

NAND3X1 _7444_ (
    .A(_952_),
    .B(_963_),
    .C(_959_),
    .Y(_964_)
);

OAI21X1 _7024_ (
    .A(_584_),
    .B(_609_),
    .C(_608_),
    .Y(_616_)
);

FILL FILL_2__13171_ (
);

FILL FILL_2__6717_ (
);

FILL FILL_1__12584_ (
);

FILL FILL_1__12164_ (
);

FILL FILL_0__11997_ (
);

FILL FILL_0__9591_ (
);

FILL FILL_2__9189_ (
);

FILL FILL_0__9171_ (
);

AOI21X1 _11862_ (
    .A(_4964_),
    .B(_4959_),
    .C(_4966_),
    .Y(_4982_)
);

FILL FILL_0__11577_ (
);

NOR2X1 _11442_ (
    .A(_4627_),
    .B(_4626_),
    .Y(_4630_)
);

FILL FILL_0__11157_ (
);

OAI21X1 _11022_ (
    .A(_4763_),
    .B(_4220_),
    .C(_4212_),
    .Y(_4221_)
);

FILL FILL_2__11904_ (
);

NAND3X1 _8649_ (
    .A(_2082_),
    .B(_2084_),
    .C(_2083_),
    .Y(_2085_)
);

OAI21X1 _8229_ (
    .A(_2372_),
    .B(_1668_),
    .C(_1669_),
    .Y(_1670_)
);

FILL FILL_1__7186_ (
);

FILL FILL_0__7904_ (
);

FILL FILL_3__8893_ (
);

AOI21X1 _12647_ (
    .A(_5679_),
    .B(_5675_),
    .C(_5661_),
    .Y(_5688_)
);

FILL FILL_3__8053_ (
);

AOI21X1 _12227_ (
    .A(_5338_),
    .B(_5239_),
    .C(_5340_),
    .Y(_5341_)
);

FILL FILL_0__13303_ (
);

FILL FILL_2__6890_ (
);

FILL FILL_2__6470_ (
);

FILL FILL_2__10296_ (
);

FILL FILL_1__9752_ (
);

FILL FILL_1__9332_ (
);

FILL FILL_3__9678_ (
);

FILL FILL_1__10650_ (
);

FILL FILL_1__10230_ (
);

FILL FILL_2__7675_ (
);

FILL FILL_2__7255_ (
);

NAND2X1 _6715_ (
    .A(_306_),
    .B(_307_),
    .Y(_313_)
);

FILL FILL_2__12862_ (
);

FILL FILL_2__12442_ (
);

FILL FILL_2__12022_ (
);

NAND2X1 _9187_ (
    .A(vdd),
    .B(\X[3]_5_bF$buf2 ),
    .Y(_2547_)
);

FILL FILL_1__11855_ (
);

FILL FILL_1__11435_ (
);

FILL FILL_1__11015_ (
);

FILL FILL_0__8862_ (
);

FILL FILL_0__8442_ (
);

FILL FILL_0__10848_ (
);

FILL FILL_0__10428_ (
);

DFFPOSX1 _10713_ (
    .D(_3978_[6]),
    .CLK(clk_bF$buf21),
    .Q(\Y[5] [6])
);

FILL FILL_0__8022_ (
);

FILL FILL_0__10008_ (
);

NOR2X1 _13185_ (
    .A(\u_fir_pe7.rYin [1]),
    .B(\u_fir_pe7.mul [1]),
    .Y(_6214_)
);

FILL FILL_2__9821_ (
);

FILL FILL_2__9401_ (
);

FILL FILL_1__6877_ (
);

FILL FILL_1__6457_ (
);

FILL FILL_2__13227_ (
);

FILL FILL_0__9647_ (
);

FILL FILL_0__9227_ (
);

NOR2X1 _11918_ (
    .A(_5023_),
    .B(_5036_),
    .Y(_5037_)
);

FILL FILL_3__7324_ (
);

FILL FILL_3__10994_ (
);

FILL FILL_3__10574_ (
);

FILL FILL_0__10181_ (
);

FILL FILL_1__8603_ (
);

FILL FILL_3__8529_ (
);

INVX1 _7673_ (
    .A(_1187_),
    .Y(_1190_)
);

DFFPOSX1 _7253_ (
    .D(_796_[14]),
    .CLK(clk_bF$buf1),
    .Q(\u_fir_pe0.mul [14])
);

FILL FILL_2__6946_ (
);

FILL FILL_3__11779_ (
);

FILL FILL_2__6526_ (
);

FILL FILL_3__11359_ (
);

FILL FILL_1__12393_ (
);

OAI21X1 _11671_ (
    .A(_4786_),
    .B(_4789_),
    .C(_4783_),
    .Y(_4794_)
);

FILL FILL_0__11386_ (
);

INVX2 _11251_ (
    .A(gnd),
    .Y(_4447_)
);

FILL FILL_1__9808_ (
);

FILL FILL_3__12720_ (
);

FILL FILL_2__11713_ (
);

NAND2X1 _8878_ (
    .A(_2298_),
    .B(_2301_),
    .Y(_2384_[8])
);

AOI21X1 _8458_ (
    .A(_1860_),
    .B(_1861_),
    .C(_1818_),
    .Y(_1896_)
);

NOR2X1 _8038_ (
    .A(\u_fir_pe1.rYin [12]),
    .B(\u_fir_pe1.mul [12]),
    .Y(_1542_)
);

FILL FILL_1__10706_ (
);

FILL FILL_0__7713_ (
);

FILL FILL_1__13178_ (
);

AOI21X1 _12876_ (
    .A(_5911_),
    .B(_5913_),
    .C(_5909_),
    .Y(_5914_)
);

FILL FILL_3__8282_ (
);

NOR2X1 _12456_ (
    .A(_5558_),
    .B(_5413_),
    .Y(_5571_[0])
);

NAND3X1 _12036_ (
    .A(_5151_),
    .B(_5152_),
    .C(_5153_),
    .Y(_5154_)
);

FILL FILL_2__12918_ (
);

FILL FILL_0__13112_ (
);

FILL FILL_0__8918_ (
);

FILL FILL_1__9981_ (
);

FILL FILL_1__9561_ (
);

FILL FILL_1__9141_ (
);

FILL FILL_3__9067_ (
);

FILL FILL_2__7484_ (
);

FILL FILL_2__7064_ (
);

AOI21X1 _6944_ (
    .A(_470_),
    .B(_486_),
    .C(_538_),
    .Y(_539_)
);

NAND3X1 _6524_ (
    .A(_123_),
    .B(_124_),
    .C(_122_),
    .Y(_125_)
);

FILL FILL_2__12671_ (
);

FILL FILL_2__12251_ (
);

FILL FILL_1__11664_ (
);

FILL FILL_1__11244_ (
);

FILL FILL_2__8689_ (
);

FILL FILL_0__8671_ (
);

FILL FILL_0__8251_ (
);

FILL FILL_2__8269_ (
);

FILL FILL_0__10657_ (
);

INVX1 _10942_ (
    .A(_4141_),
    .Y(_4142_)
);

AND2X2 _10522_ (
    .A(_3791_),
    .B(_3790_),
    .Y(_3795_)
);

FILL FILL_0__10237_ (
);

OAI21X1 _10102_ (
    .A(_3381_),
    .B(_3376_),
    .C(_3304_),
    .Y(_3382_)
);

FILL FILL_2__9630_ (
);

FILL FILL_2__9210_ (
);

OAI21X1 _7729_ (
    .A(_1244_),
    .B(_1245_),
    .C(_1241_),
    .Y(_1246_)
);

INVX1 _7309_ (
    .A(_830_),
    .Y(_831_)
);

FILL FILL_1__6686_ (
);

FILL FILL_2__13036_ (
);

FILL FILL_1__12869_ (
);

FILL FILL_1__12449_ (
);

FILL FILL_1__12029_ (
);

FILL FILL_3__7973_ (
);

FILL FILL_0__9456_ (
);

FILL FILL_3__7553_ (
);

FILL FILL_0__9036_ (
);

NAND2X1 _11727_ (
    .A(_4848_),
    .B(_4842_),
    .Y(_5577_[4])
);

FILL FILL_3__7133_ (
);

NOR3X1 _11307_ (
    .A(_4290_),
    .B(_4458_),
    .C(_4401_),
    .Y(_4502_)
);

FILL FILL_0__12803_ (
);

FILL FILL254250x205350 (
);

FILL FILL_1__8832_ (
);

FILL FILL_1__8412_ (
);

FILL FILL_3__8758_ (
);

OAI21X1 _7482_ (
    .A(_926_),
    .B(_924_),
    .C(_917_),
    .Y(_1002_)
);

INVX1 _7062_ (
    .A(\u_fir_pe0.mul [3]),
    .Y(_649_)
);

FILL FILL_2__6755_ (
);

OR2X2 _11480_ (
    .A(_4657_),
    .B(_4662_),
    .Y(_4664_)
);

FILL FILL_0__11195_ (
);

OAI21X1 _11060_ (
    .A(_4258_),
    .B(_4254_),
    .C(_4194_),
    .Y(_4259_)
);

FILL FILL_1__9617_ (
);

FILL FILL_2__11942_ (
);

FILL FILL_2__11522_ (
);

FILL FILL_2__11102_ (
);

OAI21X1 _8687_ (
    .A(_2067_),
    .B(_2120_),
    .C(_2121_),
    .Y(_2122_)
);

NAND3X1 _8267_ (
    .A(_1695_),
    .B(_1699_),
    .C(_1701_),
    .Y(_1708_)
);

FILL FILL_1__10935_ (
);

FILL FILL_1__10515_ (
);

FILL FILL254550x61350 (
);

FILL FILL_0__7942_ (
);

FILL FILL_0__7522_ (
);

FILL FILL_0__7102_ (
);

OAI21X1 _12685_ (
    .A(_6357_),
    .B(_5723_),
    .C(_5724_),
    .Y(_5725_)
);

NAND2X1 _12265_ (
    .A(_5349_),
    .B(_5377_),
    .Y(_5378_)
);

FILL FILL_2__8901_ (
);

FILL FILL_3__13314_ (
);

FILL FILL_2__12727_ (
);

FILL FILL_2__12307_ (
);

FILL FILL_0__8727_ (
);

FILL FILL_0__8307_ (
);

FILL FILL_3__6404_ (
);

FILL FILL_1__9790_ (
);

FILL FILL_1__9370_ (
);

FILL FILL_3__9296_ (
);

FILL FILL_2__7293_ (
);

NAND3X1 _6753_ (
    .A(_349_),
    .B(_350_),
    .C(_348_),
    .Y(_351_)
);

FILL FILL_2__12060_ (
);

FILL FILL_3__10859_ (
);

FILL FILL_1__11893_ (
);

FILL FILL_3__10439_ (
);

FILL FILL_1__11473_ (
);

FILL FILL_3__10019_ (
);

FILL FILL_1__11053_ (
);

FILL FILL_0__8480_ (
);

FILL FILL_2__8498_ (
);

FILL FILL_0__10886_ (
);

FILL FILL_0__10466_ (
);

FILL FILL_0__8060_ (
);

DFFPOSX1 _10751_ (
    .D(_3983_[4]),
    .CLK(clk_bF$buf54),
    .Q(\u_fir_pe4.mul [4])
);

NAND2X1 _10331_ (
    .A(_3591_),
    .B(_3601_),
    .Y(_3608_)
);

FILL FILL_0__10046_ (
);

INVX1 _7958_ (
    .A(\u_fir_pe1.mul [5]),
    .Y(_1463_)
);

NAND3X1 _7538_ (
    .A(_1036_),
    .B(_1050_),
    .C(_1053_),
    .Y(_1057_)
);

NAND3X1 _7118_ (
    .A(_701_),
    .B(_698_),
    .C(_661_),
    .Y(_702_)
);

FILL FILL_1__6495_ (
);

FILL FILL_2__13265_ (
);

FILL FILL_1__12678_ (
);

FILL FILL_1__12258_ (
);

FILL FILL_0__9685_ (
);

FILL FILL_0__9265_ (
);

INVX1 _11956_ (
    .A(_5070_),
    .Y(_5075_)
);

NOR2X1 _11536_ (
    .A(_4719_),
    .B(_4718_),
    .Y(_4720_)
);

AOI21X1 _11116_ (
    .A(_4313_),
    .B(_4311_),
    .C(_4309_),
    .Y(_4314_)
);

FILL FILL253350x43350 (
);

FILL FILL_0__12612_ (
);

FILL FILL_3__10192_ (
);

FILL FILL_1__8641_ (
);

FILL FILL_1__8221_ (
);

FILL FILL_3__8147_ (
);

OAI21X1 _7291_ (
    .A(_1575_),
    .B(_812_),
    .C(_813_),
    .Y(_814_)
);

FILL FILL_2__6984_ (
);

FILL FILL_2__6564_ (
);

FILL FILL_1__9426_ (
);

FILL FILL_2__11751_ (
);

FILL FILL_2__11331_ (
);

NAND3X1 _8496_ (
    .A(_1932_),
    .B(_1933_),
    .C(_1931_),
    .Y(_1934_)
);

DFFPOSX1 _8076_ (
    .D(_1586_[0]),
    .CLK(clk_bF$buf57),
    .Q(\Y[2] [0])
);

FILL FILL_1__10324_ (
);

FILL FILL_0__7751_ (
);

FILL FILL_2__7769_ (
);

FILL FILL_2__7349_ (
);

FILL FILL_0__7331_ (
);

DFFPOSX1 _12494_ (
    .D(\Y[7] [9]),
    .CLK(clk_bF$buf46),
    .Q(\u_fir_pe6.rYin [9])
);

AOI22X1 _12074_ (
    .A(_5024_),
    .B(_5190_),
    .C(_5116_),
    .D(_5112_),
    .Y(_5191_)
);

FILL FILL_2__8710_ (
);

FILL FILL_3__13123_ (
);

AOI21X1 _6809_ (
    .A(_331_),
    .B(_405_),
    .C(_404_),
    .Y(_406_)
);

FILL FILL_2__12956_ (
);

FILL FILL_2__12536_ (
);

FILL FILL_2__12116_ (
);

FILL FILL_0__13150_ (
);

FILL FILL_1__11949_ (
);

FILL FILL_1__11529_ (
);

FILL FILL_1__11109_ (
);

FILL FILL_0__8536_ (
);

FILL FILL_3__6633_ (
);

NAND2X1 _10807_ (
    .A(\X[5] [0]),
    .B(vdd),
    .Y(_4009_)
);

INVX1 _13279_ (
    .A(\u_fir_pe7.rYin [10]),
    .Y(_6303_)
);

FILL FILL_2__9915_ (
);

FILL FILL_1__7912_ (
);

FILL FILL_3__7418_ (
);

NAND2X1 _6982_ (
    .A(_572_),
    .B(_575_),
    .Y(_576_)
);

NAND3X1 _6562_ (
    .A(_157_),
    .B(_161_),
    .C(_159_),
    .Y(_162_)
);

FILL FILL_3__10668_ (
);

FILL FILL_3__10248_ (
);

FILL FILL_1__11282_ (
);

FILL FILL_0__10695_ (
);

AOI21X1 _10980_ (
    .A(_4103_),
    .B(_4102_),
    .C(_4039_),
    .Y(_4180_)
);

OAI21X1 _10560_ (
    .A(_3820_),
    .B(_3821_),
    .C(_3825_),
    .Y(_3828_)
);

FILL FILL_0__10275_ (
);

INVX1 _10140_ (
    .A(_3418_),
    .Y(_3419_)
);

FILL FILL_2__10602_ (
);

NAND3X1 _7767_ (
    .A(_1204_),
    .B(_1282_),
    .C(_1212_),
    .Y(_1283_)
);

INVX1 _7347_ (
    .A(_867_),
    .Y(_868_)
);

FILL FILL_2__13074_ (
);

FILL FILL_0__6602_ (
);

FILL FILL_1__12067_ (
);

FILL FILL_0__9494_ (
);

FILL FILL_3__7591_ (
);

FILL FILL_0__9074_ (
);

NAND3X1 _11765_ (
    .A(_4877_),
    .B(_4873_),
    .C(_4879_),
    .Y(_4886_)
);

OAI21X1 _11345_ (
    .A(_4489_),
    .B(_4492_),
    .C(_4537_),
    .Y(_4540_)
);

FILL FILL_3__12814_ (
);

FILL FILL_2__11807_ (
);

FILL FILL_0__12841_ (
);

FILL FILL_0__12421_ (
);

FILL FILL_0__12001_ (
);

FILL FILL_1__7089_ (
);

FILL FILL_0__7807_ (
);

OAI21X1 _9913_ (
    .A(_3192_),
    .B(_3195_),
    .C(_3188_),
    .Y(_3196_)
);

FILL FILL_1__8870_ (
);

FILL FILL_1__8450_ (
);

FILL FILL_1__8030_ (
);

FILL FILL_3__8376_ (
);

FILL FILL_0__13206_ (
);

FILL FILL_2__6793_ (
);

FILL FILL_2__10199_ (
);

FILL FILL_1__9655_ (
);

FILL FILL_1__9235_ (
);

FILL FILL_2__11980_ (
);

FILL FILL_2__11560_ (
);

FILL FILL_2__11140_ (
);

FILL FILL_1__10973_ (
);

FILL FILL_1__10553_ (
);

FILL FILL_1__10133_ (
);

FILL FILL_0__7980_ (
);

FILL FILL_2__7998_ (
);

FILL FILL_2__7578_ (
);

FILL FILL_0__7560_ (
);

FILL FILL_0__7140_ (
);

FILL FILL_2__7158_ (
);

NAND3X1 _6618_ (
    .A(_143_),
    .B(_212_),
    .C(_147_),
    .Y(_217_)
);

FILL FILL_2__12765_ (
);

FILL FILL_2__12345_ (
);

FILL FILL_1__11758_ (
);

FILL FILL_1__11338_ (
);

FILL FILL_0__8765_ (
);

FILL FILL_3__6862_ (
);

FILL FILL_0__8345_ (
);

INVX1 _10616_ (
    .A(\u_fir_pe4.mul [8]),
    .Y(_3879_)
);

NAND2X1 _13088_ (
    .A(_6119_),
    .B(_6095_),
    .Y(_6123_)
);

FILL FILL_2__9724_ (
);

FILL FILL_2__9304_ (
);

FILL FILL_1__7721_ (
);

FILL FILL_1__7301_ (
);

FILL FILL_3__7647_ (
);

NAND2X1 _6791_ (
    .A(gnd),
    .B(_387_),
    .Y(_388_)
);

FILL FILL_1__11091_ (
);

FILL FILL_0__10084_ (
);

FILL FILL_1__8926_ (
);

FILL FILL_1__8506_ (
);

FILL FILL_2__10831_ (
);

FILL FILL_2__10411_ (
);

NAND2X1 _7996_ (
    .A(_1496_),
    .B(_1499_),
    .Y(_1500_)
);

NAND2X1 _7576_ (
    .A(_1093_),
    .B(_1092_),
    .Y(_1094_)
);

NAND2X1 _7156_ (
    .A(_735_),
    .B(_728_),
    .Y(_739_)
);

FILL FILL_2__6849_ (
);

FILL FILL_0__6831_ (
);

FILL FILL_0__6411_ (
);

FILL FILL_2__6429_ (
);

FILL FILL_1__12296_ (
);

INVX1 _11994_ (
    .A(_5106_),
    .Y(_5112_)
);

INVX1 _11574_ (
    .A(_4757_),
    .Y(_4758_)
);

FILL FILL_0__11289_ (
);

OAI21X1 _11154_ (
    .A(_4351_),
    .B(_4348_),
    .C(_4284_),
    .Y(_4352_)
);

FILL FILL_3__12203_ (
);

FILL FILL_0__12650_ (
);

FILL FILL_0__12230_ (
);

FILL FILL_1__10609_ (
);

FILL FILL_0__7616_ (
);

NOR2X1 _9722_ (
    .A(_3064_),
    .B(_3065_),
    .Y(_3066_)
);

AND2X2 _9302_ (
    .A(_2612_),
    .B(_2609_),
    .Y(_2661_)
);

OAI21X1 _12779_ (
    .A(_5735_),
    .B(_5739_),
    .C(_5738_),
    .Y(_5818_)
);

OAI21X1 _12359_ (
    .A(_5455_),
    .B(_5456_),
    .C(_5460_),
    .Y(_5462_)
);

FILL FILL_0__13015_ (
);

NOR2X1 _13300_ (
    .A(\u_fir_pe7.rYin [12]),
    .B(\u_fir_pe7.mul [12]),
    .Y(_6324_)
);

FILL FILL_1__9464_ (
);

FILL FILL_1__9044_ (
);

FILL FILL_1__10782_ (
);

FILL FILL_1__10362_ (
);

FILL FILL_2__7387_ (
);

FILL FILL_3__13161_ (
);

AOI21X1 _6847_ (
    .A(_300_),
    .B(_365_),
    .C(_443_),
    .Y(_444_)
);

INVX1 _6427_ (
    .A(_28_),
    .Y(_29_)
);

FILL FILL_2__12994_ (
);

FILL FILL_2__12574_ (
);

FILL FILL_2__12154_ (
);

FILL FILL_1__11987_ (
);

FILL FILL_1__11567_ (
);

FILL FILL_1__11147_ (
);

FILL FILL_0__8574_ (
);

FILL FILL_0__8154_ (
);

INVX1 _10845_ (
    .A(_4030_),
    .Y(_4047_)
);

NAND2X1 _10425_ (
    .A(_3693_),
    .B(_3697_),
    .Y(_3700_)
);

AOI21X1 _10005_ (
    .A(_3280_),
    .B(_3282_),
    .C(_3273_),
    .Y(_3286_)
);

FILL FILL_2__9953_ (
);

FILL FILL_2__9533_ (
);

FILL FILL_0__11921_ (
);

FILL FILL_2__9113_ (
);

FILL FILL_0__11501_ (
);

FILL FILL_1__6589_ (
);

FILL FILL_1__7950_ (
);

FILL FILL_1__7530_ (
);

FILL FILL_1__7110_ (
);

FILL FILL_0__9779_ (
);

FILL FILL_3__7876_ (
);

FILL FILL_0__9359_ (
);

FILL FILL_0__12706_ (
);

FILL FILL_3__10286_ (
);

FILL FILL_1__8735_ (
);

FILL FILL_1__8315_ (
);

FILL FILL_2__10640_ (
);

FILL FILL_2__10220_ (
);

AOI21X1 _7385_ (
    .A(_897_),
    .B(_893_),
    .C(_879_),
    .Y(_906_)
);

FILL FILL_3__9602_ (
);

FILL FILL_0__6640_ (
);

FILL FILL_2__6658_ (
);

FILL FILL_0__11098_ (
);

NOR2X1 _11383_ (
    .A(_4545_),
    .B(_4568_),
    .Y(_4576_)
);

FILL FILL_3__12432_ (
);

FILL FILL_2__11845_ (
);

FILL FILL_2__11425_ (
);

FILL FILL_2__11005_ (
);

FILL FILL_1__10838_ (
);

FILL FILL_1__10418_ (
);

FILL FILL_0__7845_ (
);

NAND3X1 _9951_ (
    .A(_3220_),
    .B(_3232_),
    .C(_3228_),
    .Y(_3233_)
);

FILL FILL_0__7425_ (
);

INVX1 _9531_ (
    .A(_2851_),
    .Y(_2887_)
);

FILL FILL_0__7005_ (
);

NAND3X1 _9111_ (
    .A(_2461_),
    .B(_2469_),
    .C(_2471_),
    .Y(_2472_)
);

NAND3X1 _12588_ (
    .A(_5619_),
    .B(_5623_),
    .C(_5625_),
    .Y(_5630_)
);

AOI21X1 _12168_ (
    .A(_5277_),
    .B(_5283_),
    .C(_5241_),
    .Y(_5284_)
);

FILL FILL_2__8804_ (
);

FILL FILL_3__13217_ (
);

FILL FILL_0__13244_ (
);

FILL FILL_1__6801_ (
);

FILL FILL_3__6727_ (
);

FILL FILL_1__9693_ (
);

FILL FILL_1__9273_ (
);

FILL FILL_1__10591_ (
);

FILL FILL_1__10171_ (
);

FILL FILL_2__7196_ (
);

NOR2X1 _6656_ (
    .A(_241_),
    .B(_254_),
    .Y(_255_)
);

FILL FILL_2__12383_ (
);

FILL FILL_1__11796_ (
);

FILL FILL_1__11376_ (
);

FILL FILL_0__8383_ (
);

FILL FILL_0__10789_ (
);

FILL FILL_3__6480_ (
);

OAI21X1 _10654_ (
    .A(_3914_),
    .B(_3915_),
    .C(_3910_),
    .Y(_3918_)
);

FILL FILL_0__10369_ (
);

NAND2X1 _10234_ (
    .A(vdd),
    .B(\X[4] [7]),
    .Y(_3512_)
);

FILL FILL_3__11703_ (
);

FILL FILL_2__9762_ (
);

FILL FILL_2__9342_ (
);

FILL FILL_0__11730_ (
);

FILL FILL_0__11310_ (
);

FILL FILL_1__6398_ (
);

FILL FILL_2__13168_ (
);

NAND2X1 _8802_ (
    .A(_2225_),
    .B(_2230_),
    .Y(_2231_)
);

FILL FILL_0__9588_ (
);

FILL FILL_3__7685_ (
);

FILL FILL_0__9168_ (
);

INVX1 _11859_ (
    .A(_4888_),
    .Y(_4979_)
);

FILL FILL_3__7265_ (
);

NOR2X1 _11439_ (
    .A(\u_fir_pe5.rYin [2]),
    .B(\u_fir_pe5.mul [2]),
    .Y(_4627_)
);

INVX1 _11019_ (
    .A(vdd),
    .Y(_4218_)
);

FILL FILL_3__12908_ (
);

FILL FILL_1__13102_ (
);

FILL FILL_0__12935_ (
);

NAND3X1 _12800_ (
    .A(_5818_),
    .B(_5832_),
    .C(_5835_),
    .Y(_5839_)
);

FILL FILL_1__8544_ (
);

NOR2X1 _7194_ (
    .A(_776_),
    .B(_631_),
    .Y(_789_[0])
);

FILL FILL_2__6887_ (
);

FILL FILL_2__6467_ (
);

AOI22X1 _11192_ (
    .A(vdd),
    .B(\X[5] [6]),
    .C(gnd),
    .D(\X[5] [7]),
    .Y(_4389_)
);

FILL FILL_1__9749_ (
);

FILL FILL_1__9329_ (
);

FILL FILL_3__12661_ (
);

FILL FILL_2__11654_ (
);

FILL FILL_2__11234_ (
);

OAI21X1 _8399_ (
    .A(_1683_),
    .B(_1668_),
    .C(_1752_),
    .Y(_1838_)
);

FILL FILL_1__10647_ (
);

FILL FILL_1__10227_ (
);

FILL FILL_0__7654_ (
);

NOR2X1 _9760_ (
    .A(\u_fir_pe3.rYin [9]),
    .B(\u_fir_pe3.mul [9]),
    .Y(_3104_)
);

OAI21X1 _9340_ (
    .A(_2616_),
    .B(_2621_),
    .C(_2620_),
    .Y(_2698_)
);

NOR2X1 _12397_ (
    .A(_5497_),
    .B(_5491_),
    .Y(_5500_)
);

FILL FILL_2__8613_ (
);

FILL FILL_2__12859_ (
);

FILL FILL_2__12439_ (
);

FILL FILL_2__12019_ (
);

FILL FILL_0__13053_ (
);

FILL FILL_1__6610_ (
);

FILL FILL_0__8859_ (
);

FILL FILL_3__6956_ (
);

FILL FILL_0__8439_ (
);

FILL FILL_0__8019_ (
);

FILL FILL_1__9082_ (
);

FILL FILL_2__9818_ (
);

FILL FILL_0__9800_ (
);

FILL FILL_1__7815_ (
);

AOI21X1 _6885_ (
    .A(vdd),
    .B(Xin[6]),
    .C(_412_),
    .Y(_481_)
);

NAND2X1 _6465_ (
    .A(_66_),
    .B(_60_),
    .Y(_795_[4])
);

FILL FILL_2__12192_ (
);

FILL FILL_1__11185_ (
);

FILL FILL_0__8192_ (
);

FILL FILL_0__10598_ (
);

AOI22X1 _10883_ (
    .A(gnd),
    .B(\X[5] [4]),
    .C(_4073_),
    .D(_4075_),
    .Y(_4084_)
);

OAI21X1 _10463_ (
    .A(_3684_),
    .B(_3737_),
    .C(_3680_),
    .Y(_3738_)
);

FILL FILL_0__10178_ (
);

NAND2X1 _10043_ (
    .A(_3319_),
    .B(_3321_),
    .Y(_3323_)
);

FILL FILL_3__11932_ (
);

FILL FILL_3__11512_ (
);

FILL FILL_2__10925_ (
);

FILL FILL_2__9991_ (
);

FILL FILL_2__9571_ (
);

FILL FILL_2__10505_ (
);

FILL FILL_2__9151_ (
);

FILL FILL_2__13397_ (
);

FILL FILL_0__6925_ (
);

FILL FILL_0__6505_ (
);

NAND2X1 _8611_ (
    .A(_2036_),
    .B(_2043_),
    .Y(_2047_)
);

FILL FILL_0__9397_ (
);

FILL FILL_3__7494_ (
);

NAND3X1 _11668_ (
    .A(_5522_),
    .B(_4790_),
    .C(_4788_),
    .Y(_4791_)
);

FILL FILL_3__7074_ (
);

OAI21X1 _11248_ (
    .A(_4423_),
    .B(_4425_),
    .C(_4416_),
    .Y(_4444_)
);

FILL FILL_3__12717_ (
);

FILL FILL_1__13331_ (
);

FILL FILL_0__12744_ (
);

FILL FILL_0__12324_ (
);

NAND2X1 _9816_ (
    .A(_3155_),
    .B(_3149_),
    .Y(_3159_)
);

FILL FILL_1__8773_ (
);

FILL FILL_1__8353_ (
);

FILL FILL_3__8699_ (
);

FILL FILL_3__9220_ (
);

FILL FILL_0__13109_ (
);

FILL FILL_2__6696_ (
);

FILL FILL_1__9978_ (
);

FILL FILL_3__12890_ (
);

FILL FILL_1__9558_ (
);

FILL FILL_1__9138_ (
);

FILL FILL_3__12050_ (
);

FILL FILL_2__11883_ (
);

FILL FILL_2__11463_ (
);

FILL FILL_2__11043_ (
);

FILL FILL_1__10876_ (
);

FILL FILL_1__10456_ (
);

FILL FILL_1__10036_ (
);

FILL FILL_0__7883_ (
);

FILL FILL_0__7463_ (
);

FILL FILL_0__7043_ (
);

FILL FILL_2__8842_ (
);

FILL FILL_2__8422_ (
);

FILL FILL_0__10810_ (
);

FILL FILL_3__13255_ (
);

FILL FILL_2__8002_ (
);

FILL FILL_2__12668_ (
);

FILL FILL_2__12248_ (
);

FILL FILL_0__13282_ (
);

FILL FILL_0__8668_ (
);

FILL FILL_0__8248_ (
);

AOI22X1 _10939_ (
    .A(vdd),
    .B(\X[5] [2]),
    .C(gnd),
    .D(\X[5] [3]),
    .Y(_4139_)
);

NAND2X1 _10519_ (
    .A(_3790_),
    .B(_3791_),
    .Y(_3792_)
);

FILL FILL_1__12602_ (
);

FILL FILL_2__9627_ (
);

FILL FILL_2__9207_ (
);

FILL FILL_1__7624_ (
);

INVX1 _6694_ (
    .A(_288_),
    .Y(_293_)
);

FILL FILL_3__8911_ (
);

INVX1 _10692_ (
    .A(_3950_),
    .Y(_3955_)
);

NAND3X1 _10272_ (
    .A(_3548_),
    .B(_3549_),
    .C(_3547_),
    .Y(_3550_)
);

FILL FILL_1__8829_ (
);

FILL FILL_1__8409_ (
);

FILL FILL_2__9380_ (
);

FILL FILL_2__10314_ (
);

NAND3X1 _7899_ (
    .A(_1379_),
    .B(_1381_),
    .C(_1409_),
    .Y(_1411_)
);

NAND3X1 _7479_ (
    .A(_992_),
    .B(_993_),
    .C(_998_),
    .Y(_999_)
);

NAND2X1 _7059_ (
    .A(_643_),
    .B(_646_),
    .Y(_790_[2])
);

FILL FILL_0__6734_ (
);

OR2X2 _8840_ (
    .A(_2258_),
    .B(_2263_),
    .Y(_2265_)
);

AOI21X1 _8420_ (
    .A(_1746_),
    .B(_1765_),
    .C(_1858_),
    .Y(_1859_)
);

FILL FILL_1__12199_ (
);

NAND2X1 _8000_ (
    .A(_1502_),
    .B(_1503_),
    .Y(_1504_)
);

OAI21X1 _11897_ (
    .A(_4797_),
    .B(_5015_),
    .C(_5010_),
    .Y(_5016_)
);

NOR2X1 _11477_ (
    .A(\u_fir_pe5.rYin [6]),
    .B(\u_fir_pe5.mul [6]),
    .Y(_4661_)
);

NAND3X1 _11057_ (
    .A(_4209_),
    .B(_4251_),
    .C(_4252_),
    .Y(_4256_)
);

FILL FILL_1__13140_ (
);

FILL FILL_2__11939_ (
);

FILL FILL_0__12973_ (
);

FILL FILL_2__11519_ (
);

FILL FILL_0__12553_ (
);

FILL FILL_0__12133_ (
);

FILL FILL254250x100950 (
);

FILL FILL_0__7939_ (
);

FILL FILL_0__7519_ (
);

OAI21X1 _9625_ (
    .A(_2767_),
    .B(_2978_),
    .C(_2950_),
    .Y(_2979_)
);

OAI21X1 _9205_ (
    .A(_2560_),
    .B(_2561_),
    .C(_2546_),
    .Y(_2565_)
);

FILL FILL_1__8582_ (
);

FILL FILL_1__8162_ (
);

NOR2X1 _13203_ (
    .A(\u_fir_pe7.rYin [3]),
    .B(\u_fir_pe7.mul [3]),
    .Y(_6230_)
);

FILL FILL_1__9787_ (
);

FILL FILL_1__9367_ (
);

FILL FILL_2__11692_ (
);

FILL FILL_2__11272_ (
);

FILL FILL_1__10685_ (
);

FILL FILL_1__10265_ (
);

FILL FILL_0__7692_ (
);

FILL FILL_0__7272_ (
);

FILL FILL_2__8651_ (
);

FILL FILL_2__8231_ (
);

FILL FILL_2__12897_ (
);

FILL FILL_2__12057_ (
);

FILL FILL_0__13091_ (
);

FILL FILL_0__8897_ (
);

FILL FILL_0__8477_ (
);

FILL FILL_3__6574_ (
);

DFFPOSX1 _10748_ (
    .D(_3980_[1]),
    .CLK(clk_bF$buf55),
    .Q(\u_fir_pe4.mul [1])
);

FILL FILL_0__8057_ (
);

INVX1 _10328_ (
    .A(\X[4] [4]),
    .Y(_3605_)
);

FILL FILL_1__12831_ (
);

FILL FILL_1__12411_ (
);

FILL FILL_2__9436_ (
);

FILL FILL_0__11824_ (
);

FILL FILL_2__9016_ (
);

FILL FILL_0__11404_ (
);

FILL FILL_1__7853_ (
);

FILL FILL_1__7433_ (
);

FILL FILL_1__7013_ (
);

FILL FILL_3__7359_ (
);

FILL FILL_0__12609_ (
);

FILL FILL_3__10189_ (
);

NAND2X1 _10081_ (
    .A(_3339_),
    .B(_3335_),
    .Y(_3361_)
);

FILL FILL_3__11970_ (
);

FILL FILL_1__8638_ (
);

FILL FILL_1__8218_ (
);

FILL FILL_3__11130_ (
);

FILL FILL_2__10963_ (
);

FILL FILL_2__10543_ (
);

FILL FILL_2__10123_ (
);

NAND3X1 _7288_ (
    .A(_1585_),
    .B(_810_),
    .C(_806_),
    .Y(_811_)
);

FILL FILL_0__6963_ (
);

FILL FILL_0__6543_ (
);

NAND2X1 _11286_ (
    .A(_4478_),
    .B(_4446_),
    .Y(_4482_)
);

FILL FILL_2__7922_ (
);

FILL FILL_3__12755_ (
);

FILL FILL_2__7502_ (
);

FILL FILL_2__11748_ (
);

FILL FILL_0__12782_ (
);

FILL FILL_2__11328_ (
);

FILL FILL_0__12362_ (
);

FILL FILL_0__7748_ (
);

DFFPOSX1 _9854_ (
    .D(\Y[3] [0]),
    .CLK(clk_bF$buf56),
    .Q(\u_fir_pe3.rYin [0])
);

FILL FILL_0__7328_ (
);

NOR2X1 _9434_ (
    .A(_2789_),
    .B(_2790_),
    .Y(_2791_)
);

NOR2X1 _9014_ (
    .A(_3080_),
    .B(_3122_),
    .Y(_3131_)
);

FILL FILL_1__8391_ (
);

FILL FILL_2__8707_ (
);

FILL FILL_0__13147_ (
);

NAND3X1 _13012_ (
    .A(_6046_),
    .B(_6043_),
    .C(_6047_),
    .Y(_6048_)
);

FILL FILL_1__6704_ (
);

FILL FILL_1__9596_ (
);

FILL FILL_1__9176_ (
);

FILL FILL_2__11081_ (
);

FILL FILL_1__10494_ (
);

FILL FILL_1__10074_ (
);

FILL FILL_2__7099_ (
);

FILL FILL_0__7081_ (
);

FILL FILL_1__7909_ (
);

FILL FILL_3__10401_ (
);

FILL FILL_2__8880_ (
);

FILL FILL_2__8460_ (
);

FILL FILL_2__8040_ (
);

NOR2X1 _6979_ (
    .A(_565_),
    .B(_569_),
    .Y(_573_)
);

NAND2X1 _6559_ (
    .A(_87_),
    .B(_158_),
    .Y(_159_)
);

FILL FILL_2__12286_ (
);

INVX1 _7920_ (
    .A(\u_fir_pe1.rYin [1]),
    .Y(_1429_)
);

FILL FILL_1__11699_ (
);

NAND2X1 _7500_ (
    .A(_1015_),
    .B(_1018_),
    .Y(_1019_)
);

FILL FILL_1__11279_ (
);

FILL FILL_0__8286_ (
);

NAND3X1 _10977_ (
    .A(_4121_),
    .B(_4170_),
    .C(_4171_),
    .Y(_4177_)
);

INVX1 _10557_ (
    .A(_3825_),
    .Y(_3826_)
);

AND2X2 _10137_ (
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3416_)
);

FILL FILL_1__12640_ (
);

FILL FILL_1__12220_ (
);

FILL FILL_2__9665_ (
);

FILL FILL_2__9245_ (
);

FILL FILL_0__11213_ (
);

NAND3X1 _8705_ (
    .A(_2137_),
    .B(_2139_),
    .C(_2138_),
    .Y(_2140_)
);

FILL FILL_1__7662_ (
);

FILL FILL_3__7588_ (
);

FILL FILL_3__7168_ (
);

FILL FILL_1__13005_ (
);

FILL FILL_0__12838_ (
);

NAND2X1 _12703_ (
    .A(vdd),
    .B(\X[6] [4]),
    .Y(_5743_)
);

FILL FILL_0__12418_ (
);

FILL FILL_1__8867_ (
);

FILL FILL_1__8447_ (
);

FILL FILL_1__8027_ (
);

FILL FILL_2__10772_ (
);

FILL FILL_2__10352_ (
);

OAI21X1 _7097_ (
    .A(_673_),
    .B(_674_),
    .C(_678_),
    .Y(_680_)
);

FILL FILL_3__9314_ (
);

FILL FILL_0__6772_ (
);

NOR2X1 _11095_ (
    .A(_4291_),
    .B(_4292_),
    .Y(_4293_)
);

FILL FILL_3__12984_ (
);

FILL FILL_2__7731_ (
);

FILL FILL_2__7311_ (
);

FILL FILL_3__12144_ (
);

FILL FILL_2__11977_ (
);

FILL FILL_2__11557_ (
);

FILL FILL_0__12591_ (
);

FILL FILL_2__11137_ (
);

FILL FILL_0__12171_ (
);

FILL FILL_0__7977_ (
);

FILL FILL_0__7557_ (
);

NOR3X1 _9663_ (
    .A(_3014_),
    .B(_2982_),
    .C(_3000_),
    .Y(_3015_)
);

FILL FILL_0__7137_ (
);

INVX1 _9243_ (
    .A(_2601_),
    .Y(_2602_)
);

FILL FILL_1__11911_ (
);

FILL FILL_2__8936_ (
);

FILL FILL_2__8516_ (
);

FILL FILL_0__10904_ (
);

FILL FILL254550x169350 (
);

OAI21X1 _13241_ (
    .A(_6262_),
    .B(_6263_),
    .C(_6259_),
    .Y(_6264_)
);

FILL FILL_1__6933_ (
);

FILL FILL_1__6513_ (
);

FILL FILL_3__6439_ (
);

FILL FILL_0__9703_ (
);

FILL FILL_3__7800_ (
);

FILL FILL_1__7718_ (
);

FILL FILL_3__10630_ (
);

OAI21X1 _6788_ (
    .A(_315_),
    .B(_384_),
    .C(_354_),
    .Y(_385_)
);

FILL FILL_2__12095_ (
);

FILL FILL_1__11088_ (
);

AOI22X1 _10786_ (
    .A(vdd),
    .B(\X[5] [0]),
    .C(gnd),
    .D(\X[5] [1]),
    .Y(_3989_)
);

NOR2X1 _10366_ (
    .A(_3561_),
    .B(_3641_),
    .Y(_3642_)
);

FILL FILL_2__9894_ (
);

FILL FILL_2__10828_ (
);

FILL FILL_2__9474_ (
);

FILL FILL_0__11862_ (
);

FILL FILL_2__10408_ (
);

FILL FILL_2__9054_ (
);

FILL FILL_0__11442_ (
);

FILL FILL_0__11022_ (
);

FILL FILL_0__6828_ (
);

NOR2X1 _8934_ (
    .A(_2357_),
    .B(_2356_),
    .Y(_2358_)
);

FILL FILL_0__6408_ (
);

INVX1 _8514_ (
    .A(_1865_),
    .Y(_1952_)
);

FILL FILL_1__7891_ (
);

FILL FILL_1__7471_ (
);

FILL FILL_1__7051_ (
);

FILL FILL_1__13234_ (
);

AOI21X1 _12932_ (
    .A(\X[6] [3]),
    .B(gnd),
    .C(_5966_),
    .Y(_5969_)
);

FILL FILL_0__12647_ (
);

FILL FILL_0__12227_ (
);

DFFPOSX1 _12512_ (
    .D(_5578_[11]),
    .CLK(clk_bF$buf8),
    .Q(\u_fir_pe6.mul [11])
);

OAI21X1 _9719_ (
    .A(_3056_),
    .B(_3057_),
    .C(_3061_),
    .Y(_3063_)
);

FILL FILL_1__8676_ (
);

FILL FILL_1__8256_ (
);

FILL FILL_2__10581_ (
);

FILL FILL_2__10161_ (
);

FILL FILL_3__9963_ (
);

FILL FILL_3__9543_ (
);

FILL FILL_0__6581_ (
);

FILL FILL_2__6599_ (
);

FILL FILL_2__7960_ (
);

FILL FILL_2__7540_ (
);

FILL FILL_3__12373_ (
);

FILL FILL_2__7120_ (
);

FILL FILL_2__11786_ (
);

FILL FILL_2__11366_ (
);

FILL FILL_1__10779_ (
);

FILL FILL_1__10359_ (
);

FILL FILL_0__7786_ (
);

AOI22X1 _9892_ (
    .A(\X[4] [0]),
    .B(gnd),
    .C(\X[4] [1]),
    .D(vdd),
    .Y(_3938_)
);

FILL FILL_0__7366_ (
);

INVX1 _9472_ (
    .A(_2774_),
    .Y(_2829_)
);

NOR2X1 _9052_ (
    .A(_2414_),
    .B(_2413_),
    .Y(_3185_[3])
);

FILL FILL_1__11720_ (
);

FILL FILL_1__11300_ (
);

FILL FILL_2__8745_ (
);

FILL FILL_2__8325_ (
);

FILL FILL_3__13158_ (
);

FILL FILL_0__13185_ (
);

AOI21X1 _13050_ (
    .A(_6034_),
    .B(_6037_),
    .C(_6085_),
    .Y(_6086_)
);

FILL FILL_1__6742_ (
);

FILL FILL_3__6668_ (
);

FILL FILL_1__12925_ (
);

FILL FILL_0__9932_ (
);

FILL FILL_0__11918_ (
);

FILL FILL_0__9512_ (
);

FILL FILL_1__7947_ (
);

FILL FILL_1__7527_ (
);

FILL FILL_1__7107_ (
);

INVX1 _6597_ (
    .A(_106_),
    .Y(_197_)
);

FILL FILL_3__8814_ (
);

AND2X2 _10595_ (
    .A(_3859_),
    .B(_3858_),
    .Y(_3978_[5])
);

NAND3X1 _10175_ (
    .A(_3448_),
    .B(_3447_),
    .C(_3449_),
    .Y(_3454_)
);

FILL FILL_2__6811_ (
);

FILL FILL_3__11644_ (
);

FILL FILL_3__11224_ (
);

FILL FILL253350x219750 (
);

FILL FILL_2__10637_ (
);

FILL FILL_2__9283_ (
);

FILL FILL_0__11671_ (
);

FILL FILL_2__10217_ (
);

FILL FILL_0__11251_ (
);

FILL FILL_0__6637_ (
);

OR2X2 _8743_ (
    .A(_2175_),
    .B(_2173_),
    .Y(_2177_)
);

AOI21X1 _8323_ (
    .A(_1757_),
    .B(_1759_),
    .C(_1750_),
    .Y(_1763_)
);

FILL FILL_1__7280_ (
);

FILL FILL_3__12849_ (
);

FILL FILL_3__12009_ (
);

FILL FILL_1__13043_ (
);

FILL FILL_0__12876_ (
);

NAND3X1 _12741_ (
    .A(_5774_),
    .B(_5775_),
    .C(_5780_),
    .Y(_5781_)
);

FILL FILL_0__12456_ (
);

FILL FILL_0__12036_ (
);

NAND2X1 _12321_ (
    .A(_5425_),
    .B(_5428_),
    .Y(_5572_[2])
);

NAND2X1 _9948_ (
    .A(gnd),
    .B(\X[4] [2]),
    .Y(_3230_)
);

NAND2X1 _9528_ (
    .A(_2882_),
    .B(_2878_),
    .Y(_2884_)
);

NAND3X1 _9108_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf1 ),
    .C(_2466_),
    .Y(_2469_)
);

FILL FILL_1__8485_ (
);

FILL FILL_1__8065_ (
);

FILL FILL_2__10390_ (
);

FILL FILL_3__9772_ (
);

OAI21X1 _13106_ (
    .A(_5884_),
    .B(_6058_),
    .C(_6102_),
    .Y(_6140_)
);

FILL FILL_0__6390_ (
);

FILL FILL_2__11175_ (
);

FILL FILL_1__10588_ (
);

FILL FILL_1__10168_ (
);

FILL FILL_0__7595_ (
);

FILL FILL_0__7175_ (
);

INVX1 _9281_ (
    .A(_2639_),
    .Y(_2640_)
);

FILL FILL_2__8554_ (
);

FILL FILL_0__10942_ (
);

FILL FILL_2__8134_ (
);

FILL FILL_0__10522_ (
);

FILL FILL_0__10102_ (
);

FILL FILL_1__6971_ (
);

FILL FILL_1__6551_ (
);

FILL FILL_2__13321_ (
);

FILL FILL_3__6897_ (
);

FILL FILL_1__12734_ (
);

FILL FILL_1__12314_ (
);

FILL FILL_0__9741_ (
);

FILL FILL_2__9759_ (
);

FILL FILL_2__9339_ (
);

FILL FILL_0__9321_ (
);

FILL FILL_0__11727_ (
);

FILL FILL_0__11307_ (
);

FILL FILL_1__7756_ (
);

FILL FILL_1__7336_ (
);

FILL FILL_3__8203_ (
);

FILL FILL_3__11873_ (
);

FILL FILL_2__6620_ (
);

FILL FILL_3__11453_ (
);

FILL FILL_2__10866_ (
);

FILL FILL_2__10446_ (
);

FILL FILL_2__9092_ (
);

FILL FILL_0__11480_ (
);

FILL FILL_2__10026_ (
);

FILL FILL_0__11060_ (
);

FILL FILL_1__9902_ (
);

FILL FILL_3__9408_ (
);

FILL FILL_0__6866_ (
);

DFFPOSX1 _8972_ (
    .D(\X[2] [3]),
    .CLK(clk_bF$buf28),
    .Q(\X[3] [3])
);

FILL FILL_0__6446_ (
);

AND2X2 _8552_ (
    .A(_1988_),
    .B(_1985_),
    .Y(_1989_)
);

NAND2X1 _8132_ (
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_2283_)
);

FILL FILL_1__10800_ (
);

NAND2X1 _11189_ (
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4386_)
);

FILL FILL_2__7825_ (
);

FILL FILL_3__12658_ (
);

FILL FILL_2__7405_ (
);

FILL FILL_3__12238_ (
);

FILL FILL_1__13272_ (
);

AOI21X1 _12970_ (
    .A(_5922_),
    .B(_5928_),
    .C(_6003_),
    .Y(_6007_)
);

FILL FILL_0__12685_ (
);

FILL FILL_0__12265_ (
);

NAND3X1 _12550_ (
    .A(_6367_),
    .B(_5592_),
    .C(_5588_),
    .Y(_5593_)
);

OAI22X1 _12130_ (
    .A(_5199_),
    .B(_5087_),
    .C(_4807_),
    .D(_5198_),
    .Y(_5246_)
);

INVX1 _9757_ (
    .A(_3096_),
    .Y(_3100_)
);

NAND2X1 _9337_ (
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_2695_)
);

FILL FILL_1__8294_ (
);

FILL FILL_3__9161_ (
);

NOR2X1 _13335_ (
    .A(_6356_),
    .B(_6299_),
    .Y(_6371_[1])
);

FILL FILL253650x111750 (
);

FILL FILL_1__6607_ (
);

FILL FILL_1__9499_ (
);

FILL FILL_1__9079_ (
);

FILL FILL_1__10397_ (
);

NAND3X1 _9090_ (
    .A(_2419_),
    .B(_2436_),
    .C(_2439_),
    .Y(_2452_)
);

FILL FILL_2__8783_ (
);

FILL FILL_2__8363_ (
);

FILL FILL_3__13196_ (
);

FILL FILL_0__10331_ (
);

FILL FILL_2__12189_ (
);

NAND2X1 _7823_ (
    .A(_1337_),
    .B(_1336_),
    .Y(_1338_)
);

INVX1 _7403_ (
    .A(_864_),
    .Y(_924_)
);

FILL FILL_1__6780_ (
);

FILL FILL_2__13130_ (
);

FILL FILL_0__8189_ (
);

FILL FILL_1__12963_ (
);

FILL FILL_3__11509_ (
);

FILL FILL_1__12543_ (
);

FILL FILL_1__12123_ (
);

FILL FILL_2__9988_ (
);

FILL FILL_0__9970_ (
);

FILL FILL_0__9550_ (
);

FILL FILL_2__9568_ (
);

FILL FILL_0__11956_ (
);

FILL FILL_0__9130_ (
);

FILL FILL_2__9148_ (
);

NAND2X1 _11821_ (
    .A(_4869_),
    .B(_4940_),
    .Y(_4941_)
);

FILL FILL_0__11536_ (
);

NAND2X1 _11401_ (
    .A(_4590_),
    .B(_4593_),
    .Y(_4594_)
);

FILL FILL_0__11116_ (
);

OR2X2 _8608_ (
    .A(_1974_),
    .B(_2044_),
    .Y(_2045_)
);

FILL FILL_1__7985_ (
);

FILL FILL_1__7565_ (
);

FILL FILL_1__7145_ (
);

FILL FILL_1__13328_ (
);

FILL FILL_3__8852_ (
);

FILL FILL_3__8432_ (
);

NOR3X1 _12606_ (
    .A(_5632_),
    .B(_5599_),
    .C(_5644_),
    .Y(_5647_)
);

FILL FILL_3__8012_ (
);

FILL FILL_2__10675_ (
);

FILL FILL_2__10255_ (
);

FILL FILL_1__9711_ (
);

FILL FILL_3__9637_ (
);

FILL FILL_0__6675_ (
);

OR2X2 _8781_ (
    .A(_2211_),
    .B(_2212_),
    .Y(_2213_)
);

NOR2X1 _8361_ (
    .A(_1798_),
    .B(_1800_),
    .Y(_2390_[6])
);

FILL FILL_2__7634_ (
);

FILL FILL_1__13081_ (
);

FILL FILL_0__12074_ (
);

FILL FILL253050x205350 (
);

FILL FILL_2__12821_ (
);

FILL FILL_2__12401_ (
);

NAND2X1 _9986_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf1 ),
    .Y(_3267_)
);

INVX1 _9566_ (
    .A(_2920_),
    .Y(_2921_)
);

NAND3X1 _9146_ (
    .A(_2444_),
    .B(_2502_),
    .C(_2506_),
    .Y(_2507_)
);

FILL FILL_1__11814_ (
);

FILL FILL_0__8821_ (
);

FILL FILL_2__8839_ (
);

FILL FILL_0__8401_ (
);

FILL FILL_2__8419_ (
);

FILL FILL_0__10807_ (
);

FILL FILL_3__9390_ (
);

FILL FILL_0__13279_ (
);

NAND2X1 _13144_ (
    .A(_6176_),
    .B(_6175_),
    .Y(_6177_)
);

FILL FILL_1__6836_ (
);

FILL FILL_1__6416_ (
);

FILL FILL_0__9606_ (
);

FILL FILL_3__10953_ (
);

FILL FILL_3__10113_ (
);

FILL FILL_2__8592_ (
);

FILL FILL_0__10980_ (
);

FILL FILL_2__8172_ (
);

FILL FILL_0__10560_ (
);

FILL FILL_0__10140_ (
);

FILL FILL_3__8908_ (
);

AND2X2 _7632_ (
    .A(_1111_),
    .B(_1107_),
    .Y(_1150_)
);

DFFPOSX1 _7212_ (
    .D(_790_[13]),
    .CLK(clk_bF$buf32),
    .Q(\Y[1] [13])
);

AND2X2 _10689_ (
    .A(_3946_),
    .B(_3952_),
    .Y(_3953_)
);

AOI21X1 _10269_ (
    .A(_3458_),
    .B(_3460_),
    .C(_3546_),
    .Y(_3547_)
);

FILL FILL_2__6905_ (
);

FILL FILL_3__11738_ (
);

FILL FILL_1__12772_ (
);

FILL FILL_3__11318_ (
);

FILL FILL_1__12352_ (
);

FILL FILL_2__9797_ (
);

FILL FILL_2__9377_ (
);

FILL FILL_0__11765_ (
);

DFFPOSX1 _11630_ (
    .D(_4781_[6]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [6])
);

FILL FILL_0__11345_ (
);

NAND3X1 _11210_ (
    .A(_4404_),
    .B(_4405_),
    .C(_4406_),
    .Y(_4407_)
);

NOR2X1 _8837_ (
    .A(\u_fir_pe2.rYin [5]),
    .B(\u_fir_pe2.mul [5]),
    .Y(_2262_)
);

AOI21X1 _8417_ (
    .A(_1855_),
    .B(_1854_),
    .C(_1853_),
    .Y(_1856_)
);

FILL FILL_1__7794_ (
);

FILL FILL_1__7374_ (
);

FILL FILL_1__13137_ (
);

AND2X2 _12835_ (
    .A(_5873_),
    .B(_5869_),
    .Y(_6375_[7])
);

AND2X2 _12415_ (
    .A(_5514_),
    .B(_5517_),
    .Y(_5519_)
);

FILL FILL_1__8579_ (
);

FILL FILL_1__8159_ (
);

FILL FILL_3__11071_ (
);

FILL FILL_2__10484_ (
);

FILL FILL_2__10064_ (
);

FILL FILL_1__9940_ (
);

FILL FILL_1__9520_ (
);

FILL FILL_1__9100_ (
);

FILL FILL_3__9026_ (
);

FILL FILL_0__6484_ (
);

AOI21X1 _8590_ (
    .A(_1947_),
    .B(_1949_),
    .C(_2026_),
    .Y(_2027_)
);

NAND2X1 _8170_ (
    .A(_2375_),
    .B(_1612_),
    .Y(_1613_)
);

FILL FILL_2__7863_ (
);

FILL FILL_3__12696_ (
);

FILL FILL_2__7443_ (
);

FILL FILL_2__7023_ (
);

FILL FILL_2__11689_ (
);

FILL FILL_2__11269_ (
);

AND2X2 _6903_ (
    .A(_487_),
    .B(_491_),
    .Y(_499_)
);

FILL FILL_2__12630_ (
);

FILL FILL_2__12210_ (
);

FILL FILL_0__7689_ (
);

OR2X2 _9795_ (
    .A(_3132_),
    .B(_3137_),
    .Y(_3139_)
);

FILL FILL_0__7269_ (
);

INVX1 _9375_ (
    .A(_2713_),
    .Y(_2733_)
);

FILL FILL_1__11203_ (
);

FILL FILL_2__8648_ (
);

FILL FILL_0__8630_ (
);

FILL FILL_2__8228_ (
);

FILL FILL_0__8210_ (
);

FILL FILL_0__10616_ (
);

NAND3X1 _10901_ (
    .A(_4097_),
    .B(_4091_),
    .C(_4095_),
    .Y(_4102_)
);

FILL FILL_0__13088_ (
);

DFFPOSX1 _13373_ (
    .D(\Y[6] [11]),
    .CLK(clk_bF$buf50),
    .Q(\u_fir_pe7.rYin [11])
);

FILL FILL_1__6645_ (
);

FILL FILL_2__13415_ (
);

FILL FILL_1__12828_ (
);

FILL FILL_1__12408_ (
);

FILL FILL254550x32550 (
);

FILL FILL_0__9415_ (
);

FILL FILL_3__7512_ (
);

FILL FILL_3__10342_ (
);

NAND3X1 _7861_ (
    .A(_1359_),
    .B(_1369_),
    .C(_1372_),
    .Y(_1375_)
);

NAND2X1 _7441_ (
    .A(vdd),
    .B(\X[1] [4]),
    .Y(_961_)
);

NAND2X1 _7021_ (
    .A(_613_),
    .B(_610_),
    .Y(_796_[13])
);

OR2X2 _10498_ (
    .A(_3771_),
    .B(_3748_),
    .Y(_3772_)
);

AOI22X1 _10078_ (
    .A(vdd),
    .B(\X[4]_5_bF$buf3 ),
    .C(_3347_),
    .D(_3349_),
    .Y(_3358_)
);

FILL FILL_3__11967_ (
);

FILL FILL_2__6714_ (
);

FILL FILL_3__11547_ (
);

FILL FILL_1__12581_ (
);

FILL FILL_3__11127_ (
);

FILL FILL_1__12161_ (
);

FILL FILL_0__11994_ (
);

FILL FILL_2__9186_ (
);

FILL FILL_0__11574_ (
);

FILL FILL_0__11154_ (
);

FILL FILL_2__11901_ (
);

NAND2X1 _8646_ (
    .A(_2063_),
    .B(_2060_),
    .Y(_2082_)
);

NAND2X1 _8226_ (
    .A(_2294_),
    .B(_1666_),
    .Y(_1667_)
);

FILL FILL_1__7183_ (
);

FILL FILL_2__7919_ (
);

FILL FILL_0__7901_ (
);

FILL FILL_0__12779_ (
);

FILL FILL_3__8470_ (
);

NAND3X1 _12644_ (
    .A(_5680_),
    .B(_5684_),
    .C(_5648_),
    .Y(_5685_)
);

FILL FILL_0__12359_ (
);

NOR3X1 _12224_ (
    .A(_5284_),
    .B(_5286_),
    .C(_5334_),
    .Y(_5338_)
);

FILL FILL_0__13300_ (
);

FILL FILL_1__8388_ (
);

FILL FILL_2__10293_ (
);

FILL FILL_3__9255_ (
);

OAI22X1 _13009_ (
    .A(_5594_),
    .B(_6041_),
    .C(_6042_),
    .D(_6044_),
    .Y(_6045_)
);

FILL FILL_2__7672_ (
);

FILL FILL_3__12085_ (
);

FILL FILL_2__11498_ (
);

FILL FILL_2__11078_ (
);

OAI21X1 _6712_ (
    .A(_308_),
    .B(_309_),
    .C(_304_),
    .Y(_310_)
);

FILL FILL_0__7498_ (
);

FILL FILL_0__7078_ (
);

NAND2X1 _9184_ (
    .A(gnd),
    .B(\X[3] [3]),
    .Y(_2544_)
);

FILL FILL_3__10818_ (
);

FILL FILL_1__11852_ (
);

FILL FILL_1__11432_ (
);

FILL FILL_1__11012_ (
);

FILL FILL_2__8877_ (
);

FILL FILL_2__8457_ (
);

FILL FILL_0__10845_ (
);

DFFPOSX1 _10710_ (
    .D(_3978_[3]),
    .CLK(clk_bF$buf44),
    .Q(\Y[5] [3])
);

FILL FILL_0__10425_ (
);

FILL FILL_2__8037_ (
);

FILL FILL_0__10005_ (
);

INVX1 _13182_ (
    .A(\u_fir_pe7.rYin [1]),
    .Y(_6211_)
);

NAND2X1 _7917_ (
    .A(_1427_),
    .B(_1426_),
    .Y(_1593_[15])
);

FILL FILL_1__6874_ (
);

FILL FILL_1__6454_ (
);

FILL FILL_2__13224_ (
);

FILL FILL_1__12637_ (
);

FILL FILL_1__12217_ (
);

FILL FILL_0__9644_ (
);

FILL FILL_3__7741_ (
);

FILL FILL_0__9224_ (
);

AOI22X1 _11915_ (
    .A(_4869_),
    .B(_4940_),
    .C(_4943_),
    .D(_4939_),
    .Y(_5034_)
);

FILL FILL_1__7659_ (
);

FILL FILL_1__8600_ (
);

FILL FILL_3__8946_ (
);

FILL FILL_3__8526_ (
);

AOI21X1 _7670_ (
    .A(\X[1] [3]),
    .B(gnd),
    .C(_1184_),
    .Y(_1187_)
);

DFFPOSX1 _7250_ (
    .D(_796_[11]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.mul [11])
);

FILL FILL_2__6943_ (
);

FILL FILL_2__6523_ (
);

FILL FILL_1__12390_ (
);

FILL FILL_2__10769_ (
);

FILL FILL_2__10349_ (
);

FILL FILL_0__11383_ (
);

FILL FILL_1__9805_ (
);

FILL FILL_2__11710_ (
);

FILL FILL_0__6769_ (
);

NOR2X1 _8875_ (
    .A(_2287_),
    .B(_2286_),
    .Y(_2299_)
);

AOI21X1 _8455_ (
    .A(_1875_),
    .B(_1877_),
    .C(_1892_),
    .Y(_1893_)
);

INVX1 _8035_ (
    .A(\u_fir_pe1.rYin [12]),
    .Y(_1539_)
);

FILL FILL_1__10703_ (
);

FILL FILL_0__7710_ (
);

FILL FILL_2__7728_ (
);

FILL FILL_2__7308_ (
);

FILL FILL_1__13175_ (
);

NAND2X1 _12873_ (
    .A(_5906_),
    .B(_5910_),
    .Y(_5911_)
);

FILL FILL_0__12588_ (
);

FILL FILL_0__12168_ (
);

OAI21X1 _12453_ (
    .A(_5544_),
    .B(_5547_),
    .C(_5554_),
    .Y(_5557_)
);

OAI21X1 _12033_ (
    .A(_4917_),
    .B(_5150_),
    .C(_5064_),
    .Y(_5151_)
);

FILL FILL_2__12915_ (
);

FILL FILL_1__8197_ (
);

FILL FILL_1__11908_ (
);

FILL FILL_0__8915_ (
);

FILL FILL_3__9484_ (
);

INVX1 _13238_ (
    .A(\u_fir_pe7.mul [7]),
    .Y(_6261_)
);

FILL FILL_2__7481_ (
);

FILL FILL_2__7061_ (
);

AND2X2 _6941_ (
    .A(_535_),
    .B(_532_),
    .Y(_536_)
);

NAND3X1 _6521_ (
    .A(_121_),
    .B(_54_),
    .C(_57_),
    .Y(_122_)
);

FILL FILL_1__11661_ (
);

FILL FILL_3__10207_ (
);

FILL FILL_1__11241_ (
);

FILL FILL_2__8686_ (
);

FILL FILL_2__8266_ (
);

FILL FILL_0__10654_ (
);

FILL FILL_3__13099_ (
);

FILL FILL_0__10234_ (
);

NAND3X1 _7726_ (
    .A(_1223_),
    .B(_1227_),
    .C(_1230_),
    .Y(_1243_)
);

NAND2X1 _7306_ (
    .A(vdd),
    .B(\X[1] [1]),
    .Y(_828_)
);

FILL FILL_1__6683_ (
);

FILL FILL_2__13033_ (
);

FILL FILL_1__12866_ (
);

FILL FILL_1__12446_ (
);

FILL FILL_1__12026_ (
);

FILL FILL_3__7970_ (
);

FILL FILL_0__9453_ (
);

FILL FILL_0__11859_ (
);

FILL FILL_0__9033_ (
);

OAI21X1 _11724_ (
    .A(_4845_),
    .B(_4844_),
    .C(_4811_),
    .Y(_4846_)
);

FILL FILL_0__11439_ (
);

FILL FILL_0__11019_ (
);

AOI21X1 _11304_ (
    .A(_4445_),
    .B(_4479_),
    .C(_4498_),
    .Y(_4499_)
);

FILL FILL_0__12800_ (
);

FILL FILL_1__7888_ (
);

FILL FILL_1__7468_ (
);

FILL FILL_3__10380_ (
);

FILL FILL_1__7048_ (
);

FILL FILL_3__8755_ (
);

NOR2X1 _12929_ (
    .A(_5897_),
    .B(_5900_),
    .Y(_5966_)
);

DFFPOSX1 _12509_ (
    .D(_5578_[8]),
    .CLK(clk_bF$buf22),
    .Q(\u_fir_pe6.mul [8])
);

FILL FILL_2__6752_ (
);

FILL FILL_3__11165_ (
);

FILL FILL_2__10998_ (
);

FILL FILL_2__10578_ (
);

FILL FILL_2__10158_ (
);

FILL FILL_0__11192_ (
);

FILL FILL_1__9614_ (
);

FILL FILL_0__6998_ (
);

FILL FILL_0__6578_ (
);

NAND2X1 _8684_ (
    .A(_1925_),
    .B(_1999_),
    .Y(_2119_)
);

NAND3X1 _8264_ (
    .A(_1620_),
    .B(_1700_),
    .C(_1704_),
    .Y(_1705_)
);

FILL FILL_1__10932_ (
);

FILL FILL_1__10512_ (
);

FILL FILL_2__7957_ (
);

FILL FILL_2__7537_ (
);

FILL FILL_2__7117_ (
);

NAND2X1 _12682_ (
    .A(_5720_),
    .B(_5721_),
    .Y(_5722_)
);

FILL FILL_0__12397_ (
);

OAI21X1 _12262_ (
    .A(_5087_),
    .B(_5374_),
    .C(_5353_),
    .Y(_5375_)
);

FILL FILL_3__13311_ (
);

FILL FILL_2__12724_ (
);

FILL FILL_2__12304_ (
);

NOR2X1 _9889_ (
    .A(_3877_),
    .B(_3898_),
    .Y(_3908_)
);

AOI21X1 _9469_ (
    .A(_2816_),
    .B(_2814_),
    .C(_2786_),
    .Y(_2826_)
);

NAND3X1 _9049_ (
    .A(_2411_),
    .B(_3177_),
    .C(_2410_),
    .Y(_2412_)
);

FILL FILL_1__11717_ (
);

FILL FILL_0__8724_ (
);

FILL FILL_3__6821_ (
);

FILL FILL_0__8304_ (
);

FILL FILL_3__6401_ (
);

AOI21X1 _13047_ (
    .A(_6010_),
    .B(_6016_),
    .C(_6082_),
    .Y(_6083_)
);

FILL FILL_1__6739_ (
);

FILL FILL254250x226950 (
);

FILL FILL_2__7290_ (
);

FILL FILL_0__9929_ (
);

FILL FILL_0__9509_ (
);

FILL FILL_3__7606_ (
);

AOI21X1 _6750_ (
    .A(_259_),
    .B(_261_),
    .C(_347_),
    .Y(_348_)
);

FILL FILL_1__11890_ (
);

FILL FILL_3__10436_ (
);

FILL FILL_1__11470_ (
);

FILL FILL_1__11050_ (
);

FILL FILL_2__8495_ (
);

FILL FILL_0__10883_ (
);

FILL FILL_0__10463_ (
);

FILL FILL_2__8075_ (
);

FILL FILL_0__10043_ (
);

AND2X2 _7955_ (
    .A(_1460_),
    .B(_1459_),
    .Y(_1587_[4])
);

NAND3X1 _7535_ (
    .A(_1050_),
    .B(_1049_),
    .C(_1053_),
    .Y(_1054_)
);

AND2X2 _7115_ (
    .A(_677_),
    .B(_687_),
    .Y(_698_)
);

FILL FILL_1__6492_ (
);

FILL FILL_2__13262_ (
);

FILL FILL_2__6808_ (
);

FILL FILL_1__12675_ (
);

FILL FILL_1__12255_ (
);

FILL FILL_0__9682_ (
);

FILL FILL_0__9262_ (
);

OAI21X1 _11953_ (
    .A(_4989_),
    .B(_4986_),
    .C(_5071_),
    .Y(_5072_)
);

FILL FILL_0__11668_ (
);

OAI21X1 _11533_ (
    .A(_4709_),
    .B(_4710_),
    .C(_4714_),
    .Y(_4717_)
);

FILL FILL_0__11248_ (
);

NAND3X1 _11113_ (
    .A(gnd),
    .B(\X[5] [6]),
    .C(_4310_),
    .Y(_4311_)
);

FILL FILL_1__7697_ (
);

FILL FILL_1__7277_ (
);

FILL FILL_3__8564_ (
);

AOI21X1 _12738_ (
    .A(_5765_),
    .B(_5764_),
    .C(_5715_),
    .Y(_5778_)
);

FILL FILL_3__8144_ (
);

INVX1 _12318_ (
    .A(_5422_),
    .Y(_5426_)
);

FILL FILL_2__6981_ (
);

FILL FILL_2__6561_ (
);

FILL FILL_3__11394_ (
);

FILL FILL_2__10387_ (
);

FILL FILL_1__9423_ (
);

FILL FILL_3__9349_ (
);

FILL FILL_0__6387_ (
);

AOI21X1 _8493_ (
    .A(_1840_),
    .B(_1843_),
    .C(_1849_),
    .Y(_1931_)
);

NOR2X1 _8073_ (
    .A(_1574_),
    .B(_1517_),
    .Y(_1589_[1])
);

FILL FILL_1__10321_ (
);

FILL FILL_2__7766_ (
);

FILL FILL_2__7346_ (
);

FILL FILL_3__12179_ (
);

DFFPOSX1 _12491_ (
    .D(\Y[7] [6]),
    .CLK(clk_bF$buf8),
    .Q(\u_fir_pe6.rYin [6])
);

AOI21X1 _12071_ (
    .A(_5113_),
    .B(_5187_),
    .C(_5186_),
    .Y(_5188_)
);

OAI22X1 _6806_ (
    .A(_254_),
    .B(_401_),
    .C(_324_),
    .D(_402_),
    .Y(_403_)
);

FILL FILL_2__12953_ (
);

FILL FILL_2__12533_ (
);

FILL FILL_2__12113_ (
);

OR2X2 _9698_ (
    .A(_3038_),
    .B(_3043_),
    .Y(_3045_)
);

INVX1 _9278_ (
    .A(_2631_),
    .Y(_2637_)
);

FILL FILL_1__11946_ (
);

FILL FILL_1__11526_ (
);

FILL FILL_1__11106_ (
);

FILL FILL_0__8533_ (
);

FILL FILL_0__10939_ (
);

FILL FILL_0__10519_ (
);

INVX1 _10804_ (
    .A(_4006_),
    .Y(_4007_)
);

INVX1 _13276_ (
    .A(_6298_),
    .Y(_6300_)
);

FILL FILL_2__9912_ (
);

FILL FILL_1__6968_ (
);

FILL FILL_1__6548_ (
);

FILL FILL_2__13318_ (
);

FILL FILL_0__9738_ (
);

FILL FILL_3__7835_ (
);

FILL FILL_0__9318_ (
);

FILL FILL_3__10665_ (
);

FILL FILL_0__10692_ (
);

FILL FILL_0__10272_ (
);

AND2X2 _7764_ (
    .A(_1273_),
    .B(_1279_),
    .Y(_1280_)
);

NOR3X1 _7344_ (
    .A(_850_),
    .B(_817_),
    .C(_862_),
    .Y(_865_)
);

FILL FILL_2__13071_ (
);

FILL FILL_2__6617_ (
);

FILL FILL_1__12064_ (
);

FILL FILL_0__9491_ (
);

FILL FILL_0__11897_ (
);

FILL FILL_0__9071_ (
);

FILL FILL_2__9089_ (
);

NAND3X1 _11762_ (
    .A(_4878_),
    .B(_4864_),
    .C(_4882_),
    .Y(_4883_)
);

FILL FILL_0__11477_ (
);

FILL FILL_0__11057_ (
);

NAND2X1 _11342_ (
    .A(_4533_),
    .B(_4536_),
    .Y(_4537_)
);

FILL FILL_3__12811_ (
);

FILL FILL_2__11804_ (
);

DFFPOSX1 _8969_ (
    .D(\X[2] [0]),
    .CLK(clk_bF$buf51),
    .Q(\X[3] [0])
);

INVX1 _8549_ (
    .A(_1980_),
    .Y(_1986_)
);

DFFPOSX1 _8129_ (
    .D(_1593_[13]),
    .CLK(clk_bF$buf13),
    .Q(\u_fir_pe1.mul [13])
);

FILL FILL_1__7086_ (
);

FILL FILL_0__7804_ (
);

INVX1 _9910_ (
    .A(_3192_),
    .Y(_3193_)
);

FILL FILL_1__13269_ (
);

FILL FILL_3__8793_ (
);

NAND3X1 _12967_ (
    .A(_5922_),
    .B(_5928_),
    .C(_6003_),
    .Y(_6004_)
);

FILL FILL_3__8373_ (
);

NAND3X1 _12547_ (
    .A(_5579_),
    .B(_5584_),
    .C(_5582_),
    .Y(_5590_)
);

OAI21X1 _12127_ (
    .A(_5209_),
    .B(_5211_),
    .C(_5205_),
    .Y(_5243_)
);

FILL FILL_0__13203_ (
);

FILL FILL_2__6790_ (
);

FILL FILL_2__10196_ (
);

FILL FILL_1__9652_ (
);

FILL FILL_1__9232_ (
);

FILL FILL_3__9998_ (
);

FILL FILL_3__9578_ (
);

FILL FILL_1__10970_ (
);

FILL FILL_1__10550_ (
);

FILL FILL_1__10130_ (
);

FILL FILL_2__7995_ (
);

FILL FILL_2__7575_ (
);

FILL FILL_2__7155_ (
);

AND2X2 _6615_ (
    .A(_145_),
    .B(_149_),
    .Y(_214_)
);

FILL FILL_2__12762_ (
);

FILL FILL_2__12342_ (
);

NAND2X1 _9087_ (
    .A(_2445_),
    .B(_2448_),
    .Y(_2449_)
);

FILL FILL_1__11755_ (
);

FILL FILL_1__11335_ (
);

FILL FILL_0__8762_ (
);

FILL FILL_0__8342_ (
);

FILL FILL_0__10328_ (
);

NAND2X1 _10613_ (
    .A(_3875_),
    .B(_3874_),
    .Y(_3876_)
);

NAND2X1 _13085_ (
    .A(_6119_),
    .B(_6118_),
    .Y(_6120_)
);

FILL FILL_2__9721_ (
);

FILL FILL_2__9301_ (
);

FILL FILL_1__6777_ (
);

FILL FILL_2__13127_ (
);

FILL FILL_0__9967_ (
);

FILL FILL_0__9547_ (
);

FILL FILL_0__9127_ (
);

NAND2X1 _11818_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf1 ),
    .Y(_4938_)
);

FILL FILL_3__10894_ (
);

FILL FILL_3__10054_ (
);

FILL FILL_0__10081_ (
);

FILL FILL_1__8923_ (
);

FILL FILL_1__8503_ (
);

FILL FILL_3__8849_ (
);

AOI21X1 _7993_ (
    .A(_1492_),
    .B(_1495_),
    .C(_1494_),
    .Y(_1496_)
);

AND2X2 _7573_ (
    .A(_1091_),
    .B(_1087_),
    .Y(_1593_[7])
);

AND2X2 _7153_ (
    .A(_732_),
    .B(_735_),
    .Y(_737_)
);

FILL FILL_2__6846_ (
);

FILL FILL_3__11679_ (
);

FILL FILL_2__6426_ (
);

FILL FILL_3__11259_ (
);

FILL FILL_1__12293_ (
);

AND2X2 _11991_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf3 ),
    .Y(_5109_)
);

NAND2X1 _11571_ (
    .A(\u_fir_pe5.rYin [15]),
    .B(\u_fir_pe5.mul [15]),
    .Y(_4754_)
);

FILL FILL_0__11286_ (
);

NAND3X1 _11151_ (
    .A(_4288_),
    .B(_4345_),
    .C(_4346_),
    .Y(_4349_)
);

FILL FILL_1__9708_ (
);

OAI21X1 _8778_ (
    .A(_2178_),
    .B(_2203_),
    .C(_2202_),
    .Y(_2210_)
);

AOI21X1 _8358_ (
    .A(_1714_),
    .B(_1720_),
    .C(_1797_),
    .Y(_1798_)
);

FILL FILL_1__10606_ (
);

FILL FILL_0__7613_ (
);

FILL FILL_1__13078_ (
);

FILL FILL254550x205350 (
);

OAI21X1 _12776_ (
    .A(_6357_),
    .B(_5814_),
    .C(_5806_),
    .Y(_5815_)
);

FILL FILL_3__8182_ (
);

NAND2X1 _12356_ (
    .A(_5459_),
    .B(_5454_),
    .Y(_5460_)
);

FILL FILL_3__13405_ (
);

FILL FILL_2__12818_ (
);

FILL FILL_0__13012_ (
);

FILL FILL_0__8818_ (
);

FILL FILL_3__6915_ (
);

FILL FILL_1__9461_ (
);

FILL FILL_1__9041_ (
);

FILL FILL_2__7384_ (
);

OAI21X1 _6844_ (
    .A(_440_),
    .B(_439_),
    .C(_438_),
    .Y(_441_)
);

NOR2X1 _6424_ (
    .A(_24_),
    .B(_25_),
    .Y(_26_)
);

FILL FILL_2__12991_ (
);

FILL FILL_2__12571_ (
);

FILL FILL_2__12151_ (
);

FILL FILL_1__11984_ (
);

FILL FILL_1__11564_ (
);

FILL FILL_1__11144_ (
);

FILL FILL_0__8571_ (
);

FILL FILL_2__8589_ (
);

FILL FILL_0__10977_ (
);

FILL FILL_0__8151_ (
);

FILL FILL_2__8169_ (
);

FILL FILL_0__10557_ (
);

OAI21X1 _10842_ (
    .A(_4766_),
    .B(_4003_),
    .C(_4006_),
    .Y(_4044_)
);

NOR2X1 _10422_ (
    .A(_3693_),
    .B(_3697_),
    .Y(_3698_)
);

FILL FILL_0__10137_ (
);

NAND3X1 _10002_ (
    .A(_3273_),
    .B(_3280_),
    .C(_3282_),
    .Y(_3283_)
);

FILL FILL_2__9950_ (
);

FILL FILL_2__9530_ (
);

FILL FILL_2__9110_ (
);

NAND3X1 _7629_ (
    .A(_1119_),
    .B(_1137_),
    .C(_1133_),
    .Y(_1147_)
);

DFFPOSX1 _7209_ (
    .D(_790_[10]),
    .CLK(clk_bF$buf1),
    .Q(\Y[1] [10])
);

FILL FILL_1__6586_ (
);

FILL FILL_1__12769_ (
);

FILL FILL_1__12349_ (
);

FILL FILL_0__9776_ (
);

FILL FILL_0__9356_ (
);

FILL FILL_3__7453_ (
);

DFFPOSX1 _11627_ (
    .D(_4779_[3]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.mul [3])
);

FILL FILL_3__7033_ (
);

OAI21X1 _11207_ (
    .A(_4010_),
    .B(_4401_),
    .C(_4403_),
    .Y(_4404_)
);

FILL FILL_0__12703_ (
);

FILL FILL_3__10283_ (
);

FILL FILL_1__8732_ (
);

FILL FILL_1__8312_ (
);

FILL FILL_3__8238_ (
);

NAND3X1 _7382_ (
    .A(_898_),
    .B(_902_),
    .C(_866_),
    .Y(_903_)
);

FILL FILL_2__6655_ (
);

FILL FILL_3__11488_ (
);

INVX1 _11380_ (
    .A(_4570_),
    .Y(_4574_)
);

FILL FILL_0__11095_ (
);

FILL FILL_1__9937_ (
);

FILL FILL_1__9517_ (
);

FILL FILL_2__11842_ (
);

FILL FILL_2__11422_ (
);

FILL FILL_2__11002_ (
);

OAI21X1 _8587_ (
    .A(_2023_),
    .B(_2022_),
    .C(_2021_),
    .Y(_2024_)
);

NAND2X1 _8167_ (
    .A(_1607_),
    .B(_1603_),
    .Y(_1610_)
);

FILL FILL_1__10835_ (
);

FILL FILL_1__10415_ (
);

FILL FILL_0__7842_ (
);

FILL FILL_0__7422_ (
);

FILL FILL_0__7002_ (
);

NAND2X1 _12585_ (
    .A(_5625_),
    .B(_5626_),
    .Y(_5627_)
);

AND2X2 _12165_ (
    .A(_5269_),
    .B(_5273_),
    .Y(_5281_)
);

FILL FILL_2__8801_ (
);

FILL FILL_2__12627_ (
);

FILL FILL_2__12207_ (
);

FILL FILL_0__13241_ (
);

FILL FILL_0__8627_ (
);

FILL FILL_0__8207_ (
);

FILL FILL_1__9690_ (
);

FILL FILL_1__9270_ (
);

FILL FILL_3__9196_ (
);

FILL FILL_2__7193_ (
);

FILL FILL_3__7929_ (
);

AOI22X1 _6653_ (
    .A(_87_),
    .B(_158_),
    .C(_161_),
    .D(_157_),
    .Y(_252_)
);

FILL FILL_2__12380_ (
);

FILL FILL_1__11793_ (
);

FILL FILL_1__11373_ (
);

FILL FILL_0__8380_ (
);

FILL FILL_2__8398_ (
);

FILL FILL_0__10786_ (
);

NOR2X1 _10651_ (
    .A(\u_fir_pe4.rYin [10]),
    .B(\u_fir_pe4.mul [10]),
    .Y(_3915_)
);

FILL FILL_0__10366_ (
);

NAND2X1 _10231_ (
    .A(\X[4] [4]),
    .B(vdd),
    .Y(_3509_)
);

OAI21X1 _7858_ (
    .A(_1370_),
    .B(_1371_),
    .C(_1323_),
    .Y(_1372_)
);

INVX1 _7438_ (
    .A(_957_),
    .Y(_958_)
);

NAND2X1 _7018_ (
    .A(_589_),
    .B(_588_),
    .Y(_611_)
);

FILL FILL_1__6395_ (
);

FILL FILL_2__13165_ (
);

FILL FILL_1__12998_ (
);

FILL FILL_1__12578_ (
);

FILL FILL_1__12158_ (
);

FILL FILL_0__9585_ (
);

FILL FILL_3__7682_ (
);

FILL FILL_0__9165_ (
);

OAI21X1 _11856_ (
    .A(_4975_),
    .B(_4970_),
    .C(_4898_),
    .Y(_4976_)
);

NOR2X1 _11436_ (
    .A(_4624_),
    .B(_4623_),
    .Y(_4775_[1])
);

AOI22X1 _11016_ (
    .A(vdd),
    .B(\X[5] [7]),
    .C(\X[5] [3]),
    .D(vdd),
    .Y(_4215_)
);

FILL FILL_3__12905_ (
);

FILL FILL_0__12932_ (
);

FILL FILL_1__8541_ (
);

FILL FILL_3__8887_ (
);

FILL FILL_3__8467_ (
);

FILL FILL_3__8047_ (
);

OAI21X1 _7191_ (
    .A(_762_),
    .B(_765_),
    .C(_772_),
    .Y(_775_)
);

FILL FILL_2__6884_ (
);

FILL FILL_2__6464_ (
);

FILL FILL_1__9746_ (
);

FILL FILL_1__9326_ (
);

FILL FILL_2__11651_ (
);

FILL FILL_2__11231_ (
);

NAND2X1 _8396_ (
    .A(vdd),
    .B(\X[2] [4]),
    .Y(_1835_)
);

FILL FILL_1__10644_ (
);

FILL FILL_1__10224_ (
);

CLKBUF1 CLKBUF1_insert50 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert51 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert52 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert53 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert54 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf15)
);

FILL FILL_2__7669_ (
);

FILL FILL_0__7651_ (
);

CLKBUF1 CLKBUF1_insert55 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert56 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert57 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert58 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert59 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf10)
);

OR2X2 _12394_ (
    .A(_5493_),
    .B(_5497_),
    .Y(_5498_)
);

FILL FILL_2__8610_ (
);

FILL FILL_3__13023_ (
);

OAI21X1 _6709_ (
    .A(_225_),
    .B(_230_),
    .C(_229_),
    .Y(_307_)
);

FILL FILL_2__12856_ (
);

FILL FILL_2__12436_ (
);

FILL FILL_2__12016_ (
);

FILL FILL_0__13050_ (
);

FILL FILL_1__11849_ (
);

FILL FILL_1__11429_ (
);

FILL FILL_1__11009_ (
);

FILL FILL_0__8856_ (
);

FILL FILL_0__8436_ (
);

FILL FILL_3__6533_ (
);

DFFPOSX1 _10707_ (
    .D(_3977_[0]),
    .CLK(clk_bF$buf45),
    .Q(\Y[5] [0])
);

FILL FILL_0__8016_ (
);

NAND2X1 _13179_ (
    .A(_6209_),
    .B(_6208_),
    .Y(_6375_[15])
);

FILL FILL_2__9815_ (
);

FILL FILL_1__7812_ (
);

FILL FILL_3__7318_ (
);

AND2X2 _6882_ (
    .A(Xin_5_bF$buf3),
    .B(gnd),
    .Y(_478_)
);

OAI21X1 _6462_ (
    .A(_63_),
    .B(_62_),
    .C(_29_),
    .Y(_64_)
);

FILL FILL_3__10988_ (
);

FILL FILL_3__10148_ (
);

FILL FILL_1__11182_ (
);

FILL FILL_0__10595_ (
);

NAND3X1 _10880_ (
    .A(_4069_),
    .B(_4080_),
    .C(_4076_),
    .Y(_4081_)
);

NAND2X1 _10460_ (
    .A(_3730_),
    .B(_3734_),
    .Y(_3735_)
);

FILL FILL_0__10175_ (
);

NAND2X1 _10040_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf0 ),
    .Y(_3320_)
);

FILL FILL_2__10922_ (
);

FILL FILL_2__10502_ (
);

NOR2X1 _7667_ (
    .A(_1115_),
    .B(_1118_),
    .Y(_1184_)
);

DFFPOSX1 _7247_ (
    .D(_796_[8]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.mul [8])
);

FILL FILL_2__13394_ (
);

FILL FILL_0__6922_ (
);

FILL FILL_0__6502_ (
);

FILL FILL_1__12387_ (
);

FILL FILL_0__9394_ (
);

NAND3X1 _11665_ (
    .A(_4783_),
    .B(_4787_),
    .C(_4785_),
    .Y(_4788_)
);

AOI21X1 _11245_ (
    .A(_4426_),
    .B(_4422_),
    .C(_4367_),
    .Y(_4441_)
);

FILL FILL_2__11707_ (
);

FILL FILL_0__12741_ (
);

FILL FILL_0__12321_ (
);

FILL FILL_0__7707_ (
);

NOR2X1 _9813_ (
    .A(_3155_),
    .B(_3149_),
    .Y(_3157_)
);

FILL FILL_1__8770_ (
);

FILL FILL_1__8350_ (
);

FILL FILL_0__13106_ (
);

FILL FILL_2__6693_ (
);

FILL FILL_2__10099_ (
);

FILL FILL_1__9975_ (
);

FILL FILL_1__9555_ (
);

FILL FILL_1__9135_ (
);

FILL FILL_2__11880_ (
);

FILL FILL_2__11460_ (
);

FILL FILL_2__11040_ (
);

FILL FILL_1__10873_ (
);

FILL FILL_1__10453_ (
);

FILL FILL_1__10033_ (
);

FILL FILL_2__7898_ (
);

FILL FILL_0__7880_ (
);

FILL FILL_0__7460_ (
);

FILL FILL_2__7478_ (
);

FILL FILL_2__7058_ (
);

FILL FILL_0__7040_ (
);

FILL FILL_3__13252_ (
);

AND2X2 _6938_ (
    .A(_523_),
    .B(_519_),
    .Y(_533_)
);

NAND3X1 _6518_ (
    .A(_54_),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

FILL FILL_2__12665_ (
);

FILL FILL_2__12245_ (
);

FILL FILL_1__11658_ (
);

FILL FILL_1__11238_ (
);

FILL FILL_0__8665_ (
);

FILL FILL_3__6762_ (
);

FILL FILL_0__8245_ (
);

NAND3X1 _10936_ (
    .A(_4124_),
    .B(_4133_),
    .C(_4135_),
    .Y(_4136_)
);

NAND2X1 _10516_ (
    .A(_3787_),
    .B(_3788_),
    .Y(_3789_)
);

FILL FILL_2__9624_ (
);

FILL FILL_2__9204_ (
);

FILL FILL_1__7621_ (
);

FILL FILL_3__7547_ (
);

OAI21X1 _6691_ (
    .A(_207_),
    .B(_204_),
    .C(_289_),
    .Y(_290_)
);

FILL FILL_3__10377_ (
);

FILL FILL_1__8826_ (
);

FILL FILL_1__8406_ (
);

FILL FILL_2__10311_ (
);

AND2X2 _7896_ (
    .A(_1405_),
    .B(_1402_),
    .Y(_1409_)
);

AOI21X1 _7476_ (
    .A(_983_),
    .B(_982_),
    .C(_933_),
    .Y(_996_)
);

INVX1 _7056_ (
    .A(_640_),
    .Y(_644_)
);

FILL FILL_0__6731_ (
);

FILL FILL_2__6749_ (
);

FILL FILL_1__12196_ (
);

INVX1 _11894_ (
    .A(_5012_),
    .Y(_5013_)
);

INVX1 _11474_ (
    .A(\u_fir_pe5.rYin [6]),
    .Y(_4658_)
);

FILL FILL_0__11189_ (
);

NAND3X1 _11054_ (
    .A(_4251_),
    .B(_4252_),
    .C(_4250_),
    .Y(_4253_)
);

FILL FILL_3__12523_ (
);

FILL FILL_3__12103_ (
);

FILL FILL_2__11936_ (
);

FILL FILL_0__12970_ (
);

FILL FILL_2__11516_ (
);

FILL FILL_0__12550_ (
);

FILL FILL_0__12130_ (
);

FILL FILL_1__10929_ (
);

FILL FILL_1__10509_ (
);

FILL FILL_0__7936_ (
);

FILL FILL_0__7516_ (
);

NAND2X1 _9622_ (
    .A(_2973_),
    .B(_2975_),
    .Y(_2976_)
);

OAI21X1 _9202_ (
    .A(_2560_),
    .B(_2561_),
    .C(_2559_),
    .Y(_2562_)
);

INVX1 _12679_ (
    .A(_5718_),
    .Y(_5719_)
);

NOR2X1 _12259_ (
    .A(_5368_),
    .B(_5372_),
    .Y(_5578_[12])
);

FILL FILL_0__13335_ (
);

INVX1 _13200_ (
    .A(\u_fir_pe7.rYin [3]),
    .Y(_6227_)
);

FILL FILL_3__6818_ (
);

FILL FILL_1__9784_ (
);

FILL FILL_1__9364_ (
);

FILL FILL_1__10682_ (
);

FILL FILL_1__10262_ (
);

FILL FILL_2__7287_ (
);

AOI21X1 _6747_ (
    .A(_344_),
    .B(_343_),
    .C(_342_),
    .Y(_345_)
);

FILL FILL_2__12894_ (
);

FILL FILL_2__12054_ (
);

FILL FILL_1__11887_ (
);

FILL FILL_1__11467_ (
);

FILL FILL_1__11047_ (
);

FILL FILL_0__8894_ (
);

FILL FILL_3__6991_ (
);

FILL FILL_0__8474_ (
);

DFFPOSX1 _10745_ (
    .D(\Y[4] [14]),
    .CLK(clk_bF$buf26),
    .Q(\u_fir_pe4.rYin [14])
);

FILL FILL_0__8054_ (
);

NAND2X1 _10325_ (
    .A(_3601_),
    .B(_3597_),
    .Y(_3602_)
);

FILL FILL_2__9433_ (
);

FILL FILL_0__11821_ (
);

FILL FILL_2__9013_ (
);

FILL FILL_0__11401_ (
);

FILL FILL_1__6489_ (
);

FILL FILL_2__13259_ (
);

FILL FILL_1__7850_ (
);

FILL FILL_1__7430_ (
);

FILL FILL_1__7010_ (
);

FILL FILL_0__9679_ (
);

FILL FILL_3__7776_ (
);

FILL FILL_0__9259_ (
);

FILL FILL_0__12606_ (
);

FILL FILL_1__8635_ (
);

FILL FILL_1__8215_ (
);

FILL FILL_2__10960_ (
);

FILL FILL_2__10540_ (
);

FILL FILL_2__10120_ (
);

NAND3X1 _7285_ (
    .A(_797_),
    .B(_802_),
    .C(_800_),
    .Y(_808_)
);

FILL FILL_3__9922_ (
);

FILL FILL_3__9502_ (
);

FILL FILL_2__6978_ (
);

FILL FILL_0__6960_ (
);

FILL FILL_2__6558_ (
);

FILL FILL_0__6540_ (
);

NAND3X1 _11283_ (
    .A(_4408_),
    .B(_4411_),
    .C(_4478_),
    .Y(_4479_)
);

FILL FILL_3__12752_ (
);

FILL FILL_3__12332_ (
);

FILL FILL_2__11745_ (
);

FILL FILL_2__11325_ (
);

FILL FILL_1__10318_ (
);

FILL FILL_0__7745_ (
);

DFFPOSX1 _9851_ (
    .D(\X[3]_5_bF$buf3 ),
    .CLK(clk_bF$buf51),
    .Q(\X[4] [5])
);

FILL FILL_0__7325_ (
);

OAI21X1 _9431_ (
    .A(_2713_),
    .B(_2787_),
    .C(_2734_),
    .Y(_2788_)
);

INVX1 _9011_ (
    .A(_3091_),
    .Y(_3101_)
);

DFFPOSX1 _12488_ (
    .D(\Y[7] [3]),
    .CLK(clk_bF$buf11),
    .Q(\u_fir_pe6.rYin [3])
);

OAI22X1 _12068_ (
    .A(_5036_),
    .B(_5183_),
    .C(_5106_),
    .D(_5184_),
    .Y(_5185_)
);

FILL FILL_2__8704_ (
);

FILL FILL_3__13117_ (
);

FILL FILL_0__13144_ (
);

FILL FILL_1__6701_ (
);

FILL FILL_1__9593_ (
);

FILL FILL_1__9173_ (
);

FILL FILL_2__9909_ (
);

FILL FILL_1__10491_ (
);

FILL FILL_1__10071_ (
);

FILL FILL_2__7096_ (
);

FILL FILL_1__7906_ (
);

FILL FILL_3__13290_ (
);

OR2X2 _6976_ (
    .A(_569_),
    .B(_565_),
    .Y(_570_)
);

NAND2X1 _6556_ (
    .A(gnd),
    .B(Xin_5_bF$buf2),
    .Y(_156_)
);

FILL FILL_2__12283_ (
);

FILL FILL_1__11696_ (
);

FILL FILL_1__11276_ (
);

FILL FILL_0__8283_ (
);

FILL FILL_0__10689_ (
);

AOI21X1 _10974_ (
    .A(_4086_),
    .B(_4090_),
    .C(_4054_),
    .Y(_4174_)
);

FILL FILL_3__6380_ (
);

NOR2X1 _10554_ (
    .A(\u_fir_pe4.rYin [1]),
    .B(\u_fir_pe4.mul [1]),
    .Y(_3823_)
);

FILL FILL_0__10269_ (
);

NAND2X1 _10134_ (
    .A(\X[4] [2]),
    .B(vdd),
    .Y(_3413_)
);

FILL FILL_2__9662_ (
);

FILL FILL_2__9242_ (
);

FILL FILL_0__11210_ (
);

FILL FILL_2__13068_ (
);

INVX1 _8702_ (
    .A(_2109_),
    .Y(_2137_)
);

FILL FILL_0__9488_ (
);

FILL FILL_0__9068_ (
);

AOI21X1 _11759_ (
    .A(_4874_),
    .B(_4876_),
    .C(_4867_),
    .Y(_4880_)
);

AOI21X1 _11339_ (
    .A(_4472_),
    .B(_4476_),
    .C(_4446_),
    .Y(_4534_)
);

FILL FILL_1__13002_ (
);

FILL FILL_0__12835_ (
);

INVX1 _12700_ (
    .A(_5739_),
    .Y(_5740_)
);

FILL FILL_0__12415_ (
);

NAND2X1 _9907_ (
    .A(gnd),
    .B(\X[4] [0]),
    .Y(_3190_)
);

FILL FILL_1__8864_ (
);

FILL FILL_1__8444_ (
);

FILL FILL_1__8024_ (
);

NAND2X1 _7094_ (
    .A(_677_),
    .B(_672_),
    .Y(_678_)
);

FILL FILL_3__9731_ (
);

FILL FILL_3__9311_ (
);

FILL FILL_2__6787_ (
);

INVX2 _11092_ (
    .A(gnd),
    .Y(_4290_)
);

FILL FILL_1__9649_ (
);

FILL FILL_1__9229_ (
);

FILL FILL_2__11974_ (
);

FILL FILL_2__11554_ (
);

FILL FILL_2__11134_ (
);

NAND2X1 _8299_ (
    .A(\X[2] [2]),
    .B(vdd),
    .Y(_1739_)
);

FILL FILL_1__10967_ (
);

FILL FILL_1__10547_ (
);

FILL FILL_1__10127_ (
);

FILL FILL_0__7974_ (
);

FILL FILL_0__7554_ (
);

NAND2X1 _9660_ (
    .A(_3011_),
    .B(_3010_),
    .Y(_3012_)
);

FILL FILL_0__7134_ (
);

AOI21X1 _9240_ (
    .A(_2563_),
    .B(_2567_),
    .C(_2529_),
    .Y(_2599_)
);

INVX1 _12297_ (
    .A(_5403_),
    .Y(_5409_)
);

FILL FILL_2__8933_ (
);

FILL FILL_2__8513_ (
);

FILL FILL_0__10901_ (
);

FILL FILL_2__12759_ (
);

FILL FILL_2__12339_ (
);

FILL FILL_1__6930_ (
);

FILL FILL_1__6510_ (
);

FILL FILL_0__8759_ (
);

FILL FILL_3__6856_ (
);

FILL FILL_0__8339_ (
);

FILL FILL_3__6436_ (
);

FILL FILL_0__9700_ (
);

FILL FILL_2__9718_ (
);

FILL FILL_1__7715_ (
);

OAI21X1 _6785_ (
    .A(_301_),
    .B(_381_),
    .C(_364_),
    .Y(_382_)
);

FILL FILL_2__12092_ (
);

FILL FILL_1__11085_ (
);

FILL FILL_0__10498_ (
);

INVX1 _10783_ (
    .A(_3985_),
    .Y(_3986_)
);

NAND2X1 _10363_ (
    .A(_3638_),
    .B(_3568_),
    .Y(_3640_)
);

FILL FILL_0__10078_ (
);

FILL FILL_3__11832_ (
);

FILL FILL_2__10825_ (
);

FILL FILL_2__9891_ (
);

FILL FILL_2__9471_ (
);

FILL FILL_2__10405_ (
);

FILL FILL_2__9051_ (
);

FILL FILL_2__13297_ (
);

FILL FILL_0__6825_ (
);

INVX1 _8931_ (
    .A(\u_fir_pe2.mul [14]),
    .Y(_2355_)
);

FILL FILL_0__6405_ (
);

OAI21X1 _8511_ (
    .A(_1935_),
    .B(_1939_),
    .C(_1942_),
    .Y(_1949_)
);

FILL FILL_0__9297_ (
);

NAND2X1 _11988_ (
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5106_)
);

FILL FILL_3__7394_ (
);

NOR2X1 _11568_ (
    .A(_4751_),
    .B(_4750_),
    .Y(_4775_[14])
);

NAND3X1 _11148_ (
    .A(_4300_),
    .B(_4331_),
    .C(_4336_),
    .Y(_4346_)
);

FILL FILL_3__12617_ (
);

FILL FILL_1__13231_ (
);

FILL FILL_0__12644_ (
);

FILL FILL_0__12224_ (
);

NAND2X1 _9716_ (
    .A(_3060_),
    .B(_3055_),
    .Y(_3061_)
);

FILL FILL_1__8673_ (
);

FILL FILL_1__8253_ (
);

FILL FILL_3__8179_ (
);

FILL FILL_0__13009_ (
);

FILL FILL_2__6596_ (
);

FILL FILL_1__9458_ (
);

FILL FILL_3__12790_ (
);

FILL FILL_1__9038_ (
);

FILL FILL_2__11783_ (
);

FILL FILL_2__11363_ (
);

FILL FILL_1__10776_ (
);

FILL FILL_1__10356_ (
);

FILL FILL_0__7783_ (
);

FILL FILL_0__7363_ (
);

FILL FILL254550x100950 (
);

FILL FILL_2__8742_ (
);

FILL FILL_2__8322_ (
);

FILL FILL_2__12988_ (
);

FILL FILL_2__12568_ (
);

FILL FILL_2__12148_ (
);

FILL FILL_0__13182_ (
);

FILL FILL_0__8568_ (
);

FILL FILL_0__8148_ (
);

NAND2X1 _10839_ (
    .A(_4034_),
    .B(_4037_),
    .Y(_4041_)
);

AOI21X1 _10419_ (
    .A(_3643_),
    .B(_3646_),
    .C(_3694_),
    .Y(_3695_)
);

FILL FILL_1__12922_ (
);

FILL FILL_2__9947_ (
);

FILL FILL_2__9527_ (
);

FILL FILL_0__11915_ (
);

FILL FILL_2__9107_ (
);

FILL FILL_1__7944_ (
);

FILL FILL_1__7524_ (
);

FILL FILL_1__7104_ (
);

OAI21X1 _6594_ (
    .A(_193_),
    .B(_188_),
    .C(_116_),
    .Y(_194_)
);

NOR2X1 _10592_ (
    .A(_3856_),
    .B(_3855_),
    .Y(_3857_)
);

OAI21X1 _10172_ (
    .A(_3446_),
    .B(_3450_),
    .C(_3412_),
    .Y(_3451_)
);

FILL FILL_1__8729_ (
);

FILL FILL_1__8309_ (
);

FILL FILL_3__11221_ (
);

FILL FILL_2__10634_ (
);

FILL FILL_2__9280_ (
);

FILL FILL_2__10214_ (
);

NOR3X1 _7799_ (
    .A(_1102_),
    .B(_1270_),
    .C(_1213_),
    .Y(_1314_)
);

OAI21X1 _7379_ (
    .A(_895_),
    .B(_896_),
    .C(_881_),
    .Y(_900_)
);

FILL FILL_0__6634_ (
);

NAND3X1 _8740_ (
    .A(_2155_),
    .B(_2172_),
    .C(_2171_),
    .Y(_2174_)
);

NAND3X1 _8320_ (
    .A(_1750_),
    .B(_1757_),
    .C(_1759_),
    .Y(_1760_)
);

FILL FILL_1__12099_ (
);

NAND2X1 _11797_ (
    .A(_4913_),
    .B(_4915_),
    .Y(_4917_)
);

AOI21X1 _11377_ (
    .A(_4542_),
    .B(_4544_),
    .C(_4570_),
    .Y(_4571_)
);

FILL FILL_3__12846_ (
);

FILL FILL_3__12426_ (
);

FILL FILL_3__12006_ (
);

FILL FILL_1__13040_ (
);

FILL FILL_2__11839_ (
);

FILL FILL_0__12873_ (
);

FILL FILL_2__11419_ (
);

FILL FILL_0__12453_ (
);

FILL FILL_0__12033_ (
);

FILL FILL_0__7839_ (
);

INVX1 _9945_ (
    .A(_3226_),
    .Y(_3227_)
);

FILL FILL_0__7419_ (
);

NAND3X1 _9525_ (
    .A(_2798_),
    .B(_2874_),
    .C(_2806_),
    .Y(_2881_)
);

NAND2X1 _9105_ (
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_2466_)
);

FILL FILL_1__8482_ (
);

FILL FILL_1__8062_ (
);

FILL FILL_0__13238_ (
);

OAI21X1 _13103_ (
    .A(_6090_),
    .B(_6131_),
    .C(_6130_),
    .Y(_6137_)
);

FILL FILL_1__9687_ (
);

FILL FILL_1__9267_ (
);

FILL FILL_2__11172_ (
);

FILL FILL_1__10585_ (
);

FILL FILL_1__10165_ (
);

FILL FILL_0__7592_ (
);

FILL FILL_0__7172_ (
);

FILL FILL_3__10912_ (
);

FILL FILL_2__8551_ (
);

FILL FILL_2__12797_ (
);

FILL FILL_2__12377_ (
);

FILL FILL_0__8797_ (
);

FILL FILL_0__8377_ (
);

FILL FILL_3__6474_ (
);

INVX1 _10648_ (
    .A(\u_fir_pe4.rYin [10]),
    .Y(_3912_)
);

NAND2X1 _10228_ (
    .A(\X[4] [3]),
    .B(gnd),
    .Y(_3506_)
);

FILL FILL_1__12731_ (
);

FILL FILL_1__12311_ (
);

FILL FILL_2__9756_ (
);

FILL FILL_2__9336_ (
);

FILL FILL_0__11724_ (
);

FILL FILL_0__11304_ (
);

FILL FILL_1__7753_ (
);

FILL FILL_1__7333_ (
);

FILL FILL_3__7259_ (
);

FILL FILL_0__12929_ (
);

FILL FILL_3__8620_ (
);

FILL FILL_3__10089_ (
);

FILL FILL_1__8538_ (
);

FILL FILL_2__10863_ (
);

FILL FILL_2__10443_ (
);

FILL FILL_2__10023_ (
);

NAND2X1 _7188_ (
    .A(_769_),
    .B(_771_),
    .Y(_772_)
);

FILL FILL_3__9825_ (
);

FILL FILL_3__9405_ (
);

FILL FILL_0__6863_ (
);

FILL FILL_0__6443_ (
);

NOR2X1 _11186_ (
    .A(_4117_),
    .B(_4306_),
    .Y(_4383_)
);

FILL FILL_2__7822_ (
);

FILL FILL_2__7402_ (
);

FILL FILL_2__11648_ (
);

FILL FILL_0__12682_ (
);

FILL FILL_2__11228_ (
);

FILL FILL_0__12262_ (
);

FILL FILL_0__7648_ (
);

NAND2X1 _9754_ (
    .A(_3096_),
    .B(_3097_),
    .Y(_3098_)
);

INVX1 _9334_ (
    .A(_2691_),
    .Y(_2692_)
);

FILL FILL_1__8291_ (
);

FILL FILL_2__8607_ (
);

FILL FILL_0__13047_ (
);

NOR2X1 _13332_ (
    .A(\u_fir_pe7.rYin [0]),
    .B(\u_fir_pe7.mul [0]),
    .Y(_6355_)
);

FILL FILL_1__6604_ (
);

FILL FILL254250x176550 (
);

FILL FILL_1__9496_ (
);

FILL FILL_1__9076_ (
);

FILL FILL_1__10394_ (
);

FILL FILL_1__7809_ (
);

FILL FILL_3__10301_ (
);

FILL FILL_2__8780_ (
);

FILL FILL_2__8360_ (
);

FILL FILL_3__13193_ (
);

AND2X2 _6879_ (
    .A(_473_),
    .B(_416_),
    .Y(_475_)
);

NAND3X1 _6459_ (
    .A(_28_),
    .B(_45_),
    .C(_48_),
    .Y(_61_)
);

FILL FILL_2__12186_ (
);

AOI21X1 _7820_ (
    .A(_1212_),
    .B(_1204_),
    .C(_1282_),
    .Y(_1335_)
);

NAND3X1 _7400_ (
    .A(_850_),
    .B(_914_),
    .C(_915_),
    .Y(_921_)
);

FILL FILL_1__11179_ (
);

FILL FILL_0__8186_ (
);

NAND2X1 _10877_ (
    .A(gnd),
    .B(\X[5] [3]),
    .Y(_4078_)
);

NAND2X1 _10457_ (
    .A(_3728_),
    .B(_3704_),
    .Y(_3732_)
);

OAI21X1 _10037_ (
    .A(_3316_),
    .B(_3317_),
    .C(_3315_),
    .Y(_3318_)
);

FILL FILL_3__11926_ (
);

FILL FILL_1__12960_ (
);

FILL FILL_1__12540_ (
);

FILL FILL_1__12120_ (
);

FILL FILL_2__9985_ (
);

FILL FILL_2__10919_ (
);

FILL FILL_2__9565_ (
);

FILL FILL_0__11953_ (
);

FILL FILL_2__9145_ (
);

FILL FILL_0__11533_ (
);

FILL FILL_0__11113_ (
);

FILL FILL_0__6919_ (
);

AOI21X1 _8605_ (
    .A(_2030_),
    .B(_2025_),
    .C(_1977_),
    .Y(_2042_)
);

FILL FILL_1__7982_ (
);

FILL FILL_1__7562_ (
);

FILL FILL_1__7142_ (
);

FILL FILL_3__7488_ (
);

FILL FILL_1__13325_ (
);

FILL FILL_0__12738_ (
);

OAI21X1 _12603_ (
    .A(_5632_),
    .B(_5644_),
    .C(_5638_),
    .Y(_5645_)
);

FILL FILL_0__12318_ (
);

FILL FILL_1__8767_ (
);

FILL FILL_1__8347_ (
);

FILL FILL_2__10672_ (
);

FILL FILL_2__10252_ (
);

FILL FILL_0__6672_ (
);

FILL FILL_3__12884_ (
);

FILL FILL_2__7631_ (
);

FILL FILL_3__12044_ (
);

FILL FILL_2__11877_ (
);

FILL FILL_2__11457_ (
);

FILL FILL_2__11037_ (
);

FILL FILL_0__12071_ (
);

FILL FILL_0__7877_ (
);

OAI21X1 _9983_ (
    .A(_3966_),
    .B(_3262_),
    .C(_3263_),
    .Y(_3264_)
);

FILL FILL_0__7457_ (
);

OAI22X1 _9563_ (
    .A(_2624_),
    .B(_2626_),
    .C(_2710_),
    .D(_2535_),
    .Y(_2918_)
);

FILL FILL_0__7037_ (
);

OAI21X1 _9143_ (
    .A(_2499_),
    .B(_2500_),
    .C(_2460_),
    .Y(_2504_)
);

FILL FILL_1__11811_ (
);

FILL FILL_2__8836_ (
);

FILL FILL_2__8416_ (
);

FILL FILL_0__10804_ (
);

FILL FILL_0__13276_ (
);

NOR2X1 _13141_ (
    .A(_5814_),
    .B(_6041_),
    .Y(_6174_)
);

FILL FILL_1__6833_ (
);

FILL FILL_1__6413_ (
);

FILL FILL_3__6759_ (
);

FILL FILL_0__9603_ (
);

FILL FILL_3__7700_ (
);

FILL FILL_1__7618_ (
);

FILL FILL_3__10530_ (
);

NAND3X1 _6688_ (
    .A(_135_),
    .B(_274_),
    .C(_279_),
    .Y(_287_)
);

NOR2X1 _10686_ (
    .A(_3947_),
    .B(_3949_),
    .Y(_3950_)
);

AOI21X1 _10266_ (
    .A(_3543_),
    .B(_3542_),
    .C(_3541_),
    .Y(_3544_)
);

FILL FILL_2__6902_ (
);

FILL FILL_3__11315_ (
);

FILL FILL_2__9794_ (
);

FILL FILL_2__9374_ (
);

FILL FILL_0__11762_ (
);

FILL FILL_2__10308_ (
);

FILL FILL_0__11342_ (
);

FILL FILL_0__6728_ (
);

INVX1 _8834_ (
    .A(\u_fir_pe2.rYin [5]),
    .Y(_2259_)
);

AND2X2 _8414_ (
    .A(_1831_),
    .B(_1826_),
    .Y(_1853_)
);

FILL FILL_1__7791_ (
);

FILL FILL_1__7371_ (
);

FILL FILL_1__13134_ (
);

FILL FILL_0__12967_ (
);

AOI21X1 _12832_ (
    .A(_5866_),
    .B(_5865_),
    .C(_5767_),
    .Y(_5871_)
);

FILL FILL_0__12547_ (
);

FILL FILL_0__12127_ (
);

NOR2X1 _12412_ (
    .A(\u_fir_pe6.rYin [11]),
    .B(\u_fir_pe6.mul [11]),
    .Y(_5516_)
);

OAI21X1 _9619_ (
    .A(_2970_),
    .B(_2972_),
    .C(_2951_),
    .Y(_2973_)
);

FILL FILL_1__8576_ (
);

FILL FILL_1__8156_ (
);

FILL FILL_2__10481_ (
);

FILL FILL_2__10061_ (
);

FILL FILL_3__9443_ (
);

FILL FILL_3__9023_ (
);

FILL FILL253650x219750 (
);

FILL FILL_2__6499_ (
);

FILL FILL_0__6481_ (
);

FILL FILL_2__7860_ (
);

FILL FILL_3__12693_ (
);

FILL FILL_2__7440_ (
);

FILL FILL_3__12273_ (
);

FILL FILL_2__7020_ (
);

FILL FILL_2__11686_ (
);

FILL FILL_2__11266_ (
);

INVX1 _6900_ (
    .A(_460_),
    .Y(_496_)
);

FILL FILL_1__10679_ (
);

FILL FILL_1__10259_ (
);

FILL FILL_0__7686_ (
);

NOR2X1 _9792_ (
    .A(\u_fir_pe3.rYin [12]),
    .B(\u_fir_pe3.mul [12]),
    .Y(_3136_)
);

FILL FILL_0__7266_ (
);

NAND3X1 _9372_ (
    .A(_2715_),
    .B(_2717_),
    .C(_2719_),
    .Y(_2730_)
);

FILL FILL_1__11200_ (
);

FILL FILL_2__8645_ (
);

FILL FILL_2__8225_ (
);

FILL FILL_0__10613_ (
);

FILL FILL_3__13058_ (
);

FILL FILL_0__13085_ (
);

DFFPOSX1 _13370_ (
    .D(\Y[6] [8]),
    .CLK(clk_bF$buf5),
    .Q(\u_fir_pe7.rYin [8])
);

FILL FILL_1__6642_ (
);

FILL FILL_2__13412_ (
);

FILL FILL_3__6568_ (
);

FILL FILL_1__12825_ (
);

FILL FILL_1__12405_ (
);

FILL FILL_0__9412_ (
);

FILL FILL_0__11818_ (
);

FILL FILL_1__7847_ (
);

FILL FILL_1__7427_ (
);

FILL FILL_1__7007_ (
);

AOI21X1 _6497_ (
    .A(_92_),
    .B(_94_),
    .C(_85_),
    .Y(_98_)
);

FILL FILL_3__8714_ (
);

INVX1 _10495_ (
    .A(_3768_),
    .Y(_3769_)
);

NAND3X1 _10075_ (
    .A(_3343_),
    .B(_3354_),
    .C(_3350_),
    .Y(_3355_)
);

FILL FILL_2__6711_ (
);

FILL FILL_3__11544_ (
);

FILL FILL_2__10957_ (
);

FILL FILL_0__11991_ (
);

FILL FILL_2__10537_ (
);

FILL FILL_2__9183_ (
);

FILL FILL_0__11571_ (
);

FILL FILL_2__10117_ (
);

FILL FILL_0__11151_ (
);

FILL FILL_0__6957_ (
);

FILL FILL_0__6537_ (
);

NAND2X1 _8643_ (
    .A(_2076_),
    .B(_2070_),
    .Y(_2079_)
);

NAND2X1 _8223_ (
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1664_)
);

FILL FILL_1__7180_ (
);

FILL FILL_2__7916_ (
);

FILL FILL_0__12776_ (
);

OAI21X1 _12641_ (
    .A(_5677_),
    .B(_5678_),
    .C(_5663_),
    .Y(_5682_)
);

FILL FILL_0__12356_ (
);

NAND3X1 _12221_ (
    .A(_5293_),
    .B(_5335_),
    .C(_5294_),
    .Y(_5336_)
);

DFFPOSX1 _9848_ (
    .D(\X[3] [2]),
    .CLK(clk_bF$buf42),
    .Q(\X[4] [2])
);

NAND3X1 _9428_ (
    .A(_2783_),
    .B(_2779_),
    .C(_2784_),
    .Y(_2785_)
);

DFFPOSX1 _9008_ (
    .D(_2390_[15]),
    .CLK(clk_bF$buf28),
    .Q(\u_fir_pe2.mul [15])
);

FILL FILL_1__8385_ (
);

FILL FILL_2__10290_ (
);

FILL FILL_3__9672_ (
);

FILL FILL_3__9252_ (
);

NOR3X1 _13006_ (
    .A(_5884_),
    .B(_5711_),
    .C(_5900_),
    .Y(_6042_)
);

FILL FILL_2__11495_ (
);

FILL FILL_2__11075_ (
);

FILL FILL_1__10488_ (
);

FILL FILL_1__10068_ (
);

FILL FILL_0__7495_ (
);

FILL FILL_0__7075_ (
);

NAND2X1 _9181_ (
    .A(_2540_),
    .B(_2532_),
    .Y(_2541_)
);

FILL FILL_3__10815_ (
);

FILL FILL_2__8874_ (
);

FILL FILL_2__8454_ (
);

FILL FILL_0__10842_ (
);

FILL FILL_3__13287_ (
);

FILL FILL_0__10422_ (
);

FILL FILL_2__8034_ (
);

FILL FILL_0__10002_ (
);

NAND2X1 _7914_ (
    .A(_1425_),
    .B(_1419_),
    .Y(_1593_[14])
);

FILL FILL_1__6871_ (
);

FILL FILL_1__6451_ (
);

FILL FILL_2__13221_ (
);

FILL FILL_3__6797_ (
);

FILL FILL_1__12634_ (
);

FILL FILL_1__12214_ (
);

FILL FILL253950x111750 (
);

FILL FILL_0__9641_ (
);

FILL FILL_2__9659_ (
);

FILL FILL_0__9221_ (
);

INVX1 _11912_ (
    .A(_5030_),
    .Y(_5031_)
);

FILL FILL_2__9239_ (
);

FILL FILL_0__11207_ (
);

FILL FILL_1__7656_ (
);

FILL FILL_3__8943_ (
);

FILL FILL_2__6940_ (
);

FILL FILL_3__11773_ (
);

FILL FILL_2__6520_ (
);

FILL FILL_2__10766_ (
);

FILL FILL_2__10346_ (
);

FILL FILL_0__11380_ (
);

FILL FILL_1__9802_ (
);

FILL FILL_3__9728_ (
);

FILL FILL_0__6766_ (
);

NAND3X1 _8872_ (
    .A(_2295_),
    .B(_2292_),
    .C(_2255_),
    .Y(_2296_)
);

AOI21X1 _8452_ (
    .A(_1801_),
    .B(_1879_),
    .C(_1887_),
    .Y(_1890_)
);

AOI21X1 _8032_ (
    .A(_1532_),
    .B(_1523_),
    .C(_1530_),
    .Y(_1535_)
);

FILL FILL_1__10700_ (
);

AOI21X1 _11089_ (
    .A(_4251_),
    .B(_4252_),
    .C(_4209_),
    .Y(_4287_)
);

FILL FILL_2__7725_ (
);

FILL FILL_3__12558_ (
);

FILL FILL_2__7305_ (
);

FILL FILL_3__12138_ (
);

FILL FILL_1__13172_ (
);

AOI21X1 _12870_ (
    .A(_5907_),
    .B(_5905_),
    .C(_5903_),
    .Y(_5908_)
);

FILL FILL_0__12585_ (
);

FILL FILL_0__12165_ (
);

NAND2X1 _12450_ (
    .A(_5551_),
    .B(_5553_),
    .Y(_5554_)
);

AOI21X1 _12030_ (
    .A(_5147_),
    .B(_5146_),
    .C(_5082_),
    .Y(_5148_)
);

FILL FILL_2__12912_ (
);

AND2X2 _9657_ (
    .A(_2987_),
    .B(_2986_),
    .Y(_3009_)
);

AOI21X1 _9237_ (
    .A(_2585_),
    .B(_2593_),
    .C(_2596_),
    .Y(_2597_)
);

FILL FILL_1__8194_ (
);

FILL FILL_1__11905_ (
);

FILL FILL_0__8912_ (
);

FILL FILL_3__9061_ (
);

AND2X2 _13235_ (
    .A(_6258_),
    .B(_6257_),
    .Y(_6369_[6])
);

FILL FILL_1__6927_ (
);

FILL FILL_1__6507_ (
);

FILL FILL_1__9399_ (
);

FILL FILL_1__10297_ (
);

FILL FILL_3__10624_ (
);

FILL FILL253350x205350 (
);

FILL FILL_2__8683_ (
);

FILL FILL_2__8263_ (
);

FILL FILL_0__10651_ (
);

FILL FILL_0__10231_ (
);

FILL FILL_2__12089_ (
);

INVX1 _7723_ (
    .A(_1161_),
    .Y(_1240_)
);

NOR2X1 _7303_ (
    .A(_824_),
    .B(_823_),
    .Y(_825_)
);

FILL FILL_1__6680_ (
);

FILL FILL_2__13030_ (
);

FILL FILL_1__12863_ (
);

FILL FILL_3__11409_ (
);

FILL FILL_1__12443_ (
);

FILL FILL_1__12023_ (
);

FILL FILL_2__9888_ (
);

FILL FILL_2__9468_ (
);

FILL FILL_0__9450_ (
);

FILL FILL_0__11856_ (
);

FILL FILL_0__9030_ (
);

FILL FILL_2__9048_ (
);

NAND3X1 _11721_ (
    .A(_4810_),
    .B(_4827_),
    .C(_4830_),
    .Y(_4843_)
);

FILL FILL_0__11436_ (
);

NAND3X1 _11301_ (
    .A(_4480_),
    .B(_4486_),
    .C(_4444_),
    .Y(_4496_)
);

FILL FILL_0__11016_ (
);

AND2X2 _8928_ (
    .A(_2351_),
    .B(_2350_),
    .Y(_2384_[13])
);

AOI21X1 _8508_ (
    .A(_1945_),
    .B(_1940_),
    .C(_1909_),
    .Y(_1946_)
);

FILL FILL_1__7885_ (
);

FILL FILL_1__7465_ (
);

FILL FILL_1__7045_ (
);

FILL FILL_1__13228_ (
);

AOI21X1 _12926_ (
    .A(_5928_),
    .B(_5929_),
    .C(_5896_),
    .Y(_5963_)
);

FILL FILL_3__8332_ (
);

DFFPOSX1 _12506_ (
    .D(_5578_[5]),
    .CLK(clk_bF$buf22),
    .Q(\u_fir_pe6.mul [5])
);

FILL FILL_3__11582_ (
);

FILL FILL_3__11162_ (
);

FILL FILL_2__10995_ (
);

FILL FILL_2__10575_ (
);

FILL FILL_2__10155_ (
);

FILL FILL_1__9611_ (
);

FILL FILL_3__9957_ (
);

FILL FILL_3__9117_ (
);

FILL FILL_0__6995_ (
);

FILL FILL_0__6575_ (
);

OAI21X1 _8681_ (
    .A(_1668_),
    .B(_1899_),
    .C(_2073_),
    .Y(_2116_)
);

AOI21X1 _8261_ (
    .A(_1697_),
    .B(_1698_),
    .C(_1696_),
    .Y(_1702_)
);

FILL FILL_2__7954_ (
);

FILL FILL_3__12787_ (
);

FILL FILL_2__7534_ (
);

FILL FILL_3__12367_ (
);

FILL FILL_2__7114_ (
);

FILL FILL_0__12394_ (
);

FILL FILL_2__12721_ (
);

FILL FILL_2__12301_ (
);

NAND2X1 _9886_ (
    .A(\X[4] [0]),
    .B(vdd),
    .Y(_3877_)
);

INVX1 _9466_ (
    .A(_2745_),
    .Y(_2823_)
);

NAND2X1 _9046_ (
    .A(_2405_),
    .B(_2408_),
    .Y(_2409_)
);

FILL FILL_1__11714_ (
);

FILL FILL_2__8739_ (
);

FILL FILL_0__8721_ (
);

FILL FILL_2__8319_ (
);

FILL FILL_0__8301_ (
);

FILL FILL_3__9290_ (
);

FILL FILL_0__13179_ (
);

NAND3X1 _13044_ (
    .A(_6075_),
    .B(_6076_),
    .C(_6079_),
    .Y(_6080_)
);

FILL FILL_1__6736_ (
);

FILL FILL_1__12919_ (
);

FILL FILL_0__9926_ (
);

FILL FILL_0__9506_ (
);

FILL FILL_3__10853_ (
);

FILL FILL254250x108150 (
);

FILL FILL_3__10013_ (
);

FILL FILL_2__8492_ (
);

FILL FILL_0__10880_ (
);

FILL FILL_0__10460_ (
);

FILL FILL_2__8072_ (
);

FILL FILL_0__10040_ (
);

FILL FILL_3__8808_ (
);

OAI21X1 _7952_ (
    .A(_1448_),
    .B(_1444_),
    .C(_1457_),
    .Y(_1458_)
);

NAND2X1 _7532_ (
    .A(vdd),
    .B(\X[1]_5_bF$buf2 ),
    .Y(_1051_)
);

OAI21X1 _7112_ (
    .A(_665_),
    .B(_666_),
    .C(_694_),
    .Y(_695_)
);

INVX1 _10589_ (
    .A(\u_fir_pe4.mul [5]),
    .Y(_3854_)
);

NAND3X1 _10169_ (
    .A(_3427_),
    .B(_3441_),
    .C(_3444_),
    .Y(_3448_)
);

FILL FILL_2__6805_ (
);

FILL FILL_1__12672_ (
);

FILL FILL_1__12252_ (
);

FILL FILL_2__9697_ (
);

FILL FILL_2__9277_ (
);

NAND3X1 _11950_ (
    .A(_4917_),
    .B(_5056_),
    .C(_5061_),
    .Y(_5069_)
);

FILL FILL_0__11665_ (
);

NAND2X1 _11530_ (
    .A(_4713_),
    .B(_4708_),
    .Y(_4714_)
);

FILL FILL_0__11245_ (
);

OAI21X1 _11110_ (
    .A(_4225_),
    .B(_4233_),
    .C(_4232_),
    .Y(_4308_)
);

NAND2X1 _8737_ (
    .A(_2157_),
    .B(_2170_),
    .Y(_2171_)
);

NAND3X1 _8317_ (
    .A(gnd),
    .B(\X[2] [4]),
    .C(_1747_),
    .Y(_1757_)
);

FILL FILL_1__7694_ (
);

FILL FILL_1__7274_ (
);

FILL FILL_1__13037_ (
);

FILL FILL_3__8561_ (
);

NAND3X1 _12735_ (
    .A(_5769_),
    .B(_5770_),
    .C(_5771_),
    .Y(_5775_)
);

AND2X2 _12315_ (
    .A(\u_fir_pe6.rYin [2]),
    .B(\u_fir_pe6.mul [2]),
    .Y(_5423_)
);

FILL FILL_1__8899_ (
);

FILL FILL_1__8479_ (
);

FILL FILL_1__8059_ (
);

FILL FILL_2__10384_ (
);

FILL FILL_1__9420_ (
);

FILL FILL_3__9766_ (
);

FILL FILL_3__9346_ (
);

FILL FILL_0__6384_ (
);

NAND2X1 _8490_ (
    .A(_1919_),
    .B(_1927_),
    .Y(_1928_)
);

NOR2X1 _8070_ (
    .A(\u_fir_pe1.rYin [0]),
    .B(\u_fir_pe1.mul [0]),
    .Y(_1573_)
);

FILL FILL_2__7763_ (
);

FILL FILL_2__7343_ (
);

FILL FILL_2__11169_ (
);

NOR2X1 _6803_ (
    .A(_398_),
    .B(_399_),
    .Y(_400_)
);

FILL FILL_2__12950_ (
);

FILL FILL_2__12530_ (
);

FILL FILL_2__12110_ (
);

FILL FILL_0__7589_ (
);

NOR2X1 _9695_ (
    .A(\u_fir_pe3.rYin [3]),
    .B(\u_fir_pe3.mul [3]),
    .Y(_3042_)
);

FILL FILL_0__7169_ (
);

NAND2X1 _9275_ (
    .A(_2632_),
    .B(_2633_),
    .Y(_2634_)
);

FILL FILL_3__10909_ (
);

FILL FILL_1__11943_ (
);

FILL FILL_1__11523_ (
);

FILL FILL_1__11103_ (
);

FILL FILL_0__8950_ (
);

FILL FILL_2__8548_ (
);

FILL FILL_0__8530_ (
);

FILL FILL_0__10936_ (
);

FILL FILL_0__10516_ (
);

NAND2X1 _10801_ (
    .A(_4766_),
    .B(_4003_),
    .Y(_4004_)
);

NAND2X1 _13273_ (
    .A(_6296_),
    .B(_6295_),
    .Y(_6369_[9])
);

FILL FILL_1__6965_ (
);

FILL FILL_1__6545_ (
);

FILL FILL_2__13315_ (
);

FILL FILL_1__12728_ (
);

FILL FILL_1__12308_ (
);

FILL FILL_0__9735_ (
);

FILL FILL_0__9315_ (
);

FILL FILL_3__7412_ (
);

FILL FILL_3__10242_ (
);

OAI21X1 _7761_ (
    .A(_871_),
    .B(_1116_),
    .C(_1270_),
    .Y(_1277_)
);

OAI21X1 _7341_ (
    .A(_850_),
    .B(_862_),
    .C(_856_),
    .Y(_863_)
);

NAND3X1 _10398_ (
    .A(_3595_),
    .B(_3673_),
    .C(_3603_),
    .Y(_3674_)
);

FILL FILL_3__11867_ (
);

FILL FILL_2__6614_ (
);

FILL FILL_3__11027_ (
);

FILL FILL_1__12061_ (
);

FILL FILL_0__11894_ (
);

FILL FILL_2__9086_ (
);

FILL FILL_0__11474_ (
);

FILL FILL_0__11054_ (
);

FILL FILL_2__11801_ (
);

DFFPOSX1 _8966_ (
    .D(_2384_[13]),
    .CLK(clk_bF$buf55),
    .Q(\Y[3] [13])
);

INVX1 _8546_ (
    .A(_1982_),
    .Y(_1983_)
);

DFFPOSX1 _8126_ (
    .D(_1593_[10]),
    .CLK(clk_bF$buf13),
    .Q(\u_fir_pe1.mul [10])
);

FILL FILL_1__7083_ (
);

FILL FILL_2__7819_ (
);

FILL FILL_0__7801_ (
);

FILL FILL_1__13266_ (
);

FILL FILL_3__8790_ (
);

FILL FILL_0__12679_ (
);

NAND3X1 _12964_ (
    .A(_5998_),
    .B(_5999_),
    .C(_6000_),
    .Y(_6001_)
);

FILL FILL_0__12259_ (
);

OAI21X1 _12544_ (
    .A(_5583_),
    .B(_5586_),
    .C(_5579_),
    .Y(_5587_)
);

INVX1 _12124_ (
    .A(_5239_),
    .Y(_5240_)
);

FILL FILL_0__13200_ (
);

FILL FILL_1__8288_ (
);

FILL FILL_2__10193_ (
);

NAND3X1 _13329_ (
    .A(_6346_),
    .B(_6352_),
    .C(_6347_),
    .Y(_6353_)
);

FILL FILL_2__7992_ (
);

FILL FILL_2__7572_ (
);

FILL FILL_2__7152_ (
);

FILL FILL_2__11398_ (
);

INVX1 _6612_ (
    .A(_210_),
    .Y(_211_)
);

FILL FILL_0__7398_ (
);

NAND2X1 _9084_ (
    .A(_2400_),
    .B(_2405_),
    .Y(_2446_)
);

FILL FILL_1__11752_ (
);

FILL FILL_1__11332_ (
);

FILL FILL_2__8777_ (
);

FILL FILL_2__8357_ (
);

FILL FILL_0__10325_ (
);

OAI21X1 _10610_ (
    .A(_3871_),
    .B(_3872_),
    .C(_3868_),
    .Y(_3873_)
);

AOI21X1 _13082_ (
    .A(_5994_),
    .B(_5986_),
    .C(_6064_),
    .Y(_6117_)
);

NAND3X1 _7817_ (
    .A(_1326_),
    .B(_1331_),
    .C(_1330_),
    .Y(_1332_)
);

FILL FILL_1__6774_ (
);

FILL FILL_2__13124_ (
);

FILL FILL_1__12957_ (
);

FILL FILL_1__12537_ (
);

FILL FILL_1__12117_ (
);

FILL FILL_0__9964_ (
);

FILL FILL_0__9544_ (
);

FILL FILL_3__7641_ (
);

FILL FILL_0__9124_ (
);

NAND2X1 _11815_ (
    .A(gnd),
    .B(\X[7] [3]),
    .Y(_4935_)
);

FILL FILL_1__7979_ (
);

FILL FILL_1__7559_ (
);

FILL FILL_3__10471_ (
);

FILL FILL_1__7139_ (
);

FILL FILL_1__8920_ (
);

FILL FILL_1__8500_ (
);

FILL FILL_3__8426_ (
);

NAND2X1 _7990_ (
    .A(_1472_),
    .B(_1484_),
    .Y(_1493_)
);

AOI21X1 _7570_ (
    .A(_1084_),
    .B(_1083_),
    .C(_985_),
    .Y(_1089_)
);

NOR2X1 _7150_ (
    .A(\u_fir_pe0.rYin [11]),
    .B(\u_fir_pe0.mul [11]),
    .Y(_734_)
);

FILL FILL_2__6843_ (
);

FILL FILL_2__6423_ (
);

FILL FILL_3__11256_ (
);

FILL FILL_1__12290_ (
);

FILL FILL_2__10669_ (
);

FILL FILL_2__10249_ (
);

FILL FILL_0__11283_ (
);

FILL FILL_1__9705_ (
);

FILL FILL_0__6669_ (
);

NAND2X1 _8775_ (
    .A(_2207_),
    .B(_2204_),
    .Y(_2390_[13])
);

OAI21X1 _8355_ (
    .A(_1793_),
    .B(_1794_),
    .C(_1792_),
    .Y(_1795_)
);

FILL FILL_1__10603_ (
);

FILL FILL_0__7610_ (
);

FILL FILL_2__7628_ (
);

FILL FILL_1__13075_ (
);

INVX1 _12773_ (
    .A(gnd),
    .Y(_5812_)
);

FILL FILL_0__12068_ (
);

NOR2X1 _12353_ (
    .A(_5455_),
    .B(_5456_),
    .Y(_5457_)
);

FILL FILL_3__13402_ (
);

FILL FILL_2__12815_ (
);

FILL FILL_1__11808_ (
);

FILL FILL_0__8815_ (
);

FILL FILL_3__6912_ (
);

FILL FILL_3__9384_ (
);

INVX1 _13138_ (
    .A(_6145_),
    .Y(_6171_)
);

FILL FILL_2__7381_ (
);

INVX1 _6841_ (
    .A(_383_),
    .Y(_438_)
);

NOR2X1 _6421_ (
    .A(_23_),
    .B(_22_),
    .Y(_794_[3])
);

FILL FILL_1__11981_ (
);

FILL FILL_1__11561_ (
);

FILL FILL_3__10107_ (
);

FILL FILL_1__11141_ (
);

FILL FILL_2__8586_ (
);

FILL FILL_0__10974_ (
);

FILL FILL_2__8166_ (
);

FILL FILL_0__10554_ (
);

FILL FILL_0__10134_ (
);

INVX1 _7626_ (
    .A(_1057_),
    .Y(_1144_)
);

DFFPOSX1 _7206_ (
    .D(_790_[7]),
    .CLK(clk_bF$buf32),
    .Q(\Y[1] [7])
);

FILL FILL_1__6583_ (
);

FILL FILL_1__12766_ (
);

FILL FILL_1__12346_ (
);

FILL FILL_0__9773_ (
);

FILL FILL_3__7870_ (
);

FILL FILL_0__9353_ (
);

FILL FILL_0__11759_ (
);

DFFPOSX1 _11624_ (
    .D(_4776_[0]),
    .CLK(clk_bF$buf50),
    .Q(\u_fir_pe5.mul [0])
);

FILL FILL_3__7030_ (
);

FILL FILL_0__11339_ (
);

NAND2X1 _11204_ (
    .A(\X[5]_5_bF$buf0 ),
    .B(gnd),
    .Y(_4401_)
);

FILL FILL254550x226950 (
);

FILL FILL_0__12700_ (
);

FILL FILL_1__7788_ (
);

FILL FILL_1__7368_ (
);

FILL FILL_3__8655_ (
);

AND2X2 _12829_ (
    .A(_5864_),
    .B(_5867_),
    .Y(_5868_)
);

AND2X2 _12409_ (
    .A(_5511_),
    .B(_5512_),
    .Y(_5572_[10])
);

FILL FILL_2__6652_ (
);

FILL FILL_3__11485_ (
);

FILL FILL_2__10898_ (
);

FILL FILL_2__10478_ (
);

FILL FILL_2__10058_ (
);

FILL FILL_0__11092_ (
);

FILL FILL_1__9934_ (
);

FILL FILL_1__9514_ (
);

FILL FILL_0__6898_ (
);

FILL FILL_0__6478_ (
);

NAND2X1 _8584_ (
    .A(_1985_),
    .B(_1988_),
    .Y(_2021_)
);

NAND3X1 _8164_ (
    .A(_1604_),
    .B(_1606_),
    .C(_1605_),
    .Y(_1607_)
);

FILL FILL_1__10832_ (
);

FILL FILL_1__10412_ (
);

FILL FILL_2__7857_ (
);

FILL FILL_2__7437_ (
);

FILL FILL_2__7017_ (
);

FILL FILL_0__12297_ (
);

NAND3X1 _12582_ (
    .A(_5611_),
    .B(_5623_),
    .C(_5619_),
    .Y(_5624_)
);

INVX1 _12162_ (
    .A(_5242_),
    .Y(_5278_)
);

FILL FILL_3__13211_ (
);

FILL FILL_2__12624_ (
);

FILL FILL_2__12204_ (
);

INVX1 _9789_ (
    .A(\u_fir_pe3.rYin [12]),
    .Y(_3133_)
);

OAI21X1 _9369_ (
    .A(_2726_),
    .B(_2720_),
    .C(_2714_),
    .Y(_2727_)
);

FILL FILL_0__8624_ (
);

FILL FILL_0__8204_ (
);

DFFPOSX1 _13367_ (
    .D(\Y[6] [5]),
    .CLK(clk_bF$buf39),
    .Q(\u_fir_pe7.rYin [5])
);

FILL FILL_1__6639_ (
);

FILL FILL_2__13409_ (
);

FILL FILL_2__7190_ (
);

FILL FILL_0__9829_ (
);

FILL FILL_0__9409_ (
);

FILL FILL_3__7506_ (
);

INVX1 _6650_ (
    .A(_248_),
    .Y(_249_)
);

FILL FILL_1__11790_ (
);

FILL FILL_3__10336_ (
);

FILL FILL_1__11370_ (
);

FILL FILL_2__8395_ (
);

FILL FILL_0__10783_ (
);

FILL FILL_0__10363_ (
);

NAND3X1 _7855_ (
    .A(_1361_),
    .B(_1368_),
    .C(_1367_),
    .Y(_1369_)
);

AND2X2 _7435_ (
    .A(vdd),
    .B(\X[1] [4]),
    .Y(_955_)
);

NAND2X1 _7015_ (
    .A(_606_),
    .B(_607_),
    .Y(_608_)
);

FILL FILL_1__6392_ (
);

FILL FILL_2__13162_ (
);

FILL FILL_2__6708_ (
);

FILL FILL_1__12995_ (
);

FILL FILL_1__12575_ (
);

FILL FILL_1__12155_ (
);

FILL FILL_0__11988_ (
);

FILL FILL_0__9582_ (
);

FILL FILL_0__9162_ (
);

NAND3X1 _11853_ (
    .A(_4966_),
    .B(_4959_),
    .C(_4964_),
    .Y(_4973_)
);

FILL FILL_0__11568_ (
);

NAND2X1 _11433_ (
    .A(_4616_),
    .B(_4621_),
    .Y(_4622_)
);

FILL FILL_0__11148_ (
);

AND2X2 _11013_ (
    .A(\X[5] [3]),
    .B(vdd),
    .Y(_4212_)
);

FILL FILL_1__7597_ (
);

FILL FILL_1__7177_ (
);

FILL FILL_3__8884_ (
);

OAI21X1 _12638_ (
    .A(_5677_),
    .B(_5678_),
    .C(_5676_),
    .Y(_5679_)
);

NAND3X1 _12218_ (
    .A(_5324_),
    .B(_5328_),
    .C(_5332_),
    .Y(_5333_)
);

FILL FILL_2__6881_ (
);

FILL FILL_2__6461_ (
);

FILL FILL_3__11294_ (
);

FILL FILL_2__10287_ (
);

FILL FILL_1__9743_ (
);

FILL FILL_1__9323_ (
);

FILL FILL_3__9669_ (
);

NAND2X1 _8393_ (
    .A(_1826_),
    .B(_1831_),
    .Y(_1832_)
);

FILL FILL_1__10641_ (
);

FILL FILL_1__10221_ (
);

CLKBUF1 CLKBUF1_insert20 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert21 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert22 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert23 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert24 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf45)
);

FILL FILL_2__7666_ (
);

CLKBUF1 CLKBUF1_insert25 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf44)
);

FILL FILL_3__12079_ (
);

CLKBUF1 CLKBUF1_insert26 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert27 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert28 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert29 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf40)
);

NOR2X1 _12391_ (
    .A(\u_fir_pe6.rYin [9]),
    .B(\u_fir_pe6.mul [9]),
    .Y(_5495_)
);

NAND2X1 _6706_ (
    .A(Xin[1]),
    .B(gnd),
    .Y(_304_)
);

FILL FILL_2__12853_ (
);

FILL FILL_2__12433_ (
);

FILL FILL_2__12013_ (
);

OAI21X1 _9598_ (
    .A(_2696_),
    .B(_2870_),
    .C(_2914_),
    .Y(_2952_)
);

NAND3X1 _9178_ (
    .A(_2537_),
    .B(_2531_),
    .C(_2534_),
    .Y(_2538_)
);

FILL FILL_1__11846_ (
);

FILL FILL_1__11426_ (
);

FILL FILL_1__11006_ (
);

FILL FILL_0__8853_ (
);

FILL FILL_3__6950_ (
);

FILL FILL_0__8433_ (
);

FILL FILL_0__10839_ (
);

FILL FILL_3__6530_ (
);

FILL FILL_0__10419_ (
);

NOR2X1 _10704_ (
    .A(_3965_),
    .B(_3908_),
    .Y(_3980_[1])
);

FILL FILL_0__8013_ (
);

NAND2X1 _13176_ (
    .A(_6207_),
    .B(_6201_),
    .Y(_6375_[14])
);

FILL FILL_2__9812_ (
);

FILL FILL_1__6868_ (
);

FILL FILL_1__6448_ (
);

FILL FILL_2__13218_ (
);

FILL FILL_0__9638_ (
);

FILL FILL_3__7735_ (
);

FILL FILL_0__9218_ (
);

INVX1 _11909_ (
    .A(_5022_),
    .Y(_5028_)
);

FILL FILL_3__7315_ (
);

FILL FILL_3__10565_ (
);

FILL FILL_0__10592_ (
);

FILL FILL_0__10172_ (
);

AOI21X1 _7664_ (
    .A(_1146_),
    .B(_1147_),
    .C(_1114_),
    .Y(_1181_)
);

DFFPOSX1 _7244_ (
    .D(_796_[5]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.mul [5])
);

FILL FILL_2__6937_ (
);

FILL FILL_2__6517_ (
);

FILL FILL_1__12384_ (
);

FILL FILL_0__9391_ (
);

FILL FILL_0__11797_ (
);

OR2X2 _11662_ (
    .A(_5513_),
    .B(_4784_),
    .Y(_4785_)
);

FILL FILL_0__11377_ (
);

NAND2X1 _11242_ (
    .A(_4427_),
    .B(_4434_),
    .Y(_4438_)
);

FILL FILL_3__12711_ (
);

FILL FILL_2__11704_ (
);

AND2X2 _8869_ (
    .A(_2271_),
    .B(_2281_),
    .Y(_2292_)
);

OAI21X1 _8449_ (
    .A(_1886_),
    .B(_1887_),
    .C(_1885_),
    .Y(_1888_)
);

NOR2X1 _8029_ (
    .A(_1532_),
    .B(_1529_),
    .Y(_1533_)
);

FILL FILL_0__7704_ (
);

NOR2X1 _9810_ (
    .A(\u_fir_pe3.rYin [14]),
    .B(\u_fir_pe3.mul [14]),
    .Y(_3154_)
);

FILL FILL_1__13169_ (
);

NAND3X1 _12867_ (
    .A(vdd),
    .B(\X[6] [6]),
    .C(_5904_),
    .Y(_5905_)
);

FILL FILL_3__8273_ (
);

NAND2X1 _12447_ (
    .A(_5546_),
    .B(_5540_),
    .Y(_5550_)
);

AOI21X1 _12027_ (
    .A(_5139_),
    .B(_5144_),
    .C(_5083_),
    .Y(_5145_)
);

FILL FILL_2__12909_ (
);

FILL FILL_0__13103_ (
);

FILL FILL254250x212550 (
);

FILL FILL_2__6690_ (
);

FILL FILL_0__8909_ (
);

FILL FILL_2__10096_ (
);

FILL FILL_1__9972_ (
);

FILL FILL_1__9552_ (
);

FILL FILL_1__9132_ (
);

FILL FILL_3__9898_ (
);

FILL FILL_3__9478_ (
);

FILL FILL_3__9058_ (
);

FILL FILL_1__10870_ (
);

FILL FILL_1__10450_ (
);

FILL FILL_1__10030_ (
);

FILL FILL_2__7895_ (
);

FILL FILL_2__7475_ (
);

FILL FILL_2__7055_ (
);

INVX1 _6935_ (
    .A(_529_),
    .Y(_530_)
);

NAND3X1 _6515_ (
    .A(_53_),
    .B(_111_),
    .C(_115_),
    .Y(_116_)
);

FILL FILL_2__12662_ (
);

FILL FILL_2__12242_ (
);

FILL FILL_1__11655_ (
);

FILL FILL_1__11235_ (
);

FILL FILL_0__8662_ (
);

FILL FILL_0__8242_ (
);

FILL FILL_0__10648_ (
);

NAND3X1 _10933_ (
    .A(vdd),
    .B(\X[5] [6]),
    .C(_4130_),
    .Y(_4133_)
);

NAND2X1 _10513_ (
    .A(_3785_),
    .B(_3784_),
    .Y(_3786_)
);

FILL FILL_0__10228_ (
);

FILL FILL_2__9621_ (
);

FILL FILL_2__9201_ (
);

FILL FILL_1__6677_ (
);

FILL FILL_2__13027_ (
);

FILL FILL_3__7964_ (
);

FILL FILL_0__9447_ (
);

FILL FILL_0__9027_ (
);

NAND2X1 _11718_ (
    .A(_4836_),
    .B(_4839_),
    .Y(_4840_)
);

FILL FILL_3__7124_ (
);

FILL FILL_3__10794_ (
);

FILL FILL_1__8823_ (
);

FILL FILL_1__8403_ (
);

FILL FILL_3__8749_ (
);

NAND2X1 _7893_ (
    .A(_1402_),
    .B(_1405_),
    .Y(_1406_)
);

NAND3X1 _7473_ (
    .A(_987_),
    .B(_988_),
    .C(_989_),
    .Y(_993_)
);

AND2X2 _7053_ (
    .A(\u_fir_pe0.rYin [2]),
    .B(\u_fir_pe0.mul [2]),
    .Y(_641_)
);

FILL FILL_2__6746_ (
);

FILL FILL_3__11579_ (
);

FILL FILL_1__12193_ (
);

AND2X2 _11891_ (
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5010_)
);

OR2X2 _11471_ (
    .A(_4649_),
    .B(_4654_),
    .Y(_4656_)
);

FILL FILL_0__11186_ (
);

AOI21X1 _11051_ (
    .A(_4137_),
    .B(_4156_),
    .C(_4249_),
    .Y(_4250_)
);

FILL FILL_3__12940_ (
);

FILL FILL_1__9608_ (
);

FILL FILL_3__12100_ (
);

FILL FILL_2__11933_ (
);

FILL FILL_2__11513_ (
);

OAI22X1 _8678_ (
    .A(_2011_),
    .B(_2056_),
    .C(_2112_),
    .D(_2111_),
    .Y(_2113_)
);

NAND3X1 _8258_ (
    .A(_1696_),
    .B(_1698_),
    .C(_1697_),
    .Y(_1699_)
);

FILL FILL_1__10926_ (
);

FILL FILL_1__10506_ (
);

FILL FILL_0__7933_ (
);

FILL FILL_0__7513_ (
);

FILL FILL_1__13398_ (
);

AOI21X1 _12676_ (
    .A(_5670_),
    .B(_5674_),
    .C(_5663_),
    .Y(_5716_)
);

OAI21X1 _12256_ (
    .A(_5158_),
    .B(_5369_),
    .C(_5341_),
    .Y(_5370_)
);

FILL FILL_3__13305_ (
);

FILL FILL_2__12718_ (
);

FILL FILL_0__13332_ (
);

FILL FILL_0__8718_ (
);

FILL FILL_1__9781_ (
);

FILL FILL_1__9361_ (
);

FILL FILL_3__9287_ (
);

FILL FILL_2__7284_ (
);

INVX1 _6744_ (
    .A(_322_),
    .Y(_342_)
);

FILL FILL_2__12891_ (
);

FILL FILL_2__12051_ (
);

FILL FILL_1__11884_ (
);

FILL FILL_1__11464_ (
);

FILL FILL_1__11044_ (
);

FILL FILL_0__8891_ (
);

FILL FILL_2__8489_ (
);

FILL FILL_0__8471_ (
);

FILL FILL_0__10877_ (
);

FILL FILL_0__10457_ (
);

DFFPOSX1 _10742_ (
    .D(\Y[4] [11]),
    .CLK(clk_bF$buf44),
    .Q(\u_fir_pe4.rYin [11])
);

FILL FILL_2__8069_ (
);

FILL FILL_0__8051_ (
);

NAND2X1 _10322_ (
    .A(_3589_),
    .B(_3598_),
    .Y(_3599_)
);

FILL FILL_0__10037_ (
);

FILL FILL_2__9430_ (
);

FILL FILL_2__9010_ (
);

NOR2X1 _7949_ (
    .A(\u_fir_pe1.rYin [4]),
    .B(\u_fir_pe1.mul [4]),
    .Y(_1455_)
);

OAI21X1 _7529_ (
    .A(_1047_),
    .B(_1042_),
    .C(_1036_),
    .Y(_1048_)
);

NOR2X1 _7109_ (
    .A(_690_),
    .B(_691_),
    .Y(_692_)
);

FILL FILL_1__6486_ (
);

FILL FILL_2__13256_ (
);

FILL FILL_1__12669_ (
);

FILL FILL_1__12249_ (
);

FILL FILL_0__9676_ (
);

FILL FILL_0__9256_ (
);

AOI21X1 _11947_ (
    .A(_5065_),
    .B(_5064_),
    .C(_5063_),
    .Y(_5066_)
);

FILL FILL_3__7353_ (
);

NOR2X1 _11527_ (
    .A(_4709_),
    .B(_4710_),
    .Y(_4711_)
);

OAI21X1 _11107_ (
    .A(_4000_),
    .B(_4304_),
    .C(_4010_),
    .Y(_4305_)
);

FILL FILL_0__12603_ (
);

FILL FILL_3__10183_ (
);

FILL FILL_1__8632_ (
);

FILL FILL_1__8212_ (
);

FILL FILL_3__8138_ (
);

OAI21X1 _7282_ (
    .A(_801_),
    .B(_804_),
    .C(_797_),
    .Y(_805_)
);

FILL FILL_2__6975_ (
);

FILL FILL_2__6555_ (
);

NAND3X1 _11280_ (
    .A(_4473_),
    .B(_4475_),
    .C(_4474_),
    .Y(_4476_)
);

FILL FILL_1__9417_ (
);

FILL FILL_2__11742_ (
);

FILL FILL_2__11322_ (
);

AND2X2 _8487_ (
    .A(gnd),
    .B(\X[2] [6]),
    .Y(_1925_)
);

NAND3X1 _8067_ (
    .A(_1564_),
    .B(_1570_),
    .C(_1565_),
    .Y(_1571_)
);

FILL FILL_1__10315_ (
);

FILL FILL_0__7742_ (
);

FILL FILL_0__7322_ (
);

DFFPOSX1 _12485_ (
    .D(\Y[7] [0]),
    .CLK(clk_bF$buf49),
    .Q(\u_fir_pe6.rYin [0])
);

NOR2X1 _12065_ (
    .A(_5180_),
    .B(_5181_),
    .Y(_5182_)
);

FILL FILL_2__8701_ (
);

FILL FILL_2__12947_ (
);

FILL FILL_2__12527_ (
);

FILL FILL_2__12107_ (
);

FILL FILL_0__13141_ (
);

FILL FILL_0__8947_ (
);

FILL FILL_0__8527_ (
);

FILL FILL_3__6624_ (
);

FILL FILL_1__9590_ (
);

FILL FILL_1__9170_ (
);

FILL FILL_2__9906_ (
);

FILL FILL_2__7093_ (
);

FILL FILL_1__7903_ (
);

FILL FILL_3__7829_ (
);

FILL FILL_3__7409_ (
);

NOR2X1 _6973_ (
    .A(_144_),
    .B(_305_),
    .Y(_567_)
);

NAND2X1 _6553_ (
    .A(gnd),
    .B(Xin[3]),
    .Y(_153_)
);

FILL FILL_2__12280_ (
);

FILL FILL_3__10659_ (
);

FILL FILL_1__11693_ (
);

FILL FILL_1__11273_ (
);

FILL FILL_2__8298_ (
);

FILL FILL_0__8280_ (
);

FILL FILL_0__10686_ (
);

NAND3X1 _10971_ (
    .A(_4157_),
    .B(_4161_),
    .C(_4164_),
    .Y(_4171_)
);

INVX1 _10551_ (
    .A(\u_fir_pe4.rYin [1]),
    .Y(_3820_)
);

FILL FILL_0__10266_ (
);

NAND2X1 _10131_ (
    .A(_3406_),
    .B(_3409_),
    .Y(_3410_)
);

AND2X2 _7758_ (
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_1274_)
);

AOI21X1 _7338_ (
    .A(_837_),
    .B(_841_),
    .C(_829_),
    .Y(_860_)
);

FILL FILL_2__13065_ (
);

FILL FILL_1__12898_ (
);

FILL FILL_1__12058_ (
);

FILL FILL_0__9485_ (
);

FILL FILL_3__7582_ (
);

FILL FILL_0__9065_ (
);

NAND3X1 _11756_ (
    .A(_4867_),
    .B(_4874_),
    .C(_4876_),
    .Y(_4877_)
);

NAND3X1 _11336_ (
    .A(_4528_),
    .B(_4530_),
    .C(_4529_),
    .Y(_4531_)
);

FILL FILL_3__12805_ (
);

FILL FILL_0__12832_ (
);

FILL FILL_0__12412_ (
);

INVX1 _9904_ (
    .A(_3975_),
    .Y(_3976_)
);

FILL FILL_1__8861_ (
);

FILL FILL_1__8441_ (
);

FILL FILL_1__8021_ (
);

FILL FILL_3__8367_ (
);

NOR2X1 _7091_ (
    .A(_673_),
    .B(_674_),
    .Y(_675_)
);

FILL FILL_2__6784_ (
);

FILL FILL_3__11197_ (
);

FILL FILL_1__9646_ (
);

FILL FILL_1__9226_ (
);

FILL FILL_2__11971_ (
);

FILL FILL_2__11551_ (
);

FILL FILL_2__11131_ (
);

AND2X2 _8296_ (
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_1736_)
);

FILL FILL_1__10964_ (
);

FILL FILL_1__10544_ (
);

FILL FILL_1__10124_ (
);

FILL FILL_2__7989_ (
);

FILL FILL_0__7971_ (
);

FILL FILL_2__7569_ (
);

FILL FILL_0__7551_ (
);

FILL FILL_2__7149_ (
);

FILL FILL_0__7131_ (
);

NOR3X1 _12294_ (
    .A(_5405_),
    .B(_5373_),
    .C(_5391_),
    .Y(_5406_)
);

FILL FILL_2__8930_ (
);

FILL FILL_2__8510_ (
);

AOI21X1 _6609_ (
    .A(_172_),
    .B(_176_),
    .C(_138_),
    .Y(_208_)
);

FILL FILL_2__12756_ (
);

FILL FILL_2__12336_ (
);

FILL FILL_1__11749_ (
);

FILL FILL_1__11329_ (
);

FILL FILL_0__8756_ (
);

FILL FILL_3__6853_ (
);

FILL FILL_0__8336_ (
);

INVX1 _10607_ (
    .A(\u_fir_pe4.mul [7]),
    .Y(_3870_)
);

NAND3X1 _13079_ (
    .A(_6108_),
    .B(_6113_),
    .C(_6112_),
    .Y(_6114_)
);

FILL FILL_2__9715_ (
);

FILL FILL_1__7712_ (
);

FILL FILL_3__7638_ (
);

INVX1 _6782_ (
    .A(_372_),
    .Y(_379_)
);

FILL FILL_3__10048_ (
);

FILL FILL_1__11082_ (
);

FILL FILL_0__10495_ (
);

NAND2X1 _10780_ (
    .A(vdd),
    .B(\X[5] [3]),
    .Y(_4772_)
);

OAI21X1 _10360_ (
    .A(_3635_),
    .B(_3636_),
    .C(_3632_),
    .Y(_3637_)
);

FILL FILL_0__10075_ (
);

FILL FILL_1__8917_ (
);

FILL FILL_2__10822_ (
);

FILL FILL_2__10402_ (
);

NOR2X1 _7987_ (
    .A(\u_fir_pe1.rYin [8]),
    .B(\u_fir_pe1.mul [8]),
    .Y(_1490_)
);

AND2X2 _7567_ (
    .A(_1082_),
    .B(_1085_),
    .Y(_1086_)
);

AND2X2 _7147_ (
    .A(_729_),
    .B(_730_),
    .Y(_790_[10])
);

FILL FILL_2__13294_ (
);

FILL FILL_0__6822_ (
);

FILL FILL_0__6402_ (
);

FILL FILL_1__12287_ (
);

FILL FILL_0__9294_ (
);

NAND2X1 _11985_ (
    .A(\X[7] [4]),
    .B(gnd),
    .Y(_5103_)
);

NOR2X1 _11565_ (
    .A(_4748_),
    .B(_4747_),
    .Y(_4749_)
);

INVX1 _11145_ (
    .A(_4256_),
    .Y(_4343_)
);

FILL FILL_0__12641_ (
);

FILL FILL_0__12221_ (
);

FILL FILL_0__7607_ (
);

NOR2X1 _9713_ (
    .A(_3056_),
    .B(_3057_),
    .Y(_3058_)
);

FILL FILL_1__8670_ (
);

FILL FILL_1__8250_ (
);

FILL FILL_3__8596_ (
);

FILL FILL_0__13006_ (
);

FILL FILL_2__6593_ (
);

FILL FILL253650x93750 (
);

FILL FILL_1__9455_ (
);

FILL FILL_1__9035_ (
);

FILL FILL_2__11780_ (
);

FILL FILL_2__11360_ (
);

FILL FILL_1__10773_ (
);

FILL FILL_1__10353_ (
);

FILL FILL_2__7798_ (
);

FILL FILL_0__7780_ (
);

FILL FILL_2__7378_ (
);

FILL FILL_0__7360_ (
);

FILL FILL_3__13152_ (
);

AOI21X1 _6838_ (
    .A(_425_),
    .B(_423_),
    .C(_395_),
    .Y(_435_)
);

NAND3X1 _6418_ (
    .A(_20_),
    .B(_786_),
    .C(_19_),
    .Y(_21_)
);

FILL FILL_2__12985_ (
);

FILL FILL_2__12565_ (
);

FILL FILL_2__12145_ (
);

FILL FILL_1__11978_ (
);

FILL FILL_1__11558_ (
);

FILL FILL_1__11138_ (
);

FILL FILL_0__8565_ (
);

FILL FILL_0__8145_ (
);

AOI22X1 _10836_ (
    .A(_3994_),
    .B(_3999_),
    .C(_4034_),
    .D(_4037_),
    .Y(_4038_)
);

AOI21X1 _10416_ (
    .A(_3619_),
    .B(_3625_),
    .C(_3691_),
    .Y(_3692_)
);

FILL FILL_2__9944_ (
);

FILL FILL_0__11912_ (
);

FILL FILL_2__9524_ (
);

FILL FILL_2__9104_ (
);

FILL FILL_1__7941_ (
);

FILL FILL_1__7521_ (
);

FILL FILL_1__7101_ (
);

FILL FILL_3__7447_ (
);

NAND3X1 _6591_ (
    .A(_184_),
    .B(_177_),
    .C(_182_),
    .Y(_191_)
);

FILL FILL_3__10277_ (
);

FILL FILL_1__8726_ (
);

FILL FILL_1__8306_ (
);

FILL FILL_2__10631_ (
);

FILL FILL_2__10211_ (
);

AOI21X1 _7796_ (
    .A(_1257_),
    .B(_1291_),
    .C(_1310_),
    .Y(_1311_)
);

OAI21X1 _7376_ (
    .A(_895_),
    .B(_896_),
    .C(_894_),
    .Y(_897_)
);

FILL FILL_0__6631_ (
);

FILL FILL_2__6649_ (
);

FILL FILL_1__12096_ (
);

NAND2X1 _11794_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf2 ),
    .Y(_4914_)
);

FILL FILL_0__11089_ (
);

OR2X2 _11374_ (
    .A(_4566_),
    .B(_4564_),
    .Y(_4568_)
);

FILL FILL_3__12423_ (
);

FILL FILL_2__11836_ (
);

FILL FILL_0__12870_ (
);

FILL FILL_2__11416_ (
);

FILL FILL_0__12450_ (
);

FILL FILL_0__12030_ (
);

FILL FILL_1__10829_ (
);

FILL FILL_1__10409_ (
);

FILL FILL_0__7836_ (
);

AND2X2 _9942_ (
    .A(gnd),
    .B(\X[4] [2]),
    .Y(_3224_)
);

FILL FILL_0__7416_ (
);

NAND3X1 _9522_ (
    .A(_2861_),
    .B(_2877_),
    .C(_2875_),
    .Y(_2878_)
);

AND2X2 _9102_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf1 ),
    .Y(_2463_)
);

AOI21X1 _12999_ (
    .A(_6020_),
    .B(_6016_),
    .C(_5961_),
    .Y(_6035_)
);

NAND2X1 _12579_ (
    .A(vdd),
    .B(\X[6] [2]),
    .Y(_5621_)
);

NAND2X1 _12159_ (
    .A(_5273_),
    .B(_5269_),
    .Y(_5275_)
);

FILL FILL_0__13235_ (
);

NAND2X1 _13100_ (
    .A(_6133_),
    .B(_6134_),
    .Y(_6375_[11])
);

FILL FILL_3__6718_ (
);

FILL FILL_1__9684_ (
);

FILL FILL_1__9264_ (
);

FILL FILL_1__10582_ (
);

FILL FILL_1__10162_ (
);

FILL FILL_2__7187_ (
);

INVX1 _6647_ (
    .A(_240_),
    .Y(_246_)
);

FILL FILL_2__12794_ (
);

FILL FILL_2__12374_ (
);

FILL FILL_1__11787_ (
);

FILL FILL_1__11367_ (
);

FILL FILL_0__8794_ (
);

FILL FILL_3__6891_ (
);

FILL FILL_0__8374_ (
);

FILL FILL_3__6471_ (
);

INVX1 _10645_ (
    .A(_3907_),
    .Y(_3909_)
);

NAND2X1 _10225_ (
    .A(_3498_),
    .B(_3502_),
    .Y(_3503_)
);

FILL FILL_2__9753_ (
);

FILL FILL_2__9333_ (
);

FILL FILL_0__11721_ (
);

FILL FILL_0__11301_ (
);

FILL FILL_1__6389_ (
);

FILL FILL_2__13159_ (
);

FILL FILL_1__7750_ (
);

FILL FILL_1__7330_ (
);

FILL FILL_0__9999_ (
);

FILL FILL_0__9579_ (
);

FILL FILL_3__7676_ (
);

FILL FILL_0__9159_ (
);

FILL FILL_3__7256_ (
);

FILL FILL_0__12926_ (
);

FILL FILL_1__8535_ (
);

FILL FILL_2__10860_ (
);

FILL FILL_2__10440_ (
);

FILL FILL_2__10020_ (
);

NAND2X1 _7185_ (
    .A(_764_),
    .B(_758_),
    .Y(_768_)
);

FILL FILL_3__9822_ (
);

FILL FILL_2__6878_ (
);

FILL FILL_0__6860_ (
);

FILL FILL_0__6440_ (
);

FILL FILL_2__6458_ (
);

AND2X2 _11183_ (
    .A(_4379_),
    .B(_4376_),
    .Y(_4380_)
);

FILL FILL_3__12652_ (
);

FILL FILL_3__12232_ (
);

FILL FILL_2__11645_ (
);

FILL FILL_2__11225_ (
);

FILL FILL_1__10638_ (
);

FILL FILL_1__10218_ (
);

FILL FILL_0__7645_ (
);

OAI21X1 _9751_ (
    .A(_3083_),
    .B(_3084_),
    .C(_3094_),
    .Y(_3095_)
);

INVX1 _9331_ (
    .A(_2673_),
    .Y(_2689_)
);

INVX1 _12388_ (
    .A(_5487_),
    .Y(_5491_)
);

FILL FILL_2__8604_ (
);

FILL FILL_3__13017_ (
);

FILL FILL_0__13044_ (
);

FILL FILL_1__6601_ (
);

FILL FILL_3__6947_ (
);

FILL FILL_1__9493_ (
);

FILL FILL_1__9073_ (
);

FILL FILL_2__9809_ (
);

FILL FILL_1__10391_ (
);

FILL FILL_1__7806_ (
);

OAI21X1 _6876_ (
    .A(_419_),
    .B(_471_),
    .C(_407_),
    .Y(_472_)
);

NAND2X1 _6456_ (
    .A(_54_),
    .B(_57_),
    .Y(_58_)
);

FILL FILL_2__12183_ (
);

FILL FILL_1__11176_ (
);

FILL FILL_0__8183_ (
);

FILL FILL_0__10589_ (
);

OAI21X1 _10874_ (
    .A(_4074_),
    .B(_4000_),
    .C(_4068_),
    .Y(_4075_)
);

NAND2X1 _10454_ (
    .A(_3728_),
    .B(_3727_),
    .Y(_3729_)
);

FILL FILL_0__10169_ (
);

INVX1 _10034_ (
    .A(_3255_),
    .Y(_3315_)
);

FILL FILL_3__11503_ (
);

FILL FILL_2__9982_ (
);

FILL FILL_2__10916_ (
);

FILL FILL_2__9562_ (
);

FILL FILL_0__11950_ (
);

FILL FILL_2__9142_ (
);

FILL FILL_0__11530_ (
);

FILL FILL_0__11110_ (
);

FILL FILL_0__6916_ (
);

OAI21X1 _8602_ (
    .A(_2029_),
    .B(_2028_),
    .C(_1979_),
    .Y(_2039_)
);

FILL FILL_0__9388_ (
);

NAND2X1 _11659_ (
    .A(gnd),
    .B(\X[7] [2]),
    .Y(_4782_)
);

FILL FILL_3__7065_ (
);

OR2X2 _11239_ (
    .A(_4365_),
    .B(_4435_),
    .Y(_4436_)
);

FILL FILL_1__13322_ (
);

FILL FILL_0__12735_ (
);

AOI21X1 _12600_ (
    .A(_5619_),
    .B(_5623_),
    .C(_5611_),
    .Y(_5642_)
);

FILL FILL_0__12315_ (
);

INVX1 _9807_ (
    .A(\u_fir_pe3.rYin [14]),
    .Y(_3150_)
);

FILL FILL_1__8764_ (
);

FILL FILL_1__8344_ (
);

FILL FILL_3__9211_ (
);

FILL FILL_2__6687_ (
);

FILL FILL_1__9969_ (
);

FILL FILL_3__12881_ (
);

FILL FILL_1__9549_ (
);

FILL FILL_1__9129_ (
);

FILL FILL_3__12041_ (
);

FILL FILL_2__11874_ (
);

FILL FILL_2__11454_ (
);

FILL FILL_2__11034_ (
);

NAND2X1 _8199_ (
    .A(_1638_),
    .B(_1634_),
    .Y(_1641_)
);

FILL FILL_1__10867_ (
);

FILL FILL_1__10447_ (
);

FILL FILL_1__10027_ (
);

FILL FILL_0__7874_ (
);

NAND2X1 _9980_ (
    .A(_3888_),
    .B(_3260_),
    .Y(_3261_)
);

FILL FILL_0__7454_ (
);

NAND2X1 _9560_ (
    .A(_2910_),
    .B(_2914_),
    .Y(_2915_)
);

FILL FILL_0__7034_ (
);

OAI21X1 _9140_ (
    .A(_2499_),
    .B(_2500_),
    .C(_2498_),
    .Y(_2501_)
);

INVX1 _12197_ (
    .A(_5311_),
    .Y(_5312_)
);

FILL FILL_2__8833_ (
);

FILL FILL_2__8413_ (
);

FILL FILL_0__10801_ (
);

FILL FILL_3__13246_ (
);

FILL FILL_2__12659_ (
);

FILL FILL_2__12239_ (
);

FILL FILL_0__13273_ (
);

FILL FILL_1__6830_ (
);

FILL FILL_1__6410_ (
);

FILL FILL_0__8659_ (
);

FILL FILL_0__8239_ (
);

FILL FILL_0__9600_ (
);

FILL FILL_2__9618_ (
);

FILL FILL_1__7615_ (
);

AOI21X1 _6685_ (
    .A(_283_),
    .B(_282_),
    .C(_281_),
    .Y(_284_)
);

FILL FILL_3__8902_ (
);

FILL FILL_0__10398_ (
);

OAI21X1 _10683_ (
    .A(_3939_),
    .B(_3940_),
    .C(_3944_),
    .Y(_3946_)
);

AND2X2 _10263_ (
    .A(_3502_),
    .B(_3498_),
    .Y(_3541_)
);

FILL FILL_3__11732_ (
);

FILL FILL_2__9791_ (
);

FILL FILL_2__9371_ (
);

FILL FILL_2__10305_ (
);

FILL FILL_2__13197_ (
);

FILL FILL_0__6725_ (
);

OR2X2 _8831_ (
    .A(_2255_),
    .B(_2253_),
    .Y(_2257_)
);

OAI21X1 _8411_ (
    .A(_1842_),
    .B(_1849_),
    .C(_1834_),
    .Y(_1850_)
);

FILL FILL_0__9197_ (
);

NAND2X1 _11888_ (
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_5007_)
);

FILL FILL_3__7294_ (
);

NOR2X1 _11468_ (
    .A(\u_fir_pe5.rYin [5]),
    .B(\u_fir_pe5.mul [5]),
    .Y(_4653_)
);

AOI21X1 _11048_ (
    .A(_4246_),
    .B(_4245_),
    .C(_4244_),
    .Y(_4247_)
);

FILL FILL_3__12517_ (
);

FILL FILL_1__13131_ (
);

FILL FILL_0__12964_ (
);

FILL FILL_0__12544_ (
);

FILL FILL_0__12124_ (
);

AOI21X1 _9616_ (
    .A(_2968_),
    .B(_2969_),
    .C(_2952_),
    .Y(_2970_)
);

FILL FILL_1__8573_ (
);

FILL FILL_1__8153_ (
);

FILL FILL_3__9440_ (
);

FILL FILL_0__13329_ (
);

FILL FILL_2__6496_ (
);

FILL FILL_1__9778_ (
);

FILL FILL_1__9358_ (
);

FILL FILL_2__11683_ (
);

FILL FILL_2__11263_ (
);

FILL FILL_1__10676_ (
);

FILL FILL_1__10256_ (
);

FILL FILL_0__7683_ (
);

FILL FILL_0__7263_ (
);

FILL FILL_2__8642_ (
);

FILL FILL_2__8222_ (
);

FILL FILL_0__10610_ (
);

FILL FILL_2__12888_ (
);

FILL FILL_2__12048_ (
);

FILL FILL_0__13082_ (
);

FILL FILL_0__8888_ (
);

FILL FILL_3__6985_ (
);

FILL FILL_0__8468_ (
);

FILL FILL_3__6565_ (
);

DFFPOSX1 _10739_ (
    .D(\Y[4] [8]),
    .CLK(clk_bF$buf55),
    .Q(\u_fir_pe4.rYin [8])
);

FILL FILL_0__8048_ (
);

AND2X2 _10319_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3596_)
);

FILL FILL_1__12822_ (
);

FILL FILL_1__12402_ (
);

FILL FILL_2__9427_ (
);

FILL FILL_0__11815_ (
);

FILL FILL_3_CLKBUF1_insert91 (
);

FILL FILL_3_CLKBUF1_insert93 (
);

FILL FILL_3_CLKBUF1_insert95 (
);

FILL FILL_3_CLKBUF1_insert96 (
);

FILL FILL_1__7844_ (
);

FILL FILL_1__7424_ (
);

FILL FILL_1__7004_ (
);

NAND3X1 _6494_ (
    .A(_85_),
    .B(_92_),
    .C(_94_),
    .Y(_95_)
);

NAND3X1 _10492_ (
    .A(_3750_),
    .B(_3760_),
    .C(_3763_),
    .Y(_3766_)
);

NAND2X1 _10072_ (
    .A(gnd),
    .B(\X[4] [4]),
    .Y(_3352_)
);

FILL FILL_1__8629_ (
);

FILL FILL_3__11961_ (
);

FILL FILL_1__8209_ (
);

FILL FILL_3__11121_ (
);

FILL FILL_2__10954_ (
);

FILL FILL_2__10534_ (
);

FILL FILL_2__9180_ (
);

FILL FILL_2__10114_ (
);

OAI21X1 _7699_ (
    .A(_822_),
    .B(_1213_),
    .C(_1215_),
    .Y(_1216_)
);

INVX1 _7279_ (
    .A(_801_),
    .Y(_802_)
);

FILL FILL_3__9916_ (
);

FILL FILL_0__6954_ (
);

FILL FILL_0__6534_ (
);

NAND3X1 _8640_ (
    .A(_2074_),
    .B(_2075_),
    .C(_2073_),
    .Y(_2076_)
);

NOR2X1 _8220_ (
    .A(_1615_),
    .B(_1652_),
    .Y(_1661_)
);

NAND2X1 _11697_ (
    .A(_4817_),
    .B(_4818_),
    .Y(_4819_)
);

NAND2X1 _11277_ (
    .A(_4454_),
    .B(_4451_),
    .Y(_4473_)
);

FILL FILL_2__7913_ (
);

FILL FILL_3__12746_ (
);

FILL FILL_2__11739_ (
);

FILL FILL_0__12773_ (
);

FILL FILL_2__11319_ (
);

FILL FILL_0__12353_ (
);

FILL FILL_0__7739_ (
);

DFFPOSX1 _9845_ (
    .D(_3181_[15]),
    .CLK(clk_bF$buf26),
    .Q(\Y[4] [15])
);

FILL FILL_0__7319_ (
);

OAI21X1 _9425_ (
    .A(_2781_),
    .B(_2780_),
    .C(_2777_),
    .Y(_2782_)
);

DFFPOSX1 _9005_ (
    .D(_2390_[12]),
    .CLK(clk_bF$buf15),
    .Q(\u_fir_pe2.mul [12])
);

FILL FILL_1__8382_ (
);

FILL FILL_0__13138_ (
);

OAI21X1 _13003_ (
    .A(_5965_),
    .B(_5969_),
    .C(_5967_),
    .Y(_6039_)
);

FILL FILL_1__9587_ (
);

FILL FILL_1__9167_ (
);

FILL FILL_2__11492_ (
);

FILL FILL_2__11072_ (
);

FILL FILL_1__10485_ (
);

FILL FILL_1__10065_ (
);

FILL FILL253650x25350 (
);

FILL FILL_0__7492_ (
);

FILL FILL_0__7072_ (
);

FILL FILL_2__8871_ (
);

FILL FILL_2__8451_ (
);

FILL FILL_2__8031_ (
);

FILL FILL_2__12697_ (
);

FILL FILL_2__12277_ (
);

INVX1 _7911_ (
    .A(_1413_),
    .Y(_1423_)
);

FILL FILL_0__8697_ (
);

FILL FILL_3__6794_ (
);

FILL FILL_0__8277_ (
);

NAND3X1 _10968_ (
    .A(_4121_),
    .B(_4162_),
    .C(_4167_),
    .Y(_4168_)
);

NAND2X1 _10548_ (
    .A(_3818_),
    .B(_3817_),
    .Y(_3984_[15])
);

AOI21X1 _10128_ (
    .A(_3335_),
    .B(_3331_),
    .C(_3400_),
    .Y(_3407_)
);

FILL FILL_1__12631_ (
);

FILL FILL_1__12211_ (
);

FILL FILL_2__9656_ (
);

FILL FILL_2__9236_ (
);

FILL FILL_0__11204_ (
);

FILL FILL254550x176550 (
);

FILL FILL_1__7653_ (
);

FILL FILL_3__7999_ (
);

FILL FILL_3__7159_ (
);

FILL FILL_1__13416_ (
);

FILL FILL_0__12829_ (
);

FILL FILL_3__8520_ (
);

FILL FILL_0__12409_ (
);

FILL FILL_1__8858_ (
);

FILL FILL_1__8438_ (
);

FILL FILL_1__8018_ (
);

FILL FILL_3__11350_ (
);

FILL FILL_2__10763_ (
);

FILL FILL_2__10343_ (
);

OAI21X1 _7088_ (
    .A(_665_),
    .B(_666_),
    .C(_670_),
    .Y(_672_)
);

FILL FILL_3__9305_ (
);

FILL FILL_0__6763_ (
);

AOI21X1 _11086_ (
    .A(_4266_),
    .B(_4268_),
    .C(_4283_),
    .Y(_4284_)
);

FILL FILL_3__12975_ (
);

FILL FILL_2__7722_ (
);

FILL FILL_2__7302_ (
);

FILL FILL_3__12135_ (
);

FILL FILL_2__11968_ (
);

FILL FILL_2__11548_ (
);

FILL FILL_0__12582_ (
);

FILL FILL_2__11128_ (
);

FILL FILL_0__12162_ (
);

FILL FILL_0__7968_ (
);

FILL FILL_0__7548_ (
);

AOI21X1 _9654_ (
    .A(_2948_),
    .B(_2950_),
    .C(_3005_),
    .Y(_3006_)
);

FILL FILL_0__7128_ (
);

NAND2X1 _9234_ (
    .A(_2593_),
    .B(_2585_),
    .Y(_2594_)
);

FILL FILL_1__8191_ (
);

FILL FILL_1__11902_ (
);

FILL FILL_2__8927_ (
);

FILL FILL_2__8507_ (
);

NOR2X1 _13232_ (
    .A(_6255_),
    .B(_6254_),
    .Y(_6256_)
);

FILL FILL_1__6924_ (
);

FILL FILL_1__6504_ (
);

FILL FILL_1__9396_ (
);

FILL FILL_1__10294_ (
);

FILL FILL_1__7709_ (
);

FILL FILL_3__10201_ (
);

FILL FILL_2__8680_ (
);

FILL FILL_2__8260_ (
);

FILL FILL_3__13093_ (
);

AND2X2 _6779_ (
    .A(_367_),
    .B(_372_),
    .Y(_377_)
);

FILL FILL_2__12086_ (
);

AOI21X1 _7720_ (
    .A(_1227_),
    .B(_1223_),
    .C(_1182_),
    .Y(_1237_)
);

FILL FILL_1__11499_ (
);

NAND2X1 _7300_ (
    .A(\X[1] [4]),
    .B(gnd),
    .Y(_822_)
);

FILL FILL_1__11079_ (
);

NOR2X1 _10777_ (
    .A(_4768_),
    .B(_4767_),
    .Y(_4769_)
);

NAND3X1 _10357_ (
    .A(_3614_),
    .B(_3618_),
    .C(_3621_),
    .Y(_3634_)
);

FILL FILL_1__12860_ (
);

FILL FILL_1__12440_ (
);

FILL FILL_1__12020_ (
);

FILL FILL_2__10819_ (
);

FILL FILL_2__9465_ (
);

FILL FILL_0__11853_ (
);

FILL FILL_2__9045_ (
);

FILL FILL_0__11433_ (
);

FILL FILL_0__11013_ (
);

FILL FILL_0__6819_ (
);

NOR2X1 _8925_ (
    .A(_2348_),
    .B(_2347_),
    .Y(_2349_)
);

NAND3X1 _8505_ (
    .A(_1936_),
    .B(_1937_),
    .C(_1938_),
    .Y(_1943_)
);

FILL FILL_1__7882_ (
);

FILL FILL_1__7462_ (
);

FILL FILL_1__7042_ (
);

FILL FILL_3__7388_ (
);

FILL FILL_1__13225_ (
);

AOI21X1 _12923_ (
    .A(_5940_),
    .B(_5939_),
    .C(_5882_),
    .Y(_5960_)
);

FILL FILL_0__12638_ (
);

FILL FILL_0__12218_ (
);

DFFPOSX1 _12503_ (
    .D(_5575_[2]),
    .CLK(clk_bF$buf49),
    .Q(\u_fir_pe6.mul [2])
);

FILL FILL_1__8667_ (
);

FILL FILL_1__8247_ (
);

FILL FILL_2__10992_ (
);

FILL FILL_2__10572_ (
);

FILL FILL_2__10152_ (
);

FILL FILL_3__9534_ (
);

FILL FILL_0__6992_ (
);

FILL FILL_0__6572_ (
);

FILL FILL_2__7951_ (
);

FILL FILL_2__7531_ (
);

FILL FILL_2__7111_ (
);

FILL FILL_2__11777_ (
);

FILL FILL_2__11357_ (
);

FILL FILL_0__12391_ (
);

FILL FILL_0__7777_ (
);

DFFPOSX1 _9883_ (
    .D(_3187_[13]),
    .CLK(clk_bF$buf36),
    .Q(\u_fir_pe3.mul [13])
);

FILL FILL_0__7357_ (
);

AOI21X1 _9463_ (
    .A(_2806_),
    .B(_2813_),
    .C(_2788_),
    .Y(_2820_)
);

INVX2 _9043_ (
    .A(\X[3] [3]),
    .Y(_2406_)
);

FILL FILL_1__11711_ (
);

FILL FILL_2__8736_ (
);

FILL FILL_2__8316_ (
);

FILL FILL_0__10704_ (
);

FILL FILL_0__13176_ (
);

AOI21X1 _13041_ (
    .A(_5974_),
    .B(_6004_),
    .C(_6007_),
    .Y(_6077_)
);

FILL FILL_1__6733_ (
);

FILL FILL_3__6659_ (
);

FILL FILL_1__12916_ (
);

FILL FILL253950x219750 (
);

FILL FILL_0__9923_ (
);

FILL FILL_0__11909_ (
);

FILL FILL_0__9503_ (
);

FILL FILL_1__7938_ (
);

FILL FILL_3__10850_ (
);

FILL FILL_1__7518_ (
);

FILL FILL_3__10430_ (
);

FILL FILL_3__10010_ (
);

BUFX2 BUFX2_insert0 (
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf3 )
);

BUFX2 BUFX2_insert1 (
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf2 )
);

AOI22X1 _6588_ (
    .A(_111_),
    .B(_106_),
    .C(_183_),
    .D(_187_),
    .Y(_188_)
);

BUFX2 BUFX2_insert2 (
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf1 )
);

BUFX2 BUFX2_insert3 (
    .A(\X[1] [5]),
    .Y(\X[1]_5_bF$buf0 )
);

BUFX2 BUFX2_insert4 (
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf3 )
);

BUFX2 BUFX2_insert5 (
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf2 )
);

BUFX2 BUFX2_insert6 (
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf1 )
);

BUFX2 BUFX2_insert7 (
    .A(\X[3] [5]),
    .Y(\X[3]_5_bF$buf0 )
);

BUFX2 BUFX2_insert8 (
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf3 )
);

BUFX2 BUFX2_insert9 (
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf2 )
);

AND2X2 _10586_ (
    .A(_3851_),
    .B(_3850_),
    .Y(_3978_[4])
);

NAND3X1 _10166_ (
    .A(_3441_),
    .B(_3440_),
    .C(_3444_),
    .Y(_3445_)
);

FILL FILL_2__6802_ (
);

FILL FILL_3__11215_ (
);

FILL FILL_2__9694_ (
);

FILL FILL_2__10628_ (
);

FILL FILL_2__9274_ (
);

FILL FILL_0__11662_ (
);

FILL FILL_2__10208_ (
);

FILL FILL_0__11242_ (
);

FILL FILL_0__6628_ (
);

INVX1 _8734_ (
    .A(_2165_),
    .Y(_2168_)
);

AOI22X1 _8314_ (
    .A(vdd),
    .B(\X[2] [3]),
    .C(gnd),
    .D(\X[2] [4]),
    .Y(_1754_)
);

FILL FILL_1__7691_ (
);

FILL FILL_1__7271_ (
);

FILL FILL_1__13034_ (
);

FILL FILL_0__12867_ (
);

AOI21X1 _12732_ (
    .A(_5771_),
    .B(_5770_),
    .C(_5769_),
    .Y(_5772_)
);

FILL FILL_0__12447_ (
);

FILL FILL_0__12027_ (
);

NOR2X1 _12312_ (
    .A(_5413_),
    .B(_5418_),
    .Y(_5421_)
);

NAND2X1 _9939_ (
    .A(vdd),
    .B(\X[4] [3]),
    .Y(_3221_)
);

NAND2X1 _9519_ (
    .A(_2874_),
    .B(_2863_),
    .Y(_2875_)
);

FILL FILL_1__8896_ (
);

FILL FILL_1__8476_ (
);

FILL FILL_1__8056_ (
);

FILL FILL_2__10381_ (
);

FILL FILL_3__9763_ (
);

FILL FILL_0__6381_ (
);

FILL FILL_2__6399_ (
);

FILL FILL_2__7760_ (
);

FILL FILL254250x129750 (
);

FILL FILL_3__12593_ (
);

FILL FILL_2__7340_ (
);

FILL FILL_3__12173_ (
);

FILL FILL_2__11166_ (
);

FILL FILL_1__10999_ (
);

OAI21X1 _6800_ (
    .A(_322_),
    .B(_396_),
    .C(_343_),
    .Y(_397_)
);

FILL FILL_1__10579_ (
);

FILL FILL_1__10159_ (
);

FILL FILL_0__7586_ (
);

INVX1 _9692_ (
    .A(\u_fir_pe3.rYin [3]),
    .Y(_3039_)
);

FILL FILL_0__7166_ (
);

NAND2X1 _9272_ (
    .A(vdd),
    .B(\X[3] [6]),
    .Y(_2631_)
);

FILL FILL_1__11940_ (
);

FILL FILL_1__11520_ (
);

FILL FILL_1__11100_ (
);

FILL FILL_2__8545_ (
);

FILL FILL_0__10933_ (
);

FILL FILL_0__10513_ (
);

INVX1 _13270_ (
    .A(_6293_),
    .Y(_6294_)
);

FILL FILL_1__6962_ (
);

FILL FILL_1__6542_ (
);

FILL FILL_2__13312_ (
);

FILL FILL_3__6888_ (
);

FILL FILL_1__12725_ (
);

FILL FILL_1__12305_ (
);

FILL FILL_0__9732_ (
);

FILL FILL_0__9312_ (
);

FILL FILL_0__11718_ (
);

FILL FILL_1__7747_ (
);

FILL FILL_1__7327_ (
);

NAND2X1 _6397_ (
    .A(gnd),
    .B(Xin[2]),
    .Y(_0_)
);

FILL FILL_3__8614_ (
);

AND2X2 _10395_ (
    .A(_3664_),
    .B(_3670_),
    .Y(_3671_)
);

FILL FILL_2__6611_ (
);

FILL FILL_3__11444_ (
);

FILL FILL_2__10857_ (
);

FILL FILL_0__11891_ (
);

FILL FILL_2__10437_ (
);

FILL FILL_2__9083_ (
);

FILL FILL_0__11471_ (
);

FILL FILL_2__10017_ (
);

FILL FILL_0__11051_ (
);

FILL FILL_0__6857_ (
);

DFFPOSX1 _8963_ (
    .D(_2384_[10]),
    .CLK(clk_bF$buf17),
    .Q(\Y[3] [10])
);

FILL FILL_0__6437_ (
);

NAND2X1 _8543_ (
    .A(\X[2] [2]),
    .B(gnd),
    .Y(_1980_)
);

DFFPOSX1 _8123_ (
    .D(_1593_[7]),
    .CLK(clk_bF$buf52),
    .Q(\u_fir_pe1.mul [7])
);

FILL FILL_1__7080_ (
);

FILL FILL_2__7816_ (
);

FILL FILL_3__12229_ (
);

FILL FILL_1__13263_ (
);

OAI21X1 _12961_ (
    .A(_5604_),
    .B(_5995_),
    .C(_5997_),
    .Y(_5998_)
);

FILL FILL_0__12676_ (
);

FILL FILL_0__12256_ (
);

INVX1 _12541_ (
    .A(_5583_),
    .Y(_5584_)
);

NAND2X1 _12121_ (
    .A(_5236_),
    .B(_5079_),
    .Y(_5237_)
);

AND2X2 _9748_ (
    .A(_3050_),
    .B(_3060_),
    .Y(_3092_)
);

NAND3X1 _9328_ (
    .A(_2676_),
    .B(_2679_),
    .C(_2595_),
    .Y(_2686_)
);

FILL FILL_1__8285_ (
);

FILL FILL_2__10190_ (
);

FILL FILL_3__9992_ (
);

FILL FILL_3__9152_ (
);

OR2X2 _13326_ (
    .A(\u_fir_pe7.rYin [15]),
    .B(\u_fir_pe7.mul [15]),
    .Y(_6350_)
);

FILL FILL_2__11395_ (
);

FILL FILL_1__10388_ (
);

FILL FILL_0__7395_ (
);

NAND3X1 _9081_ (
    .A(_2419_),
    .B(_2442_),
    .C(_2441_),
    .Y(_2443_)
);

FILL FILL_2__8774_ (
);

FILL FILL_2__8354_ (
);

FILL FILL_3__13187_ (
);

FILL FILL_0__10322_ (
);

OAI21X1 _7814_ (
    .A(_1328_),
    .B(_1327_),
    .C(_1321_),
    .Y(_1329_)
);

FILL FILL_1__6771_ (
);

FILL FILL_2__13121_ (
);

FILL FILL_1__12954_ (
);

FILL FILL_1__12534_ (
);

FILL FILL_1__12114_ (
);

FILL FILL_2__9979_ (
);

FILL FILL_0__9961_ (
);

FILL FILL_0__9541_ (
);

FILL FILL_2__9559_ (
);

FILL FILL_0__11947_ (
);

FILL FILL_0__9121_ (
);

FILL FILL_2__9139_ (
);

NAND2X1 _11812_ (
    .A(_4931_),
    .B(_4923_),
    .Y(_4932_)
);

FILL FILL_0__11527_ (
);

FILL FILL_0__11107_ (
);

FILL FILL_1__7976_ (
);

FILL FILL_1__7556_ (
);

FILL FILL_1__7136_ (
);

FILL FILL_1__13319_ (
);

FILL FILL_3__8843_ (
);

FILL FILL_3__8003_ (
);

FILL FILL253650x205350 (
);

FILL FILL_2__6840_ (
);

FILL FILL_3__11673_ (
);

FILL FILL_2__6420_ (
);

FILL FILL_2__10666_ (
);

FILL FILL_2__10246_ (
);

FILL FILL_0__11280_ (
);

FILL FILL_1__9702_ (
);

FILL FILL_3__9628_ (
);

FILL FILL_0__6666_ (
);

NAND2X1 _8772_ (
    .A(_2183_),
    .B(_2182_),
    .Y(_2205_)
);

AOI21X1 _8352_ (
    .A(_1620_),
    .B(_1704_),
    .C(_1791_),
    .Y(_1792_)
);

FILL FILL_1__10600_ (
);

FILL FILL_2__7625_ (
);

FILL FILL_3__12458_ (
);

FILL FILL_1__13072_ (
);

AOI22X1 _12770_ (
    .A(gnd),
    .B(\X[6] [7]),
    .C(\X[6] [3]),
    .D(gnd),
    .Y(_5809_)
);

FILL FILL_0__12065_ (
);

OAI21X1 _12350_ (
    .A(_5447_),
    .B(_5448_),
    .C(_5452_),
    .Y(_5454_)
);

FILL FILL_2__12812_ (
);

NAND2X1 _9977_ (
    .A(\X[4] [0]),
    .B(vdd),
    .Y(_3258_)
);

NAND2X1 _9557_ (
    .A(gnd),
    .B(_2865_),
    .Y(_2912_)
);

AOI21X1 _9137_ (
    .A(_2419_),
    .B(_2439_),
    .C(_2453_),
    .Y(_2498_)
);

FILL FILL_1__11805_ (
);

FILL FILL_0__8812_ (
);

FILL FILL_3__9381_ (
);

NOR2X1 _13135_ (
    .A(_6168_),
    .B(_6167_),
    .Y(_6169_)
);

FILL FILL_1__6827_ (
);

FILL FILL_1__6407_ (
);

FILL FILL_1__9299_ (
);

FILL FILL_1__10197_ (
);

FILL FILL_3__10944_ (
);

FILL FILL_3__10524_ (
);

FILL FILL_3__10104_ (
);

FILL FILL_2__8583_ (
);

FILL FILL_0__10971_ (
);

FILL FILL_2__8163_ (
);

FILL FILL_0__10551_ (
);

FILL FILL_0__10131_ (
);

OAI21X1 _7623_ (
    .A(_1132_),
    .B(_1126_),
    .C(_1134_),
    .Y(_1141_)
);

DFFPOSX1 _7203_ (
    .D(_790_[4]),
    .CLK(clk_bF$buf52),
    .Q(\Y[1] [4])
);

FILL FILL_1__6580_ (
);

FILL FILL_3__11729_ (
);

FILL FILL_1__12763_ (
);

FILL FILL_3__11309_ (
);

FILL FILL_1__12343_ (
);

FILL FILL_2__9788_ (
);

FILL FILL_0__9770_ (
);

FILL FILL_0__9350_ (
);

FILL FILL_2__9368_ (
);

FILL FILL_0__11756_ (
);

DFFPOSX1 _11621_ (
    .D(\Y[5] [13]),
    .CLK(clk_bF$buf57),
    .Q(\u_fir_pe5.rYin [13])
);

FILL FILL_0__11336_ (
);

OAI21X1 _11201_ (
    .A(_4318_),
    .B(_4397_),
    .C(_4396_),
    .Y(_4398_)
);

INVX1 _8828_ (
    .A(_2244_),
    .Y(_2254_)
);

NAND3X1 _8408_ (
    .A(_1840_),
    .B(_1843_),
    .C(_1841_),
    .Y(_1847_)
);

FILL FILL_1__7785_ (
);

FILL FILL_1__7365_ (
);

FILL FILL_1__13128_ (
);

FILL FILL254550x108150 (
);

NAND3X1 _12826_ (
    .A(_5860_),
    .B(_5861_),
    .C(_5862_),
    .Y(_5865_)
);

FILL FILL_3__8232_ (
);

NOR2X1 _12406_ (
    .A(_5509_),
    .B(_5508_),
    .Y(_5510_)
);

FILL FILL_3__11062_ (
);

FILL FILL_2__10895_ (
);

FILL FILL_2__10475_ (
);

FILL FILL_2__10055_ (
);

FILL FILL_1__9931_ (
);

FILL FILL_1__9511_ (
);

FILL FILL_3__9017_ (
);

FILL FILL_0__6895_ (
);

FILL FILL_0__6475_ (
);

NAND2X1 _8581_ (
    .A(_2009_),
    .B(_2016_),
    .Y(_2018_)
);

INVX1 _8161_ (
    .A(_2334_),
    .Y(_1604_)
);

FILL FILL_2__7854_ (
);

FILL FILL_3__12687_ (
);

FILL FILL_2__7434_ (
);

FILL FILL_2__7014_ (
);

FILL FILL_0__12294_ (
);

FILL FILL_2__12621_ (
);

FILL FILL_2__12201_ (
);

AOI21X1 _9786_ (
    .A(_3126_),
    .B(_3117_),
    .C(_3124_),
    .Y(_3129_)
);

NAND2X1 _9366_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2724_)
);

FILL FILL_0__8621_ (
);

FILL FILL_2__8639_ (
);

FILL FILL_0__8201_ (
);

FILL FILL_2__8219_ (
);

FILL FILL_0__10607_ (
);

FILL FILL_0__13079_ (
);

DFFPOSX1 _13364_ (
    .D(\Y[6] [2]),
    .CLK(clk_bF$buf11),
    .Q(\u_fir_pe7.rYin [2])
);

FILL FILL_1__6636_ (
);

FILL FILL_2__13406_ (
);

FILL FILL_1__12819_ (
);

FILL FILL_0__9826_ (
);

FILL FILL_0__9406_ (
);

FILL FILL_3__7503_ (
);

FILL FILL_2__8392_ (
);

FILL FILL_0__10780_ (
);

FILL FILL_0__10360_ (
);

FILL FILL_3__8708_ (
);

AOI21X1 _7852_ (
    .A(gnd),
    .B(_1363_),
    .C(_1365_),
    .Y(_1366_)
);

OAI22X1 _7432_ (
    .A(_839_),
    .B(_950_),
    .C(_882_),
    .D(_951_),
    .Y(_952_)
);

NAND3X1 _7012_ (
    .A(_578_),
    .B(_580_),
    .C(_604_),
    .Y(_605_)
);

OAI21X1 _10489_ (
    .A(_3761_),
    .B(_3762_),
    .C(_3714_),
    .Y(_3763_)
);

INVX1 _10069_ (
    .A(_3348_),
    .Y(_3349_)
);

FILL FILL_3__11958_ (
);

FILL FILL_2__6705_ (
);

FILL FILL_1__12992_ (
);

FILL FILL_3__11538_ (
);

FILL FILL_1__12572_ (
);

FILL FILL_1__12152_ (
);

FILL FILL_0__11985_ (
);

FILL FILL_2__9597_ (
);

FILL FILL_2__9177_ (
);

AOI22X1 _11850_ (
    .A(_4893_),
    .B(_4888_),
    .C(_4965_),
    .D(_4969_),
    .Y(_4970_)
);

FILL FILL_0__11565_ (
);

NOR2X1 _11430_ (
    .A(_4617_),
    .B(_4618_),
    .Y(_4619_)
);

FILL FILL_0__11145_ (
);

OAI21X1 _11010_ (
    .A(_4158_),
    .B(_4208_),
    .C(_4152_),
    .Y(_4209_)
);

NAND2X1 _8637_ (
    .A(_2071_),
    .B(_2072_),
    .Y(_2073_)
);

AOI21X1 _8217_ (
    .A(_1655_),
    .B(_1658_),
    .C(_1649_),
    .Y(_1659_)
);

FILL FILL_1__7594_ (
);

FILL FILL_1__7174_ (
);

FILL FILL_3__8461_ (
);

INVX1 _12635_ (
    .A(_5663_),
    .Y(_5676_)
);

NAND2X1 _12215_ (
    .A(_5329_),
    .B(_5296_),
    .Y(_5330_)
);

FILL FILL_1__8799_ (
);

FILL FILL_1__8379_ (
);

FILL FILL_3__11291_ (
);

FILL FILL_2__10284_ (
);

FILL FILL_1__9740_ (
);

FILL FILL_1__9320_ (
);

FILL FILL_3__9246_ (
);

INVX1 _8390_ (
    .A(\X[2] [7]),
    .Y(_1829_)
);

FILL FILL_2__7663_ (
);

FILL FILL_3__12076_ (
);

FILL FILL_2__11489_ (
);

FILL FILL_2__11069_ (
);

INVX1 _6703_ (
    .A(_300_),
    .Y(_301_)
);

FILL FILL_2__12850_ (
);

FILL FILL_2__12430_ (
);

FILL FILL_2__12010_ (
);

FILL FILL_0__7489_ (
);

OAI21X1 _9595_ (
    .A(_2902_),
    .B(_2943_),
    .C(_2942_),
    .Y(_2949_)
);

FILL FILL_0__7069_ (
);

INVX2 _9175_ (
    .A(\X[3] [6]),
    .Y(_2535_)
);

FILL FILL_3__10809_ (
);

FILL FILL_1__11843_ (
);

FILL FILL_1__11423_ (
);

FILL FILL_1__11003_ (
);

FILL FILL_0__8850_ (
);

FILL FILL_2__8868_ (
);

FILL FILL_0__8430_ (
);

FILL FILL_2__8448_ (
);

FILL FILL_0__10836_ (
);

NOR2X1 _10701_ (
    .A(\u_fir_pe4.rYin [0]),
    .B(\u_fir_pe4.mul [0]),
    .Y(_3964_)
);

FILL FILL_0__10416_ (
);

FILL FILL_0__8010_ (
);

FILL FILL_2__8028_ (
);

INVX1 _13173_ (
    .A(_6195_),
    .Y(_6205_)
);

INVX1 _7908_ (
    .A(_1379_),
    .Y(_1420_)
);

FILL FILL_1__6865_ (
);

FILL FILL_1__6445_ (
);

FILL FILL_2__13215_ (
);

FILL FILL_1__12628_ (
);

FILL FILL_1__12208_ (
);

FILL FILL_0__9635_ (
);

FILL FILL_3__7732_ (
);

FILL FILL_0__9215_ (
);

NAND2X1 _11906_ (
    .A(_5023_),
    .B(_5024_),
    .Y(_5025_)
);

FILL FILL_3__10142_ (
);

FILL FILL_3__8937_ (
);

AOI21X1 _7661_ (
    .A(_1158_),
    .B(_1157_),
    .C(_1100_),
    .Y(_1178_)
);

DFFPOSX1 _7241_ (
    .D(_793_[2]),
    .CLK(clk_bF$buf16),
    .Q(\u_fir_pe0.mul [2])
);

NOR2X1 _10298_ (
    .A(_3506_),
    .B(_3509_),
    .Y(_3575_)
);

FILL FILL_2__6934_ (
);

FILL FILL_3__11767_ (
);

FILL FILL_2__6514_ (
);

FILL FILL_1__12381_ (
);

FILL FILL_0__11794_ (
);

FILL FILL_0__11374_ (
);

FILL FILL_2__11701_ (
);

OAI21X1 _8866_ (
    .A(_2259_),
    .B(_2260_),
    .C(_2288_),
    .Y(_2289_)
);

NOR2X1 _8446_ (
    .A(_1801_),
    .B(_1798_),
    .Y(_1885_)
);

AND2X2 _8026_ (
    .A(\u_fir_pe1.rYin [11]),
    .B(\u_fir_pe1.mul [11]),
    .Y(_1530_)
);

FILL FILL_0__7701_ (
);

FILL FILL_2__7719_ (
);

FILL FILL_1__13166_ (
);

FILL FILL_0__12999_ (
);

FILL FILL_3__8690_ (
);

OAI21X1 _12864_ (
    .A(_5819_),
    .B(_5827_),
    .C(_5826_),
    .Y(_5902_)
);

FILL FILL_0__12579_ (
);

FILL FILL_0__12159_ (
);

NOR2X1 _12444_ (
    .A(_5546_),
    .B(_5540_),
    .Y(_5548_)
);

NAND3X1 _12024_ (
    .A(_5135_),
    .B(_5136_),
    .C(_5137_),
    .Y(_5142_)
);

FILL FILL_2__12906_ (
);

FILL FILL_0__13100_ (
);

FILL FILL_1__8188_ (
);

FILL FILL_0__8906_ (
);

FILL FILL_2__10093_ (
);

FILL FILL_3__9475_ (
);

INVX1 _13229_ (
    .A(\u_fir_pe7.mul [6]),
    .Y(_6253_)
);

FILL FILL_2__7892_ (
);

FILL FILL_2__7472_ (
);

FILL FILL_2__7052_ (
);

FILL FILL_2__11298_ (
);

OAI22X1 _6932_ (
    .A(_233_),
    .B(_235_),
    .C(_319_),
    .D(_144_),
    .Y(_527_)
);

OAI21X1 _6512_ (
    .A(_108_),
    .B(_109_),
    .C(_69_),
    .Y(_113_)
);

FILL FILL_0__7298_ (
);

FILL FILL_3__10618_ (
);

FILL FILL_1__11652_ (
);

FILL FILL_1__11232_ (
);

FILL FILL_2__8677_ (
);

FILL FILL_2__8257_ (
);

FILL FILL_0__10645_ (
);

NAND2X1 _10930_ (
    .A(\X[5] [2]),
    .B(vdd),
    .Y(_4130_)
);

NOR2X1 _10510_ (
    .A(_3423_),
    .B(_3650_),
    .Y(_3783_)
);

FILL FILL_0__10225_ (
);

NAND3X1 _7717_ (
    .A(_1180_),
    .B(_1228_),
    .C(_1233_),
    .Y(_1234_)
);

FILL FILL_1__6674_ (
);

FILL FILL_2__13024_ (
);

FILL FILL_1__12857_ (
);

FILL FILL_1__12437_ (
);

FILL FILL_1__12017_ (
);

FILL FILL_0__9444_ (
);

FILL FILL_0__9024_ (
);

NAND2X1 _11715_ (
    .A(_4791_),
    .B(_4796_),
    .Y(_4837_)
);

FILL FILL_1__7879_ (
);

FILL FILL_3__10791_ (
);

FILL FILL_1__7459_ (
);

FILL FILL_3__10371_ (
);

FILL FILL_1__7039_ (
);

FILL FILL_1__8820_ (
);

FILL FILL_1__8400_ (
);

FILL FILL_3__8326_ (
);

OAI21X1 _7890_ (
    .A(_1360_),
    .B(_1373_),
    .C(_1377_),
    .Y(_1403_)
);

AOI21X1 _7470_ (
    .A(_989_),
    .B(_988_),
    .C(_987_),
    .Y(_990_)
);

NOR2X1 _7050_ (
    .A(_631_),
    .B(_636_),
    .Y(_639_)
);

FILL FILL_3__11996_ (
);

FILL FILL_2__6743_ (
);

FILL FILL_3__11156_ (
);

FILL FILL_1__12190_ (
);

FILL FILL_2__10989_ (
);

FILL FILL_2__10569_ (
);

FILL FILL_2__10149_ (
);

FILL FILL_0__11183_ (
);

FILL FILL_1__9605_ (
);

FILL FILL_2__11930_ (
);

FILL FILL_2__11510_ (
);

FILL FILL_0__6989_ (
);

FILL FILL_0__6569_ (
);

NAND2X1 _8675_ (
    .A(_2078_),
    .B(_2081_),
    .Y(_2110_)
);

NAND2X1 _8255_ (
    .A(_1675_),
    .B(_1671_),
    .Y(_1696_)
);

FILL FILL_1__10923_ (
);

FILL FILL_1__10503_ (
);

FILL FILL_2__7948_ (
);

FILL FILL_0__7930_ (
);

FILL FILL_0__7510_ (
);

FILL FILL_2__7528_ (
);

FILL FILL_2__7108_ (
);

FILL FILL_1__13395_ (
);

OR2X2 _12673_ (
    .A(_5712_),
    .B(_5710_),
    .Y(_5713_)
);

FILL FILL_0__12388_ (
);

NAND2X1 _12253_ (
    .A(_5364_),
    .B(_5366_),
    .Y(_5367_)
);

FILL FILL_3__13302_ (
);

FILL FILL_2__12715_ (
);

FILL FILL_1__11708_ (
);

FILL FILL_0__8715_ (
);

FILL FILL_3__6812_ (
);

NAND3X1 _13038_ (
    .A(_6039_),
    .B(_6073_),
    .C(_6071_),
    .Y(_6074_)
);

FILL FILL_2__7281_ (
);

NAND3X1 _6741_ (
    .A(_324_),
    .B(_326_),
    .C(_328_),
    .Y(_339_)
);

FILL FILL_1__11881_ (
);

FILL FILL_3__10427_ (
);

FILL FILL_1__11461_ (
);

FILL FILL_1__11041_ (
);

FILL FILL_2__8486_ (
);

FILL FILL_0__10874_ (
);

FILL FILL_0__10454_ (
);

FILL FILL_2__8066_ (
);

FILL FILL_0__10034_ (
);

INVX1 _7946_ (
    .A(\u_fir_pe1.rYin [4]),
    .Y(_1452_)
);

AOI22X1 _7526_ (
    .A(vdd),
    .B(\X[1] [4]),
    .C(vdd),
    .D(\X[1]_5_bF$buf3 ),
    .Y(_1045_)
);

NAND2X1 _7106_ (
    .A(_685_),
    .B(_688_),
    .Y(_790_[7])
);

FILL FILL_1__6483_ (
);

FILL FILL_2__13253_ (
);

FILL FILL_1__12666_ (
);

FILL FILL_1__12246_ (
);

FILL FILL_0__9673_ (
);

FILL FILL_3__7770_ (
);

FILL FILL_0__9253_ (
);

INVX1 _11944_ (
    .A(_4917_),
    .Y(_5063_)
);

FILL FILL_0__11659_ (
);

FILL FILL_3__7350_ (
);

INVX1 _11524_ (
    .A(_4707_),
    .Y(_4708_)
);

FILL FILL_0__11239_ (
);

OAI21X1 _11104_ (
    .A(_4223_),
    .B(_4301_),
    .C(_4245_),
    .Y(_4302_)
);

FILL FILL_0__12600_ (
);

FILL FILL_1__7688_ (
);

FILL FILL_1__7268_ (
);

FILL FILL_3__8555_ (
);

OAI21X1 _12729_ (
    .A(_5691_),
    .B(_5768_),
    .C(_5685_),
    .Y(_5769_)
);

FILL FILL_3__8135_ (
);

NOR2X1 _12309_ (
    .A(_5417_),
    .B(_5416_),
    .Y(_5418_)
);

FILL FILL_2__6972_ (
);

FILL FILL_2__6552_ (
);

FILL FILL_3__11385_ (
);

FILL FILL_2__10798_ (
);

FILL FILL_2__10378_ (
);

FILL FILL_1__9414_ (
);

FILL FILL_0__6798_ (
);

FILL FILL_0__6378_ (
);

OAI21X1 _8484_ (
    .A(_1683_),
    .B(_1738_),
    .C(_1921_),
    .Y(_1922_)
);

OR2X2 _8064_ (
    .A(\u_fir_pe1.rYin [15]),
    .B(\u_fir_pe1.mul [15]),
    .Y(_1568_)
);

FILL FILL_1__10312_ (
);

FILL FILL_2__7757_ (
);

FILL FILL_2__7337_ (
);

FILL FILL_0__12197_ (
);

DFFPOSX1 _12482_ (
    .D(\X[7]_5_bF$buf1 ),
    .CLK(clk_bF$buf37),
    .Q(_6376_[5])
);

OAI21X1 _12062_ (
    .A(_5104_),
    .B(_5178_),
    .C(_5125_),
    .Y(_5179_)
);

FILL FILL_3__13111_ (
);

FILL FILL_2__12944_ (
);

FILL FILL_2__12524_ (
);

FILL FILL_2__12104_ (
);

NAND2X1 _9689_ (
    .A(_3036_),
    .B(_3035_),
    .Y(_3037_)
);

NAND3X1 _9269_ (
    .A(_2616_),
    .B(_2625_),
    .C(_2627_),
    .Y(_2628_)
);

FILL FILL_1__11937_ (
);

FILL FILL_1__11517_ (
);

FILL FILL_0__8944_ (
);

FILL FILL_0__8524_ (
);

FILL FILL_3__9093_ (
);

AND2X2 _13267_ (
    .A(\u_fir_pe7.rYin [9]),
    .B(\u_fir_pe7.mul [9]),
    .Y(_6291_)
);

FILL FILL_2__9903_ (
);

FILL FILL_1__6959_ (
);

FILL FILL_1__6539_ (
);

FILL FILL_2__13309_ (
);

FILL FILL_2__7090_ (
);

FILL FILL_1__7900_ (
);

FILL FILL_0__9729_ (
);

FILL FILL_3__7826_ (
);

FILL FILL_0__9309_ (
);

INVX1 _6970_ (
    .A(_526_),
    .Y(_564_)
);

NAND2X1 _6550_ (
    .A(_149_),
    .B(_141_),
    .Y(_150_)
);

FILL FILL_1__11690_ (
);

FILL FILL_3__10236_ (
);

FILL FILL_1__11270_ (
);

FILL FILL_2__8295_ (
);

FILL FILL_0__10683_ (
);

FILL FILL_0__10263_ (
);

NOR2X1 _7755_ (
    .A(_1270_),
    .B(_1213_),
    .Y(_1271_)
);

OR2X2 _7335_ (
    .A(_856_),
    .B(_855_),
    .Y(_857_)
);

FILL FILL_2__13062_ (
);

FILL FILL_2__6608_ (
);

FILL FILL_1__12895_ (
);

FILL FILL_1__12055_ (
);

FILL FILL_0__9482_ (
);

FILL FILL_0__11888_ (
);

FILL FILL_0__9062_ (
);

NAND3X1 _11753_ (
    .A(vdd),
    .B(\X[7] [3]),
    .C(_4865_),
    .Y(_4874_)
);

FILL FILL_0__11468_ (
);

FILL FILL_0__11048_ (
);

INVX1 _11333_ (
    .A(_4500_),
    .Y(_4528_)
);

FILL FILL_1__7497_ (
);

FILL FILL_1__7077_ (
);

NAND2X1 _9901_ (
    .A(_3908_),
    .B(_3972_),
    .Y(_3973_)
);

FILL FILL_3__8784_ (
);

NAND2X1 _12958_ (
    .A(\X[6]_5_bF$buf2 ),
    .B(gnd),
    .Y(_5995_)
);

NAND2X1 _12538_ (
    .A(vdd),
    .B(\X[6] [0]),
    .Y(_5581_)
);

NAND2X1 _12118_ (
    .A(_5234_),
    .B(_5233_),
    .Y(_5578_[9])
);

FILL FILL_2__6781_ (
);

FILL FILL_2__10187_ (
);

FILL FILL_1__9643_ (
);

FILL FILL_1__9223_ (
);

FILL FILL_3__9569_ (
);

NAND2X1 _8293_ (
    .A(\X[2] [1]),
    .B(gnd),
    .Y(_1733_)
);

FILL FILL_1__10961_ (
);

FILL FILL_1__10541_ (
);

FILL FILL_1__10121_ (
);

FILL FILL_2__7986_ (
);

FILL FILL_2__7566_ (
);

FILL FILL_3__12399_ (
);

FILL FILL_2__7146_ (
);

NAND2X1 _12291_ (
    .A(_5402_),
    .B(_5401_),
    .Y(_5403_)
);

AOI21X1 _6606_ (
    .A(_194_),
    .B(_202_),
    .C(_205_),
    .Y(_206_)
);

FILL FILL_2__12753_ (
);

FILL FILL_2__12333_ (
);

NOR3X1 _9498_ (
    .A(_2696_),
    .B(_2523_),
    .C(_2712_),
    .Y(_2854_)
);

NAND3X1 _9078_ (
    .A(_2420_),
    .B(_2436_),
    .C(_2439_),
    .Y(_2440_)
);

FILL FILL_1__11746_ (
);

FILL FILL_1__11326_ (
);

FILL FILL_0__8753_ (
);

FILL FILL_0__8333_ (
);

FILL FILL_3__6430_ (
);

FILL FILL_0__10319_ (
);

AND2X2 _10604_ (
    .A(_3867_),
    .B(_3866_),
    .Y(_3978_[6])
);

FILL FILL_0_BUFX2_insert70 (
);

FILL FILL_0_BUFX2_insert71 (
);

FILL FILL_0_BUFX2_insert72 (
);

FILL FILL_0_BUFX2_insert73 (
);

FILL FILL254550x212550 (
);

FILL FILL_0_BUFX2_insert74 (
);

FILL FILL_0_BUFX2_insert75 (
);

FILL FILL_0_BUFX2_insert76 (
);

FILL FILL_0_BUFX2_insert77 (
);

FILL FILL_0_BUFX2_insert78 (
);

OAI21X1 _13076_ (
    .A(_6110_),
    .B(_6109_),
    .C(_6103_),
    .Y(_6111_)
);

FILL FILL_0_BUFX2_insert79 (
);

FILL FILL_2__9712_ (
);

FILL FILL_1__6768_ (
);

FILL FILL_2__13118_ (
);

FILL FILL_0__9958_ (
);

FILL FILL_0__9538_ (
);

FILL FILL_0__9118_ (
);

NAND3X1 _11809_ (
    .A(_4928_),
    .B(_4922_),
    .C(_4925_),
    .Y(_4929_)
);

FILL FILL_3__10885_ (
);

FILL FILL_3__10465_ (
);

FILL FILL_3__10045_ (
);

FILL FILL_0__10492_ (
);

FILL FILL_0__10072_ (
);

FILL FILL_1__8914_ (
);

INVX1 _7984_ (
    .A(\u_fir_pe1.rYin [8]),
    .Y(_1487_)
);

NAND3X1 _7564_ (
    .A(_1078_),
    .B(_1079_),
    .C(_1080_),
    .Y(_1083_)
);

NOR2X1 _7144_ (
    .A(_727_),
    .B(_726_),
    .Y(_728_)
);

FILL FILL_2__13291_ (
);

FILL FILL_2__6837_ (
);

FILL FILL_2__6417_ (
);

FILL FILL_1__12284_ (
);

NAND2X1 _11982_ (
    .A(\X[7] [3]),
    .B(gnd),
    .Y(_5100_)
);

FILL FILL_0__9291_ (
);

FILL FILL_0__11697_ (
);

INVX1 _11562_ (
    .A(\u_fir_pe5.mul [14]),
    .Y(_4746_)
);

FILL FILL_0__11277_ (
);

OAI21X1 _11142_ (
    .A(_4326_),
    .B(_4330_),
    .C(_4333_),
    .Y(_4340_)
);

FILL FILL_3__12611_ (
);

NAND2X1 _8769_ (
    .A(_2200_),
    .B(_2201_),
    .Y(_2202_)
);

AOI21X1 _8349_ (
    .A(_1712_),
    .B(_1711_),
    .C(_1648_),
    .Y(_1789_)
);

FILL FILL_0__7604_ (
);

OAI21X1 _9710_ (
    .A(_3046_),
    .B(_3047_),
    .C(_3053_),
    .Y(_3055_)
);

FILL FILL_1__13069_ (
);

AND2X2 _12767_ (
    .A(\X[6] [3]),
    .B(gnd),
    .Y(_5806_)
);

FILL FILL_3__8173_ (
);

NAND2X1 _12347_ (
    .A(_5451_),
    .B(_5446_),
    .Y(_5452_)
);

FILL FILL_2__12809_ (
);

FILL FILL_0__13003_ (
);

FILL FILL_2__6590_ (
);

FILL FILL_0__8809_ (
);

FILL FILL_3__6906_ (
);

FILL FILL_1__9452_ (
);

FILL FILL_1__9032_ (
);

FILL FILL_3__9798_ (
);

FILL FILL_1__10770_ (
);

FILL FILL_1__10350_ (
);

FILL FILL_2__7795_ (
);

FILL FILL_2__7375_ (
);

INVX1 _6835_ (
    .A(_354_),
    .Y(_432_)
);

NAND2X1 _6415_ (
    .A(_14_),
    .B(_17_),
    .Y(_18_)
);

FILL FILL_2__12982_ (
);

FILL FILL_2__12562_ (
);

FILL FILL_2__12142_ (
);

FILL FILL_1__11975_ (
);

FILL FILL_1__11555_ (
);

FILL FILL_1__11135_ (
);

FILL FILL_0__8562_ (
);

FILL FILL_0__10968_ (
);

FILL FILL_0__8142_ (
);

FILL FILL_0__10548_ (
);

NAND2X1 _10833_ (
    .A(_4017_),
    .B(_4032_),
    .Y(_4035_)
);

NAND3X1 _10413_ (
    .A(_3684_),
    .B(_3685_),
    .C(_3688_),
    .Y(_3689_)
);

FILL FILL_0__10128_ (
);

FILL FILL_2__9941_ (
);

FILL FILL_2__9521_ (
);

FILL FILL_2__9101_ (
);

FILL FILL_1__6997_ (
);

FILL FILL_1__6577_ (
);

FILL FILL_0__9767_ (
);

FILL FILL_3__7864_ (
);

FILL FILL_0__9347_ (
);

FILL FILL_3__7444_ (
);

DFFPOSX1 _11618_ (
    .D(\Y[5] [10]),
    .CLK(clk_bF$buf18),
    .Q(\u_fir_pe5.rYin [10])
);

FILL FILL_3__7024_ (
);

FILL FILL_3__10694_ (
);

FILL FILL_1__8723_ (
);

FILL FILL_1__8303_ (
);

FILL FILL_3__8649_ (
);

FILL FILL_3__8229_ (
);

NAND3X1 _7793_ (
    .A(_1292_),
    .B(_1298_),
    .C(_1256_),
    .Y(_1308_)
);

INVX1 _7373_ (
    .A(_881_),
    .Y(_894_)
);

FILL FILL_2__6646_ (
);

FILL FILL_3__11479_ (
);

FILL FILL_1__12093_ (
);

OAI21X1 _11791_ (
    .A(_4910_),
    .B(_4911_),
    .C(_4909_),
    .Y(_4912_)
);

FILL FILL_0__11086_ (
);

NAND3X1 _11371_ (
    .A(_4546_),
    .B(_4563_),
    .C(_4562_),
    .Y(_4565_)
);

FILL FILL_1__9928_ (
);

FILL FILL_3__12840_ (
);

FILL FILL_1__9508_ (
);

FILL FILL_3__12000_ (
);

FILL FILL_2__11833_ (
);

FILL FILL_2__11413_ (
);

DFFPOSX1 _8998_ (
    .D(_2390_[5]),
    .CLK(clk_bF$buf51),
    .Q(\u_fir_pe2.mul [5])
);

NAND2X1 _8578_ (
    .A(_2000_),
    .B(_2003_),
    .Y(_2015_)
);

NOR2X1 _8158_ (
    .A(_2325_),
    .B(_1596_),
    .Y(_1601_)
);

FILL FILL_1__10826_ (
);

FILL FILL_1__10406_ (
);

FILL FILL_0__7833_ (
);

FILL FILL_0__7413_ (
);

FILL FILL_1__13298_ (
);

NAND2X1 _12996_ (
    .A(_6021_),
    .B(_6028_),
    .Y(_6032_)
);

INVX1 _12576_ (
    .A(_5617_),
    .Y(_5618_)
);

NAND3X1 _12156_ (
    .A(_5189_),
    .B(_5265_),
    .C(_5197_),
    .Y(_5272_)
);

FILL FILL_2__12618_ (
);

FILL FILL_0__13232_ (
);

FILL FILL_0__8618_ (
);

FILL FILL_1__9681_ (
);

FILL FILL_1__9261_ (
);

FILL FILL_3__9187_ (
);

FILL FILL_2__7184_ (
);

NAND2X1 _6644_ (
    .A(_241_),
    .B(_242_),
    .Y(_243_)
);

FILL FILL_2__12791_ (
);

FILL FILL_2__12371_ (
);

FILL FILL_1__11784_ (
);

FILL FILL_1__11364_ (
);

FILL FILL_0__8791_ (
);

FILL FILL_2__8389_ (
);

FILL FILL_0__8371_ (
);

FILL FILL_0__10777_ (
);

FILL FILL_0__10357_ (
);

NAND2X1 _10642_ (
    .A(_3905_),
    .B(_3904_),
    .Y(_3978_[9])
);

OR2X2 _10222_ (
    .A(_3495_),
    .B(_3494_),
    .Y(_3500_)
);

FILL FILL_2__9750_ (
);

FILL FILL_2__9330_ (
);

NOR2X1 _7849_ (
    .A(_1270_),
    .B(_1323_),
    .Y(_1363_)
);

AND2X2 _7429_ (
    .A(_944_),
    .B(_948_),
    .Y(_949_)
);

NAND2X1 _7009_ (
    .A(_594_),
    .B(_601_),
    .Y(_602_)
);

FILL FILL_1__6386_ (
);

FILL FILL_2__13156_ (
);

FILL FILL_1__12989_ (
);

FILL FILL_1__12569_ (
);

FILL FILL_1__12149_ (
);

FILL FILL_0__9996_ (
);

FILL FILL_0__9576_ (
);

FILL FILL_3__7673_ (
);

FILL FILL_0__9156_ (
);

OAI21X1 _11847_ (
    .A(_4962_),
    .B(_4963_),
    .C(_4920_),
    .Y(_4967_)
);

AND2X2 _11427_ (
    .A(\u_fir_pe5.rYin [0]),
    .B(\u_fir_pe5.mul [0]),
    .Y(_4616_)
);

OAI21X1 _11007_ (
    .A(_4204_),
    .B(_4205_),
    .C(_4195_),
    .Y(_4206_)
);

FILL FILL_0__12923_ (
);

FILL FILL_3__10083_ (
);

FILL FILL_1__8952_ (
);

FILL FILL_1__8532_ (
);

FILL FILL_3__8878_ (
);

FILL FILL_3__8038_ (
);

NOR2X1 _7182_ (
    .A(_764_),
    .B(_758_),
    .Y(_766_)
);

FILL FILL_2__6875_ (
);

FILL FILL_2__6455_ (
);

INVX1 _11180_ (
    .A(_4371_),
    .Y(_4377_)
);

FILL FILL_1__9737_ (
);

FILL FILL_1__9317_ (
);

FILL FILL_2__11642_ (
);

FILL FILL_2__11222_ (
);

NAND3X1 _8387_ (
    .A(_1820_),
    .B(_1825_),
    .C(_1823_),
    .Y(_1826_)
);

FILL FILL_1__10635_ (
);

FILL FILL_1__10215_ (
);

FILL FILL_0__7642_ (
);

NAND2X1 _12385_ (
    .A(_5487_),
    .B(_5488_),
    .Y(_5489_)
);

FILL FILL_2__8601_ (
);

FILL FILL_3__13014_ (
);

FILL FILL_2__12847_ (
);

FILL FILL_2__12427_ (
);

FILL FILL_2__12007_ (
);

FILL FILL_0__13041_ (
);

FILL FILL_0__8847_ (
);

FILL FILL_0__8427_ (
);

FILL FILL_3__6524_ (
);

FILL FILL_0__8007_ (
);

FILL FILL_1__9490_ (
);

FILL FILL_1__9070_ (
);

FILL FILL_2__9806_ (
);

FILL FILL_1__7803_ (
);

FILL FILL_3__7309_ (
);

NAND3X1 _6873_ (
    .A(_467_),
    .B(_464_),
    .C(_468_),
    .Y(_469_)
);

NAND2X1 _6453_ (
    .A(_9_),
    .B(_14_),
    .Y(_55_)
);

FILL FILL_2__12180_ (
);

FILL FILL_3__10979_ (
);

FILL FILL_3__10559_ (
);

FILL FILL_3__10139_ (
);

FILL FILL_1__11173_ (
);

FILL FILL_2__8198_ (
);

FILL FILL_0__8180_ (
);

FILL FILL_0__10586_ (
);

AND2X2 _10871_ (
    .A(gnd),
    .B(\X[5] [3]),
    .Y(_4072_)
);

AOI21X1 _10451_ (
    .A(_3603_),
    .B(_3595_),
    .C(_3673_),
    .Y(_3726_)
);

FILL FILL_0__10166_ (
);

NAND3X1 _10031_ (
    .A(_3241_),
    .B(_3305_),
    .C(_3306_),
    .Y(_3312_)
);

BUFX2 BUFX2_insert80 (
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf1 )
);

BUFX2 BUFX2_insert81 (
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf0 )
);

BUFX2 BUFX2_insert82 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf3)
);

BUFX2 BUFX2_insert83 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf2)
);

BUFX2 BUFX2_insert84 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf1)
);

BUFX2 BUFX2_insert85 (
    .A(Xin[5]),
    .Y(Xin_5_bF$buf0)
);

BUFX2 BUFX2_insert86 (
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf3 )
);

BUFX2 BUFX2_insert87 (
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf2 )
);

FILL FILL_2__10913_ (
);

BUFX2 BUFX2_insert88 (
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf1 )
);

BUFX2 BUFX2_insert89 (
    .A(\X[7] [5]),
    .Y(\X[7]_5_bF$buf0 )
);

NAND2X1 _7658_ (
    .A(_1171_),
    .B(_1175_),
    .Y(_1593_[8])
);

DFFPOSX1 _7238_ (
    .D(Yin[15]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.rYin [15])
);

FILL FILL_0__6913_ (
);

FILL FILL_1__12798_ (
);

FILL FILL_1__12378_ (
);

FILL FILL_0__9385_ (
);

INVX1 _11656_ (
    .A(_5567_),
    .Y(_5568_)
);

AOI21X1 _11236_ (
    .A(_4421_),
    .B(_4416_),
    .C(_4368_),
    .Y(_4433_)
);

FILL FILL_0__12732_ (
);

FILL FILL_0__12312_ (
);

OR2X2 _9804_ (
    .A(_3140_),
    .B(_3146_),
    .Y(_3148_)
);

FILL FILL_1__8761_ (
);

FILL FILL_1__8341_ (
);

FILL FILL_3__8267_ (
);

FILL FILL_2__6684_ (
);

FILL FILL_3__11097_ (
);

FILL FILL_1__9966_ (
);

FILL FILL_1__9546_ (
);

FILL FILL_1__9126_ (
);

FILL FILL_2__11871_ (
);

FILL FILL_2__11451_ (
);

FILL FILL_2__11031_ (
);

NAND3X1 _8196_ (
    .A(_1627_),
    .B(_1635_),
    .C(_1637_),
    .Y(_1638_)
);

FILL FILL_1__10864_ (
);

FILL FILL_1__10444_ (
);

FILL FILL_1__10024_ (
);

FILL FILL_2__7889_ (
);

FILL FILL_0__7871_ (
);

FILL FILL_2__7469_ (
);

FILL FILL_0__7451_ (
);

FILL FILL_2__7049_ (
);

FILL FILL_0__7031_ (
);

OAI22X1 _12194_ (
    .A(_5015_),
    .B(_5017_),
    .C(_5101_),
    .D(_4926_),
    .Y(_5309_)
);

FILL FILL_2__8830_ (
);

FILL FILL_2__8410_ (
);

NAND2X1 _6929_ (
    .A(_519_),
    .B(_523_),
    .Y(_524_)
);

OAI21X1 _6509_ (
    .A(_108_),
    .B(_109_),
    .C(_107_),
    .Y(_110_)
);

FILL FILL_2__12656_ (
);

FILL FILL_2__12236_ (
);

FILL FILL_0__13270_ (
);

FILL FILL_1__11649_ (
);

FILL FILL_1__11229_ (
);

FILL FILL_0__8656_ (
);

FILL FILL_3__6753_ (
);

FILL FILL_0__8236_ (
);

AND2X2 _10927_ (
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4127_)
);

INVX1 _10507_ (
    .A(_3754_),
    .Y(_3780_)
);

BUFX2 _13399_ (
    .A(_6376_[5]),
    .Y(Xout[5])
);

FILL FILL_2__9615_ (
);

FILL FILL_1__7612_ (
);

FILL FILL_3__7538_ (
);

FILL FILL_3__7118_ (
);

INVX1 _6682_ (
    .A(_135_),
    .Y(_281_)
);

FILL FILL_3__10368_ (
);

FILL FILL_0__10395_ (
);

NAND2X1 _10680_ (
    .A(_3943_),
    .B(_3937_),
    .Y(_3944_)
);

NAND3X1 _10260_ (
    .A(_3510_),
    .B(_3528_),
    .C(_3524_),
    .Y(_3538_)
);

FILL FILL_1__8817_ (
);

FILL FILL_2__10302_ (
);

OR2X2 _7887_ (
    .A(_1398_),
    .B(_1391_),
    .Y(_1400_)
);

OAI21X1 _7467_ (
    .A(_909_),
    .B(_986_),
    .C(_903_),
    .Y(_987_)
);

NOR2X1 _7047_ (
    .A(_635_),
    .B(_634_),
    .Y(_636_)
);

FILL FILL_2__13194_ (
);

FILL FILL_0__6722_ (
);

FILL FILL_1__12187_ (
);

FILL FILL_0__9194_ (
);

NAND2X1 _11885_ (
    .A(_5000_),
    .B(_5003_),
    .Y(_5004_)
);

FILL FILL_3__7291_ (
);

INVX1 _11465_ (
    .A(\u_fir_pe5.rYin [5]),
    .Y(_4650_)
);

AND2X2 _11045_ (
    .A(_4222_),
    .B(_4217_),
    .Y(_4244_)
);

FILL FILL_3__12934_ (
);

FILL FILL_2__11927_ (
);

FILL FILL_0__12961_ (
);

FILL FILL_2__11507_ (
);

FILL FILL_0__12541_ (
);

FILL FILL_0__12121_ (
);

FILL FILL_0__7927_ (
);

FILL FILL_0__7507_ (
);

NAND2X1 _9613_ (
    .A(_2963_),
    .B(_2966_),
    .Y(_2967_)
);

FILL FILL_1__8570_ (
);

FILL FILL_1__8150_ (
);

FILL FILL_3__8496_ (
);

FILL FILL_0__13326_ (
);

FILL FILL_2__6493_ (
);

FILL FILL_1__9775_ (
);

FILL FILL_1__9355_ (
);

FILL FILL_2__11680_ (
);

FILL FILL_2__11260_ (
);

FILL FILL_1__10673_ (
);

FILL FILL_1__10253_ (
);

FILL FILL_2__7698_ (
);

FILL FILL_0__7680_ (
);

FILL FILL_0__7260_ (
);

FILL FILL_2__7278_ (
);

FILL FILL_3__13052_ (
);

OAI21X1 _6738_ (
    .A(_335_),
    .B(_329_),
    .C(_323_),
    .Y(_336_)
);

FILL FILL_2__12885_ (
);

FILL FILL_2__12045_ (
);

FILL FILL_1__11878_ (
);

FILL FILL_1__11458_ (
);

FILL FILL_1__11038_ (
);

FILL FILL_0__8885_ (
);

FILL FILL_3__6982_ (
);

FILL FILL_0__8465_ (
);

DFFPOSX1 _10736_ (
    .D(\Y[4] [5]),
    .CLK(clk_bF$buf10),
    .Q(\u_fir_pe4.rYin [5])
);

FILL FILL_0__8045_ (
);

AND2X2 _10316_ (
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3593_)
);

FILL FILL_2__9424_ (
);

FILL FILL_0__11812_ (
);

FILL FILL_3_CLKBUF1_insert60 (
);

FILL FILL_3_CLKBUF1_insert61 (
);

FILL FILL_3_CLKBUF1_insert63 (
);

FILL FILL_3_CLKBUF1_insert65 (
);

FILL FILL_1__7841_ (
);

FILL FILL_3_CLKBUF1_insert67 (
);

FILL FILL_1__7421_ (
);

FILL FILL_1__7001_ (
);

FILL FILL_3_CLKBUF1_insert69 (
);

FILL FILL_3__7767_ (
);

NAND3X1 _6491_ (
    .A(vdd),
    .B(Xin[3]),
    .C(_83_),
    .Y(_92_)
);

FILL FILL_3__10177_ (
);

FILL FILL_1__8626_ (
);

FILL FILL_1__8206_ (
);

FILL FILL_2__10951_ (
);

FILL FILL_2__10531_ (
);

FILL FILL_2__10111_ (
);

NAND2X1 _7696_ (
    .A(\X[1]_5_bF$buf0 ),
    .B(gnd),
    .Y(_1213_)
);

NAND2X1 _7276_ (
    .A(vdd),
    .B(\X[1] [0]),
    .Y(_799_)
);

FILL FILL_3__9913_ (
);

FILL FILL_2__6969_ (
);

FILL FILL_0__6951_ (
);

FILL FILL_2__6549_ (
);

FILL FILL_0__6531_ (
);

INVX1 _11694_ (
    .A(_4815_),
    .Y(_4816_)
);

NAND2X1 _11274_ (
    .A(_4467_),
    .B(_4461_),
    .Y(_4470_)
);

FILL FILL_2__7910_ (
);

FILL FILL_3__12323_ (
);

FILL FILL_2__11736_ (
);

FILL FILL_0__12770_ (
);

FILL FILL_2__11316_ (
);

FILL FILL_0__12350_ (
);

FILL FILL_1__10309_ (
);

FILL FILL_0__7736_ (
);

DFFPOSX1 _9842_ (
    .D(_3181_[12]),
    .CLK(clk_bF$buf12),
    .Q(\Y[4] [12])
);

FILL FILL_0__7316_ (
);

NAND2X1 _9422_ (
    .A(gnd),
    .B(_2778_),
    .Y(_2779_)
);

DFFPOSX1 _9002_ (
    .D(_2390_[9]),
    .CLK(clk_bF$buf51),
    .Q(\u_fir_pe2.mul [9])
);

INVX1 _12899_ (
    .A(_5850_),
    .Y(_5937_)
);

DFFPOSX1 _12479_ (
    .D(\X[7] [2]),
    .CLK(clk_bF$buf37),
    .Q(_6376_[2])
);

NAND3X1 _12059_ (
    .A(_5174_),
    .B(_5170_),
    .C(_5175_),
    .Y(_5176_)
);

FILL FILL_3__13108_ (
);

FILL FILL_0__13135_ (
);

AOI21X1 _13000_ (
    .A(_5951_),
    .B(_6021_),
    .C(_6035_),
    .Y(_6036_)
);

FILL FILL_3__6618_ (
);

FILL FILL_1__9584_ (
);

FILL FILL_1__9164_ (
);

FILL FILL_1__10482_ (
);

FILL FILL_1__10062_ (
);

FILL FILL_2__7087_ (
);

FILL FILL_3__13281_ (
);

OAI21X1 _6967_ (
    .A(_305_),
    .B(_479_),
    .C(_523_),
    .Y(_561_)
);

NAND3X1 _6547_ (
    .A(_146_),
    .B(_140_),
    .C(_143_),
    .Y(_147_)
);

FILL FILL_2__12694_ (
);

FILL FILL_2__12274_ (
);

FILL FILL_1__11687_ (
);

FILL FILL_1__11267_ (
);

FILL FILL_0__8694_ (
);

FILL FILL_0__8274_ (
);

AOI21X1 _10965_ (
    .A(_4159_),
    .B(_4160_),
    .C(_4158_),
    .Y(_4165_)
);

NAND2X1 _10545_ (
    .A(_3816_),
    .B(_3810_),
    .Y(_3984_[14])
);

NAND2X1 _10125_ (
    .A(_3401_),
    .B(_3403_),
    .Y(_3404_)
);

FILL FILL_2__9653_ (
);

FILL FILL_2__9233_ (
);

FILL FILL_0__11201_ (
);

FILL FILL_2__13059_ (
);

FILL FILL_1__7650_ (
);

FILL FILL_0__9899_ (
);

FILL FILL_0__9479_ (
);

FILL FILL_0__9059_ (
);

FILL FILL_1__13413_ (
);

FILL FILL_0__12826_ (
);

FILL FILL_0__12406_ (
);

FILL FILL_1__8855_ (
);

FILL FILL_1__8435_ (
);

FILL FILL_1__8015_ (
);

FILL FILL_2__10340_ (
);

NAND2X1 _7085_ (
    .A(_669_),
    .B(_664_),
    .Y(_670_)
);

FILL FILL_3__9722_ (
);

FILL FILL_2__6778_ (
);

FILL FILL_0__6760_ (
);

AOI21X1 _11083_ (
    .A(_4192_),
    .B(_4270_),
    .C(_4278_),
    .Y(_4281_)
);

FILL FILL_3__12552_ (
);

FILL FILL_2__11965_ (
);

FILL FILL_2__11545_ (
);

FILL FILL_2__11125_ (
);

FILL FILL_1__10958_ (
);

FILL FILL_1__10538_ (
);

FILL FILL_1__10118_ (
);

FILL FILL_0__7965_ (
);

FILL FILL_0__7545_ (
);

NAND3X1 _9651_ (
    .A(_2975_),
    .B(_3003_),
    .C(_3002_),
    .Y(_3004_)
);

FILL FILL_0__7125_ (
);

AOI21X1 _9231_ (
    .A(_2573_),
    .B(_2568_),
    .C(_2575_),
    .Y(_2591_)
);

AND2X2 _12288_ (
    .A(_5378_),
    .B(_5377_),
    .Y(_5400_)
);

FILL FILL_2__8924_ (
);

FILL FILL_2__8504_ (
);

FILL FILL_3__13337_ (
);

FILL FILL_1__6921_ (
);

FILL FILL_1__6501_ (
);

FILL FILL_3__6847_ (
);

FILL FILL_1__9393_ (
);

FILL FILL_2__9709_ (
);

FILL FILL_1__10291_ (
);

FILL FILL_1__7706_ (
);

NAND2X1 _6776_ (
    .A(_373_),
    .B(_297_),
    .Y(_374_)
);

FILL FILL_2__12083_ (
);

FILL FILL_1__11496_ (
);

FILL FILL_1__11076_ (
);

FILL FILL_0__10489_ (
);

NAND2X1 _10774_ (
    .A(_4765_),
    .B(_4745_),
    .Y(_4766_)
);

INVX1 _10354_ (
    .A(_3552_),
    .Y(_3631_)
);

FILL FILL_0__10069_ (
);

FILL FILL_3__11823_ (
);

FILL FILL_3__11403_ (
);

FILL FILL_2__10816_ (
);

FILL FILL_2__9462_ (
);

FILL FILL_0__11850_ (
);

FILL FILL_2__9042_ (
);

FILL FILL_0__11430_ (
);

FILL FILL_0__11010_ (
);

FILL FILL_2__13288_ (
);

FILL FILL_0__6816_ (
);

INVX1 _8922_ (
    .A(\u_fir_pe2.mul [13]),
    .Y(_2346_)
);

OAI21X1 _8502_ (
    .A(_1935_),
    .B(_1939_),
    .C(_1911_),
    .Y(_1940_)
);

FILL FILL_0__9288_ (
);

NAND2X1 _11979_ (
    .A(_5092_),
    .B(_5096_),
    .Y(_5097_)
);

FILL FILL_3__7385_ (
);

AND2X2 _11559_ (
    .A(_4742_),
    .B(_4741_),
    .Y(_4775_[13])
);

AOI21X1 _11139_ (
    .A(_4336_),
    .B(_4331_),
    .C(_4300_),
    .Y(_4337_)
);

FILL FILL_3__12608_ (
);

FILL FILL_1__13222_ (
);

FILL FILL_0__12635_ (
);

NAND2X1 _12920_ (
    .A(_5953_),
    .B(_5957_),
    .Y(_6375_[8])
);

FILL FILL_0__12215_ (
);

DFFPOSX1 _12500_ (
    .D(\Y[7] [15]),
    .CLK(clk_bF$buf11),
    .Q(\u_fir_pe6.rYin [15])
);

NAND2X1 _9707_ (
    .A(_3050_),
    .B(_3052_),
    .Y(_3053_)
);

FILL FILL_1__8664_ (
);

FILL FILL_1__8244_ (
);

FILL FILL_3__9111_ (
);

FILL FILL_2__6587_ (
);

FILL FILL_3__12781_ (
);

FILL FILL_1__9449_ (
);

FILL FILL_1__9029_ (
);

FILL FILL_2__11774_ (
);

FILL FILL_2__11354_ (
);

DFFPOSX1 _8099_ (
    .D(\X[1] [7]),
    .CLK(clk_bF$buf54),
    .Q(\X[2] [7])
);

FILL FILL_1__10767_ (
);

FILL FILL_1__10347_ (
);

FILL FILL_0__7774_ (
);

DFFPOSX1 _9880_ (
    .D(_3187_[10]),
    .CLK(clk_bF$buf36),
    .Q(\u_fir_pe3.mul [10])
);

FILL FILL_0__7354_ (
);

NAND3X1 _9460_ (
    .A(_2786_),
    .B(_2814_),
    .C(_2816_),
    .Y(_2817_)
);

OAI21X1 _9040_ (
    .A(_2395_),
    .B(_2398_),
    .C(_2392_),
    .Y(_2403_)
);

INVX1 _12097_ (
    .A(_5136_),
    .Y(_5214_)
);

FILL FILL_2__8733_ (
);

FILL FILL_2__8313_ (
);

FILL FILL_0__10701_ (
);

FILL FILL_2__12979_ (
);

FILL FILL_2__12559_ (
);

FILL FILL_2__12139_ (
);

FILL FILL_0__13173_ (
);

FILL FILL_1__6730_ (
);

FILL FILL_0__8559_ (
);

FILL FILL_0__8139_ (
);

FILL FILL_1__12913_ (
);

FILL FILL_0__9920_ (
);

FILL FILL_2__9938_ (
);

FILL FILL_0__11906_ (
);

FILL FILL_0__9500_ (
);

FILL FILL_2__9518_ (
);

FILL FILL_1__7935_ (
);

FILL FILL_1__7515_ (
);

OAI21X1 _6585_ (
    .A(_180_),
    .B(_181_),
    .C(_138_),
    .Y(_185_)
);

FILL FILL_3__8802_ (
);

FILL FILL_0__10298_ (
);

OAI21X1 _10583_ (
    .A(_3839_),
    .B(_3835_),
    .C(_3848_),
    .Y(_3849_)
);

NAND2X1 _10163_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf3 ),
    .Y(_3442_)
);

FILL FILL_2__9691_ (
);

FILL FILL_2__10625_ (
);

FILL FILL_2__9271_ (
);

FILL FILL_2__10205_ (
);

FILL FILL_2__13097_ (
);

FILL FILL_0__6625_ (
);

NAND2X1 _8731_ (
    .A(_2159_),
    .B(_2163_),
    .Y(_2165_)
);

INVX1 _8311_ (
    .A(_1750_),
    .Y(_1751_)
);

FILL FILL_0__9097_ (
);

INVX1 _11788_ (
    .A(_4849_),
    .Y(_4909_)
);

FILL FILL_3__7194_ (
);

NAND2X1 _11368_ (
    .A(_4548_),
    .B(_4561_),
    .Y(_4562_)
);

FILL FILL_3__12837_ (
);

FILL FILL_3__12417_ (
);

FILL FILL_1__13031_ (
);

FILL FILL_0__12864_ (
);

FILL FILL_0__12444_ (
);

FILL FILL_0__12024_ (
);

NAND2X1 _9936_ (
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3218_)
);

AOI21X1 _9516_ (
    .A(gnd),
    .B(\X[3] [6]),
    .C(_2803_),
    .Y(_2872_)
);

FILL FILL_1__8893_ (
);

FILL FILL_1__8473_ (
);

FILL FILL_1__8053_ (
);

FILL FILL_3__9340_ (
);

FILL FILL_0__13229_ (
);

FILL FILL_2__6396_ (
);

FILL FILL_1__9678_ (
);

FILL FILL_1__9258_ (
);

FILL FILL_3__12170_ (
);

FILL FILL_2__11583_ (
);

FILL FILL_2__11163_ (
);

FILL FILL_1__10996_ (
);

FILL FILL_1__10576_ (
);

FILL FILL_1__10156_ (
);

FILL FILL_0__7583_ (
);

FILL FILL_0__7163_ (
);

FILL FILL_3__10903_ (
);

FILL FILL_2__8542_ (
);

FILL FILL_0__10930_ (
);

FILL FILL_0__10510_ (
);

FILL FILL_2__12788_ (
);

FILL FILL_2__12368_ (
);

FILL FILL_0__8788_ (
);

FILL FILL_0__8368_ (
);

FILL FILL_3__6465_ (
);

INVX1 _10639_ (
    .A(_3902_),
    .Y(_3903_)
);

AND2X2 _10219_ (
    .A(_3495_),
    .B(_3494_),
    .Y(_3497_)
);

FILL FILL_1__12722_ (
);

FILL FILL_1__12302_ (
);

FILL FILL_2__9747_ (
);

FILL FILL_2__9327_ (
);

FILL FILL_0__11715_ (
);

FILL FILL_1__7744_ (
);

FILL FILL_1__7324_ (
);

FILL FILL254250x183750 (
);

INVX1 _6394_ (
    .A(_785_),
    .Y(_786_)
);

FILL FILL_3__8611_ (
);

OAI21X1 _10392_ (
    .A(_3262_),
    .B(_3507_),
    .C(_3661_),
    .Y(_3668_)
);

FILL FILL_1__8949_ (
);

FILL FILL_1__8529_ (
);

FILL FILL_3__11021_ (
);

FILL FILL_2__10854_ (
);

FILL FILL_2__10434_ (
);

FILL FILL_2__9080_ (
);

FILL FILL_2__10014_ (
);

OAI21X1 _7599_ (
    .A(_812_),
    .B(_1116_),
    .C(_822_),
    .Y(_1117_)
);

NOR2X1 _7179_ (
    .A(\u_fir_pe0.rYin [14]),
    .B(\u_fir_pe0.mul [14]),
    .Y(_763_)
);

FILL FILL_3__9816_ (
);

FILL FILL_0__6854_ (
);

DFFPOSX1 _8960_ (
    .D(_2384_[7]),
    .CLK(clk_bF$buf47),
    .Q(\Y[3] [7])
);

FILL FILL_0__6434_ (
);

OAI21X1 _8540_ (
    .A(_1898_),
    .B(_1902_),
    .C(_1907_),
    .Y(_1977_)
);

DFFPOSX1 _8120_ (
    .D(_1592_[4]),
    .CLK(clk_bF$buf43),
    .Q(\u_fir_pe1.mul [4])
);

DFFPOSX1 _11597_ (
    .D(_4775_[13]),
    .CLK(clk_bF$buf6),
    .Q(\Y[6] [13])
);

INVX1 _11177_ (
    .A(_4373_),
    .Y(_4374_)
);

FILL FILL_2__7813_ (
);

FILL FILL_3__12646_ (
);

FILL FILL_1__13260_ (
);

FILL FILL_0__12673_ (
);

FILL FILL_2__11219_ (
);

FILL FILL_0__12253_ (
);

FILL FILL_0__7639_ (
);

OAI21X1 _9745_ (
    .A(_3072_),
    .B(_3073_),
    .C(_3087_),
    .Y(_3088_)
);

INVX1 _9325_ (
    .A(_2679_),
    .Y(_2684_)
);

FILL FILL_1__8282_ (
);

FILL FILL_0__13038_ (
);

INVX1 _13323_ (
    .A(_6341_),
    .Y(_6346_)
);

FILL FILL_1__9487_ (
);

FILL FILL_1__9067_ (
);

FILL FILL_2__11392_ (
);

FILL FILL_1__10385_ (
);

FILL FILL_0__7392_ (
);

FILL FILL_2__8771_ (
);

FILL FILL_2__8351_ (
);

FILL FILL_2__12597_ (
);

FILL FILL_2__12177_ (
);

NAND3X1 _7811_ (
    .A(_1322_),
    .B(_1325_),
    .C(_1279_),
    .Y(_1326_)
);

FILL FILL_0__8597_ (
);

FILL FILL_3__6694_ (
);

FILL FILL_0__8177_ (
);

OAI22X1 _10868_ (
    .A(_4716_),
    .B(_4068_),
    .C(_4018_),
    .D(_4023_),
    .Y(_4069_)
);

NAND3X1 _10448_ (
    .A(_3717_),
    .B(_3722_),
    .C(_3721_),
    .Y(_3723_)
);

INVX1 _10028_ (
    .A(_3208_),
    .Y(_3309_)
);

FILL FILL_3__11917_ (
);

FILL FILL_1__12951_ (
);

FILL FILL_1__12531_ (
);

FILL FILL_1__12111_ (
);

FILL FILL_2__9976_ (
);

FILL FILL_2__9556_ (
);

FILL FILL_0__11944_ (
);

FILL FILL_2__9136_ (
);

FILL FILL_0__11524_ (
);

FILL FILL_0__11104_ (
);

FILL FILL_1__7973_ (
);

FILL FILL_1__7553_ (
);

FILL FILL_1__7133_ (
);

FILL FILL_3__7479_ (
);

FILL FILL_3__7059_ (
);

FILL FILL_1__13316_ (
);

FILL FILL_0__12729_ (
);

FILL FILL_0__12309_ (
);

FILL FILL_1__8758_ (
);

FILL FILL_3__11670_ (
);

FILL FILL_1__8338_ (
);

FILL FILL_3__11250_ (
);

FILL FILL_2__10663_ (
);

FILL FILL_2__10243_ (
);

FILL FILL_3__9205_ (
);

FILL FILL_0__6663_ (
);

FILL FILL_3__12875_ (
);

FILL FILL_2__7622_ (
);

FILL FILL_3__12035_ (
);

FILL FILL_2__11868_ (
);

FILL FILL_2__11448_ (
);

FILL FILL_2__11028_ (
);

FILL FILL_0__12062_ (
);

FILL FILL_0__7868_ (
);

NOR2X1 _9974_ (
    .A(_3209_),
    .B(_3246_),
    .Y(_3255_)
);

FILL FILL_0__7448_ (
);

AOI22X1 _9554_ (
    .A(\X[3]_5_bF$buf3 ),
    .B(gnd),
    .C(_2868_),
    .D(_2869_),
    .Y(_2909_)
);

FILL FILL_0__7028_ (
);

NAND3X1 _9134_ (
    .A(_2486_),
    .B(_2482_),
    .C(_2488_),
    .Y(_2495_)
);

FILL FILL_1__11802_ (
);

FILL FILL_2__8827_ (
);

FILL FILL_2__8407_ (
);

FILL FILL_0__13267_ (
);

NAND3X1 _13132_ (
    .A(_5956_),
    .B(_6029_),
    .C(_6135_),
    .Y(_6166_)
);

FILL FILL_1__6824_ (
);

FILL FILL_1__6404_ (
);

FILL FILL_1__9296_ (
);

FILL FILL_1__10194_ (
);

FILL FILL_1__7609_ (
);

FILL FILL_3__10521_ (
);

FILL FILL_2__8580_ (
);

FILL FILL_2__8160_ (
);

NAND3X1 _6679_ (
    .A(_222_),
    .B(_263_),
    .C(_268_),
    .Y(_278_)
);

AOI21X1 _7620_ (
    .A(_1133_),
    .B(_1137_),
    .C(_1119_),
    .Y(_1138_)
);

DFFPOSX1 _7200_ (
    .D(_790_[1]),
    .CLK(clk_bF$buf19),
    .Q(\Y[1] [1])
);

FILL FILL_1__11399_ (
);

NOR2X1 _10677_ (
    .A(_3939_),
    .B(_3940_),
    .Y(_3941_)
);

INVX1 _10257_ (
    .A(_3448_),
    .Y(_3535_)
);

FILL FILL_1__12760_ (
);

FILL FILL_3__11306_ (
);

FILL FILL_1__12340_ (
);

FILL FILL_2__9785_ (
);

FILL FILL_2__9365_ (
);

FILL FILL_0__11753_ (
);

FILL FILL_0__11333_ (
);

FILL FILL_0__6719_ (
);

NOR2X1 _8825_ (
    .A(_2249_),
    .B(_2250_),
    .Y(_2251_)
);

AOI21X1 _8405_ (
    .A(_1841_),
    .B(_1843_),
    .C(_1840_),
    .Y(_1844_)
);

FILL FILL_1__7782_ (
);

FILL FILL_1__7362_ (
);

FILL FILL_1__13125_ (
);

FILL FILL_0__12958_ (
);

OAI21X1 _12823_ (
    .A(_5848_),
    .B(_5852_),
    .C(_5855_),
    .Y(_5862_)
);

FILL FILL_0__12538_ (
);

FILL FILL_0__12118_ (
);

INVX1 _12403_ (
    .A(\u_fir_pe6.mul [10]),
    .Y(_5507_)
);

FILL FILL_1__8567_ (
);

FILL FILL_1__8147_ (
);

FILL FILL_2__10892_ (
);

FILL FILL_2__10472_ (
);

FILL FILL_2__10052_ (
);

FILL FILL_3__9434_ (
);

FILL FILL_0__6892_ (
);

FILL FILL_0__6472_ (
);

FILL FILL_2__7851_ (
);

FILL FILL_2__7431_ (
);

FILL FILL_3__12264_ (
);

FILL FILL_2__7011_ (
);

FILL FILL_2__11677_ (
);

FILL FILL_2__11257_ (
);

FILL FILL_0__12291_ (
);

FILL FILL_0__7677_ (
);

NOR2X1 _9783_ (
    .A(_3126_),
    .B(_3123_),
    .Y(_3127_)
);

FILL FILL_0__7257_ (
);

INVX1 _9363_ (
    .A(_2715_),
    .Y(_2721_)
);

FILL FILL_2__8636_ (
);

FILL FILL_2__8216_ (
);

FILL FILL_0__10604_ (
);

FILL FILL_3__13049_ (
);

DFFPOSX1 _13361_ (
    .D(\X[6] [7]),
    .CLK(clk_bF$buf37),
    .Q(\X[7] [7])
);

FILL FILL_0__13076_ (
);

FILL FILL_1__6633_ (
);

FILL FILL_2__13403_ (
);

FILL FILL_3__6559_ (
);

FILL FILL_1__12816_ (
);

FILL FILL_0__9823_ (
);

FILL FILL_3__7920_ (
);

FILL FILL_0__9403_ (
);

FILL FILL_0__11809_ (
);

FILL FILL254550x129750 (
);

FILL FILL_1__7838_ (
);

FILL FILL_1__7418_ (
);

INVX1 _6488_ (
    .A(vdd),
    .Y(_89_)
);

FILL FILL_3__8705_ (
);

NAND3X1 _10486_ (
    .A(_3752_),
    .B(_3759_),
    .C(_3758_),
    .Y(_3760_)
);

AND2X2 _10066_ (
    .A(gnd),
    .B(\X[4] [4]),
    .Y(_3346_)
);

FILL FILL_2__6702_ (
);

FILL FILL_3__11115_ (
);

FILL FILL_2__10948_ (
);

FILL FILL_0__11982_ (
);

FILL FILL_2__9594_ (
);

FILL FILL_2__10528_ (
);

FILL FILL_2__9174_ (
);

FILL FILL_0__11562_ (
);

FILL FILL_2__10108_ (
);

FILL FILL_0__11142_ (
);

FILL FILL_0__6948_ (
);

FILL FILL_0__6528_ (
);

OAI22X1 _8634_ (
    .A(_1925_),
    .B(_2006_),
    .C(_2068_),
    .D(_2069_),
    .Y(_2070_)
);

INVX1 _8214_ (
    .A(_1639_),
    .Y(_1656_)
);

FILL FILL_1__7591_ (
);

FILL FILL_1__7171_ (
);

FILL FILL_2__7907_ (
);

FILL FILL_0__12767_ (
);

NAND3X1 _12632_ (
    .A(vdd),
    .B(\X[6] [2]),
    .C(_5672_),
    .Y(_5673_)
);

FILL FILL_0__12347_ (
);

NAND2X1 _12212_ (
    .A(_5321_),
    .B(_5318_),
    .Y(_5327_)
);

DFFPOSX1 _9839_ (
    .D(_3181_[9]),
    .CLK(clk_bF$buf17),
    .Q(\Y[4] [9])
);

OAI21X1 _9419_ (
    .A(_2706_),
    .B(_2775_),
    .C(_2745_),
    .Y(_2776_)
);

FILL FILL_1__8796_ (
);

FILL FILL_1__8376_ (
);

FILL FILL_2__10281_ (
);

FILL FILL_3__9663_ (
);

BUFX2 _13417_ (
    .A(_6377_[9]),
    .Y(Yout[9])
);

FILL FILL_2__7660_ (
);

FILL FILL_2__11486_ (
);

FILL FILL_2__11066_ (
);

FILL FILL_1__10899_ (
);

INVX1 _6700_ (
    .A(_282_),
    .Y(_298_)
);

FILL FILL_1__10479_ (
);

FILL FILL_1__10059_ (
);

FILL FILL_0__7486_ (
);

NAND2X1 _9592_ (
    .A(_2945_),
    .B(_2946_),
    .Y(_3187_[11])
);

FILL FILL_0__7066_ (
);

AND2X2 _9172_ (
    .A(\X[3] [2]),
    .B(gnd),
    .Y(_2532_)
);

FILL FILL_1__11840_ (
);

FILL FILL_1__11420_ (
);

FILL FILL_1__11000_ (
);

FILL FILL_2__8865_ (
);

FILL FILL_2__8445_ (
);

FILL FILL_0__10833_ (
);

FILL FILL_3__13278_ (
);

FILL FILL_0__10413_ (
);

FILL FILL_2__8025_ (
);

INVX1 _13170_ (
    .A(_6161_),
    .Y(_6202_)
);

NAND2X1 _7905_ (
    .A(_1415_),
    .B(_1414_),
    .Y(_1417_)
);

FILL FILL_1__6862_ (
);

FILL FILL_1__6442_ (
);

FILL FILL_2__13212_ (
);

FILL FILL_3__6788_ (
);

FILL FILL_1__12625_ (
);

FILL FILL_1__12205_ (
);

FILL FILL_0__9632_ (
);

FILL FILL_0__9212_ (
);

NAND2X1 _11903_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5022_)
);

FILL FILL_1__7647_ (
);

FILL FILL_3__8934_ (
);

AOI21X1 _10295_ (
    .A(_3537_),
    .B(_3538_),
    .C(_3505_),
    .Y(_3572_)
);

FILL FILL_2__6931_ (
);

FILL FILL_3__11764_ (
);

FILL FILL_2__6511_ (
);

FILL FILL_3__11344_ (
);

FILL FILL_0__11791_ (
);

FILL FILL_2__10337_ (
);

FILL FILL_0__11371_ (
);

FILL FILL_0__6757_ (
);

NOR2X1 _8863_ (
    .A(_2284_),
    .B(_2285_),
    .Y(_2286_)
);

NAND3X1 _8443_ (
    .A(_1782_),
    .B(_1880_),
    .C(_1881_),
    .Y(_1882_)
);

OAI21X1 _8023_ (
    .A(_1523_),
    .B(_1524_),
    .C(_1519_),
    .Y(_1527_)
);

FILL FILL_3__12969_ (
);

FILL FILL_2__7716_ (
);

FILL FILL_3__12549_ (
);

FILL FILL_3__12129_ (
);

FILL FILL_1__13163_ (
);

FILL FILL_0__12996_ (
);

OAI21X1 _12861_ (
    .A(_5594_),
    .B(_5898_),
    .C(_5604_),
    .Y(_5899_)
);

FILL FILL_0__12576_ (
);

FILL FILL_0__12156_ (
);

NOR2X1 _12441_ (
    .A(\u_fir_pe6.rYin [14]),
    .B(\u_fir_pe6.mul [14]),
    .Y(_5545_)
);

OAI21X1 _12021_ (
    .A(_5138_),
    .B(_5134_),
    .C(_5085_),
    .Y(_5139_)
);

FILL FILL_2__12903_ (
);

OAI21X1 _9648_ (
    .A(_2982_),
    .B(_2977_),
    .C(_3000_),
    .Y(_3001_)
);

INVX1 _9228_ (
    .A(_2497_),
    .Y(_2588_)
);

FILL FILL_1__8185_ (
);

FILL FILL253950x205350 (
);

FILL FILL_0__8903_ (
);

FILL FILL_2__10090_ (
);

FILL FILL_3__9892_ (
);

FILL FILL_3__9052_ (
);

AND2X2 _13226_ (
    .A(_6250_),
    .B(_6249_),
    .Y(_6369_[5])
);

FILL FILL_1__6918_ (
);

FILL FILL_2__11295_ (
);

FILL FILL_1__10288_ (
);

FILL FILL_0__7295_ (
);

FILL FILL_3__10615_ (
);

FILL FILL_2__8674_ (
);

FILL FILL_2__8254_ (
);

FILL FILL_0__10642_ (
);

FILL FILL_3__13087_ (
);

FILL FILL_0__10222_ (
);

INVX1 _7714_ (
    .A(_1223_),
    .Y(_1231_)
);

FILL FILL_1__6671_ (
);

FILL FILL_2__13021_ (
);

FILL FILL_1__12854_ (
);

FILL FILL_1__12434_ (
);

FILL FILL_1__12014_ (
);

FILL FILL_2__9459_ (
);

FILL FILL_0__9441_ (
);

FILL FILL_0__11847_ (
);

FILL FILL_2__9039_ (
);

FILL FILL_0__9021_ (
);

NAND3X1 _11712_ (
    .A(_4810_),
    .B(_4833_),
    .C(_4832_),
    .Y(_4834_)
);

FILL FILL_0__11427_ (
);

FILL FILL_0__11007_ (
);

AND2X2 _8919_ (
    .A(_2342_),
    .B(_2341_),
    .Y(_2384_[12])
);

FILL FILL_1__7876_ (
);

FILL FILL_1__7456_ (
);

FILL FILL_1__7036_ (
);

FILL FILL_1__13219_ (
);

FILL FILL_3__8743_ (
);

AOI21X1 _12917_ (
    .A(_5868_),
    .B(_5783_),
    .C(_5954_),
    .Y(_5955_)
);

FILL FILL_3__8323_ (
);

FILL FILL_3__11993_ (
);

FILL FILL_2__6740_ (
);

FILL FILL_3__11573_ (
);

FILL FILL254250x115350 (
);

FILL FILL_2__10986_ (
);

FILL FILL_2__10566_ (
);

FILL FILL_2__10146_ (
);

FILL FILL_0__11180_ (
);

FILL FILL_1__9602_ (
);

FILL FILL_3__9948_ (
);

FILL FILL_3__9528_ (
);

FILL FILL_3__9108_ (
);

FILL FILL_0__6986_ (
);

FILL FILL_0__6566_ (
);

NOR2X1 _8672_ (
    .A(_2087_),
    .B(_2092_),
    .Y(_2107_)
);

AOI22X1 _8252_ (
    .A(gnd),
    .B(\X[2] [4]),
    .C(_1682_),
    .D(_1684_),
    .Y(_1693_)
);

FILL FILL_1__10920_ (
);

FILL FILL_1__10500_ (
);

FILL FILL_2__7945_ (
);

FILL FILL253950x54150 (
);

FILL FILL_2__7525_ (
);

FILL FILL_3__12358_ (
);

FILL FILL_2__7105_ (
);

AND2X2 _12670_ (
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5710_)
);

FILL FILL_0__12385_ (
);

OAI21X1 _12250_ (
    .A(_5361_),
    .B(_5363_),
    .C(_5342_),
    .Y(_5364_)
);

FILL FILL_2__12712_ (
);

DFFPOSX1 _9877_ (
    .D(_3187_[7]),
    .CLK(clk_bF$buf42),
    .Q(\u_fir_pe3.mul [7])
);

NAND3X1 _9457_ (
    .A(_2806_),
    .B(_2813_),
    .C(_2788_),
    .Y(_2814_)
);

NAND3X1 _9037_ (
    .A(_3131_),
    .B(_2399_),
    .C(_2397_),
    .Y(_2400_)
);

FILL FILL_1__11705_ (
);

FILL FILL_0__8712_ (
);

FILL FILL_3__9281_ (
);

NAND3X1 _13035_ (
    .A(_6066_),
    .B(_6070_),
    .C(_6040_),
    .Y(_6071_)
);

FILL FILL_1__6727_ (
);

FILL FILL_1__9199_ (
);

FILL FILL_0__9917_ (
);

FILL FILL_1__10097_ (
);

FILL FILL_3__10844_ (
);

FILL FILL_3__10004_ (
);

FILL FILL_2__8483_ (
);

FILL FILL_0__10871_ (
);

FILL FILL_0__10451_ (
);

FILL FILL_2__8063_ (
);

FILL FILL_0__10031_ (
);

NAND2X1 _7943_ (
    .A(_1449_),
    .B(_1444_),
    .Y(_1450_)
);

AOI21X1 _7523_ (
    .A(_1041_),
    .B(_1040_),
    .C(_1037_),
    .Y(_1042_)
);

INVX1 _7103_ (
    .A(_680_),
    .Y(_686_)
);

FILL FILL_1__6480_ (
);

FILL FILL_2__13250_ (
);

FILL FILL_1__12663_ (
);

FILL FILL_1__12243_ (
);

FILL FILL_0__9670_ (
);

FILL FILL_2__9688_ (
);

FILL FILL_0__9250_ (
);

FILL FILL_2__9268_ (
);

NAND3X1 _11941_ (
    .A(_5004_),
    .B(_5045_),
    .C(_5050_),
    .Y(_5060_)
);

FILL FILL_0__11656_ (
);

AOI21X1 _11521_ (
    .A(_4699_),
    .B(_4677_),
    .C(_4697_),
    .Y(_4704_)
);

FILL FILL_0__11236_ (
);

NAND3X1 _11101_ (
    .A(_4296_),
    .B(_4298_),
    .C(_4297_),
    .Y(_4299_)
);

NOR2X1 _8728_ (
    .A(_2161_),
    .B(_2160_),
    .Y(_2162_)
);

AOI22X1 _8308_ (
    .A(vdd),
    .B(\X[2] [2]),
    .C(gnd),
    .D(\X[2] [3]),
    .Y(_1748_)
);

FILL FILL_1__7685_ (
);

FILL FILL_1__7265_ (
);

FILL FILL_1__13028_ (
);

FILL FILL_3__8552_ (
);

NAND3X1 _12726_ (
    .A(_5763_),
    .B(_5764_),
    .C(_5765_),
    .Y(_5766_)
);

INVX1 _12306_ (
    .A(\u_fir_pe6.mul [1]),
    .Y(_5415_)
);

FILL FILL_2__10795_ (
);

FILL FILL_2__10375_ (
);

FILL FILL_1__9411_ (
);

FILL FILL_3__9757_ (
);

FILL FILL_0__6795_ (
);

NAND2X1 _8481_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf0 ),
    .Y(_1919_)
);

INVX1 _8061_ (
    .A(_1559_),
    .Y(_1564_)
);

FILL FILL_2__7754_ (
);

FILL FILL_3__12587_ (
);

FILL FILL_2__7334_ (
);

FILL FILL_0__12194_ (
);

FILL FILL_2__12941_ (
);

FILL FILL_2__12521_ (
);

FILL FILL_2__12101_ (
);

OAI21X1 _9686_ (
    .A(_3032_),
    .B(_3033_),
    .C(_3031_),
    .Y(_3034_)
);

OAI21X1 _9266_ (
    .A(_2406_),
    .B(_2624_),
    .C(_2619_),
    .Y(_2625_)
);

FILL FILL_1__11934_ (
);

FILL FILL_1__11514_ (
);

FILL FILL_0__8941_ (
);

FILL FILL_2__8539_ (
);

FILL FILL_0__8521_ (
);

FILL FILL_0__10927_ (
);

FILL FILL_0__10507_ (
);

FILL FILL_0__13399_ (
);

INVX1 _13264_ (
    .A(_6271_),
    .Y(_6287_)
);

FILL FILL_2__9900_ (
);

FILL FILL_1__6956_ (
);

FILL FILL_1__6536_ (
);

FILL FILL_2__13306_ (
);

FILL FILL_1__12719_ (
);

FILL FILL_0__9726_ (
);

FILL FILL_0__9306_ (
);

FILL FILL_3__7403_ (
);

FILL FILL_3__10233_ (
);

FILL FILL_2__8292_ (
);

FILL FILL_0__10680_ (
);

FILL FILL_0__10260_ (
);

NOR2X1 _7752_ (
    .A(_1203_),
    .B(_1200_),
    .Y(_1268_)
);

OR2X2 _7332_ (
    .A(_853_),
    .B(_852_),
    .Y(_854_)
);

AND2X2 _10389_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3665_)
);

FILL FILL_3__11858_ (
);

FILL FILL_2__6605_ (
);

FILL FILL_1__12892_ (
);

FILL FILL_3__11438_ (
);

FILL FILL_3__11018_ (
);

FILL FILL_1__12052_ (
);

FILL FILL_0__11885_ (
);

FILL FILL_2__9497_ (
);

FILL FILL_2__9077_ (
);

INVX1 _11750_ (
    .A(vdd),
    .Y(_4871_)
);

FILL FILL_0__11465_ (
);

FILL FILL_0__11045_ (
);

NAND2X1 _11330_ (
    .A(_4517_),
    .B(_4520_),
    .Y(_4525_)
);

DFFPOSX1 _8957_ (
    .D(_2384_[4]),
    .CLK(clk_bF$buf47),
    .Q(\Y[3] [4])
);

AOI21X1 _8537_ (
    .A(_1891_),
    .B(_1961_),
    .C(_1973_),
    .Y(_1974_)
);

DFFPOSX1 _8117_ (
    .D(_1589_[1]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.mul [1])
);

FILL FILL_1__7494_ (
);

FILL FILL_1__7074_ (
);

FILL FILL_1__13257_ (
);

OAI21X1 _12955_ (
    .A(_5912_),
    .B(_5991_),
    .C(_5990_),
    .Y(_5992_)
);

FILL FILL_3__8361_ (
);

INVX1 _12535_ (
    .A(_6366_),
    .Y(_6367_)
);

AND2X2 _12115_ (
    .A(_5231_),
    .B(_5224_),
    .Y(_5232_)
);

FILL FILL_1__8699_ (
);

FILL FILL_1__8279_ (
);

FILL FILL_3__11191_ (
);

FILL FILL_2__10184_ (
);

FILL FILL_1__9640_ (
);

FILL FILL_1__9220_ (
);

FILL FILL_3__9146_ (
);

NAND2X1 _8290_ (
    .A(_1729_),
    .B(_1728_),
    .Y(_1730_)
);

FILL FILL_2__7983_ (
);

FILL FILL_2__7563_ (
);

FILL FILL_2__7143_ (
);

FILL FILL_2__11389_ (
);

NAND2X1 _6603_ (
    .A(_202_),
    .B(_194_),
    .Y(_203_)
);

FILL FILL_2__12750_ (
);

FILL FILL_2__12330_ (
);

FILL FILL_0__7389_ (
);

OAI21X1 _9495_ (
    .A(_2777_),
    .B(_2781_),
    .C(_2779_),
    .Y(_2851_)
);

INVX1 _9075_ (
    .A(_2423_),
    .Y(_2437_)
);

FILL FILL_1__11743_ (
);

FILL FILL_1__11323_ (
);

FILL FILL_2__8768_ (
);

FILL FILL_0__8750_ (
);

FILL FILL_0__8330_ (
);

FILL FILL_2__8348_ (
);

FILL FILL_0__10316_ (
);

NOR2X1 _10601_ (
    .A(_3864_),
    .B(_3863_),
    .Y(_3865_)
);

NAND3X1 _13073_ (
    .A(_6104_),
    .B(_6107_),
    .C(_6061_),
    .Y(_6108_)
);

NAND2X1 _7808_ (
    .A(gnd),
    .B(\X[1] [7]),
    .Y(_1323_)
);

FILL FILL_1__6765_ (
);

FILL FILL_2__13115_ (
);

FILL FILL_1__12948_ (
);

FILL FILL_1__12528_ (
);

FILL FILL_1__12108_ (
);

FILL FILL_0__9955_ (
);

FILL FILL_0__9535_ (
);

FILL FILL_3__7632_ (
);

FILL FILL_0__9115_ (
);

INVX2 _11806_ (
    .A(\X[7] [6]),
    .Y(_4926_)
);

FILL FILL_3__10462_ (
);

FILL FILL_1__8911_ (
);

FILL FILL_3__8417_ (
);

NOR2X1 _7981_ (
    .A(_1481_),
    .B(_1480_),
    .Y(_1484_)
);

OAI21X1 _7561_ (
    .A(_1066_),
    .B(_1070_),
    .C(_1073_),
    .Y(_1080_)
);

INVX1 _7141_ (
    .A(\u_fir_pe0.mul [10]),
    .Y(_725_)
);

AND2X2 _10198_ (
    .A(_3473_),
    .B(_3476_),
    .Y(_3477_)
);

FILL FILL_2__6834_ (
);

FILL FILL_2__6414_ (
);

FILL FILL_1__12281_ (
);

FILL FILL_0__11694_ (
);

FILL FILL_0__11274_ (
);

NAND3X1 _8766_ (
    .A(_2172_),
    .B(_2174_),
    .C(_2198_),
    .Y(_2199_)
);

NAND3X1 _8346_ (
    .A(_1730_),
    .B(_1779_),
    .C(_1780_),
    .Y(_1786_)
);

FILL FILL_0__7601_ (
);

FILL FILL_2__7619_ (
);

FILL FILL_1__13066_ (
);

FILL FILL_0__12899_ (
);

FILL FILL_3__8590_ (
);

OAI21X1 _12764_ (
    .A(_5752_),
    .B(_5802_),
    .C(_5746_),
    .Y(_5803_)
);

FILL FILL_3__8170_ (
);

FILL FILL_0__12059_ (
);

NOR2X1 _12344_ (
    .A(_5447_),
    .B(_5448_),
    .Y(_5449_)
);

FILL FILL_2__12806_ (
);

FILL FILL_0__13000_ (
);

FILL FILL_0__8806_ (
);

FILL FILL_3__9375_ (
);

OR2X2 _13129_ (
    .A(_6162_),
    .B(_6139_),
    .Y(_6163_)
);

FILL FILL_2__7792_ (
);

FILL FILL_2__7372_ (
);

FILL FILL_2__11198_ (
);

AOI21X1 _6832_ (
    .A(_415_),
    .B(_422_),
    .C(_397_),
    .Y(_429_)
);

INVX2 _6412_ (
    .A(Xin[3]),
    .Y(_15_)
);

FILL FILL_0__7198_ (
);

FILL FILL_3__10938_ (
);

FILL FILL_1__11972_ (
);

FILL FILL_1__11552_ (
);

FILL FILL_1__11132_ (
);

FILL FILL_2__8577_ (
);

FILL FILL_0__10965_ (
);

FILL FILL_2__8157_ (
);

FILL FILL_0__10545_ (
);

NAND2X1 _10830_ (
    .A(_4029_),
    .B(_4025_),
    .Y(_4032_)
);

AOI21X1 _10410_ (
    .A(_3583_),
    .B(_3613_),
    .C(_3616_),
    .Y(_3686_)
);

FILL FILL_0__10125_ (
);

NAND3X1 _7617_ (
    .A(_1127_),
    .B(_1131_),
    .C(_1129_),
    .Y(_1135_)
);

FILL FILL_1__6994_ (
);

FILL FILL_1__6574_ (
);

FILL FILL_1__12757_ (
);

FILL FILL_1__12337_ (
);

FILL FILL_0__9764_ (
);

FILL FILL_3__7861_ (
);

FILL FILL_0__9344_ (
);

DFFPOSX1 _11615_ (
    .D(\Y[5] [7]),
    .CLK(clk_bF$buf18),
    .Q(\u_fir_pe5.rYin [7])
);

FILL FILL_3__7021_ (
);

FILL FILL_1__7779_ (
);

FILL FILL_1__7359_ (
);

FILL FILL_1__8720_ (
);

FILL FILL_1__8300_ (
);

FILL FILL_3__8646_ (
);

OAI21X1 _7790_ (
    .A(_1305_),
    .B(_1173_),
    .C(_1255_),
    .Y(_1306_)
);

NAND3X1 _7370_ (
    .A(vdd),
    .B(\X[1] [2]),
    .C(_890_),
    .Y(_891_)
);

FILL FILL_2__6643_ (
);

FILL FILL_3__11056_ (
);

FILL FILL_1__12090_ (
);

FILL FILL_2__10889_ (
);

FILL FILL_2__10469_ (
);

FILL FILL_2__10049_ (
);

FILL FILL_0__11083_ (
);

FILL FILL_1__9925_ (
);

FILL FILL_1__9505_ (
);

FILL FILL_2__11830_ (
);

FILL FILL_0__6889_ (
);

FILL FILL_2__11410_ (
);

DFFPOSX1 _8995_ (
    .D(_2387_[2]),
    .CLK(clk_bF$buf53),
    .Q(\u_fir_pe2.mul [2])
);

FILL FILL_0__6469_ (
);

OAI21X1 _8575_ (
    .A(_2011_),
    .B(_1913_),
    .C(_1726_),
    .Y(_2012_)
);

AOI22X1 _8155_ (
    .A(vdd),
    .B(\X[2] [0]),
    .C(gnd),
    .D(\X[2] [1]),
    .Y(_1598_)
);

FILL FILL_1__10823_ (
);

FILL FILL_1__10403_ (
);

FILL FILL_2__7848_ (
);

FILL FILL_0__7830_ (
);

FILL FILL_0__7410_ (
);

FILL FILL_2__7428_ (
);

FILL FILL_2__7008_ (
);

FILL FILL_1__13295_ (
);

OR2X2 _12993_ (
    .A(_5959_),
    .B(_6029_),
    .Y(_6030_)
);

AND2X2 _12573_ (
    .A(vdd),
    .B(\X[6] [2]),
    .Y(_5615_)
);

FILL FILL_0__12288_ (
);

NAND3X1 _12153_ (
    .A(_5252_),
    .B(_5268_),
    .C(_5266_),
    .Y(_5269_)
);

FILL FILL_3__13202_ (
);

FILL FILL_2__12615_ (
);

FILL FILL_0__8615_ (
);

FILL FILL_3__6712_ (
);

DFFPOSX1 _13358_ (
    .D(\X[6] [4]),
    .CLK(clk_bF$buf2),
    .Q(\X[7] [4])
);

FILL FILL_2__7181_ (
);

NAND2X1 _6641_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_240_)
);

FILL FILL_1__11781_ (
);

FILL FILL_3__10327_ (
);

FILL FILL_1__11361_ (
);

FILL FILL_2__8386_ (
);

FILL FILL_0__10774_ (
);

FILL FILL_0__10354_ (
);

INVX1 _7846_ (
    .A(_1359_),
    .Y(_1360_)
);

NAND2X1 _7426_ (
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_946_)
);

NAND2X1 _7006_ (
    .A(_598_),
    .B(_572_),
    .Y(_599_)
);

FILL FILL_1__6383_ (
);

FILL FILL_2__13153_ (
);

FILL FILL_1__12986_ (
);

FILL FILL_1__12566_ (
);

FILL FILL_1__12146_ (
);

FILL FILL_0__9993_ (
);

FILL FILL_0__9573_ (
);

FILL FILL_0__11979_ (
);

FILL FILL_0__9153_ (
);

OAI21X1 _11844_ (
    .A(_4962_),
    .B(_4963_),
    .C(_4961_),
    .Y(_4964_)
);

FILL FILL_0__11559_ (
);

OAI21X1 _11424_ (
    .A(_4552_),
    .B(_4602_),
    .C(_4580_),
    .Y(_4615_)
);

FILL FILL_0__11139_ (
);

NAND3X1 _11004_ (
    .A(_4196_),
    .B(_4202_),
    .C(_4201_),
    .Y(_4203_)
);

FILL FILL_0__12920_ (
);

FILL FILL_1__7588_ (
);

FILL FILL_1__7168_ (
);

FILL FILL_3__10080_ (
);

NAND3X1 _12629_ (
    .A(_5665_),
    .B(_5669_),
    .C(_5667_),
    .Y(_5670_)
);

NAND3X1 _12209_ (
    .A(_5297_),
    .B(_5323_),
    .C(_5319_),
    .Y(_5324_)
);

FILL FILL_2__6872_ (
);

FILL FILL_2__6452_ (
);

FILL FILL_3__11285_ (
);

FILL FILL_2__10698_ (
);

FILL FILL_2__10278_ (
);

FILL FILL_1__9734_ (
);

FILL FILL_1__9314_ (
);

FILL FILL_0__6698_ (
);

NAND2X1 _8384_ (
    .A(_1821_),
    .B(_1822_),
    .Y(_1823_)
);

FILL FILL_1__10632_ (
);

FILL FILL_1__10212_ (
);

FILL FILL253650x126150 (
);

FILL FILL_2__7657_ (
);

FILL FILL_0__12097_ (
);

OAI21X1 _12382_ (
    .A(_5474_),
    .B(_5475_),
    .C(_5485_),
    .Y(_5486_)
);

FILL FILL_2__12844_ (
);

FILL FILL_2__12424_ (
);

FILL FILL_2__12004_ (
);

INVX1 _9589_ (
    .A(_2943_),
    .Y(_2944_)
);

OAI21X1 _9169_ (
    .A(_2493_),
    .B(_2528_),
    .C(_2487_),
    .Y(_2529_)
);

FILL FILL_1__11837_ (
);

FILL FILL_1__11417_ (
);

FILL FILL_0__8844_ (
);

FILL FILL_3__6941_ (
);

FILL FILL_0__8424_ (
);

FILL FILL_0__8004_ (
);

NAND2X1 _13167_ (
    .A(_6197_),
    .B(_6196_),
    .Y(_6199_)
);

FILL FILL_2__9803_ (
);

FILL FILL_1__6859_ (
);

FILL FILL_1__6439_ (
);

FILL FILL_2__13209_ (
);

FILL FILL_1__7800_ (
);

FILL FILL_0__9629_ (
);

FILL FILL_3__7726_ (
);

FILL FILL_0__9209_ (
);

OAI22X1 _6870_ (
    .A(_15_),
    .B(_462_),
    .C(_463_),
    .D(_465_),
    .Y(_466_)
);

NAND3X1 _6450_ (
    .A(_28_),
    .B(_51_),
    .C(_50_),
    .Y(_52_)
);

FILL FILL_3__10556_ (
);

FILL FILL_1__11170_ (
);

FILL FILL_2__8195_ (
);

FILL FILL_0__10583_ (
);

FILL FILL_0__10163_ (
);

FILL FILL_2__10910_ (
);

AOI21X1 _7655_ (
    .A(_1086_),
    .B(_1001_),
    .C(_1172_),
    .Y(_1173_)
);

DFFPOSX1 _7235_ (
    .D(Yin[12]),
    .CLK(clk_bF$buf16),
    .Q(\u_fir_pe0.rYin [12])
);

FILL FILL_2__6928_ (
);

FILL FILL_0__6910_ (
);

FILL FILL_2__6508_ (
);

FILL FILL_1__12795_ (
);

FILL FILL_1__12375_ (
);

FILL FILL_0__9382_ (
);

FILL FILL_0__11788_ (
);

NOR2X1 _11653_ (
    .A(_5562_),
    .B(_5542_),
    .Y(_5565_)
);

FILL FILL_0__11368_ (
);

OAI21X1 _11233_ (
    .A(_4420_),
    .B(_4419_),
    .C(_4370_),
    .Y(_4430_)
);

FILL FILL_3__12702_ (
);

FILL FILL_1__7397_ (
);

NOR2X1 _9801_ (
    .A(\u_fir_pe3.rYin [13]),
    .B(\u_fir_pe3.mul [13]),
    .Y(_3145_)
);

FILL FILL_3__8684_ (
);

OAI21X1 _12858_ (
    .A(_5817_),
    .B(_5895_),
    .C(_5839_),
    .Y(_5896_)
);

FILL FILL_3__8264_ (
);

INVX1 _12438_ (
    .A(\u_fir_pe6.rYin [14]),
    .Y(_5541_)
);

NAND3X1 _12018_ (
    .A(_5131_),
    .B(_5132_),
    .C(_5099_),
    .Y(_5136_)
);

FILL FILL_2__6681_ (
);

FILL FILL_2__10087_ (
);

FILL FILL_1__9963_ (
);

FILL FILL_1__9543_ (
);

FILL FILL_1__9123_ (
);

FILL FILL_3__9889_ (
);

FILL FILL_3__9469_ (
);

FILL FILL_3__9049_ (
);

NAND3X1 _8193_ (
    .A(gnd),
    .B(\X[2] [2]),
    .C(_1625_),
    .Y(_1635_)
);

FILL FILL_1__10861_ (
);

FILL FILL_1__10441_ (
);

FILL FILL_1__10021_ (
);

FILL FILL_2__7886_ (
);

FILL FILL_2__7466_ (
);

FILL FILL_3__12299_ (
);

FILL FILL_2__7046_ (
);

NAND2X1 _12191_ (
    .A(_5301_),
    .B(_5305_),
    .Y(_5306_)
);

NAND2X1 _6926_ (
    .A(gnd),
    .B(_474_),
    .Y(_521_)
);

AOI21X1 _6506_ (
    .A(_28_),
    .B(_48_),
    .C(_62_),
    .Y(_107_)
);

FILL FILL_2__12653_ (
);

FILL FILL_2__12233_ (
);

OAI21X1 _9398_ (
    .A(_2747_),
    .B(_2743_),
    .C(_2750_),
    .Y(_2756_)
);

FILL FILL_1__11646_ (
);

FILL FILL_1__11226_ (
);

FILL FILL_0__8653_ (
);

FILL FILL_0__8233_ (
);

FILL FILL_0__10639_ (
);

NAND2X1 _10924_ (
    .A(\X[5] [1]),
    .B(gnd),
    .Y(_4124_)
);

NOR2X1 _10504_ (
    .A(_3777_),
    .B(_3776_),
    .Y(_3778_)
);

FILL FILL_0__10219_ (
);

BUFX2 _13396_ (
    .A(_6376_[2]),
    .Y(Xout[2])
);

FILL FILL_2__9612_ (
);

FILL FILL_1__6668_ (
);

FILL FILL_2__13018_ (
);

FILL FILL_3__7955_ (
);

FILL FILL_0__9438_ (
);

FILL FILL_0__9018_ (
);

NAND3X1 _11709_ (
    .A(_4811_),
    .B(_4827_),
    .C(_4830_),
    .Y(_4831_)
);

FILL FILL_3__7115_ (
);

FILL FILL_3__10785_ (
);

FILL FILL_0__10392_ (
);

FILL FILL_1__8814_ (
);

OR2X2 _7884_ (
    .A(_1369_),
    .B(_1395_),
    .Y(_1397_)
);

NAND3X1 _7464_ (
    .A(_981_),
    .B(_982_),
    .C(_983_),
    .Y(_984_)
);

INVX1 _7044_ (
    .A(\u_fir_pe0.mul [1]),
    .Y(_633_)
);

FILL FILL_2__13191_ (
);

FILL FILL_2__6737_ (
);

FILL FILL_1__12184_ (
);

FILL FILL_0__9191_ (
);

AOI21X1 _11882_ (
    .A(_4929_),
    .B(_4925_),
    .C(_4994_),
    .Y(_5001_)
);

OR2X2 _11462_ (
    .A(_4646_),
    .B(_4644_),
    .Y(_4648_)
);

FILL FILL_0__11177_ (
);

OAI21X1 _11042_ (
    .A(_4233_),
    .B(_4240_),
    .C(_4225_),
    .Y(_4241_)
);

FILL FILL_3__12931_ (
);

FILL FILL_2__11924_ (
);

FILL FILL_2__11504_ (
);

NOR2X1 _8669_ (
    .A(_2101_),
    .B(_2104_),
    .Y(_2390_[10])
);

NAND3X1 _8249_ (
    .A(_1678_),
    .B(_1689_),
    .C(_1685_),
    .Y(_1690_)
);

FILL FILL_1__10917_ (
);

FILL FILL_0__7924_ (
);

FILL FILL_0__7504_ (
);

NOR2X1 _9610_ (
    .A(_2956_),
    .B(_2960_),
    .Y(_2964_)
);

INVX1 _12667_ (
    .A(_5704_),
    .Y(_5708_)
);

FILL FILL_3__8073_ (
);

AOI21X1 _12247_ (
    .A(_5359_),
    .B(_5360_),
    .C(_5343_),
    .Y(_5361_)
);

FILL FILL_2__12709_ (
);

FILL FILL_0__13323_ (
);

FILL FILL_2__6490_ (
);

FILL FILL_0__8709_ (
);

FILL FILL_1__9772_ (
);

FILL FILL_1__9352_ (
);

FILL FILL_3__9698_ (
);

FILL FILL_1__10670_ (
);

FILL FILL_1__10250_ (
);

FILL FILL_2__7695_ (
);

FILL FILL_2__7275_ (
);

NAND2X1 _6735_ (
    .A(vdd),
    .B(Xin[6]),
    .Y(_333_)
);

FILL FILL_2__12882_ (
);

FILL FILL_2__12042_ (
);

FILL FILL_1__11875_ (
);

FILL FILL_1__11455_ (
);

FILL FILL_1__11035_ (
);

FILL FILL_0__8882_ (
);

FILL FILL_0__8462_ (
);

FILL FILL_0__10868_ (
);

FILL FILL_0__10448_ (
);

DFFPOSX1 _10733_ (
    .D(\Y[4] [2]),
    .CLK(clk_bF$buf55),
    .Q(\u_fir_pe4.rYin [2])
);

FILL FILL_0__8042_ (
);

AOI22X1 _10313_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf2 ),
    .C(gnd),
    .D(\X[4] [6]),
    .Y(_3590_)
);

FILL FILL_0__10028_ (
);

FILL FILL_2__9421_ (
);

FILL FILL_1__6897_ (
);

FILL FILL_1__6477_ (
);

FILL FILL_2__13247_ (
);

FILL FILL_3_CLKBUF1_insert30 (
);

FILL FILL_3_CLKBUF1_insert32 (
);

FILL FILL_3_CLKBUF1_insert34 (
);

FILL FILL_3_CLKBUF1_insert36 (
);

FILL FILL_3_CLKBUF1_insert37 (
);

FILL FILL254250x54150 (
);

FILL FILL_3_CLKBUF1_insert39 (
);

FILL FILL_0__9667_ (
);

FILL FILL_0__9247_ (
);

INVX1 _11938_ (
    .A(_4959_),
    .Y(_5057_)
);

FILL FILL_3__7344_ (
);

OAI21X1 _11518_ (
    .A(_4697_),
    .B(_4698_),
    .C(_4696_),
    .Y(_4702_)
);

FILL FILL_3__10594_ (
);

FILL FILL_3__10174_ (
);

FILL FILL_1__8623_ (
);

FILL FILL_1__8203_ (
);

OAI21X1 _7693_ (
    .A(_1130_),
    .B(_1209_),
    .C(_1208_),
    .Y(_1210_)
);

INVX1 _7273_ (
    .A(_1584_),
    .Y(_1585_)
);

FILL FILL_2__6966_ (
);

FILL FILL_3__11799_ (
);

FILL FILL_2__6546_ (
);

FILL FILL_3__11379_ (
);

NAND2X1 _11691_ (
    .A(gnd),
    .B(\X[7] [1]),
    .Y(_4813_)
);

NAND3X1 _11271_ (
    .A(_4465_),
    .B(_4466_),
    .C(_4464_),
    .Y(_4467_)
);

FILL FILL_1__9828_ (
);

FILL FILL_1__9408_ (
);

FILL FILL_0_CLKBUF1_insert90 (
);

FILL FILL_0_CLKBUF1_insert91 (
);

FILL FILL_0_CLKBUF1_insert92 (
);

FILL FILL_2__11733_ (
);

FILL FILL_0_CLKBUF1_insert93 (
);

FILL FILL_0_CLKBUF1_insert94 (
);

FILL FILL_2__11313_ (
);

NOR2X1 _8898_ (
    .A(_2321_),
    .B(_2320_),
    .Y(_2322_)
);

FILL FILL_0_CLKBUF1_insert95 (
);

OAI21X1 _8478_ (
    .A(_1912_),
    .B(_1915_),
    .C(_1914_),
    .Y(_1916_)
);

FILL FILL_0_CLKBUF1_insert96 (
);

AND2X2 _8058_ (
    .A(_1555_),
    .B(_1561_),
    .Y(_1562_)
);

FILL FILL_1__10306_ (
);

FILL FILL_0__7733_ (
);

FILL FILL_0__7313_ (
);

FILL FILL_1__13198_ (
);

OAI21X1 _12896_ (
    .A(_5920_),
    .B(_5924_),
    .C(_5927_),
    .Y(_5934_)
);

DFFPOSX1 _12476_ (
    .D(_5572_[15]),
    .CLK(clk_bF$buf22),
    .Q(_6377_[15])
);

OAI21X1 _12056_ (
    .A(_5172_),
    .B(_5171_),
    .C(_5168_),
    .Y(_5173_)
);

FILL FILL_2__12938_ (
);

FILL FILL_2__12518_ (
);

FILL FILL_0__13132_ (
);

FILL FILL_0__8938_ (
);

FILL FILL_0__8518_ (
);

FILL FILL_3__6615_ (
);

FILL FILL_1__9581_ (
);

FILL FILL_1__9161_ (
);

FILL FILL_3__9087_ (
);

FILL FILL_2__7084_ (
);

OAI21X1 _6964_ (
    .A(_511_),
    .B(_552_),
    .C(_551_),
    .Y(_558_)
);

INVX2 _6544_ (
    .A(Xin[6]),
    .Y(_144_)
);

FILL FILL_2__12691_ (
);

FILL FILL_2__12271_ (
);

FILL FILL_1__11684_ (
);

FILL FILL_1__11264_ (
);

FILL FILL_0__8691_ (
);

FILL FILL_0__8271_ (
);

FILL FILL_2__8289_ (
);

FILL FILL_0__10677_ (
);

NAND3X1 _10962_ (
    .A(_4157_),
    .B(_4123_),
    .C(_4161_),
    .Y(_4162_)
);

INVX1 _10542_ (
    .A(_3804_),
    .Y(_3814_)
);

FILL FILL_0__10257_ (
);

INVX1 _10122_ (
    .A(_3400_),
    .Y(_3401_)
);

FILL FILL_2__9650_ (
);

FILL FILL_2__9230_ (
);

NAND2X1 _7749_ (
    .A(gnd),
    .B(_1195_),
    .Y(_1265_)
);

INVX1 _7329_ (
    .A(_850_),
    .Y(_851_)
);

FILL FILL_2__13056_ (
);

FILL FILL_1__12889_ (
);

FILL FILL_1__12049_ (
);

FILL FILL_0__9896_ (
);

FILL FILL_0__9476_ (
);

FILL FILL_3__7573_ (
);

FILL FILL_0__9056_ (
);

INVX1 _11747_ (
    .A(_4867_),
    .Y(_4868_)
);

FILL FILL_3__7153_ (
);

NAND2X1 _11327_ (
    .A(_4521_),
    .B(_4501_),
    .Y(_4522_)
);

FILL FILL_1__13410_ (
);

FILL FILL_0__12823_ (
);

FILL FILL_0__12403_ (
);

FILL FILL_1__8852_ (
);

FILL FILL_1__8432_ (
);

FILL FILL_1__8012_ (
);

FILL FILL_3__8358_ (
);

NOR2X1 _7082_ (
    .A(_665_),
    .B(_666_),
    .Y(_667_)
);

FILL FILL_2__6775_ (
);

OAI21X1 _11080_ (
    .A(_4277_),
    .B(_4278_),
    .C(_4276_),
    .Y(_4279_)
);

FILL FILL_1__9637_ (
);

FILL FILL_1__9217_ (
);

FILL FILL_2__11962_ (
);

FILL FILL_2__11542_ (
);

FILL FILL_2__11122_ (
);

OAI21X1 _8287_ (
    .A(_2304_),
    .B(_1726_),
    .C(_1671_),
    .Y(_1727_)
);

FILL FILL_1__10955_ (
);

FILL FILL_1__10535_ (
);

FILL FILL_1__10115_ (
);

FILL FILL_0__7962_ (
);

FILL FILL_0__7542_ (
);

FILL FILL_0__7122_ (
);

AOI21X1 _12285_ (
    .A(_5339_),
    .B(_5341_),
    .C(_5396_),
    .Y(_5397_)
);

FILL FILL_2__8921_ (
);

FILL FILL_2__8501_ (
);

FILL FILL_2__12747_ (
);

FILL FILL_2__12327_ (
);

FILL FILL_0__8747_ (
);

FILL FILL_0__8327_ (
);

FILL FILL_1__9390_ (
);

FILL FILL_2__9706_ (
);

FILL FILL_1__7703_ (
);

NAND3X1 _6773_ (
    .A(_301_),
    .B(_362_),
    .C(_357_),
    .Y(_371_)
);

FILL FILL_2__12080_ (
);

FILL FILL_3__10879_ (
);

FILL FILL_3__10039_ (
);

FILL FILL_1__11493_ (
);

FILL FILL_1__11073_ (
);

FILL FILL_0__10486_ (
);

INVX1 _10771_ (
    .A(\X[5] [2]),
    .Y(_4755_)
);

AOI21X1 _10351_ (
    .A(_3618_),
    .B(_3614_),
    .C(_3573_),
    .Y(_3628_)
);

FILL FILL_0__10066_ (
);

FILL FILL_1__8908_ (
);

FILL FILL_3__11400_ (
);

FILL FILL_2__10813_ (
);

NOR2X1 _7978_ (
    .A(\u_fir_pe1.rYin [7]),
    .B(\u_fir_pe1.mul [7]),
    .Y(_1481_)
);

AOI21X1 _7558_ (
    .A(_1076_),
    .B(_1071_),
    .C(_932_),
    .Y(_1077_)
);

AOI21X1 _7138_ (
    .A(_703_),
    .B(_718_),
    .C(_721_),
    .Y(_722_)
);

FILL FILL_2__13285_ (
);

FILL FILL_0__6813_ (
);

FILL FILL_1__12698_ (
);

FILL FILL_1__12278_ (
);

FILL FILL_0__9285_ (
);

OR2X2 _11976_ (
    .A(_5089_),
    .B(_5088_),
    .Y(_5094_)
);

NOR2X1 _11556_ (
    .A(_4739_),
    .B(_4738_),
    .Y(_4740_)
);

NAND3X1 _11136_ (
    .A(_4327_),
    .B(_4328_),
    .C(_4329_),
    .Y(_4334_)
);

FILL FILL_0__12632_ (
);

FILL FILL_0__12212_ (
);

NOR2X1 _9704_ (
    .A(_3049_),
    .B(_3048_),
    .Y(_3050_)
);

FILL FILL_1__8661_ (
);

FILL FILL_1__8241_ (
);

FILL FILL_3__8587_ (
);

FILL FILL_0__13417_ (
);

FILL FILL_2__6584_ (
);

FILL FILL_1__9446_ (
);

FILL FILL_1__9026_ (
);

FILL FILL_2__11771_ (
);

FILL FILL_2__11351_ (
);

DFFPOSX1 _8096_ (
    .D(\X[1] [4]),
    .CLK(clk_bF$buf1),
    .Q(\X[2] [4])
);

FILL FILL_1__10764_ (
);

FILL FILL_1__10344_ (
);

FILL FILL_2__7789_ (
);

FILL FILL_0__7771_ (
);

FILL FILL_0__7351_ (
);

FILL FILL_2__7369_ (
);

AOI21X1 _12094_ (
    .A(_5197_),
    .B(_5204_),
    .C(_5179_),
    .Y(_5211_)
);

FILL FILL_2__8730_ (
);

FILL FILL_2__8310_ (
);

FILL FILL_3__13143_ (
);

NAND3X1 _6829_ (
    .A(_395_),
    .B(_423_),
    .C(_425_),
    .Y(_426_)
);

OAI21X1 _6409_ (
    .A(_4_),
    .B(_7_),
    .C(_1_),
    .Y(_12_)
);

FILL FILL_2__12976_ (
);

FILL FILL_2__12556_ (
);

FILL FILL_2__12136_ (
);

FILL FILL_0__13170_ (
);

FILL FILL_1__11969_ (
);

FILL FILL_1__11549_ (
);

FILL FILL_1__11129_ (
);

FILL FILL_0__8556_ (
);

FILL FILL_3__6653_ (
);

FILL FILL_0__8136_ (
);

NAND3X1 _10827_ (
    .A(_4018_),
    .B(_4026_),
    .C(_4028_),
    .Y(_4029_)
);

NAND3X1 _10407_ (
    .A(_3648_),
    .B(_3682_),
    .C(_3680_),
    .Y(_3683_)
);

FILL FILL_1__12910_ (
);

NOR2X1 _13299_ (
    .A(_6321_),
    .B(_6322_),
    .Y(_6323_)
);

FILL FILL_2__9935_ (
);

FILL FILL_0__11903_ (
);

FILL FILL_2__9515_ (
);

FILL FILL_1__7932_ (
);

FILL FILL_1__7512_ (
);

FILL FILL_3__7438_ (
);

OAI21X1 _6582_ (
    .A(_180_),
    .B(_181_),
    .C(_179_),
    .Y(_182_)
);

FILL FILL254550x97350 (
);

FILL FILL_3__10268_ (
);

FILL FILL_0__10295_ (
);

NOR2X1 _10580_ (
    .A(\u_fir_pe4.rYin [4]),
    .B(\u_fir_pe4.mul [4]),
    .Y(_3846_)
);

OAI21X1 _10160_ (
    .A(_3438_),
    .B(_3433_),
    .C(_3427_),
    .Y(_3439_)
);

FILL FILL_1__8717_ (
);

FILL FILL_2__10622_ (
);

FILL FILL_2__10202_ (
);

INVX1 _7787_ (
    .A(_1302_),
    .Y(_1303_)
);

NAND3X1 _7367_ (
    .A(_883_),
    .B(_887_),
    .C(_885_),
    .Y(_888_)
);

FILL FILL_2__13094_ (
);

FILL FILL_0__6622_ (
);

FILL FILL_1__12087_ (
);

FILL FILL_0__9094_ (
);

NAND3X1 _11785_ (
    .A(_4835_),
    .B(_4899_),
    .C(_4900_),
    .Y(_4906_)
);

INVX1 _11365_ (
    .A(_4556_),
    .Y(_4559_)
);

FILL FILL_2__11827_ (
);

FILL FILL_0__12861_ (
);

FILL FILL_2__11407_ (
);

FILL FILL_0__12441_ (
);

FILL FILL_0__12021_ (
);

FILL FILL_0__7827_ (
);

AOI22X1 _9933_ (
    .A(\X[4] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[4] [4]),
    .Y(_3215_)
);

FILL FILL_0__7407_ (
);

AND2X2 _9513_ (
    .A(\X[3]_5_bF$buf3 ),
    .B(vdd),
    .Y(_2869_)
);

FILL FILL_1__8890_ (
);

FILL FILL_1__8470_ (
);

FILL FILL_1__8050_ (
);

FILL FILL_0__13226_ (
);

FILL FILL_2__6393_ (
);

FILL FILL_3__6709_ (
);

FILL FILL_1__9675_ (
);

FILL FILL_1__9255_ (
);

FILL FILL_2__11580_ (
);

FILL FILL_2__11160_ (
);

FILL FILL_1__10993_ (
);

FILL FILL_1__10573_ (
);

FILL FILL_1__10153_ (
);

FILL FILL_2__7598_ (
);

FILL FILL_0__7580_ (
);

FILL FILL_2__7178_ (
);

FILL FILL_0__7160_ (
);

FILL FILL_3__10900_ (
);

NAND3X1 _6638_ (
    .A(_225_),
    .B(_234_),
    .C(_236_),
    .Y(_237_)
);

FILL FILL_2__12785_ (
);

FILL FILL_2__12365_ (
);

FILL FILL_1__11778_ (
);

FILL FILL_1__11358_ (
);

FILL FILL_0__8785_ (
);

FILL FILL_3__6882_ (
);

FILL FILL_0__8365_ (
);

AND2X2 _10636_ (
    .A(\u_fir_pe4.rYin [9]),
    .B(\u_fir_pe4.mul [9]),
    .Y(_3900_)
);

NOR2X1 _10216_ (
    .A(_3958_),
    .B(_3493_),
    .Y(_3494_)
);

FILL FILL_2__9744_ (
);

FILL FILL_2__9324_ (
);

FILL FILL_0__11712_ (
);

FILL FILL_1__7741_ (
);

FILL FILL_1__7321_ (
);

FILL FILL_3__7667_ (
);

NOR2X1 _6391_ (
    .A(_780_),
    .B(_760_),
    .Y(_783_)
);

FILL FILL_0__12917_ (
);

FILL FILL_3__10497_ (
);

FILL FILL_1__8946_ (
);

FILL FILL_1__8526_ (
);

FILL FILL_2__10851_ (
);

FILL FILL_2__10431_ (
);

FILL FILL_2__10011_ (
);

OAI21X1 _7596_ (
    .A(_1035_),
    .B(_1113_),
    .C(_1057_),
    .Y(_1114_)
);

INVX1 _7176_ (
    .A(\u_fir_pe0.rYin [14]),
    .Y(_759_)
);

FILL FILL_2__6869_ (
);

FILL FILL_0__6851_ (
);

FILL FILL_0__6431_ (
);

FILL FILL_2__6449_ (
);

DFFPOSX1 _11594_ (
    .D(_4775_[10]),
    .CLK(clk_bF$buf50),
    .Q(\Y[6] [10])
);

NAND2X1 _11174_ (
    .A(\X[5] [2]),
    .B(gnd),
    .Y(_4371_)
);

FILL FILL_2__7810_ (
);

FILL FILL_3__12643_ (
);

FILL FILL_3__12223_ (
);

FILL FILL_0__12670_ (
);

FILL FILL_2__11216_ (
);

FILL FILL_0__12250_ (
);

FILL FILL_1__10629_ (
);

FILL FILL_1__10209_ (
);

FILL FILL_0__7636_ (
);

NAND2X1 _9742_ (
    .A(_3048_),
    .B(_3060_),
    .Y(_3085_)
);

OAI21X1 _9322_ (
    .A(_2598_),
    .B(_2595_),
    .C(_2680_),
    .Y(_2681_)
);

AND2X2 _12799_ (
    .A(_5816_),
    .B(_5811_),
    .Y(_5838_)
);

AND2X2 _12379_ (
    .A(_5441_),
    .B(_5451_),
    .Y(_5483_)
);

FILL FILL_3__13008_ (
);

FILL FILL_0__13035_ (
);

AND2X2 _13320_ (
    .A(_6337_),
    .B(_6343_),
    .Y(_6344_)
);

FILL FILL_3__6938_ (
);

FILL FILL_1__9484_ (
);

FILL FILL_1__9064_ (
);

FILL FILL_1__10382_ (
);

NOR3X1 _6867_ (
    .A(_305_),
    .B(_132_),
    .C(_321_),
    .Y(_463_)
);

NAND3X1 _6447_ (
    .A(_29_),
    .B(_45_),
    .C(_48_),
    .Y(_49_)
);

FILL FILL_2__12594_ (
);

FILL FILL_2__12174_ (
);

FILL FILL_1__11167_ (
);

FILL FILL_0__8594_ (
);

FILL FILL_0__8174_ (
);

NAND3X1 _10865_ (
    .A(_4055_),
    .B(_4063_),
    .C(_4065_),
    .Y(_4066_)
);

OAI21X1 _10445_ (
    .A(_3719_),
    .B(_3718_),
    .C(_3712_),
    .Y(_3720_)
);

NAND3X1 _10025_ (
    .A(_3214_),
    .B(_3301_),
    .C(_3302_),
    .Y(_3306_)
);

FILL FILL_2__10907_ (
);

FILL FILL_2__9973_ (
);

FILL FILL_2__9553_ (
);

FILL FILL_0__11941_ (
);

FILL FILL_2__9133_ (
);

FILL FILL_0__11521_ (
);

FILL FILL_0__11101_ (
);

FILL FILL_0__6907_ (
);

FILL FILL_1__7970_ (
);

FILL FILL_1__7550_ (
);

FILL FILL_1__7130_ (
);

FILL FILL_0__9799_ (
);

FILL FILL_3__7896_ (
);

FILL FILL_0__9379_ (
);

FILL FILL_3__7056_ (
);

FILL FILL_1__13313_ (
);

FILL FILL_0__12726_ (
);

FILL FILL_0__12306_ (
);

FILL FILL_1__8755_ (
);

FILL FILL_1__8335_ (
);

FILL FILL_2__10660_ (
);

FILL FILL_2__10240_ (
);

FILL FILL_3__9622_ (
);

FILL FILL_3__9202_ (
);

FILL FILL_0__6660_ (
);

FILL FILL_2__6678_ (
);

FILL FILL_3__12872_ (
);

FILL FILL_3__12452_ (
);

FILL FILL_2__11865_ (
);

FILL FILL_2__11445_ (
);

FILL FILL_2__11025_ (
);

FILL FILL_1__10858_ (
);

FILL FILL_1__10438_ (
);

FILL FILL_1__10018_ (
);

FILL FILL_0__7865_ (
);

AOI21X1 _9971_ (
    .A(_3249_),
    .B(_3252_),
    .C(_3243_),
    .Y(_3253_)
);

FILL FILL_0__7445_ (
);

NAND2X1 _9551_ (
    .A(_2859_),
    .B(_2860_),
    .Y(_2906_)
);

FILL FILL_0__7025_ (
);

NAND3X1 _9131_ (
    .A(_2487_),
    .B(_2473_),
    .C(_2491_),
    .Y(_2492_)
);

NAND2X1 _12188_ (
    .A(gnd),
    .B(_5256_),
    .Y(_5303_)
);

FILL FILL_2__8824_ (
);

FILL FILL_2__8404_ (
);

FILL FILL_3__13237_ (
);

FILL FILL_0__13264_ (
);

FILL FILL_1__6821_ (
);

FILL FILL_1__6401_ (
);

FILL FILL_3__6747_ (
);

FILL FILL_1__9293_ (
);

FILL FILL_2_CLKBUF1_insert40 (
);

FILL FILL_2_CLKBUF1_insert41 (
);

FILL FILL_2__9609_ (
);

FILL FILL_2_CLKBUF1_insert42 (
);

FILL FILL_2_CLKBUF1_insert43 (
);

FILL FILL_2_CLKBUF1_insert44 (
);

FILL FILL_2_CLKBUF1_insert45 (
);

FILL FILL_2_CLKBUF1_insert46 (
);

FILL FILL_2_CLKBUF1_insert47 (
);

FILL FILL_2_CLKBUF1_insert48 (
);

FILL FILL_1__10191_ (
);

FILL FILL_2_CLKBUF1_insert49 (
);

FILL FILL_1__7606_ (
);

INVX1 _6676_ (
    .A(_177_),
    .Y(_275_)
);

FILL FILL_1__11396_ (
);

FILL FILL_0__10389_ (
);

OAI21X1 _10674_ (
    .A(_3930_),
    .B(_3931_),
    .C(_3935_),
    .Y(_3937_)
);

OAI21X1 _10254_ (
    .A(_3523_),
    .B(_3517_),
    .C(_3525_),
    .Y(_3532_)
);

FILL FILL_3__11723_ (
);

FILL FILL_2__9782_ (
);

FILL FILL_2__9362_ (
);

FILL FILL_0__11750_ (
);

FILL FILL_0__11330_ (
);

FILL FILL_2__13188_ (
);

FILL FILL_0__6716_ (
);

NAND2X1 _8822_ (
    .A(_2247_),
    .B(_2248_),
    .Y(_2384_[3])
);

NAND2X1 _8402_ (
    .A(_1752_),
    .B(_1836_),
    .Y(_1841_)
);

FILL FILL_0__9188_ (
);

NAND2X1 _11879_ (
    .A(_4995_),
    .B(_4997_),
    .Y(_4998_)
);

FILL FILL_3__7285_ (
);

INVX1 _11459_ (
    .A(_4635_),
    .Y(_4645_)
);

NAND3X1 _11039_ (
    .A(_4231_),
    .B(_4234_),
    .C(_4232_),
    .Y(_4238_)
);

FILL FILL_1__13122_ (
);

FILL FILL_0__12955_ (
);

AOI21X1 _12820_ (
    .A(_5858_),
    .B(_5853_),
    .C(_5714_),
    .Y(_5859_)
);

FILL FILL_0__12535_ (
);

FILL FILL_0__12115_ (
);

AOI21X1 _12400_ (
    .A(_5485_),
    .B(_5500_),
    .C(_5503_),
    .Y(_5504_)
);

OR2X2 _9607_ (
    .A(_2960_),
    .B(_2956_),
    .Y(_2961_)
);

FILL FILL_1__8564_ (
);

FILL FILL_1__8144_ (
);

FILL FILL_3__9431_ (
);

FILL FILL_2__6487_ (
);

FILL FILL_1__9769_ (
);

FILL FILL_1__9349_ (
);

FILL FILL_2__11674_ (
);

FILL FILL_2__11254_ (
);

FILL FILL_1__10667_ (
);

FILL FILL_1__10247_ (
);

FILL FILL_0__7674_ (
);

AND2X2 _9780_ (
    .A(\u_fir_pe3.rYin [11]),
    .B(\u_fir_pe3.mul [11]),
    .Y(_3124_)
);

AND2X2 _9360_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .Y(_2718_)
);

FILL FILL_2__8633_ (
);

FILL FILL_2__8213_ (
);

FILL FILL_0__10601_ (
);

FILL FILL_2__12879_ (
);

FILL FILL_2__12459_ (
);

FILL FILL_2__12039_ (
);

FILL FILL_0__13073_ (
);

FILL FILL_1__6630_ (
);

FILL FILL_2__13400_ (
);

FILL FILL_0__8879_ (
);

FILL FILL_3__6976_ (
);

FILL FILL_0__8459_ (
);

FILL FILL_3__6556_ (
);

FILL FILL_0__8039_ (
);

FILL FILL_1__12813_ (
);

FILL FILL_0__9820_ (
);

FILL FILL_2__9418_ (
);

FILL FILL_0__9400_ (
);

FILL FILL_0__11806_ (
);

FILL FILL_1__7835_ (
);

FILL FILL_1__7415_ (
);

INVX1 _6485_ (
    .A(_85_),
    .Y(_86_)
);

AOI21X1 _10483_ (
    .A(gnd),
    .B(_3754_),
    .C(_3756_),
    .Y(_3757_)
);

FILL FILL_0__10198_ (
);

OAI22X1 _10063_ (
    .A(_3230_),
    .B(_3341_),
    .C(_3273_),
    .D(_3342_),
    .Y(_3343_)
);

FILL FILL_3__11952_ (
);

FILL FILL_3__11532_ (
);

FILL FILL_3__11112_ (
);

FILL FILL_2__10945_ (
);

FILL FILL_2__9591_ (
);

FILL FILL_2__10525_ (
);

FILL FILL_2__9171_ (
);

FILL FILL_2__10105_ (
);

FILL FILL_3__9907_ (
);

FILL FILL_0__6945_ (
);

FILL FILL_0__6525_ (
);

NAND2X1 _8631_ (
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_2067_)
);

OAI21X1 _8211_ (
    .A(_2375_),
    .B(_1612_),
    .C(_1615_),
    .Y(_1653_)
);

NOR2X1 _11688_ (
    .A(_4809_),
    .B(_4808_),
    .Y(_4810_)
);

FILL FILL_3__7094_ (
);

NAND2X1 _11268_ (
    .A(_4462_),
    .B(_4463_),
    .Y(_4464_)
);

FILL FILL_2__7904_ (
);

FILL FILL_3__12737_ (
);

FILL FILL_3__12317_ (
);

FILL FILL_0__12764_ (
);

FILL FILL_0__12344_ (
);

FILL FILL254550x183750 (
);

DFFPOSX1 _9836_ (
    .D(_3181_[6]),
    .CLK(clk_bF$buf15),
    .Q(\Y[4] [6])
);

OAI21X1 _9416_ (
    .A(_2692_),
    .B(_2772_),
    .C(_2755_),
    .Y(_2773_)
);

FILL FILL_1__8793_ (
);

FILL FILL_1__8373_ (
);

FILL FILL_3__8299_ (
);

FILL FILL_3__9240_ (
);

FILL FILL_0__13129_ (
);

BUFX2 _13414_ (
    .A(_6377_[6]),
    .Y(Yout[6])
);

FILL FILL_1__9998_ (
);

FILL FILL_1__9578_ (
);

FILL FILL_1__9158_ (
);

FILL FILL_3__12070_ (
);

FILL FILL_2__11483_ (
);

FILL FILL_2__11063_ (
);

FILL FILL_1__10896_ (
);

FILL FILL_1__10476_ (
);

FILL FILL_1__10056_ (
);

FILL FILL_0__7483_ (
);

FILL FILL_0__7063_ (
);

FILL FILL_2__8862_ (
);

FILL FILL_2__8442_ (
);

FILL FILL_0__10830_ (
);

FILL FILL_0__10410_ (
);

FILL FILL_2__8022_ (
);

FILL FILL_2__12688_ (
);

FILL FILL_2__12268_ (
);

OAI21X1 _7902_ (
    .A(_1391_),
    .B(_1398_),
    .C(_1397_),
    .Y(_1414_)
);

FILL FILL_0__8688_ (
);

FILL FILL_0__8268_ (
);

OAI21X1 _10959_ (
    .A(_4154_),
    .B(_4155_),
    .C(_4140_),
    .Y(_4159_)
);

INVX1 _10539_ (
    .A(_3770_),
    .Y(_3811_)
);

NAND2X1 _10119_ (
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3398_)
);

FILL FILL_1__12622_ (
);

FILL FILL_1__12202_ (
);

FILL FILL_2__9647_ (
);

FILL FILL_2__9227_ (
);

NAND3X1 _11900_ (
    .A(_5007_),
    .B(_5016_),
    .C(_5018_),
    .Y(_5019_)
);

FILL FILL_1__7644_ (
);

FILL FILL_1__13407_ (
);

FILL FILL_3__8511_ (
);

AOI21X1 _10292_ (
    .A(_3549_),
    .B(_3548_),
    .C(_3491_),
    .Y(_3569_)
);

FILL FILL_1__8849_ (
);

FILL FILL_1__8429_ (
);

FILL FILL_1__8009_ (
);

FILL FILL_3__11341_ (
);

FILL FILL_2__10334_ (
);

OAI21X1 _7499_ (
    .A(_1016_),
    .B(_1017_),
    .C(_1007_),
    .Y(_1018_)
);

OAI21X1 _7079_ (
    .A(_655_),
    .B(_656_),
    .C(_662_),
    .Y(_664_)
);

FILL FILL_0__6754_ (
);

NAND2X1 _8860_ (
    .A(_2279_),
    .B(_2282_),
    .Y(_2384_[7])
);

OAI21X1 _8440_ (
    .A(_1878_),
    .B(_1874_),
    .C(_1790_),
    .Y(_1879_)
);

NOR2X1 _8020_ (
    .A(\u_fir_pe1.rYin [10]),
    .B(\u_fir_pe1.mul [10]),
    .Y(_1524_)
);

OAI21X1 _11497_ (
    .A(_4650_),
    .B(_4651_),
    .C(_4679_),
    .Y(_4680_)
);

NOR2X1 _11077_ (
    .A(_4192_),
    .B(_4189_),
    .Y(_4276_)
);

FILL FILL_3__12966_ (
);

FILL FILL_2__7713_ (
);

FILL FILL_1__13160_ (
);

FILL FILL_2__11959_ (
);

FILL FILL_0__12993_ (
);

FILL FILL_2__11539_ (
);

FILL FILL_0__12573_ (
);

FILL FILL_2__11119_ (
);

FILL FILL_0__12153_ (
);

FILL FILL_2__12900_ (
);

FILL FILL_0__7959_ (
);

FILL FILL_0__7539_ (
);

AND2X2 _9645_ (
    .A(_2994_),
    .B(_2993_),
    .Y(_2998_)
);

FILL FILL_0__7119_ (
);

OAI21X1 _9225_ (
    .A(_2584_),
    .B(_2579_),
    .C(_2507_),
    .Y(_2585_)
);

FILL FILL_1__8182_ (
);

FILL FILL_0__8900_ (
);

FILL FILL_2__8918_ (
);

NOR2X1 _13223_ (
    .A(_6247_),
    .B(_6246_),
    .Y(_6248_)
);

FILL FILL_1__6915_ (
);

FILL FILL_1__9387_ (
);

FILL FILL_2__11292_ (
);

FILL FILL_1__10285_ (
);

FILL FILL_0__7292_ (
);

FILL FILL_2__8671_ (
);

FILL FILL_2__8251_ (
);

FILL FILL_3__13084_ (
);

FILL FILL_2__12077_ (
);

NAND3X1 _7711_ (
    .A(_1223_),
    .B(_1227_),
    .C(_1182_),
    .Y(_1228_)
);

FILL FILL_0__8497_ (
);

FILL FILL_3__6594_ (
);

NOR2X1 _10768_ (
    .A(_4674_),
    .B(_4716_),
    .Y(_4725_)
);

NAND3X1 _10348_ (
    .A(_3571_),
    .B(_3619_),
    .C(_3624_),
    .Y(_3625_)
);

FILL FILL_3__11817_ (
);

FILL FILL_1__12851_ (
);

FILL FILL_1__12431_ (
);

FILL FILL_1__12011_ (
);

FILL FILL_2__9456_ (
);

FILL FILL_0__11844_ (
);

FILL FILL_2__9036_ (
);

FILL FILL_0__11424_ (
);

FILL FILL_0__11004_ (
);

NOR2X1 _8916_ (
    .A(_2339_),
    .B(_2338_),
    .Y(_2340_)
);

FILL FILL_1__7873_ (
);

FILL FILL_1__7453_ (
);

FILL FILL_1__7033_ (
);

FILL FILL_3__7379_ (
);

FILL FILL_1__13216_ (
);

FILL FILL_3__8740_ (
);

FILL FILL_0__12629_ (
);

NAND2X1 _12914_ (
    .A(_5951_),
    .B(_5946_),
    .Y(_5952_)
);

FILL FILL_0__12209_ (
);

FILL FILL_1__8658_ (
);

FILL FILL_1__8238_ (
);

FILL FILL_2__10983_ (
);

FILL FILL_2__10563_ (
);

FILL FILL_2__10143_ (
);

FILL FILL_3__9525_ (
);

FILL FILL_0__6983_ (
);

FILL FILL_0__6563_ (
);

FILL FILL_2__7942_ (
);

FILL FILL_2__7522_ (
);

FILL FILL_2__7102_ (
);

FILL FILL_2__11768_ (
);

FILL FILL_2__11348_ (
);

FILL FILL_0__12382_ (
);

FILL FILL_0__7768_ (
);

DFFPOSX1 _9874_ (
    .D(_3186_[4]),
    .CLK(clk_bF$buf14),
    .Q(\u_fir_pe3.mul [4])
);

FILL FILL_0__7348_ (
);

NAND2X1 _9454_ (
    .A(_2794_),
    .B(_2804_),
    .Y(_2811_)
);

NAND3X1 _9034_ (
    .A(_2392_),
    .B(_2396_),
    .C(_2394_),
    .Y(_2397_)
);

FILL FILL_1__11702_ (
);

FILL FILL_2__8727_ (
);

FILL FILL_2__8307_ (
);

FILL FILL_0__13167_ (
);

NAND2X1 _13032_ (
    .A(_6064_),
    .B(_6051_),
    .Y(_6068_)
);

FILL FILL_1__6724_ (
);

FILL FILL_1__9196_ (
);

FILL FILL_1__12907_ (
);

FILL FILL_0__9914_ (
);

FILL FILL_1__10094_ (
);

FILL FILL_1__7929_ (
);

FILL FILL_3__10841_ (
);

FILL FILL_1__7509_ (
);

FILL FILL_3__10421_ (
);

FILL FILL_2__8480_ (
);

FILL FILL_2__8060_ (
);

INVX1 _6999_ (
    .A(_566_),
    .Y(_592_)
);

AOI21X1 _6579_ (
    .A(_82_),
    .B(_100_),
    .C(_178_),
    .Y(_179_)
);

NOR2X1 _7940_ (
    .A(_1445_),
    .B(_1446_),
    .Y(_1447_)
);

AND2X2 _7520_ (
    .A(vdd),
    .B(\X[1]_5_bF$buf3 ),
    .Y(_1039_)
);

FILL FILL_1__11299_ (
);

NOR2X1 _7100_ (
    .A(_681_),
    .B(_682_),
    .Y(_683_)
);

INVX1 _10997_ (
    .A(_4195_),
    .Y(_4196_)
);

INVX1 _10577_ (
    .A(\u_fir_pe4.rYin [4]),
    .Y(_3843_)
);

AOI22X1 _10157_ (
    .A(gnd),
    .B(\X[4] [4]),
    .C(gnd),
    .D(\X[4]_5_bF$buf3 ),
    .Y(_3436_)
);

FILL FILL_1__12660_ (
);

FILL FILL_3__11206_ (
);

FILL FILL_1__12240_ (
);

FILL FILL253950x75750 (
);

FILL FILL_2__9685_ (
);

FILL FILL_2__10619_ (
);

FILL FILL_2__9265_ (
);

FILL FILL_0__11653_ (
);

FILL FILL_0__11233_ (
);

FILL FILL_0__6619_ (
);

NOR2X1 _8725_ (
    .A(_1668_),
    .B(_2056_),
    .Y(_2159_)
);

NAND3X1 _8305_ (
    .A(_1733_),
    .B(_1742_),
    .C(_1744_),
    .Y(_1745_)
);

FILL FILL_1__7682_ (
);

FILL FILL_1__7262_ (
);

FILL FILL_3__7188_ (
);

FILL FILL_1__13025_ (
);

FILL FILL_0__12858_ (
);

AND2X2 _12723_ (
    .A(_5713_),
    .B(_5714_),
    .Y(_5763_)
);

FILL FILL_0__12438_ (
);

FILL FILL_0__12018_ (
);

INVX1 _12303_ (
    .A(_4806_),
    .Y(_5573_[0])
);

FILL FILL_1__8887_ (
);

FILL FILL_1__8467_ (
);

FILL FILL_1__8047_ (
);

FILL FILL_2__10792_ (
);

FILL FILL_2__10372_ (
);

FILL FILL_0__6792_ (
);

FILL FILL_2__7751_ (
);

FILL FILL_3__12584_ (
);

FILL FILL_2__7331_ (
);

FILL FILL_3__12164_ (
);

FILL FILL_2__11997_ (
);

FILL FILL_2__11577_ (
);

FILL FILL_2__11157_ (
);

FILL FILL_0__12191_ (
);

FILL FILL_0__7997_ (
);

FILL FILL_0__7577_ (
);

OAI21X1 _9683_ (
    .A(_3023_),
    .B(_3024_),
    .C(_3028_),
    .Y(_3031_)
);

FILL FILL_0__7157_ (
);

INVX1 _9263_ (
    .A(_2621_),
    .Y(_2622_)
);

FILL FILL_1__11931_ (
);

FILL FILL_1__11511_ (
);

FILL FILL_2__8536_ (
);

FILL FILL_0__10924_ (
);

FILL FILL_0__10504_ (
);

FILL FILL_0__13396_ (
);

INVX1 _13261_ (
    .A(_6282_),
    .Y(_6285_)
);

FILL FILL_1__6953_ (
);

FILL FILL_1__6533_ (
);

FILL FILL_2__13303_ (
);

FILL FILL_1__12716_ (
);

FILL FILL_0__9723_ (
);

FILL FILL_3__7820_ (
);

FILL FILL_0__9303_ (
);

FILL FILL_0__11709_ (
);

FILL FILL_1__7738_ (
);

FILL FILL_3__10650_ (
);

FILL FILL_1__7318_ (
);

NOR2X1 _6388_ (
    .A(_770_),
    .B(_778_),
    .Y(_780_)
);

FILL FILL_3__8605_ (
);

NOR2X1 _10386_ (
    .A(_3661_),
    .B(_3604_),
    .Y(_3662_)
);

FILL FILL_2__6602_ (
);

FILL FILL_3__11435_ (
);

FILL FILL_2__10848_ (
);

FILL FILL_2__9494_ (
);

FILL FILL_0__11882_ (
);

FILL FILL_2__10428_ (
);

FILL FILL_2__9074_ (
);

FILL FILL_0__11462_ (
);

FILL FILL_2__10008_ (
);

FILL FILL_0__11042_ (
);

FILL FILL_0__6848_ (
);

DFFPOSX1 _8954_ (
    .D(_2384_[1]),
    .CLK(clk_bF$buf56),
    .Q(\Y[3] [1])
);

FILL FILL_0__6428_ (
);

NAND2X1 _8534_ (
    .A(_1971_),
    .B(_1970_),
    .Y(_1972_)
);

DFFPOSX1 _8114_ (
    .D(\Y[1] [14]),
    .CLK(clk_bF$buf25),
    .Q(\u_fir_pe1.rYin [14])
);

FILL FILL_1__7491_ (
);

FILL FILL_1__7071_ (
);

FILL FILL_2__7807_ (
);

FILL FILL_1__13254_ (
);

NAND2X1 _12952_ (
    .A(vdd),
    .B(\X[6] [7]),
    .Y(_5989_)
);

FILL FILL_0__12667_ (
);

FILL FILL_0__12247_ (
);

NAND2X1 _12532_ (
    .A(_6299_),
    .B(_6363_),
    .Y(_6364_)
);

AOI21X1 _12112_ (
    .A(_5228_),
    .B(_5227_),
    .C(_5220_),
    .Y(_5229_)
);

INVX1 _9739_ (
    .A(\u_fir_pe3.mul [8]),
    .Y(_3082_)
);

NAND3X1 _9319_ (
    .A(_2526_),
    .B(_2665_),
    .C(_2670_),
    .Y(_2678_)
);

FILL FILL_1__8696_ (
);

FILL FILL_1__8276_ (
);

FILL FILL_2__10181_ (
);

FILL FILL_3__9983_ (
);

FILL FILL_3__9563_ (
);

FILL FILL_3__9143_ (
);

NOR2X1 _13317_ (
    .A(_6338_),
    .B(_6340_),
    .Y(_6341_)
);

FILL FILL253650x212550 (
);

FILL FILL_1_CLKBUF1_insert50 (
);

FILL FILL_1_CLKBUF1_insert51 (
);

FILL FILL_1_CLKBUF1_insert52 (
);

FILL FILL_1_CLKBUF1_insert53 (
);

FILL FILL_1_CLKBUF1_insert54 (
);

FILL FILL_2__7980_ (
);

FILL FILL_1_CLKBUF1_insert55 (
);

FILL FILL_2__7560_ (
);

FILL FILL_3__12393_ (
);

FILL FILL_1_CLKBUF1_insert56 (
);

FILL FILL_2__7140_ (
);

FILL FILL_1_CLKBUF1_insert57 (
);

FILL FILL_1_CLKBUF1_insert58 (
);

FILL FILL_1_CLKBUF1_insert59 (
);

FILL FILL_2__11386_ (
);

FILL FILL_1__10799_ (
);

AOI21X1 _6600_ (
    .A(_182_),
    .B(_177_),
    .C(_184_),
    .Y(_200_)
);

FILL FILL_1__10379_ (
);

FILL FILL_0__7386_ (
);

AOI21X1 _9492_ (
    .A(_2763_),
    .B(_2833_),
    .C(_2847_),
    .Y(_2848_)
);

NAND3X1 _9072_ (
    .A(gnd),
    .B(\X[3] [1]),
    .C(_2433_),
    .Y(_2434_)
);

FILL FILL_1__11740_ (
);

FILL FILL_1__11320_ (
);

FILL FILL_2__8765_ (
);

FILL FILL_2__8345_ (
);

FILL FILL_3__13178_ (
);

FILL FILL_0__10313_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

NAND2X1 _13070_ (
    .A(gnd),
    .B(\X[6] [7]),
    .Y(_6105_)
);

NAND3X1 _7805_ (
    .A(_1317_),
    .B(_1318_),
    .C(_1319_),
    .Y(_1320_)
);

FILL FILL_1__6762_ (
);

FILL FILL_2__13112_ (
);

FILL FILL_3__6688_ (
);

FILL FILL_1__12945_ (
);

FILL FILL_1__12525_ (
);

FILL FILL_1__12105_ (
);

FILL FILL_0__9952_ (
);

FILL FILL_0__9532_ (
);

FILL FILL_0__11938_ (
);

FILL FILL_0__9112_ (
);

AND2X2 _11803_ (
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_4923_)
);

FILL FILL_0__11518_ (
);

FILL FILL_1__7967_ (
);

FILL FILL_1__7547_ (
);

FILL FILL_1__7127_ (
);

FILL FILL_3__8834_ (
);

NAND3X1 _10195_ (
    .A(_3469_),
    .B(_3470_),
    .C(_3471_),
    .Y(_3474_)
);

FILL FILL_2__6831_ (
);

FILL FILL_3__11664_ (
);

FILL FILL_2__6411_ (
);

FILL FILL_2__10657_ (
);

FILL FILL_0__11691_ (
);

FILL FILL_2__10237_ (
);

FILL FILL_0__11271_ (
);

FILL FILL_3__9619_ (
);

FILL FILL_0__6657_ (
);

NAND2X1 _8763_ (
    .A(_2188_),
    .B(_2195_),
    .Y(_2196_)
);

AOI21X1 _8343_ (
    .A(_1695_),
    .B(_1699_),
    .C(_1663_),
    .Y(_1783_)
);

FILL FILL_2__7616_ (
);

FILL FILL_1__13063_ (
);

FILL FILL_0__12896_ (
);

OAI21X1 _12761_ (
    .A(_5798_),
    .B(_5799_),
    .C(_5789_),
    .Y(_5800_)
);

FILL FILL_0__12056_ (
);

OAI21X1 _12341_ (
    .A(_5437_),
    .B(_5438_),
    .C(_5444_),
    .Y(_5446_)
);

FILL FILL_2__12803_ (
);

INVX1 _9968_ (
    .A(_3233_),
    .Y(_3250_)
);

NAND2X1 _9548_ (
    .A(_2896_),
    .B(_2900_),
    .Y(_2903_)
);

AOI21X1 _9128_ (
    .A(_2483_),
    .B(_2485_),
    .C(_2476_),
    .Y(_2489_)
);

FILL FILL_0__8803_ (
);

FILL FILL_3__9792_ (
);

FILL FILL254550x115350 (
);

INVX1 _13126_ (
    .A(_6159_),
    .Y(_6160_)
);

FILL FILL_1__6818_ (
);

FILL FILL_2__11195_ (
);

FILL FILL_1__10188_ (
);

FILL FILL_0__7195_ (
);

FILL FILL_3__10935_ (
);

FILL FILL_3__10515_ (
);

FILL FILL_2__8574_ (
);

FILL FILL_0__10962_ (
);

FILL FILL_2__8154_ (
);

FILL FILL_0__10542_ (
);

FILL FILL_0__10122_ (
);

AOI21X1 _7614_ (
    .A(_1129_),
    .B(_1131_),
    .C(_1127_),
    .Y(_1132_)
);

FILL FILL_1__6991_ (
);

FILL FILL_1__6571_ (
);

FILL FILL_3__6497_ (
);

FILL FILL_1__12754_ (
);

FILL FILL_1__12334_ (
);

FILL FILL_0__9761_ (
);

FILL FILL_2__9779_ (
);

FILL FILL_2__9359_ (
);

FILL FILL_0__9341_ (
);

FILL FILL_0__11747_ (
);

DFFPOSX1 _11612_ (
    .D(\Y[5] [4]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.rYin [4])
);

FILL FILL_0__11327_ (
);

NOR2X1 _8819_ (
    .A(_2245_),
    .B(_2244_),
    .Y(_2246_)
);

FILL FILL_1__7776_ (
);

FILL FILL_1__7356_ (
);

FILL FILL_1__13119_ (
);

NAND3X1 _12817_ (
    .A(_5850_),
    .B(_5849_),
    .C(_5851_),
    .Y(_5856_)
);

FILL FILL_3__8223_ (
);

FILL FILL_3__11893_ (
);

FILL FILL_2__6640_ (
);

FILL FILL_3__11473_ (
);

FILL FILL_3__11053_ (
);

FILL FILL_2__10886_ (
);

FILL FILL_2__10466_ (
);

FILL FILL_2__10046_ (
);

FILL FILL_0__11080_ (
);

FILL FILL_1__9922_ (
);

FILL FILL_1__9502_ (
);

FILL FILL_0__6886_ (
);

DFFPOSX1 _8992_ (
    .D(\Y[2] [15]),
    .CLK(clk_bF$buf42),
    .Q(\u_fir_pe2.rYin [15])
);

FILL FILL_0__6466_ (
);

NAND3X1 _8572_ (
    .A(_1994_),
    .B(_2001_),
    .C(_2008_),
    .Y(_2009_)
);

INVX1 _8152_ (
    .A(_1594_),
    .Y(_1595_)
);

FILL FILL_1__10820_ (
);

FILL FILL_1__10400_ (
);

FILL FILL_2__7845_ (
);

FILL FILL_3__12678_ (
);

FILL FILL_2__7425_ (
);

FILL FILL_3__12258_ (
);

FILL FILL_2__7005_ (
);

FILL FILL_1__13292_ (
);

AOI21X1 _12990_ (
    .A(_6015_),
    .B(_6010_),
    .C(_5962_),
    .Y(_6027_)
);

FILL FILL_0__12285_ (
);

NAND2X1 _12570_ (
    .A(gnd),
    .B(\X[6] [3]),
    .Y(_5612_)
);

NAND2X1 _12150_ (
    .A(_5265_),
    .B(_5254_),
    .Y(_5266_)
);

FILL FILL_2__12612_ (
);

OAI21X1 _9777_ (
    .A(_3117_),
    .B(_3118_),
    .C(_3113_),
    .Y(_3121_)
);

NAND2X1 _9357_ (
    .A(vdd),
    .B(\X[3] [7]),
    .Y(_2715_)
);

FILL FILL_0__8612_ (
);

FILL FILL_3__9181_ (
);

DFFPOSX1 _13355_ (
    .D(\X[6] [1]),
    .CLK(clk_bF$buf2),
    .Q(\X[7] [1])
);

FILL FILL_1__6627_ (
);

FILL FILL_1__9099_ (
);

FILL FILL_0__9817_ (
);

FILL FILL_3__7914_ (
);

FILL FILL_2__8383_ (
);

FILL FILL_0__10771_ (
);

FILL FILL_0__10351_ (
);

AND2X2 _7843_ (
    .A(_1339_),
    .B(_1334_),
    .Y(_1357_)
);

OAI21X1 _7423_ (
    .A(_1575_),
    .B(_941_),
    .C(_942_),
    .Y(_943_)
);

NAND2X1 _7003_ (
    .A(_567_),
    .B(_595_),
    .Y(_596_)
);

FILL FILL_1__6380_ (
);

FILL FILL_2__13150_ (
);

FILL FILL_1__12983_ (
);

FILL FILL_3__11529_ (
);

FILL FILL_1__12563_ (
);

FILL FILL_1__12143_ (
);

FILL FILL_0__9990_ (
);

FILL FILL_0__11976_ (
);

FILL FILL_2__9588_ (
);

FILL FILL_0__9570_ (
);

FILL FILL_2__9168_ (
);

FILL FILL_0__9150_ (
);

AOI21X1 _11841_ (
    .A(_4864_),
    .B(_4882_),
    .C(_4960_),
    .Y(_4961_)
);

FILL FILL_0__11556_ (
);

NAND3X1 _11421_ (
    .A(_4611_),
    .B(_4612_),
    .C(_4610_),
    .Y(_4613_)
);

FILL FILL_0__11136_ (
);

OAI21X1 _11001_ (
    .A(_4124_),
    .B(_4199_),
    .C(_4128_),
    .Y(_4200_)
);

AND2X2 _8628_ (
    .A(_2060_),
    .B(_2063_),
    .Y(_2064_)
);

NAND2X1 _8208_ (
    .A(_1643_),
    .B(_1646_),
    .Y(_1650_)
);

FILL FILL_1__7585_ (
);

FILL FILL_1__7165_ (
);

FILL FILL_3__8452_ (
);

NAND2X1 _12626_ (
    .A(_5615_),
    .B(_5666_),
    .Y(_5667_)
);

FILL FILL_3__8032_ (
);

AOI21X1 _12206_ (
    .A(_5252_),
    .B(_5268_),
    .C(_5320_),
    .Y(_5321_)
);

FILL FILL_3__11282_ (
);

FILL FILL_2__10695_ (
);

FILL FILL_2__10275_ (
);

FILL FILL_1__9731_ (
);

FILL FILL_1__9311_ (
);

FILL FILL_3__9657_ (
);

FILL FILL_3__9237_ (
);

FILL FILL_0__6695_ (
);

INVX1 _8381_ (
    .A(_1819_),
    .Y(_1820_)
);

FILL FILL_2__7654_ (
);

FILL FILL_0__12094_ (
);

FILL FILL_2__12841_ (
);

FILL FILL_2__12421_ (
);

FILL FILL_2__12001_ (
);

OAI21X1 _9586_ (
    .A(_2887_),
    .B(_2940_),
    .C(_2883_),
    .Y(_2941_)
);

NAND2X1 _9166_ (
    .A(_2522_),
    .B(_2524_),
    .Y(_2526_)
);

FILL FILL_1__11834_ (
);

FILL FILL_1__11414_ (
);

FILL FILL_0__8841_ (
);

FILL FILL_2__8859_ (
);

FILL FILL_0__8421_ (
);

FILL FILL_2__8439_ (
);

FILL FILL_0__10827_ (
);

FILL FILL_0__10407_ (
);

FILL FILL_0__8001_ (
);

FILL FILL_2__8019_ (
);

FILL FILL_0__13299_ (
);

OAI21X1 _13164_ (
    .A(_6173_),
    .B(_6180_),
    .C(_6179_),
    .Y(_6196_)
);

FILL FILL_2__9800_ (
);

FILL FILL_1__6856_ (
);

FILL FILL_1__6436_ (
);

FILL FILL_2__13206_ (
);

FILL FILL_1__12619_ (
);

FILL FILL_0__9626_ (
);

FILL FILL_0__9206_ (
);

FILL FILL_3__10973_ (
);

FILL FILL_3__10133_ (
);

FILL FILL_2__8192_ (
);

FILL FILL_0__10580_ (
);

FILL FILL_0__10160_ (
);

FILL FILL_3__8928_ (
);

NAND2X1 _7652_ (
    .A(_1169_),
    .B(_1164_),
    .Y(_1170_)
);

DFFPOSX1 _7232_ (
    .D(Yin[9]),
    .CLK(clk_bF$buf41),
    .Q(\u_fir_pe0.rYin [9])
);

NAND2X1 _10289_ (
    .A(_3562_),
    .B(_3566_),
    .Y(_3984_[8])
);

FILL FILL_2__6925_ (
);

FILL FILL_3__11758_ (
);

FILL FILL_2__6505_ (
);

FILL FILL_1__12792_ (
);

FILL FILL_1__12372_ (
);

FILL FILL_2__9397_ (
);

FILL FILL_0__11785_ (
);

NOR2X1 _11650_ (
    .A(_5552_),
    .B(_5560_),
    .Y(_5562_)
);

FILL FILL_0__11365_ (
);

NAND3X1 _11230_ (
    .A(_4367_),
    .B(_4422_),
    .C(_4426_),
    .Y(_4427_)
);

INVX1 _8857_ (
    .A(_2274_),
    .Y(_2280_)
);

NAND3X1 _8437_ (
    .A(_1803_),
    .B(_1871_),
    .C(_1872_),
    .Y(_1876_)
);

INVX1 _8017_ (
    .A(\u_fir_pe1.rYin [10]),
    .Y(_1521_)
);

FILL FILL_1__7394_ (
);

FILL FILL_1__13157_ (
);

FILL FILL_3__8681_ (
);

NAND3X1 _12855_ (
    .A(_5890_),
    .B(_5892_),
    .C(_5891_),
    .Y(_5893_)
);

OR2X2 _12435_ (
    .A(_5531_),
    .B(_5537_),
    .Y(_5539_)
);

NAND3X1 _12015_ (
    .A(_5131_),
    .B(_5132_),
    .C(_5130_),
    .Y(_5133_)
);

FILL FILL_1__8599_ (
);

FILL FILL_1__8179_ (
);

FILL FILL_3__11091_ (
);

FILL FILL_2__10084_ (
);

FILL FILL_1__9960_ (
);

FILL FILL_1__9540_ (
);

FILL FILL_1__9120_ (
);

FILL FILL_3__9466_ (
);

AOI22X1 _8190_ (
    .A(vdd),
    .B(\X[2] [1]),
    .C(gnd),
    .D(\X[2] [2]),
    .Y(_1632_)
);

FILL FILL_2__7883_ (
);

FILL FILL_2__7463_ (
);

FILL FILL_2__7043_ (
);

FILL FILL_2__11289_ (
);

AOI22X1 _6923_ (
    .A(Xin_5_bF$buf3),
    .B(gnd),
    .C(_477_),
    .D(_478_),
    .Y(_518_)
);

NAND3X1 _6503_ (
    .A(_95_),
    .B(_91_),
    .C(_97_),
    .Y(_104_)
);

FILL FILL_2__12650_ (
);

FILL FILL_2__12230_ (
);

FILL FILL_0__7289_ (
);

NAND3X1 _9395_ (
    .A(_2751_),
    .B(_2752_),
    .C(_2750_),
    .Y(_2753_)
);

FILL FILL_3__10609_ (
);

FILL FILL_1__11643_ (
);

FILL FILL_1__11223_ (
);

FILL FILL_0__8650_ (
);

FILL FILL_2__8668_ (
);

FILL FILL_0__8230_ (
);

FILL FILL_2__8248_ (
);

FILL FILL_0__10636_ (
);

NAND2X1 _10921_ (
    .A(_4120_),
    .B(_4119_),
    .Y(_4121_)
);

NAND3X1 _10501_ (
    .A(_3565_),
    .B(_3638_),
    .C(_3744_),
    .Y(_3775_)
);

FILL FILL_0__10216_ (
);

DFFPOSX1 _13393_ (
    .D(_6375_[15]),
    .CLK(clk_bF$buf56),
    .Q(\u_fir_pe7.mul [15])
);

AOI21X1 _7708_ (
    .A(_1140_),
    .B(_1146_),
    .C(_1221_),
    .Y(_1225_)
);

FILL FILL_1__6665_ (
);

FILL FILL_2__13015_ (
);

FILL FILL_1__12848_ (
);

FILL FILL_1__12428_ (
);

FILL FILL_1__12008_ (
);

FILL FILL_0__9435_ (
);

FILL FILL_3__7532_ (
);

FILL FILL_0__9015_ (
);

INVX1 _11706_ (
    .A(_4814_),
    .Y(_4828_)
);

FILL FILL_3__10362_ (
);

FILL FILL_1__8811_ (
);

FILL FILL_3__8317_ (
);

OAI22X1 _7881_ (
    .A(_941_),
    .B(_1259_),
    .C(_1102_),
    .D(_1032_),
    .Y(_1394_)
);

AND2X2 _7461_ (
    .A(_931_),
    .B(_932_),
    .Y(_981_)
);

INVX1 _7041_ (
    .A(_24_),
    .Y(_791_[0])
);

OAI21X1 _10098_ (
    .A(_3300_),
    .B(_3377_),
    .C(_3294_),
    .Y(_3378_)
);

FILL FILL_3__11987_ (
);

FILL FILL_2__6734_ (
);

FILL FILL_3__11147_ (
);

FILL FILL_1__12181_ (
);

FILL FILL_0__11174_ (
);

FILL FILL_2__11921_ (
);

FILL FILL_2__11501_ (
);

NAND2X1 _8666_ (
    .A(_1971_),
    .B(_2044_),
    .Y(_2102_)
);

NAND2X1 _8246_ (
    .A(gnd),
    .B(\X[2] [3]),
    .Y(_1687_)
);

FILL FILL_1__10914_ (
);

FILL FILL_0__7921_ (
);

FILL FILL_2__7939_ (
);

FILL FILL_2__7519_ (
);

FILL FILL_0__7501_ (
);

FILL FILL_0__12799_ (
);

NAND3X1 _12664_ (
    .A(_5699_),
    .B(_5704_),
    .C(_5646_),
    .Y(_5705_)
);

FILL FILL_0__12379_ (
);

NAND2X1 _12244_ (
    .A(_5354_),
    .B(_5357_),
    .Y(_5358_)
);

FILL FILL_2__12706_ (
);

FILL FILL_0__13320_ (
);

FILL FILL_0__8706_ (
);

FILL FILL_3__6803_ (
);

NAND3X1 _13029_ (
    .A(_5986_),
    .B(_6064_),
    .C(_5994_),
    .Y(_6065_)
);

FILL FILL_2__7692_ (
);

FILL FILL_2__7272_ (
);

FILL FILL_2__11098_ (
);

INVX1 _6732_ (
    .A(_324_),
    .Y(_330_)
);

FILL FILL_0__7098_ (
);

FILL FILL_1__11872_ (
);

FILL FILL_1__11452_ (
);

FILL FILL_1__11032_ (
);

FILL FILL_2__8897_ (
);

FILL FILL_2__8477_ (
);

FILL FILL_0__10865_ (
);

DFFPOSX1 _10730_ (
    .D(\X[4] [7]),
    .CLK(clk_bF$buf45),
    .Q(\X[5] [7])
);

FILL FILL_0__10445_ (
);

FILL FILL_2__8057_ (
);

AND2X2 _10310_ (
    .A(_3320_),
    .B(_3509_),
    .Y(_3587_)
);

FILL FILL_0__10025_ (
);

AOI21X1 _7937_ (
    .A(_1437_),
    .B(_1442_),
    .C(_1438_),
    .Y(_1444_)
);

OAI21X1 _7517_ (
    .A(_953_),
    .B(_957_),
    .C(_956_),
    .Y(_1036_)
);

FILL FILL_1__6894_ (
);

FILL FILL_1__6474_ (
);

FILL FILL_2__13244_ (
);

FILL FILL_1__12657_ (
);

FILL FILL_1__12237_ (
);

FILL FILL_0__9664_ (
);

FILL FILL_3__7761_ (
);

FILL FILL_0__9244_ (
);

OAI21X1 _11935_ (
    .A(_5040_),
    .B(_5044_),
    .C(_5047_),
    .Y(_5054_)
);

NOR2X1 _11515_ (
    .A(_4698_),
    .B(_4697_),
    .Y(_4699_)
);

FILL FILL_1__7679_ (
);

FILL FILL_3__10591_ (
);

FILL FILL_1__7259_ (
);

FILL FILL_1__8620_ (
);

FILL FILL_1__8200_ (
);

FILL FILL_3__8546_ (
);

NAND2X1 _7690_ (
    .A(vdd),
    .B(\X[1] [7]),
    .Y(_1207_)
);

FILL FILL_1_BUFX2_insert80 (
);

NAND2X1 _7270_ (
    .A(_1517_),
    .B(_1581_),
    .Y(_1582_)
);

FILL FILL_1_BUFX2_insert81 (
);

FILL FILL_1_BUFX2_insert82 (
);

FILL FILL_1_BUFX2_insert83 (
);

FILL FILL_1_BUFX2_insert84 (
);

FILL FILL_1_BUFX2_insert85 (
);

FILL FILL_1_BUFX2_insert86 (
);

FILL FILL_1_BUFX2_insert87 (
);

FILL FILL_1_BUFX2_insert88 (
);

FILL FILL_1_BUFX2_insert89 (
);

FILL FILL_2__6963_ (
);

FILL FILL_2__6543_ (
);

FILL FILL_3__11376_ (
);

FILL FILL_2__10789_ (
);

FILL FILL_2__10369_ (
);

FILL FILL_1__9825_ (
);

FILL FILL_1__9405_ (
);

FILL FILL_0_CLKBUF1_insert60 (
);

FILL FILL_0_CLKBUF1_insert61 (
);

FILL FILL_0_CLKBUF1_insert62 (
);

FILL FILL_2__11730_ (
);

FILL FILL_0_CLKBUF1_insert63 (
);

FILL FILL_0_CLKBUF1_insert64 (
);

FILL FILL_0__6789_ (
);

FILL FILL_2__11310_ (
);

FILL FILL_0_CLKBUF1_insert65 (
);

INVX1 _8895_ (
    .A(\u_fir_pe2.mul [10]),
    .Y(_2319_)
);

INVX1 _8475_ (
    .A(gnd),
    .Y(_1913_)
);

FILL FILL_0_CLKBUF1_insert66 (
);

FILL FILL_0_CLKBUF1_insert67 (
);

NOR2X1 _8055_ (
    .A(_1556_),
    .B(_1558_),
    .Y(_1559_)
);

FILL FILL_0_CLKBUF1_insert68 (
);

FILL FILL_0_CLKBUF1_insert69 (
);

FILL FILL_1__10303_ (
);

FILL FILL_2__7748_ (
);

FILL FILL_0__7730_ (
);

FILL FILL_2__7328_ (
);

FILL FILL_0__7310_ (
);

FILL FILL_1__13195_ (
);

AOI21X1 _12893_ (
    .A(_5930_),
    .B(_5925_),
    .C(_5894_),
    .Y(_5931_)
);

FILL FILL_0__12188_ (
);

DFFPOSX1 _12473_ (
    .D(_5572_[12]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[12])
);

NAND2X1 _12053_ (
    .A(gnd),
    .B(_5169_),
    .Y(_5170_)
);

FILL FILL_3__13102_ (
);

FILL FILL_2__12935_ (
);

FILL FILL_1__11928_ (
);

FILL FILL_1__11508_ (
);

FILL FILL_0__8935_ (
);

FILL FILL_0__8515_ (
);

FILL FILL254250x75750 (
);

FILL FILL_3__9084_ (
);

NAND2X1 _13258_ (
    .A(_6278_),
    .B(_6281_),
    .Y(_6282_)
);

FILL FILL_2__7081_ (
);

NAND2X1 _6961_ (
    .A(_554_),
    .B(_555_),
    .Y(_796_[11])
);

AND2X2 _6541_ (
    .A(Xin[2]),
    .B(gnd),
    .Y(_141_)
);

FILL FILL253950x126150 (
);

FILL FILL_1__11681_ (
);

FILL FILL_3__10227_ (
);

FILL FILL_1__11261_ (
);

FILL FILL_2__8286_ (
);

FILL FILL_0__10674_ (
);

FILL FILL_0__10254_ (
);

INVX1 _7746_ (
    .A(_1261_),
    .Y(_1262_)
);

NAND3X1 _7326_ (
    .A(_837_),
    .B(_841_),
    .C(_843_),
    .Y(_848_)
);

FILL FILL_2__13053_ (
);

FILL FILL_1__12886_ (
);

FILL FILL_1__12046_ (
);

FILL FILL_0__9893_ (
);

FILL FILL_3__7990_ (
);

FILL FILL_0__9473_ (
);

FILL FILL_0__11879_ (
);

FILL FILL_0__9053_ (
);

NAND2X1 _11744_ (
    .A(gnd),
    .B(\X[7] [2]),
    .Y(_4865_)
);

FILL FILL_0__11459_ (
);

FILL FILL_3__7150_ (
);

FILL FILL_0__11039_ (
);

INVX1 _11324_ (
    .A(_4516_),
    .Y(_4519_)
);

FILL FILL_0__12820_ (
);

FILL FILL_0__12400_ (
);

FILL FILL_1__7488_ (
);

FILL FILL_1__7068_ (
);

FILL FILL_3__8775_ (
);

NAND2X1 _12949_ (
    .A(_5985_),
    .B(_5982_),
    .Y(_5986_)
);

INVX1 _12529_ (
    .A(_6360_),
    .Y(_6361_)
);

AOI21X1 _12109_ (
    .A(_5082_),
    .B(_5147_),
    .C(_5225_),
    .Y(_5226_)
);

FILL FILL_2__6772_ (
);

FILL FILL_2__10598_ (
);

FILL FILL_2__10178_ (
);

FILL FILL_1__9634_ (
);

FILL FILL_1__9214_ (
);

FILL FILL_0__6598_ (
);

AND2X2 _8284_ (
    .A(_1724_),
    .B(_1720_),
    .Y(_2390_[5])
);

FILL FILL_1__10952_ (
);

FILL FILL_1__10532_ (
);

FILL FILL_1__10112_ (
);

FILL FILL_2__7977_ (
);

FILL FILL_2__7557_ (
);

FILL FILL_2__7137_ (
);

NAND3X1 _12282_ (
    .A(_5366_),
    .B(_5394_),
    .C(_5393_),
    .Y(_5395_)
);

FILL FILL_3__13331_ (
);

FILL FILL_2__12744_ (
);

FILL FILL_2__12324_ (
);

NOR2X1 _9489_ (
    .A(_2764_),
    .B(_2844_),
    .Y(_2845_)
);

NAND3X1 _9069_ (
    .A(_2425_),
    .B(_2430_),
    .C(_2428_),
    .Y(_2431_)
);

FILL FILL_1__11737_ (
);

FILL FILL_1__11317_ (
);

FILL FILL_0__8744_ (
);

FILL FILL_0__8324_ (
);

FILL FILL_3__6421_ (
);

NAND3X1 _13067_ (
    .A(_6099_),
    .B(_6100_),
    .C(_6101_),
    .Y(_6102_)
);

FILL FILL_2__9703_ (
);

FILL FILL_1__6759_ (
);

FILL FILL_2__13109_ (
);

FILL FILL_1__7700_ (
);

FILL FILL_0__9949_ (
);

FILL FILL_0__9529_ (
);

FILL FILL_3__7626_ (
);

FILL FILL_0__9109_ (
);

AOI21X1 _6770_ (
    .A(_278_),
    .B(_277_),
    .C(_209_),
    .Y(_368_)
);

FILL FILL_3__10876_ (
);

FILL FILL_3__10456_ (
);

FILL FILL_1__11490_ (
);

FILL FILL_1__11070_ (
);

FILL FILL_0__10483_ (
);

FILL FILL_0__10063_ (
);

FILL FILL_1__8905_ (
);

FILL FILL_2__10810_ (
);

INVX1 _7975_ (
    .A(\u_fir_pe1.rYin [7]),
    .Y(_1478_)
);

NAND3X1 _7555_ (
    .A(_1068_),
    .B(_1067_),
    .C(_1069_),
    .Y(_1074_)
);

NOR2X1 _7135_ (
    .A(_715_),
    .B(_709_),
    .Y(_718_)
);

FILL FILL_2__13282_ (
);

FILL FILL_0__6810_ (
);

FILL FILL_2__6828_ (
);

FILL FILL_2__6408_ (
);

FILL FILL_1__12695_ (
);

FILL FILL_1__12275_ (
);

FILL FILL_0__9282_ (
);

AND2X2 _11973_ (
    .A(_5089_),
    .B(_5088_),
    .Y(_5091_)
);

FILL FILL_0__11688_ (
);

INVX1 _11553_ (
    .A(\u_fir_pe5.mul [13]),
    .Y(_4737_)
);

FILL FILL_0__11268_ (
);

OAI21X1 _11133_ (
    .A(_4326_),
    .B(_4330_),
    .C(_4302_),
    .Y(_4331_)
);

FILL FILL_3__12602_ (
);

FILL FILL_1__7297_ (
);

INVX1 _9701_ (
    .A(\u_fir_pe3.mul [4]),
    .Y(_3047_)
);

NAND3X1 _12758_ (
    .A(_5790_),
    .B(_5796_),
    .C(_5795_),
    .Y(_5797_)
);

FILL FILL_3__8164_ (
);

NAND2X1 _12338_ (
    .A(_5441_),
    .B(_5443_),
    .Y(_5444_)
);

FILL FILL_0__13414_ (
);

FILL FILL_2__6581_ (
);

FILL FILL_1__9443_ (
);

FILL FILL_1__9023_ (
);

DFFPOSX1 _8093_ (
    .D(\X[1] [1]),
    .CLK(clk_bF$buf21),
    .Q(\X[2] [1])
);

FILL FILL_1__10341_ (
);

FILL FILL_2__7786_ (
);

FILL FILL_2__7366_ (
);

FILL FILL_3__12199_ (
);

NAND3X1 _12091_ (
    .A(_5177_),
    .B(_5205_),
    .C(_5207_),
    .Y(_5208_)
);

NAND3X1 _6826_ (
    .A(_415_),
    .B(_422_),
    .C(_397_),
    .Y(_423_)
);

NAND3X1 _6406_ (
    .A(_740_),
    .B(_8_),
    .C(_6_),
    .Y(_9_)
);

FILL FILL_2__12973_ (
);

FILL FILL_2__12553_ (
);

FILL FILL_2__12133_ (
);

NAND3X1 _9298_ (
    .A(_2651_),
    .B(_2650_),
    .C(_2652_),
    .Y(_2657_)
);

FILL FILL_1__11966_ (
);

FILL FILL_1__11546_ (
);

FILL FILL_1__11126_ (
);

FILL FILL_0__8553_ (
);

FILL FILL_0__10959_ (
);

FILL FILL_3__6650_ (
);

FILL FILL_0__8133_ (
);

FILL FILL_0__10539_ (
);

NAND3X1 _10824_ (
    .A(gnd),
    .B(\X[5] [2]),
    .C(_4016_),
    .Y(_4026_)
);

NAND3X1 _10404_ (
    .A(_3675_),
    .B(_3679_),
    .C(_3649_),
    .Y(_3680_)
);

FILL FILL_0__10119_ (
);

OAI21X1 _13296_ (
    .A(_6318_),
    .B(_6301_),
    .C(_6317_),
    .Y(_6320_)
);

FILL FILL_2__9932_ (
);

FILL FILL_0__11900_ (
);

FILL FILL_2__9512_ (
);

FILL FILL_1__6988_ (
);

FILL FILL_1__6568_ (
);

FILL FILL_0__9758_ (
);

FILL FILL_3__7855_ (
);

FILL FILL_0__9338_ (
);

FILL FILL_3__7435_ (
);

DFFPOSX1 _11609_ (
    .D(\Y[5] [1]),
    .CLK(clk_bF$buf6),
    .Q(\u_fir_pe5.rYin [1])
);

FILL FILL_3__7015_ (
);

FILL FILL_3__10685_ (
);

FILL FILL_0__10292_ (
);

FILL FILL_1__8714_ (
);

NAND2X1 _7784_ (
    .A(_1292_),
    .B(_1298_),
    .Y(_1300_)
);

NAND2X1 _7364_ (
    .A(_833_),
    .B(_884_),
    .Y(_885_)
);

FILL FILL_2__13091_ (
);

FILL FILL_2__6637_ (
);

FILL FILL_1__12084_ (
);

FILL FILL_0__9091_ (
);

INVX1 _11782_ (
    .A(_4802_),
    .Y(_4903_)
);

FILL FILL_0__11497_ (
);

FILL FILL_0__11077_ (
);

NAND2X1 _11362_ (
    .A(_4550_),
    .B(_4554_),
    .Y(_4556_)
);

FILL FILL_1__9919_ (
);

FILL FILL_3__12831_ (
);

FILL FILL_3__12411_ (
);

FILL FILL_2__11824_ (
);

FILL FILL_2__11404_ (
);

DFFPOSX1 _8989_ (
    .D(\Y[2] [12]),
    .CLK(clk_bF$buf10),
    .Q(\u_fir_pe2.rYin [12])
);

NAND2X1 _8569_ (
    .A(vdd),
    .B(\X[2] [7]),
    .Y(_2006_)
);

NAND2X1 _8149_ (
    .A(vdd),
    .B(\X[2] [3]),
    .Y(_2381_)
);

FILL FILL_1__10817_ (
);

FILL FILL_0__7824_ (
);

NAND2X1 _9930_ (
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3212_)
);

FILL FILL_0__7404_ (
);

AND2X2 _9510_ (
    .A(_2864_),
    .B(_2807_),
    .Y(_2866_)
);

FILL FILL_1__13289_ (
);

OAI21X1 _12987_ (
    .A(_6014_),
    .B(_6013_),
    .C(_5964_),
    .Y(_6024_)
);

FILL FILL_3__8393_ (
);

NAND2X1 _12567_ (
    .A(\X[6] [0]),
    .B(vdd),
    .Y(_5609_)
);

AOI21X1 _12147_ (
    .A(vdd),
    .B(\X[7] [6]),
    .C(_5194_),
    .Y(_5263_)
);

FILL FILL_2__12609_ (
);

FILL FILL_0__13223_ (
);

FILL FILL_2__6390_ (
);

FILL FILL_0__8609_ (
);

FILL FILL_1__9672_ (
);

FILL FILL_1__9252_ (
);

FILL FILL_3__9598_ (
);

FILL FILL_3__9178_ (
);

FILL FILL_1__10990_ (
);

FILL FILL_1__10570_ (
);

FILL FILL_1__10150_ (
);

FILL FILL_2__7595_ (
);

FILL FILL_2__7175_ (
);

OAI21X1 _6635_ (
    .A(_15_),
    .B(_233_),
    .C(_228_),
    .Y(_234_)
);

FILL FILL_2__12782_ (
);

FILL FILL_2__12362_ (
);

FILL FILL_1__11775_ (
);

FILL FILL_1__11355_ (
);

FILL FILL_0__8782_ (
);

FILL FILL_0__8362_ (
);

FILL FILL_0__10768_ (
);

FILL FILL_0__10348_ (
);

INVX1 _10633_ (
    .A(_3880_),
    .Y(_3896_)
);

OAI21X1 _10213_ (
    .A(_3410_),
    .B(_3490_),
    .C(_3459_),
    .Y(_3491_)
);

FILL FILL_2__9741_ (
);

FILL FILL_2__9321_ (
);

FILL FILL_1__6797_ (
);

FILL FILL_2__13147_ (
);

FILL FILL_0__9987_ (
);

FILL FILL_0__9567_ (
);

FILL FILL_0__9147_ (
);

NAND3X1 _11838_ (
    .A(_4955_),
    .B(_4957_),
    .C(_4956_),
    .Y(_4958_)
);

NAND2X1 _11418_ (
    .A(_4609_),
    .B(_4573_),
    .Y(_4610_)
);

FILL FILL_0__12914_ (
);

FILL FILL_3__10074_ (
);

FILL FILL_1__8943_ (
);

FILL FILL_1__8523_ (
);

FILL FILL_3__8869_ (
);

FILL FILL_3__8029_ (
);

NAND3X1 _7593_ (
    .A(_1108_),
    .B(_1110_),
    .C(_1109_),
    .Y(_1111_)
);

OR2X2 _7173_ (
    .A(_749_),
    .B(_755_),
    .Y(_757_)
);

FILL FILL_2__6866_ (
);

FILL FILL_3__11699_ (
);

FILL FILL_2__6446_ (
);

DFFPOSX1 _11591_ (
    .D(_4775_[7]),
    .CLK(clk_bF$buf48),
    .Q(\Y[6] [7])
);

OAI21X1 _11171_ (
    .A(_4289_),
    .B(_4293_),
    .C(_4298_),
    .Y(_4368_)
);

FILL FILL_1__9728_ (
);

FILL FILL_1__9308_ (
);

FILL FILL_3__12220_ (
);

FILL FILL_2__11213_ (
);

INVX1 _8798_ (
    .A(\u_fir_pe2.mul [1]),
    .Y(_2227_)
);

AOI21X1 _8378_ (
    .A(_1756_),
    .B(_1760_),
    .C(_1749_),
    .Y(_1817_)
);

FILL FILL_1__10626_ (
);

FILL FILL_1__10206_ (
);

FILL FILL_0__7633_ (
);

FILL FILL_1__13098_ (
);

OAI21X1 _12796_ (
    .A(_5827_),
    .B(_5834_),
    .C(_5819_),
    .Y(_5835_)
);

OAI21X1 _12376_ (
    .A(_5463_),
    .B(_5464_),
    .C(_5478_),
    .Y(_5479_)
);

FILL FILL_2__12838_ (
);

FILL FILL_2__12418_ (
);

FILL FILL_0__13032_ (
);

FILL FILL_0__8838_ (
);

FILL FILL_0__8418_ (
);

FILL FILL_3__6515_ (
);

FILL FILL_1__9481_ (
);

FILL FILL_1__9061_ (
);

FILL FILL253350x10950 (
);

OAI21X1 _6864_ (
    .A(_386_),
    .B(_390_),
    .C(_388_),
    .Y(_460_)
);

INVX1 _6444_ (
    .A(_32_),
    .Y(_46_)
);

FILL FILL_2__12591_ (
);

FILL FILL_2__12171_ (
);

FILL FILL_1__11164_ (
);

FILL FILL_0__8591_ (
);

FILL FILL_0__10997_ (
);

FILL FILL_2__8189_ (
);

FILL FILL_0__8171_ (
);

FILL FILL_0__10577_ (
);

NAND3X1 _10862_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf2 ),
    .C(_4060_),
    .Y(_4063_)
);

NAND3X1 _10442_ (
    .A(_3713_),
    .B(_3716_),
    .C(_3670_),
    .Y(_3717_)
);

FILL FILL_0__10157_ (
);

NAND3X1 _10022_ (
    .A(_3300_),
    .B(_3301_),
    .C(_3302_),
    .Y(_3303_)
);

FILL FILL_3__11911_ (
);

FILL FILL_2__10904_ (
);

FILL FILL_2__9970_ (
);

FILL FILL_2__9550_ (
);

FILL FILL_2__9130_ (
);

NAND3X1 _7649_ (
    .A(_1097_),
    .B(_1161_),
    .C(_1162_),
    .Y(_1167_)
);

DFFPOSX1 _7229_ (
    .D(Yin[6]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [6])
);

FILL FILL_0__6904_ (
);

FILL FILL_1__12789_ (
);

FILL FILL_1__12369_ (
);

FILL FILL_0__9796_ (
);

FILL FILL_0__9376_ (
);

FILL FILL_3__7473_ (
);

NOR2X1 _11647_ (
    .A(_5532_),
    .B(_5522_),
    .Y(_5542_)
);

INVX1 _11227_ (
    .A(_4416_),
    .Y(_4424_)
);

FILL FILL_1__13310_ (
);

FILL FILL_0__12723_ (
);

FILL FILL_0__12303_ (
);

FILL FILL_1__8752_ (
);

FILL FILL_1__8332_ (
);

FILL FILL_3__8258_ (
);

FILL FILL_2__6675_ (
);

FILL FILL_3__11088_ (
);

FILL FILL_1__9957_ (
);

FILL FILL_1__9537_ (
);

FILL FILL_1__9117_ (
);

FILL FILL_2__11862_ (
);

FILL FILL_2__11442_ (
);

FILL FILL_2__11022_ (
);

AND2X2 _8187_ (
    .A(gnd),
    .B(\X[2] [1]),
    .Y(_1629_)
);

FILL FILL_1__10855_ (
);

FILL FILL_1__10435_ (
);

FILL FILL_1__10015_ (
);

FILL FILL_0__7862_ (
);

FILL FILL_0__7442_ (
);

FILL FILL_0__7022_ (
);

AOI22X1 _12185_ (
    .A(\X[7]_5_bF$buf0 ),
    .B(gnd),
    .C(_5259_),
    .D(_5260_),
    .Y(_5300_)
);

FILL FILL_2__8821_ (
);

FILL FILL_2__8401_ (
);

FILL FILL_2__12647_ (
);

FILL FILL_2__12227_ (
);

FILL FILL_0__13261_ (
);

FILL FILL_0__8647_ (
);

FILL FILL_3__6744_ (
);

FILL FILL_0__8227_ (
);

OAI21X1 _10918_ (
    .A(_4695_),
    .B(_4117_),
    .C(_4062_),
    .Y(_4118_)
);

FILL FILL_1__9290_ (
);

FILL FILL_2__9606_ (
);

FILL FILL_2_CLKBUF1_insert12 (
);

FILL FILL_2_CLKBUF1_insert13 (
);

FILL FILL_2_CLKBUF1_insert14 (
);

FILL FILL_2_CLKBUF1_insert15 (
);

FILL FILL_2_CLKBUF1_insert16 (
);

FILL FILL_2_CLKBUF1_insert17 (
);

FILL FILL_2_CLKBUF1_insert18 (
);

FILL FILL_2_CLKBUF1_insert19 (
);

FILL FILL_1__7603_ (
);

FILL FILL_3__7949_ (
);

FILL FILL_3__7529_ (
);

FILL FILL_3__7109_ (
);

OAI21X1 _6673_ (
    .A(_258_),
    .B(_262_),
    .C(_265_),
    .Y(_272_)
);

FILL FILL_1__11393_ (
);

FILL FILL_0__10386_ (
);

NAND2X1 _10671_ (
    .A(_3934_),
    .B(_3929_),
    .Y(_3935_)
);

AOI21X1 _10251_ (
    .A(_3524_),
    .B(_3528_),
    .C(_3510_),
    .Y(_3529_)
);

FILL FILL_1__8808_ (
);

FILL FILL_3__11720_ (
);

FILL FILL_3__11300_ (
);

INVX1 _7878_ (
    .A(_1390_),
    .Y(_1391_)
);

AOI21X1 _7458_ (
    .A(_968_),
    .B(_964_),
    .C(_949_),
    .Y(_978_)
);

OAI21X1 _7038_ (
    .A(_616_),
    .B(_615_),
    .C(_627_),
    .Y(_629_)
);

FILL FILL_2__13185_ (
);

FILL FILL_0__6713_ (
);

FILL FILL_1__12598_ (
);

FILL FILL_1__12178_ (
);

FILL FILL_0__9185_ (
);

INVX1 _11876_ (
    .A(_4994_),
    .Y(_4995_)
);

NOR2X1 _11456_ (
    .A(_4640_),
    .B(_4641_),
    .Y(_4642_)
);

AOI21X1 _11036_ (
    .A(_4232_),
    .B(_4234_),
    .C(_4231_),
    .Y(_4235_)
);

FILL FILL_3__12925_ (
);

FILL FILL_2__11918_ (
);

FILL FILL_0__12952_ (
);

FILL FILL_0__12532_ (
);

FILL FILL_0__12112_ (
);

FILL FILL_0__7918_ (
);

NOR2X1 _9604_ (
    .A(_2535_),
    .B(_2696_),
    .Y(_2958_)
);

FILL FILL_1__8561_ (
);

FILL FILL_1__8141_ (
);

FILL FILL_3__8487_ (
);

FILL FILL_3__8067_ (
);

FILL FILL_0__13317_ (
);

FILL FILL_2__6484_ (
);

FILL FILL_1__9766_ (
);

FILL FILL_1__9346_ (
);

FILL FILL_2__11671_ (
);

FILL FILL_2__11251_ (
);

FILL FILL_1__10664_ (
);

FILL FILL_1__10244_ (
);

FILL FILL_0__7671_ (
);

FILL FILL_2__7689_ (
);

FILL FILL_2__7269_ (
);

FILL FILL_2__8630_ (
);

FILL FILL_2__8210_ (
);

FILL FILL_3__13043_ (
);

AND2X2 _6729_ (
    .A(gnd),
    .B(Xin_5_bF$buf0),
    .Y(_327_)
);

FILL FILL_2__12876_ (
);

FILL FILL_2__12456_ (
);

FILL FILL_2__12036_ (
);

FILL FILL_0__13070_ (
);

FILL FILL_1__11869_ (
);

FILL FILL_1__11449_ (
);

FILL FILL_1__11029_ (
);

FILL FILL_0__8876_ (
);

FILL FILL_3__6973_ (
);

FILL FILL_0__8456_ (
);

DFFPOSX1 _10727_ (
    .D(\X[4] [4]),
    .CLK(clk_bF$buf7),
    .Q(\X[5] [4])
);

FILL FILL_0__8036_ (
);

AOI21X1 _10307_ (
    .A(_3527_),
    .B(_3526_),
    .C(_3511_),
    .Y(_3584_)
);

FILL FILL_1__12810_ (
);

AOI21X1 _13199_ (
    .A(_6219_),
    .B(_6224_),
    .C(_6220_),
    .Y(_6226_)
);

FILL FILL_2__9415_ (
);

FILL FILL_0__11803_ (
);

FILL FILL_1__7832_ (
);

FILL FILL_1__7412_ (
);

NAND2X1 _6482_ (
    .A(gnd),
    .B(Xin[2]),
    .Y(_83_)
);

FILL FILL_3__10168_ (
);

NOR2X1 _10480_ (
    .A(_3661_),
    .B(_3714_),
    .Y(_3754_)
);

FILL FILL_0__10195_ (
);

AND2X2 _10060_ (
    .A(_3335_),
    .B(_3339_),
    .Y(_3340_)
);

FILL FILL_1__8617_ (
);

FILL FILL_2__10942_ (
);

FILL FILL_2__10522_ (
);

FILL FILL_2__10102_ (
);

NAND2X1 _7687_ (
    .A(_1203_),
    .B(_1200_),
    .Y(_1204_)
);

INVX1 _7267_ (
    .A(_1578_),
    .Y(_1579_)
);

FILL FILL_3__9904_ (
);

FILL FILL_0__6942_ (
);

FILL FILL_0__6522_ (
);

NAND2X1 _11685_ (
    .A(\X[7] [4]),
    .B(gnd),
    .Y(_4807_)
);

FILL FILL_3__7091_ (
);

OAI22X1 _11265_ (
    .A(_4316_),
    .B(_4397_),
    .C(_4459_),
    .D(_4460_),
    .Y(_4461_)
);

FILL FILL_2__7901_ (
);

FILL FILL_3__12314_ (
);

FILL FILL_2__11727_ (
);

FILL FILL_0__12761_ (
);

FILL FILL_2__11307_ (
);

FILL FILL_0__12341_ (
);

FILL FILL_0__7727_ (
);

DFFPOSX1 _9833_ (
    .D(_3181_[3]),
    .CLK(clk_bF$buf0),
    .Q(\Y[4] [3])
);

FILL FILL_0__7307_ (
);

INVX1 _9413_ (
    .A(_2763_),
    .Y(_2770_)
);

FILL FILL_1__8790_ (
);

FILL FILL_1__8370_ (
);

FILL FILL_0__13126_ (
);

BUFX2 _13411_ (
    .A(_6377_[3]),
    .Y(Yout[3])
);

FILL FILL_3__6609_ (
);

FILL FILL_1__9995_ (
);

FILL FILL_1__9575_ (
);

FILL FILL_1__9155_ (
);

FILL FILL_2__11480_ (
);

FILL FILL_2__11060_ (
);

FILL FILL_1__10893_ (
);

FILL FILL_1__10473_ (
);

FILL FILL_1__10053_ (
);

FILL FILL_0__7480_ (
);

FILL FILL_2__7498_ (
);

FILL FILL_0__7060_ (
);

FILL FILL_2__7078_ (
);

FILL FILL_3__10800_ (
);

FILL FILL_3__13272_ (
);

INVX1 _6958_ (
    .A(_552_),
    .Y(_553_)
);

OAI21X1 _6538_ (
    .A(_102_),
    .B(_137_),
    .C(_96_),
    .Y(_138_)
);

FILL FILL_2__12685_ (
);

FILL FILL_2__12265_ (
);

FILL FILL_1__11678_ (
);

FILL FILL_1__11258_ (
);

FILL FILL_0__8685_ (
);

FILL FILL_0__8265_ (
);

OAI21X1 _10956_ (
    .A(_4154_),
    .B(_4155_),
    .C(_4153_),
    .Y(_4156_)
);

NAND2X1 _10536_ (
    .A(_3806_),
    .B(_3805_),
    .Y(_3808_)
);

INVX1 _10116_ (
    .A(_3390_),
    .Y(_3395_)
);

FILL FILL_2__9644_ (
);

FILL FILL_2__9224_ (
);

FILL FILL_1__7641_ (
);

FILL FILL_3__7567_ (
);

FILL FILL_1__13404_ (
);

FILL FILL_0__12817_ (
);

FILL FILL_3__10397_ (
);

FILL FILL_1__8846_ (
);

FILL FILL_1__8426_ (
);

FILL FILL_1__8006_ (
);

FILL FILL_2__10331_ (
);

NAND3X1 _7496_ (
    .A(_1008_),
    .B(_1014_),
    .C(_1013_),
    .Y(_1015_)
);

NAND2X1 _7076_ (
    .A(_659_),
    .B(_661_),
    .Y(_662_)
);

FILL FILL_3__9713_ (
);

FILL FILL_0__6751_ (
);

FILL FILL_2__6769_ (
);

NOR2X1 _11494_ (
    .A(_4675_),
    .B(_4676_),
    .Y(_4677_)
);

NAND3X1 _11074_ (
    .A(_4173_),
    .B(_4271_),
    .C(_4272_),
    .Y(_4273_)
);

FILL FILL_2__7710_ (
);

FILL FILL_3__12543_ (
);

FILL FILL_2__11956_ (
);

FILL FILL_0__12990_ (
);

FILL FILL_2__11536_ (
);

FILL FILL_0__12570_ (
);

FILL FILL_2__11116_ (
);

FILL FILL_0__12150_ (
);

FILL FILL_1__10949_ (
);

FILL FILL_1__10529_ (
);

FILL FILL_1__10109_ (
);

FILL FILL_0__7956_ (
);

FILL FILL_0__7536_ (
);

NAND2X1 _9642_ (
    .A(_2993_),
    .B(_2994_),
    .Y(_2995_)
);

FILL FILL_0__7116_ (
);

NAND3X1 _9222_ (
    .A(_2575_),
    .B(_2568_),
    .C(_2573_),
    .Y(_2582_)
);

AOI22X1 _12699_ (
    .A(vdd),
    .B(\X[6] [3]),
    .C(vdd),
    .D(\X[6] [4]),
    .Y(_5739_)
);

OAI21X1 _12279_ (
    .A(_5373_),
    .B(_5368_),
    .C(_5391_),
    .Y(_5392_)
);

FILL FILL_2__8915_ (
);

INVX1 _13220_ (
    .A(\u_fir_pe7.mul [5]),
    .Y(_6245_)
);

FILL FILL_1__6912_ (
);

FILL FILL_3__6838_ (
);

FILL FILL_1__9384_ (
);

FILL FILL_1__10282_ (
);

OAI21X1 _6767_ (
    .A(_356_),
    .B(_352_),
    .C(_359_),
    .Y(_365_)
);

FILL FILL_2__12074_ (
);

FILL FILL_1__11487_ (
);

FILL FILL_1__11067_ (
);

FILL FILL_0__8494_ (
);

FILL FILL_3__6591_ (
);

INVX1 _10765_ (
    .A(_4685_),
    .Y(_4695_)
);

FILL FILL_0__8074_ (
);

INVX1 _10345_ (
    .A(_3614_),
    .Y(_3622_)
);

FILL FILL_3__11814_ (
);

FILL FILL_2__10807_ (
);

FILL FILL_2__9453_ (
);

FILL FILL_0__11841_ (
);

FILL FILL_2__9033_ (
);

FILL FILL_0__11421_ (
);

FILL FILL_0__11001_ (
);

FILL FILL_2__13279_ (
);

FILL FILL_0__6807_ (
);

INVX1 _8913_ (
    .A(\u_fir_pe2.mul [12]),
    .Y(_2337_)
);

FILL FILL_1__7870_ (
);

FILL FILL_1__7450_ (
);

FILL FILL_1__7030_ (
);

FILL FILL_0__9699_ (
);

FILL FILL_3__7796_ (
);

FILL FILL_0__9279_ (
);

FILL FILL_1__13213_ (
);

NAND3X1 _12911_ (
    .A(_5879_),
    .B(_5943_),
    .C(_5944_),
    .Y(_5949_)
);

FILL FILL_0__12626_ (
);

FILL FILL_0__12206_ (
);

FILL FILL_1__8655_ (
);

FILL FILL_1__8235_ (
);

FILL FILL_2__10980_ (
);

FILL FILL_2__10560_ (
);

FILL FILL_2__10140_ (
);

FILL FILL_3__9942_ (
);

FILL FILL_3__9102_ (
);

FILL FILL_2__6998_ (
);

FILL FILL_0__6980_ (
);

FILL FILL_0__6560_ (
);

FILL FILL_2__6578_ (
);

FILL FILL_3__12772_ (
);

FILL FILL_3__12352_ (
);

FILL FILL_2__11765_ (
);

FILL FILL_2__11345_ (
);

FILL FILL_1__10338_ (
);

FILL FILL_0__7765_ (
);

DFFPOSX1 _9871_ (
    .D(_3183_[1]),
    .CLK(clk_bF$buf14),
    .Q(\u_fir_pe3.mul [1])
);

FILL FILL_0__7345_ (
);

INVX1 _9451_ (
    .A(\X[3] [4]),
    .Y(_2808_)
);

OR2X2 _9031_ (
    .A(_3122_),
    .B(_2393_),
    .Y(_2394_)
);

NAND3X1 _12088_ (
    .A(_5197_),
    .B(_5204_),
    .C(_5179_),
    .Y(_5205_)
);

FILL FILL_2__8724_ (
);

FILL FILL_2__8304_ (
);

FILL FILL_3__13137_ (
);

FILL FILL_0__13164_ (
);

FILL FILL_1__6721_ (
);

FILL FILL_1__9193_ (
);

FILL FILL_1__12904_ (
);

FILL FILL_2__9929_ (
);

FILL FILL_0__9911_ (
);

FILL FILL_2__9509_ (
);

FILL FILL_1__10091_ (
);

FILL FILL_1__7926_ (
);

FILL FILL_1__7506_ (
);

NOR2X1 _6996_ (
    .A(_589_),
    .B(_588_),
    .Y(_590_)
);

NAND3X1 _6576_ (
    .A(_173_),
    .B(_175_),
    .C(_174_),
    .Y(_176_)
);

FILL FILL_1__11296_ (
);

AOI21X1 _10994_ (
    .A(_4157_),
    .B(_4161_),
    .C(_4123_),
    .Y(_4193_)
);

NAND2X1 _10574_ (
    .A(_3840_),
    .B(_3835_),
    .Y(_3841_)
);

FILL FILL_0__10289_ (
);

AOI21X1 _10154_ (
    .A(_3432_),
    .B(_3431_),
    .C(_3428_),
    .Y(_3433_)
);

FILL FILL_2__9682_ (
);

FILL FILL_2__10616_ (
);

FILL FILL_2__9262_ (
);

FILL FILL_0__11650_ (
);

FILL FILL_0__11230_ (
);

FILL FILL_2__13088_ (
);

FILL FILL_0__6616_ (
);

OAI21X1 _8722_ (
    .A(_2124_),
    .B(_2118_),
    .C(_2128_),
    .Y(_2156_)
);

NAND3X1 _8302_ (
    .A(vdd),
    .B(\X[2] [6]),
    .C(_1739_),
    .Y(_1742_)
);

FILL FILL_0__9088_ (
);

NAND3X1 _11779_ (
    .A(_4808_),
    .B(_4895_),
    .C(_4896_),
    .Y(_4900_)
);

FILL FILL_3__7185_ (
);

NOR2X1 _11359_ (
    .A(_4552_),
    .B(_4551_),
    .Y(_4553_)
);

FILL FILL_3__12408_ (
);

FILL FILL_1__13022_ (
);

FILL FILL_0__12855_ (
);

AOI21X1 _12720_ (
    .A(_5750_),
    .B(_5746_),
    .C(_5731_),
    .Y(_5760_)
);

FILL FILL_0__12435_ (
);

FILL FILL_0__12015_ (
);

OAI21X1 _12300_ (
    .A(_5398_),
    .B(_5397_),
    .C(_5409_),
    .Y(_5411_)
);

INVX1 _9927_ (
    .A(_3209_),
    .Y(_3210_)
);

OAI21X1 _9507_ (
    .A(_2810_),
    .B(_2862_),
    .C(_2798_),
    .Y(_2863_)
);

FILL FILL_1__8884_ (
);

FILL FILL_1__8464_ (
);

FILL FILL_1__8044_ (
);

FILL FILL254250x190950 (
);

FILL FILL_3__9331_ (
);

FILL FILL_2__6387_ (
);

FILL FILL_1__9669_ (
);

FILL FILL_1__9249_ (
);

FILL FILL_3__12161_ (
);

FILL FILL_2__11994_ (
);

FILL FILL_2__11574_ (
);

FILL FILL_2__11154_ (
);

FILL FILL_1__10987_ (
);

FILL FILL_1__10567_ (
);

FILL FILL_1__10147_ (
);

FILL FILL_0__7994_ (
);

FILL FILL_0__7574_ (
);

INVX1 _9680_ (
    .A(_3028_),
    .Y(_3029_)
);

FILL FILL_0__7154_ (
);

AND2X2 _9260_ (
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2619_)
);

FILL FILL_2__8533_ (
);

FILL FILL_0__10921_ (
);

FILL FILL_0__10501_ (
);

FILL FILL_2__12779_ (
);

FILL FILL_2__12359_ (
);

FILL FILL_1__6950_ (
);

FILL FILL_1__6530_ (
);

FILL FILL_0__8779_ (
);

FILL FILL_2__13300_ (
);

FILL FILL_0__8359_ (
);

FILL FILL_3__6456_ (
);

FILL FILL_1__12713_ (
);

FILL FILL_0__9720_ (
);

FILL FILL_2__9738_ (
);

FILL FILL_0__9300_ (
);

FILL FILL_2__9318_ (
);

FILL FILL_0__11706_ (
);

FILL FILL_1__7735_ (
);

FILL FILL_1__7315_ (
);

NOR2X1 _6385_ (
    .A(_750_),
    .B(_740_),
    .Y(_760_)
);

NOR2X1 _10383_ (
    .A(_3594_),
    .B(_3591_),
    .Y(_3659_)
);

FILL FILL_0__10098_ (
);

FILL FILL_3__11852_ (
);

FILL FILL_3__11012_ (
);

FILL FILL_2__10845_ (
);

FILL FILL_2__9491_ (
);

FILL FILL_2__10425_ (
);

FILL FILL_2__9071_ (
);

FILL FILL_2__10005_ (
);

FILL FILL_3__9807_ (
);

FILL FILL_0__6845_ (
);

NOR2X1 _8951_ (
    .A(_2314_),
    .B(_2378_),
    .Y(_2373_)
);

FILL FILL_0__6425_ (
);

OAI21X1 _8531_ (
    .A(_1796_),
    .B(_1886_),
    .C(_1882_),
    .Y(_1969_)
);

DFFPOSX1 _8111_ (
    .D(\Y[1] [11]),
    .CLK(clk_bF$buf54),
    .Q(\u_fir_pe1.rYin [11])
);

DFFPOSX1 _11588_ (
    .D(_4775_[4]),
    .CLK(clk_bF$buf39),
    .Q(\Y[6] [4])
);

AOI21X1 _11168_ (
    .A(_4282_),
    .B(_4352_),
    .C(_4364_),
    .Y(_4365_)
);

FILL FILL_2__7804_ (
);

FILL FILL_3__12637_ (
);

FILL FILL_1__13251_ (
);

FILL FILL_0__12664_ (
);

FILL FILL_0__12244_ (
);

NAND2X1 _9736_ (
    .A(_3078_),
    .B(_3077_),
    .Y(_3079_)
);

AOI21X1 _9316_ (
    .A(_2674_),
    .B(_2673_),
    .C(_2672_),
    .Y(_2675_)
);

FILL FILL_1__8693_ (
);

FILL FILL_1__8273_ (
);

FILL FILL_3__8199_ (
);

FILL FILL_3__9560_ (
);

FILL FILL_0__13029_ (
);

OAI21X1 _13314_ (
    .A(_6330_),
    .B(_6331_),
    .C(_6335_),
    .Y(_6337_)
);

FILL FILL_1_CLKBUF1_insert20 (
);

FILL FILL_1_CLKBUF1_insert21 (
);

FILL FILL_1_CLKBUF1_insert22 (
);

FILL FILL_1_CLKBUF1_insert23 (
);

FILL FILL_1_CLKBUF1_insert24 (
);

FILL FILL_1__9898_ (
);

FILL FILL_1__9478_ (
);

FILL FILL_1_CLKBUF1_insert25 (
);

FILL FILL_1__9058_ (
);

FILL FILL_1_CLKBUF1_insert26 (
);

FILL FILL_1_CLKBUF1_insert27 (
);

FILL FILL_1_CLKBUF1_insert28 (
);

FILL FILL_1_CLKBUF1_insert29 (
);

FILL FILL_2__11383_ (
);

FILL FILL_1__10796_ (
);

FILL FILL_1__10376_ (
);

FILL FILL_0__7383_ (
);

FILL FILL_3__10703_ (
);

FILL FILL_2__8762_ (
);

FILL FILL_2__8342_ (
);

FILL FILL_0__10310_ (
);

FILL FILL_2__12588_ (
);

FILL FILL_2__12168_ (
);

NOR2X1 _7802_ (
    .A(_1214_),
    .B(_1259_),
    .Y(_1317_)
);

FILL FILL_0__8588_ (
);

FILL FILL_3__6685_ (
);

FILL FILL_0__8168_ (
);

NAND2X1 _10859_ (
    .A(\X[5] [1]),
    .B(vdd),
    .Y(_4060_)
);

NAND2X1 _10439_ (
    .A(vdd),
    .B(\X[4] [7]),
    .Y(_3714_)
);

INVX1 _10019_ (
    .A(_3214_),
    .Y(_3300_)
);

FILL FILL_3__11908_ (
);

FILL FILL_1__12942_ (
);

FILL FILL_1__12522_ (
);

FILL FILL_1__12102_ (
);

FILL FILL_2__9967_ (
);

FILL FILL_2__9547_ (
);

FILL FILL_0__11935_ (
);

FILL FILL_2__9127_ (
);

OAI21X1 _11800_ (
    .A(_4884_),
    .B(_4919_),
    .C(_4878_),
    .Y(_4920_)
);

FILL FILL_0__11515_ (
);

FILL FILL_1__7964_ (
);

FILL FILL_1__7544_ (
);

FILL FILL_1__7124_ (
);

FILL FILL_1__13307_ (
);

FILL FILL_3__8411_ (
);

OAI21X1 _10192_ (
    .A(_3457_),
    .B(_3461_),
    .C(_3464_),
    .Y(_3471_)
);

FILL FILL_1__8749_ (
);

FILL FILL_1__8329_ (
);

FILL FILL_3__11241_ (
);

FILL FILL_2__10654_ (
);

FILL FILL_2__10234_ (
);

NAND3X1 _7399_ (
    .A(_851_),
    .B(_908_),
    .C(_912_),
    .Y(_920_)
);

FILL FILL_0__6654_ (
);

NAND2X1 _8760_ (
    .A(_2192_),
    .B(_2166_),
    .Y(_2193_)
);

NAND3X1 _8340_ (
    .A(_1766_),
    .B(_1770_),
    .C(_1773_),
    .Y(_1780_)
);

NAND3X1 _11397_ (
    .A(_4563_),
    .B(_4565_),
    .C(_4589_),
    .Y(_4590_)
);

FILL FILL_3__12866_ (
);

FILL FILL_2__7613_ (
);

FILL FILL_3__12026_ (
);

FILL FILL_1__13060_ (
);

FILL FILL_2__11859_ (
);

FILL FILL_0__12893_ (
);

FILL FILL_2__11439_ (
);

FILL FILL_2__11019_ (
);

FILL FILL_0__12053_ (
);

FILL FILL_2__12800_ (
);

FILL FILL_0__7859_ (
);

OAI21X1 _9965_ (
    .A(_3969_),
    .B(_3206_),
    .C(_3209_),
    .Y(_3247_)
);

FILL FILL_0__7439_ (
);

NOR2X1 _9545_ (
    .A(_2896_),
    .B(_2900_),
    .Y(_2901_)
);

FILL FILL_0__7019_ (
);

NAND3X1 _9125_ (
    .A(_2476_),
    .B(_2483_),
    .C(_2485_),
    .Y(_2486_)
);

FILL FILL_0__8800_ (
);

FILL FILL_2__8818_ (
);

FILL FILL_0__13258_ (
);

NAND3X1 _13123_ (
    .A(_6141_),
    .B(_6151_),
    .C(_6154_),
    .Y(_6157_)
);

FILL FILL_1__6815_ (
);

FILL FILL_1__9287_ (
);

FILL FILL_2__11192_ (
);

FILL FILL_1__10185_ (
);

FILL FILL_0__7192_ (
);

FILL FILL_2__8571_ (
);

FILL FILL_2__8151_ (
);

FILL FILL_2__12397_ (
);

NAND2X1 _7611_ (
    .A(_1124_),
    .B(_1128_),
    .Y(_1129_)
);

FILL FILL_0__8397_ (
);

NOR2X1 _10668_ (
    .A(_3930_),
    .B(_3931_),
    .Y(_3932_)
);

NAND3X1 _10248_ (
    .A(_3518_),
    .B(_3522_),
    .C(_3520_),
    .Y(_3526_)
);

FILL FILL_1__12751_ (
);

FILL FILL_1__12331_ (
);

FILL FILL_2__9776_ (
);

FILL FILL_2__9356_ (
);

FILL FILL_0__11744_ (
);

FILL FILL_0__11324_ (
);

INVX1 _8816_ (
    .A(\u_fir_pe2.mul [3]),
    .Y(_2243_)
);

FILL FILL_1__7773_ (
);

FILL FILL_1__7353_ (
);

FILL FILL_1__13116_ (
);

FILL FILL_0__12949_ (
);

FILL FILL_3__8640_ (
);

OAI21X1 _12814_ (
    .A(_5852_),
    .B(_5848_),
    .C(_5788_),
    .Y(_5853_)
);

FILL FILL_0__12529_ (
);

FILL FILL_0__12109_ (
);

FILL FILL254550x136950 (
);

FILL FILL_1__8558_ (
);

FILL FILL_1__8138_ (
);

FILL FILL_3__11470_ (
);

FILL FILL_2__10883_ (
);

FILL FILL_2__10463_ (
);

FILL FILL_2__10043_ (
);

FILL FILL_3__9425_ (
);

FILL FILL_0__6883_ (
);

FILL FILL_0__6463_ (
);

FILL FILL_2__7842_ (
);

FILL FILL_2__7422_ (
);

FILL FILL_3__12255_ (
);

FILL FILL_2__7002_ (
);

FILL FILL_2__11668_ (
);

FILL FILL_2__11248_ (
);

FILL FILL_0__12282_ (
);

FILL FILL_0__7668_ (
);

NOR2X1 _9774_ (
    .A(\u_fir_pe3.rYin [10]),
    .B(\u_fir_pe3.mul [10]),
    .Y(_3118_)
);

NAND2X1 _9354_ (
    .A(\X[3] [4]),
    .B(vdd),
    .Y(_2712_)
);

FILL FILL_2__8627_ (
);

FILL FILL_2__8207_ (
);

FILL FILL_0__13067_ (
);

DFFPOSX1 _13352_ (
    .D(_6369_[14]),
    .CLK(clk_bF$buf9),
    .Q(\Y[7] [14])
);

FILL FILL_1__6624_ (
);

FILL FILL_1__9096_ (
);

FILL FILL_1__12807_ (
);

FILL FILL_0__9814_ (
);

FILL FILL_3__7911_ (
);

FILL FILL_1__7829_ (
);

FILL FILL_1__7409_ (
);

FILL FILL_3__10321_ (
);

FILL FILL_2__8380_ (
);

NAND3X1 _6899_ (
    .A(_460_),
    .B(_494_),
    .C(_492_),
    .Y(_495_)
);

NAND3X1 _6479_ (
    .A(Xin[1]),
    .B(gnd),
    .C(_79_),
    .Y(_80_)
);

NAND3X1 _7840_ (
    .A(_1251_),
    .B(_1353_),
    .C(_1094_),
    .Y(_1354_)
);

NAND2X1 _7420_ (
    .A(_938_),
    .B(_939_),
    .Y(_940_)
);

OAI21X1 _7000_ (
    .A(_305_),
    .B(_592_),
    .C(_571_),
    .Y(_593_)
);

FILL FILL_1__11199_ (
);

OAI21X1 _10897_ (
    .A(_4093_),
    .B(_4094_),
    .C(_4054_),
    .Y(_4098_)
);

INVX1 _10477_ (
    .A(_3750_),
    .Y(_3751_)
);

NAND2X1 _10057_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3337_)
);

FILL FILL_3__11946_ (
);

FILL FILL_1__12980_ (
);

FILL FILL_1__12560_ (
);

FILL FILL_3__11106_ (
);

FILL FILL_1__12140_ (
);

FILL FILL_2__10939_ (
);

FILL FILL_2__9585_ (
);

FILL FILL_0__11973_ (
);

FILL FILL_2__10519_ (
);

FILL FILL_2__9165_ (
);

FILL FILL_0__11553_ (
);

FILL FILL_0__11133_ (
);

FILL FILL_0__6939_ (
);

FILL FILL_0__6519_ (
);

NOR2X1 _8625_ (
    .A(_1609_),
    .B(_2056_),
    .Y(_2061_)
);

AOI22X1 _8205_ (
    .A(_1603_),
    .B(_1608_),
    .C(_1643_),
    .D(_1646_),
    .Y(_1647_)
);

FILL FILL_1__7582_ (
);

FILL FILL_1__7162_ (
);

FILL FILL_0__12758_ (
);

NAND2X1 _12623_ (
    .A(gnd),
    .B(\X[6] [4]),
    .Y(_5664_)
);

FILL FILL_0__12338_ (
);

AND2X2 _12203_ (
    .A(_5317_),
    .B(_5314_),
    .Y(_5318_)
);

FILL FILL_1__8787_ (
);

FILL FILL_1__8367_ (
);

FILL FILL_2__10692_ (
);

FILL FILL_2__10272_ (
);

FILL FILL_3__9654_ (
);

BUFX2 _13408_ (
    .A(_6377_[14]),
    .Y(Yout[14])
);

FILL FILL_0__6692_ (
);

FILL FILL_2__7651_ (
);

FILL FILL_2__11897_ (
);

FILL FILL_2__11477_ (
);

FILL FILL_2__11057_ (
);

FILL FILL_0__12091_ (
);

FILL FILL_0__7897_ (
);

FILL FILL_0__7477_ (
);

NAND2X1 _9583_ (
    .A(_2933_),
    .B(_2937_),
    .Y(_2938_)
);

FILL FILL_0__7057_ (
);

NAND2X1 _9163_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf1 ),
    .Y(_2523_)
);

FILL FILL_1__11831_ (
);

FILL FILL_1__11411_ (
);

FILL FILL_2__8856_ (
);

FILL FILL_2__8436_ (
);

FILL FILL_0__10824_ (
);

FILL FILL_0__10404_ (
);

FILL FILL_2__8016_ (
);

FILL FILL_0__13296_ (
);

NAND3X1 _13161_ (
    .A(_6161_),
    .B(_6163_),
    .C(_6191_),
    .Y(_6193_)
);

FILL FILL_1__6853_ (
);

FILL FILL_1__6433_ (
);

FILL FILL_2__13203_ (
);

FILL FILL_3__6779_ (
);

FILL FILL_1__12616_ (
);

FILL FILL253950x212550 (
);

FILL FILL_0__9623_ (
);

FILL FILL_0__9203_ (
);

FILL FILL_3__7300_ (
);

FILL FILL_3__10970_ (
);

FILL FILL_1__7638_ (
);

FILL FILL_3__10550_ (
);

FILL FILL_3__8505_ (
);

AOI21X1 _10286_ (
    .A(_3477_),
    .B(_3392_),
    .C(_3563_),
    .Y(_3564_)
);

FILL FILL_2__6922_ (
);

FILL FILL_3__11755_ (
);

FILL FILL_2__6502_ (
);

FILL FILL_3__11335_ (
);

FILL FILL_2__9394_ (
);

FILL FILL_0__11782_ (
);

FILL FILL_2__10328_ (
);

FILL FILL_0__11362_ (
);

FILL FILL_0__6748_ (
);

NOR2X1 _8854_ (
    .A(_2275_),
    .B(_2276_),
    .Y(_2277_)
);

NAND3X1 _8434_ (
    .A(_1871_),
    .B(_1872_),
    .C(_1870_),
    .Y(_1873_)
);

INVX1 _8014_ (
    .A(_1516_),
    .Y(_1518_)
);

FILL FILL_1__7391_ (
);

FILL FILL_2__7707_ (
);

FILL FILL_1__13154_ (
);

FILL FILL_0__12987_ (
);

INVX1 _12852_ (
    .A(_5883_),
    .Y(_5890_)
);

FILL FILL_0__12567_ (
);

FILL FILL_0__12147_ (
);

NOR2X1 _12432_ (
    .A(\u_fir_pe6.rYin [13]),
    .B(\u_fir_pe6.mul [13]),
    .Y(_5536_)
);

AOI21X1 _12012_ (
    .A(_5041_),
    .B(_5043_),
    .C(_5129_),
    .Y(_5130_)
);

NAND2X1 _9639_ (
    .A(_2990_),
    .B(_2991_),
    .Y(_2992_)
);

AOI22X1 _9219_ (
    .A(_2502_),
    .B(_2497_),
    .C(_2574_),
    .D(_2578_),
    .Y(_2579_)
);

FILL FILL_1__8596_ (
);

FILL FILL_1__8176_ (
);

FILL FILL_2__10081_ (
);

FILL FILL_3__9043_ (
);

AND2X2 _13217_ (
    .A(_6242_),
    .B(_6241_),
    .Y(_6369_[4])
);

FILL FILL_1__6909_ (
);

FILL FILL_2__7880_ (
);

FILL FILL_2__7460_ (
);

FILL FILL_3__12293_ (
);

FILL FILL_2__7040_ (
);

FILL FILL_2__11286_ (
);

NAND2X1 _6920_ (
    .A(_468_),
    .B(_469_),
    .Y(_515_)
);

FILL FILL_1__10699_ (
);

NAND3X1 _6500_ (
    .A(_96_),
    .B(_82_),
    .C(_100_),
    .Y(_101_)
);

FILL FILL_1__10279_ (
);

FILL FILL_0__7286_ (
);

AOI21X1 _9392_ (
    .A(_2661_),
    .B(_2663_),
    .C(_2749_),
    .Y(_2750_)
);

FILL FILL_3__10606_ (
);

FILL FILL_1__11640_ (
);

FILL FILL_1__11220_ (
);

FILL FILL_2__8665_ (
);

FILL FILL253950x61350 (
);

FILL FILL_2__8245_ (
);

FILL FILL_0__10633_ (
);

FILL FILL_3__13078_ (
);

FILL FILL_0__10213_ (
);

DFFPOSX1 _13390_ (
    .D(_6375_[12]),
    .CLK(clk_bF$buf24),
    .Q(\u_fir_pe7.mul [12])
);

NAND3X1 _7705_ (
    .A(_1140_),
    .B(_1146_),
    .C(_1221_),
    .Y(_1222_)
);

FILL FILL_1__6662_ (
);

FILL FILL_2__13012_ (
);

FILL FILL_1__12845_ (
);

FILL FILL_1__12425_ (
);

FILL FILL_1__12005_ (
);

FILL FILL_0__9432_ (
);

FILL FILL_0__11838_ (
);

FILL FILL_0__9012_ (
);

NAND3X1 _11703_ (
    .A(gnd),
    .B(\X[7] [1]),
    .C(_4824_),
    .Y(_4825_)
);

FILL FILL_0__11418_ (
);

FILL FILL_1__7867_ (
);

FILL FILL_1__7447_ (
);

FILL FILL_1__7027_ (
);

FILL FILL_3__8734_ (
);

OAI21X1 _12908_ (
    .A(_5945_),
    .B(_5942_),
    .C(_5878_),
    .Y(_5946_)
);

FILL FILL_3__8314_ (
);

NAND3X1 _10095_ (
    .A(_3372_),
    .B(_3373_),
    .C(_3374_),
    .Y(_3375_)
);

FILL FILL_2__6731_ (
);

FILL FILL_3__11564_ (
);

FILL FILL_2__10977_ (
);

FILL FILL_2__10557_ (
);

FILL FILL_2__10137_ (
);

FILL FILL_0__11171_ (
);

FILL FILL_3__9939_ (
);

FILL FILL_3__9519_ (
);

FILL FILL_0__6977_ (
);

FILL FILL_0__6557_ (
);

NOR2X1 _8663_ (
    .A(_2096_),
    .B(_2098_),
    .Y(_2099_)
);

OAI21X1 _8243_ (
    .A(_1683_),
    .B(_1609_),
    .C(_1677_),
    .Y(_1684_)
);

FILL FILL_1__10911_ (
);

FILL FILL_2__7936_ (
);

FILL FILL_2__7516_ (
);

FILL FILL_3__12349_ (
);

FILL FILL_0__12796_ (
);

NAND3X1 _12661_ (
    .A(_5633_),
    .B(_5690_),
    .C(_5694_),
    .Y(_5702_)
);

FILL FILL_0__12376_ (
);

NOR2X1 _12241_ (
    .A(_5347_),
    .B(_5351_),
    .Y(_5355_)
);

FILL FILL_2__12703_ (
);

DFFPOSX1 _9868_ (
    .D(\Y[3] [14]),
    .CLK(clk_bF$buf36),
    .Q(\u_fir_pe3.rYin [14])
);

NAND2X1 _9448_ (
    .A(_2804_),
    .B(_2800_),
    .Y(_2805_)
);

NAND2X1 _9028_ (
    .A(vdd),
    .B(\X[3] [2]),
    .Y(_2391_)
);

FILL FILL_0__8703_ (
);

FILL FILL_3__9272_ (
);

AND2X2 _13026_ (
    .A(_6055_),
    .B(_6061_),
    .Y(_6062_)
);

FILL FILL_1__6718_ (
);

FILL FILL_0__9908_ (
);

FILL FILL_2__11095_ (
);

FILL FILL_1__10088_ (
);

FILL FILL_0__7095_ (
);

FILL FILL_3__10835_ (
);

FILL FILL_3__10415_ (
);

FILL FILL_2__8894_ (
);

FILL FILL_2__8474_ (
);

FILL FILL_0__10862_ (
);

FILL FILL_0__10442_ (
);

FILL FILL_2__8054_ (
);

FILL FILL_0__10022_ (
);

NOR2X1 _7934_ (
    .A(_1439_),
    .B(_1438_),
    .Y(_1442_)
);

OAI21X1 _7514_ (
    .A(_1575_),
    .B(_1032_),
    .C(_1024_),
    .Y(_1033_)
);

FILL FILL_1__6891_ (
);

FILL FILL_1__6471_ (
);

FILL FILL_2__13241_ (
);

FILL FILL_3__6397_ (
);

FILL FILL_1__12654_ (
);

FILL FILL_1__12234_ (
);

FILL FILL_0__9661_ (
);

FILL FILL_2__9679_ (
);

FILL FILL_0__9241_ (
);

FILL FILL_2__9259_ (
);

AOI21X1 _11932_ (
    .A(_5050_),
    .B(_5045_),
    .C(_5004_),
    .Y(_5051_)
);

FILL FILL_0__11647_ (
);

OAI21X1 _11512_ (
    .A(_4694_),
    .B(_4691_),
    .C(_4693_),
    .Y(_4696_)
);

FILL FILL_0__11227_ (
);

AOI21X1 _8719_ (
    .A(_2150_),
    .B(_2051_),
    .C(_2152_),
    .Y(_2153_)
);

FILL FILL_1__7676_ (
);

FILL FILL_1__7256_ (
);

FILL FILL_1__13019_ (
);

INVX1 _12717_ (
    .A(_5675_),
    .Y(_5757_)
);

FILL FILL_2__6960_ (
);

FILL FILL_3__11793_ (
);

FILL FILL_2__6540_ (
);

FILL FILL_2__10786_ (
);

FILL FILL_2__10366_ (
);

FILL FILL_1__9822_ (
);

FILL FILL_1__9402_ (
);

FILL FILL_3__9748_ (
);

FILL FILL_0_CLKBUF1_insert30 (
);

FILL FILL_0_CLKBUF1_insert31 (
);

FILL FILL_0_CLKBUF1_insert32 (
);

FILL FILL_0_CLKBUF1_insert33 (
);

FILL FILL_0_CLKBUF1_insert34 (
);

FILL FILL_0__6786_ (
);

AOI21X1 _8892_ (
    .A(_2297_),
    .B(_2312_),
    .C(_2315_),
    .Y(_2316_)
);

FILL FILL_0_CLKBUF1_insert35 (
);

AOI21X1 _8472_ (
    .A(_1850_),
    .B(_1847_),
    .C(_1833_),
    .Y(_1910_)
);

FILL FILL_0_CLKBUF1_insert36 (
);

OAI21X1 _8052_ (
    .A(_1548_),
    .B(_1549_),
    .C(_1553_),
    .Y(_1555_)
);

FILL FILL_0_CLKBUF1_insert37 (
);

FILL FILL_0_CLKBUF1_insert38 (
);

FILL FILL_0_CLKBUF1_insert39 (
);

FILL FILL_1__10300_ (
);

FILL FILL_2__7745_ (
);

FILL FILL_3__12578_ (
);

FILL FILL_2__7325_ (
);

FILL FILL_1__13192_ (
);

NAND3X1 _12890_ (
    .A(_5921_),
    .B(_5922_),
    .C(_5923_),
    .Y(_5928_)
);

FILL FILL_0__12185_ (
);

DFFPOSX1 _12470_ (
    .D(_5572_[9]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[9])
);

OAI21X1 _12050_ (
    .A(_5097_),
    .B(_5166_),
    .C(_5136_),
    .Y(_5167_)
);

FILL FILL_2__12932_ (
);

NOR2X1 _9677_ (
    .A(\u_fir_pe3.rYin [1]),
    .B(\u_fir_pe3.mul [1]),
    .Y(_3026_)
);

NAND2X1 _9257_ (
    .A(\X[3] [2]),
    .B(vdd),
    .Y(_2616_)
);

FILL FILL_1__11925_ (
);

FILL FILL_1__11505_ (
);

FILL FILL_0__8932_ (
);

FILL FILL_0__8512_ (
);

FILL FILL_0__10918_ (
);

AOI21X1 _13255_ (
    .A(_6274_),
    .B(_6277_),
    .C(_6276_),
    .Y(_6278_)
);

FILL FILL_1__6947_ (
);

FILL FILL_1__6527_ (
);

FILL FILL_0__9717_ (
);

FILL FILL_3__10644_ (
);

FILL FILL_3__10224_ (
);

FILL FILL_2__8283_ (
);

FILL FILL_0__10671_ (
);

FILL FILL_0__10251_ (
);

INVX2 _7743_ (
    .A(gnd),
    .Y(_1259_)
);

NAND2X1 _7323_ (
    .A(_843_),
    .B(_844_),
    .Y(_845_)
);

FILL FILL_2__13050_ (
);

FILL FILL_3__11849_ (
);

FILL FILL_1__12883_ (
);

FILL FILL_3__11429_ (
);

FILL FILL_1__12043_ (
);

FILL FILL_0__9890_ (
);

FILL FILL_0__9470_ (
);

FILL FILL_2__9488_ (
);

FILL FILL_0__11876_ (
);

FILL FILL_2__9068_ (
);

FILL FILL_0__9050_ (
);

NAND3X1 _11741_ (
    .A(\X[7] [1]),
    .B(gnd),
    .C(_4861_),
    .Y(_4862_)
);

FILL FILL_0__11456_ (
);

FILL FILL_0__11036_ (
);

AOI21X1 _11321_ (
    .A(_4467_),
    .B(_4510_),
    .C(_4513_),
    .Y(_4516_)
);

NOR2X1 _8948_ (
    .A(_2370_),
    .B(_2225_),
    .Y(_2383_[0])
);

NAND3X1 _8528_ (
    .A(_1963_),
    .B(_1964_),
    .C(_1965_),
    .Y(_1966_)
);

DFFPOSX1 _8108_ (
    .D(\Y[1] [8]),
    .CLK(clk_bF$buf52),
    .Q(\u_fir_pe1.rYin [8])
);

FILL FILL_1__7485_ (
);

FILL FILL_1__7065_ (
);

FILL FILL_1__13248_ (
);

AOI22X1 _12946_ (
    .A(vdd),
    .B(\X[6] [6]),
    .C(vdd),
    .D(\X[6] [7]),
    .Y(_5983_)
);

FILL FILL_3__8352_ (
);

INVX2 _12526_ (
    .A(gnd),
    .Y(_6357_)
);

OAI21X1 _12106_ (
    .A(_5222_),
    .B(_5221_),
    .C(_5220_),
    .Y(_5223_)
);

FILL FILL_3__11182_ (
);

FILL FILL_2__10595_ (
);

FILL FILL_2__10175_ (
);

FILL FILL_1__9631_ (
);

FILL FILL_1__9211_ (
);

FILL FILL_3__9977_ (
);

FILL FILL_3__9137_ (
);

FILL FILL_0__6595_ (
);

INVX1 _8281_ (
    .A(_1714_),
    .Y(_1722_)
);

FILL FILL_2__7974_ (
);

FILL FILL_2__7554_ (
);

FILL FILL_3__12387_ (
);

FILL FILL_2__7134_ (
);

FILL FILL_2__12741_ (
);

FILL FILL_2__12321_ (
);

NAND2X1 _9486_ (
    .A(_2841_),
    .B(_2771_),
    .Y(_2843_)
);

NAND2X1 _9066_ (
    .A(_2426_),
    .B(_2427_),
    .Y(_2428_)
);

FILL FILL_1__11734_ (
);

FILL FILL_1__11314_ (
);

FILL FILL_2__8759_ (
);

FILL FILL_0__8741_ (
);

FILL FILL_0__8321_ (
);

FILL FILL_2__8339_ (
);

FILL FILL_0__10307_ (
);

FILL FILL_0__13199_ (
);

NOR2X1 _13064_ (
    .A(_5996_),
    .B(_6041_),
    .Y(_6099_)
);

FILL FILL_2__9700_ (
);

FILL FILL_1__6756_ (
);

FILL FILL_2__13106_ (
);

FILL FILL_1__12939_ (
);

FILL FILL_1__12519_ (
);

FILL FILL_0__9946_ (
);

FILL FILL_0__9526_ (
);

FILL FILL_3__7623_ (
);

FILL FILL_0__9106_ (
);

FILL FILL_0__10480_ (
);

FILL FILL_0__10060_ (
);

FILL FILL_1__8902_ (
);

FILL FILL_3__8828_ (
);

FILL FILL_3__8408_ (
);

OR2X2 _7972_ (
    .A(_1469_),
    .B(_1474_),
    .Y(_1476_)
);

OAI21X1 _7552_ (
    .A(_1070_),
    .B(_1066_),
    .C(_1006_),
    .Y(_1071_)
);

OR2X2 _7132_ (
    .A(_711_),
    .B(_715_),
    .Y(_716_)
);

AOI21X1 _10189_ (
    .A(_3467_),
    .B(_3462_),
    .C(_3323_),
    .Y(_3468_)
);

FILL FILL_2__6825_ (
);

FILL FILL_2__6405_ (
);

FILL FILL_1__12692_ (
);

FILL FILL_1__12272_ (
);

FILL FILL_2__9297_ (
);

NOR2X1 _11970_ (
    .A(_5552_),
    .B(_5087_),
    .Y(_5088_)
);

FILL FILL_0__11685_ (
);

AND2X2 _11550_ (
    .A(_4733_),
    .B(_4732_),
    .Y(_4775_[12])
);

FILL FILL_0__11265_ (
);

NAND3X1 _11130_ (
    .A(_4308_),
    .B(_4323_),
    .C(_4324_),
    .Y(_4328_)
);

NAND2X1 _8757_ (
    .A(_2161_),
    .B(_2189_),
    .Y(_2190_)
);

NAND3X1 _8337_ (
    .A(_1730_),
    .B(_1771_),
    .C(_1776_),
    .Y(_1777_)
);

FILL FILL_1__7294_ (
);

FILL FILL_1__13057_ (
);

FILL FILL_3__8581_ (
);

OAI21X1 _12755_ (
    .A(_5718_),
    .B(_5793_),
    .C(_5722_),
    .Y(_5794_)
);

NOR2X1 _12335_ (
    .A(_5440_),
    .B(_5439_),
    .Y(_5441_)
);

FILL FILL_0__13411_ (
);

FILL FILL_1__8499_ (
);

FILL FILL_1__9440_ (
);

FILL FILL_1__9020_ (
);

FILL FILL_3__9366_ (
);

DFFPOSX1 _8090_ (
    .D(_1587_[14]),
    .CLK(clk_bF$buf3),
    .Q(\Y[2] [14])
);

FILL FILL_2__7783_ (
);

FILL FILL_2__7363_ (
);

FILL FILL_3__12196_ (
);

FILL FILL_2__11189_ (
);

NAND2X1 _6823_ (
    .A(_403_),
    .B(_413_),
    .Y(_420_)
);

NAND3X1 _6403_ (
    .A(_1_),
    .B(_5_),
    .C(_3_),
    .Y(_6_)
);

FILL FILL_2__12970_ (
);

FILL FILL_2__12550_ (
);

FILL FILL_2__12130_ (
);

FILL FILL_0__7189_ (
);

OAI21X1 _9295_ (
    .A(_2649_),
    .B(_2653_),
    .C(_2615_),
    .Y(_2654_)
);

FILL FILL_3__10929_ (
);

FILL FILL_1__11963_ (
);

FILL FILL_1__11543_ (
);

FILL FILL_1__11123_ (
);

FILL FILL_0__8550_ (
);

FILL FILL_2__8568_ (
);

FILL FILL_0__10956_ (
);

FILL FILL_2__8148_ (
);

FILL FILL_0__10536_ (
);

AOI22X1 _10821_ (
    .A(vdd),
    .B(\X[5] [1]),
    .C(gnd),
    .D(\X[5] [2]),
    .Y(_4023_)
);

NAND2X1 _10401_ (
    .A(_3673_),
    .B(_3660_),
    .Y(_3677_)
);

FILL FILL_0__10116_ (
);

NOR2X1 _13293_ (
    .A(_6315_),
    .B(_6316_),
    .Y(_6369_[11])
);

AOI21X1 _7608_ (
    .A(_1125_),
    .B(_1123_),
    .C(_1121_),
    .Y(_1126_)
);

FILL FILL_1__6985_ (
);

FILL FILL_1__6565_ (
);

FILL FILL_2__13335_ (
);

FILL FILL_1__12748_ (
);

FILL FILL_1__12328_ (
);

FILL FILL_0__9755_ (
);

FILL FILL_3__7852_ (
);

FILL FILL_0__9335_ (
);

DFFPOSX1 _11606_ (
    .D(\X[5] [6]),
    .CLK(clk_bF$buf45),
    .Q(\X[6] [6])
);

FILL FILL_3__10262_ (
);

FILL FILL_1__8711_ (
);

NAND2X1 _7781_ (
    .A(_1295_),
    .B(_1296_),
    .Y(_1297_)
);

NAND2X1 _7361_ (
    .A(gnd),
    .B(\X[1] [4]),
    .Y(_882_)
);

FILL FILL_3__11887_ (
);

FILL FILL_2__6634_ (
);

FILL FILL_3__11047_ (
);

FILL FILL_1__12081_ (
);

FILL FILL_0__11494_ (
);

FILL FILL_0__11074_ (
);

FILL FILL_1__9916_ (
);

FILL FILL_2__11821_ (
);

FILL FILL_2__11401_ (
);

DFFPOSX1 _8986_ (
    .D(\Y[2] [9]),
    .CLK(clk_bF$buf44),
    .Q(\u_fir_pe2.rYin [9])
);

AOI22X1 _8566_ (
    .A(_1836_),
    .B(_2002_),
    .C(_1928_),
    .D(_1924_),
    .Y(_2003_)
);

NOR2X1 _8146_ (
    .A(_2377_),
    .B(_2376_),
    .Y(_2378_)
);

FILL FILL_1__10814_ (
);

FILL FILL_2__7839_ (
);

FILL FILL_0__7821_ (
);

FILL FILL_0__7401_ (
);

FILL FILL_2__7419_ (
);

FILL FILL_1__13286_ (
);

NAND3X1 _12984_ (
    .A(_5961_),
    .B(_6016_),
    .C(_6020_),
    .Y(_6021_)
);

FILL FILL_0__12699_ (
);

FILL FILL_0__12279_ (
);

AOI22X1 _12564_ (
    .A(\X[6] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[6] [4]),
    .Y(_5606_)
);

AND2X2 _12144_ (
    .A(\X[7]_5_bF$buf0 ),
    .B(gnd),
    .Y(_5260_)
);

FILL FILL_2__12606_ (
);

FILL FILL_0__13220_ (
);

FILL FILL_0__8606_ (
);

FILL FILL_3__6703_ (
);

FILL FILL_3__9595_ (
);

DFFPOSX1 _13349_ (
    .D(_6369_[11]),
    .CLK(clk_bF$buf9),
    .Q(\Y[7] [11])
);

FILL FILL_2__7592_ (
);

FILL FILL_2__7172_ (
);

INVX1 _6632_ (
    .A(_230_),
    .Y(_231_)
);

FILL FILL_1__11772_ (
);

FILL FILL_3__10318_ (
);

FILL FILL_1__11352_ (
);

FILL FILL_2__8797_ (
);

FILL FILL_2__8377_ (
);

FILL FILL_0__10765_ (
);

FILL FILL_0__10345_ (
);

INVX1 _10630_ (
    .A(_3891_),
    .Y(_3894_)
);

OAI21X1 _10210_ (
    .A(_3398_),
    .B(_3408_),
    .C(_3404_),
    .Y(_3488_)
);

OAI21X1 _7837_ (
    .A(_1301_),
    .B(_1304_),
    .C(_1349_),
    .Y(_1352_)
);

INVX1 _7417_ (
    .A(_936_),
    .Y(_937_)
);

FILL FILL_1__6794_ (
);

FILL FILL_2__13144_ (
);

FILL FILL_1__12977_ (
);

FILL FILL_1__12557_ (
);

FILL FILL_1__12137_ (
);

FILL FILL_0__9984_ (
);

FILL FILL_0__9564_ (
);

FILL FILL_3__7661_ (
);

FILL FILL_0__9144_ (
);

NAND2X1 _11835_ (
    .A(_4933_),
    .B(_4929_),
    .Y(_4955_)
);

OAI21X1 _11415_ (
    .A(_4601_),
    .B(_4600_),
    .C(_4606_),
    .Y(_4607_)
);

FILL FILL_0__12911_ (
);

FILL FILL_1__7999_ (
);

FILL FILL_1__7579_ (
);

FILL FILL_3__10491_ (
);

FILL FILL_1__7159_ (
);

FILL FILL_1__8940_ (
);

FILL FILL_1__8520_ (
);

FILL FILL_3__8446_ (
);

INVX1 _7590_ (
    .A(_1101_),
    .Y(_1108_)
);

NOR2X1 _7170_ (
    .A(\u_fir_pe0.rYin [13]),
    .B(\u_fir_pe0.mul [13]),
    .Y(_754_)
);

FILL FILL_2__6863_ (
);

FILL FILL_3__11696_ (
);

FILL FILL_2__6443_ (
);

FILL FILL_3__11276_ (
);

FILL FILL_2__10689_ (
);

FILL FILL_2__10269_ (
);

FILL FILL_1__9725_ (
);

FILL FILL_1__9305_ (
);

FILL FILL_2__11210_ (
);

FILL FILL_0__6689_ (
);

INVX1 _8795_ (
    .A(_1618_),
    .Y(_2385_[0])
);

NOR2X1 _8375_ (
    .A(_1807_),
    .B(_1809_),
    .Y(_1814_)
);

FILL FILL_1__10623_ (
);

FILL FILL_1__10203_ (
);

FILL FILL_0__7630_ (
);

FILL FILL_2__7648_ (
);

FILL FILL_1__13095_ (
);

NAND3X1 _12793_ (
    .A(_5825_),
    .B(_5828_),
    .C(_5826_),
    .Y(_5832_)
);

FILL FILL_0__12088_ (
);

NAND2X1 _12373_ (
    .A(_5439_),
    .B(_5451_),
    .Y(_5476_)
);

FILL FILL_2__12835_ (
);

FILL FILL_2__12415_ (
);

FILL FILL_1__11828_ (
);

FILL FILL_1__11408_ (
);

FILL FILL_0__8835_ (
);

FILL FILL_3__6932_ (
);

FILL FILL_0__8415_ (
);

AND2X2 _13158_ (
    .A(_6187_),
    .B(_6184_),
    .Y(_6191_)
);

FILL FILL_3__7717_ (
);

AOI21X1 _6861_ (
    .A(_372_),
    .B(_442_),
    .C(_456_),
    .Y(_457_)
);

NAND3X1 _6441_ (
    .A(gnd),
    .B(Xin[1]),
    .C(_42_),
    .Y(_43_)
);

FILL FILL_1__11581_ (
);

FILL FILL_1__11161_ (
);

FILL FILL_0__10994_ (
);

FILL FILL_2__8186_ (
);

FILL FILL_0__10574_ (
);

FILL FILL_0__10154_ (
);

FILL FILL_2__10901_ (
);

OAI21X1 _7646_ (
    .A(_1163_),
    .B(_1160_),
    .C(_1096_),
    .Y(_1164_)
);

DFFPOSX1 _7226_ (
    .D(Yin[3]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [3])
);

FILL FILL_0__6901_ (
);

FILL FILL_2__6919_ (
);

FILL FILL_1__12786_ (
);

FILL FILL_1__12366_ (
);

FILL FILL_0__9793_ (
);

FILL FILL_3__7890_ (
);

FILL FILL_0__9373_ (
);

FILL FILL_0__11779_ (
);

FILL FILL_3__7470_ (
);

NAND2X1 _11644_ (
    .A(vdd),
    .B(\X[7] [1]),
    .Y(_5513_)
);

FILL FILL_3__7050_ (
);

FILL FILL_0__11359_ (
);

OAI21X1 _11224_ (
    .A(_4420_),
    .B(_4419_),
    .C(_4418_),
    .Y(_4421_)
);

FILL FILL_0__12720_ (
);

FILL FILL_0__12300_ (
);

FILL FILL_1__7388_ (
);

FILL FILL_3__8675_ (
);

NOR2X1 _12849_ (
    .A(_5885_),
    .B(_5886_),
    .Y(_5887_)
);

INVX1 _12429_ (
    .A(\u_fir_pe6.rYin [13]),
    .Y(_5533_)
);

AOI21X1 _12009_ (
    .A(_5126_),
    .B(_5125_),
    .C(_5124_),
    .Y(_5127_)
);

FILL FILL_2__6672_ (
);

FILL FILL_2__10498_ (
);

FILL FILL_2__10078_ (
);

FILL FILL_1__9954_ (
);

FILL FILL_1__9534_ (
);

FILL FILL_1__9114_ (
);

FILL FILL_0__6498_ (
);

OAI22X1 _8184_ (
    .A(_1624_),
    .B(_1625_),
    .C(_1594_),
    .D(_1598_),
    .Y(_1626_)
);

FILL FILL_1__10852_ (
);

FILL FILL_1__10432_ (
);

FILL FILL_1__10012_ (
);

FILL FILL_2__7877_ (
);

FILL FILL_2__7457_ (
);

FILL FILL_2__7037_ (
);

NAND2X1 _12182_ (
    .A(_5250_),
    .B(_5251_),
    .Y(_5297_)
);

FILL FILL_3__13231_ (
);

NAND2X1 _6917_ (
    .A(_505_),
    .B(_509_),
    .Y(_512_)
);

FILL FILL_2__12644_ (
);

FILL FILL_2__12224_ (
);

AOI21X1 _9389_ (
    .A(_2746_),
    .B(_2745_),
    .C(_2744_),
    .Y(_2747_)
);

FILL FILL_1__11217_ (
);

FILL FILL_0__8644_ (
);

FILL FILL_0__8224_ (
);

AND2X2 _10915_ (
    .A(_4115_),
    .B(_4111_),
    .Y(_4781_[5])
);

DFFPOSX1 _13387_ (
    .D(_6375_[9]),
    .CLK(clk_bF$buf9),
    .Q(\u_fir_pe7.mul [9])
);

FILL FILL_2__9603_ (
);

FILL FILL_1__6659_ (
);

FILL FILL_2__13009_ (
);

FILL FILL_1__7600_ (
);

FILL FILL_3__7946_ (
);

FILL FILL_0__9429_ (
);

FILL FILL_0__9009_ (
);

AOI21X1 _6670_ (
    .A(_268_),
    .B(_263_),
    .C(_222_),
    .Y(_269_)
);

FILL FILL_3__10776_ (
);

FILL FILL_3__10356_ (
);

FILL FILL_1__11390_ (
);

FILL FILL_0__10383_ (
);

FILL FILL_1__8805_ (
);

NOR2X1 _7875_ (
    .A(_1357_),
    .B(_1380_),
    .Y(_1388_)
);

INVX1 _7455_ (
    .A(_893_),
    .Y(_975_)
);

INVX1 _7035_ (
    .A(_621_),
    .Y(_627_)
);

FILL FILL254550x54150 (
);

FILL FILL_2__13182_ (
);

FILL FILL_2__6728_ (
);

FILL FILL_0__6710_ (
);

FILL FILL_1__12595_ (
);

FILL FILL_1__12175_ (
);

FILL FILL_0__9182_ (
);

NAND2X1 _11873_ (
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4992_)
);

NAND2X1 _11453_ (
    .A(_4638_),
    .B(_4639_),
    .Y(_4775_[3])
);

FILL FILL_0__11168_ (
);

NAND2X1 _11033_ (
    .A(_4143_),
    .B(_4227_),
    .Y(_4232_)
);

FILL FILL_2__11915_ (
);

FILL FILL_1__7197_ (
);

FILL FILL_1__10908_ (
);

FILL FILL_0__7915_ (
);

INVX1 _9601_ (
    .A(_2917_),
    .Y(_2955_)
);

FILL FILL254250x61350 (
);

NAND3X1 _12658_ (
    .A(_5695_),
    .B(_5698_),
    .C(_5647_),
    .Y(_5699_)
);

FILL FILL_3__8064_ (
);

OR2X2 _12238_ (
    .A(_5351_),
    .B(_5347_),
    .Y(_5352_)
);

FILL FILL_0__13314_ (
);

FILL FILL_2__6481_ (
);

FILL FILL_1__9763_ (
);

FILL FILL_1__9343_ (
);

FILL FILL_3__9689_ (
);

FILL FILL_1__10661_ (
);

FILL FILL_1__10241_ (
);

FILL FILL_2__7686_ (
);

FILL FILL_2__7266_ (
);

NAND2X1 _6726_ (
    .A(gnd),
    .B(Xin[7]),
    .Y(_324_)
);

FILL FILL_2__12873_ (
);

FILL FILL_2__12453_ (
);

FILL FILL_2__12033_ (
);

NAND3X1 _9198_ (
    .A(_2546_),
    .B(_2557_),
    .C(_2553_),
    .Y(_2558_)
);

FILL FILL_1__11866_ (
);

FILL FILL_1__11446_ (
);

FILL FILL_1__11026_ (
);

FILL FILL_0__8873_ (
);

FILL FILL_0__8453_ (
);

FILL FILL_0__10859_ (
);

FILL FILL_3__6550_ (
);

FILL FILL_0__10439_ (
);

FILL FILL_0__8033_ (
);

DFFPOSX1 _10724_ (
    .D(\X[4] [1]),
    .CLK(clk_bF$buf25),
    .Q(\X[5] [1])
);

INVX1 _10304_ (
    .A(_3578_),
    .Y(_3581_)
);

FILL FILL_0__10019_ (
);

NOR2X1 _13196_ (
    .A(_6221_),
    .B(_6220_),
    .Y(_6224_)
);

FILL FILL_2__9412_ (
);

FILL FILL_0__11800_ (
);

FILL FILL_1__6888_ (
);

FILL FILL_1__6468_ (
);

FILL FILL_2__13238_ (
);

FILL FILL_0__9658_ (
);

NAND3X1 _11929_ (
    .A(_5042_),
    .B(_5041_),
    .C(_5043_),
    .Y(_5048_)
);

FILL FILL_0__9238_ (
);

FILL FILL_3__7335_ (
);

NAND2X1 _11509_ (
    .A(_4689_),
    .B(_4692_),
    .Y(_4775_[8])
);

FILL FILL253050x43350 (
);

FILL FILL_3__10585_ (
);

FILL FILL_3__10165_ (
);

FILL FILL_0__10192_ (
);

FILL FILL_1__8614_ (
);

AOI22X1 _7684_ (
    .A(vdd),
    .B(\X[1] [6]),
    .C(vdd),
    .D(\X[1] [7]),
    .Y(_1201_)
);

INVX2 _7264_ (
    .A(gnd),
    .Y(_1575_)
);

FILL FILL_2__6957_ (
);

FILL FILL_2__6537_ (
);

AOI21X1 _11682_ (
    .A(_4801_),
    .B(_4802_),
    .C(_5568_),
    .Y(_4805_)
);

FILL FILL_0__11397_ (
);

NAND2X1 _11262_ (
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4458_)
);

FILL FILL_1__9819_ (
);

FILL FILL_3__12731_ (
);

FILL FILL_2__11724_ (
);

FILL FILL_2__11304_ (
);

NOR2X1 _8889_ (
    .A(_2309_),
    .B(_2303_),
    .Y(_2312_)
);

NAND2X1 _8469_ (
    .A(_1900_),
    .B(_1901_),
    .Y(_1907_)
);

NAND2X1 _8049_ (
    .A(_1552_),
    .B(_1546_),
    .Y(_1553_)
);

FILL FILL_0__7724_ (
);

DFFPOSX1 _9830_ (
    .D(_3180_[0]),
    .CLK(clk_bF$buf56),
    .Q(\Y[4] [0])
);

FILL FILL_0__7304_ (
);

AND2X2 _9410_ (
    .A(_2758_),
    .B(_2763_),
    .Y(_2768_)
);

FILL FILL_1__13189_ (
);

OAI21X1 _12887_ (
    .A(_5920_),
    .B(_5924_),
    .C(_5896_),
    .Y(_5925_)
);

FILL FILL_3__8293_ (
);

DFFPOSX1 _12467_ (
    .D(_5572_[6]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[6])
);

OAI21X1 _12047_ (
    .A(_5083_),
    .B(_5163_),
    .C(_5146_),
    .Y(_5164_)
);

FILL FILL_2__12929_ (
);

FILL FILL_0__13123_ (
);

FILL FILL_0__8929_ (
);

FILL FILL_0__8509_ (
);

FILL FILL_1__9992_ (
);

FILL FILL_1__9572_ (
);

FILL FILL_1__9152_ (
);

FILL FILL_3__9078_ (
);

FILL FILL_1__10890_ (
);

FILL FILL_1__10470_ (
);

FILL FILL_1__10050_ (
);

FILL FILL_2__7495_ (
);

FILL FILL_2__7075_ (
);

OAI21X1 _6955_ (
    .A(_496_),
    .B(_549_),
    .C(_492_),
    .Y(_550_)
);

NAND2X1 _6535_ (
    .A(_131_),
    .B(_133_),
    .Y(_135_)
);

FILL FILL_2__12682_ (
);

FILL FILL_2__12262_ (
);

FILL FILL_1__11675_ (
);

FILL FILL_1__11255_ (
);

FILL FILL_0__8682_ (
);

FILL FILL_0__8262_ (
);

FILL FILL_0__10668_ (
);

INVX1 _10953_ (
    .A(_4140_),
    .Y(_4153_)
);

OAI21X1 _10533_ (
    .A(_3782_),
    .B(_3789_),
    .C(_3788_),
    .Y(_3805_)
);

FILL FILL_0__10248_ (
);

OAI21X1 _10113_ (
    .A(_3317_),
    .B(_3315_),
    .C(_3308_),
    .Y(_3393_)
);

FILL FILL_2__9641_ (
);

FILL FILL_2__9221_ (
);

FILL FILL_1__6697_ (
);

FILL FILL_2__13047_ (
);

FILL FILL_0__9887_ (
);

FILL FILL_3__7984_ (
);

FILL FILL_0__9467_ (
);

FILL FILL_3__7564_ (
);

FILL FILL_0__9047_ (
);

NAND3X1 _11738_ (
    .A(_4858_),
    .B(_4853_),
    .C(_4855_),
    .Y(_4859_)
);

FILL FILL_3__7144_ (
);

OAI21X1 _11318_ (
    .A(_4458_),
    .B(_4511_),
    .C(_4512_),
    .Y(_4513_)
);

FILL FILL_1__13401_ (
);

FILL FILL_0__12814_ (
);

FILL FILL_1__8843_ (
);

FILL FILL_1__8423_ (
);

FILL FILL_1__8003_ (
);

FILL FILL_3__8769_ (
);

FILL FILL_3__8349_ (
);

OAI21X1 _7493_ (
    .A(_936_),
    .B(_1011_),
    .C(_940_),
    .Y(_1012_)
);

NOR2X1 _7073_ (
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

FILL FILL_2__6766_ (
);

NAND2X1 _11491_ (
    .A(_4670_),
    .B(_4673_),
    .Y(_4775_[7])
);

OAI21X1 _11071_ (
    .A(_4269_),
    .B(_4265_),
    .C(_4181_),
    .Y(_4270_)
);

FILL FILL_3__12960_ (
);

FILL FILL_1__9628_ (
);

FILL FILL_1__9208_ (
);

FILL FILL_3__12120_ (
);

FILL FILL_2__11953_ (
);

FILL FILL_2__11533_ (
);

FILL FILL_2__11113_ (
);

AOI21X1 _8698_ (
    .A(_2064_),
    .B(_2080_),
    .C(_2132_),
    .Y(_2133_)
);

NAND3X1 _8278_ (
    .A(_1717_),
    .B(_1718_),
    .C(_1716_),
    .Y(_1719_)
);

FILL FILL_1__10946_ (
);

FILL FILL_1__10526_ (
);

FILL FILL_1__10106_ (
);

FILL FILL_0__7953_ (
);

FILL FILL_0__7533_ (
);

FILL FILL_0__7113_ (
);

INVX1 _12696_ (
    .A(_5735_),
    .Y(_5736_)
);

AND2X2 _12276_ (
    .A(_5385_),
    .B(_5384_),
    .Y(_5389_)
);

FILL FILL_2__8912_ (
);

FILL FILL_2__12738_ (
);

FILL FILL_2__12318_ (
);

FILL FILL_0__8738_ (
);

FILL FILL_0__8318_ (
);

FILL FILL_3__6415_ (
);

FILL FILL_1__9381_ (
);

NAND3X1 _6764_ (
    .A(_360_),
    .B(_361_),
    .C(_359_),
    .Y(_362_)
);

FILL FILL_2__12071_ (
);

FILL FILL_1__11484_ (
);

FILL FILL_1__11064_ (
);

FILL FILL_0__8491_ (
);

FILL FILL_0__10897_ (
);

FILL FILL_0__10477_ (
);

DFFPOSX1 _10762_ (
    .D(_3984_[15]),
    .CLK(clk_bF$buf38),
    .Q(\u_fir_pe4.mul [15])
);

FILL FILL_0__8071_ (
);

NAND3X1 _10342_ (
    .A(_3614_),
    .B(_3618_),
    .C(_3573_),
    .Y(_3619_)
);

FILL FILL_0__10057_ (
);

FILL FILL254250x248550 (
);

FILL FILL_2__10804_ (
);

FILL FILL_2__9450_ (
);

FILL FILL_2__9030_ (
);

NOR2X1 _7969_ (
    .A(\u_fir_pe1.rYin [6]),
    .B(\u_fir_pe1.mul [6]),
    .Y(_1473_)
);

NAND3X1 _7549_ (
    .A(_1021_),
    .B(_1063_),
    .C(_1064_),
    .Y(_1068_)
);

NOR2X1 _7129_ (
    .A(\u_fir_pe0.rYin [9]),
    .B(\u_fir_pe0.mul [9]),
    .Y(_713_)
);

FILL FILL_2__13276_ (
);

FILL FILL_0__6804_ (
);

NAND2X1 _8910_ (
    .A(_2329_),
    .B(_2322_),
    .Y(_2333_)
);

FILL FILL_1__12689_ (
);

FILL FILL_1__12269_ (
);

FILL FILL_0__9696_ (
);

FILL FILL_3__7793_ (
);

FILL FILL_0__9276_ (
);

OAI21X1 _11967_ (
    .A(_5004_),
    .B(_5084_),
    .C(_5053_),
    .Y(_5085_)
);

NOR2X1 _11547_ (
    .A(_4730_),
    .B(_4729_),
    .Y(_4731_)
);

NAND3X1 _11127_ (
    .A(_4323_),
    .B(_4324_),
    .C(_4322_),
    .Y(_4325_)
);

FILL FILL_1__13210_ (
);

FILL FILL_0__12623_ (
);

FILL FILL_0__12203_ (
);

FILL FILL_1__8652_ (
);

FILL FILL_1__8232_ (
);

FILL FILL_0__13408_ (
);

FILL FILL_2__6995_ (
);

FILL FILL_2__6575_ (
);

FILL FILL_1__9437_ (
);

FILL FILL_1__9017_ (
);

FILL FILL_2__11762_ (
);

FILL FILL_2__11342_ (
);

DFFPOSX1 _8087_ (
    .D(_1587_[11]),
    .CLK(clk_bF$buf7),
    .Q(\Y[2] [11])
);

FILL FILL_1__10335_ (
);

FILL FILL_0__7762_ (
);

FILL FILL_0__7342_ (
);

NAND2X1 _12085_ (
    .A(_5185_),
    .B(_5195_),
    .Y(_5202_)
);

FILL FILL_2__8721_ (
);

FILL FILL_2__8301_ (
);

FILL FILL_3__13134_ (
);

FILL FILL_2__12967_ (
);

FILL FILL_2__12547_ (
);

FILL FILL_2__12127_ (
);

FILL FILL_0__13161_ (
);

FILL FILL_0__8547_ (
);

FILL FILL_3__6644_ (
);

AND2X2 _10818_ (
    .A(gnd),
    .B(\X[5] [1]),
    .Y(_4020_)
);

FILL FILL_1__9190_ (
);

FILL FILL_1__12901_ (
);

FILL FILL_2__9926_ (
);

FILL FILL_2__9506_ (
);

FILL FILL_1__7923_ (
);

FILL FILL_1__7503_ (
);

FILL FILL_3__7429_ (
);

FILL FILL_3__7009_ (
);

NAND3X1 _6993_ (
    .A(_377_),
    .B(_450_),
    .C(_556_),
    .Y(_587_)
);

NAND2X1 _6573_ (
    .A(_151_),
    .B(_147_),
    .Y(_173_)
);

FILL FILL_3__10679_ (
);

FILL FILL_3__10259_ (
);

FILL FILL_1__11293_ (
);

AOI21X1 _10991_ (
    .A(_4179_),
    .B(_4187_),
    .C(_4190_),
    .Y(_4191_)
);

NOR2X1 _10571_ (
    .A(_3836_),
    .B(_3837_),
    .Y(_3838_)
);

FILL FILL_0__10286_ (
);

AND2X2 _10151_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf3 ),
    .Y(_3430_)
);

FILL FILL_1__8708_ (
);

FILL FILL_3__11200_ (
);

FILL FILL_2__10613_ (
);

NAND2X1 _7778_ (
    .A(_1290_),
    .B(_1258_),
    .Y(_1294_)
);

AND2X2 _7358_ (
    .A(_874_),
    .B(_878_),
    .Y(_879_)
);

FILL FILL_2__13085_ (
);

FILL FILL_0__6613_ (
);

FILL FILL_1__12078_ (
);

FILL FILL_0__9085_ (
);

NAND3X1 _11776_ (
    .A(_4894_),
    .B(_4895_),
    .C(_4896_),
    .Y(_4897_)
);

NOR2X1 _11356_ (
    .A(_4059_),
    .B(_4447_),
    .Y(_4550_)
);

FILL FILL_3__12825_ (
);

FILL FILL_2__11818_ (
);

FILL FILL_0__12852_ (
);

FILL FILL_0__12432_ (
);

FILL FILL_0__12012_ (
);

FILL FILL_0__7818_ (
);

NAND2X1 _9924_ (
    .A(_3969_),
    .B(_3206_),
    .Y(_3207_)
);

NAND3X1 _9504_ (
    .A(_2858_),
    .B(_2855_),
    .C(_2859_),
    .Y(_2860_)
);

FILL FILL_1__8881_ (
);

FILL FILL_1__8461_ (
);

FILL FILL_1__8041_ (
);

FILL FILL_3__8387_ (
);

FILL FILL_0__13217_ (
);

FILL FILL_2__6384_ (
);

FILL FILL_1__9666_ (
);

FILL FILL_1__9246_ (
);

FILL FILL_2__11991_ (
);

FILL FILL_2__11571_ (
);

FILL FILL_2__11151_ (
);

FILL FILL_1__10984_ (
);

FILL FILL_1__10564_ (
);

FILL FILL_1__10144_ (
);

FILL FILL_0__7991_ (
);

FILL FILL_0__7571_ (
);

FILL FILL_2__7589_ (
);

FILL FILL_2__7169_ (
);

FILL FILL_0__7151_ (
);

FILL FILL_2__8950_ (
);

FILL FILL_2__8530_ (
);

AND2X2 _6629_ (
    .A(gnd),
    .B(Xin[7]),
    .Y(_228_)
);

FILL FILL_2__12776_ (
);

FILL FILL_2__12356_ (
);

FILL FILL_1__11769_ (
);

FILL FILL_1__11349_ (
);

FILL FILL_0__8776_ (
);

FILL FILL_3__6873_ (
);

FILL FILL_0__8356_ (
);

NAND2X1 _10627_ (
    .A(_3887_),
    .B(_3890_),
    .Y(_3891_)
);

NAND2X1 _10207_ (
    .A(_3484_),
    .B(_3483_),
    .Y(_3485_)
);

FILL FILL_1__12710_ (
);

OAI21X1 _13099_ (
    .A(_6083_),
    .B(_6086_),
    .C(_6131_),
    .Y(_6134_)
);

FILL FILL_2__9735_ (
);

FILL FILL_2__9315_ (
);

FILL FILL_0__11703_ (
);

FILL FILL_1__7732_ (
);

FILL FILL_1__7312_ (
);

FILL FILL_3__7658_ (
);

NAND2X1 _6382_ (
    .A(vdd),
    .B(Xin[1]),
    .Y(_731_)
);

FILL FILL_0__12908_ (
);

NAND2X1 _10380_ (
    .A(gnd),
    .B(_3586_),
    .Y(_3656_)
);

FILL FILL_0__10095_ (
);

FILL FILL_1__8937_ (
);

FILL FILL_1__8517_ (
);

FILL FILL_2__10842_ (
);

FILL FILL_2__10422_ (
);

FILL FILL_2__10002_ (
);

NOR2X1 _7587_ (
    .A(_1103_),
    .B(_1104_),
    .Y(_1105_)
);

INVX1 _7167_ (
    .A(\u_fir_pe0.rYin [13]),
    .Y(_751_)
);

FILL FILL_0__6842_ (
);

FILL FILL_0__6422_ (
);

DFFPOSX1 _11585_ (
    .D(_4775_[1]),
    .CLK(clk_bF$buf40),
    .Q(\Y[6] [1])
);

NAND2X1 _11165_ (
    .A(_4362_),
    .B(_4361_),
    .Y(_4363_)
);

FILL FILL_2__7801_ (
);

FILL FILL_3__12634_ (
);

FILL FILL_3__12214_ (
);

FILL FILL_0__12661_ (
);

FILL FILL_2__11207_ (
);

FILL FILL_0__12241_ (
);

FILL FILL_0__7627_ (
);

OAI21X1 _9733_ (
    .A(_3074_),
    .B(_3075_),
    .C(_3071_),
    .Y(_3076_)
);

INVX1 _9313_ (
    .A(_2526_),
    .Y(_2672_)
);

FILL FILL_1__8690_ (
);

FILL FILL_1__8270_ (
);

FILL FILL_0__13026_ (
);

NAND2X1 _13311_ (
    .A(_6334_),
    .B(_6328_),
    .Y(_6335_)
);

FILL FILL_3__6509_ (
);

FILL FILL_1__9895_ (
);

FILL FILL_1__9475_ (
);

FILL FILL_1__9055_ (
);

FILL FILL_2__11380_ (
);

FILL FILL_1__10793_ (
);

FILL FILL_1__10373_ (
);

FILL FILL_2__7398_ (
);

FILL FILL_0__7380_ (
);

FILL FILL_3__10700_ (
);

FILL FILL_3__13172_ (
);

NOR2X1 _6858_ (
    .A(_373_),
    .B(_453_),
    .Y(_454_)
);

NAND3X1 _6438_ (
    .A(_34_),
    .B(_39_),
    .C(_37_),
    .Y(_40_)
);

FILL FILL_2__12585_ (
);

FILL FILL_2__12165_ (
);

FILL FILL_1__11998_ (
);

FILL FILL_1__11578_ (
);

FILL FILL_1__11158_ (
);

FILL FILL_0__8585_ (
);

FILL FILL_0__8165_ (
);

AND2X2 _10856_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf2 ),
    .Y(_4057_)
);

NAND3X1 _10436_ (
    .A(_3708_),
    .B(_3709_),
    .C(_3710_),
    .Y(_3711_)
);

AOI21X1 _10016_ (
    .A(_3288_),
    .B(_3284_),
    .C(_3270_),
    .Y(_3297_)
);

FILL FILL_2__9964_ (
);

FILL FILL_2__9544_ (
);

FILL FILL_0__11932_ (
);

FILL FILL_2__9124_ (
);

FILL FILL_0__11512_ (
);

FILL FILL_1__7961_ (
);

FILL FILL_1__7541_ (
);

FILL FILL_1__7121_ (
);

FILL FILL_3__7887_ (
);

FILL FILL_1__13304_ (
);

FILL FILL_0__12717_ (
);

FILL FILL_3__10297_ (
);

FILL FILL_1__8746_ (
);

FILL FILL_1__8326_ (
);

FILL FILL_2__10651_ (
);

FILL FILL_2__10231_ (
);

NAND3X1 _7396_ (
    .A(_913_),
    .B(_916_),
    .C(_865_),
    .Y(_917_)
);

FILL FILL_3__9613_ (
);

FILL FILL_0__6651_ (
);

FILL FILL_2__6669_ (
);

NAND2X1 _11394_ (
    .A(_4579_),
    .B(_4586_),
    .Y(_4587_)
);

FILL FILL_2__7610_ (
);

FILL FILL_3__12443_ (
);

FILL FILL_2__11856_ (
);

FILL FILL_0__12890_ (
);

FILL FILL_2__11436_ (
);

FILL FILL_2__11016_ (
);

FILL FILL_0__12050_ (
);

FILL FILL_1__10849_ (
);

FILL FILL_1__10429_ (
);

FILL FILL_1__10009_ (
);

FILL FILL_0__7856_ (
);

NAND2X1 _9962_ (
    .A(_3237_),
    .B(_3240_),
    .Y(_3244_)
);

FILL FILL_0__7436_ (
);

AOI21X1 _9542_ (
    .A(_2846_),
    .B(_2849_),
    .C(_2897_),
    .Y(_2898_)
);

FILL FILL_0__7016_ (
);

NAND3X1 _9122_ (
    .A(gnd),
    .B(\X[3] [3]),
    .C(_2474_),
    .Y(_2483_)
);

INVX1 _12599_ (
    .A(_5624_),
    .Y(_5641_)
);

NAND2X1 _12179_ (
    .A(_5287_),
    .B(_5291_),
    .Y(_5294_)
);

FILL FILL_2__8815_ (
);

FILL FILL_3__13228_ (
);

FILL FILL_0__13255_ (
);

OAI21X1 _13120_ (
    .A(_6152_),
    .B(_6153_),
    .C(_6105_),
    .Y(_6154_)
);

FILL FILL_1__6812_ (
);

FILL FILL_3__6738_ (
);

FILL FILL_1__9284_ (
);

FILL FILL_1__10182_ (
);

NAND3X1 _6667_ (
    .A(_260_),
    .B(_259_),
    .C(_261_),
    .Y(_266_)
);

FILL FILL_2__12394_ (
);

FILL FILL_1__11387_ (
);

FILL FILL_0__8394_ (
);

FILL FILL_3__6491_ (
);

OAI21X1 _10665_ (
    .A(_3927_),
    .B(_3910_),
    .C(_3926_),
    .Y(_3929_)
);

AOI21X1 _10245_ (
    .A(_3520_),
    .B(_3522_),
    .C(_3518_),
    .Y(_3523_)
);

FILL FILL_3__11714_ (
);

FILL FILL_2__9773_ (
);

FILL FILL_2__9353_ (
);

FILL FILL_0__11741_ (
);

FILL FILL_0__11321_ (
);

FILL FILL_2__13179_ (
);

FILL FILL_0__6707_ (
);

NAND2X1 _8813_ (
    .A(_2237_),
    .B(_2240_),
    .Y(_2384_[2])
);

FILL FILL_1__7770_ (
);

FILL FILL_1__7350_ (
);

FILL FILL_0__9599_ (
);

FILL FILL_0__9179_ (
);

FILL FILL_3__7276_ (
);

FILL FILL_1__13113_ (
);

FILL FILL_0__12946_ (
);

NAND3X1 _12811_ (
    .A(_5803_),
    .B(_5845_),
    .C(_5846_),
    .Y(_5850_)
);

FILL FILL_0__12526_ (
);

FILL FILL_0__12106_ (
);

FILL FILL_1__8555_ (
);

FILL FILL_1__8135_ (
);

FILL FILL_2__10880_ (
);

FILL FILL_2__10460_ (
);

FILL FILL_2__10040_ (
);

FILL FILL_0__6880_ (
);

FILL FILL_2__6898_ (
);

FILL FILL_2__6478_ (
);

FILL FILL_0__6460_ (
);

FILL FILL_3__12672_ (
);

FILL FILL_2__11665_ (
);

FILL FILL_2__11245_ (
);

FILL FILL_1__10658_ (
);

FILL FILL_1__10238_ (
);

FILL FILL_0__7665_ (
);

INVX1 _9771_ (
    .A(\u_fir_pe3.rYin [10]),
    .Y(_3115_)
);

NAND2X1 _9351_ (
    .A(\X[3] [3]),
    .B(gnd),
    .Y(_2709_)
);

FILL FILL_2__8624_ (
);

FILL FILL_2__8204_ (
);

FILL FILL_0__13064_ (
);

FILL FILL254550x190950 (
);

FILL FILL_1__6621_ (
);

FILL FILL_3__6967_ (
);

FILL FILL_1__9093_ (
);

FILL FILL_1__12804_ (
);

FILL FILL_2__9829_ (
);

FILL FILL_0__9811_ (
);

FILL FILL_2__9409_ (
);

FILL FILL_1__7826_ (
);

FILL FILL_1__7406_ (
);

NAND3X1 _6896_ (
    .A(_487_),
    .B(_491_),
    .C(_461_),
    .Y(_492_)
);

NAND3X1 _6476_ (
    .A(_76_),
    .B(_71_),
    .C(_73_),
    .Y(_77_)
);

FILL FILL_1__11196_ (
);

OAI21X1 _10894_ (
    .A(_4093_),
    .B(_4094_),
    .C(_4092_),
    .Y(_4095_)
);

AND2X2 _10474_ (
    .A(_3730_),
    .B(_3725_),
    .Y(_3748_)
);

FILL FILL_0__10189_ (
);

OAI21X1 _10054_ (
    .A(_3966_),
    .B(_3332_),
    .C(_3333_),
    .Y(_3334_)
);

FILL FILL_3__11943_ (
);

FILL FILL_3__11523_ (
);

FILL FILL_3__11103_ (
);

FILL FILL_2__10936_ (
);

FILL FILL_2__9582_ (
);

FILL FILL_0__11970_ (
);

FILL FILL_2__10516_ (
);

FILL FILL_2__9162_ (
);

FILL FILL_0__11550_ (
);

FILL FILL_0__11130_ (
);

FILL FILL_0__6936_ (
);

FILL FILL_0__6516_ (
);

OAI22X1 _8622_ (
    .A(_2011_),
    .B(_1899_),
    .C(_1619_),
    .D(_2010_),
    .Y(_2058_)
);

NAND2X1 _8202_ (
    .A(_1626_),
    .B(_1641_),
    .Y(_1644_)
);

NAND3X1 _11679_ (
    .A(_5564_),
    .B(_4796_),
    .C(_4799_),
    .Y(_4802_)
);

FILL FILL_3__7085_ (
);

AND2X2 _11259_ (
    .A(_4451_),
    .B(_4454_),
    .Y(_4455_)
);

FILL FILL_3__12728_ (
);

FILL FILL_3__12308_ (
);

FILL FILL_0__12755_ (
);

AND2X2 _12620_ (
    .A(_5656_),
    .B(_5660_),
    .Y(_5661_)
);

FILL FILL_0__12335_ (
);

AND2X2 _12200_ (
    .A(_5305_),
    .B(_5301_),
    .Y(_5315_)
);

NOR2X1 _9827_ (
    .A(_3168_),
    .B(_3111_),
    .Y(_3183_[1])
);

NAND2X1 _9407_ (
    .A(_2764_),
    .B(_2688_),
    .Y(_2765_)
);

FILL FILL_1__8784_ (
);

FILL FILL_1__8364_ (
);

FILL FILL_3__9231_ (
);

BUFX2 _13405_ (
    .A(_6377_[11]),
    .Y(Yout[11])
);

FILL FILL_1__9989_ (
);

FILL FILL_1__9569_ (
);

FILL FILL_1__9149_ (
);

FILL FILL_3__12061_ (
);

FILL FILL_2__11894_ (
);

FILL FILL_2__11474_ (
);

FILL FILL_2__11054_ (
);

FILL FILL_1__10887_ (
);

FILL FILL_1__10467_ (
);

FILL FILL_1__10047_ (
);

FILL FILL_0__7894_ (
);

FILL FILL_0__7474_ (
);

NAND2X1 _9580_ (
    .A(_2931_),
    .B(_2907_),
    .Y(_2935_)
);

FILL FILL_0__7054_ (
);

OAI21X1 _9160_ (
    .A(_2519_),
    .B(_2520_),
    .C(_2518_),
    .Y(_2521_)
);

FILL FILL_2__8853_ (
);

FILL FILL_2__8433_ (
);

FILL FILL_0__10821_ (
);

FILL FILL_3__13266_ (
);

FILL FILL_0__10401_ (
);

FILL FILL_2__8013_ (
);

FILL FILL_2__12679_ (
);

FILL FILL_2__12259_ (
);

FILL FILL_0__13293_ (
);

FILL FILL_1__6850_ (
);

FILL FILL_1__6430_ (
);

FILL FILL_0__8679_ (
);

FILL FILL_2__13200_ (
);

FILL FILL_0__8259_ (
);

FILL FILL_1__12613_ (
);

FILL FILL_0__9620_ (
);

FILL FILL_2__9638_ (
);

FILL FILL_0__9200_ (
);

FILL FILL_2__9218_ (
);

FILL FILL_1__7635_ (
);

FILL FILL_3__8922_ (
);

FILL FILL_3__8502_ (
);

NAND2X1 _10283_ (
    .A(_3560_),
    .B(_3555_),
    .Y(_3561_)
);

FILL FILL_2__9391_ (
);

FILL FILL_2__10325_ (
);

FILL FILL_3__9707_ (
);

FILL FILL_0__6745_ (
);

OAI21X1 _8851_ (
    .A(_2267_),
    .B(_2268_),
    .C(_2272_),
    .Y(_2274_)
);

AOI21X1 _8431_ (
    .A(_1778_),
    .B(_1776_),
    .C(_1869_),
    .Y(_1870_)
);

NAND2X1 _8011_ (
    .A(_1514_),
    .B(_1513_),
    .Y(_1587_[9])
);

INVX1 _11488_ (
    .A(_4665_),
    .Y(_4671_)
);

NAND3X1 _11068_ (
    .A(_4194_),
    .B(_4262_),
    .C(_4263_),
    .Y(_4267_)
);

FILL FILL_2__7704_ (
);

FILL FILL_1__13151_ (
);

FILL FILL_0__12984_ (
);

FILL FILL_0__12564_ (
);

FILL FILL_0__12144_ (
);

NAND2X1 _9636_ (
    .A(_2988_),
    .B(_2987_),
    .Y(_2989_)
);

OAI21X1 _9216_ (
    .A(_2571_),
    .B(_2572_),
    .C(_2529_),
    .Y(_2576_)
);

FILL FILL_1__8593_ (
);

FILL FILL_1__8173_ (
);

FILL FILL_2__8909_ (
);

FILL FILL_3__9460_ (
);

OAI21X1 _13214_ (
    .A(_6230_),
    .B(_6226_),
    .C(_6239_),
    .Y(_6240_)
);

FILL FILL_1__6906_ (
);

FILL FILL_1__9798_ (
);

FILL FILL_1__9378_ (
);

FILL FILL_3__12290_ (
);

FILL FILL_2__11283_ (
);

FILL FILL_1__10696_ (
);

FILL FILL_1__10276_ (
);

FILL FILL_0__7283_ (
);

FILL FILL_2__8662_ (
);

FILL FILL_2__8242_ (
);

FILL FILL_0__10630_ (
);

FILL FILL_3__13075_ (
);

FILL FILL_0__10210_ (
);

FILL FILL_2__12068_ (
);

NAND3X1 _7702_ (
    .A(_1216_),
    .B(_1217_),
    .C(_1218_),
    .Y(_1219_)
);

FILL FILL_0__8488_ (
);

FILL FILL_3__6585_ (
);

DFFPOSX1 _10759_ (
    .D(_3984_[12]),
    .CLK(clk_bF$buf43),
    .Q(\u_fir_pe4.mul [12])
);

FILL FILL_0__8068_ (
);

AOI21X1 _10339_ (
    .A(_3531_),
    .B(_3537_),
    .C(_3612_),
    .Y(_3616_)
);

FILL FILL_3__11808_ (
);

FILL FILL_1__12842_ (
);

FILL FILL_1__12422_ (
);

FILL FILL_1__12002_ (
);

FILL FILL_2__9447_ (
);

FILL FILL_0__11835_ (
);

FILL FILL_2__9027_ (
);

NAND3X1 _11700_ (
    .A(_4816_),
    .B(_4821_),
    .C(_4819_),
    .Y(_4822_)
);

FILL FILL_0__11415_ (
);

AND2X2 _8907_ (
    .A(_2326_),
    .B(_2329_),
    .Y(_2331_)
);

FILL FILL_1__7864_ (
);

FILL FILL_1__7444_ (
);

FILL FILL_1__7024_ (
);

FILL FILL_1__13207_ (
);

FILL FILL_3__8731_ (
);

NAND3X1 _12905_ (
    .A(_5882_),
    .B(_5939_),
    .C(_5940_),
    .Y(_5943_)
);

AND2X2 _10092_ (
    .A(_3322_),
    .B(_3323_),
    .Y(_3372_)
);

FILL FILL_1__8649_ (
);

FILL FILL_1__8229_ (
);

FILL FILL_3__11141_ (
);

FILL FILL_2__10974_ (
);

FILL FILL_2__10554_ (
);

FILL FILL_2__10134_ (
);

NAND2X1 _7299_ (
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_821_)
);

FILL FILL_0__6974_ (
);

FILL FILL_0__6554_ (
);

AOI21X1 _8660_ (
    .A(_2089_),
    .B(_2095_),
    .C(_2053_),
    .Y(_2096_)
);

AND2X2 _8240_ (
    .A(gnd),
    .B(\X[2] [3]),
    .Y(_1681_)
);

NAND2X1 _11297_ (
    .A(_4362_),
    .B(_4435_),
    .Y(_4493_)
);

FILL FILL_2__7933_ (
);

FILL FILL_3__12766_ (
);

FILL FILL_2__7513_ (
);

FILL FILL_2__11759_ (
);

FILL FILL_0__12793_ (
);

FILL FILL_2__11339_ (
);

FILL FILL_0__12373_ (
);

FILL FILL_2__12700_ (
);

FILL FILL_0__7759_ (
);

DFFPOSX1 _9865_ (
    .D(\Y[3] [11]),
    .CLK(clk_bF$buf0),
    .Q(\u_fir_pe3.rYin [11])
);

FILL FILL_0__7339_ (
);

NAND2X1 _9445_ (
    .A(_2792_),
    .B(_2801_),
    .Y(_2802_)
);

INVX1 _9025_ (
    .A(_3176_),
    .Y(_3177_)
);

FILL FILL_0__8700_ (
);

FILL FILL_2__8718_ (
);

FILL FILL_0__13158_ (
);

OAI21X1 _13023_ (
    .A(_5653_),
    .B(_5898_),
    .C(_6052_),
    .Y(_6059_)
);

FILL FILL_1__6715_ (
);

FILL FILL_1__9187_ (
);

FILL FILL_0__9905_ (
);

FILL FILL_2__11092_ (
);

FILL FILL_1__10085_ (
);

FILL FILL_0__7092_ (
);

FILL FILL_3__10412_ (
);

FILL FILL_2__8891_ (
);

FILL FILL_2__8471_ (
);

FILL FILL_2__8051_ (
);

FILL FILL_2__12297_ (
);

NOR2X1 _7931_ (
    .A(\u_fir_pe1.rYin [2]),
    .B(\u_fir_pe1.mul [2]),
    .Y(_1439_)
);

INVX1 _7511_ (
    .A(gnd),
    .Y(_1030_)
);

FILL FILL_0__8297_ (
);

NAND2X1 _10988_ (
    .A(_4187_),
    .B(_4179_),
    .Y(_4188_)
);

AOI21X1 _10568_ (
    .A(_3828_),
    .B(_3833_),
    .C(_3829_),
    .Y(_3835_)
);

OAI21X1 _10148_ (
    .A(_3344_),
    .B(_3348_),
    .C(_3347_),
    .Y(_3427_)
);

FILL FILL_1__12651_ (
);

FILL FILL_1__12231_ (
);

FILL FILL_2__9676_ (
);

FILL FILL_2__9256_ (
);

FILL FILL_0__11644_ (
);

FILL FILL_0__11224_ (
);

NOR3X1 _8716_ (
    .A(_2096_),
    .B(_2098_),
    .C(_2146_),
    .Y(_2150_)
);

FILL FILL_1__7673_ (
);

FILL FILL_3__7599_ (
);

FILL FILL_3__7179_ (
);

FILL FILL_1__13016_ (
);

FILL FILL_0__12849_ (
);

FILL FILL_3__8540_ (
);

NAND3X1 _12714_ (
    .A(_5741_),
    .B(_5745_),
    .C(_5747_),
    .Y(_5754_)
);

FILL FILL_0__12429_ (
);

FILL FILL_0__12009_ (
);

FILL FILL_1__8878_ (
);

FILL FILL_3__11790_ (
);

FILL FILL_1__8458_ (
);

FILL FILL_1__8038_ (
);

FILL FILL_3__11370_ (
);

FILL FILL_2__10783_ (
);

FILL FILL_2__10363_ (
);

FILL FILL_3__9325_ (
);

FILL FILL_0__6783_ (
);

FILL FILL_3__12995_ (
);

FILL FILL_2__7742_ (
);

FILL FILL_2__7322_ (
);

FILL FILL_3__12155_ (
);

FILL FILL_2__11988_ (
);

FILL FILL_2__11568_ (
);

FILL FILL_2__11148_ (
);

FILL FILL_0__12182_ (
);

FILL FILL_0__7988_ (
);

FILL FILL_0__7568_ (
);

INVX1 _9674_ (
    .A(\u_fir_pe3.rYin [1]),
    .Y(_3023_)
);

FILL FILL_0__7148_ (
);

NAND2X1 _9254_ (
    .A(_2609_),
    .B(_2612_),
    .Y(_2613_)
);

FILL FILL_1__11922_ (
);

FILL FILL_1__11502_ (
);

FILL FILL_2__8947_ (
);

FILL FILL_2__8527_ (
);

FILL FILL_0__10915_ (
);

NAND2X1 _13252_ (
    .A(_6254_),
    .B(_6266_),
    .Y(_6275_)
);

FILL FILL_1__6944_ (
);

FILL FILL_1__6524_ (
);

FILL FILL_1__12707_ (
);

FILL FILL_0__9714_ (
);

FILL FILL_3__7811_ (
);

FILL FILL_1__7729_ (
);

FILL FILL_3__10641_ (
);

FILL FILL_1__7309_ (
);

FILL FILL_2__8280_ (
);

AOI21X1 _6799_ (
    .A(_339_),
    .B(_338_),
    .C(_323_),
    .Y(_396_)
);

AND2X2 _6379_ (
    .A(Xin[1]),
    .B(gnd),
    .Y(_700_)
);

OAI21X1 _7740_ (
    .A(_1235_),
    .B(_1237_),
    .C(_1228_),
    .Y(_1256_)
);

NAND3X1 _7320_ (
    .A(_829_),
    .B(_841_),
    .C(_837_),
    .Y(_842_)
);

FILL FILL_1__11099_ (
);

INVX2 _10797_ (
    .A(\X[5] [3]),
    .Y(_4000_)
);

INVX1 _10377_ (
    .A(_3652_),
    .Y(_3653_)
);

FILL FILL_1__12880_ (
);

FILL FILL_1__12460_ (
);

FILL FILL_1__12040_ (
);

FILL FILL_2__10839_ (
);

FILL FILL_2__9485_ (
);

FILL FILL_0__11873_ (
);

FILL FILL_2__10419_ (
);

FILL FILL_2__9065_ (
);

FILL FILL_0__11453_ (
);

FILL FILL_0__11033_ (
);

FILL FILL_0__6839_ (
);

OAI21X1 _8945_ (
    .A(_2356_),
    .B(_2359_),
    .C(_2366_),
    .Y(_2369_)
);

FILL FILL_0__6419_ (
);

OAI21X1 _8525_ (
    .A(_1729_),
    .B(_1962_),
    .C(_1876_),
    .Y(_1963_)
);

DFFPOSX1 _8105_ (
    .D(\Y[1] [5]),
    .CLK(clk_bF$buf32),
    .Q(\u_fir_pe1.rYin [5])
);

FILL FILL_1__7482_ (
);

FILL FILL_1__7062_ (
);

FILL FILL_1__13245_ (
);

NAND2X1 _12943_ (
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5980_)
);

FILL FILL_0__12658_ (
);

FILL FILL_0__12238_ (
);

AOI22X1 _12523_ (
    .A(\X[6] [0]),
    .B(vdd),
    .C(\X[6] [1]),
    .D(gnd),
    .Y(_6329_)
);

INVX1 _12103_ (
    .A(_5165_),
    .Y(_5220_)
);

FILL FILL_1__8687_ (
);

FILL FILL_1__8267_ (
);

FILL FILL_2__10592_ (
);

FILL FILL_2__10172_ (
);

FILL FILL_3__9974_ (
);

FILL FILL_3__9554_ (
);

NOR2X1 _13308_ (
    .A(_6330_),
    .B(_6331_),
    .Y(_6332_)
);

FILL FILL_0__6592_ (
);

FILL FILL_2__7971_ (
);

FILL FILL_2__7551_ (
);

FILL FILL_3__12384_ (
);

FILL FILL_2__7131_ (
);

FILL FILL_2__11797_ (
);

FILL FILL_2__11377_ (
);

FILL FILL_0__7797_ (
);

FILL FILL_0__7377_ (
);

OAI21X1 _9483_ (
    .A(_2838_),
    .B(_2839_),
    .C(_2835_),
    .Y(_2840_)
);

INVX1 _9063_ (
    .A(_2424_),
    .Y(_2425_)
);

FILL FILL_1__11731_ (
);

FILL FILL_1__11311_ (
);

FILL FILL_2__8756_ (
);

FILL FILL_2__8336_ (
);

FILL FILL_3__13169_ (
);

FILL FILL_0__10304_ (
);

FILL FILL_0__13196_ (
);

NOR3X1 _13061_ (
    .A(_5884_),
    .B(_6052_),
    .C(_5995_),
    .Y(_6096_)
);

FILL FILL_1__6753_ (
);

FILL FILL_2__13103_ (
);

FILL FILL_3__6679_ (
);

FILL FILL_1__12936_ (
);

FILL FILL_0__9943_ (
);

FILL FILL_0__9523_ (
);

FILL FILL_0__11929_ (
);

FILL FILL_0__9103_ (
);

FILL FILL_0__11509_ (
);

FILL FILL254550x122550 (
);

FILL FILL_1__7958_ (
);

FILL FILL_3__10870_ (
);

FILL FILL_1__7538_ (
);

FILL FILL_1__7118_ (
);

FILL FILL_3__10030_ (
);

FILL FILL_3__8825_ (
);

NAND3X1 _10186_ (
    .A(_3459_),
    .B(_3458_),
    .C(_3460_),
    .Y(_3465_)
);

FILL FILL_2__6822_ (
);

FILL FILL_3__11655_ (
);

FILL FILL_2__6402_ (
);

FILL FILL_3__11235_ (
);

FILL FILL_2__10648_ (
);

FILL FILL_2__9294_ (
);

FILL FILL_0__11682_ (
);

FILL FILL_2__10228_ (
);

FILL FILL_0__11262_ (
);

FILL FILL_0__6648_ (
);

OAI21X1 _8754_ (
    .A(_1899_),
    .B(_2186_),
    .C(_2165_),
    .Y(_2187_)
);

AOI21X1 _8334_ (
    .A(_1768_),
    .B(_1769_),
    .C(_1767_),
    .Y(_1774_)
);

FILL FILL_1__7291_ (
);

FILL FILL_2__7607_ (
);

FILL FILL_1__13054_ (
);

FILL FILL_0__12887_ (
);

NAND2X1 _12752_ (
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5791_)
);

FILL FILL_0__12047_ (
);

INVX1 _12332_ (
    .A(\u_fir_pe6.mul [4]),
    .Y(_5438_)
);

AOI22X1 _9959_ (
    .A(_3197_),
    .B(_3202_),
    .C(_3237_),
    .D(_3240_),
    .Y(_3241_)
);

AOI21X1 _9539_ (
    .A(_2822_),
    .B(_2828_),
    .C(_2894_),
    .Y(_2895_)
);

INVX1 _9119_ (
    .A(gnd),
    .Y(_2480_)
);

FILL FILL_1__8496_ (
);

FILL FILL_3__9783_ (
);

NAND3X1 _13117_ (
    .A(_6143_),
    .B(_6150_),
    .C(_6149_),
    .Y(_6151_)
);

FILL FILL_1__6809_ (
);

FILL FILL_2__7780_ (
);

FILL FILL_2__7360_ (
);

FILL FILL_2__11186_ (
);

INVX1 _6820_ (
    .A(Xin[4]),
    .Y(_417_)
);

FILL FILL_1__10599_ (
);

OR2X2 _6400_ (
    .A(_731_),
    .B(_2_),
    .Y(_3_)
);

FILL FILL_1__10179_ (
);

FILL FILL_2_BUFX2_insert70 (
);

FILL FILL_0__7186_ (
);

NAND3X1 _9292_ (
    .A(_2630_),
    .B(_2644_),
    .C(_2647_),
    .Y(_2651_)
);

FILL FILL_2_BUFX2_insert71 (
);

FILL FILL_2_BUFX2_insert72 (
);

FILL FILL_2_BUFX2_insert73 (
);

FILL FILL_1__11960_ (
);

FILL FILL_3__10506_ (
);

FILL FILL_2_BUFX2_insert74 (
);

FILL FILL_2_BUFX2_insert75 (
);

FILL FILL_1__11540_ (
);

FILL FILL_2_BUFX2_insert76 (
);

FILL FILL_1__11120_ (
);

FILL FILL_2_BUFX2_insert77 (
);

FILL FILL_2_BUFX2_insert78 (
);

FILL FILL_2_BUFX2_insert79 (
);

FILL FILL_2__8565_ (
);

FILL FILL_0__10953_ (
);

FILL FILL_2__8145_ (
);

FILL FILL_3__13398_ (
);

FILL FILL_0__10533_ (
);

FILL FILL_0__10113_ (
);

NOR2X1 _13290_ (
    .A(_6313_),
    .B(_6312_),
    .Y(_6314_)
);

NAND3X1 _7605_ (
    .A(vdd),
    .B(\X[1] [6]),
    .C(_1122_),
    .Y(_1123_)
);

FILL FILL_1__6982_ (
);

FILL FILL_1__6562_ (
);

FILL FILL_2__13332_ (
);

FILL FILL_1__12745_ (
);

FILL FILL_1__12325_ (
);

FILL FILL_0__9752_ (
);

FILL FILL_0__9332_ (
);

FILL FILL_0__11738_ (
);

DFFPOSX1 _11603_ (
    .D(\X[5] [3]),
    .CLK(clk_bF$buf26),
    .Q(\X[6] [3])
);

FILL FILL_0__11318_ (
);

FILL FILL_1__7767_ (
);

FILL FILL_1__7347_ (
);

NAND3X1 _12808_ (
    .A(_5845_),
    .B(_5846_),
    .C(_5844_),
    .Y(_5847_)
);

FILL FILL_3__8214_ (
);

FILL FILL_3__11884_ (
);

FILL FILL_2__6631_ (
);

FILL FILL_3__11464_ (
);

FILL FILL_3__11044_ (
);

FILL FILL_2__10877_ (
);

FILL FILL_2__10457_ (
);

FILL FILL_0__11491_ (
);

FILL FILL_2__10037_ (
);

FILL FILL_0__11071_ (
);

FILL FILL_1__9913_ (
);

FILL FILL_3__9419_ (
);

FILL FILL_0__6877_ (
);

DFFPOSX1 _8983_ (
    .D(\Y[2] [6]),
    .CLK(clk_bF$buf15),
    .Q(\u_fir_pe2.rYin [6])
);

FILL FILL_0__6457_ (
);

AOI21X1 _8563_ (
    .A(_1925_),
    .B(_1999_),
    .C(_1998_),
    .Y(_2000_)
);

NAND2X1 _8143_ (
    .A(_2374_),
    .B(_2354_),
    .Y(_2375_)
);

FILL FILL_1__10811_ (
);

FILL FILL_2__7836_ (
);

FILL FILL_3__12669_ (
);

FILL FILL_2__7416_ (
);

FILL FILL_3__12249_ (
);

FILL FILL_1__13283_ (
);

INVX1 _12981_ (
    .A(_6010_),
    .Y(_6018_)
);

FILL FILL_0__12696_ (
);

FILL FILL_0__12276_ (
);

NAND2X1 _12561_ (
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5603_)
);

AND2X2 _12141_ (
    .A(_5255_),
    .B(_5198_),
    .Y(_5257_)
);

FILL FILL_2__12603_ (
);

INVX1 _9768_ (
    .A(_3110_),
    .Y(_3112_)
);

NAND2X1 _9348_ (
    .A(_2701_),
    .B(_2705_),
    .Y(_2706_)
);

FILL FILL_0__8603_ (
);

FILL FILL_3__9172_ (
);

DFFPOSX1 _13346_ (
    .D(_6369_[8]),
    .CLK(clk_bF$buf46),
    .Q(\Y[7] [8])
);

FILL FILL_1__6618_ (
);

FILL FILL_0__9808_ (
);

FILL FILL_3__7905_ (
);

FILL FILL_2__8794_ (
);

FILL FILL_2__8374_ (
);

FILL FILL_0__10342_ (
);

FILL FILL254250x198150 (
);

NAND2X1 _7834_ (
    .A(_1345_),
    .B(_1348_),
    .Y(_1349_)
);

AOI21X1 _7414_ (
    .A(_888_),
    .B(_892_),
    .C(_881_),
    .Y(_934_)
);

FILL FILL_1__6791_ (
);

FILL FILL_2__13141_ (
);

FILL FILL_1__12974_ (
);

FILL FILL_1__12554_ (
);

FILL FILL_1__12134_ (
);

FILL FILL_0__9981_ (
);

FILL FILL_2__9999_ (
);

FILL FILL_2__9579_ (
);

FILL FILL_0__9561_ (
);

FILL FILL_0__11967_ (
);

FILL FILL_0__9141_ (
);

FILL FILL_2__9159_ (
);

AOI22X1 _11832_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf1 ),
    .C(_4941_),
    .D(_4943_),
    .Y(_4952_)
);

FILL FILL_0__11547_ (
);

OR2X2 _11412_ (
    .A(_4602_),
    .B(_4603_),
    .Y(_4604_)
);

FILL FILL_0__11127_ (
);

OAI21X1 _8619_ (
    .A(_2021_),
    .B(_2023_),
    .C(_2017_),
    .Y(_2055_)
);

FILL FILL_1__7996_ (
);

FILL FILL_1__7576_ (
);

FILL FILL_1__7156_ (
);

FILL FILL_3__8863_ (
);

FILL FILL_3__8443_ (
);

NAND2X1 _12617_ (
    .A(gnd),
    .B(\X[6]_5_bF$buf3 ),
    .Y(_5658_)
);

FILL FILL_3__8023_ (
);

FILL FILL_2__6860_ (
);

FILL FILL_2__6440_ (
);

FILL FILL_2__10686_ (
);

FILL FILL_2__10266_ (
);

FILL FILL_1__9722_ (
);

FILL FILL_1__9302_ (
);

FILL FILL_3__9648_ (
);

FILL FILL_3__9228_ (
);

FILL FILL_0__6686_ (
);

OAI21X1 _8792_ (
    .A(_2210_),
    .B(_2209_),
    .C(_2221_),
    .Y(_2223_)
);

NAND3X1 _8372_ (
    .A(_1737_),
    .B(_1806_),
    .C(_1741_),
    .Y(_1811_)
);

FILL FILL_1__10620_ (
);

FILL FILL_1__10200_ (
);

FILL FILL_2__7645_ (
);

FILL FILL_1__13092_ (
);

AOI21X1 _12790_ (
    .A(_5826_),
    .B(_5828_),
    .C(_5825_),
    .Y(_5829_)
);

FILL FILL_0__12085_ (
);

INVX1 _12370_ (
    .A(\u_fir_pe6.mul [8]),
    .Y(_5473_)
);

FILL FILL_2__12832_ (
);

FILL FILL_2__12412_ (
);

OAI21X1 _9997_ (
    .A(_3277_),
    .B(_3203_),
    .C(_3271_),
    .Y(_3278_)
);

NAND2X1 _9577_ (
    .A(_2931_),
    .B(_2930_),
    .Y(_2932_)
);

INVX1 _9157_ (
    .A(_2458_),
    .Y(_2518_)
);

FILL FILL_1__11825_ (
);

FILL FILL_1__11405_ (
);

FILL FILL_0__8832_ (
);

FILL FILL_0__8412_ (
);

FILL FILL_0__10818_ (
);

FILL FILL253950x14550 (
);

NAND2X1 _13155_ (
    .A(_6184_),
    .B(_6187_),
    .Y(_6188_)
);

FILL FILL_1__6847_ (
);

FILL FILL_1__6427_ (
);

FILL FILL_0__9617_ (
);

FILL FILL_3__10964_ (
);

FILL FILL_3__10124_ (
);

FILL FILL_0__10991_ (
);

FILL FILL_2__8183_ (
);

FILL FILL_0__10571_ (
);

FILL FILL_0__10151_ (
);

FILL FILL_3__8919_ (
);

NAND3X1 _7643_ (
    .A(_1100_),
    .B(_1157_),
    .C(_1158_),
    .Y(_1161_)
);

DFFPOSX1 _7223_ (
    .D(Yin[0]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [0])
);

FILL FILL_2__6916_ (
);

FILL FILL_3__11749_ (
);

FILL FILL_1__12783_ (
);

FILL FILL_1__12363_ (
);

FILL FILL_0__9790_ (
);

FILL FILL_2__9388_ (
);

FILL FILL_0__9370_ (
);

FILL FILL_0__11776_ (
);

AND2X2 _11641_ (
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_5482_)
);

FILL FILL_0__11356_ (
);

AOI21X1 _11221_ (
    .A(_4338_),
    .B(_4340_),
    .C(_4417_),
    .Y(_4418_)
);

NAND2X1 _8848_ (
    .A(_2271_),
    .B(_2266_),
    .Y(_2272_)
);

AOI21X1 _8428_ (
    .A(_1866_),
    .B(_1865_),
    .C(_1864_),
    .Y(_1867_)
);

INVX1 _8008_ (
    .A(_1511_),
    .Y(_1512_)
);

FILL FILL_1__7385_ (
);

FILL FILL_1__13148_ (
);

INVX2 _12846_ (
    .A(gnd),
    .Y(_5884_)
);

OR2X2 _12426_ (
    .A(_5523_),
    .B(_5528_),
    .Y(_5530_)
);

INVX1 _12006_ (
    .A(_5104_),
    .Y(_5124_)
);

FILL FILL_3__11082_ (
);

FILL FILL_2__10495_ (
);

FILL FILL253050x248550 (
);

FILL FILL_2__10075_ (
);

FILL FILL_1__9951_ (
);

FILL FILL_1__9531_ (
);

FILL FILL_1__9111_ (
);

FILL FILL_3__9037_ (
);

FILL FILL_0__6495_ (
);

INVX1 _8181_ (
    .A(_1622_),
    .Y(_1623_)
);

FILL FILL_2__7874_ (
);

FILL FILL_2__7454_ (
);

FILL FILL_2__7034_ (
);

NOR2X1 _6914_ (
    .A(_505_),
    .B(_509_),
    .Y(_510_)
);

FILL FILL_2__12641_ (
);

FILL FILL_2__12221_ (
);

AND2X2 _9386_ (
    .A(_2705_),
    .B(_2701_),
    .Y(_2744_)
);

FILL FILL_1__11214_ (
);

FILL FILL_2__8659_ (
);

FILL FILL_0__8641_ (
);

FILL FILL_2__8239_ (
);

FILL FILL_0__8221_ (
);

FILL FILL_0__10627_ (
);

INVX1 _10912_ (
    .A(_4105_),
    .Y(_4113_)
);

FILL FILL_0__10207_ (
);

FILL FILL_0__13099_ (
);

DFFPOSX1 _13384_ (
    .D(_6375_[6]),
    .CLK(clk_bF$buf11),
    .Q(\u_fir_pe7.mul [6])
);

FILL FILL_2__9600_ (
);

FILL FILL_1__6656_ (
);

FILL FILL_2__13006_ (
);

FILL FILL_1__12839_ (
);

FILL FILL_1__12419_ (
);

FILL FILL_0__9426_ (
);

FILL FILL_3__7523_ (
);

FILL FILL_3__10353_ (
);

FILL FILL_0__10380_ (
);

FILL FILL_1__8802_ (
);

FILL FILL_3__8308_ (
);

INVX1 _7872_ (
    .A(_1382_),
    .Y(_1386_)
);

NAND3X1 _7452_ (
    .A(_959_),
    .B(_963_),
    .C(_965_),
    .Y(_972_)
);

NOR3X1 _7032_ (
    .A(_623_),
    .B(_591_),
    .C(_609_),
    .Y(_624_)
);

AOI21X1 _10089_ (
    .A(_3359_),
    .B(_3355_),
    .C(_3340_),
    .Y(_3369_)
);

FILL FILL_3__11978_ (
);

FILL FILL_2__6725_ (
);

FILL FILL_3__11558_ (
);

FILL FILL_1__12592_ (
);

FILL FILL_3__11138_ (
);

FILL FILL_1__12172_ (
);

FILL FILL_2__9197_ (
);

INVX1 _11870_ (
    .A(_4984_),
    .Y(_4989_)
);

NOR2X1 _11450_ (
    .A(_4636_),
    .B(_4635_),
    .Y(_4637_)
);

FILL FILL_0__11165_ (
);

OAI21X1 _11030_ (
    .A(_4074_),
    .B(_4059_),
    .C(_4143_),
    .Y(_4229_)
);

FILL FILL_2__11912_ (
);

AND2X2 _8657_ (
    .A(_2081_),
    .B(_2085_),
    .Y(_2093_)
);

OAI22X1 _8237_ (
    .A(_2325_),
    .B(_1677_),
    .C(_1627_),
    .D(_1632_),
    .Y(_1678_)
);

FILL FILL_1__7194_ (
);

FILL FILL_1__10905_ (
);

FILL FILL_0__7912_ (
);

FILL FILL_3__8481_ (
);

NAND3X1 _12655_ (
    .A(_5691_),
    .B(_5685_),
    .C(_5689_),
    .Y(_5696_)
);

NOR2X1 _12235_ (
    .A(_4926_),
    .B(_5087_),
    .Y(_5349_)
);

FILL FILL_0__13311_ (
);

FILL FILL_1__8399_ (
);

FILL FILL_1__9760_ (
);

FILL FILL_1__9340_ (
);

FILL FILL_3__9266_ (
);

FILL FILL_2__7683_ (
);

FILL FILL_2__7263_ (
);

FILL FILL_3__12096_ (
);

FILL FILL_2__11089_ (
);

NAND2X1 _6723_ (
    .A(Xin[4]),
    .B(gnd),
    .Y(_321_)
);

FILL FILL_2__12870_ (
);

FILL FILL_2__12450_ (
);

FILL FILL_2__12030_ (
);

FILL FILL_0__7089_ (
);

NAND2X1 _9195_ (
    .A(gnd),
    .B(\X[3] [4]),
    .Y(_2555_)
);

FILL FILL_3__10829_ (
);

FILL FILL_1__11863_ (
);

FILL FILL_1__11443_ (
);

FILL FILL_1__11023_ (
);

FILL FILL_0__8870_ (
);

FILL FILL_2__8888_ (
);

FILL FILL_2__8468_ (
);

FILL FILL_0__8450_ (
);

FILL FILL_0__10856_ (
);

FILL FILL_0__10436_ (
);

DFFPOSX1 _10721_ (
    .D(_3978_[14]),
    .CLK(clk_bF$buf18),
    .Q(\Y[5] [14])
);

FILL FILL_2__8048_ (
);

FILL FILL_0__8030_ (
);

AOI21X1 _10301_ (
    .A(\X[4] [3]),
    .B(gnd),
    .C(_3575_),
    .Y(_3578_)
);

FILL FILL_0__10016_ (
);

NOR2X1 _13193_ (
    .A(\u_fir_pe7.rYin [2]),
    .B(\u_fir_pe7.mul [2]),
    .Y(_6221_)
);

NOR2X1 _7928_ (
    .A(_1436_),
    .B(_1435_),
    .Y(_1587_[1])
);

AOI22X1 _7508_ (
    .A(gnd),
    .B(\X[1] [7]),
    .C(\X[1] [3]),
    .D(gnd),
    .Y(_1027_)
);

FILL FILL_1__6885_ (
);

FILL FILL_1__6465_ (
);

FILL FILL_2__13235_ (
);

FILL FILL_1__12648_ (
);

FILL FILL_1__12228_ (
);

FILL FILL_0__9655_ (
);

FILL FILL_3__7752_ (
);

FILL FILL_0__9235_ (
);

OAI21X1 _11926_ (
    .A(_5040_),
    .B(_5044_),
    .C(_5006_),
    .Y(_5045_)
);

NOR2X1 _11506_ (
    .A(_4678_),
    .B(_4677_),
    .Y(_4690_)
);

FILL FILL_3__10582_ (
);

FILL FILL_1__8611_ (
);

FILL FILL_3__8537_ (
);

NAND2X1 _7681_ (
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1198_)
);

AOI22X1 _7261_ (
    .A(\X[1] [0]),
    .B(vdd),
    .C(\X[1] [1]),
    .D(gnd),
    .Y(_1547_)
);

FILL FILL253950x133350 (
);

FILL FILL_2__6954_ (
);

FILL FILL_2__6534_ (
);

FILL FILL_0__11394_ (
);

FILL FILL_1__9816_ (
);

FILL FILL_2__11721_ (
);

FILL FILL_2__11301_ (
);

OR2X2 _8886_ (
    .A(_2305_),
    .B(_2309_),
    .Y(_2310_)
);

OAI21X1 _8466_ (
    .A(_1902_),
    .B(_1903_),
    .C(_1898_),
    .Y(_1904_)
);

NOR2X1 _8046_ (
    .A(_1548_),
    .B(_1549_),
    .Y(_1550_)
);

FILL FILL_2__7739_ (
);

FILL FILL_0__7721_ (
);

FILL FILL_0__7301_ (
);

FILL FILL_2__7319_ (
);

FILL FILL_1__13186_ (
);

NAND3X1 _12884_ (
    .A(_5902_),
    .B(_5917_),
    .C(_5918_),
    .Y(_5922_)
);

FILL FILL_0__12599_ (
);

FILL FILL_3__8290_ (
);

FILL FILL_0__12179_ (
);

DFFPOSX1 _12464_ (
    .D(_5572_[3]),
    .CLK(clk_bF$buf29),
    .Q(_6377_[3])
);

INVX1 _12044_ (
    .A(_5154_),
    .Y(_5161_)
);

FILL FILL_2__12926_ (
);

FILL FILL_0__13120_ (
);

FILL FILL_1__11919_ (
);

FILL FILL_0__8926_ (
);

FILL FILL_0__8506_ (
);

FILL FILL_3__9495_ (
);

NOR2X1 _13249_ (
    .A(\u_fir_pe7.rYin [8]),
    .B(\u_fir_pe7.mul [8]),
    .Y(_6272_)
);

FILL FILL_2__7492_ (
);

FILL FILL_2__7072_ (
);

NAND2X1 _6952_ (
    .A(_542_),
    .B(_546_),
    .Y(_547_)
);

NAND2X1 _6532_ (
    .A(gnd),
    .B(Xin_5_bF$buf3),
    .Y(_132_)
);

FILL FILL_1__11672_ (
);

FILL FILL_3__10218_ (
);

FILL FILL_1__11252_ (
);

FILL FILL_2__8697_ (
);

FILL FILL_2__8277_ (
);

FILL FILL_0__10665_ (
);

NAND3X1 _10950_ (
    .A(vdd),
    .B(\X[5] [3]),
    .C(_4149_),
    .Y(_4150_)
);

FILL FILL_0__10245_ (
);

NAND3X1 _10530_ (
    .A(_3770_),
    .B(_3772_),
    .C(_3800_),
    .Y(_3802_)
);

NAND3X1 _10110_ (
    .A(_3383_),
    .B(_3384_),
    .C(_3389_),
    .Y(_3390_)
);

AOI21X1 _7737_ (
    .A(_1238_),
    .B(_1234_),
    .C(_1179_),
    .Y(_1253_)
);

NAND2X1 _7317_ (
    .A(vdd),
    .B(\X[1] [2]),
    .Y(_839_)
);

FILL FILL_1__6694_ (
);

FILL FILL_2__13044_ (
);

FILL FILL_1__12877_ (
);

FILL FILL_1__12457_ (
);

FILL FILL_1__12037_ (
);

FILL FILL_3__7981_ (
);

FILL FILL_0__9464_ (
);

FILL FILL_0__9044_ (
);

INVX2 _11735_ (
    .A(\X[7]_5_bF$buf2 ),
    .Y(_4856_)
);

NAND2X1 _11315_ (
    .A(_4316_),
    .B(_4390_),
    .Y(_4510_)
);

FILL FILL_0__12811_ (
);

FILL FILL_1__7899_ (
);

FILL FILL_1__7479_ (
);

FILL FILL_3__10391_ (
);

FILL FILL_1__7059_ (
);

FILL FILL_1__8840_ (
);

FILL FILL_1__8420_ (
);

FILL FILL_1__8000_ (
);

FILL FILL_3__8766_ (
);

NAND2X1 _7490_ (
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_1009_)
);

INVX1 _7070_ (
    .A(\u_fir_pe0.mul [4]),
    .Y(_656_)
);

FILL FILL_2__6763_ (
);

FILL FILL_3__11176_ (
);

FILL FILL_2__10589_ (
);

FILL FILL_2__10169_ (
);

FILL FILL_1__9625_ (
);

FILL FILL_1__9205_ (
);

FILL FILL_2__11950_ (
);

FILL FILL_2__11530_ (
);

FILL FILL_2__11110_ (
);

FILL FILL_0__6589_ (
);

AND2X2 _8695_ (
    .A(_2129_),
    .B(_2126_),
    .Y(_2130_)
);

NAND3X1 _8275_ (
    .A(_1715_),
    .B(_1648_),
    .C(_1651_),
    .Y(_1716_)
);

FILL FILL_1__10943_ (
);

FILL FILL_1__10523_ (
);

FILL FILL_1__10103_ (
);

FILL FILL_0__7950_ (
);

FILL FILL_2__7968_ (
);

FILL FILL_0__7530_ (
);

FILL FILL_2__7548_ (
);

FILL FILL_0__7110_ (
);

FILL FILL_2__7128_ (
);

AOI22X1 _12693_ (
    .A(vdd),
    .B(\X[6] [2]),
    .C(vdd),
    .D(\X[6] [3]),
    .Y(_5733_)
);

NAND2X1 _12273_ (
    .A(_5384_),
    .B(_5385_),
    .Y(_5386_)
);

FILL FILL_3__13322_ (
);

FILL FILL_2__12735_ (
);

FILL FILL_2__12315_ (
);

FILL FILL_1__11728_ (
);

FILL FILL_1__11308_ (
);

FILL FILL_0__8735_ (
);

FILL FILL_3__6832_ (
);

FILL FILL_0__8315_ (
);

FILL FILL_3__6412_ (
);

AOI21X1 _13058_ (
    .A(_6039_),
    .B(_6073_),
    .C(_6092_),
    .Y(_6093_)
);

FILL FILL_3__7617_ (
);

AOI21X1 _6761_ (
    .A(_270_),
    .B(_272_),
    .C(_358_),
    .Y(_359_)
);

FILL FILL_3__10447_ (
);

FILL FILL_1__11481_ (
);

FILL FILL_1__11061_ (
);

FILL FILL_0__10894_ (
);

FILL FILL_0__10474_ (
);

FILL FILL_0__10054_ (
);

FILL FILL_2__10801_ (
);

INVX1 _7966_ (
    .A(\u_fir_pe1.rYin [6]),
    .Y(_1470_)
);

NAND3X1 _7546_ (
    .A(_1063_),
    .B(_1064_),
    .C(_1062_),
    .Y(_1065_)
);

INVX1 _7126_ (
    .A(_705_),
    .Y(_709_)
);

FILL FILL_2__13273_ (
);

FILL FILL_2__6819_ (
);

FILL FILL_0__6801_ (
);

FILL FILL_1__12686_ (
);

FILL FILL_1__12266_ (
);

FILL FILL_0__9693_ (
);

FILL FILL_0__9273_ (
);

OAI21X1 _11964_ (
    .A(_4992_),
    .B(_5002_),
    .C(_4998_),
    .Y(_5082_)
);

FILL FILL_0__11679_ (
);

FILL FILL_3__7370_ (
);

INVX1 _11544_ (
    .A(\u_fir_pe5.mul [12]),
    .Y(_4728_)
);

FILL FILL_0__11259_ (
);

AOI21X1 _11124_ (
    .A(_4231_),
    .B(_4234_),
    .C(_4240_),
    .Y(_4322_)
);

FILL FILL_0__12620_ (
);

FILL FILL_0__12200_ (
);

FILL FILL_1__7288_ (
);

OAI21X1 _12749_ (
    .A(_5715_),
    .B(_5787_),
    .C(_5756_),
    .Y(_5788_)
);

FILL FILL_3__8155_ (
);

OR2X2 _12329_ (
    .A(_5429_),
    .B(_5434_),
    .Y(_5436_)
);

FILL FILL_0__13405_ (
);

FILL FILL_2__6992_ (
);

FILL FILL_2__6572_ (
);

FILL FILL_2__10398_ (
);

FILL FILL_1__9434_ (
);

FILL FILL_1__9014_ (
);

FILL FILL_0__6398_ (
);

DFFPOSX1 _8084_ (
    .D(_1587_[8]),
    .CLK(clk_bF$buf57),
    .Q(\Y[2] [8])
);

FILL FILL_1__10332_ (
);

FILL FILL_2__7777_ (
);

FILL FILL_2__7357_ (
);

INVX1 _12082_ (
    .A(\X[7] [4]),
    .Y(_5199_)
);

NAND2X1 _6817_ (
    .A(_413_),
    .B(_409_),
    .Y(_414_)
);

FILL FILL_2__12964_ (
);

FILL FILL_2__12544_ (
);

FILL FILL_2__12124_ (
);

NAND3X1 _9289_ (
    .A(_2644_),
    .B(_2643_),
    .C(_2647_),
    .Y(_2648_)
);

FILL FILL_1__11957_ (
);

FILL FILL_1__11537_ (
);

FILL FILL_1__11117_ (
);

FILL FILL_0__8544_ (
);

OAI22X1 _10815_ (
    .A(_4015_),
    .B(_4016_),
    .C(_3985_),
    .D(_3989_),
    .Y(_4017_)
);

OAI21X1 _13287_ (
    .A(_6303_),
    .B(_6304_),
    .C(_6308_),
    .Y(_6311_)
);

FILL FILL_2__9923_ (
);

FILL FILL_2__9503_ (
);

FILL FILL_1__6979_ (
);

FILL FILL_1__6559_ (
);

FILL FILL_2__13329_ (
);

FILL FILL_1__7920_ (
);

FILL FILL_1__7500_ (
);

FILL FILL_0__9749_ (
);

FILL FILL_3__7846_ (
);

FILL FILL_0__9329_ (
);

FILL FILL_3__7006_ (
);

OR2X2 _6990_ (
    .A(_583_),
    .B(_560_),
    .Y(_584_)
);

AOI22X1 _6570_ (
    .A(gnd),
    .B(Xin_5_bF$buf2),
    .C(_159_),
    .D(_161_),
    .Y(_170_)
);

FILL FILL_3__10676_ (
);

FILL FILL_1__11290_ (
);

FILL FILL_0__10283_ (
);

FILL FILL_1__8705_ (
);

FILL FILL_2__10610_ (
);

NAND3X1 _7775_ (
    .A(_1220_),
    .B(_1223_),
    .C(_1290_),
    .Y(_1291_)
);

NAND2X1 _7355_ (
    .A(gnd),
    .B(\X[1]_5_bF$buf1 ),
    .Y(_876_)
);

FILL FILL_2__13082_ (
);

FILL FILL_2__6628_ (
);

FILL FILL_0__6610_ (
);

FILL FILL_1__12075_ (
);

FILL FILL_0__9082_ (
);

INVX1 _11773_ (
    .A(_4808_),
    .Y(_4894_)
);

FILL FILL_0__11488_ (
);

FILL FILL_0__11068_ (
);

OAI21X1 _11353_ (
    .A(_4515_),
    .B(_4509_),
    .C(_4519_),
    .Y(_4547_)
);

FILL FILL_3__12822_ (
);

FILL FILL_3__12402_ (
);

FILL FILL_2__11815_ (
);

FILL FILL_1__7097_ (
);

FILL FILL_1__10808_ (
);

FILL FILL_0__7815_ (
);

NAND2X1 _9921_ (
    .A(_3201_),
    .B(_3197_),
    .Y(_3204_)
);

OAI22X1 _9501_ (
    .A(_2406_),
    .B(_2853_),
    .C(_2854_),
    .D(_2856_),
    .Y(_2857_)
);

OAI21X1 _12978_ (
    .A(_6014_),
    .B(_6013_),
    .C(_6012_),
    .Y(_6015_)
);

FILL FILL_3__8384_ (
);

INVX1 _12558_ (
    .A(_5600_),
    .Y(_5601_)
);

OAI21X1 _12138_ (
    .A(_5201_),
    .B(_5253_),
    .C(_5189_),
    .Y(_5254_)
);

FILL FILL_0__13214_ (
);

FILL FILL_2__6381_ (
);

FILL FILL_1__9663_ (
);

FILL FILL_1__9243_ (
);

FILL FILL_3__9589_ (
);

FILL FILL_1__10981_ (
);

FILL FILL_1__10561_ (
);

FILL FILL_1__10141_ (
);

FILL FILL_2__7586_ (
);

FILL FILL_2__7166_ (
);

NAND2X1 _6626_ (
    .A(Xin[2]),
    .B(gnd),
    .Y(_225_)
);

FILL FILL_2__12773_ (
);

FILL FILL_2__12353_ (
);

NOR3X1 _9098_ (
    .A(_2444_),
    .B(_2411_),
    .C(_2456_),
    .Y(_2459_)
);

FILL FILL_1__11766_ (
);

FILL FILL_1__11346_ (
);

FILL FILL_0__8773_ (
);

FILL FILL_0__8353_ (
);

FILL FILL_3__6450_ (
);

FILL FILL_0__10339_ (
);

AOI21X1 _10624_ (
    .A(_3883_),
    .B(_3886_),
    .C(_3885_),
    .Y(_3887_)
);

AND2X2 _10204_ (
    .A(_3482_),
    .B(_3478_),
    .Y(_3984_[7])
);

NAND2X1 _13096_ (
    .A(_6127_),
    .B(_6130_),
    .Y(_6131_)
);

FILL FILL_2__9732_ (
);

FILL FILL_2__9312_ (
);

FILL FILL_0__11700_ (
);

FILL FILL_1__6788_ (
);

FILL FILL_2__13138_ (
);

FILL FILL_0__9978_ (
);

FILL FILL_0__9558_ (
);

FILL FILL_0__9138_ (
);

NAND3X1 _11829_ (
    .A(_4937_),
    .B(_4948_),
    .C(_4944_),
    .Y(_4949_)
);

OAI21X1 _11409_ (
    .A(_4569_),
    .B(_4594_),
    .C(_4593_),
    .Y(_4601_)
);

FILL FILL_0__12905_ (
);

FILL FILL_3__10065_ (
);

FILL FILL_0__10092_ (
);

FILL FILL_1__8934_ (
);

FILL FILL_1__8514_ (
);

INVX2 _7584_ (
    .A(gnd),
    .Y(_1102_)
);

OR2X2 _7164_ (
    .A(_741_),
    .B(_746_),
    .Y(_748_)
);

FILL FILL_3__9801_ (
);

FILL FILL_2__6857_ (
);

FILL FILL_2__6437_ (
);

NOR2X1 _11582_ (
    .A(_4705_),
    .B(_4769_),
    .Y(_4764_)
);

FILL FILL_0__11297_ (
);

OAI21X1 _11162_ (
    .A(_4187_),
    .B(_4277_),
    .C(_4273_),
    .Y(_4360_)
);

FILL FILL_1__9719_ (
);

FILL FILL_2__11204_ (
);

INVX1 _8789_ (
    .A(_2215_),
    .Y(_2221_)
);

AND2X2 _8369_ (
    .A(_1739_),
    .B(_1743_),
    .Y(_1808_)
);

FILL FILL_1__10617_ (
);

FILL FILL_0__7624_ (
);

INVX1 _9730_ (
    .A(\u_fir_pe3.mul [7]),
    .Y(_3073_)
);

NAND3X1 _9310_ (
    .A(_2613_),
    .B(_2654_),
    .C(_2659_),
    .Y(_2669_)
);

FILL FILL_1__13089_ (
);

NAND2X1 _12787_ (
    .A(_5737_),
    .B(_5821_),
    .Y(_5826_)
);

NAND2X1 _12367_ (
    .A(_5469_),
    .B(_5468_),
    .Y(_5470_)
);

FILL FILL_2__12829_ (
);

FILL FILL_2__12409_ (
);

FILL FILL_0__13023_ (
);

FILL FILL_0__8829_ (
);

FILL FILL_3__6926_ (
);

FILL FILL_0__8409_ (
);

FILL FILL_3__6506_ (
);

FILL FILL_1__9892_ (
);

FILL FILL_1__9472_ (
);

FILL FILL_1__9052_ (
);

FILL FILL_1__10790_ (
);

FILL FILL_1__10370_ (
);

FILL FILL_2__7395_ (
);

NAND2X1 _6855_ (
    .A(_450_),
    .B(_380_),
    .Y(_452_)
);

NAND2X1 _6435_ (
    .A(_35_),
    .B(_36_),
    .Y(_37_)
);

FILL FILL_2__12582_ (
);

FILL FILL_2__12162_ (
);

FILL FILL_1__11995_ (
);

FILL FILL_1__11575_ (
);

FILL FILL_1__11155_ (
);

FILL FILL_0__8582_ (
);

FILL FILL_0__10988_ (
);

FILL FILL_0__8162_ (
);

FILL FILL_0__10568_ (
);

OAI21X1 _10853_ (
    .A(_4014_),
    .B(_4048_),
    .C(_4030_),
    .Y(_4054_)
);

NOR2X1 _10433_ (
    .A(_3605_),
    .B(_3650_),
    .Y(_3708_)
);

FILL FILL_0__10148_ (
);

NAND3X1 _10013_ (
    .A(_3289_),
    .B(_3293_),
    .C(_3257_),
    .Y(_3294_)
);

FILL FILL_3__11902_ (
);

FILL FILL_2__9961_ (
);

FILL FILL_2__9541_ (
);

FILL FILL_2__9121_ (
);

FILL FILL_1__6597_ (
);

FILL FILL_0__9787_ (
);

FILL FILL_0__9367_ (
);

FILL FILL_3__7464_ (
);

DFFPOSX1 _11638_ (
    .D(_4781_[14]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [14])
);

OAI21X1 _11218_ (
    .A(_4414_),
    .B(_4413_),
    .C(_4412_),
    .Y(_4415_)
);

FILL FILL_1__13301_ (
);

FILL FILL_0__12714_ (
);

FILL FILL_3__10294_ (
);

FILL FILL_1__8743_ (
);

FILL FILL_1__8323_ (
);

FILL FILL254250x14550 (
);

FILL FILL_3__8249_ (
);

NAND3X1 _7393_ (
    .A(_909_),
    .B(_903_),
    .C(_907_),
    .Y(_914_)
);

FILL FILL_3__9610_ (
);

FILL FILL_2__6666_ (
);

FILL FILL254550x248550 (
);

FILL FILL_3__11499_ (
);

FILL FILL_3__11079_ (
);

NAND2X1 _11391_ (
    .A(_4583_),
    .B(_4557_),
    .Y(_4584_)
);

FILL FILL_1__9948_ (
);

FILL FILL_1__9528_ (
);

FILL FILL_1__9108_ (
);

FILL FILL_3__12020_ (
);

FILL FILL_2__11853_ (
);

FILL FILL_2__11433_ (
);

FILL FILL_2__11013_ (
);

OAI21X1 _8598_ (
    .A(_2034_),
    .B(_2033_),
    .C(_2032_),
    .Y(_2035_)
);

NOR2X1 _8178_ (
    .A(_1618_),
    .B(_1619_),
    .Y(_1620_)
);

FILL FILL_1__10846_ (
);

FILL FILL_1__10426_ (
);

FILL FILL_1__10006_ (
);

FILL FILL_0__7853_ (
);

FILL FILL_0__7433_ (
);

FILL FILL_0__7013_ (
);

OAI21X1 _12596_ (
    .A(_6360_),
    .B(_5597_),
    .C(_5600_),
    .Y(_5638_)
);

NOR2X1 _12176_ (
    .A(_5287_),
    .B(_5291_),
    .Y(_5292_)
);

FILL FILL_2__8812_ (
);

FILL FILL_2__12638_ (
);

FILL FILL_2__12218_ (
);

FILL FILL_0__13252_ (
);

FILL FILL_0__8638_ (
);

FILL FILL_3__6735_ (
);

FILL FILL_0__8218_ (
);

NAND3X1 _10909_ (
    .A(_4108_),
    .B(_4109_),
    .C(_4107_),
    .Y(_4110_)
);

FILL FILL_1__9281_ (
);

OAI21X1 _6664_ (
    .A(_258_),
    .B(_262_),
    .C(_224_),
    .Y(_263_)
);

FILL FILL_2__12391_ (
);

FILL FILL_1__11384_ (
);

FILL FILL_0__8391_ (
);

FILL FILL_0__10797_ (
);

FILL FILL_0__10377_ (
);

NOR2X1 _10662_ (
    .A(_3924_),
    .B(_3925_),
    .Y(_3978_[11])
);

NAND2X1 _10242_ (
    .A(_3515_),
    .B(_3519_),
    .Y(_3520_)
);

FILL FILL_2__9770_ (
);

FILL FILL_2__10704_ (
);

FILL FILL_2__9350_ (
);

AOI21X1 _7869_ (
    .A(_1354_),
    .B(_1356_),
    .C(_1382_),
    .Y(_1383_)
);

NAND3X1 _7449_ (
    .A(_964_),
    .B(_949_),
    .C(_968_),
    .Y(_969_)
);

NAND2X1 _7029_ (
    .A(_620_),
    .B(_619_),
    .Y(_621_)
);

FILL FILL_2__13176_ (
);

FILL FILL_0__6704_ (
);

INVX1 _8810_ (
    .A(_2234_),
    .Y(_2238_)
);

FILL FILL_1__12589_ (
);

FILL FILL_1__12169_ (
);

FILL FILL_0__9596_ (
);

FILL FILL_3__7693_ (
);

FILL FILL_0__9176_ (
);

OAI21X1 _11867_ (
    .A(_4911_),
    .B(_4909_),
    .C(_4902_),
    .Y(_4987_)
);

INVX1 _11447_ (
    .A(\u_fir_pe5.mul [3]),
    .Y(_4634_)
);

NAND2X1 _11027_ (
    .A(vdd),
    .B(\X[5] [4]),
    .Y(_4226_)
);

FILL FILL_3__12916_ (
);

FILL FILL_1__13110_ (
);

FILL FILL_2__11909_ (
);

FILL FILL_0__12943_ (
);

FILL FILL_0__12523_ (
);

FILL FILL_0__12103_ (
);

FILL FILL_0__7909_ (
);

FILL FILL_1__8552_ (
);

FILL FILL_1__8132_ (
);

FILL FILL_3__8898_ (
);

FILL FILL_3__8478_ (
);

FILL FILL_3__8058_ (
);

FILL FILL_0__13308_ (
);

FILL FILL_2__6895_ (
);

FILL FILL_2__6475_ (
);

FILL FILL_1__9757_ (
);

FILL FILL_1__9337_ (
);

FILL FILL_2__11662_ (
);

FILL FILL_2__11242_ (
);

FILL FILL_1__10655_ (
);

FILL FILL_1__10235_ (
);

FILL FILL_0__7662_ (
);

FILL FILL_2__8621_ (
);

FILL FILL_2__8201_ (
);

FILL FILL_3__13034_ (
);

FILL FILL_2__12867_ (
);

FILL FILL_2__12447_ (
);

FILL FILL_2__12027_ (
);

FILL FILL_0__13061_ (
);

FILL FILL_0__8867_ (
);

FILL FILL_0__8447_ (
);

FILL FILL_3__6544_ (
);

DFFPOSX1 _10718_ (
    .D(_3978_[11]),
    .CLK(clk_bF$buf50),
    .Q(\Y[5] [11])
);

FILL FILL_0__8027_ (
);

FILL FILL_1__9090_ (
);

FILL FILL_1__12801_ (
);

FILL FILL_2__9826_ (
);

FILL FILL_2__9406_ (
);

FILL FILL_1__7823_ (
);

FILL FILL_1__7403_ (
);

FILL FILL_3__7329_ (
);

NAND2X1 _6893_ (
    .A(_485_),
    .B(_472_),
    .Y(_489_)
);

INVX2 _6473_ (
    .A(Xin_5_bF$buf3),
    .Y(_74_)
);

FILL FILL_3__10999_ (
);

FILL FILL_3__10159_ (
);

FILL FILL_1__11193_ (
);

AOI21X1 _10891_ (
    .A(_4013_),
    .B(_4033_),
    .C(_4047_),
    .Y(_4092_)
);

NAND3X1 _10471_ (
    .A(_3642_),
    .B(_3744_),
    .C(_3485_),
    .Y(_3745_)
);

FILL FILL_0__10186_ (
);

NAND2X1 _10051_ (
    .A(_3329_),
    .B(_3330_),
    .Y(_3331_)
);

FILL FILL_1__8608_ (
);

FILL FILL_3__11520_ (
);

FILL FILL_2__10933_ (
);

FILL FILL_2__10513_ (
);

NOR2X1 _7678_ (
    .A(_929_),
    .B(_1118_),
    .Y(_1195_)
);

NOR2X1 _7258_ (
    .A(_1486_),
    .B(_1507_),
    .Y(_1517_)
);

FILL FILL_0__6933_ (
);

FILL FILL_0__6513_ (
);

FILL FILL_1__12398_ (
);

OAI21X1 _11676_ (
    .A(_5560_),
    .B(_4797_),
    .C(_4798_),
    .Y(_4799_)
);

NOR2X1 _11256_ (
    .A(_4000_),
    .B(_4447_),
    .Y(_4452_)
);

FILL FILL_2__11718_ (
);

FILL FILL_0__12752_ (
);

FILL FILL_0__12332_ (
);

FILL FILL_0__7718_ (
);

NOR2X1 _9824_ (
    .A(\u_fir_pe3.rYin [0]),
    .B(\u_fir_pe3.mul [0]),
    .Y(_3167_)
);

NAND3X1 _9404_ (
    .A(_2692_),
    .B(_2753_),
    .C(_2748_),
    .Y(_2762_)
);

FILL FILL_1__8781_ (
);

FILL FILL_1__8361_ (
);

FILL FILL_0__13117_ (
);

BUFX2 _13402_ (
    .A(_6377_[0]),
    .Y(Yout[0])
);

FILL FILL_1__9986_ (
);

FILL FILL_1__9566_ (
);

FILL FILL_1__9146_ (
);

FILL FILL_2__11891_ (
);

FILL FILL_2__11471_ (
);

FILL FILL_2__11051_ (
);

FILL FILL_1__10884_ (
);

FILL FILL_1__10464_ (
);

FILL FILL_1__10044_ (
);

FILL FILL_0__7891_ (
);

FILL FILL_0__7471_ (
);

FILL FILL_2__7489_ (
);

FILL FILL_0__7051_ (
);

FILL FILL_2__7069_ (
);

FILL FILL254250x234150 (
);

FILL FILL_2__8850_ (
);

FILL FILL_2__8430_ (
);

FILL FILL_3__13263_ (
);

FILL FILL_2__8010_ (
);

NAND2X1 _6949_ (
    .A(_540_),
    .B(_516_),
    .Y(_544_)
);

OAI21X1 _6529_ (
    .A(_128_),
    .B(_129_),
    .C(_127_),
    .Y(_130_)
);

FILL FILL_2__12676_ (
);

FILL FILL_2__12256_ (
);

FILL FILL_0__13290_ (
);

FILL FILL_1__11669_ (
);

FILL FILL_1__11249_ (
);

FILL FILL_0__8676_ (
);

FILL FILL_3__6773_ (
);

FILL FILL_0__8256_ (
);

NAND3X1 _10947_ (
    .A(_4142_),
    .B(_4146_),
    .C(_4144_),
    .Y(_4147_)
);

AND2X2 _10527_ (
    .A(_3796_),
    .B(_3793_),
    .Y(_3800_)
);

AOI21X1 _10107_ (
    .A(_3374_),
    .B(_3373_),
    .C(_3324_),
    .Y(_3387_)
);

FILL FILL_1__12610_ (
);

FILL FILL_2__9635_ (
);

FILL FILL_2__9215_ (
);

FILL FILL_1__7632_ (
);

FILL FILL_3__7558_ (
);

FILL FILL254550x90150 (
);

FILL FILL_0__12808_ (
);

FILL FILL_3__10388_ (
);

NAND3X1 _10280_ (
    .A(_3488_),
    .B(_3552_),
    .C(_3553_),
    .Y(_3558_)
);

FILL FILL_1__8837_ (
);

FILL FILL_1__8417_ (
);

FILL FILL_2__10322_ (
);

OAI21X1 _7487_ (
    .A(_933_),
    .B(_1005_),
    .C(_974_),
    .Y(_1006_)
);

OR2X2 _7067_ (
    .A(_647_),
    .B(_652_),
    .Y(_654_)
);

FILL FILL_3__9704_ (
);

FILL FILL_0__6742_ (
);

NOR2X1 _11485_ (
    .A(_4666_),
    .B(_4667_),
    .Y(_4668_)
);

NAND3X1 _11065_ (
    .A(_4262_),
    .B(_4263_),
    .C(_4261_),
    .Y(_4264_)
);

FILL FILL_2__7701_ (
);

FILL FILL_3__12534_ (
);

FILL FILL_3__12114_ (
);

FILL FILL_2__11947_ (
);

FILL FILL_0__12981_ (
);

FILL FILL_2__11527_ (
);

FILL FILL_0__12561_ (
);

FILL FILL_2__11107_ (
);

FILL FILL_0__12141_ (
);

FILL FILL_0__7947_ (
);

FILL FILL_0__7527_ (
);

NOR2X1 _9633_ (
    .A(_2626_),
    .B(_2853_),
    .Y(_2986_)
);

FILL FILL_0__7107_ (
);

OAI21X1 _9213_ (
    .A(_2571_),
    .B(_2572_),
    .C(_2570_),
    .Y(_2573_)
);

FILL FILL_1__8590_ (
);

FILL FILL_1__8170_ (
);

FILL FILL_2__8906_ (
);

NOR2X1 _13211_ (
    .A(\u_fir_pe7.rYin [4]),
    .B(\u_fir_pe7.mul [4]),
    .Y(_6237_)
);

FILL FILL_1__6903_ (
);

FILL FILL_3__6829_ (
);

FILL FILL_1__9795_ (
);

FILL FILL_1__9375_ (
);

FILL FILL_2__11280_ (
);

FILL FILL_1__10693_ (
);

FILL FILL_1__10273_ (
);

FILL FILL_2__7298_ (
);

FILL FILL_0__7280_ (
);

FILL FILL_3__10600_ (
);

AOI21X1 _6758_ (
    .A(_355_),
    .B(_354_),
    .C(_353_),
    .Y(_356_)
);

FILL FILL_2__12065_ (
);

FILL FILL_1__11898_ (
);

FILL FILL_1__11478_ (
);

FILL FILL_1__11058_ (
);

FILL FILL_0__8485_ (
);

DFFPOSX1 _10756_ (
    .D(_3984_[9]),
    .CLK(clk_bF$buf21),
    .Q(\u_fir_pe4.mul [9])
);

FILL FILL_0__8065_ (
);

NAND3X1 _10336_ (
    .A(_3531_),
    .B(_3537_),
    .C(_3612_),
    .Y(_3613_)
);

FILL FILL_2__9444_ (
);

FILL FILL_0__11832_ (
);

FILL FILL_2__9024_ (
);

FILL FILL_0__11412_ (
);

NOR2X1 _8904_ (
    .A(\u_fir_pe2.rYin [11]),
    .B(\u_fir_pe2.mul [11]),
    .Y(_2328_)
);

FILL FILL_1__7861_ (
);

FILL FILL_1__7441_ (
);

FILL FILL_1__7021_ (
);

FILL FILL_3__7787_ (
);

FILL FILL_1__13204_ (
);

NAND3X1 _12902_ (
    .A(_5894_),
    .B(_5925_),
    .C(_5930_),
    .Y(_5940_)
);

FILL FILL_0__12617_ (
);

FILL FILL_1__8646_ (
);

FILL FILL_1__8226_ (
);

FILL FILL_2__10971_ (
);

FILL FILL_2__10551_ (
);

FILL FILL_2__10131_ (
);

INVX1 _7296_ (
    .A(_818_),
    .Y(_819_)
);

FILL FILL_3__9933_ (
);

FILL FILL_2__6989_ (
);

FILL FILL_0__6971_ (
);

FILL FILL_2__6569_ (
);

FILL FILL_0__6551_ (
);

NOR2X1 _11294_ (
    .A(_4487_),
    .B(_4489_),
    .Y(_4490_)
);

FILL FILL_2__7930_ (
);

FILL FILL_3__12763_ (
);

FILL FILL_2__7510_ (
);

FILL FILL_3__12343_ (
);

FILL FILL_2__11756_ (
);

FILL FILL_0__12790_ (
);

FILL FILL_2__11336_ (
);

FILL FILL_0__12370_ (
);

FILL FILL_1__10329_ (
);

FILL FILL_0__7756_ (
);

DFFPOSX1 _9862_ (
    .D(\Y[3] [8]),
    .CLK(clk_bF$buf36),
    .Q(\u_fir_pe3.rYin [8])
);

FILL FILL_0__7336_ (
);

AND2X2 _9442_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2799_)
);

NOR2X1 _9022_ (
    .A(_3171_),
    .B(_3151_),
    .Y(_3174_)
);

DFFPOSX1 _12499_ (
    .D(\Y[7] [14]),
    .CLK(clk_bF$buf9),
    .Q(\u_fir_pe6.rYin [14])
);

NAND2X1 _12079_ (
    .A(_5195_),
    .B(_5191_),
    .Y(_5196_)
);

FILL FILL_2__8715_ (
);

FILL FILL_3__13128_ (
);

FILL FILL_0__13155_ (
);

AND2X2 _13020_ (
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_6056_)
);

FILL FILL_1__6712_ (
);

FILL FILL_1__9184_ (
);

FILL FILL_0__9902_ (
);

FILL FILL_1__10082_ (
);

FILL FILL_1__7917_ (
);

INVX1 _6987_ (
    .A(_580_),
    .Y(_581_)
);

NAND3X1 _6567_ (
    .A(_155_),
    .B(_166_),
    .C(_162_),
    .Y(_167_)
);

FILL FILL_2__12294_ (
);

FILL FILL_1__11287_ (
);

FILL FILL_0__8294_ (
);

AOI21X1 _10985_ (
    .A(_4167_),
    .B(_4162_),
    .C(_4169_),
    .Y(_4185_)
);

FILL FILL_3__6391_ (
);

NOR2X1 _10565_ (
    .A(_3830_),
    .B(_3829_),
    .Y(_3833_)
);

OAI21X1 _10145_ (
    .A(_3966_),
    .B(_3423_),
    .C(_3415_),
    .Y(_3424_)
);

FILL FILL_2__9673_ (
);

FILL FILL_2__10607_ (
);

FILL FILL_2__9253_ (
);

FILL FILL_0__11641_ (
);

FILL FILL_0__11221_ (
);

FILL FILL_2__13079_ (
);

FILL FILL_0__6607_ (
);

NAND3X1 _8713_ (
    .A(_2105_),
    .B(_2147_),
    .C(_2106_),
    .Y(_2148_)
);

FILL FILL_1__7670_ (
);

FILL FILL_0__9499_ (
);

FILL FILL_0__9079_ (
);

FILL FILL_3__7176_ (
);

FILL FILL_1__13013_ (
);

FILL FILL_0__12846_ (
);

NAND3X1 _12711_ (
    .A(_5746_),
    .B(_5731_),
    .C(_5750_),
    .Y(_5751_)
);

FILL FILL_0__12426_ (
);

FILL FILL_0__12006_ (
);

NAND3X1 _9918_ (
    .A(_3198_),
    .B(_3200_),
    .C(_3199_),
    .Y(_3201_)
);

FILL FILL_1__8875_ (
);

FILL FILL_1__8455_ (
);

FILL FILL_1__8035_ (
);

FILL FILL_2__10780_ (
);

FILL FILL_2__10360_ (
);

FILL FILL_3__9742_ (
);

FILL FILL_3__9322_ (
);

FILL FILL_0__6780_ (
);

FILL FILL_2__6798_ (
);

FILL FILL_2__6378_ (
);

FILL FILL_3__12992_ (
);

FILL FILL_2__11985_ (
);

FILL FILL_2__11565_ (
);

FILL FILL_2__11145_ (
);

FILL FILL_1__10978_ (
);

FILL FILL_1__10558_ (
);

FILL FILL_1__10138_ (
);

FILL FILL_0__7985_ (
);

FILL FILL_0__7565_ (
);

NAND2X1 _9671_ (
    .A(_3021_),
    .B(_3020_),
    .Y(_3187_[15])
);

FILL FILL_0__7145_ (
);

AOI21X1 _9251_ (
    .A(_2538_),
    .B(_2534_),
    .C(_2603_),
    .Y(_2610_)
);

FILL FILL_2__8944_ (
);

FILL FILL_2__8524_ (
);

FILL FILL_0__10912_ (
);

FILL FILL_1__6941_ (
);

FILL FILL_1__6521_ (
);

FILL FILL_3__6867_ (
);

FILL FILL_3__6447_ (
);

FILL FILL_1__12704_ (
);

FILL FILL_2__9729_ (
);

FILL FILL_0__9711_ (
);

FILL FILL_2__9309_ (
);

FILL FILL_1__7726_ (
);

FILL FILL_1__7306_ (
);

INVX1 _6796_ (
    .A(_390_),
    .Y(_393_)
);

FILL FILL_1__11096_ (
);

OAI21X1 _10794_ (
    .A(_3989_),
    .B(_3992_),
    .C(_3986_),
    .Y(_3997_)
);

INVX2 _10374_ (
    .A(gnd),
    .Y(_3650_)
);

FILL FILL_0__10089_ (
);

FILL FILL_3__11843_ (
);

FILL FILL_3__11003_ (
);

FILL FILL_2__10836_ (
);

FILL FILL_2__9482_ (
);

FILL FILL_0__11870_ (
);

FILL FILL_2__10416_ (
);

FILL FILL_2__9062_ (
);

FILL FILL_0__11450_ (
);

FILL FILL_0__11030_ (
);

FILL FILL_0__6836_ (
);

NAND2X1 _8942_ (
    .A(_2363_),
    .B(_2365_),
    .Y(_2366_)
);

FILL FILL_0__6416_ (
);

AOI21X1 _8522_ (
    .A(_1959_),
    .B(_1958_),
    .C(_1894_),
    .Y(_1960_)
);

DFFPOSX1 _8102_ (
    .D(\Y[1] [2]),
    .CLK(clk_bF$buf52),
    .Q(\u_fir_pe1.rYin [2])
);

AOI21X1 _11999_ (
    .A(_5114_),
    .B(_5116_),
    .C(_5112_),
    .Y(_5117_)
);

NOR2X1 _11579_ (
    .A(_4761_),
    .B(_4616_),
    .Y(_4774_[0])
);

NAND3X1 _11159_ (
    .A(_4354_),
    .B(_4355_),
    .C(_4356_),
    .Y(_4357_)
);

FILL FILL_3__12628_ (
);

FILL FILL_3__12208_ (
);

FILL FILL_1__13242_ (
);

NOR2X1 _12940_ (
    .A(_5711_),
    .B(_5900_),
    .Y(_5977_)
);

FILL FILL_0__12655_ (
);

FILL FILL_0__12235_ (
);

NOR2X1 _12520_ (
    .A(_6268_),
    .B(_6289_),
    .Y(_6299_)
);

AOI21X1 _12100_ (
    .A(_5207_),
    .B(_5205_),
    .C(_5177_),
    .Y(_5217_)
);

AND2X2 _9727_ (
    .A(_3070_),
    .B(_3069_),
    .Y(_3181_[6])
);

INVX1 _9307_ (
    .A(_2568_),
    .Y(_2666_)
);

FILL FILL_1__8684_ (
);

FILL FILL_1__8264_ (
);

OAI21X1 _13305_ (
    .A(_6321_),
    .B(_6322_),
    .C(_6326_),
    .Y(_6328_)
);

FILL FILL_1__9889_ (
);

FILL FILL_1__9469_ (
);

FILL FILL_1__9049_ (
);

FILL FILL_2__11794_ (
);

FILL FILL_2__11374_ (
);

FILL FILL_1__10787_ (
);

FILL FILL_1__10367_ (
);

FILL FILL_0__7794_ (
);

FILL FILL_0__7374_ (
);

NAND3X1 _9480_ (
    .A(_2817_),
    .B(_2821_),
    .C(_2824_),
    .Y(_2837_)
);

NAND2X1 _9060_ (
    .A(gnd),
    .B(\X[3] [1]),
    .Y(_2422_)
);

FILL FILL_2__8753_ (
);

FILL FILL_2__8333_ (
);

FILL FILL_0__10301_ (
);

FILL FILL_2__12999_ (
);

FILL FILL_2__12579_ (
);

FILL FILL_2__12159_ (
);

FILL FILL_0__13193_ (
);

FILL FILL_1__6750_ (
);

FILL FILL_2__13100_ (
);

FILL FILL_0__8579_ (
);

FILL FILL_0__8159_ (
);

FILL FILL_1__12933_ (
);

FILL FILL_2__9958_ (
);

FILL FILL_0__9940_ (
);

FILL FILL_2__9538_ (
);

FILL FILL_0__9520_ (
);

FILL FILL_0__11926_ (
);

FILL FILL_2__9118_ (
);

FILL FILL_0__9100_ (
);

FILL FILL_0__11506_ (
);

FILL FILL_1__7955_ (
);

FILL FILL_1__7535_ (
);

FILL FILL_1__7115_ (
);

FILL FILL_3__8402_ (
);

OAI21X1 _10183_ (
    .A(_3461_),
    .B(_3457_),
    .C(_3397_),
    .Y(_3462_)
);

FILL FILL_3__11232_ (
);

FILL FILL_2__10645_ (
);

FILL FILL_2__9291_ (
);

FILL FILL_2__10225_ (
);

FILL FILL_0__6645_ (
);

NOR2X1 _8751_ (
    .A(_2180_),
    .B(_2184_),
    .Y(_2390_[12])
);

NAND3X1 _8331_ (
    .A(_1766_),
    .B(_1732_),
    .C(_1770_),
    .Y(_1771_)
);

NAND2X1 _11388_ (
    .A(_4552_),
    .B(_4580_),
    .Y(_4581_)
);

FILL FILL_3__12857_ (
);

FILL FILL_2__7604_ (
);

FILL FILL_3__12437_ (
);

FILL FILL_3__12017_ (
);

FILL FILL_1__13051_ (
);

FILL FILL_0__12884_ (
);

FILL FILL_0__12044_ (
);

NAND2X1 _9956_ (
    .A(_3220_),
    .B(_3235_),
    .Y(_3238_)
);

NAND3X1 _9536_ (
    .A(_2887_),
    .B(_2888_),
    .C(_2891_),
    .Y(_2892_)
);

INVX1 _9116_ (
    .A(_2476_),
    .Y(_2477_)
);

FILL FILL_1__8493_ (
);

FILL FILL_1__8073_ (
);

FILL FILL_2__8809_ (
);

FILL FILL_3__9360_ (
);

FILL FILL_0__13249_ (
);

AOI21X1 _13114_ (
    .A(gnd),
    .B(_6145_),
    .C(_6147_),
    .Y(_6148_)
);

FILL FILL_1__6806_ (
);

FILL FILL_1__9698_ (
);

FILL FILL_1__9278_ (
);

FILL FILL_3__12190_ (
);

FILL FILL_2__11183_ (
);

FILL FILL_1__10596_ (
);

FILL FILL_1__10176_ (
);

FILL FILL_0__7183_ (
);

FILL FILL_2__8562_ (
);

FILL FILL_0__10950_ (
);

FILL FILL_2__8142_ (
);

FILL FILL_0__10530_ (
);

FILL FILL_0__10110_ (
);

FILL FILL_2__12388_ (
);

OAI21X1 _7602_ (
    .A(_1037_),
    .B(_1045_),
    .C(_1044_),
    .Y(_1120_)
);

FILL FILL_0__8388_ (
);

FILL FILL_3__6485_ (
);

NOR2X1 _10659_ (
    .A(_3922_),
    .B(_3921_),
    .Y(_3923_)
);

AOI21X1 _10239_ (
    .A(_3516_),
    .B(_3514_),
    .C(_3512_),
    .Y(_3517_)
);

FILL FILL_3__11708_ (
);

FILL FILL_1__12742_ (
);

FILL FILL_1__12322_ (
);

FILL FILL_2__9767_ (
);

FILL FILL_2__9347_ (
);

FILL FILL_0__11735_ (
);

DFFPOSX1 _11600_ (
    .D(\X[5] [0]),
    .CLK(clk_bF$buf27),
    .Q(\X[6] [0])
);

FILL FILL_0__11315_ (
);

AND2X2 _8807_ (
    .A(\u_fir_pe2.rYin [2]),
    .B(\u_fir_pe2.mul [2]),
    .Y(_2235_)
);

FILL FILL_1__7764_ (
);

FILL FILL_1__7344_ (
);

FILL FILL_1__13107_ (
);

FILL FILL_3__8631_ (
);

AOI21X1 _12805_ (
    .A(_5731_),
    .B(_5750_),
    .C(_5843_),
    .Y(_5844_)
);

FILL FILL_1__8549_ (
);

FILL FILL_3__11461_ (
);

FILL FILL_2__10874_ (
);

FILL FILL_2__10454_ (
);

FILL FILL_2__10034_ (
);

FILL FILL_1__9910_ (
);

DFFPOSX1 _7199_ (
    .D(_789_[0]),
    .CLK(clk_bF$buf32),
    .Q(\Y[1] [0])
);

FILL FILL_3__9416_ (
);

FILL FILL_0__6874_ (
);

DFFPOSX1 _8980_ (
    .D(\Y[2] [3]),
    .CLK(clk_bF$buf44),
    .Q(\u_fir_pe2.rYin [3])
);

FILL FILL_0__6454_ (
);

OAI22X1 _8560_ (
    .A(_1848_),
    .B(_1995_),
    .C(_1918_),
    .D(_1996_),
    .Y(_1997_)
);

INVX1 _8140_ (
    .A(\X[2] [2]),
    .Y(_2364_)
);

AOI22X1 _11197_ (
    .A(_4227_),
    .B(_4393_),
    .C(_4319_),
    .D(_4315_),
    .Y(_4394_)
);

FILL FILL_2__7833_ (
);

FILL FILL_2__7413_ (
);

FILL FILL_1__13280_ (
);

FILL FILL_2__11659_ (
);

FILL FILL_0__12693_ (
);

FILL FILL_2__11239_ (
);

FILL FILL_0__12273_ (
);

FILL FILL_2__12600_ (
);

FILL FILL_0__7659_ (
);

NAND2X1 _9765_ (
    .A(_3108_),
    .B(_3107_),
    .Y(_3181_[9])
);

OR2X2 _9345_ (
    .A(_2698_),
    .B(_2697_),
    .Y(_2703_)
);

FILL FILL_2__8618_ (
);

FILL FILL_0__8600_ (
);

FILL FILL_0__13058_ (
);

DFFPOSX1 _13343_ (
    .D(_6369_[5]),
    .CLK(clk_bF$buf46),
    .Q(\Y[7] [5])
);

FILL FILL_1__6615_ (
);

FILL FILL_1__9087_ (
);

FILL FILL_0__9805_ (
);

FILL FILL_3__10312_ (
);

FILL FILL_2__8791_ (
);

FILL FILL_2__8371_ (
);

FILL FILL_2__12197_ (
);

AOI21X1 _7831_ (
    .A(_1284_),
    .B(_1288_),
    .C(_1258_),
    .Y(_1346_)
);

OR2X2 _7411_ (
    .A(_930_),
    .B(_928_),
    .Y(_931_)
);

FILL FILL_0__8197_ (
);

NAND3X1 _10888_ (
    .A(_4080_),
    .B(_4076_),
    .C(_4082_),
    .Y(_4089_)
);

OAI21X1 _10468_ (
    .A(_3692_),
    .B(_3695_),
    .C(_3740_),
    .Y(_3743_)
);

INVX1 _10048_ (
    .A(_3327_),
    .Y(_3328_)
);

FILL FILL_3__11937_ (
);

FILL FILL_1__12971_ (
);

FILL FILL_1__12551_ (
);

FILL FILL_1__12131_ (
);

FILL FILL_2__9996_ (
);

FILL FILL_2__9576_ (
);

FILL FILL_0__11964_ (
);

FILL FILL_2__9156_ (
);

FILL FILL_0__11544_ (
);

FILL FILL_0__11124_ (
);

INVX1 _8616_ (
    .A(_2051_),
    .Y(_2052_)
);

FILL FILL_1__7993_ (
);

FILL FILL_1__7573_ (
);

FILL FILL_1__7153_ (
);

FILL FILL_3__7499_ (
);

FILL FILL_1__13336_ (
);

FILL FILL_3__8860_ (
);

FILL FILL_0__12749_ (
);

OAI21X1 _12614_ (
    .A(_6357_),
    .B(_5653_),
    .C(_5654_),
    .Y(_5655_)
);

FILL FILL_0__12329_ (
);

FILL FILL_1__8778_ (
);

FILL FILL_3__11690_ (
);

FILL FILL_1__8358_ (
);

FILL FILL_3__11270_ (
);

FILL FILL_2__10683_ (
);

FILL FILL_2__10263_ (
);

FILL FILL_3__9645_ (
);

FILL FILL_0__6683_ (
);

FILL FILL_2__7642_ (
);

FILL FILL_3__12055_ (
);

FILL FILL_2__11888_ (
);

FILL FILL_2__11468_ (
);

FILL FILL_2__11048_ (
);

FILL FILL_0__12082_ (
);

FILL FILL_0__7888_ (
);

AND2X2 _9994_ (
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3275_)
);

FILL FILL_0__7468_ (
);

AOI21X1 _9574_ (
    .A(_2806_),
    .B(_2798_),
    .C(_2876_),
    .Y(_2929_)
);

FILL FILL_0__7048_ (
);

NAND3X1 _9154_ (
    .A(_2444_),
    .B(_2508_),
    .C(_2509_),
    .Y(_2515_)
);

FILL FILL_1__11822_ (
);

FILL FILL_1__11402_ (
);

FILL FILL_2__8847_ (
);

FILL FILL_2__8427_ (
);

FILL FILL_0__10815_ (
);

FILL FILL_2__8007_ (
);

FILL FILL_0__13287_ (
);

OAI21X1 _13152_ (
    .A(_6142_),
    .B(_6155_),
    .C(_6159_),
    .Y(_6185_)
);

FILL FILL_1__6844_ (
);

FILL FILL_1__6424_ (
);

FILL FILL_1__12607_ (
);

FILL FILL_0__9614_ (
);

FILL FILL_3__7711_ (
);

FILL FILL_1__7629_ (
);

FILL FILL_3__10541_ (
);

FILL FILL_2__8180_ (
);

NAND2X1 _6699_ (
    .A(_296_),
    .B(_295_),
    .Y(_297_)
);

NAND3X1 _7640_ (
    .A(_1112_),
    .B(_1143_),
    .C(_1148_),
    .Y(_1158_)
);

DFFPOSX1 _7220_ (
    .D(Xin_5_bF$buf1),
    .CLK(clk_bF$buf16),
    .Q(\X[1] [5])
);

INVX1 _10697_ (
    .A(_3960_),
    .Y(_3961_)
);

OAI21X1 _10277_ (
    .A(_3554_),
    .B(_3551_),
    .C(_3487_),
    .Y(_3555_)
);

FILL FILL_2__6913_ (
);

FILL FILL_1__12780_ (
);

FILL FILL_3__11326_ (
);

FILL FILL_1__12360_ (
);

FILL FILL_2__9385_ (
);

FILL FILL_0__11773_ (
);

FILL FILL_2__10319_ (
);

FILL FILL_0__11353_ (
);

FILL FILL_0__6739_ (
);

NOR2X1 _8845_ (
    .A(_2267_),
    .B(_2268_),
    .Y(_2269_)
);

AND2X2 _8425_ (
    .A(_1815_),
    .B(_1812_),
    .Y(_1864_)
);

AND2X2 _8005_ (
    .A(\u_fir_pe1.rYin [9]),
    .B(\u_fir_pe1.mul [9]),
    .Y(_1509_)
);

FILL FILL_1__7382_ (
);

FILL FILL_1__13145_ (
);

FILL FILL_0__12978_ (
);

AOI21X1 _12843_ (
    .A(_5845_),
    .B(_5846_),
    .C(_5803_),
    .Y(_5881_)
);

FILL FILL_0__12558_ (
);

FILL FILL_0__12138_ (
);

NOR2X1 _12423_ (
    .A(\u_fir_pe6.rYin [12]),
    .B(\u_fir_pe6.mul [12]),
    .Y(_5527_)
);

NAND3X1 _12003_ (
    .A(_5106_),
    .B(_5108_),
    .C(_5110_),
    .Y(_5121_)
);

FILL FILL_1__8587_ (
);

FILL FILL_1__8167_ (
);

FILL FILL_2__10492_ (
);

FILL FILL_2__10072_ (
);

FILL FILL_3__9034_ (
);

INVX1 _13208_ (
    .A(\u_fir_pe7.rYin [4]),
    .Y(_6234_)
);

FILL FILL_0__6492_ (
);

FILL FILL_2__7871_ (
);

FILL FILL_2__7451_ (
);

FILL FILL_3__12284_ (
);

FILL FILL_2__7031_ (
);

FILL FILL_2__11697_ (
);

FILL FILL_2__11277_ (
);

AOI21X1 _6911_ (
    .A(_455_),
    .B(_458_),
    .C(_506_),
    .Y(_507_)
);

FILL FILL_0__7697_ (
);

FILL FILL_0__7277_ (
);

NAND3X1 _9383_ (
    .A(_2713_),
    .B(_2731_),
    .C(_2727_),
    .Y(_2741_)
);

FILL FILL_1__11211_ (
);

FILL FILL_2__8656_ (
);

FILL FILL_2__8236_ (
);

FILL FILL_0__10624_ (
);

FILL FILL_3__13069_ (
);

FILL FILL_0__10204_ (
);

FILL FILL_0__13096_ (
);

DFFPOSX1 _13381_ (
    .D(_6373_[3]),
    .CLK(clk_bF$buf27),
    .Q(\u_fir_pe7.mul [3])
);

FILL FILL_1__6653_ (
);

FILL FILL_2__13003_ (
);

FILL FILL_1__12836_ (
);

FILL FILL_1__12416_ (
);

FILL FILL_3__7940_ (
);

FILL FILL_0__9423_ (
);

FILL FILL_0__11829_ (
);

FILL FILL_0__11409_ (
);

FILL FILL_3__7100_ (
);

FILL FILL_1__7858_ (
);

FILL FILL_3__10770_ (
);

FILL FILL_1__7438_ (
);

FILL FILL_1__7018_ (
);

FILL FILL_3__8725_ (
);

INVX1 _10086_ (
    .A(_3284_),
    .Y(_3366_)
);

FILL FILL_2__6722_ (
);

FILL FILL_3__11555_ (
);

FILL FILL_2__10968_ (
);

FILL FILL_2__10548_ (
);

FILL FILL_2__9194_ (
);

FILL FILL_0__11582_ (
);

FILL FILL_2__10128_ (
);

FILL FILL_0__11162_ (
);

FILL FILL_0__6968_ (
);

FILL FILL_0__6548_ (
);

INVX1 _8654_ (
    .A(_2054_),
    .Y(_2090_)
);

NAND3X1 _8234_ (
    .A(_1664_),
    .B(_1672_),
    .C(_1674_),
    .Y(_1675_)
);

FILL FILL_1__7191_ (
);

FILL FILL_1__10902_ (
);

FILL FILL_2__7927_ (
);

FILL FILL_2__7507_ (
);

FILL FILL_0__12787_ (
);

NAND3X1 _12652_ (
    .A(_5680_),
    .B(_5684_),
    .C(_5686_),
    .Y(_5693_)
);

FILL FILL_0__12367_ (
);

INVX1 _12232_ (
    .A(_5308_),
    .Y(_5346_)
);

DFFPOSX1 _9859_ (
    .D(\Y[3] [5]),
    .CLK(clk_bF$buf53),
    .Q(\u_fir_pe3.rYin [5])
);

AND2X2 _9439_ (
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2796_)
);

NOR2X1 _9019_ (
    .A(_3161_),
    .B(_3169_),
    .Y(_3171_)
);

FILL FILL_1__8396_ (
);

FILL FILL_3__9683_ (
);

FILL FILL_3__9263_ (
);

NOR2X1 _13017_ (
    .A(_6052_),
    .B(_5995_),
    .Y(_6053_)
);

FILL FILL_1__6709_ (
);

FILL FILL_2__7680_ (
);

FILL FILL_2__7260_ (
);

FILL FILL_2__11086_ (
);

NAND2X1 _6720_ (
    .A(Xin[3]),
    .B(gnd),
    .Y(_318_)
);

FILL FILL_1__10499_ (
);

FILL FILL_1__10079_ (
);

FILL FILL_0__7086_ (
);

INVX1 _9192_ (
    .A(_2551_),
    .Y(_2552_)
);

FILL FILL_3__10826_ (
);

FILL FILL_1__11860_ (
);

FILL FILL_3__10406_ (
);

FILL FILL_1__11440_ (
);

FILL FILL_1__11020_ (
);

FILL FILL_2__8885_ (
);

FILL FILL_2__8465_ (
);

FILL FILL_0__10853_ (
);

FILL FILL_0__10433_ (
);

FILL FILL_3__13298_ (
);

FILL FILL_2__8045_ (
);

FILL FILL_0__10013_ (
);

NOR2X1 _13190_ (
    .A(_6218_),
    .B(_6217_),
    .Y(_6369_[1])
);

NAND2X1 _7925_ (
    .A(_1428_),
    .B(_1433_),
    .Y(_1434_)
);

AND2X2 _7505_ (
    .A(\X[1] [3]),
    .B(gnd),
    .Y(_1024_)
);

FILL FILL_1__6882_ (
);

FILL FILL_1__6462_ (
);

FILL FILL_2__13232_ (
);

FILL FILL_3__6388_ (
);

FILL FILL_1__12645_ (
);

FILL FILL_1__12225_ (
);

FILL FILL_0__9652_ (
);

FILL FILL_0__9232_ (
);

NAND3X1 _11923_ (
    .A(_5021_),
    .B(_5035_),
    .C(_5038_),
    .Y(_5042_)
);

NAND3X1 _11503_ (
    .A(_4686_),
    .B(_4683_),
    .C(_4646_),
    .Y(_4687_)
);

FILL FILL_0__11218_ (
);

FILL FILL_1__7667_ (
);

AOI21X1 _12708_ (
    .A(_5742_),
    .B(_5744_),
    .C(_5735_),
    .Y(_5748_)
);

FILL FILL_2__6951_ (
);

FILL FILL254550x198150 (
);

FILL FILL_3__11784_ (
);

FILL FILL_2__6531_ (
);

FILL FILL_2__10777_ (
);

FILL FILL_2__10357_ (
);

FILL FILL_0__11391_ (
);

FILL FILL_1__9813_ (
);

FILL FILL_3__9739_ (
);

FILL FILL_0__6777_ (
);

NOR2X1 _8883_ (
    .A(\u_fir_pe2.rYin [9]),
    .B(\u_fir_pe2.mul [9]),
    .Y(_2307_)
);

OAI21X1 _8463_ (
    .A(_1819_),
    .B(_1824_),
    .C(_1823_),
    .Y(_1901_)
);

OAI21X1 _8043_ (
    .A(_1539_),
    .B(_1540_),
    .C(_1544_),
    .Y(_1546_)
);

FILL FILL_2__7736_ (
);

FILL FILL_3__12569_ (
);

FILL FILL_2__7316_ (
);

FILL FILL_3__12149_ (
);

FILL FILL_1__13183_ (
);

NAND3X1 _12881_ (
    .A(_5917_),
    .B(_5918_),
    .C(_5916_),
    .Y(_5919_)
);

FILL FILL_0__12596_ (
);

FILL FILL_0__12176_ (
);

DFFPOSX1 _12461_ (
    .D(_5571_[0]),
    .CLK(clk_bF$buf49),
    .Q(_6377_[0])
);

AND2X2 _12041_ (
    .A(_5149_),
    .B(_5154_),
    .Y(_5159_)
);

FILL FILL_2__12923_ (
);

NAND2X1 _9668_ (
    .A(_3019_),
    .B(_3013_),
    .Y(_3187_[14])
);

NAND2X1 _9248_ (
    .A(_2604_),
    .B(_2606_),
    .Y(_2607_)
);

FILL FILL_1__11916_ (
);

FILL FILL_0__8923_ (
);

FILL FILL_0__8503_ (
);

FILL FILL_0__10909_ (
);

FILL FILL_3__6600_ (
);

INVX1 _13246_ (
    .A(\u_fir_pe7.rYin [8]),
    .Y(_6269_)
);

FILL FILL_1__6938_ (
);

FILL FILL_1__6518_ (
);

FILL FILL_0__9708_ (
);

FILL FILL_3__7805_ (
);

FILL FILL_3__10635_ (
);

FILL FILL_2__8694_ (
);

FILL FILL_2__8274_ (
);

FILL FILL_0__10662_ (
);

FILL FILL_0__10242_ (
);

NAND2X1 _7734_ (
    .A(_1239_),
    .B(_1246_),
    .Y(_1250_)
);

INVX1 _7314_ (
    .A(_835_),
    .Y(_836_)
);

FILL FILL_1__6691_ (
);

FILL FILL_2__13041_ (
);

FILL FILL_1__12874_ (
);

FILL FILL_1__12454_ (
);

FILL FILL_1__12034_ (
);

FILL FILL_2__9899_ (
);

FILL FILL_2__9479_ (
);

FILL FILL_0__9461_ (
);

FILL FILL_0__11867_ (
);

FILL FILL_2__9059_ (
);

FILL FILL_0__9041_ (
);

INVX1 _11732_ (
    .A(_4852_),
    .Y(_4853_)
);

FILL FILL_0__11447_ (
);

FILL FILL_0__11027_ (
);

OAI21X1 _11312_ (
    .A(_4059_),
    .B(_4290_),
    .C(_4464_),
    .Y(_4507_)
);

NAND2X1 _8939_ (
    .A(_2358_),
    .B(_2352_),
    .Y(_2362_)
);

AOI21X1 _8519_ (
    .A(_1951_),
    .B(_1956_),
    .C(_1895_),
    .Y(_1957_)
);

FILL FILL_1__7896_ (
);

FILL FILL_1__7476_ (
);

FILL FILL_1__7056_ (
);

FILL FILL_1__13239_ (
);

AND2X2 _12937_ (
    .A(_5973_),
    .B(_5970_),
    .Y(_5974_)
);

FILL FILL_3__8343_ (
);

NAND2X1 _12517_ (
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_6268_)
);

FILL FILL_2__6760_ (
);

FILL FILL_3__11173_ (
);

FILL FILL_2__10586_ (
);

FILL FILL_2__10166_ (
);

FILL FILL_1__9622_ (
);

FILL FILL_1__9202_ (
);

FILL FILL_3__9968_ (
);

FILL FILL_3__9128_ (
);

FILL FILL_0__6586_ (
);

AND2X2 _8692_ (
    .A(_2117_),
    .B(_2113_),
    .Y(_2127_)
);

NAND3X1 _8272_ (
    .A(_1648_),
    .B(_1711_),
    .C(_1712_),
    .Y(_1713_)
);

FILL FILL_1__10940_ (
);

FILL FILL_1__10520_ (
);

FILL FILL_1__10100_ (
);

FILL FILL_2__7965_ (
);

FILL FILL_3__12798_ (
);

FILL FILL_2__7545_ (
);

FILL FILL_3__12378_ (
);

FILL FILL_2__7125_ (
);

NAND3X1 _12690_ (
    .A(_5718_),
    .B(_5727_),
    .C(_5729_),
    .Y(_5730_)
);

NAND2X1 _12270_ (
    .A(_5381_),
    .B(_5382_),
    .Y(_5383_)
);

FILL FILL_2__12732_ (
);

FILL FILL_2__12312_ (
);

NAND2X1 _9897_ (
    .A(_3968_),
    .B(_3948_),
    .Y(_3969_)
);

INVX1 _9477_ (
    .A(_2755_),
    .Y(_2834_)
);

NOR2X1 _9057_ (
    .A(_2418_),
    .B(_2417_),
    .Y(_2419_)
);

FILL FILL_1__11725_ (
);

FILL FILL_1__11305_ (
);

FILL FILL_0__8732_ (
);

FILL FILL_0__8312_ (
);

NAND3X1 _13055_ (
    .A(_6074_),
    .B(_6080_),
    .C(_6038_),
    .Y(_6090_)
);

FILL FILL_1__6747_ (
);

FILL FILL253350x248550 (
);

FILL FILL_0__9937_ (
);

FILL FILL_0__9517_ (
);

FILL FILL_3__7614_ (
);

FILL FILL_3__10024_ (
);

FILL FILL_0__10891_ (
);

FILL FILL_0__10471_ (
);

FILL FILL_0__10051_ (
);

FILL FILL_3__8819_ (
);

OR2X2 _7963_ (
    .A(_1461_),
    .B(_1466_),
    .Y(_1468_)
);

AOI21X1 _7543_ (
    .A(_949_),
    .B(_968_),
    .C(_1061_),
    .Y(_1062_)
);

NAND2X1 _7123_ (
    .A(_705_),
    .B(_706_),
    .Y(_707_)
);

FILL FILL_2__13270_ (
);

FILL FILL_2__6816_ (
);

FILL FILL_3__11649_ (
);

FILL FILL_1__12683_ (
);

FILL FILL_1__12263_ (
);

FILL FILL_0__9690_ (
);

FILL FILL_2__9288_ (
);

FILL FILL_0__9270_ (
);

NAND2X1 _11961_ (
    .A(_5078_),
    .B(_5077_),
    .Y(_5079_)
);

FILL FILL_0__11676_ (
);

NAND2X1 _11541_ (
    .A(_4720_),
    .B(_4713_),
    .Y(_4724_)
);

FILL FILL_0__11256_ (
);

NAND2X1 _11121_ (
    .A(_4310_),
    .B(_4318_),
    .Y(_4319_)
);

OAI21X1 _8748_ (
    .A(_1970_),
    .B(_2181_),
    .C(_2153_),
    .Y(_2182_)
);

OAI21X1 _8328_ (
    .A(_1763_),
    .B(_1764_),
    .C(_1749_),
    .Y(_1768_)
);

FILL FILL_1__7285_ (
);

FILL FILL_1__13048_ (
);

FILL FILL_3__8572_ (
);

NOR2X1 _12746_ (
    .A(_5783_),
    .B(_5785_),
    .Y(_6375_[6])
);

NOR2X1 _12326_ (
    .A(\u_fir_pe6.rYin [3]),
    .B(\u_fir_pe6.mul [3]),
    .Y(_5433_)
);

FILL FILL_0__13402_ (
);

FILL FILL_2__10395_ (
);

FILL FILL_1__9431_ (
);

FILL FILL_1__9011_ (
);

FILL FILL_3__9777_ (
);

FILL FILL_3__9357_ (
);

FILL FILL_0__6395_ (
);

DFFPOSX1 _8081_ (
    .D(_1587_[5]),
    .CLK(clk_bF$buf38),
    .Q(\Y[2] [5])
);

FILL FILL_2__7774_ (
);

FILL FILL_2__7354_ (
);

NAND2X1 _6814_ (
    .A(_401_),
    .B(_410_),
    .Y(_411_)
);

FILL FILL_2__12961_ (
);

FILL FILL_2__12541_ (
);

FILL FILL_2__12121_ (
);

NAND2X1 _9286_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .Y(_2645_)
);

FILL FILL_1__11954_ (
);

FILL FILL_1__11534_ (
);

FILL FILL_1__11114_ (
);

FILL FILL_2__8559_ (
);

FILL FILL_0__8541_ (
);

FILL FILL_0__10947_ (
);

FILL FILL_2__8139_ (
);

FILL FILL_0__10527_ (
);

INVX1 _10812_ (
    .A(_4013_),
    .Y(_4014_)
);

FILL FILL_0__10107_ (
);

NAND2X1 _13284_ (
    .A(_6307_),
    .B(_6302_),
    .Y(_6308_)
);

FILL FILL_2__9920_ (
);

FILL FILL_2__9500_ (
);

FILL FILL_1__6976_ (
);

FILL FILL_1__6556_ (
);

FILL FILL_2__13326_ (
);

FILL FILL_1__12739_ (
);

FILL FILL_1__12319_ (
);

FILL FILL_0__9746_ (
);

FILL FILL_0__9326_ (
);

FILL FILL_3__7423_ (
);

FILL FILL_3__10253_ (
);

FILL FILL_0__10280_ (
);

FILL FILL_1__8702_ (
);

FILL FILL_3__8208_ (
);

NAND3X1 _7772_ (
    .A(_1285_),
    .B(_1287_),
    .C(_1286_),
    .Y(_1288_)
);

OAI21X1 _7352_ (
    .A(_1575_),
    .B(_871_),
    .C(_872_),
    .Y(_873_)
);

FILL FILL_3__11878_ (
);

FILL FILL_2__6625_ (
);

FILL FILL_3__11038_ (
);

FILL FILL_1__12072_ (
);

FILL FILL_2__9097_ (
);

AOI21X1 _11770_ (
    .A(_4882_),
    .B(_4878_),
    .C(_4864_),
    .Y(_4891_)
);

FILL FILL_0__11485_ (
);

FILL FILL_0__11065_ (
);

AOI21X1 _11350_ (
    .A(_4541_),
    .B(_4442_),
    .C(_4543_),
    .Y(_4544_)
);

FILL FILL_1__9907_ (
);

FILL FILL_2__11812_ (
);

DFFPOSX1 _8977_ (
    .D(\Y[2] [0]),
    .CLK(clk_bF$buf17),
    .Q(\u_fir_pe2.rYin [0])
);

NOR2X1 _8557_ (
    .A(_1992_),
    .B(_1993_),
    .Y(_1994_)
);

NOR2X1 _8137_ (
    .A(_2283_),
    .B(_2325_),
    .Y(_2334_)
);

FILL FILL_1__7094_ (
);

FILL FILL_1__10805_ (
);

FILL FILL_0__7812_ (
);

FILL FILL_1__13277_ (
);

AOI21X1 _12975_ (
    .A(_5932_),
    .B(_5934_),
    .C(_6011_),
    .Y(_6012_)
);

NAND2X1 _12555_ (
    .A(_6360_),
    .B(_5597_),
    .Y(_5598_)
);

NAND3X1 _12135_ (
    .A(_5249_),
    .B(_5246_),
    .C(_5250_),
    .Y(_5251_)
);

FILL FILL_0__13211_ (
);

FILL FILL_1__8299_ (
);

FILL FILL_1__9660_ (
);

FILL FILL_1__9240_ (
);

FILL FILL_3__9586_ (
);

FILL FILL_2__7583_ (
);

FILL FILL_2__7163_ (
);

NAND2X1 _6623_ (
    .A(_218_),
    .B(_221_),
    .Y(_222_)
);

FILL FILL_2__12770_ (
);

FILL FILL_2__12350_ (
);

OAI21X1 _9095_ (
    .A(_2444_),
    .B(_2456_),
    .C(_2450_),
    .Y(_2457_)
);

FILL FILL_1__11763_ (
);

FILL FILL_1__11343_ (
);

FILL FILL_0__8770_ (
);

FILL FILL_2__8788_ (
);

FILL FILL_0__8350_ (
);

FILL FILL_2__8368_ (
);

FILL FILL_0__10336_ (
);

NAND2X1 _10621_ (
    .A(_3863_),
    .B(_3875_),
    .Y(_3884_)
);

AOI21X1 _10201_ (
    .A(_3475_),
    .B(_3474_),
    .C(_3376_),
    .Y(_3480_)
);

AOI21X1 _13093_ (
    .A(_6066_),
    .B(_6070_),
    .C(_6040_),
    .Y(_6128_)
);

NAND3X1 _7828_ (
    .A(_1340_),
    .B(_1342_),
    .C(_1341_),
    .Y(_1343_)
);

AND2X2 _7408_ (
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_928_)
);

FILL FILL_1__6785_ (
);

FILL FILL_2__13135_ (
);

FILL FILL_1__12968_ (
);

FILL FILL_1__12548_ (
);

FILL FILL_1__12128_ (
);

FILL FILL_0__9975_ (
);

FILL FILL_0__9555_ (
);

FILL FILL_3__7652_ (
);

FILL FILL_0__9135_ (
);

NAND2X1 _11826_ (
    .A(vdd),
    .B(\X[7] [4]),
    .Y(_4946_)
);

NAND2X1 _11406_ (
    .A(_4598_),
    .B(_4595_),
    .Y(_4781_[13])
);

FILL FILL_0__12902_ (
);

FILL FILL_3__10482_ (
);

FILL FILL_1__8931_ (
);

FILL FILL_1__8511_ (
);

FILL FILL_3__8437_ (
);

AOI21X1 _7581_ (
    .A(_1063_),
    .B(_1064_),
    .C(_1021_),
    .Y(_1099_)
);

NOR2X1 _7161_ (
    .A(\u_fir_pe0.rYin [12]),
    .B(\u_fir_pe0.mul [12]),
    .Y(_745_)
);

FILL FILL_2__6854_ (
);

FILL FILL_2__6434_ (
);

FILL FILL_3__11267_ (
);

FILL FILL_0__11294_ (
);

FILL FILL_1__9716_ (
);

FILL FILL_2__11201_ (
);

NOR3X1 _8786_ (
    .A(_2217_),
    .B(_2185_),
    .C(_2203_),
    .Y(_2218_)
);

INVX1 _8366_ (
    .A(_1804_),
    .Y(_1805_)
);

FILL FILL_1__10614_ (
);

FILL FILL_0__7621_ (
);

FILL FILL_2__7639_ (
);

FILL FILL_1__13086_ (
);

OAI21X1 _12784_ (
    .A(_5668_),
    .B(_5653_),
    .C(_5737_),
    .Y(_5823_)
);

FILL FILL_3__8190_ (
);

FILL FILL_0__12079_ (
);

OAI21X1 _12364_ (
    .A(_5465_),
    .B(_5466_),
    .C(_5462_),
    .Y(_5467_)
);

FILL FILL_3__13413_ (
);

FILL FILL_2__12826_ (
);

FILL FILL_2__12406_ (
);

FILL FILL_0__13020_ (
);

FILL FILL_1__11819_ (
);

FILL FILL_0__8826_ (
);

FILL FILL_3__6923_ (
);

FILL FILL_0__8406_ (
);

FILL FILL_3__9395_ (
);

OR2X2 _13149_ (
    .A(_6180_),
    .B(_6173_),
    .Y(_6182_)
);

FILL FILL_2__7392_ (
);

FILL FILL_3__7708_ (
);

OAI21X1 _6852_ (
    .A(_447_),
    .B(_448_),
    .C(_444_),
    .Y(_449_)
);

INVX1 _6432_ (
    .A(_33_),
    .Y(_34_)
);

FILL FILL_1__11992_ (
);

FILL FILL_1__11572_ (
);

FILL FILL_3__10118_ (
);

FILL FILL_1__11152_ (
);

FILL FILL_2__8597_ (
);

FILL FILL_0__10985_ (
);

FILL FILL_2__8177_ (
);

FILL FILL_0__10565_ (
);

NAND2X1 _10850_ (
    .A(_4051_),
    .B(_4045_),
    .Y(_4780_[4])
);

NOR3X1 _10430_ (
    .A(_3493_),
    .B(_3661_),
    .C(_3604_),
    .Y(_3705_)
);

FILL FILL_0__10145_ (
);

OAI21X1 _10010_ (
    .A(_3286_),
    .B(_3287_),
    .C(_3272_),
    .Y(_3291_)
);

INVX1 _7637_ (
    .A(_1068_),
    .Y(_1155_)
);

DFFPOSX1 _7217_ (
    .D(Xin[2]),
    .CLK(clk_bF$buf41),
    .Q(\X[1] [2])
);

FILL FILL_1__6594_ (
);

FILL FILL_1__12777_ (
);

FILL FILL_1__12357_ (
);

FILL FILL_0__9784_ (
);

FILL FILL_3__7881_ (
);

FILL FILL_0__9364_ (
);

DFFPOSX1 _11635_ (
    .D(_4781_[11]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [11])
);

FILL FILL_3__7041_ (
);

NAND2X1 _11215_ (
    .A(_4376_),
    .B(_4379_),
    .Y(_4412_)
);

FILL FILL_0__12711_ (
);

FILL FILL_1__7799_ (
);

FILL FILL_1__7379_ (
);

FILL FILL_1__8740_ (
);

FILL FILL_1__8320_ (
);

FILL FILL_3__8666_ (
);

NAND3X1 _7390_ (
    .A(_898_),
    .B(_902_),
    .C(_904_),
    .Y(_911_)
);

FILL FILL_2__6663_ (
);

FILL FILL_3__11496_ (
);

FILL FILL_2__10489_ (
);

FILL FILL_2__10069_ (
);

FILL FILL_1__9945_ (
);

FILL FILL_1__9525_ (
);

FILL FILL_1__9105_ (
);

FILL FILL_2__11850_ (
);

FILL FILL_2__11430_ (
);

FILL FILL_2__11010_ (
);

FILL FILL_0__6489_ (
);

INVX1 _8595_ (
    .A(_1977_),
    .Y(_2032_)
);

NOR2X1 _8175_ (
    .A(_1617_),
    .B(_1616_),
    .Y(_2388_[3])
);

FILL FILL_1__10843_ (
);

FILL FILL_1__10423_ (
);

FILL FILL_1__10003_ (
);

FILL FILL_2__7868_ (
);

FILL FILL_0__7850_ (
);

FILL FILL_2__7448_ (
);

FILL FILL_0__7430_ (
);

FILL FILL_0__7010_ (
);

FILL FILL_2__7028_ (
);

NAND2X1 _12593_ (
    .A(_5628_),
    .B(_5631_),
    .Y(_5635_)
);

AOI21X1 _12173_ (
    .A(_5237_),
    .B(_5240_),
    .C(_5288_),
    .Y(_5289_)
);

FILL FILL_3__13222_ (
);

AOI21X1 _6908_ (
    .A(_431_),
    .B(_437_),
    .C(_503_),
    .Y(_504_)
);

FILL FILL_2__12635_ (
);

FILL FILL_2__12215_ (
);

FILL FILL_1__11208_ (
);

FILL FILL_0__8635_ (
);

FILL FILL_0__8215_ (
);

NAND3X1 _10906_ (
    .A(_4106_),
    .B(_4039_),
    .C(_4042_),
    .Y(_4107_)
);

DFFPOSX1 _13378_ (
    .D(_6370_[0]),
    .CLK(clk_bF$buf24),
    .Q(\u_fir_pe7.mul [0])
);

NAND3X1 _6661_ (
    .A(_239_),
    .B(_253_),
    .C(_256_),
    .Y(_260_)
);

FILL FILL_3__10767_ (
);

FILL FILL_3__10347_ (
);

FILL FILL_1__11381_ (
);

FILL FILL_0__10794_ (
);

FILL FILL_0__10374_ (
);

FILL FILL_2__10701_ (
);

OR2X2 _7866_ (
    .A(_1378_),
    .B(_1376_),
    .Y(_1380_)
);

AOI21X1 _7446_ (
    .A(_960_),
    .B(_962_),
    .C(_953_),
    .Y(_966_)
);

AND2X2 _7026_ (
    .A(_596_),
    .B(_595_),
    .Y(_618_)
);

FILL FILL_2__13173_ (
);

FILL FILL_2__6719_ (
);

FILL FILL_0__6701_ (
);

FILL FILL_1__12586_ (
);

FILL FILL_1__12166_ (
);

FILL FILL_0__11999_ (
);

FILL FILL_0__9593_ (
);

FILL FILL_0__9173_ (
);

NAND3X1 _11864_ (
    .A(_4977_),
    .B(_4978_),
    .C(_4983_),
    .Y(_4984_)
);

FILL FILL_0__11579_ (
);

FILL FILL_3__7270_ (
);

NAND2X1 _11444_ (
    .A(_4628_),
    .B(_4631_),
    .Y(_4775_[2])
);

FILL FILL_0__11159_ (
);

NAND2X1 _11024_ (
    .A(_4217_),
    .B(_4222_),
    .Y(_4223_)
);

FILL FILL_2__11906_ (
);

FILL FILL_0__12940_ (
);

FILL FILL_0__12520_ (
);

FILL FILL_0__12100_ (
);

FILL FILL_1__7188_ (
);

FILL FILL_0__7906_ (
);

FILL FILL_3__8895_ (
);

NAND3X1 _12649_ (
    .A(_5605_),
    .B(_5685_),
    .C(_5689_),
    .Y(_5690_)
);

FILL FILL_3__8055_ (
);

OAI21X1 _12229_ (
    .A(_5087_),
    .B(_5261_),
    .C(_5305_),
    .Y(_5343_)
);

FILL FILL_0__13305_ (
);

FILL FILL_2__6892_ (
);

FILL FILL_2__6472_ (
);

FILL FILL_2__10298_ (
);

FILL FILL_1__9754_ (
);

FILL FILL_1__9334_ (
);

FILL FILL_1__10652_ (
);

FILL FILL_1__10232_ (
);

FILL FILL_2__7677_ (
);

FILL FILL_2__7257_ (
);

NAND2X1 _6717_ (
    .A(_310_),
    .B(_314_),
    .Y(_315_)
);

FILL FILL_2__12864_ (
);

FILL FILL_2__12444_ (
);

FILL FILL_2__12024_ (
);

AND2X2 _9189_ (
    .A(gnd),
    .B(\X[3] [4]),
    .Y(_2549_)
);

FILL FILL_1__11857_ (
);

FILL FILL_1__11437_ (
);

FILL FILL_1__11017_ (
);

FILL FILL_0__8864_ (
);

FILL FILL_0__8444_ (
);

FILL FILL_3__6541_ (
);

DFFPOSX1 _10715_ (
    .D(_3978_[8]),
    .CLK(clk_bF$buf30),
    .Q(\Y[5] [8])
);

FILL FILL_0__8024_ (
);

NAND2X1 _13187_ (
    .A(_6210_),
    .B(_6215_),
    .Y(_6216_)
);

FILL FILL_2__9823_ (
);

FILL FILL_2__9403_ (
);

FILL FILL_1__6879_ (
);

FILL FILL_1__6459_ (
);

FILL FILL_2__13229_ (
);

FILL FILL_1__7820_ (
);

FILL FILL_1__7400_ (
);

FILL FILL_0__9649_ (
);

FILL FILL_3__7746_ (
);

FILL FILL_0__9229_ (
);

FILL FILL_3__7326_ (
);

NAND3X1 _6890_ (
    .A(_407_),
    .B(_485_),
    .C(_415_),
    .Y(_486_)
);

INVX1 _6470_ (
    .A(_70_),
    .Y(_71_)
);

FILL FILL_3__10996_ (
);

FILL FILL_3__10576_ (
);

FILL FILL_1__11190_ (
);

FILL FILL_0__10183_ (
);

FILL FILL_1__8605_ (
);

FILL FILL_2__10930_ (
);

FILL FILL_2__10510_ (
);

AND2X2 _7675_ (
    .A(_1191_),
    .B(_1188_),
    .Y(_1192_)
);

NAND2X1 _7255_ (
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_1486_)
);

FILL FILL_0__6930_ (
);

FILL FILL_2__6948_ (
);

FILL FILL_2__6528_ (
);

FILL FILL_0__6510_ (
);

FILL FILL_1__12395_ (
);

NAND3X1 _11673_ (
    .A(_5570_),
    .B(_4795_),
    .C(_4791_),
    .Y(_4796_)
);

FILL FILL_0__11388_ (
);

OAI22X1 _11253_ (
    .A(_4402_),
    .B(_4290_),
    .C(_4010_),
    .D(_4401_),
    .Y(_4449_)
);

FILL FILL_3__12722_ (
);

FILL FILL_2__11715_ (
);

FILL FILL_0__7715_ (
);

NAND3X1 _9821_ (
    .A(_3158_),
    .B(_3164_),
    .C(_3159_),
    .Y(_3165_)
);

AOI21X1 _9401_ (
    .A(_2669_),
    .B(_2668_),
    .C(_2600_),
    .Y(_2759_)
);

AOI21X1 _12878_ (
    .A(_5825_),
    .B(_5828_),
    .C(_5834_),
    .Y(_5916_)
);

FILL FILL_3__8284_ (
);

NOR2X1 _12458_ (
    .A(_5559_),
    .B(_5502_),
    .Y(_5574_[1])
);

NAND2X1 _12038_ (
    .A(_5155_),
    .B(_5079_),
    .Y(_5156_)
);

FILL FILL_0__13114_ (
);

FILL FILL_1__9983_ (
);

FILL FILL_1__9563_ (
);

FILL FILL_1__9143_ (
);

FILL FILL_3__9069_ (
);

FILL FILL_1__10881_ (
);

FILL FILL_1__10461_ (
);

FILL FILL_1__10041_ (
);

FILL FILL_2__7486_ (
);

FILL FILL_2__7066_ (
);

NAND2X1 _6946_ (
    .A(_540_),
    .B(_539_),
    .Y(_541_)
);

INVX1 _6526_ (
    .A(_67_),
    .Y(_127_)
);

FILL FILL_2__12673_ (
);

FILL FILL_2__12253_ (
);

FILL FILL_1__11666_ (
);

FILL FILL_1__11246_ (
);

FILL FILL_0__8673_ (
);

FILL FILL_3__6770_ (
);

FILL FILL_0__8253_ (
);

FILL FILL_0__10659_ (
);

NAND2X1 _10944_ (
    .A(_4072_),
    .B(_4143_),
    .Y(_4144_)
);

NAND2X1 _10524_ (
    .A(_3793_),
    .B(_3796_),
    .Y(_3797_)
);

FILL FILL_0__10239_ (
);

NAND3X1 _10104_ (
    .A(_3378_),
    .B(_3379_),
    .C(_3380_),
    .Y(_3384_)
);

FILL FILL_2__9632_ (
);

FILL FILL_2__9212_ (
);

FILL FILL_1__6688_ (
);

FILL FILL_2__13038_ (
);

FILL FILL_3__7975_ (
);

FILL FILL_0__9458_ (
);

FILL FILL_0__9038_ (
);

NOR3X1 _11729_ (
    .A(_4835_),
    .B(_4802_),
    .C(_4847_),
    .Y(_4850_)
);

FILL FILL_3__7135_ (
);

OAI22X1 _11309_ (
    .A(_4402_),
    .B(_4447_),
    .C(_4503_),
    .D(_4502_),
    .Y(_4504_)
);

FILL FILL_0__12805_ (
);

FILL FILL_1__8834_ (
);

FILL FILL_1__8414_ (
);

NOR2X1 _7484_ (
    .A(_1001_),
    .B(_1003_),
    .Y(_1593_[6])
);

NOR2X1 _7064_ (
    .A(\u_fir_pe0.rYin [3]),
    .B(\u_fir_pe0.mul [3]),
    .Y(_651_)
);

FILL FILL_2__6757_ (
);

OAI21X1 _11482_ (
    .A(_4658_),
    .B(_4659_),
    .C(_4663_),
    .Y(_4665_)
);

FILL FILL_0__11197_ (
);

AOI21X1 _11062_ (
    .A(_4169_),
    .B(_4167_),
    .C(_4260_),
    .Y(_4261_)
);

FILL FILL_3__12951_ (
);

FILL FILL_1__9619_ (
);

FILL FILL_3__12111_ (
);

FILL FILL_2__11944_ (
);

FILL FILL_2__11524_ (
);

FILL FILL_2__11104_ (
);

INVX1 _8689_ (
    .A(_2123_),
    .Y(_2124_)
);

NAND3X1 _8269_ (
    .A(_1647_),
    .B(_1705_),
    .C(_1709_),
    .Y(_1710_)
);

FILL FILL_1__10937_ (
);

FILL FILL_1__10517_ (
);

FILL FILL_0__7944_ (
);

FILL FILL_0__7524_ (
);

INVX1 _9630_ (
    .A(_2957_),
    .Y(_2983_)
);

FILL FILL_0__7104_ (
);

AOI21X1 _9210_ (
    .A(_2473_),
    .B(_2491_),
    .C(_2569_),
    .Y(_2570_)
);

NAND3X1 _12687_ (
    .A(gnd),
    .B(\X[6] [6]),
    .C(_5724_),
    .Y(_5727_)
);

NAND2X1 _12267_ (
    .A(_5379_),
    .B(_5378_),
    .Y(_5380_)
);

FILL FILL_2__8903_ (
);

FILL FILL_3__13316_ (
);

FILL FILL_2__12729_ (
);

FILL FILL_2__12309_ (
);

FILL FILL_1__6900_ (
);

FILL FILL_0__8729_ (
);

FILL FILL_0__8309_ (
);

FILL FILL_3__6406_ (
);

FILL FILL_1__9792_ (
);

FILL FILL_1__9372_ (
);

FILL FILL_3__9298_ (
);

FILL FILL_1__10690_ (
);

FILL FILL_1__10270_ (
);

FILL FILL_2__7295_ (
);

AND2X2 _6755_ (
    .A(_314_),
    .B(_310_),
    .Y(_353_)
);

FILL FILL_2__12062_ (
);

FILL FILL_1__11895_ (
);

FILL FILL_1__11475_ (
);

FILL FILL_1__11055_ (
);

FILL FILL_0__8482_ (
);

FILL FILL_0__10888_ (
);

FILL FILL_0__10468_ (
);

FILL FILL_0__8062_ (
);

DFFPOSX1 _10753_ (
    .D(_3984_[6]),
    .CLK(clk_bF$buf21),
    .Q(\u_fir_pe4.mul [6])
);

NAND3X1 _10333_ (
    .A(_3607_),
    .B(_3608_),
    .C(_3609_),
    .Y(_3610_)
);

FILL FILL_0__10048_ (
);

FILL FILL_2__9441_ (
);

FILL FILL_2__9021_ (
);

FILL FILL_1__6497_ (
);

FILL FILL_2__13267_ (
);

AND2X2 _8901_ (
    .A(_2323_),
    .B(_2324_),
    .Y(_2384_[10])
);

FILL FILL_0__9687_ (
);

FILL FILL_0__9267_ (
);

AND2X2 _11958_ (
    .A(_5076_),
    .B(_5072_),
    .Y(_5578_[7])
);

FILL FILL_3__7364_ (
);

AND2X2 _11538_ (
    .A(_4717_),
    .B(_4720_),
    .Y(_4722_)
);

AND2X2 _11118_ (
    .A(gnd),
    .B(\X[5] [6]),
    .Y(_4316_)
);

FILL FILL_1__13201_ (
);

FILL FILL_0__12614_ (
);

FILL FILL_3__10194_ (
);

FILL FILL_1__8643_ (
);

FILL FILL_1__8223_ (
);

FILL FILL_3__8149_ (
);

NAND2X1 _7293_ (
    .A(_1578_),
    .B(_815_),
    .Y(_816_)
);

FILL FILL_3__9510_ (
);

FILL FILL_2__6986_ (
);

FILL FILL_2__6566_ (
);

AOI21X1 _11291_ (
    .A(_4480_),
    .B(_4486_),
    .C(_4444_),
    .Y(_4487_)
);

FILL FILL_1__9428_ (
);

FILL FILL_3__12340_ (
);

FILL FILL_2__11753_ (
);

FILL FILL_2__11333_ (
);

INVX1 _8498_ (
    .A(_1916_),
    .Y(_1936_)
);

DFFPOSX1 _8078_ (
    .D(_1587_[2]),
    .CLK(clk_bF$buf43),
    .Q(\Y[2] [2])
);

FILL FILL_1__10326_ (
);

FILL FILL_0__7753_ (
);

FILL FILL_0__7333_ (
);

DFFPOSX1 _12496_ (
    .D(\Y[7] [11]),
    .CLK(clk_bF$buf8),
    .Q(\u_fir_pe6.rYin [11])
);

NAND2X1 _12076_ (
    .A(_5183_),
    .B(_5192_),
    .Y(_5193_)
);

FILL FILL_2__8712_ (
);

FILL FILL_2__12958_ (
);

FILL FILL_2__12538_ (
);

FILL FILL_2__12118_ (
);

FILL FILL_0__13152_ (
);

FILL FILL_0__8538_ (
);

FILL FILL_3__6635_ (
);

NOR2X1 _10809_ (
    .A(_4009_),
    .B(_4010_),
    .Y(_4011_)
);

FILL FILL_1__9181_ (
);

FILL FILL_2__9917_ (
);

FILL FILL254550x7350 (
);

FILL FILL_1__7914_ (
);

NAND3X1 _6984_ (
    .A(_562_),
    .B(_572_),
    .C(_575_),
    .Y(_578_)
);

NAND2X1 _6564_ (
    .A(vdd),
    .B(Xin[4]),
    .Y(_164_)
);

FILL FILL_2__12291_ (
);

FILL FILL_1__11284_ (
);

FILL FILL_0__8291_ (
);

FILL FILL_0__10697_ (
);

INVX1 _10982_ (
    .A(_4091_),
    .Y(_4182_)
);

NOR2X1 _10562_ (
    .A(\u_fir_pe4.rYin [2]),
    .B(\u_fir_pe4.mul [2]),
    .Y(_3830_)
);

FILL FILL_0__10277_ (
);

INVX1 _10142_ (
    .A(gnd),
    .Y(_3421_)
);

FILL FILL_2__9670_ (
);

FILL FILL_2__10604_ (
);

FILL FILL_2__9250_ (
);

NAND2X1 _7769_ (
    .A(_1266_),
    .B(_1263_),
    .Y(_1285_)
);

NAND2X1 _7349_ (
    .A(_1497_),
    .B(_869_),
    .Y(_870_)
);

FILL FILL_2__13076_ (
);

FILL FILL_0__6604_ (
);

NAND3X1 _8710_ (
    .A(_2136_),
    .B(_2140_),
    .C(_2144_),
    .Y(_2145_)
);

FILL FILL_1__12069_ (
);

FILL FILL_0__9496_ (
);

FILL FILL_3__7593_ (
);

FILL FILL_0__9076_ (
);

NAND3X1 _11767_ (
    .A(_4883_),
    .B(_4887_),
    .C(_4851_),
    .Y(_4888_)
);

NOR3X1 _11347_ (
    .A(_4487_),
    .B(_4489_),
    .C(_4537_),
    .Y(_4541_)
);

FILL FILL_3__12816_ (
);

FILL FILL_1__13010_ (
);

FILL FILL_2__11809_ (
);

FILL FILL_0__12843_ (
);

FILL FILL_0__12423_ (
);

FILL FILL_0__12003_ (
);

FILL FILL_0__7809_ (
);

INVX1 _9915_ (
    .A(_3928_),
    .Y(_3198_)
);

FILL FILL_1__8872_ (
);

FILL FILL_1__8452_ (
);

FILL FILL_1__8032_ (
);

FILL FILL_3__8378_ (
);

FILL FILL_0__13208_ (
);

FILL FILL_2__6795_ (
);

FILL FILL_1__9657_ (
);

FILL FILL_1__9237_ (
);

FILL FILL_2__11982_ (
);

FILL FILL_2__11562_ (
);

FILL FILL_2__11142_ (
);

FILL FILL_1__10975_ (
);

FILL FILL_1__10555_ (
);

FILL FILL_1__10135_ (
);

FILL FILL_0__7982_ (
);

FILL FILL_0__7562_ (
);

FILL FILL_0__7142_ (
);

FILL FILL_2__8941_ (
);

FILL FILL_2__8521_ (
);

FILL FILL_2__12767_ (
);

FILL FILL_2__12347_ (
);

FILL FILL_0__8767_ (
);

FILL FILL_3__6864_ (
);

FILL FILL_0__8347_ (
);

NOR2X1 _10618_ (
    .A(\u_fir_pe4.rYin [8]),
    .B(\u_fir_pe4.mul [8]),
    .Y(_3881_)
);

FILL FILL_1__12701_ (
);

FILL FILL_2__9726_ (
);

FILL FILL_2__9306_ (
);

FILL FILL_1__7723_ (
);

FILL FILL_1__7303_ (
);

FILL FILL_3__7649_ (
);

AOI21X1 _6793_ (
    .A(Xin[3]),
    .B(gnd),
    .C(_387_),
    .Y(_390_)
);

FILL FILL254550x234150 (
);

FILL FILL_3__10059_ (
);

FILL FILL_1__11093_ (
);

NAND3X1 _10791_ (
    .A(_4725_),
    .B(_3993_),
    .C(_3991_),
    .Y(_3994_)
);

OAI21X1 _10371_ (
    .A(_3626_),
    .B(_3628_),
    .C(_3619_),
    .Y(_3647_)
);

FILL FILL_0__10086_ (
);

FILL FILL_1__8928_ (
);

FILL FILL_1__8508_ (
);

FILL FILL_3__11420_ (
);

FILL FILL_2__10833_ (
);

FILL FILL_2__10413_ (
);

NOR2X1 _7998_ (
    .A(_1490_),
    .B(_1489_),
    .Y(_1502_)
);

AOI21X1 _7578_ (
    .A(_1078_),
    .B(_1080_),
    .C(_1095_),
    .Y(_1096_)
);

INVX1 _7158_ (
    .A(\u_fir_pe0.rYin [12]),
    .Y(_742_)
);

FILL FILL_0__6833_ (
);

FILL FILL_0__6413_ (
);

FILL FILL_1__12298_ (
);

NAND2X1 _11996_ (
    .A(_5109_),
    .B(_5113_),
    .Y(_5114_)
);

OAI21X1 _11576_ (
    .A(_4747_),
    .B(_4750_),
    .C(_4757_),
    .Y(_4760_)
);

OAI21X1 _11156_ (
    .A(_4120_),
    .B(_4353_),
    .C(_4267_),
    .Y(_4354_)
);

FILL FILL_3__12205_ (
);

FILL FILL_0__12652_ (
);

FILL FILL_0__12232_ (
);

FILL FILL_0__7618_ (
);

NOR2X1 _9724_ (
    .A(_3067_),
    .B(_3066_),
    .Y(_3068_)
);

OAI21X1 _9304_ (
    .A(_2649_),
    .B(_2653_),
    .C(_2656_),
    .Y(_2663_)
);

FILL FILL_1__8681_ (
);

FILL FILL_1__8261_ (
);

FILL FILL_0__13017_ (
);

NAND2X1 _13302_ (
    .A(_6325_),
    .B(_6320_),
    .Y(_6326_)
);

FILL FILL_1__9886_ (
);

FILL FILL_1__9466_ (
);

FILL FILL_1__9046_ (
);

FILL FILL_2__11791_ (
);

FILL FILL_2__11371_ (
);

FILL FILL_1__10784_ (
);

FILL FILL_1__10364_ (
);

FILL FILL_0__7791_ (
);

FILL FILL_2__7389_ (
);

FILL FILL_0__7371_ (
);

FILL FILL_2__8750_ (
);

FILL FILL_2__8330_ (
);

FILL FILL_3__13163_ (
);

NAND3X1 _6849_ (
    .A(_426_),
    .B(_430_),
    .C(_433_),
    .Y(_446_)
);

NAND2X1 _6429_ (
    .A(gnd),
    .B(Xin[1]),
    .Y(_31_)
);

FILL FILL_2__12996_ (
);

FILL FILL_2__12576_ (
);

FILL FILL_2__12156_ (
);

FILL FILL_0__13190_ (
);

FILL FILL_1__11989_ (
);

FILL FILL_1__11569_ (
);

FILL FILL_1__11149_ (
);

FILL FILL_0__8576_ (
);

FILL FILL_0__8156_ (
);

OAI21X1 _10847_ (
    .A(_4048_),
    .B(_4047_),
    .C(_4014_),
    .Y(_4049_)
);

AOI21X1 _10427_ (
    .A(_3648_),
    .B(_3682_),
    .C(_3701_),
    .Y(_3702_)
);

OAI21X1 _10007_ (
    .A(_3286_),
    .B(_3287_),
    .C(_3285_),
    .Y(_3288_)
);

FILL FILL_1__12930_ (
);

FILL FILL_2__9955_ (
);

FILL FILL_2__9535_ (
);

FILL FILL_0__11923_ (
);

FILL FILL_2__9115_ (
);

FILL FILL_0__11503_ (
);

FILL FILL_1__7952_ (
);

FILL FILL_1__7532_ (
);

FILL FILL_1__7112_ (
);

FILL FILL_0__12708_ (
);

FILL FILL_3__10288_ (
);

NAND3X1 _10180_ (
    .A(_3412_),
    .B(_3454_),
    .C(_3455_),
    .Y(_3459_)
);

FILL FILL_1__8737_ (
);

FILL FILL_1__8317_ (
);

FILL FILL_2__10642_ (
);

FILL FILL_2__10222_ (
);

NAND3X1 _7387_ (
    .A(_823_),
    .B(_903_),
    .C(_907_),
    .Y(_908_)
);

FILL FILL_3__9604_ (
);

FILL FILL_0__6642_ (
);

OAI21X1 _11385_ (
    .A(_4290_),
    .B(_4577_),
    .C(_4556_),
    .Y(_4578_)
);

FILL FILL_2__7601_ (
);

FILL FILL_3__12434_ (
);

FILL FILL_2__11847_ (
);

FILL FILL_0__12881_ (
);

FILL FILL_2__11427_ (
);

FILL FILL_2__11007_ (
);

FILL FILL_0__12041_ (
);

FILL FILL_0__7847_ (
);

NAND2X1 _9953_ (
    .A(_3232_),
    .B(_3228_),
    .Y(_3235_)
);

FILL FILL_0__7427_ (
);

AOI21X1 _9533_ (
    .A(_2786_),
    .B(_2816_),
    .C(_2819_),
    .Y(_2889_)
);

FILL FILL_0__7007_ (
);

NAND2X1 _9113_ (
    .A(gnd),
    .B(\X[3] [2]),
    .Y(_2474_)
);

FILL FILL_1__8490_ (
);

FILL FILL_1__8070_ (
);

FILL FILL_2__8806_ (
);

FILL FILL_0__13246_ (
);

NOR2X1 _13111_ (
    .A(_6052_),
    .B(_6105_),
    .Y(_6145_)
);

FILL FILL_1__6803_ (
);

FILL FILL_3__6729_ (
);

FILL FILL_1__9695_ (
);

FILL FILL_1__9275_ (
);

FILL FILL_2__11180_ (
);

FILL FILL_1__10593_ (
);

FILL FILL_1__10173_ (
);

FILL FILL_0__7180_ (
);

FILL FILL_2_BUFX2_insert10 (
);

FILL FILL_2__7198_ (
);

FILL FILL_2_BUFX2_insert11 (
);

FILL FILL_3__10920_ (
);

FILL FILL_3__10500_ (
);

NAND3X1 _6658_ (
    .A(_253_),
    .B(_252_),
    .C(_256_),
    .Y(_257_)
);

FILL FILL_2__12385_ (
);

FILL FILL_1__11798_ (
);

FILL FILL_1__11378_ (
);

FILL FILL_0__8385_ (
);

FILL FILL_3__6482_ (
);

OAI21X1 _10656_ (
    .A(_3912_),
    .B(_3913_),
    .C(_3917_),
    .Y(_3920_)
);

NAND3X1 _10236_ (
    .A(gnd),
    .B(\X[4] [6]),
    .C(_3513_),
    .Y(_3514_)
);

FILL FILL_3__11705_ (
);

FILL FILL_2__9764_ (
);

FILL FILL_2__9344_ (
);

FILL FILL_0__11732_ (
);

FILL FILL_0__11312_ (
);

NOR2X1 _8804_ (
    .A(_2225_),
    .B(_2230_),
    .Y(_2233_)
);

FILL FILL_1__7761_ (
);

FILL FILL_1__7341_ (
);

FILL FILL_3__7687_ (
);

FILL FILL_3__7267_ (
);

FILL FILL_1__13104_ (
);

FILL FILL_0__12937_ (
);

AOI21X1 _12802_ (
    .A(_5840_),
    .B(_5839_),
    .C(_5838_),
    .Y(_5841_)
);

FILL FILL_0__12517_ (
);

FILL FILL_1__8546_ (
);

FILL FILL_2__10871_ (
);

FILL FILL_2__10451_ (
);

FILL FILL_2__10031_ (
);

NOR2X1 _7196_ (
    .A(_777_),
    .B(_720_),
    .Y(_792_[1])
);

FILL FILL_2__6889_ (
);

FILL FILL_0__6871_ (
);

FILL FILL_2__6469_ (
);

FILL FILL_0__6451_ (
);

AOI21X1 _11194_ (
    .A(_4316_),
    .B(_4390_),
    .C(_4389_),
    .Y(_4391_)
);

FILL FILL_2__7830_ (
);

FILL FILL_3__12663_ (
);

FILL FILL_2__7410_ (
);

FILL FILL_2__11656_ (
);

FILL FILL_0__12690_ (
);

FILL FILL_2__11236_ (
);

FILL FILL_0__12270_ (
);

FILL FILL_1__10649_ (
);

FILL FILL_1__10229_ (
);

FILL FILL_0__7656_ (
);

INVX1 _9762_ (
    .A(_3105_),
    .Y(_3106_)
);

AND2X2 _9342_ (
    .A(_2698_),
    .B(_2697_),
    .Y(_2700_)
);

INVX1 _12399_ (
    .A(_5501_),
    .Y(_5503_)
);

FILL FILL_2__8615_ (
);

FILL FILL_3__13028_ (
);

FILL FILL_0__13055_ (
);

DFFPOSX1 _13340_ (
    .D(_6369_[2]),
    .CLK(clk_bF$buf27),
    .Q(\Y[7] [2])
);

FILL FILL_1__6612_ (
);

FILL FILL_3__6958_ (
);

FILL FILL_1__9084_ (
);

FILL FILL_0__9802_ (
);

FILL FILL_1__7817_ (
);

AND2X2 _6887_ (
    .A(_476_),
    .B(_482_),
    .Y(_483_)
);

NOR3X1 _6467_ (
    .A(_53_),
    .B(_20_),
    .C(_65_),
    .Y(_68_)
);

FILL FILL_2__12194_ (
);

FILL FILL_1__11187_ (
);

FILL FILL_0__8194_ (
);

NAND3X1 _10885_ (
    .A(_4081_),
    .B(_4067_),
    .C(_4085_),
    .Y(_4086_)
);

NAND2X1 _10465_ (
    .A(_3736_),
    .B(_3739_),
    .Y(_3740_)
);

AOI21X1 _10045_ (
    .A(_3279_),
    .B(_3283_),
    .C(_3272_),
    .Y(_3325_)
);

FILL FILL_3__11934_ (
);

FILL FILL_3__11514_ (
);

FILL FILL_2__10927_ (
);

FILL FILL_2__9993_ (
);

FILL FILL_2__9573_ (
);

FILL FILL_0__11961_ (
);

FILL FILL_2__10507_ (
);

FILL FILL_2__9153_ (
);

FILL FILL_0__11541_ (
);

FILL FILL_0__11121_ (
);

FILL FILL_2__13399_ (
);

FILL FILL_0__6927_ (
);

FILL FILL_0__6507_ (
);

NAND2X1 _8613_ (
    .A(_2048_),
    .B(_1891_),
    .Y(_2049_)
);

FILL FILL_1__7990_ (
);

FILL FILL_1__7570_ (
);

FILL FILL_1__7150_ (
);

FILL FILL_0__9399_ (
);

FILL FILL_3__7076_ (
);

FILL FILL_1__13333_ (
);

FILL FILL_0__12746_ (
);

NAND2X1 _12611_ (
    .A(_6279_),
    .B(_5651_),
    .Y(_5652_)
);

FILL FILL_0__12326_ (
);

OR2X2 _9818_ (
    .A(\u_fir_pe3.rYin [15]),
    .B(\u_fir_pe3.mul [15]),
    .Y(_3162_)
);

FILL FILL_1__8775_ (
);

FILL FILL_1__8355_ (
);

FILL FILL_2__10680_ (
);

FILL FILL_2__10260_ (
);

FILL FILL_3__9222_ (
);

FILL FILL_2__6698_ (
);

FILL FILL_0__6680_ (
);

FILL FILL_3__12892_ (
);

FILL FILL_3__12052_ (
);

FILL FILL_2__11885_ (
);

FILL FILL_2__11465_ (
);

FILL FILL_2__11045_ (
);

FILL FILL_1__10878_ (
);

FILL FILL_1__10458_ (
);

FILL FILL_1__10038_ (
);

FILL FILL_0__7885_ (
);

OAI22X1 _9991_ (
    .A(_3919_),
    .B(_3271_),
    .C(_3221_),
    .D(_3226_),
    .Y(_3272_)
);

FILL FILL_0__7465_ (
);

NAND3X1 _9571_ (
    .A(_2920_),
    .B(_2925_),
    .C(_2924_),
    .Y(_2926_)
);

FILL FILL_0__7045_ (
);

INVX1 _9151_ (
    .A(_2411_),
    .Y(_2512_)
);

FILL FILL_2__8844_ (
);

FILL FILL_2__8424_ (
);

FILL FILL_0__10812_ (
);

FILL FILL_3__13257_ (
);

FILL FILL_2__8004_ (
);

FILL FILL_0__13284_ (
);

FILL FILL_1__6841_ (
);

FILL FILL_1__6421_ (
);

FILL FILL_1__12604_ (
);

FILL FILL_2__9629_ (
);

FILL FILL_0__9611_ (
);

FILL FILL_2__9209_ (
);

FILL FILL_1__7626_ (
);

AND2X2 _6696_ (
    .A(_294_),
    .B(_290_),
    .Y(_796_[7])
);

FILL FILL_3__8913_ (
);

NAND2X1 _10694_ (
    .A(\u_fir_pe4.rYin [15]),
    .B(\u_fir_pe4.mul [15]),
    .Y(_3957_)
);

NAND3X1 _10274_ (
    .A(_3491_),
    .B(_3548_),
    .C(_3549_),
    .Y(_3552_)
);

FILL FILL_2__6910_ (
);

FILL FILL_3__11743_ (
);

FILL FILL_2__9382_ (
);

FILL FILL_0__11770_ (
);

FILL FILL_2__10316_ (
);

FILL FILL_0__11350_ (
);

FILL FILL_0__6736_ (
);

OAI21X1 _8842_ (
    .A(_2259_),
    .B(_2260_),
    .C(_2264_),
    .Y(_2266_)
);

NAND3X1 _8422_ (
    .A(_1832_),
    .B(_1851_),
    .C(_1845_),
    .Y(_1861_)
);

INVX1 _8002_ (
    .A(_1489_),
    .Y(_1505_)
);

OAI21X1 _11899_ (
    .A(_5560_),
    .B(_5017_),
    .C(_5009_),
    .Y(_5018_)
);

NAND2X1 _11479_ (
    .A(_4662_),
    .B(_4657_),
    .Y(_4663_)
);

AOI21X1 _11059_ (
    .A(_4257_),
    .B(_4256_),
    .C(_4255_),
    .Y(_4258_)
);

FILL FILL_3__12528_ (
);

FILL FILL_1__13142_ (
);

FILL FILL_0__12975_ (
);

AOI21X1 _12840_ (
    .A(_5860_),
    .B(_5862_),
    .C(_5877_),
    .Y(_5878_)
);

FILL FILL_0__12555_ (
);

FILL FILL_0__12135_ (
);

INVX1 _12420_ (
    .A(\u_fir_pe6.rYin [12]),
    .Y(_5524_)
);

OAI21X1 _12000_ (
    .A(_5117_),
    .B(_5111_),
    .C(_5105_),
    .Y(_5118_)
);

NOR2X1 _9627_ (
    .A(_2980_),
    .B(_2979_),
    .Y(_2981_)
);

NAND3X1 _9207_ (
    .A(_2564_),
    .B(_2566_),
    .C(_2565_),
    .Y(_2567_)
);

FILL FILL_1__8584_ (
);

FILL FILL_1__8164_ (
);

FILL FILL_3__9451_ (
);

NAND2X1 _13205_ (
    .A(_6231_),
    .B(_6226_),
    .Y(_6232_)
);

FILL FILL_1__9789_ (
);

FILL FILL_1__9369_ (
);

FILL FILL_2__11694_ (
);

FILL FILL_2__11274_ (
);

FILL FILL_1__10687_ (
);

FILL FILL_1__10267_ (
);

FILL FILL_0__7694_ (
);

FILL FILL_0__7274_ (
);

INVX1 _9380_ (
    .A(_2651_),
    .Y(_2738_)
);

FILL FILL_2__8653_ (
);

FILL FILL_2__8233_ (
);

FILL FILL_0__10621_ (
);

FILL FILL_0__10201_ (
);

FILL FILL_2__12899_ (
);

FILL FILL_2__12059_ (
);

FILL FILL_0__13093_ (
);

FILL FILL_1__6650_ (
);

FILL FILL_0__8899_ (
);

FILL FILL_2__13000_ (
);

FILL FILL_0__8479_ (
);

FILL FILL_3__6576_ (
);

FILL FILL_0__8059_ (
);

FILL FILL_1__12833_ (
);

FILL FILL_1__12413_ (
);

FILL FILL_0__9420_ (
);

FILL FILL_2__9438_ (
);

FILL FILL_0__11826_ (
);

FILL FILL_2__9018_ (
);

FILL FILL_0__11406_ (
);

FILL FILL_1__7855_ (
);

FILL FILL_1__7435_ (
);

FILL FILL_1__7015_ (
);

FILL FILL_3__8302_ (
);

NAND3X1 _10083_ (
    .A(_3350_),
    .B(_3354_),
    .C(_3356_),
    .Y(_3363_)
);

FILL FILL_3__11972_ (
);

FILL FILL_3__11132_ (
);

FILL FILL_2__10965_ (
);

FILL FILL_2__10545_ (
);

FILL FILL_2__9191_ (
);

FILL FILL_2__10125_ (
);

FILL FILL_0__6965_ (
);

FILL FILL_0__6545_ (
);

NAND2X1 _8651_ (
    .A(_2085_),
    .B(_2081_),
    .Y(_2087_)
);

NAND3X1 _8231_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf1 ),
    .C(_1669_),
    .Y(_1672_)
);

AND2X2 _11288_ (
    .A(_4472_),
    .B(_4476_),
    .Y(_4484_)
);

FILL FILL_2__7924_ (
);

FILL FILL_3__12757_ (
);

FILL FILL_2__7504_ (
);

FILL FILL_0__12784_ (
);

FILL FILL_0__12364_ (
);

DFFPOSX1 _9856_ (
    .D(\Y[3] [2]),
    .CLK(clk_bF$buf36),
    .Q(\u_fir_pe3.rYin [2])
);

AOI22X1 _9436_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf0 ),
    .C(gnd),
    .D(\X[3] [6]),
    .Y(_2793_)
);

NOR2X1 _9016_ (
    .A(_3141_),
    .B(_3131_),
    .Y(_3151_)
);

FILL FILL_1__8393_ (
);

FILL FILL_2__8709_ (
);

FILL FILL_3__9680_ (
);

FILL FILL_0__13149_ (
);

NOR2X1 _13014_ (
    .A(_5985_),
    .B(_5982_),
    .Y(_6050_)
);

FILL FILL_1__6706_ (
);

FILL FILL_1__9598_ (
);

FILL FILL_1__9178_ (
);

FILL FILL_3__12090_ (
);

FILL FILL_2__11083_ (
);

FILL FILL_1__10496_ (
);

FILL FILL_1__10076_ (
);

FILL FILL_0__7083_ (
);

FILL FILL_3__10403_ (
);

FILL FILL_2__8882_ (
);

FILL FILL_2__8462_ (
);

FILL FILL_0__10850_ (
);

FILL FILL_0__10430_ (
);

FILL FILL_2__8042_ (
);

FILL FILL_0__10010_ (
);

FILL FILL_2__12288_ (
);

NOR2X1 _7922_ (
    .A(_1429_),
    .B(_1430_),
    .Y(_1431_)
);

OAI21X1 _7502_ (
    .A(_970_),
    .B(_1020_),
    .C(_964_),
    .Y(_1021_)
);

FILL FILL_0__8288_ (
);

OAI21X1 _10979_ (
    .A(_4178_),
    .B(_4173_),
    .C(_4101_),
    .Y(_4179_)
);

NOR2X1 _10559_ (
    .A(_3827_),
    .B(_3826_),
    .Y(_3978_[1])
);

AOI22X1 _10139_ (
    .A(gnd),
    .B(\X[4] [7]),
    .C(\X[4] [3]),
    .D(gnd),
    .Y(_3418_)
);

FILL FILL_1__12642_ (
);

FILL FILL_1__12222_ (
);

FILL FILL_2__9667_ (
);

FILL FILL_2__9247_ (
);

NAND3X1 _11920_ (
    .A(_5035_),
    .B(_5034_),
    .C(_5038_),
    .Y(_5039_)
);

AND2X2 _11500_ (
    .A(_4662_),
    .B(_4672_),
    .Y(_4683_)
);

FILL FILL_0__11215_ (
);

NAND2X1 _8707_ (
    .A(_2141_),
    .B(_2108_),
    .Y(_2142_)
);

FILL FILL_1__7664_ (
);

FILL FILL_1__13007_ (
);

FILL FILL_3__8531_ (
);

NAND3X1 _12705_ (
    .A(_5735_),
    .B(_5742_),
    .C(_5744_),
    .Y(_5745_)
);

FILL FILL_1__8869_ (
);

FILL FILL_1__8449_ (
);

FILL FILL_1__8029_ (
);

FILL FILL_3__11361_ (
);

FILL FILL_2__10774_ (
);

FILL FILL_2__10354_ (
);

FILL FILL_1__9810_ (
);

INVX1 _7099_ (
    .A(\u_fir_pe0.mul [7]),
    .Y(_682_)
);

FILL FILL_3__9316_ (
);

FILL FILL_0__6774_ (
);

INVX1 _8880_ (
    .A(_2299_),
    .Y(_2303_)
);

NAND2X1 _8460_ (
    .A(\X[2] [1]),
    .B(gnd),
    .Y(_1898_)
);

NAND2X1 _8040_ (
    .A(_1543_),
    .B(_1538_),
    .Y(_1544_)
);

OAI21X1 _11097_ (
    .A(_4293_),
    .B(_4294_),
    .C(_4289_),
    .Y(_4295_)
);

FILL FILL_3__12986_ (
);

FILL FILL_2__7733_ (
);

FILL FILL_2__7313_ (
);

FILL FILL_3__12146_ (
);

FILL FILL_1__13180_ (
);

FILL FILL_2__11979_ (
);

FILL FILL_2__11559_ (
);

FILL FILL_0__12593_ (
);

FILL FILL_2__11139_ (
);

FILL FILL_0__12173_ (
);

FILL FILL_2__12920_ (
);

FILL FILL_0__7979_ (
);

FILL FILL_0__7559_ (
);

INVX1 _9665_ (
    .A(_3007_),
    .Y(_3017_)
);

FILL FILL_0__7139_ (
);

INVX1 _9245_ (
    .A(_2603_),
    .Y(_2604_)
);

FILL FILL_1__11913_ (
);

FILL FILL_2__8938_ (
);

FILL FILL_0__8920_ (
);

FILL FILL_0__8500_ (
);

FILL FILL_2__8518_ (
);

FILL FILL_0__10906_ (
);

NOR2X1 _13243_ (
    .A(_6263_),
    .B(_6262_),
    .Y(_6266_)
);

FILL FILL_1__6935_ (
);

FILL FILL_1__6515_ (
);

FILL FILL_0__9705_ (
);

FILL FILL_3__7802_ (
);

FILL FILL_2__8691_ (
);

FILL FILL_2__8271_ (
);

FILL FILL_2__12097_ (
);

OR2X2 _7731_ (
    .A(_1177_),
    .B(_1247_),
    .Y(_1248_)
);

AND2X2 _7311_ (
    .A(vdd),
    .B(\X[1] [2]),
    .Y(_833_)
);

NAND3X1 _10788_ (
    .A(_3986_),
    .B(_3990_),
    .C(_3988_),
    .Y(_3991_)
);

AOI21X1 _10368_ (
    .A(_3629_),
    .B(_3625_),
    .C(_3570_),
    .Y(_3644_)
);

FILL FILL_1__12871_ (
);

FILL FILL_1__12451_ (
);

FILL FILL_1__12031_ (
);

FILL FILL_2__9896_ (
);

FILL FILL_2__9476_ (
);

FILL FILL_0__11864_ (
);

FILL FILL_2__9056_ (
);

FILL FILL_0__11444_ (
);

FILL FILL_0__11024_ (
);

NOR2X1 _8936_ (
    .A(_2358_),
    .B(_2352_),
    .Y(_2360_)
);

NAND3X1 _8516_ (
    .A(_1947_),
    .B(_1948_),
    .C(_1949_),
    .Y(_1954_)
);

FILL FILL_1__7893_ (
);

FILL FILL_1__7473_ (
);

FILL FILL_1__7053_ (
);

FILL FILL_3__7399_ (
);

FILL FILL_3_BUFX2_insert80 (
);

FILL FILL_1__13236_ (
);

FILL FILL_3_BUFX2_insert82 (
);

FILL FILL_3_BUFX2_insert84 (
);

FILL FILL_3_BUFX2_insert85 (
);

FILL FILL_3_BUFX2_insert87 (
);

FILL FILL_3__8760_ (
);

INVX1 _12934_ (
    .A(_5965_),
    .Y(_5971_)
);

FILL FILL_0__12649_ (
);

FILL FILL_3_BUFX2_insert89 (
);

FILL FILL_0__12229_ (
);

DFFPOSX1 _12514_ (
    .D(_5578_[13]),
    .CLK(clk_bF$buf37),
    .Q(\u_fir_pe6.mul [13])
);

FILL FILL_1__8678_ (
);

FILL FILL_1__8258_ (
);

FILL FILL_2__10583_ (
);

FILL FILL_2__10163_ (
);

FILL FILL_3__9545_ (
);

FILL FILL_0__6583_ (
);

FILL FILL_2__7962_ (
);

FILL FILL_2__7542_ (
);

FILL FILL_3__12375_ (
);

FILL FILL_2__7122_ (
);

FILL FILL_2__11788_ (
);

FILL FILL_2__11368_ (
);

FILL FILL_0__7788_ (
);

INVX1 _9894_ (
    .A(\X[4] [2]),
    .Y(_3958_)
);

FILL FILL_0__7368_ (
);

AOI21X1 _9474_ (
    .A(_2821_),
    .B(_2817_),
    .C(_2776_),
    .Y(_2831_)
);

NAND2X1 _9054_ (
    .A(\X[3] [4]),
    .B(gnd),
    .Y(_2416_)
);

FILL FILL_1__11722_ (
);

FILL FILL_1__11302_ (
);

FILL FILL_2__8747_ (
);

FILL FILL_2__8327_ (
);

FILL FILL_0__13187_ (
);

OAI21X1 _13052_ (
    .A(_6087_),
    .B(_5955_),
    .C(_6037_),
    .Y(_6088_)
);

FILL FILL_1__6744_ (
);

FILL FILL_1__12927_ (
);

FILL FILL_0__9934_ (
);

FILL FILL_0__9514_ (
);

FILL FILL_1__7949_ (
);

FILL FILL_3__10861_ (
);

FILL FILL_1__7529_ (
);

FILL FILL_3__10441_ (
);

FILL FILL_1__7109_ (
);

FILL FILL_3__10021_ (
);

AOI21X1 _6599_ (
    .A(_186_),
    .B(_185_),
    .C(_136_),
    .Y(_199_)
);

NOR2X1 _7960_ (
    .A(\u_fir_pe1.rYin [5]),
    .B(\u_fir_pe1.mul [5]),
    .Y(_1465_)
);

AOI21X1 _7540_ (
    .A(_1058_),
    .B(_1057_),
    .C(_1056_),
    .Y(_1059_)
);

OAI21X1 _7120_ (
    .A(_692_),
    .B(_693_),
    .C(_703_),
    .Y(_704_)
);

INVX1 _10597_ (
    .A(\u_fir_pe4.rYin [6]),
    .Y(_3861_)
);

NAND3X1 _10177_ (
    .A(_3454_),
    .B(_3455_),
    .C(_3453_),
    .Y(_3456_)
);

FILL FILL_2__6813_ (
);

FILL FILL_3__11646_ (
);

FILL FILL_1__12680_ (
);

FILL FILL_3__11226_ (
);

FILL FILL_1__12260_ (
);

FILL FILL_2__10639_ (
);

FILL FILL_2__9285_ (
);

FILL FILL_0__11673_ (
);

FILL FILL_2__10219_ (
);

FILL FILL_0__11253_ (
);

FILL FILL_0__6639_ (
);

NAND2X1 _8745_ (
    .A(_2176_),
    .B(_2178_),
    .Y(_2179_)
);

OAI21X1 _8325_ (
    .A(_1763_),
    .B(_1764_),
    .C(_1762_),
    .Y(_1765_)
);

FILL FILL_1__7282_ (
);

FILL FILL_1__13045_ (
);

FILL FILL_0__12878_ (
);

AOI21X1 _12743_ (
    .A(_5699_),
    .B(_5705_),
    .C(_5782_),
    .Y(_5783_)
);

FILL FILL_0__12458_ (
);

FILL FILL_0__12038_ (
);

INVX1 _12323_ (
    .A(\u_fir_pe6.rYin [3]),
    .Y(_5430_)
);

FILL FILL_1__8487_ (
);

FILL FILL_1__8067_ (
);

FILL FILL_2__10392_ (
);

FILL FILL_3__9774_ (
);

INVX1 _13108_ (
    .A(_6141_),
    .Y(_6142_)
);

FILL FILL_0__6392_ (
);

FILL FILL_2__7771_ (
);

FILL FILL_2__7351_ (
);

FILL FILL_2__11177_ (
);

AND2X2 _6811_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_408_)
);

FILL FILL_0__7597_ (
);

FILL FILL_0__7177_ (
);

OAI21X1 _9283_ (
    .A(_2641_),
    .B(_2636_),
    .C(_2630_),
    .Y(_2642_)
);

FILL FILL_1__11951_ (
);

FILL FILL_1__11531_ (
);

FILL FILL_1__11111_ (
);

FILL FILL_2__8556_ (
);

FILL FILL_0__10944_ (
);

FILL FILL_2__8136_ (
);

FILL FILL_0__10524_ (
);

FILL FILL_0__10104_ (
);

NOR2X1 _13281_ (
    .A(_6303_),
    .B(_6304_),
    .Y(_6305_)
);

FILL FILL_1__6973_ (
);

FILL FILL_1__6553_ (
);

FILL FILL_2__13323_ (
);

FILL FILL_3__6899_ (
);

FILL FILL_1__12736_ (
);

FILL FILL_1__12316_ (
);

FILL FILL_0__9743_ (
);

FILL FILL_3__7840_ (
);

FILL FILL_0__9323_ (
);

FILL FILL_0__11729_ (
);

FILL FILL_3__7420_ (
);

FILL FILL_3__7000_ (
);

FILL FILL_0__11309_ (
);

FILL FILL_1__7758_ (
);

FILL FILL_3__10670_ (
);

FILL FILL_1__7338_ (
);

FILL FILL_3__8625_ (
);

FILL FILL_3__8205_ (
);

FILL FILL_3__11875_ (
);

FILL FILL_2__6622_ (
);

FILL FILL_3__11455_ (
);

FILL FILL_2__10868_ (
);

FILL FILL_2__10448_ (
);

FILL FILL_2__9094_ (
);

FILL FILL_0__11482_ (
);

FILL FILL_2__10028_ (
);

FILL FILL_0__11062_ (
);

FILL FILL_1__9904_ (
);

FILL FILL_0__6868_ (
);

DFFPOSX1 _8974_ (
    .D(\X[2]_5_bF$buf1 ),
    .CLK(clk_bF$buf14),
    .Q(\X[3] [5])
);

FILL FILL_0__6448_ (
);

OAI21X1 _8554_ (
    .A(_1916_),
    .B(_1990_),
    .C(_1937_),
    .Y(_1991_)
);

INVX1 _8134_ (
    .A(_2294_),
    .Y(_2304_)
);

FILL FILL_1__7091_ (
);

FILL FILL_1__10802_ (
);

FILL FILL_2__7827_ (
);

FILL FILL_2__7407_ (
);

FILL FILL_1__13274_ (
);

OAI21X1 _12972_ (
    .A(_6008_),
    .B(_6007_),
    .C(_6006_),
    .Y(_6009_)
);

FILL FILL_0__12687_ (
);

FILL FILL_0__12267_ (
);

NAND2X1 _12552_ (
    .A(_5592_),
    .B(_5588_),
    .Y(_5595_)
);

OAI22X1 _12132_ (
    .A(_4797_),
    .B(_5244_),
    .C(_5245_),
    .D(_5247_),
    .Y(_5248_)
);

AND2X2 _9759_ (
    .A(\u_fir_pe3.rYin [9]),
    .B(\u_fir_pe3.mul [9]),
    .Y(_3103_)
);

NOR2X1 _9339_ (
    .A(_3161_),
    .B(_2696_),
    .Y(_2697_)
);

FILL FILL_1__8296_ (
);

FILL FILL_3__9163_ (
);

NOR2X1 _13337_ (
    .A(_6358_),
    .B(_6365_),
    .Y(_6372_[2])
);

FILL FILL_1__6609_ (
);

FILL FILL_2__7580_ (
);

FILL FILL_2__7160_ (
);

AOI21X1 _6620_ (
    .A(_147_),
    .B(_143_),
    .C(_212_),
    .Y(_219_)
);

FILL FILL_1__10399_ (
);

AOI21X1 _9092_ (
    .A(_2431_),
    .B(_2435_),
    .C(_2423_),
    .Y(_2454_)
);

FILL FILL_1__11760_ (
);

FILL FILL_1__11340_ (
);

FILL FILL_2__8785_ (
);

FILL FILL_2__8365_ (
);

FILL FILL_3__13198_ (
);

FILL FILL_0__10333_ (
);

NAND3X1 _13090_ (
    .A(_6122_),
    .B(_6124_),
    .C(_6123_),
    .Y(_6125_)
);

INVX1 _7825_ (
    .A(_1312_),
    .Y(_1340_)
);

INVX1 _7405_ (
    .A(_922_),
    .Y(_926_)
);

FILL FILL_1__6782_ (
);

FILL FILL_2__13132_ (
);

FILL FILL_1__12965_ (
);

FILL FILL_1__12545_ (
);

FILL FILL_1__12125_ (
);

FILL FILL_0__9972_ (
);

FILL FILL_0__9552_ (
);

FILL FILL_0__11958_ (
);

FILL FILL_0__9132_ (
);

INVX1 _11823_ (
    .A(_4942_),
    .Y(_4943_)
);

FILL FILL_0__11538_ (
);

NAND2X1 _11403_ (
    .A(_4574_),
    .B(_4573_),
    .Y(_4596_)
);

FILL FILL_0__11118_ (
);

FILL FILL253950x21750 (
);

FILL FILL_1__7987_ (
);

FILL FILL_1__7567_ (
);

FILL FILL_1__7147_ (
);

FILL FILL_3__8854_ (
);

NAND2X1 _12608_ (
    .A(\X[6] [0]),
    .B(gnd),
    .Y(_5649_)
);

FILL FILL_3__8014_ (
);

FILL FILL_2__6851_ (
);

FILL FILL_3__11684_ (
);

FILL FILL_2__6431_ (
);

FILL FILL_2__10677_ (
);

FILL FILL_2__10257_ (
);

FILL FILL_0__11291_ (
);

FILL FILL_1__9713_ (
);

FILL FILL_3__9639_ (
);

FILL FILL_0__6677_ (
);

NAND2X1 _8783_ (
    .A(_2214_),
    .B(_2213_),
    .Y(_2215_)
);

AOI21X1 _8363_ (
    .A(_1766_),
    .B(_1770_),
    .C(_1732_),
    .Y(_1802_)
);

FILL FILL_1__10611_ (
);

FILL FILL_2__7636_ (
);

FILL FILL_1__13083_ (
);

NAND2X1 _12781_ (
    .A(vdd),
    .B(\X[6] [4]),
    .Y(_5820_)
);

FILL FILL_0__12076_ (
);

INVX1 _12361_ (
    .A(\u_fir_pe6.mul [7]),
    .Y(_5464_)
);

FILL FILL_2__12823_ (
);

FILL FILL_2__12403_ (
);

NAND3X1 _9988_ (
    .A(_3258_),
    .B(_3266_),
    .C(_3268_),
    .Y(_3269_)
);

OAI21X1 _9568_ (
    .A(_2922_),
    .B(_2921_),
    .C(_2915_),
    .Y(_2923_)
);

NAND3X1 _9148_ (
    .A(_2417_),
    .B(_2504_),
    .C(_2505_),
    .Y(_2509_)
);

FILL FILL_1__11816_ (
);

FILL FILL_0__8823_ (
);

FILL FILL_0__8403_ (
);

FILL FILL_0__10809_ (
);

FILL FILL_3__6500_ (
);

FILL FILL_3__9392_ (
);

OR2X2 _13146_ (
    .A(_6151_),
    .B(_6177_),
    .Y(_6179_)
);

FILL FILL_1__6838_ (
);

FILL FILL_1__6418_ (
);

FILL FILL_0__9608_ (
);

FILL FILL_3__10955_ (
);

FILL FILL_3__10535_ (
);

FILL FILL_3__10115_ (
);

FILL FILL_2__8594_ (
);

FILL FILL_0__10982_ (
);

FILL FILL_2__8174_ (
);

FILL FILL_0__10562_ (
);

FILL FILL_0__10142_ (
);

OAI21X1 _7634_ (
    .A(_1138_),
    .B(_1142_),
    .C(_1145_),
    .Y(_1152_)
);

DFFPOSX1 _7214_ (
    .D(_790_[15]),
    .CLK(clk_bF$buf25),
    .Q(\Y[1] [15])
);

FILL FILL_1__6591_ (
);

FILL FILL_2__6907_ (
);

FILL FILL_1__12774_ (
);

FILL FILL_1__12354_ (
);

FILL FILL_0__9781_ (
);

FILL FILL_2__9799_ (
);

FILL FILL253650x248550 (
);

FILL FILL_2__9379_ (
);

FILL FILL_0__9361_ (
);

FILL FILL_0__11767_ (
);

DFFPOSX1 _11632_ (
    .D(_4781_[8]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [8])
);

FILL FILL_0__11347_ (
);

NAND2X1 _11212_ (
    .A(_4400_),
    .B(_4407_),
    .Y(_4409_)
);

NAND2X1 _8839_ (
    .A(_2263_),
    .B(_2258_),
    .Y(_2264_)
);

INVX1 _8419_ (
    .A(_1761_),
    .Y(_1858_)
);

FILL FILL_1__7796_ (
);

FILL FILL_1__7376_ (
);

FILL FILL_1__13139_ (
);

AOI21X1 _12837_ (
    .A(_5786_),
    .B(_5864_),
    .C(_5872_),
    .Y(_5875_)
);

FILL FILL_3__8243_ (
);

AOI21X1 _12417_ (
    .A(_5517_),
    .B(_5508_),
    .C(_5515_),
    .Y(_5520_)
);

FILL FILL_2__6660_ (
);

FILL FILL_3__11073_ (
);

FILL FILL_2__10486_ (
);

FILL FILL_2__10066_ (
);

FILL FILL_1__9942_ (
);

FILL FILL_1__9522_ (
);

FILL FILL_1__9102_ (
);

FILL FILL_3__9028_ (
);

FILL FILL_0__6486_ (
);

AOI21X1 _8592_ (
    .A(_2019_),
    .B(_2017_),
    .C(_1989_),
    .Y(_2029_)
);

NAND3X1 _8172_ (
    .A(_1614_),
    .B(_2380_),
    .C(_1613_),
    .Y(_1615_)
);

FILL FILL_1__10840_ (
);

FILL FILL_1__10420_ (
);

FILL FILL_1__10000_ (
);

FILL FILL_2__7865_ (
);

FILL FILL_3__12698_ (
);

FILL FILL_2__7445_ (
);

FILL FILL_2__7025_ (
);

AOI22X1 _12590_ (
    .A(_5588_),
    .B(_5593_),
    .C(_5628_),
    .D(_5631_),
    .Y(_5632_)
);

AOI21X1 _12170_ (
    .A(_5213_),
    .B(_5219_),
    .C(_5285_),
    .Y(_5286_)
);

NAND3X1 _6905_ (
    .A(_496_),
    .B(_497_),
    .C(_500_),
    .Y(_501_)
);

FILL FILL_2__12632_ (
);

FILL FILL_2__12212_ (
);

OAI21X1 _9797_ (
    .A(_3133_),
    .B(_3134_),
    .C(_3138_),
    .Y(_3140_)
);

OAI21X1 _9377_ (
    .A(_2726_),
    .B(_2720_),
    .C(_2728_),
    .Y(_2735_)
);

FILL FILL_1__11205_ (
);

FILL FILL_0__8632_ (
);

FILL FILL_0__8212_ (
);

FILL FILL_0__10618_ (
);

NAND3X1 _10903_ (
    .A(_4039_),
    .B(_4102_),
    .C(_4103_),
    .Y(_4104_)
);

DFFPOSX1 _13375_ (
    .D(\Y[6] [13]),
    .CLK(clk_bF$buf40),
    .Q(\u_fir_pe7.rYin [13])
);

FILL FILL_1__6647_ (
);

FILL FILL_2__13417_ (
);

FILL FILL_0__9417_ (
);

FILL FILL_3__7514_ (
);

FILL FILL_3__10344_ (
);

FILL FILL_0__10791_ (
);

FILL FILL_0__10371_ (
);

FILL FILL_3__8719_ (
);

NAND3X1 _7863_ (
    .A(_1358_),
    .B(_1375_),
    .C(_1374_),
    .Y(_1377_)
);

NAND3X1 _7443_ (
    .A(_953_),
    .B(_960_),
    .C(_962_),
    .Y(_963_)
);

AOI21X1 _7023_ (
    .A(_557_),
    .B(_559_),
    .C(_614_),
    .Y(_615_)
);

FILL FILL_2__13170_ (
);

FILL FILL_3__11969_ (
);

FILL FILL_2__6716_ (
);

FILL FILL_3__11549_ (
);

FILL FILL_1__12583_ (
);

FILL FILL_1__12163_ (
);

FILL FILL_0__11996_ (
);

FILL FILL_0__9590_ (
);

FILL FILL_2__9188_ (
);

FILL FILL_0__9170_ (
);

AOI21X1 _11861_ (
    .A(_4968_),
    .B(_4967_),
    .C(_4918_),
    .Y(_4981_)
);

FILL FILL_0__11576_ (
);

INVX1 _11441_ (
    .A(_4625_),
    .Y(_4629_)
);

FILL FILL_0__11156_ (
);

INVX1 _11021_ (
    .A(\X[5] [7]),
    .Y(_4220_)
);

FILL FILL_3__12910_ (
);

FILL FILL_2__11903_ (
);

NAND3X1 _8648_ (
    .A(_2001_),
    .B(_2077_),
    .C(_2009_),
    .Y(_2084_)
);

NAND2X1 _8228_ (
    .A(\X[2] [1]),
    .B(vdd),
    .Y(_1669_)
);

FILL FILL_1__7185_ (
);

FILL FILL_0__7903_ (
);

FILL FILL_3__8472_ (
);

AOI21X1 _12646_ (
    .A(_5682_),
    .B(_5683_),
    .C(_5681_),
    .Y(_5687_)
);

OAI21X1 _12226_ (
    .A(_5293_),
    .B(_5334_),
    .C(_5333_),
    .Y(_5340_)
);

FILL FILL_0__13302_ (
);

FILL FILL_2__10295_ (
);

FILL FILL_1__9751_ (
);

FILL FILL_1__9331_ (
);

FILL FILL_3__9257_ (
);

FILL FILL_2__7674_ (
);

FILL FILL_3__12087_ (
);

OR2X2 _6714_ (
    .A(_307_),
    .B(_306_),
    .Y(_312_)
);

FILL FILL_2__12861_ (
);

FILL FILL_2__12441_ (
);

FILL FILL_2__12021_ (
);

OAI22X1 _9186_ (
    .A(_2433_),
    .B(_2544_),
    .C(_2476_),
    .D(_2545_),
    .Y(_2546_)
);

FILL FILL_1__11854_ (
);

FILL FILL_1__11434_ (
);

FILL FILL_1__11014_ (
);

FILL FILL_2__8879_ (
);

FILL FILL_0__8861_ (
);

FILL FILL_2__8459_ (
);

FILL FILL_0__8441_ (
);

FILL FILL_0__10847_ (
);

FILL FILL_0__10427_ (
);

DFFPOSX1 _10712_ (
    .D(_3978_[5]),
    .CLK(clk_bF$buf57),
    .Q(\Y[5] [5])
);

FILL FILL_2__8039_ (
);

FILL FILL_0__8021_ (
);

FILL FILL_0__10007_ (
);

NOR2X1 _13184_ (
    .A(_6211_),
    .B(_6212_),
    .Y(_6213_)
);

FILL FILL_2__9820_ (
);

FILL FILL_2__9400_ (
);

AND2X2 _7919_ (
    .A(\u_fir_pe1.rYin [0]),
    .B(\u_fir_pe1.mul [0]),
    .Y(_1428_)
);

FILL FILL_1__6876_ (
);

FILL FILL_1__6456_ (
);

FILL FILL_2__13226_ (
);

FILL FILL_1__12639_ (
);

FILL FILL_1__12219_ (
);

FILL FILL_0__9646_ (
);

FILL FILL_3__7743_ (
);

NAND2X1 _11917_ (
    .A(vdd),
    .B(\X[7]_5_bF$buf3 ),
    .Y(_5036_)
);

FILL FILL_0__9226_ (
);

FILL FILL_3__10153_ (
);

FILL FILL_0__10180_ (
);

FILL FILL_1__8602_ (
);

FILL FILL_3__8948_ (
);

FILL FILL_3__8528_ (
);

INVX1 _7672_ (
    .A(_1183_),
    .Y(_1189_)
);

DFFPOSX1 _7252_ (
    .D(_796_[13]),
    .CLK(clk_bF$buf1),
    .Q(\u_fir_pe0.mul [13])
);

FILL FILL_2__6945_ (
);

FILL FILL_2__6525_ (
);

FILL FILL_1__12392_ (
);

NAND3X1 _11670_ (
    .A(_4782_),
    .B(_4787_),
    .C(_4785_),
    .Y(_4793_)
);

FILL FILL_0__11385_ (
);

OAI21X1 _11250_ (
    .A(_4412_),
    .B(_4414_),
    .C(_4408_),
    .Y(_4446_)
);

FILL FILL_1__9807_ (
);

FILL FILL_2__11712_ (
);

NAND2X1 _8877_ (
    .A(_2299_),
    .B(_2300_),
    .Y(_2301_)
);

INVX1 _8457_ (
    .A(_1894_),
    .Y(_1895_)
);

NOR2X1 _8037_ (
    .A(_1539_),
    .B(_1540_),
    .Y(_1541_)
);

FILL FILL_1__10705_ (
);

FILL FILL_0__7712_ (
);

FILL FILL_1__13177_ (
);

NAND2X1 _12875_ (
    .A(_5904_),
    .B(_5912_),
    .Y(_5913_)
);

NOR2X1 _12455_ (
    .A(\u_fir_pe6.rYin [0]),
    .B(\u_fir_pe6.mul [0]),
    .Y(_5558_)
);

NAND3X1 _12035_ (
    .A(_5083_),
    .B(_5144_),
    .C(_5139_),
    .Y(_5153_)
);

FILL FILL_2__12917_ (
);

FILL FILL_0__13111_ (
);

FILL FILL_1__8199_ (
);

FILL FILL_0__8917_ (
);

FILL FILL_1__9980_ (
);

FILL FILL_1__9560_ (
);

FILL FILL_1__9140_ (
);

FILL FILL_3__9486_ (
);

FILL FILL_2__7483_ (
);

FILL FILL_2__7063_ (
);

AOI21X1 _6943_ (
    .A(_415_),
    .B(_407_),
    .C(_485_),
    .Y(_538_)
);

NAND3X1 _6523_ (
    .A(_53_),
    .B(_117_),
    .C(_118_),
    .Y(_124_)
);

FILL FILL_2__12670_ (
);

FILL FILL_2__12250_ (
);

FILL FILL_1__11663_ (
);

FILL FILL_3__10209_ (
);

FILL FILL_1__11243_ (
);

FILL FILL_2__8688_ (
);

FILL FILL_0__8670_ (
);

FILL FILL_0__8250_ (
);

FILL FILL_2__8268_ (
);

FILL FILL_0__10656_ (
);

NAND2X1 _10941_ (
    .A(gnd),
    .B(\X[5]_5_bF$buf1 ),
    .Y(_4141_)
);

OAI21X1 _10521_ (
    .A(_3751_),
    .B(_3764_),
    .C(_3768_),
    .Y(_3794_)
);

FILL FILL_0__10236_ (
);

AOI21X1 _10101_ (
    .A(_3380_),
    .B(_3379_),
    .C(_3378_),
    .Y(_3381_)
);

AOI21X1 _7728_ (
    .A(_1233_),
    .B(_1228_),
    .C(_1180_),
    .Y(_1245_)
);

NAND2X1 _7308_ (
    .A(gnd),
    .B(\X[1] [3]),
    .Y(_830_)
);

FILL FILL_1__6685_ (
);

FILL FILL_2__13035_ (
);

FILL FILL_1__12868_ (
);

FILL FILL_1__12448_ (
);

FILL FILL_1__12028_ (
);

FILL FILL_0__9455_ (
);

FILL FILL_0__9035_ (
);

OAI21X1 _11726_ (
    .A(_4835_),
    .B(_4847_),
    .C(_4841_),
    .Y(_4848_)
);

NAND2X1 _11306_ (
    .A(_4469_),
    .B(_4472_),
    .Y(_4501_)
);

FILL FILL_0__12802_ (
);

FILL FILL_3__10382_ (
);

FILL FILL_1__8831_ (
);

FILL FILL_1__8411_ (
);

FILL FILL_3__8337_ (
);

AOI21X1 _7481_ (
    .A(_917_),
    .B(_923_),
    .C(_1000_),
    .Y(_1001_)
);

INVX1 _7061_ (
    .A(\u_fir_pe0.rYin [3]),
    .Y(_648_)
);

FILL FILL_2__6754_ (
);

FILL FILL_3__11167_ (
);

FILL FILL_0__11194_ (
);

FILL FILL_1__9616_ (
);

FILL FILL_2__11941_ (
);

FILL FILL_2__11521_ (
);

FILL FILL_2__11101_ (
);

OAI22X1 _8686_ (
    .A(_1827_),
    .B(_1829_),
    .C(_1913_),
    .D(_1738_),
    .Y(_2121_)
);

OAI21X1 _8266_ (
    .A(_1702_),
    .B(_1703_),
    .C(_1663_),
    .Y(_1707_)
);

FILL FILL_1__10934_ (
);

FILL FILL_1__10514_ (
);

FILL FILL_2__7959_ (
);

FILL FILL_0__7941_ (
);

FILL FILL_0__7521_ (
);

FILL FILL_2__7539_ (
);

FILL FILL_2__7119_ (
);

FILL FILL_0__7101_ (
);

NAND2X1 _12684_ (
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5724_)
);

FILL FILL_0__12399_ (
);

NOR2X1 _12264_ (
    .A(_5017_),
    .B(_5244_),
    .Y(_5377_)
);

FILL FILL_2__8900_ (
);

FILL FILL_3__13313_ (
);

FILL FILL_2__12726_ (
);

FILL FILL_2__12306_ (
);

FILL FILL_1__11719_ (
);

FILL FILL_0__8726_ (
);

FILL FILL_3__6823_ (
);

FILL FILL_0__8306_ (
);

INVX1 _13049_ (
    .A(_6084_),
    .Y(_6085_)
);

FILL FILL_2__7292_ (
);

FILL FILL_3__7608_ (
);

NAND3X1 _6752_ (
    .A(_322_),
    .B(_340_),
    .C(_336_),
    .Y(_350_)
);

FILL FILL_1__11892_ (
);

FILL FILL_3__10438_ (
);

FILL FILL_1__11472_ (
);

FILL FILL_1__11052_ (
);

FILL FILL_2__8497_ (
);

FILL FILL_0__10885_ (
);

FILL FILL_0__10465_ (
);

DFFPOSX1 _10750_ (
    .D(_3982_[3]),
    .CLK(clk_bF$buf10),
    .Q(\u_fir_pe4.mul [3])
);

OAI21X1 _10330_ (
    .A(_3213_),
    .B(_3604_),
    .C(_3606_),
    .Y(_3607_)
);

FILL FILL_0__10045_ (
);

INVX1 _7957_ (
    .A(\u_fir_pe1.rYin [5]),
    .Y(_1462_)
);

AND2X2 _7537_ (
    .A(_1034_),
    .B(_1029_),
    .Y(_1056_)
);

AND2X2 _7117_ (
    .A(_659_),
    .B(_669_),
    .Y(_701_)
);

FILL FILL_1__6494_ (
);

FILL FILL_2__13264_ (
);

FILL FILL_1__12677_ (
);

FILL FILL_1__12257_ (
);

FILL FILL_0__9684_ (
);

FILL FILL_3__7781_ (
);

FILL FILL_0__9264_ (
);

AOI21X1 _11955_ (
    .A(_5069_),
    .B(_5068_),
    .C(_4970_),
    .Y(_5074_)
);

FILL FILL_3__7361_ (
);

NOR2X1 _11535_ (
    .A(\u_fir_pe5.rYin [11]),
    .B(\u_fir_pe5.mul [11]),
    .Y(_4719_)
);

OAI21X1 _11115_ (
    .A(_4074_),
    .B(_4129_),
    .C(_4312_),
    .Y(_4313_)
);

FILL FILL_0__12611_ (
);

FILL FILL_1__7699_ (
);

FILL FILL_1__7279_ (
);

FILL FILL_1__8640_ (
);

FILL FILL_1__8220_ (
);

FILL FILL_3__8566_ (
);

FILL FILL_3__8146_ (
);

NAND2X1 _7290_ (
    .A(_810_),
    .B(_806_),
    .Y(_813_)
);

FILL FILL_2__6983_ (
);

FILL FILL_2__6563_ (
);

FILL FILL_3__11396_ (
);

FILL FILL_2__10389_ (
);

FILL FILL_1__9425_ (
);

FILL FILL_2__11750_ (
);

FILL FILL_2__11330_ (
);

FILL FILL_0__6389_ (
);

NAND3X1 _8495_ (
    .A(_1918_),
    .B(_1920_),
    .C(_1922_),
    .Y(_1933_)
);

NOR2X1 _8075_ (
    .A(_1576_),
    .B(_1583_),
    .Y(_1590_[2])
);

FILL FILL_1__10323_ (
);

FILL FILL_2__7768_ (
);

FILL FILL_0__7750_ (
);

FILL FILL_2__7348_ (
);

FILL FILL_0__7330_ (
);

DFFPOSX1 _12493_ (
    .D(\Y[7] [8]),
    .CLK(clk_bF$buf46),
    .Q(\u_fir_pe6.rYin [8])
);

AND2X2 _12073_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5190_)
);

AND2X2 _6808_ (
    .A(gnd),
    .B(Xin[7]),
    .Y(_405_)
);

FILL FILL_2__12955_ (
);

FILL FILL_2__12535_ (
);

FILL FILL_2__12115_ (
);

FILL FILL_1__11948_ (
);

FILL FILL_1__11528_ (
);

FILL FILL_1__11108_ (
);

FILL FILL_0__8535_ (
);

NOR2X1 _10806_ (
    .A(_4008_),
    .B(_4007_),
    .Y(_4779_[3])
);

INVX1 _13278_ (
    .A(_6301_),
    .Y(_6302_)
);

FILL FILL_2__9914_ (
);

FILL FILL_1__7911_ (
);

FILL FILL_3__7837_ (
);

OAI21X1 _6981_ (
    .A(_573_),
    .B(_574_),
    .C(_526_),
    .Y(_575_)
);

INVX1 _6561_ (
    .A(_160_),
    .Y(_161_)
);

FILL FILL_1__11281_ (
);

FILL FILL_0__10694_ (
);

FILL FILL_0__10274_ (
);

FILL FILL_2__10601_ (
);

NAND2X1 _7766_ (
    .A(_1279_),
    .B(_1273_),
    .Y(_1282_)
);

NAND2X1 _7346_ (
    .A(\X[1] [0]),
    .B(gnd),
    .Y(_867_)
);

FILL FILL_2__13073_ (
);

FILL FILL_2__6619_ (
);

FILL FILL_0__6601_ (
);

FILL FILL_1__12066_ (
);

FILL FILL_0__9493_ (
);

FILL FILL_0__11899_ (
);

FILL FILL_3__7590_ (
);

FILL FILL_0__9073_ (
);

OAI21X1 _11764_ (
    .A(_4880_),
    .B(_4881_),
    .C(_4866_),
    .Y(_4885_)
);

FILL FILL_0__11479_ (
);

FILL FILL_3__7170_ (
);

FILL FILL_0__11059_ (
);

NAND3X1 _11344_ (
    .A(_4496_),
    .B(_4538_),
    .C(_4497_),
    .Y(_4539_)
);

FILL FILL_3__12813_ (
);

FILL FILL_2__11806_ (
);

FILL FILL_0__12840_ (
);

FILL FILL_0__12420_ (
);

FILL FILL_0__12000_ (
);

FILL FILL_1__7088_ (
);

FILL FILL_0__7806_ (
);

NOR2X1 _9912_ (
    .A(_3919_),
    .B(_3190_),
    .Y(_3195_)
);

FILL FILL_3__8795_ (
);

NAND2X1 _12969_ (
    .A(_5970_),
    .B(_5973_),
    .Y(_6006_)
);

NAND3X1 _12549_ (
    .A(_5589_),
    .B(_5591_),
    .C(_5590_),
    .Y(_5592_)
);

NOR3X1 _12129_ (
    .A(_5087_),
    .B(_4914_),
    .C(_5103_),
    .Y(_5245_)
);

FILL FILL_0__13205_ (
);

FILL FILL_2__6792_ (
);

FILL FILL_2__10198_ (
);

FILL FILL_1__9654_ (
);

FILL FILL_1__9234_ (
);

FILL FILL_1__10972_ (
);

FILL FILL_1__10552_ (
);

FILL FILL_1__10132_ (
);

FILL FILL_2__7997_ (
);

FILL FILL_2__7577_ (
);

FILL FILL_2__7157_ (
);

NAND2X1 _6617_ (
    .A(_213_),
    .B(_215_),
    .Y(_216_)
);

FILL FILL_2__12764_ (
);

FILL FILL_2__12344_ (
);

OR2X2 _9089_ (
    .A(_2450_),
    .B(_2449_),
    .Y(_2451_)
);

FILL FILL_1__11757_ (
);

FILL FILL_1__11337_ (
);

FILL FILL_0__8764_ (
);

FILL FILL_0__8344_ (
);

FILL FILL_3__6441_ (
);

INVX1 _10615_ (
    .A(\u_fir_pe4.rYin [8]),
    .Y(_3878_)
);

INVX1 _13087_ (
    .A(_6094_),
    .Y(_6122_)
);

FILL FILL_2__9723_ (
);

FILL FILL_2__9303_ (
);

FILL FILL_1__6779_ (
);

FILL FILL_2__13129_ (
);

FILL FILL_1__7720_ (
);

FILL FILL_1__7300_ (
);

FILL FILL_0__9969_ (
);

FILL FILL_0__9549_ (
);

FILL FILL_0__9129_ (
);

NOR2X1 _6790_ (
    .A(_318_),
    .B(_321_),
    .Y(_387_)
);

FILL FILL_3__10896_ (
);

FILL FILL_3__10476_ (
);

FILL FILL_3__10056_ (
);

FILL FILL_1__11090_ (
);

FILL FILL_0__10083_ (
);

FILL FILL_1__8925_ (
);

FILL FILL_1__8505_ (
);

FILL FILL_2__10830_ (
);

FILL FILL_2__10410_ (
);

NAND3X1 _7995_ (
    .A(_1498_),
    .B(_1495_),
    .C(_1458_),
    .Y(_1499_)
);

AOI21X1 _7575_ (
    .A(_1004_),
    .B(_1082_),
    .C(_1090_),
    .Y(_1093_)
);

AOI21X1 _7155_ (
    .A(_735_),
    .B(_726_),
    .C(_733_),
    .Y(_738_)
);

FILL FILL_0__6830_ (
);

FILL FILL_2__6848_ (
);

FILL FILL_0__6410_ (
);

FILL FILL_2__6428_ (
);

FILL FILL_1__12295_ (
);

AOI21X1 _11993_ (
    .A(_5110_),
    .B(_5108_),
    .C(_5106_),
    .Y(_5111_)
);

NAND2X1 _11573_ (
    .A(_4754_),
    .B(_4756_),
    .Y(_4757_)
);

FILL FILL_0__11288_ (
);

AOI21X1 _11153_ (
    .A(_4350_),
    .B(_4349_),
    .C(_4285_),
    .Y(_4351_)
);

FILL FILL_3__12622_ (
);

FILL FILL_1__10608_ (
);

FILL FILL254550x14550 (
);

FILL FILL_0__7615_ (
);

INVX1 _9721_ (
    .A(\u_fir_pe3.mul [6]),
    .Y(_3065_)
);

AOI21X1 _9301_ (
    .A(_2659_),
    .B(_2654_),
    .C(_2613_),
    .Y(_2660_)
);

NAND2X1 _12778_ (
    .A(_5811_),
    .B(_5816_),
    .Y(_5817_)
);

FILL FILL_3__8184_ (
);

AND2X2 _12358_ (
    .A(_5461_),
    .B(_5460_),
    .Y(_5572_[6])
);

FILL FILL_3__13407_ (
);

FILL FILL_0__13014_ (
);

FILL FILL_3__6917_ (
);

FILL FILL_1__9463_ (
);

FILL FILL_1__9043_ (
);

FILL FILL254250x21750 (
);

FILL FILL_1__10781_ (
);

FILL FILL_1__10361_ (
);

FILL FILL_2__7386_ (
);

INVX1 _6846_ (
    .A(_364_),
    .Y(_443_)
);

NOR2X1 _6426_ (
    .A(_27_),
    .B(_26_),
    .Y(_28_)
);

FILL FILL_2__12993_ (
);

FILL FILL_2__12573_ (
);

FILL FILL_2__12153_ (
);

FILL FILL_1__11986_ (
);

FILL FILL_1__11566_ (
);

FILL FILL_1__11146_ (
);

FILL FILL_0__8573_ (
);

FILL FILL_0__10979_ (
);

FILL FILL_3__6670_ (
);

FILL FILL_0__8153_ (
);

FILL FILL_0__10559_ (
);

NAND3X1 _10844_ (
    .A(_4013_),
    .B(_4030_),
    .C(_4033_),
    .Y(_4046_)
);

NAND3X1 _10424_ (
    .A(_3683_),
    .B(_3689_),
    .C(_3647_),
    .Y(_3699_)
);

FILL FILL_0__10139_ (
);

INVX1 _10004_ (
    .A(_3272_),
    .Y(_3285_)
);

FILL FILL_2__9952_ (
);

FILL FILL_2__9532_ (
);

FILL FILL_0__11920_ (
);

FILL FILL_2__9112_ (
);

FILL FILL_0__11500_ (
);

FILL FILL_1__6588_ (
);

FILL FILL_0__9778_ (
);

FILL FILL_0__9358_ (
);

FILL FILL_3__7455_ (
);

DFFPOSX1 _11629_ (
    .D(_4781_[5]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.mul [5])
);

FILL FILL_3__7035_ (
);

NAND2X1 _11209_ (
    .A(_4391_),
    .B(_4394_),
    .Y(_4406_)
);

FILL FILL_0__12705_ (
);

FILL FILL_1__8734_ (
);

FILL FILL_1__8314_ (
);

AOI21X1 _7384_ (
    .A(_900_),
    .B(_901_),
    .C(_899_),
    .Y(_905_)
);

FILL FILL_2__6657_ (
);

NOR2X1 _11382_ (
    .A(_4571_),
    .B(_4575_),
    .Y(_4781_[12])
);

FILL FILL_0__11097_ (
);

FILL FILL_1__9939_ (
);

FILL FILL_3__12851_ (
);

FILL FILL_1__9519_ (
);

FILL FILL_3__12011_ (
);

FILL FILL_2__11844_ (
);

FILL FILL_2__11424_ (
);

FILL FILL_2__11004_ (
);

INVX1 _8589_ (
    .A(_1948_),
    .Y(_2026_)
);

NAND2X1 _8169_ (
    .A(_1608_),
    .B(_1611_),
    .Y(_1612_)
);

FILL FILL_1__10837_ (
);

FILL FILL_1__10417_ (
);

FILL FILL_0__7844_ (
);

NAND3X1 _9950_ (
    .A(_3221_),
    .B(_3229_),
    .C(_3231_),
    .Y(_3232_)
);

FILL FILL_0__7424_ (
);

NAND3X1 _9530_ (
    .A(_2851_),
    .B(_2885_),
    .C(_2883_),
    .Y(_2886_)
);

FILL FILL_0__7004_ (
);

NAND3X1 _9110_ (
    .A(\X[3] [1]),
    .B(gnd),
    .C(_2470_),
    .Y(_2471_)
);

NAND2X1 _12587_ (
    .A(_5611_),
    .B(_5626_),
    .Y(_5629_)
);

NAND3X1 _12167_ (
    .A(_5278_),
    .B(_5279_),
    .C(_5282_),
    .Y(_5283_)
);

FILL FILL_2__8803_ (
);

FILL FILL_2__12629_ (
);

FILL FILL_2__12209_ (
);

FILL FILL_0__13243_ (
);

FILL FILL_1__6800_ (
);

FILL FILL_0__8629_ (
);

FILL FILL_0__8209_ (
);

FILL FILL_1__9692_ (
);

FILL FILL_1__9272_ (
);

FILL FILL_3__9198_ (
);

FILL FILL_1__10590_ (
);

FILL FILL_1__10170_ (
);

FILL FILL_2__7195_ (
);

NAND2X1 _6655_ (
    .A(vdd),
    .B(Xin_5_bF$buf0),
    .Y(_254_)
);

FILL FILL_2__12382_ (
);

FILL FILL_1__11795_ (
);

FILL FILL_1__11375_ (
);

FILL FILL_0__8382_ (
);

FILL FILL_0__10788_ (
);

NAND2X1 _10653_ (
    .A(_3916_),
    .B(_3911_),
    .Y(_3917_)
);

FILL FILL_0__10368_ (
);

OAI21X1 _10233_ (
    .A(_3428_),
    .B(_3436_),
    .C(_3435_),
    .Y(_3511_)
);

FILL FILL_2__9761_ (
);

FILL FILL_2__9341_ (
);

FILL FILL_1__6397_ (
);

FILL FILL_2__13167_ (
);

NOR2X1 _8801_ (
    .A(_2229_),
    .B(_2228_),
    .Y(_2230_)
);

FILL FILL_0__9587_ (
);

FILL FILL_3__7684_ (
);

FILL FILL_0__9167_ (
);

NAND3X1 _11858_ (
    .A(_4972_),
    .B(_4973_),
    .C(_4974_),
    .Y(_4978_)
);

AND2X2 _11438_ (
    .A(\u_fir_pe5.rYin [2]),
    .B(\u_fir_pe5.mul [2]),
    .Y(_4626_)
);

NAND3X1 _11018_ (
    .A(_4211_),
    .B(_4216_),
    .C(_4214_),
    .Y(_4217_)
);

FILL FILL_3__12907_ (
);

FILL FILL_1__13101_ (
);

FILL FILL_0__12934_ (
);

FILL FILL_3__10094_ (
);

FILL FILL_1__8543_ (
);

FILL FILL_3__8889_ (
);

FILL FILL_3__8469_ (
);

FILL FILL_3__8049_ (
);

NOR2X1 _7193_ (
    .A(\u_fir_pe0.rYin [0]),
    .B(\u_fir_pe0.mul [0]),
    .Y(_776_)
);

FILL FILL_3__9410_ (
);

FILL FILL_2__6886_ (
);

FILL FILL_2__6466_ (
);

OAI22X1 _11191_ (
    .A(_4239_),
    .B(_4386_),
    .C(_4309_),
    .D(_4387_),
    .Y(_4388_)
);

FILL FILL_1__9748_ (
);

FILL FILL_1__9328_ (
);

FILL FILL_3__12240_ (
);

FILL FILL_2__11653_ (
);

FILL FILL_2__11233_ (
);

NAND2X1 _8398_ (
    .A(_1835_),
    .B(_1836_),
    .Y(_1837_)
);

FILL FILL_1__10646_ (
);

FILL FILL_1__10226_ (
);

FILL FILL_0__7653_ (
);

NAND2X1 _12396_ (
    .A(_5499_),
    .B(_5498_),
    .Y(_5572_[9])
);

FILL FILL_2__8612_ (
);

FILL FILL_3__13025_ (
);

FILL FILL_2__12858_ (
);

FILL FILL_2__12438_ (
);

FILL FILL_2__12018_ (
);

FILL FILL_0__13052_ (
);

FILL FILL_0__8858_ (
);

FILL FILL_0__8438_ (
);

FILL FILL_3__6535_ (
);

DFFPOSX1 _10709_ (
    .D(_3978_[2]),
    .CLK(clk_bF$buf6),
    .Q(\Y[5] [2])
);

FILL FILL_0__8018_ (
);

FILL FILL_1__9081_ (
);

FILL FILL_2__9817_ (
);

FILL FILL_1__7814_ (
);

OAI21X1 _6884_ (
    .A(_74_),
    .B(_319_),
    .C(_473_),
    .Y(_480_)
);

OAI21X1 _6464_ (
    .A(_53_),
    .B(_65_),
    .C(_59_),
    .Y(_66_)
);

FILL FILL_2__12191_ (
);

FILL FILL_1__11184_ (
);

FILL FILL_0__8191_ (
);

FILL FILL_0__10597_ (
);

AOI21X1 _10882_ (
    .A(_4077_),
    .B(_4079_),
    .C(_4070_),
    .Y(_4083_)
);

AOI21X1 _10462_ (
    .A(_3675_),
    .B(_3679_),
    .C(_3649_),
    .Y(_3737_)
);

FILL FILL_0__10177_ (
);

OR2X2 _10042_ (
    .A(_3321_),
    .B(_3319_),
    .Y(_3322_)
);

FILL FILL254250x241350 (
);

FILL FILL_2__10924_ (
);

FILL FILL_2__9990_ (
);

FILL FILL_2__9570_ (
);

FILL FILL_2__10504_ (
);

FILL FILL_2__9150_ (
);

INVX1 _7669_ (
    .A(_1185_),
    .Y(_1186_)
);

DFFPOSX1 _7249_ (
    .D(_796_[10]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.mul [10])
);

FILL FILL_2__13396_ (
);

FILL FILL_0__6924_ (
);

FILL FILL_0__6504_ (
);

NAND2X1 _8610_ (
    .A(_2046_),
    .B(_2045_),
    .Y(_2390_[9])
);

FILL FILL_1__12389_ (
);

FILL FILL_0__9396_ (
);

OAI21X1 _11667_ (
    .A(_4786_),
    .B(_4789_),
    .C(_4782_),
    .Y(_4790_)
);

INVX1 _11247_ (
    .A(_4442_),
    .Y(_4443_)
);

FILL FILL_1__13330_ (
);

FILL FILL_2__11709_ (
);

FILL FILL_0__12743_ (
);

FILL FILL254250x208950 (
);

FILL FILL_0__12323_ (
);

FILL FILL_0__7709_ (
);

INVX1 _9815_ (
    .A(_3153_),
    .Y(_3158_)
);

FILL FILL_1__8772_ (
);

FILL FILL_1__8352_ (
);

FILL FILL_3__8278_ (
);

FILL FILL_0__13108_ (
);

FILL FILL_2__6695_ (
);

FILL FILL_1__9977_ (
);

FILL FILL_1__9557_ (
);

FILL FILL_1__9137_ (
);

FILL FILL_2__11882_ (
);

FILL FILL_2__11462_ (
);

FILL FILL_2__11042_ (
);

FILL FILL_1__10875_ (
);

FILL FILL_1__10455_ (
);

FILL FILL_1__10035_ (
);

FILL FILL254550x64950 (
);

FILL FILL_0__7882_ (
);

FILL FILL_0__7462_ (
);

FILL FILL_0__7042_ (
);

FILL FILL_2__8841_ (
);

FILL FILL_2__8421_ (
);

FILL FILL_3__13254_ (
);

FILL FILL_2__8001_ (
);

FILL FILL_2__12667_ (
);

FILL FILL_2__12247_ (
);

FILL FILL_0__13281_ (
);

FILL FILL_0__8667_ (
);

FILL FILL_3__6764_ (
);

FILL FILL_0__8247_ (
);

NAND2X1 _10938_ (
    .A(vdd),
    .B(\X[5] [3]),
    .Y(_4138_)
);

OR2X2 _10518_ (
    .A(_3789_),
    .B(_3782_),
    .Y(_3791_)
);

FILL FILL_1__12601_ (
);

FILL FILL_2__9626_ (
);

FILL FILL_2__9206_ (
);

FILL FILL_1__7623_ (
);

FILL FILL_3__7549_ (
);

FILL FILL_3__7129_ (
);

AOI21X1 _6693_ (
    .A(_287_),
    .B(_286_),
    .C(_188_),
    .Y(_292_)
);

FILL FILL_3__8910_ (
);

FILL FILL_3__10379_ (
);

NOR2X1 _10691_ (
    .A(_3954_),
    .B(_3953_),
    .Y(_3978_[14])
);

NAND3X1 _10271_ (
    .A(_3503_),
    .B(_3534_),
    .C(_3539_),
    .Y(_3549_)
);

FILL FILL_1__8828_ (
);

FILL FILL_3__11740_ (
);

FILL FILL_1__8408_ (
);

FILL FILL_3__11320_ (
);

FILL FILL_2__10313_ (
);

NAND2X1 _7898_ (
    .A(_1410_),
    .B(_1407_),
    .Y(_1593_[13])
);

OAI21X1 _7478_ (
    .A(_996_),
    .B(_997_),
    .C(_995_),
    .Y(_998_)
);

NAND2X1 _7058_ (
    .A(_645_),
    .B(_644_),
    .Y(_646_)
);

FILL FILL_0__6733_ (
);

FILL FILL_1__12198_ (
);

INVX1 _11896_ (
    .A(gnd),
    .Y(_5015_)
);

NOR2X1 _11476_ (
    .A(_4658_),
    .B(_4659_),
    .Y(_4660_)
);

AND2X2 _11056_ (
    .A(_4206_),
    .B(_4203_),
    .Y(_4255_)
);

FILL FILL_3__12945_ (
);

FILL FILL_3__12525_ (
);

FILL FILL_3__12105_ (
);

FILL FILL_2__11938_ (
);

FILL FILL_0__12972_ (
);

FILL FILL_2__11518_ (
);

FILL FILL_0__12552_ (
);

FILL FILL_0__12132_ (
);

FILL FILL_0__7938_ (
);

FILL FILL_0__7518_ (
);

NAND3X1 _9624_ (
    .A(_2768_),
    .B(_2841_),
    .C(_2947_),
    .Y(_2978_)
);

NAND2X1 _9204_ (
    .A(_2542_),
    .B(_2538_),
    .Y(_2564_)
);

FILL FILL_1__8581_ (
);

FILL FILL_1__8161_ (
);

FILL FILL_0__13337_ (
);

NOR2X1 _13202_ (
    .A(_6227_),
    .B(_6228_),
    .Y(_6229_)
);

FILL FILL_1__9786_ (
);

FILL FILL_1__9366_ (
);

FILL FILL_2__11691_ (
);

FILL FILL_2__11271_ (
);

FILL FILL_1__10684_ (
);

FILL FILL_1__10264_ (
);

FILL FILL_0__7691_ (
);

FILL FILL_0__7271_ (
);

FILL FILL_2__7289_ (
);

FILL FILL_2__8650_ (
);

FILL FILL_2__8230_ (
);

FILL FILL_3__13063_ (
);

INVX1 _6749_ (
    .A(_260_),
    .Y(_347_)
);

FILL FILL_2__12896_ (
);

FILL FILL_2__12056_ (
);

FILL FILL_0__13090_ (
);

FILL FILL_1__11889_ (
);

FILL FILL_1__11469_ (
);

FILL FILL_1__11049_ (
);

FILL FILL_0__8896_ (
);

FILL FILL_3__6993_ (
);

FILL FILL_0__8476_ (
);

DFFPOSX1 _10747_ (
    .D(_3979_[0]),
    .CLK(clk_bF$buf38),
    .Q(\u_fir_pe4.mul [0])
);

FILL FILL_0__8056_ (
);

NAND2X1 _10327_ (
    .A(\X[4]_5_bF$buf0 ),
    .B(vdd),
    .Y(_3604_)
);

FILL FILL_1__12830_ (
);

FILL FILL_1__12410_ (
);

FILL FILL_2__9435_ (
);

FILL FILL_0__11823_ (
);

FILL FILL_2__9015_ (
);

FILL FILL_0__11403_ (
);

FILL FILL_1__7852_ (
);

FILL FILL_1__7432_ (
);

FILL FILL_1__7012_ (
);

FILL FILL_3__7778_ (
);

FILL FILL_0__12608_ (
);

NAND3X1 _10080_ (
    .A(_3355_),
    .B(_3340_),
    .C(_3359_),
    .Y(_3360_)
);

FILL FILL_1__8637_ (
);

FILL FILL_1__8217_ (
);

FILL FILL_2__10962_ (
);

FILL FILL_2__10542_ (
);

FILL FILL_2__10122_ (
);

NAND3X1 _7287_ (
    .A(_807_),
    .B(_809_),
    .C(_808_),
    .Y(_810_)
);

FILL FILL_3__9924_ (
);

FILL FILL_3__9504_ (
);

FILL FILL_0__6962_ (
);

FILL FILL_0__6542_ (
);

INVX1 _11285_ (
    .A(_4445_),
    .Y(_4481_)
);

FILL FILL_2__7921_ (
);

FILL FILL_2__7501_ (
);

FILL FILL_3__12334_ (
);

FILL FILL_2__11747_ (
);

FILL FILL_0__12781_ (
);

FILL FILL_2__11327_ (
);

FILL FILL_0__12361_ (
);

FILL FILL_0__7747_ (
);

DFFPOSX1 _9853_ (
    .D(\X[3] [7]),
    .CLK(clk_bF$buf42),
    .Q(\X[4] [7])
);

FILL FILL_0__7327_ (
);

AND2X2 _9433_ (
    .A(_2523_),
    .B(_2712_),
    .Y(_2790_)
);

NAND2X1 _9013_ (
    .A(gnd),
    .B(\X[3] [1]),
    .Y(_3122_)
);

FILL FILL_1__8390_ (
);

FILL FILL_2__8706_ (
);

FILL FILL_3__13119_ (
);

FILL FILL_0__13146_ (
);

NAND2X1 _13011_ (
    .A(gnd),
    .B(_5977_),
    .Y(_6047_)
);

FILL FILL_1__6703_ (
);

FILL FILL_3__6629_ (
);

FILL FILL_1__9595_ (
);

FILL FILL_1__9175_ (
);

FILL FILL_2__11080_ (
);

FILL FILL_1__10493_ (
);

FILL FILL_1__10073_ (
);

FILL FILL_2__7098_ (
);

FILL FILL_0__7080_ (
);

FILL FILL_1__7908_ (
);

FILL FILL_3__10820_ (
);

FILL FILL_3__13292_ (
);

NAND3X1 _6978_ (
    .A(_564_),
    .B(_571_),
    .C(_570_),
    .Y(_572_)
);

AND2X2 _6558_ (
    .A(gnd),
    .B(Xin[4]),
    .Y(_158_)
);

FILL FILL_2__12285_ (
);

FILL FILL_1__11698_ (
);

FILL FILL_1__11278_ (
);

FILL FILL_0__8285_ (
);

NAND3X1 _10976_ (
    .A(_4169_),
    .B(_4162_),
    .C(_4167_),
    .Y(_4176_)
);

FILL FILL_3__6382_ (
);

NAND2X1 _10556_ (
    .A(_3819_),
    .B(_3824_),
    .Y(_3825_)
);

AND2X2 _10136_ (
    .A(\X[4] [3]),
    .B(gnd),
    .Y(_3415_)
);

FILL FILL_2__9664_ (
);

FILL FILL_2__9244_ (
);

FILL FILL_0__11212_ (
);

NAND2X1 _8704_ (
    .A(_2133_),
    .B(_2130_),
    .Y(_2139_)
);

FILL FILL_1__7661_ (
);

FILL FILL_1__13004_ (
);

FILL FILL_0__12837_ (
);

NAND3X1 _12702_ (
    .A(vdd),
    .B(\X[6] [4]),
    .C(_5732_),
    .Y(_5742_)
);

FILL FILL_0__12417_ (
);

AOI22X1 _9909_ (
    .A(gnd),
    .B(\X[4] [0]),
    .C(gnd),
    .D(\X[4] [1]),
    .Y(_3192_)
);

FILL FILL_1__8866_ (
);

FILL FILL_1__8446_ (
);

FILL FILL_1__8026_ (
);

FILL FILL_2__10771_ (
);

FILL FILL_2__10351_ (
);

AND2X2 _7096_ (
    .A(_679_),
    .B(_678_),
    .Y(_790_[6])
);

FILL FILL_3__9733_ (
);

FILL FILL_2__6789_ (
);

FILL FILL_0__6771_ (
);

OAI21X1 _11094_ (
    .A(_4210_),
    .B(_4215_),
    .C(_4214_),
    .Y(_4292_)
);

FILL FILL_2__7730_ (
);

FILL FILL_3__12563_ (
);

FILL FILL_2__7310_ (
);

FILL FILL_2__11976_ (
);

FILL FILL_2__11556_ (
);

FILL FILL_0__12590_ (
);

FILL FILL_2__11136_ (
);

FILL FILL_0__12170_ (
);

FILL FILL_1__10969_ (
);

FILL FILL_1__10549_ (
);

FILL FILL_1__10129_ (
);

FILL FILL_0__7976_ (
);

FILL FILL_0__7556_ (
);

INVX1 _9662_ (
    .A(_2973_),
    .Y(_3014_)
);

FILL FILL_0__7136_ (
);

NAND2X1 _9242_ (
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2601_)
);

FILL FILL_1__11910_ (
);

NAND2X1 _12299_ (
    .A(_5410_),
    .B(_5404_),
    .Y(_5578_[14])
);

FILL FILL_2__8935_ (
);

FILL FILL_2__8515_ (
);

FILL FILL_0__10903_ (
);

NOR2X1 _13240_ (
    .A(\u_fir_pe7.rYin [7]),
    .B(\u_fir_pe7.mul [7]),
    .Y(_6263_)
);

FILL FILL_1__6932_ (
);

FILL FILL_1__6512_ (
);

FILL FILL_3__6858_ (
);

FILL FILL_0__9702_ (
);

FILL FILL_1__7717_ (
);

AOI21X1 _6787_ (
    .A(_349_),
    .B(_350_),
    .C(_317_),
    .Y(_384_)
);

FILL FILL_2__12094_ (
);

FILL FILL_1__11087_ (
);

OR2X2 _10785_ (
    .A(_4716_),
    .B(_3987_),
    .Y(_3988_)
);

NAND2X1 _10365_ (
    .A(_3630_),
    .B(_3637_),
    .Y(_3641_)
);

FILL FILL_3__11834_ (
);

FILL FILL_3__11414_ (
);

FILL FILL_2__10827_ (
);

FILL FILL_2__9893_ (
);

FILL FILL_2__9473_ (
);

FILL FILL_0__11861_ (
);

FILL FILL_2__10407_ (
);

FILL FILL_2__9053_ (
);

FILL FILL_0__11441_ (
);

FILL FILL_0__11021_ (
);

FILL FILL_2__13299_ (
);

FILL FILL_0__6827_ (
);

NOR2X1 _8933_ (
    .A(\u_fir_pe2.rYin [14]),
    .B(\u_fir_pe2.mul [14]),
    .Y(_2357_)
);

FILL FILL_0__6407_ (
);

OAI21X1 _8513_ (
    .A(_1950_),
    .B(_1946_),
    .C(_1897_),
    .Y(_1951_)
);

FILL FILL_1__7890_ (
);

FILL FILL_1__7470_ (
);

FILL FILL_1__7050_ (
);

FILL FILL_0__9299_ (
);

FILL FILL_3__7396_ (
);

FILL FILL_3__12619_ (
);

FILL FILL_1__13233_ (
);

INVX1 _12931_ (
    .A(_5967_),
    .Y(_5968_)
);

FILL FILL_0__12646_ (
);

FILL FILL_0__12226_ (
);

DFFPOSX1 _12511_ (
    .D(_5578_[10]),
    .CLK(clk_bF$buf23),
    .Q(\u_fir_pe6.mul [10])
);

AND2X2 _9718_ (
    .A(_3062_),
    .B(_3061_),
    .Y(_3181_[5])
);

FILL FILL_1__8675_ (
);

FILL FILL_1__8255_ (
);

FILL FILL_2__10580_ (
);

FILL FILL_2__10160_ (
);

FILL FILL_3__9122_ (
);

FILL FILL_0__6580_ (
);

FILL FILL_2__6598_ (
);

FILL FILL_3__12792_ (
);

FILL FILL_2__11785_ (
);

FILL FILL_2__11365_ (
);

FILL FILL_1__10778_ (
);

FILL FILL_1__10358_ (
);

FILL FILL_0__7785_ (
);

NOR2X1 _9891_ (
    .A(_3877_),
    .B(_3919_),
    .Y(_3928_)
);

FILL FILL_0__7365_ (
);

NAND3X1 _9471_ (
    .A(_2774_),
    .B(_2822_),
    .C(_2827_),
    .Y(_2828_)
);

AOI21X1 _9051_ (
    .A(_2410_),
    .B(_2411_),
    .C(_3177_),
    .Y(_2414_)
);

FILL FILL_2__8744_ (
);

FILL FILL_2__8324_ (
);

FILL FILL_0__13184_ (
);

FILL FILL_1__6741_ (
);

FILL FILL_1__12924_ (
);

FILL FILL_0__9931_ (
);

FILL FILL_2__9949_ (
);

FILL FILL_2__9529_ (
);

FILL FILL_0__11917_ (
);

FILL FILL_0__9511_ (
);

FILL FILL_2__9109_ (
);

FILL FILL_1__7946_ (
);

FILL FILL_1__7526_ (
);

FILL FILL_1__7106_ (
);

NAND3X1 _6596_ (
    .A(_190_),
    .B(_191_),
    .C(_192_),
    .Y(_196_)
);

OR2X2 _10594_ (
    .A(_3852_),
    .B(_3857_),
    .Y(_3859_)
);

AOI21X1 _10174_ (
    .A(_3340_),
    .B(_3359_),
    .C(_3452_),
    .Y(_3453_)
);

FILL FILL_2__6810_ (
);

FILL FILL_2__10636_ (
);

FILL FILL_2__9282_ (
);

FILL FILL_0__11670_ (
);

FILL FILL_2__10216_ (
);

FILL FILL_0__11250_ (
);

FILL FILL_0__6636_ (
);

OAI21X1 _8742_ (
    .A(_2173_),
    .B(_2175_),
    .C(_2154_),
    .Y(_2176_)
);

INVX1 _8322_ (
    .A(_1749_),
    .Y(_1762_)
);

AOI21X1 _11799_ (
    .A(_4873_),
    .B(_4877_),
    .C(_4866_),
    .Y(_4919_)
);

OAI21X1 _11379_ (
    .A(_4361_),
    .B(_4572_),
    .C(_4544_),
    .Y(_4573_)
);

FILL FILL_3__12848_ (
);

FILL FILL_3__12428_ (
);

FILL FILL_1__13042_ (
);

FILL FILL_0__12875_ (
);

OAI21X1 _12740_ (
    .A(_5778_),
    .B(_5779_),
    .C(_5777_),
    .Y(_5780_)
);

FILL FILL_0__12455_ (
);

FILL FILL_0__12035_ (
);

NAND2X1 _12320_ (
    .A(_5427_),
    .B(_5426_),
    .Y(_5428_)
);

NAND3X1 _9947_ (
    .A(gnd),
    .B(\X[4] [2]),
    .C(_3219_),
    .Y(_3229_)
);

NAND3X1 _9527_ (
    .A(_2878_),
    .B(_2882_),
    .C(_2852_),
    .Y(_2883_)
);

NAND3X1 _9107_ (
    .A(_2467_),
    .B(_2462_),
    .C(_2464_),
    .Y(_2468_)
);

FILL FILL_1__8484_ (
);

FILL FILL_1__8064_ (
);

FILL FILL_3__9351_ (
);

AND2X2 _13105_ (
    .A(_6121_),
    .B(_6116_),
    .Y(_6139_)
);

FILL FILL_1__9689_ (
);

FILL FILL_1__9269_ (
);

FILL FILL_3__12181_ (
);

FILL FILL_2__11174_ (
);

FILL FILL_1__10587_ (
);

FILL FILL_1__10167_ (
);

FILL FILL_0__7594_ (
);

FILL FILL_0__7174_ (
);

AOI22X1 _9280_ (
    .A(gnd),
    .B(\X[3] [4]),
    .C(gnd),
    .D(\X[3]_5_bF$buf2 ),
    .Y(_2639_)
);

FILL FILL_3__10914_ (
);

FILL FILL_2__8553_ (
);

FILL FILL_0__10941_ (
);

FILL FILL_2__8133_ (
);

FILL FILL_0__10521_ (
);

FILL FILL_0__10101_ (
);

FILL FILL_2__12799_ (
);

FILL FILL_2__12379_ (
);

FILL FILL_1__6970_ (
);

FILL FILL_1__6550_ (
);

FILL FILL_0__8799_ (
);

FILL FILL_2__13320_ (
);

FILL FILL_0__8379_ (
);

FILL FILL_3__6476_ (
);

FILL FILL_1__12733_ (
);

FILL FILL_1__12313_ (
);

FILL FILL_0__9740_ (
);

FILL FILL_2__9758_ (
);

FILL FILL_0__9320_ (
);

FILL FILL_2__9338_ (
);

FILL FILL_0__11726_ (
);

FILL FILL_0__11306_ (
);

FILL FILL_1__7755_ (
);

FILL FILL_1__7335_ (
);

FILL FILL_3__8622_ (
);

FILL FILL_3__11032_ (
);

FILL FILL_2__10865_ (
);

FILL FILL_2__10445_ (
);

FILL FILL_2__9091_ (
);

FILL FILL_2__10025_ (
);

FILL FILL_1__9901_ (
);

FILL FILL_3__9827_ (
);

FILL FILL_3__9407_ (
);

FILL FILL_0__6865_ (
);

DFFPOSX1 _8971_ (
    .D(\X[2] [2]),
    .CLK(clk_bF$buf28),
    .Q(\X[3] [2])
);

FILL FILL_0__6445_ (
);

NAND3X1 _8551_ (
    .A(_1986_),
    .B(_1982_),
    .C(_1987_),
    .Y(_1988_)
);

DFFPOSX1 _8131_ (
    .D(_1593_[15]),
    .CLK(clk_bF$buf43),
    .Q(\u_fir_pe1.mul [15])
);

NOR2X1 _11188_ (
    .A(_4383_),
    .B(_4384_),
    .Y(_4385_)
);

FILL FILL_2__7824_ (
);

FILL FILL_2__7404_ (
);

FILL FILL_1__13271_ (
);

FILL FILL_0__12684_ (
);

FILL FILL_0__12264_ (
);

INVX1 _9756_ (
    .A(_3083_),
    .Y(_3099_)
);

OAI21X1 _9336_ (
    .A(_2613_),
    .B(_2693_),
    .C(_2662_),
    .Y(_2694_)
);

FILL FILL_1__8293_ (
);

FILL FILL_2__8609_ (
);

FILL FILL_3__9580_ (
);

FILL FILL_0__13049_ (
);

AOI21X1 _13334_ (
    .A(\X[6] [0]),
    .B(gnd),
    .C(_6279_),
    .Y(_6356_)
);

FILL FILL_1__6606_ (
);

FILL FILL_1__9498_ (
);

FILL FILL_1__9078_ (
);

FILL FILL_1__10396_ (
);

FILL FILL_3__10303_ (
);

FILL FILL_2__8782_ (
);

FILL FILL_2__8362_ (
);

FILL FILL_0__10330_ (
);

FILL FILL_2__12188_ (
);

NAND2X1 _7822_ (
    .A(_1329_),
    .B(_1332_),
    .Y(_1337_)
);

NAND3X1 _7402_ (
    .A(_917_),
    .B(_922_),
    .C(_864_),
    .Y(_923_)
);

FILL FILL_0__8188_ (
);

NAND3X1 _10879_ (
    .A(_4070_),
    .B(_4077_),
    .C(_4079_),
    .Y(_4080_)
);

NAND3X1 _10459_ (
    .A(_3731_),
    .B(_3733_),
    .C(_3732_),
    .Y(_3734_)
);

AND2X2 _10039_ (
    .A(\X[4] [0]),
    .B(gnd),
    .Y(_3319_)
);

FILL FILL_3__11928_ (
);

FILL FILL_1__12962_ (
);

FILL FILL_1__12542_ (
);

FILL FILL_1__12122_ (
);

FILL FILL_2__9987_ (
);

FILL FILL_2__9567_ (
);

FILL FILL_0__11955_ (
);

FILL FILL_2__9147_ (
);

AND2X2 _11820_ (
    .A(gnd),
    .B(\X[7] [4]),
    .Y(_4940_)
);

FILL FILL_0__11535_ (
);

NAND2X1 _11400_ (
    .A(_4591_),
    .B(_4592_),
    .Y(_4593_)
);

FILL FILL_0__11115_ (
);

AND2X2 _8607_ (
    .A(_2043_),
    .B(_2036_),
    .Y(_2044_)
);

FILL FILL_1__7984_ (
);

FILL FILL_1__7564_ (
);

FILL FILL_1__7144_ (
);

FILL FILL_1__13327_ (
);

NOR2X1 _12605_ (
    .A(_5600_),
    .B(_5637_),
    .Y(_5646_)
);

FILL FILL_1__8769_ (
);

FILL FILL_3__11681_ (
);

FILL FILL_1__8349_ (
);

FILL FILL_3__11261_ (
);

FILL FILL_2__10674_ (
);

FILL FILL_2__10254_ (
);

FILL FILL_1__9710_ (
);

FILL FILL_3__9216_ (
);

FILL FILL_0__6674_ (
);

AND2X2 _8780_ (
    .A(_2190_),
    .B(_2189_),
    .Y(_2212_)
);

AOI21X1 _8360_ (
    .A(_1788_),
    .B(_1796_),
    .C(_1799_),
    .Y(_1800_)
);

FILL FILL_3__12886_ (
);

FILL FILL_2__7633_ (
);

FILL FILL_3__12046_ (
);

FILL FILL_1__13080_ (
);

FILL FILL_2__11879_ (
);

FILL FILL_2__11459_ (
);

FILL FILL_2__11039_ (
);

FILL FILL_0__12073_ (
);

FILL FILL_2__12820_ (
);

FILL FILL_2__12400_ (
);

FILL FILL_0__7879_ (
);

NAND3X1 _9985_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf1 ),
    .C(_3263_),
    .Y(_3266_)
);

FILL FILL_0__7459_ (
);

NAND3X1 _9565_ (
    .A(_2916_),
    .B(_2919_),
    .C(_2873_),
    .Y(_2920_)
);

FILL FILL_0__7039_ (
);

NAND3X1 _9145_ (
    .A(_2503_),
    .B(_2504_),
    .C(_2505_),
    .Y(_2506_)
);

FILL FILL_1__11813_ (
);

FILL FILL_0__8820_ (
);

FILL FILL_2__8838_ (
);

FILL FILL_0__8400_ (
);

FILL FILL_2__8418_ (
);

FILL FILL_0__10806_ (
);

FILL FILL_0__13278_ (
);

OAI22X1 _13143_ (
    .A(_5723_),
    .B(_6041_),
    .C(_5884_),
    .D(_5814_),
    .Y(_6176_)
);

FILL FILL_1__6835_ (
);

FILL FILL_1__6415_ (
);

FILL FILL_0__9605_ (
);

FILL FILL_3__7702_ (
);

FILL FILL_3__10532_ (
);

FILL FILL_2__8591_ (
);

FILL FILL_2__8171_ (
);

AOI21X1 _7631_ (
    .A(_1148_),
    .B(_1143_),
    .C(_1112_),
    .Y(_1149_)
);

DFFPOSX1 _7211_ (
    .D(_790_[12]),
    .CLK(clk_bF$buf54),
    .Q(\Y[1] [12])
);

NOR2X1 _10688_ (
    .A(_3951_),
    .B(_3950_),
    .Y(_3952_)
);

INVX1 _10268_ (
    .A(_3459_),
    .Y(_3546_)
);

FILL FILL_2__6904_ (
);

FILL FILL_1__12771_ (
);

FILL FILL_3__11317_ (
);

FILL FILL_1__12351_ (
);

FILL FILL_2__9796_ (
);

FILL FILL_2__9376_ (
);

FILL FILL_0__11764_ (
);

FILL FILL_0__11344_ (
);

NOR2X1 _8836_ (
    .A(_2259_),
    .B(_2260_),
    .Y(_2261_)
);

OAI21X1 _8416_ (
    .A(_1844_),
    .B(_1839_),
    .C(_1846_),
    .Y(_1855_)
);

FILL FILL_1__7793_ (
);

FILL FILL_1__7373_ (
);

FILL FILL_1__13136_ (
);

FILL FILL_0__12969_ (
);

FILL FILL_3__8660_ (
);

OAI21X1 _12834_ (
    .A(_5871_),
    .B(_5872_),
    .C(_5870_),
    .Y(_5873_)
);

FILL FILL_0__12549_ (
);

FILL FILL_3__8240_ (
);

FILL FILL_0__12129_ (
);

NOR2X1 _12414_ (
    .A(_5517_),
    .B(_5514_),
    .Y(_5518_)
);

FILL FILL_1__8578_ (
);

FILL FILL_1__8158_ (
);

FILL FILL_3__11490_ (
);

FILL FILL_2__10483_ (
);

FILL FILL_2__10063_ (
);

FILL FILL_3__9445_ (
);

FILL FILL_3__9025_ (
);

FILL FILL_0__6483_ (
);

FILL FILL_2__7862_ (
);

FILL FILL_2__7442_ (
);

FILL FILL_3__12275_ (
);

FILL FILL_2__7022_ (
);

FILL FILL_2__11688_ (
);

FILL FILL_2__11268_ (
);

AOI21X1 _6902_ (
    .A(_395_),
    .B(_425_),
    .C(_428_),
    .Y(_498_)
);

FILL FILL_0__7688_ (
);

NAND2X1 _9794_ (
    .A(_3137_),
    .B(_3132_),
    .Y(_3138_)
);

FILL FILL_0__7268_ (
);

AOI21X1 _9374_ (
    .A(_2727_),
    .B(_2731_),
    .C(_2713_),
    .Y(_2732_)
);

FILL FILL_1__11202_ (
);

FILL FILL_2__8647_ (
);

FILL FILL_2__8227_ (
);

FILL FILL_0__10615_ (
);

NAND3X1 _10900_ (
    .A(_4038_),
    .B(_4096_),
    .C(_4100_),
    .Y(_4101_)
);

FILL FILL_0__13087_ (
);

DFFPOSX1 _13372_ (
    .D(\Y[6] [10]),
    .CLK(clk_bF$buf50),
    .Q(\u_fir_pe7.rYin [10])
);

FILL FILL_1__6644_ (
);

FILL FILL_2__13414_ (
);

FILL FILL_1__12827_ (
);

FILL FILL_1__12407_ (
);

FILL FILL_3__7931_ (
);

FILL FILL_0__9414_ (
);

FILL FILL_1__7849_ (
);

FILL FILL_1__7429_ (
);

FILL FILL_1__7009_ (
);

OAI21X1 _6499_ (
    .A(_98_),
    .B(_99_),
    .C(_97_),
    .Y(_100_)
);

FILL FILL_3__8716_ (
);

NAND2X1 _7860_ (
    .A(_1360_),
    .B(_1373_),
    .Y(_1374_)
);

NAND3X1 _7440_ (
    .A(vdd),
    .B(\X[1] [4]),
    .C(_950_),
    .Y(_960_)
);

NAND3X1 _7020_ (
    .A(_584_),
    .B(_612_),
    .C(_611_),
    .Y(_613_)
);

OR2X2 _10497_ (
    .A(_3769_),
    .B(_3767_),
    .Y(_3771_)
);

AOI21X1 _10077_ (
    .A(_3351_),
    .B(_3353_),
    .C(_3344_),
    .Y(_3357_)
);

FILL FILL_2__6713_ (
);

FILL FILL_1__12580_ (
);

FILL FILL_1__12160_ (
);

FILL FILL_2__10959_ (
);

FILL FILL_0__11993_ (
);

FILL FILL_2__10539_ (
);

FILL FILL_2__9185_ (
);

FILL FILL_0__11573_ (
);

FILL FILL_2__10119_ (
);

FILL FILL_0__11153_ (
);

FILL FILL_2__11900_ (
);

FILL FILL_0__6959_ (
);

FILL FILL_0__6539_ (
);

NAND3X1 _8645_ (
    .A(_2064_),
    .B(_2080_),
    .C(_2078_),
    .Y(_2081_)
);

AND2X2 _8225_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf1 ),
    .Y(_1666_)
);

FILL FILL_1__7182_ (
);

FILL FILL_0__7900_ (
);

FILL FILL_2__7918_ (
);

FILL FILL253650x54150 (
);

FILL FILL_0__12778_ (
);

NAND3X1 _12643_ (
    .A(_5681_),
    .B(_5683_),
    .C(_5682_),
    .Y(_5684_)
);

FILL FILL_0__12358_ (
);

NAND2X1 _12223_ (
    .A(_5336_),
    .B(_5337_),
    .Y(_5578_[11])
);

FILL FILL_1__8387_ (
);

FILL FILL_2__10292_ (
);

FILL FILL_3__9674_ (
);

INVX1 _13008_ (
    .A(_6043_),
    .Y(_6044_)
);

FILL FILL_2__7671_ (
);

FILL FILL_2__11497_ (
);

FILL FILL_2__11077_ (
);

AND2X2 _6711_ (
    .A(_307_),
    .B(_306_),
    .Y(_309_)
);

FILL FILL_0__7497_ (
);

FILL FILL_0__7077_ (
);

AND2X2 _9183_ (
    .A(_2538_),
    .B(_2542_),
    .Y(_2543_)
);

FILL FILL_3__10817_ (
);

FILL FILL_1__11851_ (
);

FILL FILL_1__11431_ (
);

FILL FILL_1__11011_ (
);

FILL FILL_2__8876_ (
);

FILL FILL_2__8456_ (
);

FILL FILL_0__10844_ (
);

FILL FILL_3__13289_ (
);

FILL FILL_0__10424_ (
);

FILL FILL_2__8036_ (
);

FILL FILL_0__10004_ (
);

AND2X2 _13181_ (
    .A(\u_fir_pe7.rYin [0]),
    .B(\u_fir_pe7.mul [0]),
    .Y(_6210_)
);

OAI21X1 _7916_ (
    .A(_1364_),
    .B(_1414_),
    .C(_1392_),
    .Y(_1427_)
);

FILL FILL_1__6873_ (
);

FILL FILL_1__6453_ (
);

FILL FILL_2__13223_ (
);

FILL FILL_3__6799_ (
);

FILL FILL_1__12636_ (
);

FILL FILL_1__12216_ (
);

FILL FILL_0__9643_ (
);

FILL FILL_0__9223_ (
);

OAI21X1 _11914_ (
    .A(_5032_),
    .B(_5027_),
    .C(_5021_),
    .Y(_5033_)
);

FILL FILL_3__7320_ (
);

FILL FILL_0__11209_ (
);

FILL FILL_3__10990_ (
);

FILL FILL_1__7658_ (
);

FILL FILL_3__10570_ (
);

FILL FILL_3__10150_ (
);

FILL FILL_3__8945_ (
);

FILL FILL_2__6942_ (
);

FILL FILL_3__11775_ (
);

FILL FILL_2__6522_ (
);

FILL FILL_3__11355_ (
);

FILL FILL_2__10768_ (
);

FILL FILL_2__10348_ (
);

FILL FILL_0__11382_ (
);

FILL FILL_1__9804_ (
);

FILL FILL_0__6768_ (
);

OAI21X1 _8874_ (
    .A(_2286_),
    .B(_2287_),
    .C(_2297_),
    .Y(_2298_)
);

INVX1 _8454_ (
    .A(_1876_),
    .Y(_1892_)
);

OAI21X1 _8034_ (
    .A(_1536_),
    .B(_1519_),
    .C(_1535_),
    .Y(_1538_)
);

FILL FILL_1__10702_ (
);

FILL FILL_2__7727_ (
);

FILL FILL_2__7307_ (
);

FILL FILL_1__13174_ (
);

AND2X2 _12872_ (
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5910_)
);

FILL FILL_0__12587_ (
);

FILL FILL_0__12167_ (
);

NAND3X1 _12452_ (
    .A(_5549_),
    .B(_5555_),
    .C(_5550_),
    .Y(_5556_)
);

AOI21X1 _12032_ (
    .A(_5060_),
    .B(_5059_),
    .C(_4991_),
    .Y(_5150_)
);

FILL FILL_2__12914_ (
);

NAND2X1 _9659_ (
    .A(_3009_),
    .B(_3008_),
    .Y(_3011_)
);

INVX1 _9239_ (
    .A(_2593_),
    .Y(_2598_)
);

FILL FILL_1__8196_ (
);

FILL FILL_1__11907_ (
);

FILL FILL_0__8914_ (
);

FILL FILL_3__9063_ (
);

INVX1 _13237_ (
    .A(\u_fir_pe7.rYin [7]),
    .Y(_6260_)
);

FILL FILL_1__6929_ (
);

FILL FILL_1__6509_ (
);

FILL FILL_2__7480_ (
);

FILL FILL_2__7060_ (
);

NAND3X1 _6940_ (
    .A(_529_),
    .B(_534_),
    .C(_533_),
    .Y(_535_)
);

INVX1 _6520_ (
    .A(_20_),
    .Y(_121_)
);

FILL FILL_1__10299_ (
);

FILL FILL_3__10626_ (
);

FILL FILL_1__11660_ (
);

FILL FILL_1__11240_ (
);

FILL FILL_2__8685_ (
);

FILL FILL_2__8265_ (
);

FILL FILL_0__10653_ (
);

FILL FILL_0__10233_ (
);

OAI21X1 _7725_ (
    .A(_1232_),
    .B(_1231_),
    .C(_1182_),
    .Y(_1242_)
);

NAND2X1 _7305_ (
    .A(\X[1] [0]),
    .B(vdd),
    .Y(_827_)
);

FILL FILL_1__6682_ (
);

FILL FILL_2__13032_ (
);

FILL FILL_1__12865_ (
);

FILL FILL_1__12445_ (
);

FILL FILL_1__12025_ (
);

FILL FILL_0__9452_ (
);

FILL FILL_0__11858_ (
);

FILL FILL_0__9032_ (
);

AOI21X1 _11723_ (
    .A(_4822_),
    .B(_4826_),
    .C(_4814_),
    .Y(_4845_)
);

FILL FILL_0__11438_ (
);

FILL FILL_0__11018_ (
);

NOR2X1 _11303_ (
    .A(_4478_),
    .B(_4483_),
    .Y(_4498_)
);

FILL FILL_1__7887_ (
);

FILL FILL_1__7467_ (
);

FILL FILL_1__7047_ (
);

NAND2X1 _12928_ (
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5965_)
);

FILL FILL_3__8334_ (
);

DFFPOSX1 _12508_ (
    .D(_5578_[7]),
    .CLK(clk_bF$buf29),
    .Q(\u_fir_pe6.mul [7])
);

FILL FILL_2__6751_ (
);

FILL FILL_2__10997_ (
);

FILL FILL_2__10577_ (
);

FILL FILL_2__10157_ (
);

FILL FILL_0__11191_ (
);

FILL FILL_1__9613_ (
);

FILL FILL_3__9959_ (
);

FILL FILL_3__9539_ (
);

FILL FILL_3__9119_ (
);

FILL FILL_0__6997_ (
);

FILL FILL_0__6577_ (
);

NAND2X1 _8683_ (
    .A(_2113_),
    .B(_2117_),
    .Y(_2118_)
);

OAI21X1 _8263_ (
    .A(_1702_),
    .B(_1703_),
    .C(_1701_),
    .Y(_1704_)
);

FILL FILL253950x248550 (
);

FILL FILL_1__10931_ (
);

FILL FILL_1__10511_ (
);

FILL FILL_2__7956_ (
);

FILL FILL_3__12789_ (
);

FILL FILL_2__7536_ (
);

FILL FILL_3__12369_ (
);

FILL FILL_2__7116_ (
);

AND2X2 _12681_ (
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_5721_)
);

FILL FILL_0__12396_ (
);

INVX1 _12261_ (
    .A(_5348_),
    .Y(_5374_)
);

FILL FILL_2__12723_ (
);

FILL FILL_2__12303_ (
);

INVX1 _9888_ (
    .A(_3888_),
    .Y(_3898_)
);

INVX1 _9468_ (
    .A(_2817_),
    .Y(_2825_)
);

NAND3X1 _9048_ (
    .A(_3173_),
    .B(_2405_),
    .C(_2408_),
    .Y(_2411_)
);

FILL FILL_1__11716_ (
);

FILL FILL_0__8723_ (
);

FILL FILL_0__8303_ (
);

FILL FILL_3__9292_ (
);

NAND2X1 _13046_ (
    .A(_6074_),
    .B(_6080_),
    .Y(_6082_)
);

FILL FILL_1__6738_ (
);

FILL FILL_0__9928_ (
);

FILL FILL_0__9508_ (
);

FILL FILL_3__10855_ (
);

FILL FILL_3__10015_ (
);

FILL FILL_2__8494_ (
);

FILL FILL_0__10882_ (
);

FILL FILL_0__10462_ (
);

FILL FILL_2__8074_ (
);

FILL FILL_0__10042_ (
);

OR2X2 _7954_ (
    .A(_1458_),
    .B(_1456_),
    .Y(_1460_)
);

OAI21X1 _7534_ (
    .A(_1045_),
    .B(_1052_),
    .C(_1037_),
    .Y(_1053_)
);

OAI21X1 _7114_ (
    .A(_681_),
    .B(_682_),
    .C(_696_),
    .Y(_697_)
);

FILL FILL_1__6491_ (
);

FILL FILL_2__13261_ (
);

FILL FILL_2__6807_ (
);

FILL FILL_1__12674_ (
);

FILL FILL_1__12254_ (
);

FILL FILL_0__9681_ (
);

FILL FILL_2__9699_ (
);

FILL FILL_2__9279_ (
);

FILL FILL_0__9261_ (
);

AND2X2 _11952_ (
    .A(_5067_),
    .B(_5070_),
    .Y(_5071_)
);

FILL FILL_0__11667_ (
);

AND2X2 _11532_ (
    .A(_4714_),
    .B(_4715_),
    .Y(_4775_[10])
);

FILL FILL_0__11247_ (
);

NAND2X1 _11112_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf3 ),
    .Y(_4310_)
);

FILL FILL254250x158550 (
);

AOI21X1 _8739_ (
    .A(_2171_),
    .B(_2172_),
    .C(_2155_),
    .Y(_2173_)
);

NAND3X1 _8319_ (
    .A(vdd),
    .B(\X[2] [3]),
    .C(_1758_),
    .Y(_1759_)
);

FILL FILL_1__7696_ (
);

FILL FILL_1__7276_ (
);

FILL FILL_1__13039_ (
);

FILL FILL_3__8563_ (
);

AOI21X1 _12737_ (
    .A(_5605_),
    .B(_5689_),
    .C(_5776_),
    .Y(_5777_)
);

OAI21X1 _12317_ (
    .A(_5423_),
    .B(_5424_),
    .C(_5422_),
    .Y(_5425_)
);

FILL FILL_2__6980_ (
);

FILL FILL_2__6560_ (
);

FILL FILL_2__10386_ (
);

FILL FILL_1__9422_ (
);

FILL FILL_3__9768_ (
);

FILL FILL_0__6386_ (
);

OAI21X1 _8492_ (
    .A(_1929_),
    .B(_1923_),
    .C(_1917_),
    .Y(_1930_)
);

AOI21X1 _8072_ (
    .A(\X[1] [0]),
    .B(gnd),
    .C(_1497_),
    .Y(_1574_)
);

FILL FILL_1__10320_ (
);

FILL FILL_2__7765_ (
);

FILL FILL_3__12598_ (
);

FILL FILL_2__7345_ (
);

DFFPOSX1 _12490_ (
    .D(\Y[7] [5]),
    .CLK(clk_bF$buf46),
    .Q(\u_fir_pe6.rYin [5])
);

AND2X2 _12070_ (
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5187_)
);

AOI22X1 _6805_ (
    .A(gnd),
    .B(Xin_5_bF$buf0),
    .C(vdd),
    .D(Xin[6]),
    .Y(_402_)
);

FILL FILL_2__12952_ (
);

FILL FILL_2__12532_ (
);

FILL FILL_2__12112_ (
);

NAND2X1 _9697_ (
    .A(_3043_),
    .B(_3038_),
    .Y(_3044_)
);

AOI21X1 _9277_ (
    .A(_2635_),
    .B(_2634_),
    .C(_2631_),
    .Y(_2636_)
);

FILL FILL_1__11945_ (
);

FILL FILL_1__11525_ (
);

FILL FILL_1__11105_ (
);

FILL FILL_0__8952_ (
);

FILL FILL_0__8532_ (
);

FILL FILL_0__10938_ (
);

FILL FILL_0__10518_ (
);

NAND3X1 _10803_ (
    .A(_4005_),
    .B(_4771_),
    .C(_4004_),
    .Y(_4006_)
);

AOI21X1 _13275_ (
    .A(_6293_),
    .B(_6271_),
    .C(_6291_),
    .Y(_6298_)
);

FILL FILL_2__9911_ (
);

FILL FILL_1__6967_ (
);

FILL FILL_1__6547_ (
);

FILL FILL_2__13317_ (
);

FILL FILL_0__9737_ (
);

FILL FILL_0__9317_ (
);

FILL FILL_3__7414_ (
);

FILL FILL_3__10244_ (
);

FILL FILL_0__10691_ (
);

FILL FILL_0__10271_ (
);

NAND3X1 _7763_ (
    .A(_1277_),
    .B(_1278_),
    .C(_1276_),
    .Y(_1279_)
);

NOR2X1 _7343_ (
    .A(_818_),
    .B(_855_),
    .Y(_864_)
);

FILL FILL_2__13070_ (
);

FILL FILL_3__11869_ (
);

FILL FILL_2__6616_ (
);

FILL FILL_3__11449_ (
);

FILL FILL_3__11029_ (
);

FILL FILL_1__12063_ (
);

FILL FILL_0__11896_ (
);

FILL FILL_0__9490_ (
);

FILL FILL_0__9070_ (
);

FILL FILL_2__9088_ (
);

OAI21X1 _11761_ (
    .A(_4880_),
    .B(_4881_),
    .C(_4879_),
    .Y(_4882_)
);

FILL FILL_0__11476_ (
);

FILL FILL_0__11056_ (
);

NAND3X1 _11341_ (
    .A(_4527_),
    .B(_4531_),
    .C(_4535_),
    .Y(_4536_)
);

FILL FILL_2__11803_ (
);

DFFPOSX1 _8968_ (
    .D(_2384_[15]),
    .CLK(clk_bF$buf4),
    .Q(\Y[3] [15])
);

OAI21X1 _8548_ (
    .A(_1984_),
    .B(_1983_),
    .C(_1980_),
    .Y(_1985_)
);

DFFPOSX1 _8128_ (
    .D(_1593_[12]),
    .CLK(clk_bF$buf13),
    .Q(\u_fir_pe1.mul [12])
);

FILL FILL_1__7085_ (
);

FILL FILL_0__7803_ (
);

FILL FILL_1__13268_ (
);

NAND2X1 _12966_ (
    .A(_5994_),
    .B(_6001_),
    .Y(_6003_)
);

INVX1 _12546_ (
    .A(_6319_),
    .Y(_5589_)
);

OAI21X1 _12126_ (
    .A(_5168_),
    .B(_5172_),
    .C(_5170_),
    .Y(_5242_)
);

FILL FILL_0__13202_ (
);

FILL FILL_2__10195_ (
);

FILL FILL_1__9651_ (
);

FILL FILL_1__9231_ (
);

FILL FILL_3__9157_ (
);

FILL FILL_2__7994_ (
);

FILL FILL_2__7574_ (
);

FILL FILL_2__7154_ (
);

INVX1 _6614_ (
    .A(_212_),
    .Y(_213_)
);

FILL FILL_2__12761_ (
);

FILL FILL_2__12341_ (
);

OR2X2 _9086_ (
    .A(_2447_),
    .B(_2446_),
    .Y(_2448_)
);

FILL FILL_1__11754_ (
);

FILL FILL_1__11334_ (
);

FILL FILL_0__8761_ (
);

FILL FILL_2__8779_ (
);

FILL FILL_0__8341_ (
);

FILL FILL_2__8359_ (
);

FILL FILL_0__10327_ (
);

NOR2X1 _10612_ (
    .A(_3872_),
    .B(_3871_),
    .Y(_3875_)
);

NAND2X1 _13084_ (
    .A(_6111_),
    .B(_6114_),
    .Y(_6119_)
);

FILL FILL_2__9720_ (
);

FILL FILL_2__9300_ (
);

NAND2X1 _7819_ (
    .A(_1333_),
    .B(_1313_),
    .Y(_1334_)
);

FILL FILL_1__6776_ (
);

FILL FILL_2__13126_ (
);

FILL FILL_1__12959_ (
);

FILL FILL_1__12539_ (
);

FILL FILL_1__12119_ (
);

FILL FILL_0__9966_ (
);

FILL FILL_0__9546_ (
);

FILL FILL_3__7643_ (
);

FILL FILL_0__9126_ (
);

OAI22X1 _11817_ (
    .A(_4824_),
    .B(_4935_),
    .C(_4867_),
    .D(_4936_),
    .Y(_4937_)
);

FILL FILL_3__10473_ (
);

FILL FILL_0__10080_ (
);

FILL FILL_1__8922_ (
);

FILL FILL_1__8502_ (
);

FILL FILL_3__8428_ (
);

FILL FILL_3__8008_ (
);

AND2X2 _7992_ (
    .A(_1474_),
    .B(_1484_),
    .Y(_1495_)
);

OAI21X1 _7572_ (
    .A(_1089_),
    .B(_1090_),
    .C(_1088_),
    .Y(_1091_)
);

NOR2X1 _7152_ (
    .A(_735_),
    .B(_732_),
    .Y(_736_)
);

FILL FILL_2__6845_ (
);

FILL FILL_2__6425_ (
);

FILL FILL_3__11258_ (
);

FILL FILL_1__12292_ (
);

NAND3X1 _11990_ (
    .A(vdd),
    .B(\X[7] [6]),
    .C(_5107_),
    .Y(_5108_)
);

NAND2X1 _11570_ (
    .A(_4749_),
    .B(_4743_),
    .Y(_4753_)
);

FILL FILL_0__11285_ (
);

AOI21X1 _11150_ (
    .A(_4342_),
    .B(_4347_),
    .C(_4286_),
    .Y(_4348_)
);

FILL FILL_1__9707_ (
);

AOI21X1 _8777_ (
    .A(_2151_),
    .B(_2153_),
    .C(_2208_),
    .Y(_2209_)
);

NAND2X1 _8357_ (
    .A(_1796_),
    .B(_1788_),
    .Y(_1797_)
);

FILL FILL_1__10605_ (
);

FILL FILL_0__7612_ (
);

FILL FILL_1__13077_ (
);

INVX1 _12775_ (
    .A(\X[6] [7]),
    .Y(_5814_)
);

FILL FILL_3__8181_ (
);

NOR2X1 _12355_ (
    .A(_5458_),
    .B(_5457_),
    .Y(_5459_)
);

FILL FILL_3__13404_ (
);

FILL FILL_2__12817_ (
);

FILL FILL_0__13011_ (
);

FILL FILL_0__8817_ (
);

FILL FILL_3__6914_ (
);

FILL FILL_1__9460_ (
);

FILL FILL_1__9040_ (
);

FILL FILL_3__9386_ (
);

FILL FILL_2__7383_ (
);

AOI21X1 _6843_ (
    .A(_430_),
    .B(_426_),
    .C(_385_),
    .Y(_440_)
);

NAND2X1 _6423_ (
    .A(Xin[4]),
    .B(gnd),
    .Y(_25_)
);

FILL FILL_2__12990_ (
);

FILL FILL_2__12570_ (
);

FILL FILL_2__12150_ (
);

FILL FILL_3__10949_ (
);

FILL FILL_1__11983_ (
);

FILL FILL_1__11563_ (
);

FILL FILL_3__10109_ (
);

FILL FILL_1__11143_ (
);

FILL FILL_0__8570_ (
);

FILL FILL_2__8588_ (
);

FILL FILL_0__10976_ (
);

FILL FILL_2__8168_ (
);

FILL FILL_0__8150_ (
);

FILL FILL_0__10556_ (
);

NAND2X1 _10841_ (
    .A(_4039_),
    .B(_4042_),
    .Y(_4043_)
);

OAI21X1 _10421_ (
    .A(_3696_),
    .B(_3564_),
    .C(_3646_),
    .Y(_3697_)
);

FILL FILL_0__10136_ (
);

NAND3X1 _10001_ (
    .A(gnd),
    .B(\X[4] [2]),
    .C(_3281_),
    .Y(_3282_)
);

NAND3X1 _7628_ (
    .A(_1139_),
    .B(_1140_),
    .C(_1141_),
    .Y(_1146_)
);

DFFPOSX1 _7208_ (
    .D(_790_[9]),
    .CLK(clk_bF$buf16),
    .Q(\Y[1] [9])
);

FILL FILL_1__6585_ (
);

FILL FILL_1__12768_ (
);

FILL FILL_1__12348_ (
);

FILL FILL_0__9775_ (
);

FILL FILL_3__7872_ (
);

FILL FILL_0__9355_ (
);

DFFPOSX1 _11626_ (
    .D(_4778_[2]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.mul [2])
);

FILL FILL_3__7032_ (
);

OAI21X1 _11206_ (
    .A(_4402_),
    .B(_4304_),
    .C(_4117_),
    .Y(_4403_)
);

FILL FILL_0__12702_ (
);

FILL FILL_1__8731_ (
);

FILL FILL_1__8311_ (
);

FILL FILL_3__8657_ (
);

NAND3X1 _7381_ (
    .A(_899_),
    .B(_901_),
    .C(_900_),
    .Y(_902_)
);

FILL FILL_2__6654_ (
);

FILL FILL_3__11067_ (
);

FILL FILL_0__11094_ (
);

FILL FILL_1__9936_ (
);

FILL FILL_1__9516_ (
);

FILL FILL_2__11841_ (
);

FILL FILL_2__11421_ (
);

FILL FILL_2__11001_ (
);

AOI21X1 _8586_ (
    .A(_2009_),
    .B(_2016_),
    .C(_1991_),
    .Y(_2023_)
);

INVX2 _8166_ (
    .A(\X[2] [3]),
    .Y(_1609_)
);

FILL FILL_1__10834_ (
);

FILL FILL_1__10414_ (
);

FILL FILL_2__7859_ (
);

FILL FILL_0__7841_ (
);

FILL FILL_0__7421_ (
);

FILL FILL_2__7439_ (
);

FILL FILL_2__7019_ (
);

FILL FILL_0__7001_ (
);

NAND2X1 _12584_ (
    .A(_5623_),
    .B(_5619_),
    .Y(_5626_)
);

FILL FILL_0__12299_ (
);

AOI21X1 _12164_ (
    .A(_5177_),
    .B(_5207_),
    .C(_5210_),
    .Y(_5280_)
);

FILL FILL_2__8800_ (
);

FILL FILL_3__13213_ (
);

FILL FILL_2__12626_ (
);

FILL FILL_2__12206_ (
);

FILL FILL_0__13240_ (
);

FILL FILL_0__8626_ (
);

FILL FILL_3__6723_ (
);

FILL FILL_0__8206_ (
);

DFFPOSX1 _13369_ (
    .D(\Y[6] [7]),
    .CLK(clk_bF$buf48),
    .Q(\u_fir_pe7.rYin [7])
);

FILL FILL_2__7192_ (
);

FILL FILL_3__7508_ (
);

OAI21X1 _6652_ (
    .A(_250_),
    .B(_245_),
    .C(_239_),
    .Y(_251_)
);

FILL FILL_1__11792_ (
);

FILL FILL_3__10338_ (
);

FILL FILL_1__11372_ (
);

FILL FILL_2__8397_ (
);

FILL FILL_0__10785_ (
);

NOR2X1 _10650_ (
    .A(_3912_),
    .B(_3913_),
    .Y(_3914_)
);

FILL FILL_0__10365_ (
);

OAI21X1 _10230_ (
    .A(_3203_),
    .B(_3507_),
    .C(_3213_),
    .Y(_3508_)
);

INVX1 _7857_ (
    .A(_1368_),
    .Y(_1371_)
);

AOI22X1 _7437_ (
    .A(vdd),
    .B(\X[1] [3]),
    .C(vdd),
    .D(\X[1] [4]),
    .Y(_957_)
);

OAI21X1 _7017_ (
    .A(_591_),
    .B(_586_),
    .C(_609_),
    .Y(_610_)
);

FILL FILL_1__6394_ (
);

FILL FILL_2__13164_ (
);

FILL FILL_1__12997_ (
);

FILL FILL_1__12577_ (
);

FILL FILL_1__12157_ (
);

FILL FILL_0__9584_ (
);

FILL FILL_0__9164_ (
);

AOI21X1 _11855_ (
    .A(_4974_),
    .B(_4973_),
    .C(_4972_),
    .Y(_4975_)
);

FILL FILL_3__7261_ (
);

NOR2X1 _11435_ (
    .A(_4616_),
    .B(_4621_),
    .Y(_4624_)
);

NAND2X1 _11015_ (
    .A(_4212_),
    .B(_4213_),
    .Y(_4214_)
);

FILL FILL_0__12931_ (
);

FILL FILL_1__7599_ (
);

FILL FILL_1__7179_ (
);

FILL FILL_3__10091_ (
);

FILL FILL_1__8540_ (
);

FILL FILL_3__8886_ (
);

NAND3X1 _7190_ (
    .A(_767_),
    .B(_773_),
    .C(_768_),
    .Y(_774_)
);

FILL FILL_2__6883_ (
);

FILL FILL_2__6463_ (
);

FILL FILL_3__11296_ (
);

FILL FILL_2__10289_ (
);

FILL FILL_1__9745_ (
);

FILL FILL_1__9325_ (
);

FILL FILL_2__11650_ (
);

FILL FILL_2__11230_ (
);

NAND2X1 _8395_ (
    .A(gnd),
    .B(\X[2] [6]),
    .Y(_1834_)
);

FILL FILL_1__10643_ (
);

FILL FILL_1__10223_ (
);

CLKBUF1 CLKBUF1_insert40 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert41 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert42 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert43 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert44 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf25)
);

FILL FILL_2__7668_ (
);

FILL FILL_0__7650_ (
);

CLKBUF1 CLKBUF1_insert45 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert46 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert47 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert48 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert49 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf20)
);

INVX1 _12393_ (
    .A(_5496_),
    .Y(_5497_)
);

NOR2X1 _6708_ (
    .A(_770_),
    .B(_305_),
    .Y(_306_)
);

FILL FILL_2__12855_ (
);

FILL FILL_2__12435_ (
);

FILL FILL_2__12015_ (
);

FILL FILL_1__11848_ (
);

FILL FILL_1__11428_ (
);

FILL FILL_1__11008_ (
);

FILL FILL_0__8855_ (
);

FILL FILL_3__6952_ (
);

FILL FILL_0__8435_ (
);

FILL FILL_3__6532_ (
);

NOR2X1 _10706_ (
    .A(_3967_),
    .B(_3974_),
    .Y(_3981_[2])
);

FILL FILL_0__8015_ (
);

OAI21X1 _13178_ (
    .A(_6146_),
    .B(_6196_),
    .C(_6174_),
    .Y(_6209_)
);

FILL FILL_2__9814_ (
);

FILL FILL_1__7811_ (
);

FILL FILL_3__7737_ (
);

AND2X2 _6881_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_477_)
);

AOI21X1 _6461_ (
    .A(_40_),
    .B(_44_),
    .C(_32_),
    .Y(_63_)
);

FILL FILL_3__10567_ (
);

FILL FILL_1__11181_ (
);

FILL FILL_0__10594_ (
);

FILL FILL_0__10174_ (
);

FILL FILL_2__10921_ (
);

FILL FILL_2__10501_ (
);

NAND2X1 _7666_ (
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_1183_)
);

DFFPOSX1 _7246_ (
    .D(_796_[7]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.mul [7])
);

FILL FILL_2__6939_ (
);

FILL FILL_0__6921_ (
);

FILL FILL_0__6501_ (
);

FILL FILL_2__6519_ (
);

FILL FILL_1__12386_ (
);

FILL FILL_0__9393_ (
);

FILL FILL_0__11799_ (
);

FILL FILL_3__7490_ (
);

INVX1 _11664_ (
    .A(_4786_),
    .Y(_4787_)
);

FILL FILL_0__11379_ (
);

FILL FILL_3__7070_ (
);

NAND2X1 _11244_ (
    .A(_4439_),
    .B(_4282_),
    .Y(_4440_)
);

FILL FILL_3__12713_ (
);

FILL FILL_2__11706_ (
);

FILL FILL_0__12740_ (
);

FILL FILL_0__12320_ (
);

FILL FILL_0__7706_ (
);

AND2X2 _9812_ (
    .A(_3149_),
    .B(_3155_),
    .Y(_3156_)
);

FILL FILL_3__8695_ (
);

OAI21X1 _12869_ (
    .A(_5668_),
    .B(_5723_),
    .C(_5906_),
    .Y(_5907_)
);

FILL FILL_3__8275_ (
);

OR2X2 _12449_ (
    .A(\u_fir_pe6.rYin [15]),
    .B(\u_fir_pe6.mul [15]),
    .Y(_5553_)
);

OAI21X1 _12029_ (
    .A(_5138_),
    .B(_5134_),
    .C(_5141_),
    .Y(_5147_)
);

FILL FILL253650x169350 (
);

FILL FILL_0__13105_ (
);

FILL FILL_2__6692_ (
);

FILL FILL_2__10098_ (
);

FILL FILL_1__9974_ (
);

FILL FILL_1__9554_ (
);

FILL FILL_1__9134_ (
);

FILL FILL_1__10872_ (
);

FILL FILL_1__10452_ (
);

FILL FILL_1__10032_ (
);

FILL FILL_2__7897_ (
);

FILL FILL_2__7477_ (
);

FILL FILL_2__7057_ (
);

OAI21X1 _6937_ (
    .A(_531_),
    .B(_530_),
    .C(_524_),
    .Y(_532_)
);

NAND3X1 _6517_ (
    .A(_26_),
    .B(_113_),
    .C(_114_),
    .Y(_118_)
);

FILL FILL_2__12664_ (
);

FILL FILL_2__12244_ (
);

FILL FILL_1__11657_ (
);

FILL FILL_1__11237_ (
);

FILL FILL_0__8664_ (
);

FILL FILL_0__8244_ (
);

NAND2X1 _10935_ (
    .A(_4134_),
    .B(_4126_),
    .Y(_4135_)
);

OR2X2 _10515_ (
    .A(_3760_),
    .B(_3786_),
    .Y(_3788_)
);

FILL FILL_2__9623_ (
);

FILL FILL_2__9203_ (
);

FILL FILL_1__6679_ (
);

FILL FILL_2__13029_ (
);

FILL FILL_1__7620_ (
);

FILL FILL_3__7966_ (
);

FILL FILL_0__9449_ (
);

FILL FILL_0__9029_ (
);

FILL FILL_3__7126_ (
);

AND2X2 _6690_ (
    .A(_285_),
    .B(_288_),
    .Y(_289_)
);

FILL FILL_3__10796_ (
);

FILL FILL_1__8825_ (
);

FILL FILL_1__8405_ (
);

FILL FILL_2__10310_ (
);

NAND2X1 _7895_ (
    .A(_1386_),
    .B(_1385_),
    .Y(_1408_)
);

AOI21X1 _7475_ (
    .A(_823_),
    .B(_907_),
    .C(_994_),
    .Y(_995_)
);

OAI21X1 _7055_ (
    .A(_641_),
    .B(_642_),
    .C(_640_),
    .Y(_643_)
);

FILL FILL_0__6730_ (
);

FILL FILL_2__6748_ (
);

FILL FILL_1__12195_ (
);

AOI22X1 _11893_ (
    .A(gnd),
    .B(\X[7] [7]),
    .C(\X[7] [3]),
    .D(gnd),
    .Y(_5012_)
);

OAI21X1 _11473_ (
    .A(_4650_),
    .B(_4651_),
    .C(_4655_),
    .Y(_4657_)
);

FILL FILL_0__11188_ (
);

NAND3X1 _11053_ (
    .A(_4223_),
    .B(_4242_),
    .C(_4236_),
    .Y(_4252_)
);

FILL FILL_3__12942_ (
);

FILL FILL_2__11935_ (
);

FILL FILL_2__11515_ (
);

FILL FILL_1__10928_ (
);

FILL FILL_1__10508_ (
);

FILL FILL_0__7935_ (
);

FILL FILL_0__7515_ (
);

OR2X2 _9621_ (
    .A(_2974_),
    .B(_2951_),
    .Y(_2975_)
);

AOI22X1 _9201_ (
    .A(vdd),
    .B(\X[3]_5_bF$buf2 ),
    .C(_2550_),
    .D(_2552_),
    .Y(_2561_)
);

NAND2X1 _12678_ (
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5718_)
);

NOR2X1 _12258_ (
    .A(_5371_),
    .B(_5370_),
    .Y(_5372_)
);

FILL FILL_3__13307_ (
);

FILL FILL_0__13334_ (
);

FILL FILL_1__9783_ (
);

FILL FILL_1__9363_ (
);

FILL FILL_1__10681_ (
);

FILL FILL_1__10261_ (
);

FILL FILL_2__7286_ (
);

FILL FILL_3__13060_ (
);

OAI21X1 _6746_ (
    .A(_335_),
    .B(_329_),
    .C(_337_),
    .Y(_344_)
);

FILL FILL_2__12893_ (
);

FILL FILL_2__12053_ (
);

FILL FILL_1__11886_ (
);

FILL FILL_1__11466_ (
);

FILL FILL_1__11046_ (
);

FILL FILL_0__8893_ (
);

FILL FILL_0__8473_ (
);

FILL FILL_0__10879_ (
);

FILL FILL_3__6570_ (
);

FILL FILL_0__10459_ (
);

DFFPOSX1 _10744_ (
    .D(\Y[4] [13]),
    .CLK(clk_bF$buf12),
    .Q(\u_fir_pe4.rYin [13])
);

FILL FILL_0__8053_ (
);

OAI21X1 _10324_ (
    .A(_3521_),
    .B(_3600_),
    .C(_3599_),
    .Y(_3601_)
);

FILL FILL_0__10039_ (
);

FILL FILL_2__9432_ (
);

FILL FILL_0__11820_ (
);

FILL FILL_2__9012_ (
);

FILL FILL_0__11400_ (
);

FILL FILL_1__6488_ (
);

FILL FILL_2__13258_ (
);

FILL FILL_0__9678_ (
);

FILL FILL_0__9258_ (
);

NAND3X1 _11949_ (
    .A(_5063_),
    .B(_5064_),
    .C(_5065_),
    .Y(_5068_)
);

FILL FILL_3__7355_ (
);

NOR2X1 _11529_ (
    .A(_4712_),
    .B(_4711_),
    .Y(_4713_)
);

OAI21X1 _11109_ (
    .A(_4303_),
    .B(_4306_),
    .C(_4305_),
    .Y(_4307_)
);

FILL FILL_0__12605_ (
);

FILL FILL_3__10185_ (
);

FILL FILL_1__8634_ (
);

FILL FILL_1__8214_ (
);

INVX1 _7284_ (
    .A(_1537_),
    .Y(_807_)
);

FILL FILL_3__9501_ (
);

FILL FILL_2__6977_ (
);

FILL FILL_2__6557_ (
);

NAND2X1 _11282_ (
    .A(_4476_),
    .B(_4472_),
    .Y(_4478_)
);

FILL FILL_1__9419_ (
);

FILL FILL_2__11744_ (
);

FILL FILL_2__11324_ (
);

NAND2X1 _8489_ (
    .A(gnd),
    .B(\X[2] [6]),
    .Y(_1927_)
);

NAND2X1 _8069_ (
    .A(_1571_),
    .B(_1572_),
    .Y(_1587_[15])
);

FILL FILL_1__10317_ (
);

FILL FILL_0__7744_ (
);

DFFPOSX1 _9850_ (
    .D(\X[3] [4]),
    .CLK(clk_bF$buf51),
    .Q(\X[4] [4])
);

FILL FILL_0__7324_ (
);

AOI21X1 _9430_ (
    .A(_2730_),
    .B(_2729_),
    .C(_2714_),
    .Y(_2787_)
);

AND2X2 _9010_ (
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_3091_)
);

DFFPOSX1 _12487_ (
    .D(\Y[7] [2]),
    .CLK(clk_bF$buf27),
    .Q(\u_fir_pe6.rYin [2])
);

AOI22X1 _12067_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf0 ),
    .C(vdd),
    .D(\X[7] [6]),
    .Y(_5184_)
);

FILL FILL_2__8703_ (
);

FILL FILL_2__12949_ (
);

FILL FILL_2__12529_ (
);

FILL FILL_2__12109_ (
);

FILL FILL_0__13143_ (
);

FILL FILL_1__6700_ (
);

FILL FILL_0__8949_ (
);

FILL FILL_0__8529_ (
);

FILL FILL_3__6626_ (
);

FILL FILL_1__9592_ (
);

FILL FILL_1__9172_ (
);

FILL FILL_3__9098_ (
);

FILL FILL_2__9908_ (
);

FILL FILL_1__10490_ (
);

FILL FILL_1__10070_ (
);

FILL FILL_2__7095_ (
);

FILL FILL_1__7905_ (
);

AOI21X1 _6975_ (
    .A(gnd),
    .B(_566_),
    .C(_568_),
    .Y(_569_)
);

OAI22X1 _6555_ (
    .A(_42_),
    .B(_153_),
    .C(_85_),
    .D(_154_),
    .Y(_155_)
);

FILL FILL_2__12282_ (
);

FILL FILL_1__11695_ (
);

FILL FILL_1__11275_ (
);

FILL FILL_0__8282_ (
);

FILL FILL_0__10688_ (
);

AOI22X1 _10973_ (
    .A(_4096_),
    .B(_4091_),
    .C(_4168_),
    .D(_4172_),
    .Y(_4173_)
);

NOR2X1 _10553_ (
    .A(_3820_),
    .B(_3821_),
    .Y(_3822_)
);

FILL FILL_0__10268_ (
);

OAI21X1 _10133_ (
    .A(_3361_),
    .B(_3411_),
    .C(_3355_),
    .Y(_3412_)
);

FILL FILL_2__9661_ (
);

FILL FILL_2__9241_ (
);

FILL FILL_2__13067_ (
);

NAND3X1 _8701_ (
    .A(_2109_),
    .B(_2135_),
    .C(_2131_),
    .Y(_2136_)
);

FILL FILL_0__9487_ (
);

FILL FILL_3__7584_ (
);

FILL FILL_0__9067_ (
);

INVX1 _11758_ (
    .A(_4866_),
    .Y(_4879_)
);

FILL FILL_3__7164_ (
);

NAND2X1 _11338_ (
    .A(_4532_),
    .B(_4499_),
    .Y(_4533_)
);

FILL FILL_3__12807_ (
);

FILL FILL_1__13001_ (
);

FILL FILL_0__12834_ (
);

FILL FILL_0__12414_ (
);

INVX1 _9906_ (
    .A(_3188_),
    .Y(_3189_)
);

FILL FILL_1__8863_ (
);

FILL FILL_1__8443_ (
);

FILL FILL_1__8023_ (
);

FILL FILL_3__8369_ (
);

NOR2X1 _7093_ (
    .A(_676_),
    .B(_675_),
    .Y(_677_)
);

FILL FILL_2__6786_ (
);

FILL FILL_3__11199_ (
);

FILL FILL254550x241350 (
);

NAND2X1 _11091_ (
    .A(\X[5] [1]),
    .B(gnd),
    .Y(_4289_)
);

FILL FILL_3__12980_ (
);

FILL FILL_1__9648_ (
);

FILL FILL_1__9228_ (
);

FILL FILL_3__12560_ (
);

FILL FILL_3__12140_ (
);

FILL FILL_2__11973_ (
);

FILL FILL_2__11553_ (
);

FILL FILL_2__11133_ (
);

INVX2 _8298_ (
    .A(\X[2] [6]),
    .Y(_1738_)
);

FILL FILL_1__10966_ (
);

FILL FILL_1__10546_ (
);

FILL FILL_1__10126_ (
);

FILL FILL_0__7973_ (
);

FILL FILL_0__7553_ (
);

FILL FILL_0__7133_ (
);

FILL FILL254550x208950 (
);

INVX1 _12296_ (
    .A(_5398_),
    .Y(_5408_)
);

FILL FILL_2__8932_ (
);

FILL FILL_2__8512_ (
);

FILL FILL_0__10900_ (
);

FILL FILL_2__12758_ (
);

FILL FILL_2__12338_ (
);

FILL FILL_0__8758_ (
);

FILL FILL_0__8338_ (
);

NOR2X1 _10609_ (
    .A(\u_fir_pe4.rYin [7]),
    .B(\u_fir_pe4.mul [7]),
    .Y(_3872_)
);

FILL FILL_2__9717_ (
);

FILL FILL_1__7714_ (
);

AOI21X1 _6784_ (
    .A(_361_),
    .B(_360_),
    .C(_303_),
    .Y(_381_)
);

FILL FILL_2__12091_ (
);

FILL FILL_1__11084_ (
);

FILL FILL_0__10497_ (
);

NAND2X1 _10782_ (
    .A(gnd),
    .B(\X[5] [2]),
    .Y(_3985_)
);

OR2X2 _10362_ (
    .A(_3568_),
    .B(_3638_),
    .Y(_3639_)
);

FILL FILL_0__10077_ (
);

FILL FILL_1__8919_ (
);

FILL FILL_3__11411_ (
);

FILL FILL_2__10824_ (
);

FILL FILL_2__9890_ (
);

FILL FILL_2__9470_ (
);

FILL FILL_2__10404_ (
);

FILL FILL_2__9050_ (
);

OAI21X1 _7989_ (
    .A(_1462_),
    .B(_1463_),
    .C(_1491_),
    .Y(_1492_)
);

NOR2X1 _7569_ (
    .A(_1004_),
    .B(_1001_),
    .Y(_1088_)
);

AND2X2 _7149_ (
    .A(\u_fir_pe0.rYin [11]),
    .B(\u_fir_pe0.mul [11]),
    .Y(_733_)
);

FILL FILL_2__13296_ (
);

FILL FILL_0__6824_ (
);

INVX1 _8930_ (
    .A(\u_fir_pe2.rYin [14]),
    .Y(_2353_)
);

FILL FILL_0__6404_ (
);

NAND3X1 _8510_ (
    .A(_1943_),
    .B(_1944_),
    .C(_1911_),
    .Y(_1948_)
);

FILL FILL_1__12289_ (
);

FILL FILL_0__9296_ (
);

OAI21X1 _11987_ (
    .A(_5022_),
    .B(_5030_),
    .C(_5029_),
    .Y(_5105_)
);

NOR2X1 _11567_ (
    .A(_4749_),
    .B(_4743_),
    .Y(_4751_)
);

NAND3X1 _11147_ (
    .A(_4338_),
    .B(_4339_),
    .C(_4340_),
    .Y(_4345_)
);

FILL FILL_1__13230_ (
);

FILL FILL_0__12643_ (
);

FILL FILL_0__12223_ (
);

FILL FILL_0__7609_ (
);

NOR2X1 _9715_ (
    .A(_3059_),
    .B(_3058_),
    .Y(_3060_)
);

FILL FILL_1__8672_ (
);

FILL FILL_1__8252_ (
);

FILL FILL_3__8598_ (
);

FILL FILL_0__13008_ (
);

FILL FILL_2__6595_ (
);

FILL FILL_1__9457_ (
);

FILL FILL_1__9037_ (
);

FILL FILL_2__11782_ (
);

FILL FILL_2__11362_ (
);

FILL FILL_1__10775_ (
);

FILL FILL_1__10355_ (
);

FILL FILL_0__7782_ (
);

FILL FILL_0__7362_ (
);

FILL FILL_2__8741_ (
);

FILL FILL_2__8321_ (
);

FILL FILL_3__13154_ (
);

FILL FILL_2__12987_ (
);

FILL FILL_2__12567_ (
);

FILL FILL_2__12147_ (
);

FILL FILL_0__13181_ (
);

FILL FILL_0__8567_ (
);

FILL FILL_3__6664_ (
);

FILL FILL_0__8147_ (
);

NAND2X1 _10838_ (
    .A(_3994_),
    .B(_3999_),
    .Y(_4040_)
);

INVX1 _10418_ (
    .A(_3693_),
    .Y(_3694_)
);

FILL FILL_1__12921_ (
);

FILL FILL_2__9946_ (
);

FILL FILL_2__9526_ (
);

FILL FILL_0__11914_ (
);

FILL FILL_2__9106_ (
);

FILL FILL_1__7943_ (
);

FILL FILL_1__7523_ (
);

FILL FILL_1__7103_ (
);

FILL FILL_3__7449_ (
);

AOI21X1 _6593_ (
    .A(_192_),
    .B(_191_),
    .C(_190_),
    .Y(_193_)
);

FILL FILL_3__8810_ (
);

FILL FILL_3__10279_ (
);

NOR2X1 _10591_ (
    .A(\u_fir_pe4.rYin [5]),
    .B(\u_fir_pe4.mul [5]),
    .Y(_3856_)
);

AOI21X1 _10171_ (
    .A(_3449_),
    .B(_3448_),
    .C(_3447_),
    .Y(_3450_)
);

FILL FILL_1__8728_ (
);

FILL FILL_3__11640_ (
);

FILL FILL_1__8308_ (
);

FILL FILL_2__10633_ (
);

FILL FILL_2__10213_ (
);

NAND2X1 _7798_ (
    .A(_1281_),
    .B(_1284_),
    .Y(_1313_)
);

NAND2X1 _7378_ (
    .A(_878_),
    .B(_874_),
    .Y(_899_)
);

FILL FILL_0__6633_ (
);

FILL FILL_1__12098_ (
);

OR2X2 _11796_ (
    .A(_4915_),
    .B(_4913_),
    .Y(_4916_)
);

NAND2X1 _11376_ (
    .A(_4567_),
    .B(_4569_),
    .Y(_4570_)
);

FILL FILL_2__11838_ (
);

FILL FILL_0__12872_ (
);

FILL FILL_2__11418_ (
);

FILL FILL_0__12452_ (
);

FILL FILL_0__12032_ (
);

FILL FILL_0__7838_ (
);

AOI22X1 _9944_ (
    .A(gnd),
    .B(\X[4] [1]),
    .C(gnd),
    .D(\X[4] [2]),
    .Y(_3226_)
);

FILL FILL_0__7418_ (
);

NAND2X1 _9524_ (
    .A(_2876_),
    .B(_2863_),
    .Y(_2880_)
);

INVX2 _9104_ (
    .A(\X[3]_5_bF$buf3 ),
    .Y(_2465_)
);

FILL FILL_1__8481_ (
);

FILL FILL_1__8061_ (
);

FILL FILL_0__13237_ (
);

NAND3X1 _13102_ (
    .A(_6033_),
    .B(_6135_),
    .C(_5876_),
    .Y(_6136_)
);

FILL FILL_1__9686_ (
);

FILL FILL_1__9266_ (
);

FILL FILL_2__11171_ (
);

FILL FILL_1__10584_ (
);

FILL FILL_1__10164_ (
);

FILL FILL_0__7591_ (
);

FILL FILL_2__7189_ (
);

FILL FILL_0__7171_ (
);

FILL FILL_3__10911_ (
);

FILL FILL_2__8550_ (
);

AOI22X1 _6649_ (
    .A(gnd),
    .B(Xin[4]),
    .C(vdd),
    .D(Xin_5_bF$buf2),
    .Y(_248_)
);

FILL FILL_2__12796_ (
);

FILL FILL_2__12376_ (
);

FILL FILL_1__11789_ (
);

FILL FILL_1__11369_ (
);

FILL FILL_0__8796_ (
);

FILL FILL_3__6893_ (
);

FILL FILL_0__8376_ (
);

FILL FILL_3__6473_ (
);

INVX1 _10647_ (
    .A(_3910_),
    .Y(_3911_)
);

OAI21X1 _10227_ (
    .A(_3426_),
    .B(_3504_),
    .C(_3448_),
    .Y(_3505_)
);

FILL FILL_1__12730_ (
);

FILL FILL_1__12310_ (
);

FILL FILL_2__9755_ (
);

FILL FILL_2__9335_ (
);

FILL FILL_0__11723_ (
);

FILL FILL_0__11303_ (
);

FILL FILL_1__7752_ (
);

FILL FILL_1__7332_ (
);

FILL FILL_3__7678_ (
);

FILL FILL_0__12928_ (
);

FILL FILL_1__8537_ (
);

FILL FILL_2__10862_ (
);

FILL FILL_2__10442_ (
);

FILL FILL_2__10022_ (
);

OR2X2 _7187_ (
    .A(\u_fir_pe0.rYin [15]),
    .B(\u_fir_pe0.mul [15]),
    .Y(_771_)
);

FILL FILL_3__9824_ (
);

FILL FILL_0__6862_ (
);

FILL FILL_0__6442_ (
);

OAI21X1 _11185_ (
    .A(_4307_),
    .B(_4381_),
    .C(_4328_),
    .Y(_4382_)
);

FILL FILL_2__7821_ (
);

FILL FILL_3__12654_ (
);

FILL FILL_2__7401_ (
);

FILL FILL_3__12234_ (
);

FILL FILL_2__11647_ (
);

FILL FILL_0__12681_ (
);

FILL FILL_2__11227_ (
);

FILL FILL_0__12261_ (
);

FILL FILL_0__7647_ (
);

INVX1 _9753_ (
    .A(_3094_),
    .Y(_3097_)
);

OAI21X1 _9333_ (
    .A(_2601_),
    .B(_2611_),
    .C(_2607_),
    .Y(_2691_)
);

FILL FILL_1__8290_ (
);

FILL FILL_2__8606_ (
);

FILL FILL_3__13019_ (
);

FILL FILL_0__13046_ (
);

NAND2X1 _13331_ (
    .A(_6353_),
    .B(_6354_),
    .Y(_6369_[15])
);

FILL FILL_1__6603_ (
);

FILL FILL_3__6949_ (
);

FILL FILL_1__9495_ (
);

FILL FILL_1__9075_ (
);

FILL FILL_1__10393_ (
);

FILL FILL_1__7808_ (
);

NOR2X1 _6878_ (
    .A(_473_),
    .B(_416_),
    .Y(_474_)
);

OR2X2 _6458_ (
    .A(_59_),
    .B(_58_),
    .Y(_60_)
);

FILL FILL_2__12185_ (
);

FILL FILL_1__11178_ (
);

FILL FILL_0__8185_ (
);

NAND3X1 _10876_ (
    .A(gnd),
    .B(\X[5] [3]),
    .C(_4068_),
    .Y(_4077_)
);

INVX1 _10456_ (
    .A(_3703_),
    .Y(_3731_)
);

INVX1 _10036_ (
    .A(_3313_),
    .Y(_3317_)
);

FILL FILL_3__11505_ (
);

FILL FILL_2__9984_ (
);

FILL FILL_2__10918_ (
);

FILL FILL_2__9564_ (
);

FILL FILL_0__11952_ (
);

FILL FILL_2__9144_ (
);

FILL FILL_0__11532_ (
);

FILL FILL_0__11112_ (
);

FILL FILL_0__6918_ (
);

AOI21X1 _8604_ (
    .A(_2040_),
    .B(_2039_),
    .C(_2032_),
    .Y(_2041_)
);

FILL FILL_1__7981_ (
);

FILL FILL_1__7561_ (
);

FILL FILL_1__7141_ (
);

FILL FILL_3__7067_ (
);

FILL FILL_1__13324_ (
);

FILL FILL_0__12737_ (
);

AOI21X1 _12602_ (
    .A(_5640_),
    .B(_5643_),
    .C(_5634_),
    .Y(_5644_)
);

FILL FILL_0__12317_ (
);

NOR2X1 _9809_ (
    .A(_3150_),
    .B(_3152_),
    .Y(_3153_)
);

FILL FILL_1__8766_ (
);

FILL FILL_1__8346_ (
);

FILL FILL_2__10671_ (
);

FILL FILL_2__10251_ (
);

FILL FILL_3__9633_ (
);

FILL FILL_3__9213_ (
);

FILL FILL_2__6689_ (
);

FILL FILL_0__6671_ (
);

FILL FILL_3__12883_ (
);

FILL FILL_2__7630_ (
);

FILL FILL_2__11876_ (
);

FILL FILL_2__11456_ (
);

FILL FILL_2__11036_ (
);

FILL FILL_0__12070_ (
);

FILL FILL_1__10869_ (
);

FILL FILL_1__10449_ (
);

FILL FILL_1__10029_ (
);

FILL FILL_0__7876_ (
);

NAND2X1 _9982_ (
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3263_)
);

FILL FILL_0__7456_ (
);

NAND2X1 _9562_ (
    .A(vdd),
    .B(\X[3] [7]),
    .Y(_2917_)
);

FILL FILL_0__7036_ (
);

INVX1 _9142_ (
    .A(_2417_),
    .Y(_2503_)
);

FILL FILL_1__11810_ (
);

OAI21X1 _12199_ (
    .A(_5313_),
    .B(_5312_),
    .C(_5306_),
    .Y(_5314_)
);

FILL FILL_2__8835_ (
);

FILL FILL_2__8415_ (
);

FILL FILL_0__10803_ (
);

FILL FILL_3__13248_ (
);

FILL FILL_0__13275_ (
);

INVX1 _13140_ (
    .A(_6172_),
    .Y(_6173_)
);

FILL FILL_1__6832_ (
);

FILL FILL_1__6412_ (
);

FILL FILL_0__9602_ (
);

FILL FILL_1__7617_ (
);

NAND3X1 _6687_ (
    .A(_281_),
    .B(_282_),
    .C(_283_),
    .Y(_286_)
);

FILL FILL_3__8904_ (
);

INVX1 _10685_ (
    .A(\u_fir_pe4.mul [14]),
    .Y(_3949_)
);

OAI21X1 _10265_ (
    .A(_3529_),
    .B(_3533_),
    .C(_3536_),
    .Y(_3543_)
);

FILL FILL_2__6901_ (
);

FILL FILL_3__11734_ (
);

FILL FILL_2__9793_ (
);

FILL FILL_2__9373_ (
);

FILL FILL_0__11761_ (
);

FILL FILL_2__10307_ (
);

FILL FILL_0__11341_ (
);

FILL FILL_2__13199_ (
);

FILL FILL_0__6727_ (
);

OAI21X1 _8833_ (
    .A(_2249_),
    .B(_2250_),
    .C(_2256_),
    .Y(_2258_)
);

AOI21X1 _8413_ (
    .A(_1845_),
    .B(_1851_),
    .C(_1832_),
    .Y(_1852_)
);

FILL FILL_1__7790_ (
);

FILL FILL_1__7370_ (
);

FILL FILL_0__9199_ (
);

FILL FILL_3__7296_ (
);

FILL FILL_3__12519_ (
);

FILL FILL_1__13133_ (
);

FILL FILL_0__12966_ (
);

NOR2X1 _12831_ (
    .A(_5786_),
    .B(_5783_),
    .Y(_5870_)
);

FILL FILL_0__12546_ (
);

FILL FILL_0__12126_ (
);

AND2X2 _12411_ (
    .A(\u_fir_pe6.rYin [11]),
    .B(\u_fir_pe6.mul [11]),
    .Y(_5515_)
);

INVX1 _9618_ (
    .A(_2971_),
    .Y(_2972_)
);

FILL FILL_1__8575_ (
);

FILL FILL_1__8155_ (
);

FILL FILL_2__10480_ (
);

FILL FILL_2__10060_ (
);

FILL FILL_3__9442_ (
);

FILL FILL_0__6480_ (
);

FILL FILL_2__6498_ (
);

FILL FILL_2__11685_ (
);

FILL FILL_2__11265_ (
);

FILL FILL_1__10678_ (
);

FILL FILL_1__10258_ (
);

FILL FILL_0__7685_ (
);

NOR2X1 _9791_ (
    .A(_3133_),
    .B(_3134_),
    .Y(_3135_)
);

FILL FILL_0__7265_ (
);

NAND3X1 _9371_ (
    .A(_2721_),
    .B(_2725_),
    .C(_2723_),
    .Y(_2729_)
);

FILL FILL_2__8644_ (
);

FILL FILL_2__8224_ (
);

FILL FILL_0__10612_ (
);

FILL FILL_0__13084_ (
);

FILL FILL_1__6641_ (
);

FILL FILL_2__13411_ (
);

FILL FILL_3__6987_ (
);

FILL FILL_3__6567_ (
);

FILL FILL_1__12824_ (
);

FILL FILL_1__12404_ (
);

FILL FILL_2__9429_ (
);

FILL FILL_0__9411_ (
);

FILL FILL_0__11817_ (
);

FILL FILL_2__9009_ (
);

FILL FILL_1__7846_ (
);

FILL FILL_1__7426_ (
);

FILL FILL_1__7006_ (
);

INVX1 _6496_ (
    .A(_84_),
    .Y(_97_)
);

NAND3X1 _10494_ (
    .A(_3749_),
    .B(_3766_),
    .C(_3765_),
    .Y(_3768_)
);

NAND3X1 _10074_ (
    .A(_3344_),
    .B(_3351_),
    .C(_3353_),
    .Y(_3354_)
);

FILL FILL_3__11963_ (
);

FILL FILL_2__6710_ (
);

FILL FILL_3__11123_ (
);

FILL FILL_2__10956_ (
);

FILL FILL_0__11990_ (
);

FILL FILL_2__10536_ (
);

FILL FILL_2__9182_ (
);

FILL FILL_0__11570_ (
);

FILL FILL_2__10116_ (
);

FILL FILL_0__11150_ (
);

FILL FILL_3__9918_ (
);

FILL FILL_0__6956_ (
);

FILL FILL_0__6536_ (
);

NAND2X1 _8642_ (
    .A(_2077_),
    .B(_2066_),
    .Y(_2078_)
);

OAI21X1 _8222_ (
    .A(_1623_),
    .B(_1657_),
    .C(_1639_),
    .Y(_1663_)
);

INVX1 _11699_ (
    .A(_4820_),
    .Y(_4821_)
);

NAND3X1 _11279_ (
    .A(_4392_),
    .B(_4468_),
    .C(_4400_),
    .Y(_4475_)
);

FILL FILL_2__7915_ (
);

FILL FILL_3__12748_ (
);

FILL FILL_3__12328_ (
);

FILL FILL_0__12775_ (
);

NAND2X1 _12640_ (
    .A(_5660_),
    .B(_5656_),
    .Y(_5681_)
);

FILL FILL_0__12355_ (
);

INVX1 _12220_ (
    .A(_5334_),
    .Y(_5335_)
);

DFFPOSX1 _9847_ (
    .D(\X[3] [1]),
    .CLK(clk_bF$buf28),
    .Q(\X[4] [1])
);

INVX1 _9427_ (
    .A(_2781_),
    .Y(_2784_)
);

DFFPOSX1 _9007_ (
    .D(_2390_[14]),
    .CLK(clk_bF$buf42),
    .Q(\u_fir_pe2.mul [14])
);

FILL FILL_1__8384_ (
);

INVX2 _13005_ (
    .A(gnd),
    .Y(_6041_)
);

FILL FILL_1__9589_ (
);

FILL FILL_1__9169_ (
);

FILL FILL_3__12081_ (
);

FILL FILL_2__11494_ (
);

FILL FILL_2__11074_ (
);

FILL FILL_1__10487_ (
);

FILL FILL_1__10067_ (
);

FILL FILL_0__7494_ (
);

FILL FILL_0__7074_ (
);

NAND2X1 _9180_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2540_)
);

FILL FILL_2__8873_ (
);

FILL FILL_2__8453_ (
);

FILL FILL_0__10841_ (
);

FILL FILL_0__10421_ (
);

FILL FILL_2__8033_ (
);

FILL FILL_0__10001_ (
);

FILL FILL_2__12699_ (
);

FILL FILL_2__12279_ (
);

NAND3X1 _7913_ (
    .A(_1423_),
    .B(_1424_),
    .C(_1422_),
    .Y(_1425_)
);

FILL FILL_1__6870_ (
);

FILL FILL_1__6450_ (
);

FILL FILL_0__8699_ (
);

FILL FILL_2__13220_ (
);

FILL FILL_0__8279_ (
);

FILL FILL_1__12633_ (
);

FILL FILL_1__12213_ (
);

FILL FILL_0__9640_ (
);

FILL FILL_2__9658_ (
);

FILL FILL_0__9220_ (
);

AOI22X1 _11911_ (
    .A(gnd),
    .B(\X[7] [4]),
    .C(vdd),
    .D(\X[7]_5_bF$buf3 ),
    .Y(_5030_)
);

FILL FILL_2__9238_ (
);

FILL FILL_0__11206_ (
);

FILL FILL253650x75750 (
);

FILL FILL_1__7655_ (
);

FILL FILL_3__8522_ (
);

FILL FILL_3__11352_ (
);

FILL FILL_2__10765_ (
);

FILL FILL_2__10345_ (
);

FILL FILL_1__9801_ (
);

FILL FILL_3__9307_ (
);

FILL FILL_0__6765_ (
);

AND2X2 _8871_ (
    .A(_2253_),
    .B(_2263_),
    .Y(_2295_)
);

NAND3X1 _8451_ (
    .A(_1879_),
    .B(_1882_),
    .C(_1798_),
    .Y(_1889_)
);

NOR2X1 _8031_ (
    .A(_1533_),
    .B(_1534_),
    .Y(_1587_[11])
);

INVX1 _11088_ (
    .A(_4285_),
    .Y(_4286_)
);

FILL FILL_3__12977_ (
);

FILL FILL_2__7724_ (
);

FILL FILL_2__7304_ (
);

FILL FILL_3__12137_ (
);

FILL FILL_1__13171_ (
);

FILL FILL_0__12584_ (
);

FILL FILL_0__12164_ (
);

FILL FILL_2__12911_ (
);

OAI21X1 _9656_ (
    .A(_2985_),
    .B(_2992_),
    .C(_2991_),
    .Y(_3008_)
);

OAI21X1 _9236_ (
    .A(_2520_),
    .B(_2518_),
    .C(_2511_),
    .Y(_2596_)
);

FILL FILL_1__8193_ (
);

FILL FILL_1__11904_ (
);

FILL FILL_2__8929_ (
);

FILL FILL_0__8911_ (
);

FILL FILL_2__8509_ (
);

FILL FILL_3__9480_ (
);

FILL FILL_3__9060_ (
);

OR2X2 _13234_ (
    .A(_6251_),
    .B(_6256_),
    .Y(_6258_)
);

FILL FILL_1__6926_ (
);

FILL FILL_1__6506_ (
);

FILL FILL_1__9398_ (
);

FILL FILL_1__10296_ (
);

FILL FILL_3__10203_ (
);

FILL FILL_2__8682_ (
);

FILL FILL_2__8262_ (
);

FILL FILL_0__10650_ (
);

FILL FILL_3__13095_ (
);

FILL FILL_0__10230_ (
);

FILL FILL_2__12088_ (
);

NAND3X1 _7722_ (
    .A(_1179_),
    .B(_1234_),
    .C(_1238_),
    .Y(_1239_)
);

AOI22X1 _7302_ (
    .A(\X[1] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[1] [4]),
    .Y(_824_)
);

INVX1 _10779_ (
    .A(_4770_),
    .Y(_4771_)
);

AOI21X1 _10359_ (
    .A(_3624_),
    .B(_3619_),
    .C(_3571_),
    .Y(_3636_)
);

FILL FILL_3__11828_ (
);

FILL FILL_1__12862_ (
);

FILL FILL_1__12442_ (
);

FILL FILL_1__12022_ (
);

FILL FILL_2__9887_ (
);

FILL FILL_2__9467_ (
);

FILL FILL_0__11855_ (
);

FILL FILL_2__9047_ (
);

OR2X2 _11720_ (
    .A(_4841_),
    .B(_4840_),
    .Y(_4842_)
);

FILL FILL_0__11435_ (
);

NOR2X1 _11300_ (
    .A(_4492_),
    .B(_4495_),
    .Y(_4781_[10])
);

FILL FILL_0__11015_ (
);

OR2X2 _8927_ (
    .A(_2343_),
    .B(_2349_),
    .Y(_2351_)
);

NAND3X1 _8507_ (
    .A(_1943_),
    .B(_1944_),
    .C(_1942_),
    .Y(_1945_)
);

FILL FILL_1__7884_ (
);

FILL FILL_1__7464_ (
);

FILL FILL_1__7044_ (
);

FILL FILL_1__13227_ (
);

FILL FILL_3__8751_ (
);

OAI21X1 _12925_ (
    .A(_5883_),
    .B(_5887_),
    .C(_5892_),
    .Y(_5962_)
);

DFFPOSX1 _12505_ (
    .D(_5577_[4]),
    .CLK(clk_bF$buf8),
    .Q(\u_fir_pe6.mul [4])
);

FILL FILL_1__8669_ (
);

FILL FILL_1__8249_ (
);

FILL FILL_2__10994_ (
);

FILL FILL_2__10574_ (
);

FILL FILL_2__10154_ (
);

FILL FILL_1__9610_ (
);

FILL FILL_3__9536_ (
);

FILL FILL_0__6994_ (
);

FILL FILL_0__6574_ (
);

NAND2X1 _8680_ (
    .A(gnd),
    .B(_2068_),
    .Y(_2115_)
);

AOI21X1 _8260_ (
    .A(_1622_),
    .B(_1642_),
    .C(_1656_),
    .Y(_1701_)
);

FILL FILL_2__7953_ (
);

FILL FILL_2__7533_ (
);

FILL FILL_2__7113_ (
);

FILL FILL_2__11779_ (
);

FILL FILL_2__11359_ (
);

FILL FILL_0__12393_ (
);

FILL FILL_2__12720_ (
);

FILL FILL_2__12300_ (
);

FILL FILL_0__7779_ (
);

DFFPOSX1 _9885_ (
    .D(_3187_[15]),
    .CLK(clk_bF$buf4),
    .Q(\u_fir_pe3.mul [15])
);

FILL FILL_0__7359_ (
);

NAND3X1 _9465_ (
    .A(_2817_),
    .B(_2821_),
    .C(_2776_),
    .Y(_2822_)
);

OAI21X1 _9045_ (
    .A(_3169_),
    .B(_2406_),
    .C(_2407_),
    .Y(_2408_)
);

FILL FILL_1__11713_ (
);

FILL FILL_2__8738_ (
);

FILL FILL_0__8720_ (
);

FILL FILL_2__8318_ (
);

FILL FILL_0__8300_ (
);

FILL FILL_0__10706_ (
);

FILL FILL_0__13178_ (
);

NAND2X1 _13043_ (
    .A(_6077_),
    .B(_6078_),
    .Y(_6079_)
);

FILL FILL_1__6735_ (
);

FILL FILL_1__12918_ (
);

FILL FILL_0__9925_ (
);

FILL FILL_0__9505_ (
);

FILL FILL_3__7602_ (
);

FILL FILL_3__10852_ (
);

FILL FILL_3__10432_ (
);

FILL FILL_2__8491_ (
);

FILL FILL_2__8071_ (
);

INVX1 _7951_ (
    .A(_1447_),
    .Y(_1457_)
);

NAND3X1 _7531_ (
    .A(_1043_),
    .B(_1046_),
    .C(_1044_),
    .Y(_1050_)
);

NAND2X1 _7111_ (
    .A(_657_),
    .B(_669_),
    .Y(_694_)
);

INVX1 _10588_ (
    .A(\u_fir_pe4.rYin [5]),
    .Y(_3853_)
);

AND2X2 _10168_ (
    .A(_3425_),
    .B(_3420_),
    .Y(_3447_)
);

FILL FILL_2__6804_ (
);

FILL FILL_1__12671_ (
);

FILL FILL_3__11217_ (
);

FILL FILL_1__12251_ (
);

FILL FILL_2__9696_ (
);

FILL FILL_2__9276_ (
);

FILL FILL_0__11664_ (
);

FILL FILL_0__11244_ (
);

NAND2X1 _8736_ (
    .A(_2166_),
    .B(_2169_),
    .Y(_2170_)
);

NAND3X1 _8316_ (
    .A(_1751_),
    .B(_1755_),
    .C(_1753_),
    .Y(_1756_)
);

FILL FILL_1__7693_ (
);

FILL FILL_1__7273_ (
);

FILL FILL_1__13036_ (
);

FILL FILL_0__12869_ (
);

AOI21X1 _12734_ (
    .A(_5697_),
    .B(_5696_),
    .C(_5633_),
    .Y(_5774_)
);

FILL FILL_3__8140_ (
);

FILL FILL_0__12449_ (
);

FILL FILL_0__12029_ (
);

OAI21X1 _12314_ (
    .A(_5414_),
    .B(_5415_),
    .C(_5419_),
    .Y(_5422_)
);

FILL FILL_1__8898_ (
);

FILL FILL_1__8478_ (
);

FILL FILL_1__8058_ (
);

FILL FILL_3__11390_ (
);

FILL FILL_2__10383_ (
);

FILL FILL_3__9765_ (
);

FILL FILL_0__6383_ (
);

FILL FILL_2__7762_ (
);

FILL FILL_3__12595_ (
);

FILL FILL_2__7342_ (
);

FILL FILL_3__12175_ (
);

FILL FILL_2__11168_ (
);

AND2X2 _6802_ (
    .A(_132_),
    .B(_321_),
    .Y(_399_)
);

FILL FILL_0__7588_ (
);

NOR2X1 _9694_ (
    .A(_3039_),
    .B(_3040_),
    .Y(_3041_)
);

FILL FILL_0__7168_ (
);

AND2X2 _9274_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf2 ),
    .Y(_2633_)
);

FILL FILL_1__11942_ (
);

FILL FILL_1__11522_ (
);

FILL FILL_1__11102_ (
);

FILL FILL_2__8547_ (
);

FILL FILL_0__10935_ (
);

FILL FILL_0__10515_ (
);

NAND2X1 _10800_ (
    .A(_3999_),
    .B(_4002_),
    .Y(_4003_)
);

OAI21X1 _13272_ (
    .A(_6291_),
    .B(_6292_),
    .C(_6290_),
    .Y(_6296_)
);

FILL FILL_1__6964_ (
);

FILL FILL_1__6544_ (
);

FILL FILL_2__13314_ (
);

FILL FILL_1__12727_ (
);

FILL FILL_1__12307_ (
);

FILL FILL_0__9734_ (
);

FILL FILL_3__7831_ (
);

FILL FILL_0__9314_ (
);

FILL FILL_3__7411_ (
);

FILL FILL_1__7749_ (
);

FILL FILL_3__10661_ (
);

FILL FILL_1__7329_ (
);

NAND2X1 _6399_ (
    .A(gnd),
    .B(Xin[0]),
    .Y(_2_)
);

FILL FILL_3__8616_ (
);

NAND2X1 _7760_ (
    .A(_1274_),
    .B(_1275_),
    .Y(_1276_)
);

AOI21X1 _7340_ (
    .A(_858_),
    .B(_861_),
    .C(_852_),
    .Y(_862_)
);

NAND2X1 _10397_ (
    .A(_3670_),
    .B(_3664_),
    .Y(_3673_)
);

FILL FILL_2__6613_ (
);

FILL FILL_3__11446_ (
);

FILL FILL_1__12060_ (
);

FILL FILL_2__10859_ (
);

FILL FILL_0__11893_ (
);

FILL FILL_2__10439_ (
);

FILL FILL_2__9085_ (
);

FILL FILL_0__11473_ (
);

FILL FILL_2__10019_ (
);

FILL FILL_0__11053_ (
);

FILL FILL_2__11800_ (
);

FILL FILL_0__6859_ (
);

DFFPOSX1 _8965_ (
    .D(_2384_[12]),
    .CLK(clk_bF$buf55),
    .Q(\Y[3] [12])
);

FILL FILL_0__6439_ (
);

NAND2X1 _8545_ (
    .A(gnd),
    .B(_1981_),
    .Y(_1982_)
);

DFFPOSX1 _8125_ (
    .D(_1593_[9]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.mul [9])
);

FILL FILL_1__7082_ (
);

FILL FILL_2__7818_ (
);

FILL FILL_0__7800_ (
);

FILL FILL_1__13265_ (
);

FILL FILL_0__12678_ (
);

NAND2X1 _12963_ (
    .A(_5985_),
    .B(_5988_),
    .Y(_6000_)
);

FILL FILL_0__12258_ (
);

NOR2X1 _12543_ (
    .A(_6310_),
    .B(_5581_),
    .Y(_5586_)
);

AOI21X1 _12123_ (
    .A(_5154_),
    .B(_5224_),
    .C(_5238_),
    .Y(_5239_)
);

FILL FILL_1__8287_ (
);

FILL FILL_2__10192_ (
);

FILL FILL_3__9994_ (
);

FILL FILL_3__9574_ (
);

FILL FILL_3__9154_ (
);

INVX1 _13328_ (
    .A(_6351_),
    .Y(_6352_)
);

FILL FILL_2__7991_ (
);

FILL FILL_2__7571_ (
);

FILL FILL_2__7151_ (
);

FILL FILL_2__11397_ (
);

NAND2X1 _6611_ (
    .A(Xin[0]),
    .B(gnd),
    .Y(_210_)
);

FILL FILL_0__7397_ (
);

INVX1 _9083_ (
    .A(_2444_),
    .Y(_2445_)
);

FILL FILL_1__11751_ (
);

FILL FILL_1__11331_ (
);

FILL FILL_2__8776_ (
);

FILL FILL_2__8356_ (
);

FILL FILL_3__13189_ (
);

FILL FILL_0__10324_ (
);

NAND2X1 _13081_ (
    .A(_6115_),
    .B(_6095_),
    .Y(_6116_)
);

INVX1 _7816_ (
    .A(_1328_),
    .Y(_1331_)
);

FILL FILL_1__6773_ (
);

FILL FILL_2__13123_ (
);

FILL FILL_3__6699_ (
);

FILL FILL_1__12956_ (
);

FILL FILL_1__12536_ (
);

FILL FILL_1__12116_ (
);

FILL FILL_0__9963_ (
);

FILL FILL_0__9543_ (
);

FILL FILL_0__11949_ (
);

FILL FILL_0__9123_ (
);

AND2X2 _11814_ (
    .A(_4929_),
    .B(_4933_),
    .Y(_4934_)
);

FILL FILL_0__11529_ (
);

FILL FILL_0__11109_ (
);

FILL FILL_1__7978_ (
);

FILL FILL_3__10890_ (
);

FILL FILL_1__7558_ (
);

FILL FILL_1__7138_ (
);

FILL FILL_3__10050_ (
);

FILL FILL_3__8845_ (
);

FILL FILL_3__8005_ (
);

FILL FILL_2__6842_ (
);

FILL FILL_3__11675_ (
);

FILL FILL_2__6422_ (
);

FILL FILL_2__10668_ (
);

FILL FILL_2__10248_ (
);

FILL FILL_0__11282_ (
);

FILL FILL_1__9704_ (
);

FILL FILL_0__6668_ (
);

NAND3X1 _8774_ (
    .A(_2178_),
    .B(_2206_),
    .C(_2205_),
    .Y(_2207_)
);

AOI21X1 _8354_ (
    .A(_1776_),
    .B(_1771_),
    .C(_1778_),
    .Y(_1794_)
);

FILL FILL_1__10602_ (
);

FILL FILL_2__7627_ (
);

FILL FILL_1__13074_ (
);

NAND3X1 _12772_ (
    .A(_5805_),
    .B(_5810_),
    .C(_5808_),
    .Y(_5811_)
);

FILL FILL_0__12067_ (
);

INVX1 _12352_ (
    .A(\u_fir_pe6.mul [6]),
    .Y(_5456_)
);

FILL FILL_2__12814_ (
);

AND2X2 _9979_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf1 ),
    .Y(_3260_)
);

NAND3X1 _9559_ (
    .A(_2911_),
    .B(_2912_),
    .C(_2913_),
    .Y(_2914_)
);

AOI21X1 _9139_ (
    .A(_2491_),
    .B(_2487_),
    .C(_2473_),
    .Y(_2500_)
);

FILL FILL_1__11807_ (
);

FILL FILL_0__8814_ (
);

FILL FILL_3__9383_ (
);

NOR2X1 _13137_ (
    .A(_6139_),
    .B(_6162_),
    .Y(_6170_)
);

FILL FILL_1__6829_ (
);

FILL FILL_1__6409_ (
);

FILL FILL_2__7380_ (
);

NAND3X1 _6840_ (
    .A(_383_),
    .B(_431_),
    .C(_436_),
    .Y(_437_)
);

AOI21X1 _6420_ (
    .A(_19_),
    .B(_20_),
    .C(_786_),
    .Y(_23_)
);

FILL FILL_1__10199_ (
);

FILL FILL_3__10946_ (
);

FILL FILL_1__11980_ (
);

FILL FILL_3__10526_ (
);

FILL FILL_1__11560_ (
);

FILL FILL_1__11140_ (
);

FILL FILL_2__8585_ (
);

FILL FILL_0__10973_ (
);

FILL FILL_2__8165_ (
);

FILL FILL_0__10553_ (
);

FILL FILL_0__10133_ (
);

OAI21X1 _7625_ (
    .A(_1138_),
    .B(_1142_),
    .C(_1114_),
    .Y(_1143_)
);

DFFPOSX1 _7205_ (
    .D(_790_[6]),
    .CLK(clk_bF$buf16),
    .Q(\Y[1] [6])
);

FILL FILL_1__6582_ (
);

FILL FILL_1__12765_ (
);

FILL FILL_1__12345_ (
);

FILL FILL_0__9772_ (
);

FILL FILL_0__9352_ (
);

FILL FILL_0__11758_ (
);

DFFPOSX1 _11623_ (
    .D(\Y[5] [15]),
    .CLK(clk_bF$buf50),
    .Q(\u_fir_pe5.rYin [15])
);

FILL FILL_0__11338_ (
);

NAND3X1 _11203_ (
    .A(_4385_),
    .B(_4392_),
    .C(_4399_),
    .Y(_4400_)
);

FILL FILL_1__7787_ (
);

FILL FILL_1__7367_ (
);

NAND3X1 _12828_ (
    .A(_5767_),
    .B(_5865_),
    .C(_5866_),
    .Y(_5867_)
);

FILL FILL_3__8234_ (
);

OAI21X1 _12408_ (
    .A(_5508_),
    .B(_5509_),
    .C(_5504_),
    .Y(_5512_)
);

FILL FILL_2__6651_ (
);

FILL FILL_3__11064_ (
);

FILL FILL_2__10897_ (
);

FILL FILL_2__10477_ (
);

FILL FILL_2__10057_ (
);

FILL FILL_0__11091_ (
);

FILL FILL_1__9933_ (
);

FILL FILL_1__9513_ (
);

FILL FILL_3__9019_ (
);

FILL FILL_0__6897_ (
);

FILL FILL_0__6477_ (
);

NAND3X1 _8583_ (
    .A(_1989_),
    .B(_2017_),
    .C(_2019_),
    .Y(_2020_)
);

OAI21X1 _8163_ (
    .A(_1598_),
    .B(_1601_),
    .C(_1595_),
    .Y(_1606_)
);

FILL FILL_1__10831_ (
);

FILL FILL_1__10411_ (
);

FILL FILL_2__7856_ (
);

FILL FILL_3__12689_ (
);

FILL FILL_2__7436_ (
);

FILL FILL_3__12269_ (
);

FILL FILL_2__7016_ (
);

FILL FILL254550x158550 (
);

NAND3X1 _12581_ (
    .A(_5612_),
    .B(_5620_),
    .C(_5622_),
    .Y(_5623_)
);

FILL FILL_0__12296_ (
);

NAND3X1 _12161_ (
    .A(_5242_),
    .B(_5276_),
    .C(_5274_),
    .Y(_5277_)
);

FILL FILL_2__12623_ (
);

FILL FILL_2__12203_ (
);

OAI21X1 _9788_ (
    .A(_3130_),
    .B(_3113_),
    .C(_3129_),
    .Y(_3132_)
);

AOI21X1 _9368_ (
    .A(_2723_),
    .B(_2725_),
    .C(_2721_),
    .Y(_2726_)
);

FILL FILL_0__8623_ (
);

FILL FILL_3__6720_ (
);

FILL FILL_0__8203_ (
);

FILL FILL_0__10609_ (
);

FILL FILL_3__9192_ (
);

DFFPOSX1 _13366_ (
    .D(\Y[6] [4]),
    .CLK(clk_bF$buf39),
    .Q(\u_fir_pe7.rYin [4])
);

FILL FILL_1__6638_ (
);

FILL FILL_2__13408_ (
);

FILL FILL_0__9828_ (
);

FILL FILL_3__7925_ (
);

FILL FILL_0__9408_ (
);

FILL FILL_3__7505_ (
);

FILL FILL_2__8394_ (
);

FILL FILL_0__10782_ (
);

FILL FILL_0__10362_ (
);

NAND2X1 _7854_ (
    .A(_1362_),
    .B(_1366_),
    .Y(_1368_)
);

INVX1 _7434_ (
    .A(_953_),
    .Y(_954_)
);

AND2X2 _7014_ (
    .A(_603_),
    .B(_602_),
    .Y(_607_)
);

FILL FILL_1__6391_ (
);

FILL FILL_2__13161_ (
);

FILL FILL_2__6707_ (
);

FILL FILL_1__12994_ (
);

FILL FILL_1__12574_ (
);

FILL FILL_1__12154_ (
);

FILL FILL_0__11987_ (
);

FILL FILL_0__9581_ (
);

FILL FILL_2__9599_ (
);

FILL FILL_2__9179_ (
);

FILL FILL_0__9161_ (
);

OAI21X1 _11852_ (
    .A(_4894_),
    .B(_4971_),
    .C(_4888_),
    .Y(_4972_)
);

FILL FILL_0__11567_ (
);

NOR2X1 _11432_ (
    .A(_4620_),
    .B(_4619_),
    .Y(_4621_)
);

FILL FILL_0__11147_ (
);

INVX1 _11012_ (
    .A(_4210_),
    .Y(_4211_)
);

FILL FILL_3__12901_ (
);

AOI21X1 _8639_ (
    .A(gnd),
    .B(\X[2] [6]),
    .C(_2006_),
    .Y(_2075_)
);

NAND2X1 _8219_ (
    .A(_1660_),
    .B(_1654_),
    .Y(_2389_[4])
);

FILL FILL_1__7596_ (
);

FILL FILL_1__7176_ (
);

FILL FILL_3__8463_ (
);

AOI22X1 _12637_ (
    .A(gnd),
    .B(\X[6] [4]),
    .C(_5667_),
    .D(_5669_),
    .Y(_5678_)
);

FILL FILL_3__8043_ (
);

OAI21X1 _12217_ (
    .A(_5278_),
    .B(_5331_),
    .C(_5274_),
    .Y(_5332_)
);

FILL FILL_2__6880_ (
);

FILL FILL_2__6460_ (
);

FILL FILL_3__11293_ (
);

FILL FILL_2__10286_ (
);

FILL FILL_1__9742_ (
);

FILL FILL_1__9322_ (
);

FILL FILL_3__9248_ (
);

NAND3X1 _8392_ (
    .A(_1819_),
    .B(_1828_),
    .C(_1830_),
    .Y(_1831_)
);

FILL FILL_1__10640_ (
);

FILL FILL_1__10220_ (
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf55)
);

FILL FILL_2__7665_ (
);

CLKBUF1 CLKBUF1_insert15 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert16 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert17 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert18 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert19 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf50)
);

AND2X2 _12390_ (
    .A(\u_fir_pe6.rYin [9]),
    .B(\u_fir_pe6.mul [9]),
    .Y(_5494_)
);

OAI21X1 _6705_ (
    .A(_222_),
    .B(_302_),
    .C(_271_),
    .Y(_303_)
);

FILL FILL_2__12852_ (
);

FILL FILL_2__12432_ (
);

FILL FILL_2__12012_ (
);

AND2X2 _9597_ (
    .A(_2933_),
    .B(_2928_),
    .Y(_2951_)
);

OAI21X1 _9177_ (
    .A(_3169_),
    .B(_2535_),
    .C(_2536_),
    .Y(_2537_)
);

FILL FILL_1__11845_ (
);

FILL FILL_1__11425_ (
);

FILL FILL_1__11005_ (
);

FILL FILL_0__8852_ (
);

FILL FILL_0__8432_ (
);

FILL FILL_0__10838_ (
);

FILL FILL_0__10418_ (
);

AOI21X1 _10703_ (
    .A(\X[4] [0]),
    .B(vdd),
    .C(_3888_),
    .Y(_3965_)
);

FILL FILL_0__8012_ (
);

NAND3X1 _13175_ (
    .A(_6205_),
    .B(_6206_),
    .C(_6204_),
    .Y(_6207_)
);

FILL FILL_2__9811_ (
);

FILL FILL_1__6867_ (
);

FILL FILL_1__6447_ (
);

FILL FILL_2__13217_ (
);

FILL FILL_0__9637_ (
);

FILL FILL_0__9217_ (
);

AOI21X1 _11908_ (
    .A(_5026_),
    .B(_5025_),
    .C(_5022_),
    .Y(_5027_)
);

FILL FILL_3__10984_ (
);

FILL FILL_3__10144_ (
);

FILL FILL_0__10591_ (
);

FILL FILL_0__10171_ (
);

FILL FILL_3__8939_ (
);

OAI21X1 _7663_ (
    .A(_1101_),
    .B(_1105_),
    .C(_1110_),
    .Y(_1180_)
);

DFFPOSX1 _7243_ (
    .D(_795_[4]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.mul [4])
);

FILL FILL_2__6936_ (
);

FILL FILL_3__11769_ (
);

FILL FILL_2__6516_ (
);

FILL FILL_1__12383_ (
);

FILL FILL_0__9390_ (
);

FILL FILL_0__11796_ (
);

NAND2X1 _11661_ (
    .A(gnd),
    .B(\X[7] [0]),
    .Y(_4784_)
);

FILL FILL_0__11376_ (
);

NAND2X1 _11241_ (
    .A(_4437_),
    .B(_4436_),
    .Y(_4781_[9])
);

FILL FILL_2__11703_ (
);

OAI21X1 _8868_ (
    .A(_2275_),
    .B(_2276_),
    .C(_2290_),
    .Y(_2291_)
);

INVX1 _8448_ (
    .A(_1882_),
    .Y(_1887_)
);

NOR2X1 _8028_ (
    .A(_1531_),
    .B(_1530_),
    .Y(_1532_)
);

FILL FILL_0__7703_ (
);

FILL FILL_1__13168_ (
);

FILL FILL_3__8692_ (
);

NAND2X1 _12866_ (
    .A(vdd),
    .B(\X[6]_5_bF$buf0 ),
    .Y(_5904_)
);

INVX1 _12446_ (
    .A(_5544_),
    .Y(_5549_)
);

NAND3X1 _12026_ (
    .A(_5142_),
    .B(_5143_),
    .C(_5141_),
    .Y(_5144_)
);

FILL FILL_2__12908_ (
);

FILL FILL_0__13102_ (
);

FILL FILL_0__8908_ (
);

FILL FILL_2__10095_ (
);

FILL FILL_1__9971_ (
);

FILL FILL_1__9551_ (
);

FILL FILL_1__9131_ (
);

FILL FILL_3__9477_ (
);

FILL FILL_2__7894_ (
);

FILL FILL_2__7474_ (
);

FILL FILL_2__7054_ (
);

NAND3X1 _6934_ (
    .A(_525_),
    .B(_528_),
    .C(_482_),
    .Y(_529_)
);

NAND3X1 _6514_ (
    .A(_112_),
    .B(_113_),
    .C(_114_),
    .Y(_115_)
);

FILL FILL_2__12661_ (
);

FILL FILL_2__12241_ (
);

FILL FILL_1__11654_ (
);

FILL FILL_1__11234_ (
);

FILL FILL_2__8679_ (
);

FILL FILL_0__8661_ (
);

FILL FILL_0__8241_ (
);

FILL FILL_2__8259_ (
);

FILL FILL_0__10647_ (
);

NAND3X1 _10932_ (
    .A(_4131_),
    .B(_4125_),
    .C(_4128_),
    .Y(_4132_)
);

OAI22X1 _10512_ (
    .A(_3332_),
    .B(_3650_),
    .C(_3493_),
    .D(_3423_),
    .Y(_3785_)
);

FILL FILL_0__10227_ (
);

FILL FILL_2__9620_ (
);

FILL FILL_2__9200_ (
);

FILL FILL254250x144150 (
);

INVX1 _7719_ (
    .A(_1228_),
    .Y(_1236_)
);

FILL FILL_1__6676_ (
);

FILL FILL_2__13026_ (
);

FILL FILL_1__12859_ (
);

FILL FILL_1__12439_ (
);

FILL FILL_1__12019_ (
);

FILL FILL_0__9446_ (
);

FILL FILL_3__7543_ (
);

FILL FILL_0__9026_ (
);

OR2X2 _11717_ (
    .A(_4838_),
    .B(_4837_),
    .Y(_4839_)
);

FILL FILL_3__10793_ (
);

FILL FILL_3__10373_ (
);

FILL FILL_1__8822_ (
);

FILL FILL_1__8402_ (
);

FILL FILL_3__8328_ (
);

NAND2X1 _7892_ (
    .A(_1403_),
    .B(_1404_),
    .Y(_1405_)
);

AOI21X1 _7472_ (
    .A(_915_),
    .B(_914_),
    .C(_851_),
    .Y(_992_)
);

OAI21X1 _7052_ (
    .A(_632_),
    .B(_633_),
    .C(_637_),
    .Y(_640_)
);

FILL FILL_3__11998_ (
);

FILL FILL_2__6745_ (
);

FILL FILL_3__11158_ (
);

FILL FILL_1__12192_ (
);

AND2X2 _11890_ (
    .A(\X[7] [3]),
    .B(gnd),
    .Y(_5009_)
);

NAND2X1 _11470_ (
    .A(_4654_),
    .B(_4649_),
    .Y(_4655_)
);

FILL FILL_0__11185_ (
);

INVX1 _11050_ (
    .A(_4152_),
    .Y(_4249_)
);

FILL FILL_1__9607_ (
);

FILL FILL_2__11932_ (
);

FILL FILL_2__11512_ (
);

AOI22X1 _8677_ (
    .A(\X[2]_5_bF$buf2 ),
    .B(gnd),
    .C(_2071_),
    .D(_2072_),
    .Y(_2112_)
);

NAND3X1 _8257_ (
    .A(_1689_),
    .B(_1685_),
    .C(_1691_),
    .Y(_1698_)
);

FILL FILL_1__10925_ (
);

FILL FILL_1__10505_ (
);

FILL FILL_0__7932_ (
);

FILL FILL_0__7512_ (
);

FILL FILL_1__13397_ (
);

NAND2X1 _12675_ (
    .A(_5714_),
    .B(_5713_),
    .Y(_5715_)
);

NAND3X1 _12255_ (
    .A(_5159_),
    .B(_5232_),
    .C(_5338_),
    .Y(_5369_)
);

FILL FILL_2__12717_ (
);

FILL FILL_0__13331_ (
);

FILL FILL_0__8717_ (
);

FILL FILL_3__6814_ (
);

FILL FILL_1__9780_ (
);

FILL FILL_1__9360_ (
);

FILL FILL_2__7283_ (
);

AOI21X1 _6743_ (
    .A(_336_),
    .B(_340_),
    .C(_322_),
    .Y(_341_)
);

FILL FILL_2__12890_ (
);

FILL FILL_2__12050_ (
);

FILL FILL_1__11883_ (
);

FILL FILL_1__11463_ (
);

FILL FILL_1__11043_ (
);

FILL FILL_0__8890_ (
);

FILL FILL_2__8488_ (
);

FILL FILL_0__8470_ (
);

FILL FILL_0__10876_ (
);

DFFPOSX1 _10741_ (
    .D(\Y[4] [10]),
    .CLK(clk_bF$buf45),
    .Q(\u_fir_pe4.rYin [10])
);

FILL FILL_0__10456_ (
);

FILL FILL_2__8068_ (
);

FILL FILL_0__8050_ (
);

NAND2X1 _10321_ (
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3598_)
);

FILL FILL_0__10036_ (
);

NOR2X1 _7948_ (
    .A(_1452_),
    .B(_1453_),
    .Y(_1454_)
);

AOI21X1 _7528_ (
    .A(_1044_),
    .B(_1046_),
    .C(_1043_),
    .Y(_1047_)
);

INVX1 _7108_ (
    .A(\u_fir_pe0.mul [8]),
    .Y(_691_)
);

FILL FILL_1__6485_ (
);

FILL FILL_2__13255_ (
);

FILL FILL_1__12668_ (
);

FILL FILL_1__12248_ (
);

FILL FILL_0__9675_ (
);

FILL FILL_3__7772_ (
);

FILL FILL_0__9255_ (
);

OAI21X1 _11946_ (
    .A(_5051_),
    .B(_5055_),
    .C(_5058_),
    .Y(_5065_)
);

INVX1 _11526_ (
    .A(\u_fir_pe5.mul [10]),
    .Y(_4710_)
);

INVX1 _11106_ (
    .A(gnd),
    .Y(_4304_)
);

FILL FILL_0__12602_ (
);

FILL FILL_1__8631_ (
);

FILL FILL_1__8211_ (
);

FILL FILL_3__8557_ (
);

NOR2X1 _7281_ (
    .A(_1528_),
    .B(_799_),
    .Y(_804_)
);

FILL FILL_2__6974_ (
);

FILL FILL_2__6554_ (
);

FILL FILL_3__11387_ (
);

FILL FILL_1__9416_ (
);

FILL FILL_2__11741_ (
);

FILL FILL_2__11321_ (
);

INVX1 _8486_ (
    .A(_1918_),
    .Y(_1924_)
);

INVX1 _8066_ (
    .A(_1569_),
    .Y(_1570_)
);

FILL FILL_1__10314_ (
);

FILL FILL_2__7759_ (
);

FILL FILL_0__7741_ (
);

FILL FILL_0__7321_ (
);

FILL FILL_2__7339_ (
);

DFFPOSX1 _12484_ (
    .D(\X[7] [7]),
    .CLK(clk_bF$buf37),
    .Q(_6376_[7])
);

FILL FILL_0__12199_ (
);

AND2X2 _12064_ (
    .A(_4914_),
    .B(_5103_),
    .Y(_5181_)
);

FILL FILL_2__8700_ (
);

FILL FILL_3__13113_ (
);

FILL FILL_2__12946_ (
);

FILL FILL_2__12526_ (
);

FILL FILL_2__12106_ (
);

FILL FILL_0__13140_ (
);

FILL FILL_1__11939_ (
);

FILL FILL_1__11519_ (
);

FILL FILL_0__8946_ (
);

FILL FILL_0__8526_ (
);

FILL FILL_3__9095_ (
);

NOR2X1 _13269_ (
    .A(_6292_),
    .B(_6291_),
    .Y(_6293_)
);

FILL FILL_2__9905_ (
);

FILL FILL_2__7092_ (
);

FILL FILL_1__7902_ (
);

FILL FILL_3__7828_ (
);

NOR2X1 _6972_ (
    .A(_473_),
    .B(_526_),
    .Y(_566_)
);

AND2X2 _6552_ (
    .A(_147_),
    .B(_151_),
    .Y(_152_)
);

FILL FILL_1__11692_ (
);

FILL FILL_3__10238_ (
);

FILL FILL_1__11272_ (
);

FILL FILL_2__8297_ (
);

FILL FILL_0__10685_ (
);

OAI21X1 _10970_ (
    .A(_4165_),
    .B(_4166_),
    .C(_4123_),
    .Y(_4170_)
);

AND2X2 _10550_ (
    .A(\u_fir_pe4.rYin [0]),
    .B(\u_fir_pe4.mul [0]),
    .Y(_3819_)
);

FILL FILL_0__10265_ (
);

OAI21X1 _10130_ (
    .A(_3407_),
    .B(_3408_),
    .C(_3398_),
    .Y(_3409_)
);

OAI22X1 _7757_ (
    .A(_1128_),
    .B(_1209_),
    .C(_1271_),
    .D(_1272_),
    .Y(_1273_)
);

INVX1 _7337_ (
    .A(_842_),
    .Y(_859_)
);

FILL FILL_2__13064_ (
);

FILL FILL_1__12897_ (
);

FILL FILL_1__12057_ (
);

FILL FILL_0__9484_ (
);

FILL FILL_0__9064_ (
);

NAND3X1 _11755_ (
    .A(gnd),
    .B(\X[7] [2]),
    .C(_4875_),
    .Y(_4876_)
);

FILL FILL_3__7161_ (
);

NAND2X1 _11335_ (
    .A(_4524_),
    .B(_4521_),
    .Y(_4530_)
);

FILL FILL_0__12831_ (
);

FILL FILL_0__12411_ (
);

FILL FILL_1__7499_ (
);

FILL FILL_1__7079_ (
);

NAND2X1 _9903_ (
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3975_)
);

FILL FILL_1__8860_ (
);

FILL FILL_1__8440_ (
);

FILL FILL_1__8020_ (
);

FILL FILL_3__8786_ (
);

INVX1 _7090_ (
    .A(\u_fir_pe0.mul [6]),
    .Y(_674_)
);

FILL FILL_2__6783_ (
);

FILL FILL_2__10189_ (
);

FILL FILL_1__9645_ (
);

FILL FILL_1__9225_ (
);

FILL FILL_2__11970_ (
);

FILL FILL_2__11550_ (
);

FILL FILL_2__11130_ (
);

AND2X2 _8295_ (
    .A(\X[2] [2]),
    .B(vdd),
    .Y(_1735_)
);

FILL FILL_1__10963_ (
);

FILL FILL_1__10543_ (
);

FILL FILL_1__10123_ (
);

FILL FILL_2__7988_ (
);

FILL FILL_0__7970_ (
);

FILL FILL_2__7568_ (
);

FILL FILL_0__7550_ (
);

FILL FILL_2__7148_ (
);

FILL FILL_0__7130_ (
);

INVX1 _12293_ (
    .A(_5364_),
    .Y(_5405_)
);

INVX1 _6608_ (
    .A(_202_),
    .Y(_207_)
);

FILL FILL_2__12755_ (
);

FILL FILL_2__12335_ (
);

FILL FILL_1__11748_ (
);

FILL FILL_1__11328_ (
);

FILL FILL254550x21750 (
);

FILL FILL_0__8755_ (
);

FILL FILL_0__8335_ (
);

FILL FILL_3__6432_ (
);

INVX1 _10606_ (
    .A(\u_fir_pe4.rYin [7]),
    .Y(_3869_)
);

FILL FILL253950x169350 (
);

INVX1 _13078_ (
    .A(_6110_),
    .Y(_6113_)
);

FILL FILL_2__9714_ (
);

FILL FILL_1__7711_ (
);

NAND2X1 _6781_ (
    .A(_374_),
    .B(_378_),
    .Y(_796_[8])
);

FILL FILL_3__10887_ (
);

FILL FILL_3__10467_ (
);

FILL FILL_1__11081_ (
);

FILL FILL_0__10494_ (
);

FILL FILL_0__10074_ (
);

FILL FILL_1__8916_ (
);

FILL FILL_2__10821_ (
);

FILL FILL_2__10401_ (
);

NOR2X1 _7986_ (
    .A(_1487_),
    .B(_1488_),
    .Y(_1489_)
);

NAND3X1 _7566_ (
    .A(_985_),
    .B(_1083_),
    .C(_1084_),
    .Y(_1085_)
);

OAI21X1 _7146_ (
    .A(_726_),
    .B(_727_),
    .C(_722_),
    .Y(_730_)
);

FILL FILL_2__13293_ (
);

FILL FILL_0__6821_ (
);

FILL FILL_2__6839_ (
);

FILL FILL_2__6419_ (
);

FILL FILL_0__6401_ (
);

FILL FILL_1__12286_ (
);

FILL FILL_0__9293_ (
);

OAI21X1 _11984_ (
    .A(_4797_),
    .B(_5101_),
    .C(_4807_),
    .Y(_5102_)
);

FILL FILL_0__11699_ (
);

FILL FILL_3__7390_ (
);

NOR2X1 _11564_ (
    .A(\u_fir_pe5.rYin [14]),
    .B(\u_fir_pe5.mul [14]),
    .Y(_4748_)
);

FILL FILL_0__11279_ (
);

OAI21X1 _11144_ (
    .A(_4341_),
    .B(_4337_),
    .C(_4288_),
    .Y(_4342_)
);

FILL FILL_3__12613_ (
);

FILL FILL_0__12640_ (
);

FILL FILL_0__12220_ (
);

FILL FILL_0__7606_ (
);

INVX1 _9712_ (
    .A(\u_fir_pe3.mul [5]),
    .Y(_3057_)
);

NAND2X1 _12769_ (
    .A(_5806_),
    .B(_5807_),
    .Y(_5808_)
);

FILL FILL_3__8175_ (
);

AND2X2 _12349_ (
    .A(_5453_),
    .B(_5452_),
    .Y(_5572_[5])
);

FILL FILL_0__13005_ (
);

FILL FILL_2__6592_ (
);

FILL FILL_3__6908_ (
);

FILL FILL_1__9454_ (
);

FILL FILL_1__9034_ (
);

FILL FILL_1__10772_ (
);

FILL FILL_1__10352_ (
);

FILL FILL_2__7797_ (
);

FILL FILL_2__7377_ (
);

INVX1 _6837_ (
    .A(_426_),
    .Y(_434_)
);

NAND3X1 _6417_ (
    .A(_782_),
    .B(_14_),
    .C(_17_),
    .Y(_20_)
);

FILL FILL_2__12984_ (
);

FILL FILL_2__12564_ (
);

FILL FILL_2__12144_ (
);

FILL FILL_1__11977_ (
);

FILL FILL_1__11557_ (
);

FILL FILL_1__11137_ (
);

FILL FILL_0__8564_ (
);

FILL FILL_3__6661_ (
);

FILL FILL_0__8144_ (
);

NAND3X1 _10835_ (
    .A(_4013_),
    .B(_4036_),
    .C(_4035_),
    .Y(_4037_)
);

NAND2X1 _10415_ (
    .A(_3683_),
    .B(_3689_),
    .Y(_3691_)
);

FILL FILL_2__9943_ (
);

FILL FILL_0__11911_ (
);

FILL FILL_2__9523_ (
);

FILL FILL_2__9103_ (
);

FILL FILL_1__6999_ (
);

FILL FILL_1__6579_ (
);

FILL FILL_1__7940_ (
);

FILL FILL_1__7520_ (
);

FILL FILL_1__7100_ (
);

FILL FILL_0__9769_ (
);

FILL FILL_3__7866_ (
);

FILL FILL_0__9349_ (
);

FILL FILL_3__7446_ (
);

FILL FILL_3__7026_ (
);

OAI21X1 _6590_ (
    .A(_112_),
    .B(_189_),
    .C(_106_),
    .Y(_190_)
);

FILL FILL_3__10696_ (
);

FILL FILL_1__8725_ (
);

FILL FILL_1__8305_ (
);

FILL FILL_2__10630_ (
);

FILL FILL_2__10210_ (
);

NOR2X1 _7795_ (
    .A(_1290_),
    .B(_1295_),
    .Y(_1310_)
);

AOI22X1 _7375_ (
    .A(gnd),
    .B(\X[1] [4]),
    .C(_885_),
    .D(_887_),
    .Y(_896_)
);

FILL FILL_0__6630_ (
);

FILL FILL_2__6648_ (
);

FILL FILL_1__12095_ (
);

AND2X2 _11793_ (
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4913_)
);

FILL FILL_0__11088_ (
);

OAI21X1 _11373_ (
    .A(_4564_),
    .B(_4566_),
    .C(_4545_),
    .Y(_4567_)
);

FILL FILL_3__12842_ (
);

FILL FILL_3__12002_ (
);

FILL FILL_2__11835_ (
);

FILL FILL_2__11415_ (
);

FILL FILL_1__10828_ (
);

FILL FILL_1__10408_ (
);

FILL FILL_0__7835_ (
);

AND2X2 _9941_ (
    .A(gnd),
    .B(\X[4] [1]),
    .Y(_3223_)
);

FILL FILL_0__7415_ (
);

NAND3X1 _9521_ (
    .A(_2798_),
    .B(_2876_),
    .C(_2806_),
    .Y(_2877_)
);

INVX1 _9101_ (
    .A(_2461_),
    .Y(_2462_)
);

NAND2X1 _12998_ (
    .A(_6033_),
    .B(_5876_),
    .Y(_6034_)
);

NAND3X1 _12578_ (
    .A(vdd),
    .B(\X[6] [2]),
    .C(_5610_),
    .Y(_5620_)
);

NAND3X1 _12158_ (
    .A(_5269_),
    .B(_5273_),
    .C(_5243_),
    .Y(_5274_)
);

FILL FILL_3__13207_ (
);

FILL FILL_0__13234_ (
);

FILL FILL_1__9683_ (
);

FILL FILL_1__9263_ (
);

FILL FILL_3__9189_ (
);

FILL FILL_1__10581_ (
);

FILL FILL_1__10161_ (
);

FILL FILL_2__7186_ (
);

AOI21X1 _6646_ (
    .A(_244_),
    .B(_243_),
    .C(_240_),
    .Y(_245_)
);

FILL FILL_2__12793_ (
);

FILL FILL_2__12373_ (
);

FILL FILL_1__11786_ (
);

FILL FILL_1__11366_ (
);

FILL FILL_0__8793_ (
);

FILL FILL_3__6890_ (
);

FILL FILL_0__8373_ (
);

FILL FILL_0__10779_ (
);

FILL FILL_0__10359_ (
);

AOI21X1 _10644_ (
    .A(_3902_),
    .B(_3880_),
    .C(_3900_),
    .Y(_3907_)
);

NAND3X1 _10224_ (
    .A(_3499_),
    .B(_3501_),
    .C(_3500_),
    .Y(_3502_)
);

FILL FILL_2__9752_ (
);

FILL FILL_2__9332_ (
);

FILL FILL_0__11720_ (
);

FILL FILL_0__11300_ (
);

FILL FILL_1__6388_ (
);

FILL FILL_2__13158_ (
);

FILL FILL_0__9998_ (
);

FILL FILL_0__9578_ (
);

FILL FILL_0__9158_ (
);

NAND3X1 _11849_ (
    .A(_4966_),
    .B(_4967_),
    .C(_4968_),
    .Y(_4969_)
);

INVX1 _11429_ (
    .A(\u_fir_pe5.mul [1]),
    .Y(_4618_)
);

AOI21X1 _11009_ (
    .A(_4147_),
    .B(_4151_),
    .C(_4140_),
    .Y(_4208_)
);

FILL FILL_0__12925_ (
);

FILL FILL_3__10085_ (
);

FILL FILL_1__8534_ (
);

INVX1 _7184_ (
    .A(_762_),
    .Y(_767_)
);

FILL FILL_3__9401_ (
);

FILL FILL_2__6877_ (
);

FILL FILL_2__6457_ (
);

NAND3X1 _11182_ (
    .A(_4377_),
    .B(_4373_),
    .C(_4378_),
    .Y(_4379_)
);

FILL FILL_1__9739_ (
);

FILL FILL_1__9319_ (
);

FILL FILL_3__12231_ (
);

FILL FILL_2__11644_ (
);

FILL FILL_2__11224_ (
);

OAI21X1 _8389_ (
    .A(_1609_),
    .B(_1827_),
    .C(_1822_),
    .Y(_1828_)
);

FILL FILL_1__10637_ (
);

FILL FILL_1__10217_ (
);

FILL FILL_0__7644_ (
);

NAND2X1 _9750_ (
    .A(_3090_),
    .B(_3093_),
    .Y(_3094_)
);

NAND2X1 _9330_ (
    .A(_2687_),
    .B(_2686_),
    .Y(_2688_)
);

INVX1 _12387_ (
    .A(_5474_),
    .Y(_5490_)
);

FILL FILL_2__8603_ (
);

FILL FILL_3__13016_ (
);

FILL FILL_2__12849_ (
);

FILL FILL_2__12429_ (
);

FILL FILL_2__12009_ (
);

FILL FILL_0__13043_ (
);

FILL FILL_1__6600_ (
);

FILL FILL_0__8849_ (
);

FILL FILL_0__8429_ (
);

FILL FILL_3__6526_ (
);

FILL FILL_0__8009_ (
);

FILL FILL_1__9492_ (
);

FILL FILL_1__9072_ (
);

FILL FILL_2__9808_ (
);

FILL FILL_1__10390_ (
);

FILL FILL_1__7805_ (
);

NOR2X1 _6875_ (
    .A(_406_),
    .B(_403_),
    .Y(_471_)
);

OR2X2 _6455_ (
    .A(_56_),
    .B(_55_),
    .Y(_57_)
);

FILL FILL_2__12182_ (
);

FILL FILL_1__11175_ (
);

FILL FILL_0__8182_ (
);

FILL FILL_0__10588_ (
);

INVX1 _10873_ (
    .A(gnd),
    .Y(_4074_)
);

NAND2X1 _10453_ (
    .A(_3720_),
    .B(_3723_),
    .Y(_3728_)
);

FILL FILL_0__10168_ (
);

NAND3X1 _10033_ (
    .A(_3308_),
    .B(_3313_),
    .C(_3255_),
    .Y(_3314_)
);

FILL FILL_3__11922_ (
);

FILL FILL_2__9981_ (
);

FILL FILL_2__10915_ (
);

FILL FILL_2__9561_ (
);

FILL FILL_2__9141_ (
);

FILL FILL_0__6915_ (
);

AOI21X1 _8601_ (
    .A(_1894_),
    .B(_1959_),
    .C(_2037_),
    .Y(_2038_)
);

FILL FILL_0__9387_ (
);

FILL FILL_3__7484_ (
);

INVX1 _11658_ (
    .A(_5569_),
    .Y(_5570_)
);

AND2X2 _11238_ (
    .A(_4434_),
    .B(_4427_),
    .Y(_4435_)
);

FILL FILL_3__12707_ (
);

FILL FILL_1__13321_ (
);

FILL FILL_0__12734_ (
);

FILL FILL_0__12314_ (
);

OAI21X1 _9806_ (
    .A(_3142_),
    .B(_3143_),
    .C(_3147_),
    .Y(_3149_)
);

FILL FILL_1__8763_ (
);

FILL FILL_1__8343_ (
);

FILL FILL_3__8269_ (
);

FILL FILL_3__9630_ (
);

FILL FILL_2__6686_ (
);

FILL FILL_3__11099_ (
);

FILL FILL_1__9968_ (
);

FILL FILL_1__9548_ (
);

FILL FILL_1__9128_ (
);

FILL FILL_2__11873_ (
);

FILL FILL_2__11453_ (
);

FILL FILL_2__11033_ (
);

INVX1 _8198_ (
    .A(_1626_),
    .Y(_1640_)
);

FILL FILL_1__10866_ (
);

FILL FILL_1__10446_ (
);

FILL FILL_1__10026_ (
);

FILL FILL_0__7873_ (
);

FILL FILL_0__7453_ (
);

FILL FILL_0__7033_ (
);

NAND3X1 _12196_ (
    .A(_5307_),
    .B(_5310_),
    .C(_5264_),
    .Y(_5311_)
);

FILL FILL_2__8832_ (
);

FILL FILL_2__8412_ (
);

FILL FILL_0__10800_ (
);

FILL FILL_2__12658_ (
);

FILL FILL_2__12238_ (
);

FILL FILL_0__13272_ (
);

FILL FILL_0__8658_ (
);

FILL FILL_3__6755_ (
);

FILL FILL_0__8238_ (
);

INVX2 _10929_ (
    .A(\X[5] [6]),
    .Y(_4129_)
);

INVX1 _10509_ (
    .A(_3781_),
    .Y(_3782_)
);

FILL FILL_2__9617_ (
);

FILL FILL_1__7614_ (
);

OAI21X1 _6684_ (
    .A(_269_),
    .B(_273_),
    .C(_276_),
    .Y(_283_)
);

FILL FILL_0__10397_ (
);

AND2X2 _10682_ (
    .A(_3945_),
    .B(_3944_),
    .Y(_3978_[13])
);

AOI21X1 _10262_ (
    .A(_3539_),
    .B(_3534_),
    .C(_3503_),
    .Y(_3540_)
);

FILL FILL_1__8819_ (
);

FILL FILL_3__11731_ (
);

FILL FILL_3__11311_ (
);

FILL FILL_2__9790_ (
);

FILL FILL_2__9370_ (
);

FILL FILL_2__10304_ (
);

NAND3X1 _7889_ (
    .A(_1375_),
    .B(_1377_),
    .C(_1401_),
    .Y(_1402_)
);

NAND3X1 _7469_ (
    .A(_933_),
    .B(_982_),
    .C(_983_),
    .Y(_989_)
);

INVX1 _7049_ (
    .A(_637_),
    .Y(_638_)
);

FILL FILL_2__13196_ (
);

FILL FILL_0__6724_ (
);

NAND2X1 _8830_ (
    .A(_2253_),
    .B(_2255_),
    .Y(_2256_)
);

NOR2X1 _8410_ (
    .A(_1835_),
    .B(_1848_),
    .Y(_1849_)
);

FILL FILL_1__12189_ (
);

FILL FILL_0__9196_ (
);

OAI21X1 _11887_ (
    .A(_4955_),
    .B(_5005_),
    .C(_4949_),
    .Y(_5006_)
);

NOR2X1 _11467_ (
    .A(_4650_),
    .B(_4651_),
    .Y(_4652_)
);

OAI21X1 _11047_ (
    .A(_4235_),
    .B(_4230_),
    .C(_4237_),
    .Y(_4246_)
);

FILL FILL_3__12936_ (
);

FILL FILL_1__13130_ (
);

FILL FILL_2__11929_ (
);

FILL FILL_0__12963_ (
);

FILL FILL_2__11509_ (
);

FILL FILL_0__12543_ (
);

FILL FILL_0__12123_ (
);

FILL FILL_0__7929_ (
);

FILL FILL_0__7509_ (
);

NAND3X1 _9615_ (
    .A(_2953_),
    .B(_2963_),
    .C(_2966_),
    .Y(_2969_)
);

FILL FILL_1__8572_ (
);

FILL FILL_1__8152_ (
);

FILL FILL_3__8498_ (
);

FILL FILL_0__13328_ (
);

FILL FILL_2__6495_ (
);

FILL FILL_1__9777_ (
);

FILL FILL_1__9357_ (
);

FILL FILL_2__11682_ (
);

FILL FILL_2__11262_ (
);

FILL FILL_1__10675_ (
);

FILL FILL_1__10255_ (
);

FILL FILL_0__7682_ (
);

FILL FILL_0__7262_ (
);

FILL FILL_2__8641_ (
);

FILL FILL_2__8221_ (
);

FILL FILL_3__13054_ (
);

FILL FILL_2__12887_ (
);

FILL FILL_2__12047_ (
);

FILL FILL_0__13081_ (
);

FILL FILL_0__8887_ (
);

FILL FILL_3__6984_ (
);

FILL FILL_0__8467_ (
);

DFFPOSX1 _10738_ (
    .D(\Y[4] [7]),
    .CLK(clk_bF$buf7),
    .Q(\u_fir_pe4.rYin [7])
);

FILL FILL_0__8047_ (
);

NAND2X1 _10318_ (
    .A(_3594_),
    .B(_3591_),
    .Y(_3595_)
);

FILL FILL_1__12821_ (
);

FILL FILL_1__12401_ (
);

FILL FILL_2__9426_ (
);

FILL FILL_0__11814_ (
);

FILL FILL_1__7843_ (
);

FILL FILL_1__7423_ (
);

FILL FILL_1__7003_ (
);

FILL FILL_3__7769_ (
);

NAND3X1 _6493_ (
    .A(gnd),
    .B(Xin[2]),
    .C(_93_),
    .Y(_94_)
);

FILL FILL_3__8710_ (
);

FILL FILL_3__10179_ (
);

NAND2X1 _10491_ (
    .A(_3751_),
    .B(_3764_),
    .Y(_3765_)
);

NAND3X1 _10071_ (
    .A(gnd),
    .B(\X[4] [4]),
    .C(_3341_),
    .Y(_3351_)
);

FILL FILL_1__8628_ (
);

FILL FILL_1__8208_ (
);

FILL FILL_3__11540_ (
);

FILL FILL_2__10953_ (
);

FILL FILL_2__10533_ (
);

FILL FILL_2__10113_ (
);

OAI21X1 _7698_ (
    .A(_1214_),
    .B(_1116_),
    .C(_929_),
    .Y(_1215_)
);

AOI22X1 _7278_ (
    .A(vdd),
    .B(\X[1] [0]),
    .C(vdd),
    .D(\X[1] [1]),
    .Y(_801_)
);

FILL FILL_3__9915_ (
);

FILL FILL_0__6953_ (
);

FILL FILL_0__6533_ (
);

AND2X2 _11696_ (
    .A(gnd),
    .B(\X[7] [2]),
    .Y(_4818_)
);

NAND3X1 _11276_ (
    .A(_4455_),
    .B(_4471_),
    .C(_4469_),
    .Y(_4472_)
);

FILL FILL_2__7912_ (
);

FILL FILL_3__12325_ (
);

FILL FILL_2__11738_ (
);

FILL FILL_0__12772_ (
);

FILL FILL_2__11318_ (
);

FILL FILL_0__12352_ (
);

FILL FILL_0__7738_ (
);

DFFPOSX1 _9844_ (
    .D(_3181_[14]),
    .CLK(clk_bF$buf26),
    .Q(\Y[4] [14])
);

FILL FILL_0__7318_ (
);

AOI21X1 _9424_ (
    .A(\X[3] [3]),
    .B(gnd),
    .C(_2778_),
    .Y(_2781_)
);

DFFPOSX1 _9004_ (
    .D(_2390_[11]),
    .CLK(clk_bF$buf15),
    .Q(\u_fir_pe2.mul [11])
);

FILL FILL_1__8381_ (
);

FILL FILL_0__13137_ (
);

OAI21X1 _13002_ (
    .A(_6017_),
    .B(_6019_),
    .C(_6010_),
    .Y(_6038_)
);

FILL FILL_1__9586_ (
);

FILL FILL_1__9166_ (
);

FILL FILL_2__11491_ (
);

FILL FILL_2__11071_ (
);

FILL FILL_1__10484_ (
);

FILL FILL_1__10064_ (
);

FILL FILL_0__7491_ (
);

FILL FILL_2__7089_ (
);

FILL FILL_0__7071_ (
);

FILL FILL_3__10811_ (
);

FILL FILL_2__8870_ (
);

FILL FILL_2__8450_ (
);

FILL FILL_3__13283_ (
);

FILL FILL_2__8030_ (
);

INVX1 _6969_ (
    .A(_562_),
    .Y(_563_)
);

NAND2X1 _6549_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_149_)
);

FILL FILL_2__12696_ (
);

FILL FILL_2__12276_ (
);

NAND2X1 _7910_ (
    .A(_1421_),
    .B(_1385_),
    .Y(_1422_)
);

FILL FILL_1__11689_ (
);

FILL FILL_1__11269_ (
);

FILL FILL_0__8696_ (
);

FILL FILL_0__8276_ (
);

OAI21X1 _10967_ (
    .A(_4165_),
    .B(_4166_),
    .C(_4164_),
    .Y(_4167_)
);

OAI21X1 _10547_ (
    .A(_3755_),
    .B(_3805_),
    .C(_3783_),
    .Y(_3818_)
);

NAND3X1 _10127_ (
    .A(_3399_),
    .B(_3405_),
    .C(_3404_),
    .Y(_3406_)
);

FILL FILL_1__12630_ (
);

FILL FILL_1__12210_ (
);

FILL FILL_2__9655_ (
);

FILL FILL_2__9235_ (
);

FILL FILL_0__11203_ (
);

FILL FILL_1__7652_ (
);

FILL FILL_3__7578_ (
);

FILL FILL_1__13415_ (
);

FILL FILL_0__12828_ (
);

FILL FILL_0__12408_ (
);

FILL FILL_1__8857_ (
);

FILL FILL_1__8437_ (
);

FILL FILL_1__8017_ (
);

FILL FILL_2__10342_ (
);

AND2X2 _7087_ (
    .A(_671_),
    .B(_670_),
    .Y(_790_[5])
);

FILL FILL_3__9724_ (
);

FILL FILL_0__6762_ (
);

INVX1 _11085_ (
    .A(_4267_),
    .Y(_4283_)
);

FILL FILL_2__7721_ (
);

FILL FILL_3__12554_ (
);

FILL FILL_2__7301_ (
);

FILL FILL_2__11967_ (
);

FILL FILL_2__11547_ (
);

FILL FILL_0__12581_ (
);

FILL FILL_2__11127_ (
);

FILL FILL_0__12161_ (
);

FILL FILL_0__7967_ (
);

FILL FILL_0__7547_ (
);

NAND3X1 _9653_ (
    .A(_2973_),
    .B(_2975_),
    .C(_3003_),
    .Y(_3005_)
);

FILL FILL_0__7127_ (
);

NAND3X1 _9233_ (
    .A(_2586_),
    .B(_2587_),
    .C(_2592_),
    .Y(_2593_)
);

FILL FILL_1__8190_ (
);

FILL FILL_1__11901_ (
);

FILL FILL_2__8926_ (
);

FILL FILL_2__8506_ (
);

NOR2X1 _13231_ (
    .A(\u_fir_pe7.rYin [6]),
    .B(\u_fir_pe7.mul [6]),
    .Y(_6255_)
);

FILL FILL_1__6923_ (
);

FILL FILL_1__6503_ (
);

FILL FILL_3__6849_ (
);

FILL FILL_1__9395_ (
);

FILL FILL_1__10293_ (
);

FILL FILL_1__7708_ (
);

FILL FILL_3__10620_ (
);

FILL FILL_3__10200_ (
);

AOI21X1 _6778_ (
    .A(_289_),
    .B(_204_),
    .C(_375_),
    .Y(_376_)
);

FILL FILL_2__12085_ (
);

FILL FILL_1__11498_ (
);

FILL FILL_1__11078_ (
);

NOR2X1 _10776_ (
    .A(_4765_),
    .B(_4745_),
    .Y(_4768_)
);

OAI21X1 _10356_ (
    .A(_3623_),
    .B(_3622_),
    .C(_3573_),
    .Y(_3633_)
);

FILL FILL_3__11825_ (
);

FILL FILL_3__11405_ (
);

FILL FILL_2__10818_ (
);

FILL FILL_2__9464_ (
);

FILL FILL_0__11852_ (
);

FILL FILL_2__9044_ (
);

FILL FILL_0__11432_ (
);

FILL FILL_0__11012_ (
);

FILL FILL_0__6818_ (
);

NOR2X1 _8924_ (
    .A(\u_fir_pe2.rYin [13]),
    .B(\u_fir_pe2.mul [13]),
    .Y(_2348_)
);

AOI21X1 _8504_ (
    .A(_1853_),
    .B(_1855_),
    .C(_1941_),
    .Y(_1942_)
);

FILL FILL_1__7881_ (
);

FILL FILL_1__7461_ (
);

FILL FILL_1__7041_ (
);

FILL FILL_3__7387_ (
);

FILL FILL_1__13224_ (
);

FILL FILL_0__12637_ (
);

AOI21X1 _12922_ (
    .A(_5876_),
    .B(_5946_),
    .C(_5958_),
    .Y(_5959_)
);

FILL FILL_0__12217_ (
);

DFFPOSX1 _12502_ (
    .D(_5574_[1]),
    .CLK(clk_bF$buf49),
    .Q(\u_fir_pe6.mul [1])
);

AND2X2 _9709_ (
    .A(_3054_),
    .B(_3053_),
    .Y(_3181_[4])
);

FILL FILL_1__8666_ (
);

FILL FILL_1__8246_ (
);

FILL FILL_2__10991_ (
);

FILL FILL_2__10571_ (
);

FILL FILL_2__10151_ (
);

FILL FILL_3__9953_ (
);

FILL FILL_3__9113_ (
);

FILL FILL_0__6991_ (
);

FILL FILL_0__6571_ (
);

FILL FILL_2__6589_ (
);

FILL FILL_2__7950_ (
);

FILL FILL_3__12783_ (
);

FILL FILL_2__7530_ (
);

FILL FILL_3__12363_ (
);

FILL FILL_2__7110_ (
);

FILL FILL_2__11776_ (
);

FILL FILL_2__11356_ (
);

FILL FILL_0__12390_ (
);

FILL FILL_1__10769_ (
);

FILL FILL_1__10349_ (
);

FILL FILL_0__7776_ (
);

DFFPOSX1 _9882_ (
    .D(_3187_[12]),
    .CLK(clk_bF$buf4),
    .Q(\u_fir_pe3.mul [12])
);

FILL FILL_0__7356_ (
);

AOI21X1 _9462_ (
    .A(_2734_),
    .B(_2740_),
    .C(_2815_),
    .Y(_2819_)
);

NAND3X1 _9042_ (
    .A(_3179_),
    .B(_2404_),
    .C(_2400_),
    .Y(_2405_)
);

FILL FILL_1__11710_ (
);

INVX1 _12099_ (
    .A(_5208_),
    .Y(_5216_)
);

FILL FILL_2__8735_ (
);

FILL FILL_2__8315_ (
);

FILL FILL_0__10703_ (
);

FILL FILL_3__13148_ (
);

FILL FILL_0__13175_ (
);

NAND2X1 _13040_ (
    .A(_6072_),
    .B(_6040_),
    .Y(_6076_)
);

FILL FILL_1__6732_ (
);

FILL FILL_1__12915_ (
);

FILL FILL_0__9922_ (
);

FILL FILL_0__11908_ (
);

FILL FILL_0__9502_ (
);

FILL FILL_1__7937_ (
);

FILL FILL_1__7517_ (
);

NAND3X1 _6587_ (
    .A(_184_),
    .B(_185_),
    .C(_186_),
    .Y(_187_)
);

FILL FILL_3__8804_ (
);

OR2X2 _10585_ (
    .A(_3849_),
    .B(_3847_),
    .Y(_3851_)
);

OAI21X1 _10165_ (
    .A(_3436_),
    .B(_3443_),
    .C(_3428_),
    .Y(_3444_)
);

FILL FILL_2__6801_ (
);

FILL FILL_2__9693_ (
);

FILL FILL_2__10627_ (
);

FILL FILL_2__9273_ (
);

FILL FILL_0__11661_ (
);

FILL FILL_2__10207_ (
);

FILL FILL_0__11241_ (
);

FILL FILL_2__13099_ (
);

FILL FILL_0__6627_ (
);

NOR2X1 _8733_ (
    .A(_2159_),
    .B(_2163_),
    .Y(_2167_)
);

NAND2X1 _8313_ (
    .A(_1681_),
    .B(_1752_),
    .Y(_1753_)
);

FILL FILL_1__7690_ (
);

FILL FILL_1__7270_ (
);

FILL FILL_0__9099_ (
);

FILL FILL_3__7196_ (
);

FILL FILL_3__12419_ (
);

FILL FILL_1__13033_ (
);

FILL FILL_0__12866_ (
);

NAND3X1 _12731_ (
    .A(_5715_),
    .B(_5764_),
    .C(_5765_),
    .Y(_5771_)
);

FILL FILL_0__12446_ (
);

FILL FILL_0__12026_ (
);

INVX1 _12311_ (
    .A(_5419_),
    .Y(_5420_)
);

OAI22X1 _9938_ (
    .A(_3218_),
    .B(_3219_),
    .C(_3188_),
    .D(_3192_),
    .Y(_3220_)
);

AND2X2 _9518_ (
    .A(_2867_),
    .B(_2873_),
    .Y(_2874_)
);

FILL FILL_1__8895_ (
);

FILL FILL_1__8475_ (
);

FILL FILL_1__8055_ (
);

FILL FILL_2__10380_ (
);

FILL FILL_3__9342_ (
);

FILL FILL_0__6380_ (
);

FILL FILL_2__6398_ (
);

FILL FILL_3__12172_ (
);

FILL FILL_2__11165_ (
);

FILL FILL_1__10998_ (
);

FILL FILL_1__10578_ (
);

FILL FILL_1__10158_ (
);

FILL FILL_0__7585_ (
);

AOI21X1 _9691_ (
    .A(_3031_),
    .B(_3036_),
    .C(_3032_),
    .Y(_3038_)
);

FILL FILL_0__7165_ (
);

OAI21X1 _9271_ (
    .A(_2547_),
    .B(_2551_),
    .C(_2550_),
    .Y(_2630_)
);

FILL FILL_3__10905_ (
);

FILL FILL_2__8544_ (
);

FILL FILL_0__10932_ (
);

FILL FILL_0__10512_ (
);

FILL FILL_1__6961_ (
);

FILL FILL_1__6541_ (
);

FILL FILL_2__13311_ (
);

FILL FILL_3__6467_ (
);

FILL FILL_1__12724_ (
);

FILL FILL_1__12304_ (
);

FILL FILL_0__9731_ (
);

FILL FILL_2__9749_ (
);

FILL FILL_0__9311_ (
);

FILL FILL_2__9329_ (
);

FILL FILL_0__11717_ (
);

FILL FILL_1__7746_ (
);

FILL FILL_1__7326_ (
);

INVX1 _6396_ (
    .A(_787_),
    .Y(_788_)
);

NAND3X1 _10394_ (
    .A(_3668_),
    .B(_3669_),
    .C(_3667_),
    .Y(_3670_)
);

FILL FILL_3__11863_ (
);

FILL FILL_2__6610_ (
);

FILL FILL_3__11023_ (
);

FILL FILL_2__10856_ (
);

FILL FILL_0__11890_ (
);

FILL FILL_2__10436_ (
);

FILL FILL_2__9082_ (
);

FILL FILL_0__11470_ (
);

FILL FILL_2__10016_ (
);

FILL FILL_0__11050_ (
);

FILL FILL_3__9818_ (
);

FILL FILL_0__6856_ (
);

DFFPOSX1 _8962_ (
    .D(_2384_[9]),
    .CLK(clk_bF$buf17),
    .Q(\Y[3] [9])
);

FILL FILL_0__6436_ (
);

OAI21X1 _8542_ (
    .A(_1909_),
    .B(_1978_),
    .C(_1948_),
    .Y(_1979_)
);

DFFPOSX1 _8122_ (
    .D(_1593_[6]),
    .CLK(clk_bF$buf52),
    .Q(\u_fir_pe1.mul [6])
);

DFFPOSX1 _11599_ (
    .D(_4775_[15]),
    .CLK(clk_bF$buf6),
    .Q(\Y[6] [15])
);

OAI21X1 _11179_ (
    .A(_4375_),
    .B(_4374_),
    .C(_4371_),
    .Y(_4376_)
);

FILL FILL_2__7815_ (
);

FILL FILL_3__12648_ (
);

FILL FILL_1__13262_ (
);

OAI21X1 _12960_ (
    .A(_5996_),
    .B(_5898_),
    .C(_5711_),
    .Y(_5997_)
);

FILL FILL_0__12675_ (
);

FILL FILL_0__12255_ (
);

AOI22X1 _12540_ (
    .A(vdd),
    .B(\X[6] [0]),
    .C(vdd),
    .D(\X[6] [1]),
    .Y(_5583_)
);

NOR2X1 _12120_ (
    .A(_5155_),
    .B(_5235_),
    .Y(_5236_)
);

AOI21X1 _9747_ (
    .A(_3086_),
    .B(_3089_),
    .C(_3088_),
    .Y(_3090_)
);

AND2X2 _9327_ (
    .A(_2685_),
    .B(_2681_),
    .Y(_3187_[7])
);

FILL FILL_1__8284_ (
);

FILL FILL_3__9571_ (
);

NAND2X1 _13325_ (
    .A(\u_fir_pe7.rYin [15]),
    .B(\u_fir_pe7.mul [15]),
    .Y(_6348_)
);

FILL FILL_1__9489_ (
);

FILL FILL_1__9069_ (
);

FILL FILL_2__11394_ (
);

FILL FILL_1__10387_ (
);

FILL FILL_0__7394_ (
);

NAND3X1 _9080_ (
    .A(_2431_),
    .B(_2435_),
    .C(_2437_),
    .Y(_2442_)
);

FILL FILL_2__8773_ (
);

FILL FILL_2__8353_ (
);

FILL FILL_0__10321_ (
);

FILL FILL_2__12599_ (
);

FILL FILL_2__12179_ (
);

AOI21X1 _7813_ (
    .A(_1279_),
    .B(_1322_),
    .C(_1325_),
    .Y(_1328_)
);

FILL FILL_1__6770_ (
);

FILL FILL_2__13120_ (
);

FILL FILL_0__8599_ (
);

FILL FILL_3__6696_ (
);

FILL FILL_0__8179_ (
);

FILL FILL_3__11919_ (
);

FILL FILL_1__12953_ (
);

FILL FILL_1__12533_ (
);

FILL FILL_1__12113_ (
);

FILL FILL_2__9978_ (
);

FILL FILL_0__9960_ (
);

FILL FILL_0__9540_ (
);

FILL FILL_2__9558_ (
);

FILL FILL_0__11946_ (
);

FILL FILL_0__9120_ (
);

FILL FILL_2__9138_ (
);

NAND2X1 _11811_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_4931_)
);

FILL FILL_0__11526_ (
);

FILL FILL_0__11106_ (
);

FILL FILL_1__7975_ (
);

FILL FILL_1__7555_ (
);

FILL FILL_1__7135_ (
);

FILL FILL_1__13318_ (
);

FILL FILL_3__8422_ (
);

FILL FILL_3__11672_ (
);

FILL FILL_3__11252_ (
);

FILL FILL_2__10665_ (
);

FILL FILL_2__10245_ (
);

FILL FILL_1__9701_ (
);

FILL FILL_3__9207_ (
);

FILL FILL_0__6665_ (
);

OAI21X1 _8771_ (
    .A(_2185_),
    .B(_2180_),
    .C(_2203_),
    .Y(_2204_)
);

INVX1 _8351_ (
    .A(_1700_),
    .Y(_1791_)
);

FILL FILL_3__12877_ (
);

FILL FILL_2__7624_ (
);

FILL FILL_3__12037_ (
);

FILL FILL_1__13071_ (
);

FILL FILL_0__12064_ (
);

FILL FILL_2__12811_ (
);

OAI21X1 _9976_ (
    .A(_3217_),
    .B(_3251_),
    .C(_3233_),
    .Y(_3257_)
);

NOR2X1 _9556_ (
    .A(_2808_),
    .B(_2853_),
    .Y(_2911_)
);

NAND3X1 _9136_ (
    .A(_2492_),
    .B(_2496_),
    .C(_2460_),
    .Y(_2497_)
);

FILL FILL_1__11804_ (
);

FILL FILL_0__8811_ (
);

FILL FILL_2__8829_ (
);

FILL FILL_2__8409_ (
);

FILL FILL_0__13269_ (
);

INVX1 _13134_ (
    .A(_6164_),
    .Y(_6168_)
);

FILL FILL_1__6826_ (
);

FILL FILL_1__6406_ (
);

FILL FILL_1__9298_ (
);

FILL FILL_2_CLKBUF1_insert90 (
);

FILL FILL_2_CLKBUF1_insert91 (
);

FILL FILL_2_CLKBUF1_insert92 (
);

FILL FILL_2_CLKBUF1_insert93 (
);

FILL FILL_2_CLKBUF1_insert94 (
);

FILL FILL_2_CLKBUF1_insert95 (
);

FILL FILL_2_CLKBUF1_insert96 (
);

FILL FILL_1__10196_ (
);

FILL FILL_3__10523_ (
);

FILL FILL_2__8582_ (
);

FILL FILL_0__10970_ (
);

FILL FILL_2__8162_ (
);

FILL FILL_0__10550_ (
);

FILL FILL_0__10130_ (
);

NAND3X1 _7622_ (
    .A(_1120_),
    .B(_1135_),
    .C(_1136_),
    .Y(_1140_)
);

DFFPOSX1 _7202_ (
    .D(_790_[3]),
    .CLK(clk_bF$buf52),
    .Q(\Y[1] [3])
);

NOR2X1 _10679_ (
    .A(_3942_),
    .B(_3941_),
    .Y(_3943_)
);

NAND3X1 _10259_ (
    .A(_3530_),
    .B(_3531_),
    .C(_3532_),
    .Y(_3537_)
);

FILL FILL_1__12762_ (
);

FILL FILL_1__12342_ (
);

FILL FILL_2__9787_ (
);

FILL FILL_2__9367_ (
);

FILL FILL_0__11755_ (
);

DFFPOSX1 _11620_ (
    .D(\Y[5] [12]),
    .CLK(clk_bF$buf18),
    .Q(\u_fir_pe5.rYin [12])
);

FILL FILL_0__11335_ (
);

NAND2X1 _11200_ (
    .A(vdd),
    .B(\X[5] [7]),
    .Y(_4397_)
);

NOR2X1 _8827_ (
    .A(_2252_),
    .B(_2251_),
    .Y(_2253_)
);

AOI22X1 _8407_ (
    .A(_1681_),
    .B(_1752_),
    .C(_1755_),
    .D(_1751_),
    .Y(_1846_)
);

FILL FILL_1__7784_ (
);

FILL FILL_1__7364_ (
);

FILL FILL_1__13127_ (
);

FILL FILL_3__8651_ (
);

OAI21X1 _12825_ (
    .A(_5863_),
    .B(_5859_),
    .C(_5775_),
    .Y(_5864_)
);

NOR2X1 _12405_ (
    .A(\u_fir_pe6.rYin [10]),
    .B(\u_fir_pe6.mul [10]),
    .Y(_5509_)
);

FILL FILL_1__8569_ (
);

FILL FILL_1__8149_ (
);

FILL FILL_3__11481_ (
);

FILL FILL_2__10894_ (
);

FILL FILL_2__10474_ (
);

FILL FILL_2__10054_ (
);

FILL FILL_1__9930_ (
);

FILL FILL_1__9510_ (
);

FILL FILL_3__9436_ (
);

FILL FILL_0__6894_ (
);

FILL FILL_0__6474_ (
);

NAND3X1 _8580_ (
    .A(_2009_),
    .B(_2016_),
    .C(_1991_),
    .Y(_2017_)
);

NAND3X1 _8160_ (
    .A(_2334_),
    .B(_1602_),
    .C(_1600_),
    .Y(_1603_)
);

FILL FILL_2__7853_ (
);

FILL FILL_2__7433_ (
);

FILL FILL_3__12266_ (
);

FILL FILL_2__7013_ (
);

FILL FILL_2__11679_ (
);

FILL FILL_2__11259_ (
);

FILL FILL_0__12293_ (
);

FILL FILL_2__12620_ (
);

FILL FILL_2__12200_ (
);

FILL FILL_0__7679_ (
);

NOR2X1 _9785_ (
    .A(_3127_),
    .B(_3128_),
    .Y(_3181_[11])
);

FILL FILL_0__7259_ (
);

NAND2X1 _9365_ (
    .A(_2718_),
    .B(_2722_),
    .Y(_2723_)
);

FILL FILL_0__8620_ (
);

FILL FILL_2__8638_ (
);

FILL FILL_0__8200_ (
);

FILL FILL_2__8218_ (
);

FILL FILL_0__10606_ (
);

FILL FILL253650x61350 (
);

FILL FILL_0__13078_ (
);

DFFPOSX1 _13363_ (
    .D(\Y[6] [1]),
    .CLK(clk_bF$buf40),
    .Q(\u_fir_pe7.rYin [1])
);

FILL FILL_1__6635_ (
);

FILL FILL_2__13405_ (
);

FILL FILL_1__12818_ (
);

FILL FILL_0__9825_ (
);

FILL FILL_3__7922_ (
);

FILL FILL_0__9405_ (
);

FILL FILL_3__10332_ (
);

FILL FILL_2__8391_ (
);

FILL FILL_3__8707_ (
);

NOR2X1 _7851_ (
    .A(_1364_),
    .B(_1363_),
    .Y(_1365_)
);

AOI22X1 _7431_ (
    .A(vdd),
    .B(\X[1] [2]),
    .C(vdd),
    .D(\X[1] [3]),
    .Y(_951_)
);

NAND2X1 _7011_ (
    .A(_602_),
    .B(_603_),
    .Y(_604_)
);

INVX1 _10488_ (
    .A(_3759_),
    .Y(_3762_)
);

AOI22X1 _10068_ (
    .A(gnd),
    .B(\X[4] [3]),
    .C(gnd),
    .D(\X[4] [4]),
    .Y(_3348_)
);

FILL FILL_2__6704_ (
);

FILL FILL_1__12991_ (
);

FILL FILL_1__12571_ (
);

FILL FILL_3__11117_ (
);

FILL FILL_1__12151_ (
);

FILL FILL_0__11984_ (
);

FILL FILL_2__9596_ (
);

FILL FILL_2__9176_ (
);

FILL FILL_0__11564_ (
);

FILL FILL_0__11144_ (
);

AND2X2 _8636_ (
    .A(\X[2]_5_bF$buf2 ),
    .B(gnd),
    .Y(_2072_)
);

OAI21X1 _8216_ (
    .A(_1657_),
    .B(_1656_),
    .C(_1623_),
    .Y(_1658_)
);

FILL FILL_1__7593_ (
);

FILL FILL_1__7173_ (
);

FILL FILL_2__7909_ (
);

FILL FILL_3__8880_ (
);

FILL FILL_0__12769_ (
);

NAND3X1 _12634_ (
    .A(_5663_),
    .B(_5674_),
    .C(_5670_),
    .Y(_5675_)
);

FILL FILL_0__12349_ (
);

FILL FILL_3__8040_ (
);

NAND2X1 _12214_ (
    .A(_5324_),
    .B(_5328_),
    .Y(_5329_)
);

FILL FILL_1__8798_ (
);

FILL FILL_1__8378_ (
);

FILL FILL_2__10283_ (
);

FILL FILL_3__9665_ (
);

FILL FILL_2__7662_ (
);

FILL FILL_2__11488_ (
);

FILL FILL_2__11068_ (
);

OAI21X1 _6702_ (
    .A(_210_),
    .B(_220_),
    .C(_216_),
    .Y(_300_)
);

FILL FILL_0__7488_ (
);

NAND3X1 _9594_ (
    .A(_2845_),
    .B(_2947_),
    .C(_2688_),
    .Y(_2948_)
);

FILL FILL_0__7068_ (
);

NAND2X1 _9174_ (
    .A(_2532_),
    .B(_2533_),
    .Y(_2534_)
);

FILL FILL_1__11842_ (
);

FILL FILL_1__11422_ (
);

FILL FILL_1__11002_ (
);

FILL FILL_2__8867_ (
);

FILL FILL_2__8447_ (
);

FILL FILL_0__10835_ (
);

NAND2X1 _10700_ (
    .A(_3962_),
    .B(_3963_),
    .Y(_3978_[15])
);

FILL FILL_0__10415_ (
);

FILL FILL_2__8027_ (
);

NAND2X1 _13172_ (
    .A(_6203_),
    .B(_6167_),
    .Y(_6204_)
);

OAI21X1 _7907_ (
    .A(_1413_),
    .B(_1412_),
    .C(_1418_),
    .Y(_1419_)
);

FILL FILL_1__6864_ (
);

FILL FILL_1__6444_ (
);

FILL FILL_2__13214_ (
);

FILL FILL_1__12627_ (
);

FILL FILL_1__12207_ (
);

FILL FILL_0__9634_ (
);

FILL FILL_0__9214_ (
);

AND2X2 _11905_ (
    .A(vdd),
    .B(\X[7]_5_bF$buf3 ),
    .Y(_5024_)
);

FILL FILL_3__7311_ (
);

FILL FILL_3__10981_ (
);

FILL FILL_1__7649_ (
);

FILL FILL_3__10561_ (
);

FILL FILL_3__10141_ (
);

FILL FILL_3__8516_ (
);

AOI21X1 _7660_ (
    .A(_1094_),
    .B(_1164_),
    .C(_1176_),
    .Y(_1177_)
);

DFFPOSX1 _7240_ (
    .D(_792_[1]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.mul [1])
);

NAND2X1 _10297_ (
    .A(\X[4] [2]),
    .B(gnd),
    .Y(_3574_)
);

FILL FILL_2__6933_ (
);

FILL FILL_3__11766_ (
);

FILL FILL_2__6513_ (
);

FILL FILL_3__11346_ (
);

FILL FILL_1__12380_ (
);

FILL FILL_0__11793_ (
);

FILL FILL_2__10339_ (
);

FILL FILL_0__11373_ (
);

FILL FILL_2__11700_ (
);

FILL FILL_0__6759_ (
);

NAND2X1 _8865_ (
    .A(_2251_),
    .B(_2263_),
    .Y(_2288_)
);

OAI21X1 _8445_ (
    .A(_1801_),
    .B(_1798_),
    .C(_1883_),
    .Y(_1884_)
);

OAI21X1 _8025_ (
    .A(_1521_),
    .B(_1522_),
    .C(_1526_),
    .Y(_1529_)
);

FILL FILL_0__7700_ (
);

FILL FILL_2__7718_ (
);

FILL FILL_1__13165_ (
);

FILL FILL_0__12998_ (
);

OAI21X1 _12863_ (
    .A(_5897_),
    .B(_5900_),
    .C(_5899_),
    .Y(_5901_)
);

FILL FILL_0__12578_ (
);

FILL FILL_0__12158_ (
);

AND2X2 _12443_ (
    .A(_5540_),
    .B(_5546_),
    .Y(_5547_)
);

AOI21X1 _12023_ (
    .A(_5052_),
    .B(_5054_),
    .C(_5140_),
    .Y(_5141_)
);

FILL FILL_2__12905_ (
);

FILL FILL_1__8187_ (
);

FILL FILL_0__8905_ (
);

FILL FILL_2__10092_ (
);

FILL FILL_3__9894_ (
);

FILL FILL_3__9054_ (
);

INVX1 _13228_ (
    .A(\u_fir_pe7.rYin [6]),
    .Y(_6252_)
);

FILL FILL_2__7891_ (
);

FILL FILL_2__7471_ (
);

FILL FILL_2__7051_ (
);

FILL FILL_2__11297_ (
);

NAND2X1 _6931_ (
    .A(gnd),
    .B(Xin[7]),
    .Y(_526_)
);

INVX1 _6511_ (
    .A(_26_),
    .Y(_112_)
);

FILL FILL_0__7297_ (
);

FILL FILL_3__10617_ (
);

FILL FILL_1__11651_ (
);

FILL FILL_1__11231_ (
);

FILL FILL_2__8676_ (
);

FILL FILL_2__8256_ (
);

FILL FILL_0__10644_ (
);

FILL FILL_3__13089_ (
);

FILL FILL_0__10224_ (
);

OAI21X1 _7716_ (
    .A(_1232_),
    .B(_1231_),
    .C(_1230_),
    .Y(_1233_)
);

FILL FILL_1__6673_ (
);

FILL FILL_2__13023_ (
);

FILL FILL_1__12856_ (
);

FILL FILL_1__12436_ (
);

FILL FILL_1__12016_ (
);

FILL FILL_3__7960_ (
);

FILL FILL_0__9443_ (
);

FILL FILL_0__11849_ (
);

FILL FILL_3__7540_ (
);

FILL FILL_0__9023_ (
);

INVX1 _11714_ (
    .A(_4835_),
    .Y(_4836_)
);

FILL FILL_0__11429_ (
);

FILL FILL_3__7120_ (
);

FILL FILL_0__11009_ (
);

FILL FILL_1__7878_ (
);

FILL FILL_1__7458_ (
);

FILL FILL_1__7038_ (
);

FILL FILL_3__8745_ (
);

NAND2X1 _12919_ (
    .A(_5956_),
    .B(_5955_),
    .Y(_5957_)
);

FILL FILL_3__8325_ (
);

FILL FILL_2__6742_ (
);

FILL FILL_3__11575_ (
);

FILL FILL_2__10988_ (
);

FILL FILL_2__10568_ (
);

FILL FILL_2__10148_ (
);

FILL FILL_0__11182_ (
);

FILL FILL_1__9604_ (
);

FILL FILL_0__6988_ (
);

FILL FILL_0__6568_ (
);

NAND2X1 _8674_ (
    .A(_2062_),
    .B(_2063_),
    .Y(_2109_)
);

NAND3X1 _8254_ (
    .A(_1690_),
    .B(_1676_),
    .C(_1694_),
    .Y(_1695_)
);

FILL FILL_1__10922_ (
);

FILL FILL_1__10502_ (
);

FILL FILL_2__7947_ (
);

FILL FILL_2__7527_ (
);

FILL FILL_2__7107_ (
);

FILL FILL_1__13394_ (
);

OAI21X1 _12672_ (
    .A(_6289_),
    .B(_5711_),
    .C(_5656_),
    .Y(_5712_)
);

FILL FILL_0__12387_ (
);

OR2X2 _12252_ (
    .A(_5365_),
    .B(_5342_),
    .Y(_5366_)
);

FILL FILL_2__12714_ (
);

FILL FILL254250x165750 (
);

DFFPOSX1 _9879_ (
    .D(_3187_[9]),
    .CLK(clk_bF$buf4),
    .Q(\u_fir_pe3.mul [9])
);

NAND3X1 _9459_ (
    .A(_2734_),
    .B(_2740_),
    .C(_2815_),
    .Y(_2816_)
);

NAND3X1 _9039_ (
    .A(_2391_),
    .B(_2396_),
    .C(_2394_),
    .Y(_2402_)
);

FILL FILL_1__11707_ (
);

FILL FILL_0__8714_ (
);

FILL FILL_3__9283_ (
);

NAND3X1 _13037_ (
    .A(_6002_),
    .B(_6005_),
    .C(_6072_),
    .Y(_6073_)
);

FILL FILL_1__6729_ (
);

FILL FILL_2__7280_ (
);

FILL FILL_0__9919_ (
);

NAND3X1 _6740_ (
    .A(_330_),
    .B(_334_),
    .C(_332_),
    .Y(_338_)
);

FILL FILL_1__10099_ (
);

FILL FILL_3__10846_ (
);

FILL FILL_1__11880_ (
);

FILL FILL_1__11460_ (
);

FILL FILL_3__10006_ (
);

FILL FILL_1__11040_ (
);

FILL FILL_2__8485_ (
);

FILL FILL_0__10873_ (
);

FILL FILL_0__10453_ (
);

FILL FILL_2__8065_ (
);

FILL FILL_0__10033_ (
);

NAND2X1 _7945_ (
    .A(_1450_),
    .B(_1451_),
    .Y(_1587_[3])
);

NAND2X1 _7525_ (
    .A(_955_),
    .B(_1039_),
    .Y(_1044_)
);

NAND2X1 _7105_ (
    .A(_687_),
    .B(_686_),
    .Y(_688_)
);

FILL FILL_1__6482_ (
);

FILL FILL_2__13252_ (
);

FILL FILL_1__12665_ (
);

FILL FILL_1__12245_ (
);

FILL FILL_0__9672_ (
);

FILL FILL_0__9252_ (
);

AOI21X1 _11943_ (
    .A(_5061_),
    .B(_5056_),
    .C(_4917_),
    .Y(_5062_)
);

FILL FILL_0__11658_ (
);

AOI21X1 _11523_ (
    .A(_4688_),
    .B(_4703_),
    .C(_4706_),
    .Y(_4707_)
);

FILL FILL_0__11238_ (
);

AOI21X1 _11103_ (
    .A(_4241_),
    .B(_4238_),
    .C(_4224_),
    .Y(_4301_)
);

FILL FILL_1__7687_ (
);

FILL FILL_1__7267_ (
);

AOI21X1 _12728_ (
    .A(_5680_),
    .B(_5684_),
    .C(_5648_),
    .Y(_5768_)
);

NOR2X1 _12308_ (
    .A(\u_fir_pe6.rYin [1]),
    .B(\u_fir_pe6.mul [1]),
    .Y(_5417_)
);

FILL FILL_2__6971_ (
);

FILL FILL_2__6551_ (
);

FILL FILL_2__10797_ (
);

FILL FILL_2__10377_ (
);

FILL FILL_1__9413_ (
);

FILL FILL_3__9759_ (
);

FILL FILL_0__6797_ (
);

AND2X2 _8483_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf0 ),
    .Y(_1921_)
);

NAND2X1 _8063_ (
    .A(\u_fir_pe1.rYin [15]),
    .B(\u_fir_pe1.mul [15]),
    .Y(_1566_)
);

FILL FILL_1__10311_ (
);

FILL FILL_2__7756_ (
);

FILL FILL_3__12589_ (
);

FILL FILL_2__7336_ (
);

FILL FILL_0__12196_ (
);

DFFPOSX1 _12481_ (
    .D(\X[7] [4]),
    .CLK(clk_bF$buf29),
    .Q(_6376_[4])
);

AOI21X1 _12061_ (
    .A(_5121_),
    .B(_5120_),
    .C(_5105_),
    .Y(_5178_)
);

FILL FILL_3__13110_ (
);

FILL FILL_2__12943_ (
);

FILL FILL_2__12523_ (
);

FILL FILL_2__12103_ (
);

NOR2X1 _9688_ (
    .A(_3033_),
    .B(_3032_),
    .Y(_3036_)
);

OAI21X1 _9268_ (
    .A(_3169_),
    .B(_2626_),
    .C(_2618_),
    .Y(_2627_)
);

FILL FILL_1__11936_ (
);

FILL FILL_1__11516_ (
);

FILL FILL_0__8943_ (
);

FILL FILL_0__8523_ (
);

FILL FILL_0__10929_ (
);

FILL FILL_3__6620_ (
);

FILL FILL_0__10509_ (
);

OAI21X1 _13266_ (
    .A(_6288_),
    .B(_6285_),
    .C(_6287_),
    .Y(_6290_)
);

FILL FILL_2__9902_ (
);

FILL FILL_1__6958_ (
);

FILL FILL_1__6538_ (
);

FILL FILL_2__13308_ (
);

FILL FILL_0__9728_ (
);

FILL FILL_0__9308_ (
);

FILL FILL_3__7405_ (
);

FILL FILL_3__10655_ (
);

FILL FILL_3__10235_ (
);

FILL FILL_2__8294_ (
);

FILL FILL_0__10682_ (
);

FILL FILL_0__10262_ (
);

NAND2X1 _7754_ (
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_1270_)
);

OAI21X1 _7334_ (
    .A(_1578_),
    .B(_815_),
    .C(_818_),
    .Y(_856_)
);

FILL FILL_2__13061_ (
);

FILL FILL_2__6607_ (
);

FILL FILL_1__12894_ (
);

FILL FILL_1__12054_ (
);

FILL FILL_0__9481_ (
);

FILL FILL_2__9499_ (
);

FILL FILL_0__11887_ (
);

FILL FILL_2__9079_ (
);

FILL FILL_0__9061_ (
);

NAND3X1 _11752_ (
    .A(_4868_),
    .B(_4872_),
    .C(_4870_),
    .Y(_4873_)
);

FILL FILL_0__11467_ (
);

FILL FILL253650x241350 (
);

FILL FILL_0__11047_ (
);

NAND3X1 _11332_ (
    .A(_4500_),
    .B(_4526_),
    .C(_4522_),
    .Y(_4527_)
);

FILL FILL_3__12801_ (
);

DFFPOSX1 _8959_ (
    .D(_2384_[6]),
    .CLK(clk_bF$buf53),
    .Q(\Y[3] [6])
);

OAI21X1 _8539_ (
    .A(_1895_),
    .B(_1975_),
    .C(_1958_),
    .Y(_1976_)
);

DFFPOSX1 _8119_ (
    .D(_1591_[3]),
    .CLK(clk_bF$buf43),
    .Q(\u_fir_pe1.mul [3])
);

FILL FILL_1__7496_ (
);

FILL FILL_1__7076_ (
);

NOR2X1 _9900_ (
    .A(_3971_),
    .B(_3970_),
    .Y(_3972_)
);

FILL FILL_1__13259_ (
);

NAND3X1 _12957_ (
    .A(_5979_),
    .B(_5986_),
    .C(_5993_),
    .Y(_5994_)
);

FILL FILL_3__8363_ (
);

INVX1 _12537_ (
    .A(_5579_),
    .Y(_5580_)
);

NAND2X1 _12117_ (
    .A(_5232_),
    .B(_5162_),
    .Y(_5234_)
);

FILL FILL_2__6780_ (
);

FILL FILL_3__11193_ (
);

FILL FILL_2__10186_ (
);

FILL FILL_1__9642_ (
);

FILL FILL_1__9222_ (
);

FILL FILL_3__9988_ (
);

FILL FILL_3__9148_ (
);

OAI21X1 _8292_ (
    .A(_1696_),
    .B(_1731_),
    .C(_1690_),
    .Y(_1732_)
);

FILL FILL_1__10960_ (
);

FILL FILL_1__10540_ (
);

FILL FILL_1__10120_ (
);

FILL FILL_2__7985_ (
);

FILL FILL_2__7565_ (
);

FILL FILL_2__7145_ (
);

NAND2X1 _12290_ (
    .A(_5400_),
    .B(_5399_),
    .Y(_5402_)
);

OAI21X1 _6605_ (
    .A(_129_),
    .B(_127_),
    .C(_120_),
    .Y(_205_)
);

FILL FILL_2__12752_ (
);

FILL FILL_2__12332_ (
);

INVX2 _9497_ (
    .A(gnd),
    .Y(_2853_)
);

NAND2X1 _9077_ (
    .A(_2437_),
    .B(_2438_),
    .Y(_2439_)
);

FILL FILL_1__11745_ (
);

FILL FILL_1__11325_ (
);

FILL FILL_0__8752_ (
);

FILL FILL_0__8332_ (
);

FILL FILL_0__10318_ (
);

OR2X2 _10603_ (
    .A(_3860_),
    .B(_3865_),
    .Y(_3867_)
);

AOI21X1 _13075_ (
    .A(_6061_),
    .B(_6104_),
    .C(_6107_),
    .Y(_6110_)
);

FILL FILL_2__9711_ (
);

FILL FILL_1__6767_ (
);

FILL FILL_2__13117_ (
);

FILL FILL_0__9957_ (
);

FILL FILL_0__9537_ (
);

FILL FILL_3__7634_ (
);

FILL FILL_0__9117_ (
);

OAI21X1 _11808_ (
    .A(_5560_),
    .B(_4926_),
    .C(_4927_),
    .Y(_4928_)
);

FILL FILL253950x7350 (
);

FILL FILL_0__10491_ (
);

FILL FILL_0__10071_ (
);

FILL FILL_1__8913_ (
);

FILL FILL_3__8839_ (
);

FILL FILL_3__8419_ (
);

NAND2X1 _7983_ (
    .A(_1482_),
    .B(_1485_),
    .Y(_1587_[7])
);

OAI21X1 _7563_ (
    .A(_1081_),
    .B(_1077_),
    .C(_993_),
    .Y(_1082_)
);

NOR2X1 _7143_ (
    .A(\u_fir_pe0.rYin [10]),
    .B(\u_fir_pe0.mul [10]),
    .Y(_727_)
);

FILL FILL_2__13290_ (
);

FILL FILL_2__6836_ (
);

FILL FILL_2__6416_ (
);

FILL FILL_1__12283_ (
);

FILL FILL254550x144150 (
);

FILL FILL_0__9290_ (
);

OAI21X1 _11981_ (
    .A(_5020_),
    .B(_5098_),
    .C(_5042_),
    .Y(_5099_)
);

FILL FILL_0__11696_ (
);

INVX1 _11561_ (
    .A(\u_fir_pe5.rYin [14]),
    .Y(_4744_)
);

FILL FILL_0__11276_ (
);

NAND3X1 _11141_ (
    .A(_4334_),
    .B(_4335_),
    .C(_4302_),
    .Y(_4339_)
);

FILL FILL_3__12610_ (
);

AND2X2 _8768_ (
    .A(_2197_),
    .B(_2196_),
    .Y(_2201_)
);

OAI21X1 _8348_ (
    .A(_1787_),
    .B(_1782_),
    .C(_1710_),
    .Y(_1788_)
);

FILL FILL_0__7603_ (
);

FILL FILL_1__13068_ (
);

FILL FILL_3__8592_ (
);

INVX1 _12766_ (
    .A(_5804_),
    .Y(_5805_)
);

NOR2X1 _12346_ (
    .A(_5450_),
    .B(_5449_),
    .Y(_5451_)
);

FILL FILL_2__12808_ (
);

FILL FILL_0__13002_ (
);

FILL FILL_0__8808_ (
);

FILL FILL_1__9451_ (
);

FILL FILL_1__9031_ (
);

FILL FILL_3__9377_ (
);

FILL FILL_2__7794_ (
);

FILL FILL_2__7374_ (
);

NAND3X1 _6834_ (
    .A(_426_),
    .B(_430_),
    .C(_385_),
    .Y(_431_)
);

OAI21X1 _6414_ (
    .A(_778_),
    .B(_15_),
    .C(_16_),
    .Y(_17_)
);

FILL FILL_2__12981_ (
);

FILL FILL_2__12561_ (
);

FILL FILL_2__12141_ (
);

FILL FILL_1__11974_ (
);

FILL FILL_1__11554_ (
);

FILL FILL_1__11134_ (
);

FILL FILL253950x100950 (
);

FILL FILL_2__8579_ (
);

FILL FILL_0__8561_ (
);

FILL FILL_0__10967_ (
);

FILL FILL_0__8141_ (
);

FILL FILL_2__8159_ (
);

FILL FILL_0__10547_ (
);

NAND3X1 _10832_ (
    .A(_4014_),
    .B(_4030_),
    .C(_4033_),
    .Y(_4034_)
);

NAND2X1 _10412_ (
    .A(_3686_),
    .B(_3687_),
    .Y(_3688_)
);

FILL FILL_0__10127_ (
);

FILL FILL_2__9940_ (
);

FILL FILL_2__9520_ (
);

FILL FILL_2__9100_ (
);

NAND3X1 _7619_ (
    .A(_1135_),
    .B(_1136_),
    .C(_1134_),
    .Y(_1137_)
);

FILL FILL_1__6996_ (
);

FILL FILL_1__6576_ (
);

FILL FILL_1__12759_ (
);

FILL FILL_1__12339_ (
);

FILL FILL_0__9766_ (
);

FILL FILL_3__7863_ (
);

FILL FILL_0__9346_ (
);

DFFPOSX1 _11617_ (
    .D(\Y[5] [9]),
    .CLK(clk_bF$buf35),
    .Q(\u_fir_pe5.rYin [9])
);

FILL FILL_3__10273_ (
);

FILL FILL_1__8722_ (
);

FILL FILL_1__8302_ (
);

NOR2X1 _7792_ (
    .A(_1304_),
    .B(_1307_),
    .Y(_1593_[10])
);

NAND3X1 _7372_ (
    .A(_881_),
    .B(_892_),
    .C(_888_),
    .Y(_893_)
);

FILL FILL_3__11898_ (
);

FILL FILL_2__6645_ (
);

FILL FILL_3__11058_ (
);

FILL FILL_1__12092_ (
);

INVX1 _11790_ (
    .A(_4907_),
    .Y(_4911_)
);

FILL FILL_0__11085_ (
);

AOI21X1 _11370_ (
    .A(_4562_),
    .B(_4563_),
    .C(_4546_),
    .Y(_4564_)
);

FILL FILL_1__9927_ (
);

FILL FILL_1__9507_ (
);

FILL FILL_2__11832_ (
);

FILL FILL_2__11412_ (
);

DFFPOSX1 _8997_ (
    .D(_2389_[4]),
    .CLK(clk_bF$buf53),
    .Q(\u_fir_pe2.mul [4])
);

NAND2X1 _8577_ (
    .A(_1997_),
    .B(_2007_),
    .Y(_2014_)
);

NAND3X1 _8157_ (
    .A(_1595_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1600_)
);

FILL FILL_1__10825_ (
);

FILL FILL_1__10405_ (
);

FILL FILL_0__7832_ (
);

FILL FILL_0__7412_ (
);

FILL FILL_1__13297_ (
);

NAND2X1 _12995_ (
    .A(_6031_),
    .B(_6030_),
    .Y(_6375_[9])
);

AOI22X1 _12575_ (
    .A(vdd),
    .B(\X[6] [1]),
    .C(vdd),
    .D(\X[6] [2]),
    .Y(_5617_)
);

NAND2X1 _12155_ (
    .A(_5267_),
    .B(_5254_),
    .Y(_5271_)
);

FILL FILL_3__13204_ (
);

FILL FILL_2__12617_ (
);

FILL FILL_0__13231_ (
);

FILL FILL_0__8617_ (
);

FILL FILL_3__6714_ (
);

FILL FILL_1__9680_ (
);

FILL FILL_1__9260_ (
);

FILL FILL_2__7183_ (
);

AND2X2 _6643_ (
    .A(vdd),
    .B(Xin_5_bF$buf2),
    .Y(_242_)
);

FILL FILL_2__12790_ (
);

FILL FILL_2__12370_ (
);

FILL FILL_1__11783_ (
);

FILL FILL_3__10329_ (
);

FILL FILL_1__11363_ (
);

FILL FILL_0__8790_ (
);

FILL FILL_2__8388_ (
);

FILL FILL_0__8370_ (
);

FILL FILL_0__10776_ (
);

FILL FILL_0__10356_ (
);

OAI21X1 _10641_ (
    .A(_3900_),
    .B(_3901_),
    .C(_3899_),
    .Y(_3905_)
);

INVX1 _10221_ (
    .A(_3492_),
    .Y(_3499_)
);

NOR2X1 _7848_ (
    .A(_871_),
    .B(_1259_),
    .Y(_1362_)
);

NAND3X1 _7428_ (
    .A(_936_),
    .B(_945_),
    .C(_947_),
    .Y(_948_)
);

NAND2X1 _7008_ (
    .A(_599_),
    .B(_600_),
    .Y(_601_)
);

FILL FILL_1__6385_ (
);

FILL FILL_2__13155_ (
);

FILL FILL_1__12988_ (
);

FILL FILL_1__12568_ (
);

FILL FILL_1__12148_ (
);

FILL FILL_0__9995_ (
);

FILL FILL_0__9575_ (
);

FILL FILL_0__9155_ (
);

AND2X2 _11846_ (
    .A(_4916_),
    .B(_4917_),
    .Y(_4966_)
);

INVX1 _11426_ (
    .A(_4009_),
    .Y(_4776_[0])
);

NOR2X1 _11006_ (
    .A(_4198_),
    .B(_4200_),
    .Y(_4205_)
);

FILL FILL_0__12922_ (
);

FILL FILL_1__8951_ (
);

FILL FILL_1__8531_ (
);

FILL FILL_3__8457_ (
);

AND2X2 _7181_ (
    .A(_758_),
    .B(_764_),
    .Y(_765_)
);

FILL FILL_2__6874_ (
);

FILL FILL_2__6454_ (
);

FILL FILL_3__11287_ (
);

FILL FILL_1__9736_ (
);

FILL FILL_1__9316_ (
);

FILL FILL_2__11641_ (
);

FILL FILL_2__11221_ (
);

INVX1 _8386_ (
    .A(_1824_),
    .Y(_1825_)
);

FILL FILL_1__10634_ (
);

FILL FILL_1__10214_ (
);

FILL FILL_2__7659_ (
);

FILL FILL_0__7641_ (
);

FILL FILL_0__12099_ (
);

INVX1 _12384_ (
    .A(_5485_),
    .Y(_5488_)
);

FILL FILL_2__8600_ (
);

FILL FILL_2__12846_ (
);

FILL FILL_2__12426_ (
);

FILL FILL_2__12006_ (
);

FILL FILL_0__13040_ (
);

FILL FILL_1__11839_ (
);

FILL FILL_1__11419_ (
);

FILL FILL_0__8846_ (
);

FILL FILL_3__6943_ (
);

FILL FILL_0__8426_ (
);

FILL FILL_0__8006_ (
);

OAI21X1 _13169_ (
    .A(_6195_),
    .B(_6194_),
    .C(_6200_),
    .Y(_6201_)
);

FILL FILL_2__9805_ (
);

FILL FILL_1__7802_ (
);

FILL FILL_3__7728_ (
);

NAND2X1 _6872_ (
    .A(gnd),
    .B(_398_),
    .Y(_468_)
);

INVX1 _6452_ (
    .A(_53_),
    .Y(_54_)
);

FILL FILL_3__10558_ (
);

FILL FILL_1__11172_ (
);

FILL FILL_2__8197_ (
);

FILL FILL_0__10585_ (
);

INVX1 _10870_ (
    .A(_4070_),
    .Y(_4071_)
);

NAND2X1 _10450_ (
    .A(_3724_),
    .B(_3704_),
    .Y(_3725_)
);

FILL FILL_0__10165_ (
);

NAND3X1 _10030_ (
    .A(_3242_),
    .B(_3299_),
    .C(_3303_),
    .Y(_3311_)
);

BUFX2 BUFX2_insert70 (
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf3 )
);

BUFX2 BUFX2_insert71 (
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf2 )
);

BUFX2 BUFX2_insert72 (
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf1 )
);

BUFX2 BUFX2_insert73 (
    .A(\X[2] [5]),
    .Y(\X[2]_5_bF$buf0 )
);

BUFX2 BUFX2_insert74 (
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf3 )
);

BUFX2 BUFX2_insert75 (
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf2 )
);

BUFX2 BUFX2_insert76 (
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf1 )
);

BUFX2 BUFX2_insert77 (
    .A(\X[4] [5]),
    .Y(\X[4]_5_bF$buf0 )
);

FILL FILL_2__10912_ (
);

BUFX2 BUFX2_insert78 (
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf3 )
);

BUFX2 BUFX2_insert79 (
    .A(\X[6] [5]),
    .Y(\X[6]_5_bF$buf2 )
);

NAND2X1 _7657_ (
    .A(_1174_),
    .B(_1173_),
    .Y(_1175_)
);

DFFPOSX1 _7237_ (
    .D(Yin[14]),
    .CLK(clk_bF$buf41),
    .Q(\u_fir_pe0.rYin [14])
);

FILL FILL_0__6912_ (
);

FILL FILL_1__12797_ (
);

FILL FILL_1__12377_ (
);

FILL FILL_0__9384_ (
);

FILL FILL_3__7481_ (
);

NAND2X1 _11655_ (
    .A(_5502_),
    .B(_5566_),
    .Y(_5567_)
);

FILL FILL_3__7061_ (
);

AOI21X1 _11235_ (
    .A(_4431_),
    .B(_4430_),
    .C(_4423_),
    .Y(_4432_)
);

FILL FILL_3__12704_ (
);

FILL FILL_0__12731_ (
);

FILL FILL_0__12311_ (
);

FILL FILL_1__7399_ (
);

NAND2X1 _9803_ (
    .A(_3146_),
    .B(_3140_),
    .Y(_3147_)
);

FILL FILL_1__8760_ (
);

FILL FILL_1__8340_ (
);

FILL FILL_3__8686_ (
);

FILL FILL_3__8266_ (
);

FILL FILL_2__6683_ (
);

FILL FILL_2__10089_ (
);

FILL FILL_1__9965_ (
);

FILL FILL_1__9545_ (
);

FILL FILL_1__9125_ (
);

FILL FILL_2__11870_ (
);

FILL FILL_2__11450_ (
);

FILL FILL_2__11030_ (
);

NAND3X1 _8195_ (
    .A(vdd),
    .B(\X[2] [1]),
    .C(_1636_),
    .Y(_1637_)
);

FILL FILL_1__10863_ (
);

FILL FILL_1__10443_ (
);

FILL FILL_1__10023_ (
);

FILL FILL_2__7888_ (
);

FILL FILL_0__7870_ (
);

FILL FILL_2__7468_ (
);

FILL FILL_0__7450_ (
);

FILL FILL_2__7048_ (
);

FILL FILL_0__7030_ (
);

NAND2X1 _12193_ (
    .A(gnd),
    .B(\X[7] [7]),
    .Y(_5308_)
);

FILL FILL_3__13242_ (
);

NAND3X1 _6928_ (
    .A(_520_),
    .B(_521_),
    .C(_522_),
    .Y(_523_)
);

AOI21X1 _6508_ (
    .A(_100_),
    .B(_96_),
    .C(_82_),
    .Y(_109_)
);

FILL FILL_2__12655_ (
);

FILL FILL_2__12235_ (
);

FILL FILL_1__11648_ (
);

FILL FILL_1__11228_ (
);

FILL FILL_0__8655_ (
);

FILL FILL_0__8235_ (
);

AND2X2 _10926_ (
    .A(\X[5] [2]),
    .B(vdd),
    .Y(_4126_)
);

NOR2X1 _10506_ (
    .A(_3748_),
    .B(_3771_),
    .Y(_3779_)
);

BUFX2 _13398_ (
    .A(_6376_[4]),
    .Y(Xout[4])
);

FILL FILL_2__9614_ (
);

FILL FILL_1__7611_ (
);

FILL FILL_3__7957_ (
);

FILL FILL_3__7117_ (
);

AOI21X1 _6681_ (
    .A(_279_),
    .B(_274_),
    .C(_135_),
    .Y(_280_)
);

FILL FILL_3__10787_ (
);

FILL FILL_0__10394_ (
);

FILL FILL_1__8816_ (
);

FILL FILL_2__10301_ (
);

NAND2X1 _7886_ (
    .A(_1391_),
    .B(_1398_),
    .Y(_1399_)
);

AOI21X1 _7466_ (
    .A(_898_),
    .B(_902_),
    .C(_866_),
    .Y(_986_)
);

NOR2X1 _7046_ (
    .A(\u_fir_pe0.rYin [1]),
    .B(\u_fir_pe0.mul [1]),
    .Y(_635_)
);

FILL FILL_2__13193_ (
);

FILL FILL_0__6721_ (
);

FILL FILL_2__6739_ (
);

FILL FILL_1__12186_ (
);

FILL FILL_0__9193_ (
);

OAI21X1 _11884_ (
    .A(_5001_),
    .B(_5002_),
    .C(_4992_),
    .Y(_5003_)
);

OAI21X1 _11464_ (
    .A(_4640_),
    .B(_4641_),
    .C(_4647_),
    .Y(_4649_)
);

FILL FILL_0__11179_ (
);

AOI21X1 _11044_ (
    .A(_4236_),
    .B(_4242_),
    .C(_4223_),
    .Y(_4243_)
);

FILL FILL_2__11926_ (
);

FILL FILL_0__12960_ (
);

FILL FILL_2__11506_ (
);

FILL FILL_0__12540_ (
);

FILL FILL_0__12120_ (
);

FILL FILL_1__10919_ (
);

FILL FILL_0__7926_ (
);

FILL FILL_0__7506_ (
);

OAI21X1 _9612_ (
    .A(_2964_),
    .B(_2965_),
    .C(_2917_),
    .Y(_2966_)
);

AND2X2 _12669_ (
    .A(_5709_),
    .B(_5705_),
    .Y(_6375_[5])
);

FILL FILL_3__8075_ (
);

INVX1 _12249_ (
    .A(_5362_),
    .Y(_5363_)
);

FILL FILL_0__13325_ (
);

FILL FILL_2__6492_ (
);

FILL FILL_3__6808_ (
);

FILL FILL_1__9774_ (
);

FILL FILL_1__9354_ (
);

FILL FILL_1__10672_ (
);

FILL FILL_1__10252_ (
);

FILL FILL_2__7697_ (
);

FILL FILL_2__7277_ (
);

FILL FILL_3__13051_ (
);

AOI21X1 _6737_ (
    .A(_332_),
    .B(_334_),
    .C(_330_),
    .Y(_335_)
);

FILL FILL_2__12884_ (
);

FILL FILL_2__12044_ (
);

FILL FILL_1__11877_ (
);

FILL FILL_1__11457_ (
);

FILL FILL_1__11037_ (
);

FILL FILL_0__8884_ (
);

FILL FILL_0__8464_ (
);

FILL FILL_3__6561_ (
);

DFFPOSX1 _10735_ (
    .D(\Y[4] [4]),
    .CLK(clk_bF$buf38),
    .Q(\u_fir_pe4.rYin [4])
);

FILL FILL_0__8044_ (
);

AOI22X1 _10315_ (
    .A(gnd),
    .B(\X[4] [6]),
    .C(gnd),
    .D(\X[4] [7]),
    .Y(_3592_)
);

FILL FILL_2__9423_ (
);

FILL FILL_0__11811_ (
);

FILL FILL_1__6899_ (
);

FILL FILL_1__6479_ (
);

FILL FILL_2__13249_ (
);

FILL FILL_3_CLKBUF1_insert50 (
);

FILL FILL_3_CLKBUF1_insert52 (
);

FILL FILL_3_CLKBUF1_insert54 (
);

FILL FILL_3_CLKBUF1_insert56 (
);

FILL FILL_1__7840_ (
);

FILL FILL_1__7420_ (
);

FILL FILL_3_CLKBUF1_insert58 (
);

FILL FILL_1__7000_ (
);

FILL FILL_0__9669_ (
);

FILL FILL_0__9249_ (
);

FILL FILL_3__7346_ (
);

NAND3X1 _6490_ (
    .A(_86_),
    .B(_90_),
    .C(_88_),
    .Y(_91_)
);

FILL FILL_3__10596_ (
);

FILL FILL_3__10176_ (
);

FILL FILL_1__8625_ (
);

FILL FILL_1__8205_ (
);

FILL FILL_2__10950_ (
);

FILL FILL_2__10530_ (
);

FILL FILL_2__10110_ (
);

NAND3X1 _7695_ (
    .A(_1197_),
    .B(_1204_),
    .C(_1211_),
    .Y(_1212_)
);

INVX1 _7275_ (
    .A(_797_),
    .Y(_798_)
);

FILL FILL_2__6968_ (
);

FILL FILL_0__6950_ (
);

FILL FILL_2__6548_ (
);

FILL FILL_0__6530_ (
);

NAND2X1 _11693_ (
    .A(gnd),
    .B(\X[7] [3]),
    .Y(_4815_)
);

NAND2X1 _11273_ (
    .A(_4468_),
    .B(_4457_),
    .Y(_4469_)
);

FILL FILL_3__12742_ (
);

FILL FILL_2__11735_ (
);

FILL FILL_2__11315_ (
);

FILL FILL_1__10308_ (
);

FILL FILL_0__7735_ (
);

DFFPOSX1 _9841_ (
    .D(_3181_[11]),
    .CLK(clk_bF$buf17),
    .Q(\Y[4] [11])
);

FILL FILL_0__7315_ (
);

NOR2X1 _9421_ (
    .A(_2709_),
    .B(_2712_),
    .Y(_2778_)
);

DFFPOSX1 _9001_ (
    .D(_2390_[8]),
    .CLK(clk_bF$buf53),
    .Q(\u_fir_pe2.mul [8])
);

OAI21X1 _12898_ (
    .A(_5935_),
    .B(_5931_),
    .C(_5882_),
    .Y(_5936_)
);

DFFPOSX1 _12478_ (
    .D(\X[7] [1]),
    .CLK(clk_bF$buf29),
    .Q(_6376_[1])
);

INVX1 _12058_ (
    .A(_5172_),
    .Y(_5175_)
);

FILL FILL_0__13134_ (
);

FILL FILL_1__9583_ (
);

FILL FILL_1__9163_ (
);

FILL FILL_3__9089_ (
);

FILL FILL_1__10481_ (
);

FILL FILL_1__10061_ (
);

FILL FILL_2__7086_ (
);

AND2X2 _6966_ (
    .A(_542_),
    .B(_537_),
    .Y(_560_)
);

OAI21X1 _6546_ (
    .A(_778_),
    .B(_144_),
    .C(_145_),
    .Y(_146_)
);

FILL FILL_2__12693_ (
);

FILL FILL_2__12273_ (
);

FILL FILL_1__11686_ (
);

FILL FILL_1__11266_ (
);

FILL FILL_0__8693_ (
);

FILL FILL_3__6790_ (
);

FILL FILL_0__8273_ (
);

FILL FILL_0__10679_ (
);

AOI21X1 _10964_ (
    .A(_4067_),
    .B(_4085_),
    .C(_4163_),
    .Y(_4164_)
);

NAND3X1 _10544_ (
    .A(_3814_),
    .B(_3815_),
    .C(_3813_),
    .Y(_3816_)
);

FILL FILL_0__10259_ (
);

OAI21X1 _10124_ (
    .A(_3327_),
    .B(_3402_),
    .C(_3331_),
    .Y(_3403_)
);

FILL FILL_2__9652_ (
);

FILL FILL_2__9232_ (
);

FILL FILL_0__11200_ (
);

FILL FILL_2__13058_ (
);

FILL FILL_3__7995_ (
);

FILL FILL_0__9898_ (
);

FILL FILL_0__9478_ (
);

FILL FILL_3__7575_ (
);

FILL FILL_0__9058_ (
);

NAND2X1 _11749_ (
    .A(_4818_),
    .B(_4869_),
    .Y(_4870_)
);

FILL FILL_3__7155_ (
);

AOI21X1 _11329_ (
    .A(_4455_),
    .B(_4471_),
    .C(_4523_),
    .Y(_4524_)
);

FILL FILL_1__13412_ (
);

FILL FILL_0__12825_ (
);

FILL FILL_0__12405_ (
);

FILL FILL_1__8854_ (
);

FILL FILL_1__8434_ (
);

FILL FILL_1__8014_ (
);

NOR2X1 _7084_ (
    .A(_668_),
    .B(_667_),
    .Y(_669_)
);

FILL FILL_3__9301_ (
);

FILL FILL_2__6777_ (
);

NAND3X1 _11082_ (
    .A(_4270_),
    .B(_4273_),
    .C(_4189_),
    .Y(_4280_)
);

FILL FILL_3__12971_ (
);

FILL FILL_1__9639_ (
);

FILL FILL_1__9219_ (
);

FILL FILL_3__12551_ (
);

FILL FILL_3__12131_ (
);

FILL FILL_2__11964_ (
);

FILL FILL_2__11544_ (
);

FILL FILL_2__11124_ (
);

NAND2X1 _8289_ (
    .A(_1725_),
    .B(_1727_),
    .Y(_1729_)
);

FILL FILL_1__10957_ (
);

FILL FILL_1__10537_ (
);

FILL FILL_1__10117_ (
);

FILL FILL_0__7964_ (
);

FILL FILL_0__7544_ (
);

AND2X2 _9650_ (
    .A(_2999_),
    .B(_2996_),
    .Y(_3003_)
);

FILL FILL_0__7124_ (
);

AOI21X1 _9230_ (
    .A(_2577_),
    .B(_2576_),
    .C(_2527_),
    .Y(_2590_)
);

OAI21X1 _12287_ (
    .A(_5376_),
    .B(_5383_),
    .C(_5382_),
    .Y(_5399_)
);

FILL FILL_2__8923_ (
);

FILL FILL_2__8503_ (
);

FILL FILL_2__12749_ (
);

FILL FILL_2__12329_ (
);

FILL FILL_1__6920_ (
);

FILL FILL_1__6500_ (
);

FILL FILL_0__8749_ (
);

FILL FILL_0__8329_ (
);

FILL FILL_3__6426_ (
);

FILL FILL_1__9392_ (
);

FILL FILL_2__9708_ (
);

FILL FILL_1__10290_ (
);

FILL FILL_1__7705_ (
);

NAND2X1 _6775_ (
    .A(_372_),
    .B(_367_),
    .Y(_373_)
);

FILL FILL_2__12082_ (
);

FILL FILL_1__11495_ (
);

FILL FILL_1__11075_ (
);

FILL FILL_0__10488_ (
);

NOR2X1 _10773_ (
    .A(_4755_),
    .B(_4763_),
    .Y(_4765_)
);

NAND3X1 _10353_ (
    .A(_3570_),
    .B(_3625_),
    .C(_3629_),
    .Y(_3630_)
);

FILL FILL_0__10068_ (
);

FILL FILL_2__10815_ (
);

FILL FILL_2__9461_ (
);

FILL FILL_2__9041_ (
);

FILL FILL_2__13287_ (
);

FILL FILL_0__6815_ (
);

INVX1 _8921_ (
    .A(\u_fir_pe2.rYin [13]),
    .Y(_2345_)
);

AOI21X1 _8501_ (
    .A(_1938_),
    .B(_1937_),
    .C(_1936_),
    .Y(_1939_)
);

FILL FILL_0__9287_ (
);

NAND3X1 _11978_ (
    .A(_5093_),
    .B(_5095_),
    .C(_5094_),
    .Y(_5096_)
);

OR2X2 _11558_ (
    .A(_4734_),
    .B(_4740_),
    .Y(_4742_)
);

NAND3X1 _11138_ (
    .A(_4334_),
    .B(_4335_),
    .C(_4333_),
    .Y(_4336_)
);

FILL FILL_1__13221_ (
);

FILL FILL_0__12634_ (
);

FILL FILL_0__12214_ (
);

OAI21X1 _9706_ (
    .A(_3042_),
    .B(_3038_),
    .C(_3051_),
    .Y(_3052_)
);

FILL FILL_1__8663_ (
);

FILL FILL_1__8243_ (
);

FILL FILL_3__9950_ (
);

FILL FILL_3__9530_ (
);

FILL FILL_2__6586_ (
);

FILL FILL_1__9448_ (
);

FILL FILL_1__9028_ (
);

FILL FILL_3__12360_ (
);

FILL FILL_2__11773_ (
);

FILL FILL_2__11353_ (
);

DFFPOSX1 _8098_ (
    .D(\X[1] [6]),
    .CLK(clk_bF$buf15),
    .Q(\X[2] [6])
);

FILL FILL_1__10766_ (
);

FILL FILL_1__10346_ (
);

FILL FILL_0__7773_ (
);

FILL FILL_0__7353_ (
);

NAND3X1 _12096_ (
    .A(_5208_),
    .B(_5212_),
    .C(_5167_),
    .Y(_5213_)
);

FILL FILL_2__8732_ (
);

FILL FILL_2__8312_ (
);

FILL FILL_0__10700_ (
);

FILL FILL_3__13145_ (
);

FILL FILL_2__12978_ (
);

FILL FILL_2__12558_ (
);

FILL FILL_2__12138_ (
);

FILL FILL_0__13172_ (
);

FILL FILL_0__8558_ (
);

FILL FILL_3__6655_ (
);

FILL FILL_0__8138_ (
);

INVX1 _10829_ (
    .A(_4017_),
    .Y(_4031_)
);

NAND2X1 _10409_ (
    .A(_3681_),
    .B(_3649_),
    .Y(_3685_)
);

FILL FILL_1__12912_ (
);

FILL FILL_2__9937_ (
);

FILL FILL_0__11905_ (
);

FILL FILL_2__9517_ (
);

FILL FILL_1__7934_ (
);

FILL FILL_1__7514_ (
);

AND2X2 _6584_ (
    .A(_134_),
    .B(_135_),
    .Y(_184_)
);

FILL FILL_3__8801_ (
);

FILL FILL253650x108150 (
);

FILL FILL_0__10297_ (
);

INVX1 _10582_ (
    .A(_3838_),
    .Y(_3848_)
);

NAND3X1 _10162_ (
    .A(_3434_),
    .B(_3437_),
    .C(_3435_),
    .Y(_3441_)
);

FILL FILL_1__8719_ (
);

FILL FILL_3__11211_ (
);

FILL FILL_2__9690_ (
);

FILL FILL_2__10624_ (
);

FILL FILL_2__9270_ (
);

FILL FILL_2__10204_ (
);

NAND2X1 _7789_ (
    .A(_1174_),
    .B(_1247_),
    .Y(_1305_)
);

NAND2X1 _7369_ (
    .A(vdd),
    .B(\X[1] [3]),
    .Y(_890_)
);

FILL FILL_2__13096_ (
);

FILL FILL_0__6624_ (
);

OR2X2 _8730_ (
    .A(_2163_),
    .B(_2159_),
    .Y(_2164_)
);

NAND2X1 _8310_ (
    .A(gnd),
    .B(\X[2]_5_bF$buf3 ),
    .Y(_1750_)
);

FILL FILL_1__12089_ (
);

FILL FILL_0__9096_ (
);

NAND3X1 _11787_ (
    .A(_4902_),
    .B(_4907_),
    .C(_4849_),
    .Y(_4908_)
);

NAND2X1 _11367_ (
    .A(_4557_),
    .B(_4560_),
    .Y(_4561_)
);

FILL FILL_1__13030_ (
);

FILL FILL_2__11829_ (
);

FILL FILL_0__12863_ (
);

FILL FILL_2__11409_ (
);

FILL FILL_0__12443_ (
);

FILL FILL_0__12023_ (
);

FILL FILL254250x201750 (
);

FILL FILL_0__7829_ (
);

INVX1 _9935_ (
    .A(_3216_),
    .Y(_3217_)
);

FILL FILL_0__7409_ (
);

OAI21X1 _9515_ (
    .A(_2465_),
    .B(_2710_),
    .C(_2864_),
    .Y(_2871_)
);

FILL FILL_1__8892_ (
);

FILL FILL_1__8472_ (
);

FILL FILL_1__8052_ (
);

FILL FILL_3__8398_ (
);

FILL FILL_0__13228_ (
);

FILL FILL_2__6395_ (
);

FILL FILL_1__9677_ (
);

FILL FILL_1__9257_ (
);

FILL FILL_2__11582_ (
);

FILL FILL_2__11162_ (
);

FILL FILL_1__10995_ (
);

FILL FILL_1__10575_ (
);

FILL FILL_1__10155_ (
);

FILL FILL_0__7582_ (
);

FILL FILL_0__7162_ (
);

FILL FILL_2__8541_ (
);

FILL FILL_2__12787_ (
);

FILL FILL_2__12367_ (
);

FILL FILL_0__8787_ (
);

FILL FILL_3__6884_ (
);

FILL FILL_0__8367_ (
);

NOR2X1 _10638_ (
    .A(_3901_),
    .B(_3900_),
    .Y(_3902_)
);

NOR2X1 _10218_ (
    .A(_3494_),
    .B(_3495_),
    .Y(_3496_)
);

FILL FILL_1__12721_ (
);

FILL FILL_1__12301_ (
);

FILL FILL_2__9746_ (
);

FILL FILL_2__9326_ (
);

FILL FILL_0__11714_ (
);

FILL FILL_1__7743_ (
);

FILL FILL_1__7323_ (
);

FILL FILL_3__7669_ (
);

NAND2X1 _6393_ (
    .A(_720_),
    .B(_784_),
    .Y(_785_)
);

FILL FILL_0__12919_ (
);

FILL FILL_3__10499_ (
);

NAND2X1 _10391_ (
    .A(_3665_),
    .B(_3666_),
    .Y(_3667_)
);

FILL FILL_1__8948_ (
);

FILL FILL_3__11860_ (
);

FILL FILL_1__8528_ (
);

FILL FILL_3__11440_ (
);

FILL FILL_3__11020_ (
);

FILL FILL_2__10853_ (
);

FILL FILL_2__10433_ (
);

FILL FILL_2__10013_ (
);

INVX1 _7598_ (
    .A(gnd),
    .Y(_1116_)
);

NOR2X1 _7178_ (
    .A(_759_),
    .B(_761_),
    .Y(_762_)
);

FILL FILL_0__6853_ (
);

FILL FILL_0__6433_ (
);

DFFPOSX1 _11596_ (
    .D(_4775_[12]),
    .CLK(clk_bF$buf35),
    .Q(\Y[6] [12])
);

NAND2X1 _11176_ (
    .A(gnd),
    .B(_4372_),
    .Y(_4373_)
);

FILL FILL_2__7812_ (
);

FILL FILL_3__12645_ (
);

FILL FILL_3__12225_ (
);

FILL FILL_0__12672_ (
);

FILL FILL_2__11218_ (
);

FILL FILL_0__12252_ (
);

FILL FILL_0__7638_ (
);

NAND2X1 _9744_ (
    .A(_3066_),
    .B(_3078_),
    .Y(_3087_)
);

AOI21X1 _9324_ (
    .A(_2678_),
    .B(_2677_),
    .C(_2579_),
    .Y(_2683_)
);

FILL FILL_1__8281_ (
);

FILL FILL_0__13037_ (
);

NOR2X1 _13322_ (
    .A(_6345_),
    .B(_6344_),
    .Y(_6369_[14])
);

FILL FILL_1__9486_ (
);

FILL FILL_1__9066_ (
);

FILL FILL_2__11391_ (
);

FILL FILL_1__10384_ (
);

FILL FILL_0__7391_ (
);

FILL FILL_2__8770_ (
);

FILL FILL_2__8350_ (
);

FILL FILL_3__13183_ (
);

INVX1 _6869_ (
    .A(_464_),
    .Y(_465_)
);

NAND3X1 _6449_ (
    .A(_40_),
    .B(_44_),
    .C(_46_),
    .Y(_51_)
);

FILL FILL_2__12596_ (
);

FILL FILL_2__12176_ (
);

OAI21X1 _7810_ (
    .A(_1270_),
    .B(_1323_),
    .C(_1324_),
    .Y(_1325_)
);

FILL FILL_1__11169_ (
);

FILL FILL_0__8596_ (
);

FILL FILL_0__8176_ (
);

NAND2X1 _10867_ (
    .A(vdd),
    .B(\X[5] [2]),
    .Y(_4068_)
);

INVX1 _10447_ (
    .A(_3719_),
    .Y(_3722_)
);

NAND3X1 _10027_ (
    .A(_3304_),
    .B(_3307_),
    .C(_3256_),
    .Y(_3308_)
);

FILL FILL_1__12950_ (
);

FILL FILL_1__12530_ (
);

FILL FILL_1__12110_ (
);

FILL FILL_2__10909_ (
);

FILL FILL_2__9975_ (
);

FILL FILL_2__9555_ (
);

FILL FILL_0__11943_ (
);

FILL FILL_2__9135_ (
);

FILL FILL_0__11523_ (
);

FILL FILL_0__11103_ (
);

FILL FILL_0__6909_ (
);

FILL FILL_1__7972_ (
);

FILL FILL_1__7552_ (
);

FILL FILL_1__7132_ (
);

FILL FILL_3__7898_ (
);

FILL FILL_1__13315_ (
);

FILL FILL_0__12728_ (
);

FILL FILL_0__12308_ (
);

FILL FILL_1__8757_ (
);

FILL FILL_1__8337_ (
);

FILL FILL_2__10662_ (
);

FILL FILL_2__10242_ (
);

FILL FILL_3__9624_ (
);

FILL FILL_3__9204_ (
);

FILL FILL_0__6662_ (
);

FILL FILL_2__7621_ (
);

FILL FILL_3__12454_ (
);

FILL FILL_2__11867_ (
);

FILL FILL_2__11447_ (
);

FILL FILL_2__11027_ (
);

FILL FILL_0__12061_ (
);

FILL FILL_0__7867_ (
);

NAND2X1 _9973_ (
    .A(_3254_),
    .B(_3248_),
    .Y(_3983_[4])
);

FILL FILL_0__7447_ (
);

NOR3X1 _9553_ (
    .A(_2696_),
    .B(_2864_),
    .C(_2807_),
    .Y(_2908_)
);

FILL FILL_0__7027_ (
);

OAI21X1 _9133_ (
    .A(_2489_),
    .B(_2490_),
    .C(_2475_),
    .Y(_2494_)
);

FILL FILL_1__11801_ (
);

FILL FILL_2__8826_ (
);

FILL FILL_2__8406_ (
);

FILL FILL_3__13239_ (
);

FILL FILL_0__13266_ (
);

AOI21X1 _13131_ (
    .A(_6136_),
    .B(_6138_),
    .C(_6164_),
    .Y(_6165_)
);

FILL FILL_1__6823_ (
);

FILL FILL_1__6403_ (
);

FILL FILL_3__6749_ (
);

FILL FILL_1__9295_ (
);

FILL FILL_2_CLKBUF1_insert60 (
);

FILL FILL_2_CLKBUF1_insert61 (
);

FILL FILL_2_CLKBUF1_insert62 (
);

FILL FILL_2_CLKBUF1_insert63 (
);

FILL FILL_2_CLKBUF1_insert64 (
);

FILL FILL_2_CLKBUF1_insert65 (
);

FILL FILL_2_CLKBUF1_insert66 (
);

FILL FILL_2_CLKBUF1_insert67 (
);

FILL FILL_2_CLKBUF1_insert68 (
);

FILL FILL_2_CLKBUF1_insert69 (
);

FILL FILL_1__10193_ (
);

FILL FILL_3__10940_ (
);

FILL FILL_1__7608_ (
);

FILL FILL_3__10100_ (
);

NAND3X1 _6678_ (
    .A(_271_),
    .B(_270_),
    .C(_272_),
    .Y(_277_)
);

FILL FILL_1__11398_ (
);

INVX1 _10676_ (
    .A(\u_fir_pe4.mul [13]),
    .Y(_3940_)
);

OAI21X1 _10256_ (
    .A(_3529_),
    .B(_3533_),
    .C(_3505_),
    .Y(_3534_)
);

FILL FILL_3__11725_ (
);

FILL FILL_2__9784_ (
);

FILL FILL_2__9364_ (
);

FILL FILL_0__11752_ (
);

FILL FILL_0__11332_ (
);

FILL FILL_0__6718_ (
);

INVX1 _8824_ (
    .A(\u_fir_pe2.mul [4]),
    .Y(_2250_)
);

INVX1 _8404_ (
    .A(_1842_),
    .Y(_1843_)
);

FILL FILL_1__7781_ (
);

FILL FILL_1__7361_ (
);

FILL FILL_3__7287_ (
);

FILL FILL_1__13124_ (
);

FILL FILL_0__12957_ (
);

NAND3X1 _12822_ (
    .A(_5788_),
    .B(_5856_),
    .C(_5857_),
    .Y(_5861_)
);

FILL FILL_0__12537_ (
);

FILL FILL_0__12117_ (
);

INVX1 _12402_ (
    .A(\u_fir_pe6.rYin [10]),
    .Y(_5506_)
);

NAND3X1 _9609_ (
    .A(_2955_),
    .B(_2962_),
    .C(_2961_),
    .Y(_2963_)
);

FILL FILL_1__8566_ (
);

FILL FILL_1__8146_ (
);

FILL FILL_2__10891_ (
);

FILL FILL_2__10471_ (
);

FILL FILL_2__10051_ (
);

FILL FILL_3__9013_ (
);

FILL FILL_0__6891_ (
);

FILL FILL_0__6471_ (
);

FILL FILL_2__6489_ (
);

FILL FILL_2__7850_ (
);

FILL FILL_3__12683_ (
);

FILL FILL_2__7430_ (
);

FILL FILL_2__7010_ (
);

FILL FILL_2__11676_ (
);

FILL FILL_2__11256_ (
);

FILL FILL_0__12290_ (
);

FILL FILL_1__10669_ (
);

FILL FILL_1__10249_ (
);

FILL FILL_0__7676_ (
);

NOR2X1 _9782_ (
    .A(_3125_),
    .B(_3124_),
    .Y(_3126_)
);

FILL FILL_0__7256_ (
);

AOI21X1 _9362_ (
    .A(_2719_),
    .B(_2717_),
    .C(_2715_),
    .Y(_2720_)
);

FILL FILL_2__8635_ (
);

FILL FILL_2__8215_ (
);

FILL FILL_0__10603_ (
);

DFFPOSX1 _13360_ (
    .D(\X[6] [6]),
    .CLK(clk_bF$buf37),
    .Q(\X[7] [6])
);

FILL FILL_0__13075_ (
);

FILL FILL_1__6632_ (
);

FILL FILL_2__13402_ (
);

FILL FILL_3__6978_ (
);

FILL FILL_1__12815_ (
);

FILL FILL_0__9822_ (
);

FILL FILL_0__9402_ (
);

FILL FILL_0__11808_ (
);

FILL FILL_1__7837_ (
);

FILL FILL_1__7417_ (
);

NAND2X1 _6487_ (
    .A(_36_),
    .B(_87_),
    .Y(_88_)
);

NAND2X1 _10485_ (
    .A(_3753_),
    .B(_3757_),
    .Y(_3759_)
);

INVX1 _10065_ (
    .A(_3344_),
    .Y(_3345_)
);

FILL FILL_3__11954_ (
);

FILL FILL_2__6701_ (
);

FILL FILL_3__11534_ (
);

FILL FILL_3__11114_ (
);

FILL FILL_2__10947_ (
);

FILL FILL_2__9593_ (
);

FILL FILL_0__11981_ (
);

FILL FILL_2__10527_ (
);

FILL FILL_2__9173_ (
);

FILL FILL_0__11561_ (
);

FILL FILL_2__10107_ (
);

FILL FILL_0__11141_ (
);

FILL FILL_3__9909_ (
);

FILL FILL_0__6947_ (
);

FILL FILL_0__6527_ (
);

AND2X2 _8633_ (
    .A(_2067_),
    .B(_2010_),
    .Y(_2069_)
);

NAND3X1 _8213_ (
    .A(_1622_),
    .B(_1639_),
    .C(_1642_),
    .Y(_1655_)
);

FILL FILL_1__7590_ (
);

FILL FILL_1__7170_ (
);

FILL FILL_3__7096_ (
);

FILL FILL_2__7906_ (
);

FILL FILL_3__12739_ (
);

FILL FILL_3__12319_ (
);

FILL FILL_0__12766_ (
);

NAND2X1 _12631_ (
    .A(vdd),
    .B(\X[6] [3]),
    .Y(_5672_)
);

FILL FILL_0__12346_ (
);

NAND2X1 _12211_ (
    .A(_5322_),
    .B(_5298_),
    .Y(_5326_)
);

DFFPOSX1 _9838_ (
    .D(_3181_[8]),
    .CLK(clk_bF$buf0),
    .Q(\Y[4] [8])
);

AOI21X1 _9418_ (
    .A(_2740_),
    .B(_2741_),
    .C(_2708_),
    .Y(_2775_)
);

FILL FILL_1__8795_ (
);

FILL FILL_1__8375_ (
);

FILL FILL_2__10280_ (
);

FILL FILL_3__9242_ (
);

BUFX2 _13416_ (
    .A(_6377_[8]),
    .Y(Yout[8])
);

FILL FILL_3__12072_ (
);

FILL FILL_2__11485_ (
);

FILL FILL_2__11065_ (
);

FILL FILL_1__10898_ (
);

FILL FILL_1__10478_ (
);

FILL FILL_1__10058_ (
);

FILL FILL_0__7485_ (
);

OAI21X1 _9591_ (
    .A(_2895_),
    .B(_2898_),
    .C(_2943_),
    .Y(_2946_)
);

FILL FILL_0__7065_ (
);

INVX1 _9171_ (
    .A(_2530_),
    .Y(_2531_)
);

FILL FILL_3__10805_ (
);

FILL FILL_2__8864_ (
);

FILL FILL_2__8444_ (
);

FILL FILL_0__10832_ (
);

FILL FILL_0__10412_ (
);

FILL FILL_2__8024_ (
);

OR2X2 _7904_ (
    .A(_1414_),
    .B(_1415_),
    .Y(_1416_)
);

FILL FILL_1__6861_ (
);

FILL FILL_1__6441_ (
);

FILL FILL_2__13211_ (
);

FILL FILL_1__12624_ (
);

FILL FILL_1__12204_ (
);

FILL FILL_2__9649_ (
);

FILL FILL_0__9631_ (
);

FILL FILL_0__9211_ (
);

FILL FILL_2__9229_ (
);

OAI21X1 _11902_ (
    .A(_4938_),
    .B(_4942_),
    .C(_4941_),
    .Y(_5021_)
);

FILL FILL_1__7646_ (
);

FILL FILL_1__13409_ (
);

FILL FILL_3__8513_ (
);

OAI21X1 _10294_ (
    .A(_3492_),
    .B(_3496_),
    .C(_3501_),
    .Y(_3571_)
);

FILL FILL_2__6930_ (
);

FILL FILL_2__6510_ (
);

FILL FILL_0__11790_ (
);

FILL FILL_2__10336_ (
);

FILL FILL_0__11370_ (
);

FILL FILL_3__9718_ (
);

FILL FILL_0__6756_ (
);

INVX1 _8862_ (
    .A(\u_fir_pe2.mul [8]),
    .Y(_2285_)
);

NAND3X1 _8442_ (
    .A(_1729_),
    .B(_1868_),
    .C(_1873_),
    .Y(_1881_)
);

NAND2X1 _8022_ (
    .A(_1525_),
    .B(_1520_),
    .Y(_1526_)
);

OAI21X1 _11499_ (
    .A(_4666_),
    .B(_4667_),
    .C(_4681_),
    .Y(_4682_)
);

INVX1 _11079_ (
    .A(_4273_),
    .Y(_4278_)
);

FILL FILL_3__12968_ (
);

FILL FILL_2__7715_ (
);

FILL FILL_1__13162_ (
);

FILL FILL_0__12995_ (
);

INVX1 _12860_ (
    .A(gnd),
    .Y(_5898_)
);

FILL FILL_0__12575_ (
);

FILL FILL_0__12155_ (
);

NOR2X1 _12440_ (
    .A(_5541_),
    .B(_5543_),
    .Y(_5544_)
);

AOI21X1 _12020_ (
    .A(_5137_),
    .B(_5136_),
    .C(_5135_),
    .Y(_5138_)
);

FILL FILL_2__12902_ (
);

NAND2X1 _9647_ (
    .A(_2996_),
    .B(_2999_),
    .Y(_3000_)
);

NAND3X1 _9227_ (
    .A(_2581_),
    .B(_2582_),
    .C(_2583_),
    .Y(_2587_)
);

FILL FILL_1__8184_ (
);

FILL FILL254550x79350 (
);

FILL FILL_0__8902_ (
);

FILL FILL_3__9891_ (
);

FILL FILL_3__9471_ (
);

OR2X2 _13225_ (
    .A(_6243_),
    .B(_6248_),
    .Y(_6250_)
);

FILL FILL_1__6917_ (
);

FILL FILL_1__9389_ (
);

FILL FILL_2__11294_ (
);

FILL FILL_1__10287_ (
);

FILL FILL_0__7294_ (
);

FILL FILL_2__8673_ (
);

FILL FILL_2__8253_ (
);

FILL FILL_0__10641_ (
);

FILL FILL_3__13086_ (
);

FILL FILL_0__10221_ (
);

FILL FILL_2__12079_ (
);

AOI21X1 _7713_ (
    .A(_1150_),
    .B(_1152_),
    .C(_1229_),
    .Y(_1230_)
);

FILL FILL_1__6670_ (
);

FILL FILL_2__13020_ (
);

FILL FILL_0__8499_ (
);

FILL FILL_3__6596_ (
);

FILL FILL_3__11819_ (
);

FILL FILL_1__12853_ (
);

FILL FILL_1__12433_ (
);

FILL FILL_1__12013_ (
);

FILL FILL_2__9458_ (
);

FILL FILL_0__9440_ (
);

FILL FILL_0__11846_ (
);

FILL FILL_2__9038_ (
);

FILL FILL_0__9020_ (
);

NAND3X1 _11711_ (
    .A(_4822_),
    .B(_4826_),
    .C(_4828_),
    .Y(_4833_)
);

FILL FILL_0__11426_ (
);

FILL FILL_0__11006_ (
);

OR2X2 _8918_ (
    .A(_2335_),
    .B(_2340_),
    .Y(_2342_)
);

FILL FILL_1__7875_ (
);

FILL FILL_1__7455_ (
);

FILL FILL_1__7035_ (
);

FILL FILL_1__13218_ (
);

FILL FILL_3__8742_ (
);

OAI21X1 _12916_ (
    .A(_5781_),
    .B(_5871_),
    .C(_5867_),
    .Y(_5954_)
);

FILL FILL_3__11152_ (
);

FILL FILL_2__10985_ (
);

FILL FILL_2__10565_ (
);

FILL FILL_2__10145_ (
);

FILL FILL_1__9601_ (
);

FILL FILL_0__6985_ (
);

FILL FILL_0__6565_ (
);

NAND2X1 _8671_ (
    .A(_2099_),
    .B(_2103_),
    .Y(_2106_)
);

AOI21X1 _8251_ (
    .A(_1686_),
    .B(_1688_),
    .C(_1679_),
    .Y(_1692_)
);

FILL FILL_2__7944_ (
);

FILL FILL_3__12777_ (
);

FILL FILL_2__7524_ (
);

FILL FILL_2__7104_ (
);

FILL FILL_0__12384_ (
);

FILL FILL_2__12711_ (
);

DFFPOSX1 _9876_ (
    .D(_3187_[6]),
    .CLK(clk_bF$buf14),
    .Q(\u_fir_pe3.mul [6])
);

NAND3X1 _9456_ (
    .A(_2810_),
    .B(_2811_),
    .C(_2812_),
    .Y(_2813_)
);

OAI21X1 _9036_ (
    .A(_2395_),
    .B(_2398_),
    .C(_2391_),
    .Y(_2399_)
);

FILL FILL_1__11704_ (
);

FILL FILL_2__8729_ (
);

FILL FILL_0__8711_ (
);

FILL FILL_2__8309_ (
);

FILL FILL_0__13169_ (
);

NAND3X1 _13034_ (
    .A(_6067_),
    .B(_6069_),
    .C(_6068_),
    .Y(_6070_)
);

FILL FILL_1__6726_ (
);

FILL FILL_1__9198_ (
);

FILL FILL_1__12909_ (
);

FILL FILL_0__9916_ (
);

FILL FILL_1__10096_ (
);

FILL FILL_3__10423_ (
);

FILL FILL_2__8482_ (
);

FILL FILL_0__10870_ (
);

FILL FILL_0__10450_ (
);

FILL FILL_2__8062_ (
);

FILL FILL_0__10030_ (
);

NOR2X1 _7942_ (
    .A(_1448_),
    .B(_1447_),
    .Y(_1449_)
);

OAI21X1 _7522_ (
    .A(_886_),
    .B(_871_),
    .C(_955_),
    .Y(_1041_)
);

OAI21X1 _7102_ (
    .A(_683_),
    .B(_684_),
    .C(_680_),
    .Y(_685_)
);

INVX1 _10999_ (
    .A(_4197_),
    .Y(_4198_)
);

NOR2X1 _10579_ (
    .A(_3843_),
    .B(_3844_),
    .Y(_3845_)
);

AOI21X1 _10159_ (
    .A(_3435_),
    .B(_3437_),
    .C(_3434_),
    .Y(_3438_)
);

FILL FILL_1__12662_ (
);

FILL FILL_3__11208_ (
);

FILL FILL_1__12242_ (
);

FILL FILL_2__9687_ (
);

NAND3X1 _11940_ (
    .A(_5053_),
    .B(_5052_),
    .C(_5054_),
    .Y(_5059_)
);

FILL FILL_2__9267_ (
);

FILL FILL_0__11655_ (
);

NOR2X1 _11520_ (
    .A(_4700_),
    .B(_4694_),
    .Y(_4703_)
);

FILL FILL_0__11235_ (
);

NAND2X1 _11100_ (
    .A(_4291_),
    .B(_4292_),
    .Y(_4298_)
);

NOR2X1 _8727_ (
    .A(_1738_),
    .B(_1899_),
    .Y(_2161_)
);

NAND2X1 _8307_ (
    .A(vdd),
    .B(\X[2] [3]),
    .Y(_1747_)
);

FILL FILL_1__7684_ (
);

FILL FILL_1__7264_ (
);

FILL FILL_1__13027_ (
);

NAND3X1 _12725_ (
    .A(_5751_),
    .B(_5755_),
    .C(_5758_),
    .Y(_5765_)
);

INVX1 _12305_ (
    .A(\u_fir_pe6.rYin [1]),
    .Y(_5414_)
);

FILL FILL_1__8889_ (
);

FILL FILL_1__8469_ (
);

FILL FILL_1__8049_ (
);

FILL FILL_3__11381_ (
);

FILL FILL_2__10794_ (
);

FILL FILL_2__10374_ (
);

FILL FILL_1__9410_ (
);

FILL FILL_3__9336_ (
);

FILL FILL_0__6794_ (
);

NAND2X1 _8480_ (
    .A(gnd),
    .B(\X[2] [7]),
    .Y(_1918_)
);

NOR2X1 _8060_ (
    .A(_1563_),
    .B(_1562_),
    .Y(_1587_[14])
);

FILL FILL_2__7753_ (
);

FILL FILL_3__12586_ (
);

FILL FILL_2__7333_ (
);

FILL FILL_3__12166_ (
);

FILL FILL_2__11999_ (
);

FILL FILL_2__11579_ (
);

FILL FILL_2__11159_ (
);

FILL FILL_0__12193_ (
);

FILL FILL_2__12940_ (
);

FILL FILL_2__12520_ (
);

FILL FILL_0__7999_ (
);

FILL FILL_2__12100_ (
);

FILL FILL_0__7579_ (
);

NOR2X1 _9685_ (
    .A(\u_fir_pe3.rYin [2]),
    .B(\u_fir_pe3.mul [2]),
    .Y(_3033_)
);

FILL FILL_0__7159_ (
);

INVX1 _9265_ (
    .A(gnd),
    .Y(_2624_)
);

FILL FILL_1__11933_ (
);

FILL FILL_1__11513_ (
);

FILL FILL_0__8940_ (
);

FILL FILL_2__8538_ (
);

FILL FILL_0__8520_ (
);

FILL FILL_0__10926_ (
);

FILL FILL_0__10506_ (
);

FILL FILL_0__13398_ (
);

NAND2X1 _13263_ (
    .A(_6283_),
    .B(_6286_),
    .Y(_6369_[8])
);

FILL FILL_1__6955_ (
);

FILL FILL_1__6535_ (
);

FILL FILL_2__13305_ (
);

FILL FILL_1__12718_ (
);

FILL FILL_0__9725_ (
);

FILL FILL_3__7822_ (
);

FILL FILL_0__9305_ (
);

FILL FILL_3__10652_ (
);

FILL FILL_2__8291_ (
);

FILL FILL_3__8607_ (
);

AND2X2 _7751_ (
    .A(_1263_),
    .B(_1266_),
    .Y(_1267_)
);

NAND2X1 _7331_ (
    .A(_846_),
    .B(_849_),
    .Y(_853_)
);

OAI22X1 _10388_ (
    .A(_3519_),
    .B(_3600_),
    .C(_3662_),
    .D(_3663_),
    .Y(_3664_)
);

FILL FILL_2__6604_ (
);

FILL FILL_1__12891_ (
);

FILL FILL_3__11437_ (
);

FILL FILL_1__12051_ (
);

FILL FILL_2__9496_ (
);

FILL FILL_0__11884_ (
);

FILL FILL_2__9076_ (
);

FILL FILL_0__11464_ (
);

FILL FILL_0__11044_ (
);

DFFPOSX1 _8956_ (
    .D(_2384_[3]),
    .CLK(clk_bF$buf47),
    .Q(\Y[3] [3])
);

INVX1 _8536_ (
    .A(_1966_),
    .Y(_1973_)
);

DFFPOSX1 _8116_ (
    .D(_1588_[0]),
    .CLK(clk_bF$buf13),
    .Q(\u_fir_pe1.mul [0])
);

FILL FILL_1__7493_ (
);

FILL FILL_1__7073_ (
);

FILL FILL_2__7809_ (
);

FILL FILL_1__13256_ (
);

FILL FILL_3__8780_ (
);

NAND2X1 _12954_ (
    .A(vdd),
    .B(\X[6] [7]),
    .Y(_5991_)
);

FILL FILL_0__12669_ (
);

FILL FILL_3__8360_ (
);

FILL FILL_0__12249_ (
);

NAND2X1 _12534_ (
    .A(gnd),
    .B(\X[6] [3]),
    .Y(_6366_)
);

OAI21X1 _12114_ (
    .A(_5229_),
    .B(_5230_),
    .C(_5226_),
    .Y(_5231_)
);

FILL FILL_1__8698_ (
);

FILL FILL_1__8278_ (
);

FILL FILL_2__10183_ (
);

FILL FILL_3__9985_ (
);

FILL FILL_3__9565_ (
);

FILL FILL_3__9145_ (
);

NOR2X1 _13319_ (
    .A(_6342_),
    .B(_6341_),
    .Y(_6343_)
);

FILL FILL_2__7982_ (
);

FILL FILL_2__7562_ (
);

FILL FILL_3__12395_ (
);

FILL FILL_2__7142_ (
);

FILL FILL_2__11388_ (
);

NAND3X1 _6602_ (
    .A(_195_),
    .B(_196_),
    .C(_201_),
    .Y(_202_)
);

FILL FILL_0__7388_ (
);

OAI21X1 _9494_ (
    .A(_2829_),
    .B(_2831_),
    .C(_2822_),
    .Y(_2850_)
);

NAND3X1 _9074_ (
    .A(_2423_),
    .B(_2435_),
    .C(_2431_),
    .Y(_2436_)
);

FILL FILL_1__11742_ (
);

FILL FILL_1__11322_ (
);

FILL FILL_2__8767_ (
);

FILL FILL_2__8347_ (
);

FILL FILL_0__10315_ (
);

NOR2X1 _10600_ (
    .A(\u_fir_pe4.rYin [6]),
    .B(\u_fir_pe4.mul [6]),
    .Y(_3864_)
);

OAI21X1 _13072_ (
    .A(_6052_),
    .B(_6105_),
    .C(_6106_),
    .Y(_6107_)
);

NAND2X1 _7807_ (
    .A(_1128_),
    .B(_1202_),
    .Y(_1322_)
);

FILL FILL_1__6764_ (
);

FILL FILL_2__13114_ (
);

FILL FILL_1__12947_ (
);

FILL FILL_1__12527_ (
);

FILL FILL_1__12107_ (
);

FILL FILL_0__9954_ (
);

FILL FILL_0__9534_ (
);

FILL FILL_0__9114_ (
);

NAND2X1 _11805_ (
    .A(_4923_),
    .B(_4924_),
    .Y(_4925_)
);

FILL FILL_1__7969_ (
);

FILL FILL_3__10881_ (
);

FILL FILL_1__7549_ (
);

FILL FILL_1__7129_ (
);

FILL FILL_3__10041_ (
);

FILL FILL_1__8910_ (
);

FILL FILL_3__8836_ (
);

INVX1 _7980_ (
    .A(_1477_),
    .Y(_1483_)
);

NAND3X1 _7560_ (
    .A(_1006_),
    .B(_1074_),
    .C(_1075_),
    .Y(_1079_)
);

INVX1 _7140_ (
    .A(\u_fir_pe0.rYin [10]),
    .Y(_724_)
);

NAND3X1 _10197_ (
    .A(_3376_),
    .B(_3474_),
    .C(_3475_),
    .Y(_3476_)
);

FILL FILL_2__6833_ (
);

FILL FILL_3__11666_ (
);

FILL FILL_2__6413_ (
);

FILL FILL_3__11246_ (
);

FILL FILL_1__12280_ (
);

FILL FILL_2__10659_ (
);

FILL FILL_0__11693_ (
);

FILL FILL_2__10239_ (
);

FILL FILL_0__11273_ (
);

FILL FILL_0__6659_ (
);

NAND2X1 _8765_ (
    .A(_2196_),
    .B(_2197_),
    .Y(_2198_)
);

NAND3X1 _8345_ (
    .A(_1778_),
    .B(_1771_),
    .C(_1776_),
    .Y(_1785_)
);

FILL FILL_0__7600_ (
);

FILL FILL_2__7618_ (
);

FILL FILL_1__13065_ (
);

FILL FILL_0__12898_ (
);

AOI21X1 _12763_ (
    .A(_5741_),
    .B(_5745_),
    .C(_5734_),
    .Y(_5802_)
);

FILL FILL_0__12058_ (
);

INVX1 _12343_ (
    .A(\u_fir_pe6.mul [5]),
    .Y(_5448_)
);

FILL FILL_2__12805_ (
);

FILL FILL_0__8805_ (
);

FILL FILL_3__6902_ (
);

FILL FILL_3__9794_ (
);

OR2X2 _13128_ (
    .A(_6160_),
    .B(_6158_),
    .Y(_6162_)
);

FILL FILL_2__7791_ (
);

FILL FILL_2__7371_ (
);

FILL FILL_2__11197_ (
);

AOI21X1 _6831_ (
    .A(_343_),
    .B(_349_),
    .C(_424_),
    .Y(_428_)
);

NAND3X1 _6411_ (
    .A(_788_),
    .B(_13_),
    .C(_9_),
    .Y(_14_)
);

FILL FILL_0__7197_ (
);

FILL FILL_1__11971_ (
);

FILL FILL_3__10517_ (
);

FILL FILL_1__11551_ (
);

FILL FILL_1__11131_ (
);

FILL FILL_2__8576_ (
);

FILL FILL_0__10964_ (
);

FILL FILL_2__8156_ (
);

FILL FILL_0__10544_ (
);

FILL FILL_0__10124_ (
);

FILL FILL254550x165750 (
);

AOI21X1 _7616_ (
    .A(_1043_),
    .B(_1046_),
    .C(_1052_),
    .Y(_1134_)
);

FILL FILL_1__6993_ (
);

FILL FILL_1__6573_ (
);

FILL FILL_1__12756_ (
);

FILL FILL_1__12336_ (
);

FILL FILL_0__9763_ (
);

FILL FILL_0__9343_ (
);

FILL FILL_0__11749_ (
);

FILL FILL_3__7440_ (
);

DFFPOSX1 _11614_ (
    .D(\Y[5] [6]),
    .CLK(clk_bF$buf57),
    .Q(\u_fir_pe5.rYin [6])
);

FILL FILL_0__11329_ (
);

FILL FILL_1__7778_ (
);

FILL FILL_3__10690_ (
);

FILL FILL_1__7358_ (
);

FILL FILL_3__10270_ (
);

NAND3X1 _12819_ (
    .A(_5856_),
    .B(_5857_),
    .C(_5855_),
    .Y(_5858_)
);

FILL FILL_3__8225_ (
);

FILL FILL_3__11895_ (
);

FILL FILL_2__6642_ (
);

FILL FILL_3__11475_ (
);

FILL FILL_3__11055_ (
);

FILL FILL_2__10888_ (
);

FILL FILL_2__10468_ (
);

FILL FILL_2__10048_ (
);

FILL FILL_0__11082_ (
);

FILL FILL_1__9924_ (
);

FILL FILL_1__9504_ (
);

FILL FILL_0__6888_ (
);

DFFPOSX1 _8994_ (
    .D(_2386_[1]),
    .CLK(clk_bF$buf53),
    .Q(\u_fir_pe2.mul [1])
);

FILL FILL_0__6468_ (
);

INVX1 _8574_ (
    .A(\X[2] [4]),
    .Y(_2011_)
);

OR2X2 _8154_ (
    .A(_2325_),
    .B(_1596_),
    .Y(_1597_)
);

FILL FILL_1__10822_ (
);

FILL FILL_1__10402_ (
);

FILL FILL_2__7847_ (
);

FILL FILL_2__7427_ (
);

FILL FILL_2__7007_ (
);

FILL FILL_1__13294_ (
);

AND2X2 _12992_ (
    .A(_6028_),
    .B(_6021_),
    .Y(_6029_)
);

FILL FILL_0__12287_ (
);

AND2X2 _12572_ (
    .A(vdd),
    .B(\X[6] [1]),
    .Y(_5614_)
);

NAND3X1 _12152_ (
    .A(_5189_),
    .B(_5267_),
    .C(_5197_),
    .Y(_5268_)
);

FILL FILL_2__12614_ (
);

OAI21X1 _9779_ (
    .A(_3115_),
    .B(_3116_),
    .C(_3120_),
    .Y(_3123_)
);

NAND3X1 _9359_ (
    .A(gnd),
    .B(\X[3] [6]),
    .C(_2716_),
    .Y(_2717_)
);

FILL FILL_0__8614_ (
);

FILL FILL_3__6711_ (
);

FILL FILL_3__9183_ (
);

DFFPOSX1 _13357_ (
    .D(\X[6] [3]),
    .CLK(clk_bF$buf49),
    .Q(\X[7] [3])
);

FILL FILL_1__6629_ (
);

FILL FILL_2__7180_ (
);

FILL FILL_0__9819_ (
);

FILL FILL_3__7916_ (
);

OAI21X1 _6640_ (
    .A(_156_),
    .B(_160_),
    .C(_159_),
    .Y(_239_)
);

FILL FILL_1__11780_ (
);

FILL FILL_1__11360_ (
);

FILL FILL_2__8385_ (
);

FILL FILL_0__10773_ (
);

FILL FILL_0__10353_ (
);

OAI21X1 _7845_ (
    .A(_1327_),
    .B(_1321_),
    .C(_1331_),
    .Y(_1359_)
);

NAND3X1 _7425_ (
    .A(gnd),
    .B(\X[1] [6]),
    .C(_942_),
    .Y(_945_)
);

NAND2X1 _7005_ (
    .A(_597_),
    .B(_596_),
    .Y(_598_)
);

FILL FILL_1__6382_ (
);

FILL FILL_2__13152_ (
);

FILL FILL_1__12985_ (
);

FILL FILL_1__12565_ (
);

FILL FILL_1__12145_ (
);

FILL FILL_0__9992_ (
);

FILL FILL_0__11978_ (
);

FILL FILL_0__9572_ (
);

FILL FILL_0__9152_ (
);

AOI21X1 _11843_ (
    .A(_4953_),
    .B(_4949_),
    .C(_4934_),
    .Y(_4963_)
);

FILL FILL_0__11558_ (
);

OAI21X1 _11423_ (
    .A(_4601_),
    .B(_4600_),
    .C(_4612_),
    .Y(_4614_)
);

FILL FILL_0__11138_ (
);

NAND3X1 _11003_ (
    .A(_4128_),
    .B(_4197_),
    .C(_4132_),
    .Y(_4202_)
);

FILL FILL_1__7587_ (
);

FILL FILL_1__7167_ (
);

FILL FILL_3__8874_ (
);

FILL FILL_3__8454_ (
);

OAI21X1 _12628_ (
    .A(_5668_),
    .B(_5594_),
    .C(_5662_),
    .Y(_5669_)
);

FILL FILL_3__8034_ (
);

NAND2X1 _12208_ (
    .A(_5322_),
    .B(_5321_),
    .Y(_5323_)
);

FILL FILL_2__6871_ (
);

FILL FILL_2__6451_ (
);

FILL FILL_2__10697_ (
);

FILL FILL_2__10277_ (
);

FILL FILL_1__9733_ (
);

FILL FILL_1__9313_ (
);

FILL FILL_3__9659_ (
);

FILL FILL_3__9239_ (
);

FILL FILL_0__6697_ (
);

AND2X2 _8383_ (
    .A(vdd),
    .B(\X[2] [7]),
    .Y(_1822_)
);

FILL FILL253950x241350 (
);

FILL FILL_1__10631_ (
);

FILL FILL_1__10211_ (
);

FILL FILL_2__7656_ (
);

FILL FILL_0__12096_ (
);

NAND2X1 _12381_ (
    .A(_5481_),
    .B(_5484_),
    .Y(_5485_)
);

FILL FILL_3__13010_ (
);

FILL FILL_2__12843_ (
);

FILL FILL_2__12423_ (
);

FILL FILL_2__12003_ (
);

NAND2X1 _9588_ (
    .A(_2939_),
    .B(_2942_),
    .Y(_2943_)
);

AOI21X1 _9168_ (
    .A(_2482_),
    .B(_2486_),
    .C(_2475_),
    .Y(_2528_)
);

FILL FILL_1__11836_ (
);

FILL FILL_1__11416_ (
);

FILL FILL_0__8843_ (
);

FILL FILL_0__8423_ (
);

FILL FILL_0__10829_ (
);

FILL FILL_3__6520_ (
);

FILL FILL_0__10409_ (
);

FILL FILL_0__8003_ (
);

OR2X2 _13166_ (
    .A(_6196_),
    .B(_6197_),
    .Y(_6198_)
);

FILL FILL_2__9802_ (
);

FILL FILL_1__6858_ (
);

FILL FILL_1__6438_ (
);

FILL FILL_2__13208_ (
);

FILL FILL_0__9628_ (
);

FILL FILL_0__9208_ (
);

FILL FILL_3__7305_ (
);

FILL FILL_3__10975_ (
);

FILL FILL_3__10135_ (
);

FILL FILL_2__8194_ (
);

FILL FILL_0__10582_ (
);

FILL FILL_0__10162_ (
);

OAI21X1 _7654_ (
    .A(_999_),
    .B(_1089_),
    .C(_1085_),
    .Y(_1172_)
);

DFFPOSX1 _7234_ (
    .D(Yin[11]),
    .CLK(clk_bF$buf41),
    .Q(\u_fir_pe0.rYin [11])
);

FILL FILL_2__6927_ (
);

FILL FILL_2__6507_ (
);

FILL FILL_1__12794_ (
);

FILL FILL_1__12374_ (
);

FILL FILL_0__9381_ (
);

FILL FILL_2__9399_ (
);

FILL FILL_0__11787_ (
);

INVX1 _11652_ (
    .A(_5563_),
    .Y(_5564_)
);

FILL FILL_0__11367_ (
);

AOI21X1 _11232_ (
    .A(_4285_),
    .B(_4350_),
    .C(_4428_),
    .Y(_4429_)
);

NAND2X1 _8859_ (
    .A(_2281_),
    .B(_2280_),
    .Y(_2282_)
);

AOI21X1 _8439_ (
    .A(_1877_),
    .B(_1876_),
    .C(_1875_),
    .Y(_1878_)
);

NOR2X1 _8019_ (
    .A(_1521_),
    .B(_1522_),
    .Y(_1523_)
);

FILL FILL_1__7396_ (
);

NOR2X1 _9800_ (
    .A(_3142_),
    .B(_3143_),
    .Y(_3144_)
);

FILL FILL_1__13159_ (
);

FILL FILL_3__8683_ (
);

AOI21X1 _12857_ (
    .A(_5835_),
    .B(_5832_),
    .C(_5818_),
    .Y(_5895_)
);

OAI21X1 _12437_ (
    .A(_5533_),
    .B(_5534_),
    .C(_5538_),
    .Y(_5540_)
);

AND2X2 _12017_ (
    .A(_5096_),
    .B(_5092_),
    .Y(_5135_)
);

FILL FILL253950x90150 (
);

FILL FILL_2__6680_ (
);

FILL FILL_3__11093_ (
);

FILL FILL_2__10086_ (
);

FILL FILL_1__9962_ (
);

FILL FILL_1__9542_ (
);

FILL FILL_1__9122_ (
);

NAND3X1 _8192_ (
    .A(_1628_),
    .B(_1633_),
    .C(_1631_),
    .Y(_1634_)
);

FILL FILL_1__10860_ (
);

FILL FILL_1__10440_ (
);

FILL FILL_1__10020_ (
);

FILL FILL253950x57750 (
);

FILL FILL_2__7885_ (
);

FILL FILL_2__7465_ (
);

FILL FILL_2__7045_ (
);

NAND3X1 _12190_ (
    .A(_5302_),
    .B(_5303_),
    .C(_5304_),
    .Y(_5305_)
);

NOR2X1 _6925_ (
    .A(_417_),
    .B(_462_),
    .Y(_520_)
);

NAND3X1 _6505_ (
    .A(_101_),
    .B(_105_),
    .C(_69_),
    .Y(_106_)
);

FILL FILL_2__12652_ (
);

FILL FILL_2__12232_ (
);

NAND3X1 _9397_ (
    .A(_2694_),
    .B(_2751_),
    .C(_2752_),
    .Y(_2755_)
);

FILL FILL_1__11645_ (
);

FILL FILL_1__11225_ (
);

FILL FILL_0__8652_ (
);

FILL FILL_0__8232_ (
);

FILL FILL_0__10638_ (
);

OAI21X1 _10923_ (
    .A(_4087_),
    .B(_4122_),
    .C(_4081_),
    .Y(_4123_)
);

INVX1 _10503_ (
    .A(_3773_),
    .Y(_3777_)
);

FILL FILL_0__10218_ (
);

BUFX2 _13395_ (
    .A(_6376_[1]),
    .Y(Xout[1])
);

FILL FILL_2__9611_ (
);

FILL FILL_1__6667_ (
);

FILL FILL_2__13017_ (
);

FILL FILL_0__9437_ (
);

FILL FILL_3__7534_ (
);

FILL FILL_0__9017_ (
);

NAND2X1 _11708_ (
    .A(_4828_),
    .B(_4829_),
    .Y(_4830_)
);

FILL FILL_3__10364_ (
);

FILL FILL_0__10391_ (
);

FILL FILL_1__8813_ (
);

FILL FILL_3__8319_ (
);

NAND2X1 _7883_ (
    .A(_1395_),
    .B(_1369_),
    .Y(_1396_)
);

NAND3X1 _7463_ (
    .A(_969_),
    .B(_973_),
    .C(_976_),
    .Y(_983_)
);

INVX1 _7043_ (
    .A(\u_fir_pe0.rYin [1]),
    .Y(_632_)
);

FILL FILL_2__13190_ (
);

FILL FILL_3__11989_ (
);

FILL FILL_2__6736_ (
);

FILL FILL_3__11569_ (
);

FILL FILL_3__11149_ (
);

FILL FILL_1__12183_ (
);

FILL FILL_0__9190_ (
);

NAND3X1 _11881_ (
    .A(_4993_),
    .B(_4999_),
    .C(_4998_),
    .Y(_5000_)
);

NAND2X1 _11461_ (
    .A(_4644_),
    .B(_4646_),
    .Y(_4647_)
);

FILL FILL_0__11176_ (
);

NOR2X1 _11041_ (
    .A(_4226_),
    .B(_4239_),
    .Y(_4240_)
);

FILL FILL_2__11923_ (
);

FILL FILL_2__11503_ (
);

NOR2X1 _8668_ (
    .A(_2099_),
    .B(_2103_),
    .Y(_2104_)
);

NAND3X1 _8248_ (
    .A(_1679_),
    .B(_1686_),
    .C(_1688_),
    .Y(_1689_)
);

FILL FILL_1__10916_ (
);

FILL FILL_0__7923_ (
);

FILL FILL_0__7503_ (
);

FILL FILL_3__8492_ (
);

INVX1 _12666_ (
    .A(_5699_),
    .Y(_5707_)
);

NAND3X1 _12246_ (
    .A(_5344_),
    .B(_5354_),
    .C(_5357_),
    .Y(_5360_)
);

FILL FILL_2__12708_ (
);

FILL FILL_0__13322_ (
);

FILL FILL_0__8708_ (
);

FILL FILL_3__6805_ (
);

FILL FILL_1__9771_ (
);

FILL FILL_1__9351_ (
);

FILL FILL_3__9277_ (
);

FILL FILL_2__7694_ (
);

FILL FILL_2__7274_ (
);

NAND2X1 _6734_ (
    .A(_327_),
    .B(_331_),
    .Y(_332_)
);

FILL FILL_2__12881_ (
);

FILL FILL_2__12041_ (
);

FILL FILL_1__11874_ (
);

FILL FILL_1__11454_ (
);

FILL FILL_1__11034_ (
);

FILL FILL_0__8881_ (
);

FILL FILL_2__8899_ (
);

FILL FILL_0__8461_ (
);

FILL FILL_2__8479_ (
);

FILL FILL_0__10867_ (
);

FILL FILL_0__10447_ (
);

DFFPOSX1 _10732_ (
    .D(\Y[4] [1]),
    .CLK(clk_bF$buf12),
    .Q(\u_fir_pe4.rYin [1])
);

FILL FILL_2__8059_ (
);

FILL FILL_0__8041_ (
);

NAND2X1 _10312_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3589_)
);

FILL FILL_0__10027_ (
);

FILL FILL_2__9420_ (
);

INVX1 _7939_ (
    .A(\u_fir_pe1.mul [3]),
    .Y(_1446_)
);

NAND2X1 _7519_ (
    .A(vdd),
    .B(\X[1] [4]),
    .Y(_1038_)
);

FILL FILL_1__6896_ (
);

FILL FILL_1__6476_ (
);

FILL FILL_2__13246_ (
);

FILL FILL_3_CLKBUF1_insert21 (
);

FILL FILL_3_CLKBUF1_insert23 (
);

FILL FILL_1__12659_ (
);

FILL FILL_3_CLKBUF1_insert25 (
);

FILL FILL_1__12239_ (
);

FILL FILL_3_CLKBUF1_insert26 (
);

FILL FILL_3_CLKBUF1_insert28 (
);

FILL FILL_0__9666_ (
);

FILL FILL_3__7763_ (
);

FILL FILL_0__9246_ (
);

OAI21X1 _11937_ (
    .A(_5055_),
    .B(_5051_),
    .C(_4991_),
    .Y(_5056_)
);

OR2X2 _11517_ (
    .A(_4696_),
    .B(_4700_),
    .Y(_4701_)
);

FILL FILL_3__10593_ (
);

FILL FILL_1__8622_ (
);

FILL FILL_1__8202_ (
);

FILL FILL_3__8548_ (
);

NAND2X1 _7692_ (
    .A(vdd),
    .B(\X[1] [7]),
    .Y(_1209_)
);

NAND2X1 _7272_ (
    .A(gnd),
    .B(\X[1] [3]),
    .Y(_1584_)
);

FILL FILL_2__6965_ (
);

FILL FILL_2__6545_ (
);

NAND2X1 _11690_ (
    .A(\X[7] [0]),
    .B(vdd),
    .Y(_4812_)
);

AOI21X1 _11270_ (
    .A(gnd),
    .B(\X[5] [6]),
    .C(_4397_),
    .Y(_4466_)
);

FILL FILL_1__9827_ (
);

FILL FILL_1__9407_ (
);

FILL FILL_2__11732_ (
);

FILL FILL_2__11312_ (
);

NOR2X1 _8897_ (
    .A(\u_fir_pe2.rYin [10]),
    .B(\u_fir_pe2.mul [10]),
    .Y(_2321_)
);

NAND2X1 _8477_ (
    .A(\X[2] [4]),
    .B(gnd),
    .Y(_1915_)
);

NOR2X1 _8057_ (
    .A(_1560_),
    .B(_1559_),
    .Y(_1561_)
);

FILL FILL_1__10305_ (
);

FILL FILL_0__7732_ (
);

FILL FILL_0__7312_ (
);

FILL FILL_1__13197_ (
);

NAND3X1 _12895_ (
    .A(_5928_),
    .B(_5929_),
    .C(_5896_),
    .Y(_5933_)
);

DFFPOSX1 _12475_ (
    .D(_5572_[14]),
    .CLK(clk_bF$buf49),
    .Q(_6377_[14])
);

AOI21X1 _12055_ (
    .A(\X[7] [3]),
    .B(gnd),
    .C(_5169_),
    .Y(_5172_)
);

FILL FILL_3__13104_ (
);

FILL FILL_2__12937_ (
);

FILL FILL_2__12517_ (
);

FILL FILL_0__13131_ (
);

FILL FILL_0__8937_ (
);

FILL FILL_0__8517_ (
);

FILL FILL_1__9580_ (
);

FILL FILL_1__9160_ (
);

FILL FILL_2__7083_ (
);

NAND3X1 _6963_ (
    .A(_454_),
    .B(_556_),
    .C(_297_),
    .Y(_557_)
);

NAND2X1 _6543_ (
    .A(_141_),
    .B(_142_),
    .Y(_143_)
);

FILL FILL_2__12690_ (
);

FILL FILL_2__12270_ (
);

FILL FILL_1__11683_ (
);

FILL FILL_3__10229_ (
);

FILL FILL_1__11263_ (
);

FILL FILL_0__8690_ (
);

FILL FILL_0__8270_ (
);

FILL FILL_2__8288_ (
);

FILL FILL_0__10676_ (
);

NAND3X1 _10961_ (
    .A(_4158_),
    .B(_4160_),
    .C(_4159_),
    .Y(_4161_)
);

NAND2X1 _10541_ (
    .A(_3812_),
    .B(_3776_),
    .Y(_3813_)
);

FILL FILL_0__10256_ (
);

NAND2X1 _10121_ (
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3400_)
);

NOR2X1 _7748_ (
    .A(_812_),
    .B(_1259_),
    .Y(_1264_)
);

AOI22X1 _7328_ (
    .A(_806_),
    .B(_811_),
    .C(_846_),
    .D(_849_),
    .Y(_850_)
);

FILL FILL_2__13055_ (
);

FILL FILL_1__12888_ (
);

FILL FILL_1__12048_ (
);

FILL FILL_0__9895_ (
);

FILL FILL_3__7992_ (
);

FILL FILL_0__9475_ (
);

FILL FILL_0__9055_ (
);

NAND2X1 _11746_ (
    .A(gnd),
    .B(\X[7] [4]),
    .Y(_4867_)
);

FILL FILL_3__7152_ (
);

AND2X2 _11326_ (
    .A(_4520_),
    .B(_4517_),
    .Y(_4521_)
);

FILL FILL253950x176550 (
);

FILL FILL_0__12822_ (
);

FILL FILL_0__12402_ (
);

FILL FILL_1__8851_ (
);

FILL FILL_1__8431_ (
);

FILL FILL_1__8011_ (
);

FILL FILL_3__8777_ (
);

INVX1 _7081_ (
    .A(\u_fir_pe0.mul [5]),
    .Y(_666_)
);

FILL FILL_2__6774_ (
);

FILL FILL_3__11187_ (
);

FILL FILL_1__9636_ (
);

FILL FILL_1__9216_ (
);

FILL FILL_2__11961_ (
);

FILL FILL_2__11541_ (
);

FILL FILL_2__11121_ (
);

NAND2X1 _8286_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf3 ),
    .Y(_1726_)
);

FILL FILL_1__10954_ (
);

FILL FILL_1__10534_ (
);

FILL FILL_1__10114_ (
);

FILL FILL_0__7961_ (
);

FILL FILL_2__7979_ (
);

FILL FILL_2__7559_ (
);

FILL FILL_0__7541_ (
);

FILL FILL_2__7139_ (
);

FILL FILL_0__7121_ (
);

NAND3X1 _12284_ (
    .A(_5364_),
    .B(_5366_),
    .C(_5394_),
    .Y(_5396_)
);

FILL FILL_2__8920_ (
);

FILL FILL_2__8500_ (
);

FILL FILL_3__13333_ (
);

FILL FILL_2__12746_ (
);

FILL FILL_2__12326_ (
);

FILL FILL_1__11739_ (
);

FILL FILL_1__11319_ (
);

FILL FILL_0__8746_ (
);

FILL FILL_3__6843_ (
);

FILL FILL_0__8326_ (
);

FILL FILL_3__6423_ (
);

NAND2X1 _13069_ (
    .A(_5910_),
    .B(_5984_),
    .Y(_6104_)
);

FILL FILL_2__9705_ (
);

FILL FILL_1__7702_ (
);

FILL FILL_3__7628_ (
);

NAND3X1 _6772_ (
    .A(_300_),
    .B(_364_),
    .C(_365_),
    .Y(_370_)
);

FILL FILL_3__10458_ (
);

FILL FILL_1__11492_ (
);

FILL FILL_1__11072_ (
);

FILL FILL_0__10485_ (
);

NOR2X1 _10770_ (
    .A(_4735_),
    .B(_4725_),
    .Y(_4745_)
);

INVX1 _10350_ (
    .A(_3619_),
    .Y(_3627_)
);

FILL FILL_0__10065_ (
);

FILL FILL_1__8907_ (
);

FILL FILL_2__10812_ (
);

NOR2X1 _7977_ (
    .A(_1478_),
    .B(_1479_),
    .Y(_1480_)
);

NAND3X1 _7557_ (
    .A(_1074_),
    .B(_1075_),
    .C(_1073_),
    .Y(_1076_)
);

INVX1 _7137_ (
    .A(_719_),
    .Y(_721_)
);

FILL FILL_2__13284_ (
);

FILL FILL_0__6812_ (
);

FILL FILL_1__12697_ (
);

FILL FILL_1__12277_ (
);

FILL FILL_0__9284_ (
);

INVX1 _11975_ (
    .A(_5086_),
    .Y(_5093_)
);

FILL FILL_3__7381_ (
);

NOR2X1 _11555_ (
    .A(\u_fir_pe5.rYin [13]),
    .B(\u_fir_pe5.mul [13]),
    .Y(_4739_)
);

AOI21X1 _11135_ (
    .A(_4244_),
    .B(_4246_),
    .C(_4332_),
    .Y(_4333_)
);

FILL FILL_3__12604_ (
);

FILL FILL_0__12631_ (
);

FILL FILL_0__12211_ (
);

FILL FILL_1__7299_ (
);

NOR2X1 _9703_ (
    .A(\u_fir_pe3.rYin [4]),
    .B(\u_fir_pe3.mul [4]),
    .Y(_3049_)
);

FILL FILL_1__8660_ (
);

FILL FILL_1__8240_ (
);

FILL FILL_3__8166_ (
);

FILL FILL_0__13416_ (
);

FILL FILL_2__6583_ (
);

FILL FILL254250x150 (
);

FILL FILL_1__9445_ (
);

FILL FILL_1__9025_ (
);

FILL FILL_2__11770_ (
);

FILL FILL_2__11350_ (
);

DFFPOSX1 _8095_ (
    .D(\X[1] [3]),
    .CLK(clk_bF$buf1),
    .Q(\X[2] [3])
);

FILL FILL_1__10763_ (
);

FILL FILL_1__10343_ (
);

FILL FILL_2__7788_ (
);

FILL FILL_0__7770_ (
);

FILL FILL_0__7350_ (
);

FILL FILL_2__7368_ (
);

AOI21X1 _12093_ (
    .A(_5125_),
    .B(_5131_),
    .C(_5206_),
    .Y(_5210_)
);

NAND3X1 _6828_ (
    .A(_343_),
    .B(_349_),
    .C(_424_),
    .Y(_425_)
);

NAND3X1 _6408_ (
    .A(_0_),
    .B(_5_),
    .C(_3_),
    .Y(_11_)
);

FILL FILL_2__12975_ (
);

FILL FILL_2__12555_ (
);

FILL FILL_2__12135_ (
);

FILL FILL_1__11968_ (
);

FILL FILL_1__11548_ (
);

FILL FILL_1__11128_ (
);

FILL FILL_0__8555_ (
);

FILL FILL_3__6652_ (
);

FILL FILL_0__8135_ (
);

NAND3X1 _10826_ (
    .A(vdd),
    .B(\X[5] [1]),
    .C(_4027_),
    .Y(_4028_)
);

NAND3X1 _10406_ (
    .A(_3611_),
    .B(_3614_),
    .C(_3681_),
    .Y(_3682_)
);

INVX1 _13298_ (
    .A(\u_fir_pe7.mul [12]),
    .Y(_6322_)
);

FILL FILL_2__9934_ (
);

FILL FILL_2__9514_ (
);

FILL FILL_0__11902_ (
);

FILL FILL_1__7931_ (
);

FILL FILL_1__7511_ (
);

FILL FILL_3__7857_ (
);

FILL FILL_3__7017_ (
);

AOI21X1 _6581_ (
    .A(_171_),
    .B(_167_),
    .C(_152_),
    .Y(_181_)
);

FILL FILL_3__10687_ (
);

FILL FILL_0__10294_ (
);

FILL FILL_1__8716_ (
);

FILL FILL_2__10621_ (
);

FILL FILL_2__10201_ (
);

NOR2X1 _7786_ (
    .A(_1299_),
    .B(_1301_),
    .Y(_1302_)
);

OAI21X1 _7366_ (
    .A(_886_),
    .B(_812_),
    .C(_880_),
    .Y(_887_)
);

FILL FILL_2__13093_ (
);

FILL FILL_2__6639_ (
);

FILL FILL_0__6621_ (
);

FILL FILL_1__12086_ (
);

FILL FILL_0__9093_ (
);

NAND3X1 _11784_ (
    .A(_4836_),
    .B(_4893_),
    .C(_4897_),
    .Y(_4905_)
);

FILL FILL_0__11499_ (
);

FILL FILL_3__7190_ (
);

FILL FILL_0__11079_ (
);

NOR2X1 _11364_ (
    .A(_4550_),
    .B(_4554_),
    .Y(_4558_)
);

FILL FILL_3__12833_ (
);

FILL FILL_3__12413_ (
);

FILL FILL_2__11826_ (
);

FILL FILL_0__12860_ (
);

FILL FILL_2__11406_ (
);

FILL FILL_0__12440_ (
);

FILL FILL_0__12020_ (
);

FILL FILL_1__10819_ (
);

FILL FILL_0__7826_ (
);

NOR2X1 _9932_ (
    .A(_3212_),
    .B(_3213_),
    .Y(_3214_)
);

FILL FILL_0__7406_ (
);

AND2X2 _9512_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2868_)
);

AOI21X1 _12989_ (
    .A(_6025_),
    .B(_6024_),
    .C(_6017_),
    .Y(_6026_)
);

FILL FILL_3__8395_ (
);

OAI22X1 _12569_ (
    .A(_5609_),
    .B(_5610_),
    .C(_5579_),
    .D(_5583_),
    .Y(_5611_)
);

AND2X2 _12149_ (
    .A(_5258_),
    .B(_5264_),
    .Y(_5265_)
);

FILL FILL_0__13225_ (
);

FILL FILL_2__6392_ (
);

FILL FILL_1__9674_ (
);

FILL FILL_1__9254_ (
);

FILL FILL_1__10992_ (
);

FILL FILL_1__10572_ (
);

FILL FILL_1__10152_ (
);

FILL FILL_2__7597_ (
);

FILL FILL_2__7177_ (
);

OAI21X1 _6637_ (
    .A(_778_),
    .B(_235_),
    .C(_227_),
    .Y(_236_)
);

FILL FILL_2__12784_ (
);

FILL FILL_2__12364_ (
);

FILL FILL_1__11777_ (
);

FILL FILL_1__11357_ (
);

FILL FILL_0__8784_ (
);

FILL FILL_0__8364_ (
);

FILL FILL_3__6461_ (
);

OAI21X1 _10635_ (
    .A(_3897_),
    .B(_3894_),
    .C(_3896_),
    .Y(_3899_)
);

INVX2 _10215_ (
    .A(gnd),
    .Y(_3493_)
);

FILL FILL_2__9743_ (
);

FILL FILL_2__9323_ (
);

FILL FILL_0__11711_ (
);

FILL FILL_1__6799_ (
);

FILL FILL_1__6379_ (
);

FILL FILL_2__13149_ (
);

FILL FILL_1__7740_ (
);

FILL FILL_1__7320_ (
);

FILL FILL_0__9989_ (
);

FILL FILL_0__9569_ (
);

FILL FILL_0__9149_ (
);

INVX1 _6390_ (
    .A(_781_),
    .Y(_782_)
);

FILL FILL_0__12916_ (
);

FILL FILL_3__10076_ (
);

FILL FILL_1__8945_ (
);

FILL FILL_1__8525_ (
);

FILL FILL_2__10850_ (
);

FILL FILL_2__10430_ (
);

FILL FILL_2__10010_ (
);

AOI21X1 _7595_ (
    .A(_1053_),
    .B(_1050_),
    .C(_1036_),
    .Y(_1113_)
);

OAI21X1 _7175_ (
    .A(_751_),
    .B(_752_),
    .C(_756_),
    .Y(_758_)
);

FILL FILL_3__9812_ (
);

FILL FILL_2__6868_ (
);

FILL FILL_0__6850_ (
);

FILL FILL_0__6430_ (
);

FILL FILL_2__6448_ (
);

DFFPOSX1 _11593_ (
    .D(_4775_[9]),
    .CLK(clk_bF$buf35),
    .Q(\Y[6] [9])
);

OAI21X1 _11173_ (
    .A(_4300_),
    .B(_4369_),
    .C(_4339_),
    .Y(_4370_)
);

FILL FILL_2__11215_ (
);

FILL FILL_1__10628_ (
);

FILL FILL_1__10208_ (
);

FILL FILL_0__7635_ (
);

NOR2X1 _9741_ (
    .A(\u_fir_pe3.rYin [8]),
    .B(\u_fir_pe3.mul [8]),
    .Y(_3084_)
);

AND2X2 _9321_ (
    .A(_2676_),
    .B(_2679_),
    .Y(_2680_)
);

AOI21X1 _12798_ (
    .A(_5830_),
    .B(_5836_),
    .C(_5817_),
    .Y(_5837_)
);

AOI21X1 _12378_ (
    .A(_5477_),
    .B(_5480_),
    .C(_5479_),
    .Y(_5481_)
);

FILL FILL_0__13034_ (
);

FILL FILL_3__6517_ (
);

FILL FILL_1__9483_ (
);

FILL FILL_1__9063_ (
);

FILL FILL_1__10381_ (
);

FILL FILL_3__13180_ (
);

INVX2 _6866_ (
    .A(gnd),
    .Y(_462_)
);

NAND2X1 _6446_ (
    .A(_46_),
    .B(_47_),
    .Y(_48_)
);

FILL FILL_2__12593_ (
);

FILL FILL_2__12173_ (
);

FILL FILL_1__11166_ (
);

FILL FILL_0__8593_ (
);

FILL FILL_0__10999_ (
);

FILL FILL_3__6690_ (
);

FILL FILL_0__8173_ (
);

FILL FILL_0__10579_ (
);

NAND3X1 _10864_ (
    .A(\X[5] [1]),
    .B(vdd),
    .C(_4064_),
    .Y(_4065_)
);

AOI21X1 _10444_ (
    .A(_3670_),
    .B(_3713_),
    .C(_3716_),
    .Y(_3719_)
);

FILL FILL_0__10159_ (
);

NAND3X1 _10024_ (
    .A(_3300_),
    .B(_3294_),
    .C(_3298_),
    .Y(_3305_)
);

FILL FILL_3__11913_ (
);

FILL FILL_2__10906_ (
);

FILL FILL_2__9972_ (
);

FILL FILL_2__9552_ (
);

FILL FILL_0__11940_ (
);

FILL FILL_2__9132_ (
);

FILL FILL_0__11520_ (
);

FILL FILL_0__11100_ (
);

FILL FILL_0__6906_ (
);

FILL FILL_0__9798_ (
);

FILL FILL_0__9378_ (
);

FILL FILL_3__7475_ (
);

INVX2 _11649_ (
    .A(gnd),
    .Y(_5560_)
);

OAI21X1 _11229_ (
    .A(_4425_),
    .B(_4424_),
    .C(_4423_),
    .Y(_4426_)
);

FILL FILL_1__13312_ (
);

FILL FILL_0__12725_ (
);

FILL FILL_0__12305_ (
);

FILL FILL_1__8754_ (
);

FILL FILL_1__8334_ (
);

FILL FILL_3__9621_ (
);

FILL FILL_2__6677_ (
);

FILL FILL_1__9959_ (
);

FILL FILL_1__9539_ (
);

FILL FILL_1__9119_ (
);

FILL FILL_3__12031_ (
);

FILL FILL_2__11864_ (
);

FILL FILL_2__11444_ (
);

FILL FILL_2__11024_ (
);

NAND2X1 _8189_ (
    .A(_1629_),
    .B(_1630_),
    .Y(_1631_)
);

FILL FILL_1__10857_ (
);

FILL FILL_1__10437_ (
);

FILL FILL_1__10017_ (
);

FILL FILL_0__7864_ (
);

OAI21X1 _9970_ (
    .A(_3251_),
    .B(_3250_),
    .C(_3217_),
    .Y(_3252_)
);

FILL FILL_0__7444_ (
);

AOI21X1 _9550_ (
    .A(_2851_),
    .B(_2885_),
    .C(_2904_),
    .Y(_2905_)
);

FILL FILL_0__7024_ (
);

OAI21X1 _9130_ (
    .A(_2489_),
    .B(_2490_),
    .C(_2488_),
    .Y(_2491_)
);

NOR2X1 _12187_ (
    .A(_5199_),
    .B(_5244_),
    .Y(_5302_)
);

FILL FILL_2__8823_ (
);

FILL FILL_2__8403_ (
);

FILL FILL_2__12649_ (
);

FILL FILL_2__12229_ (
);

FILL FILL_0__13263_ (
);

FILL FILL_1__6820_ (
);

FILL FILL_1__6400_ (
);

FILL FILL_0__8649_ (
);

FILL FILL_3__6746_ (
);

FILL FILL_0__8229_ (
);

FILL FILL_1__9292_ (
);

FILL FILL_2_CLKBUF1_insert30 (
);

FILL FILL_2_CLKBUF1_insert31 (
);

FILL FILL_2__9608_ (
);

FILL FILL_2_CLKBUF1_insert32 (
);

FILL FILL_2_CLKBUF1_insert33 (
);

FILL FILL_2_CLKBUF1_insert34 (
);

FILL FILL_2_CLKBUF1_insert35 (
);

FILL FILL_2_CLKBUF1_insert36 (
);

FILL FILL_2_CLKBUF1_insert37 (
);

FILL FILL_2_CLKBUF1_insert38 (
);

FILL FILL_2_CLKBUF1_insert39 (
);

FILL FILL_1__10190_ (
);

FILL FILL_1__7605_ (
);

OAI21X1 _6675_ (
    .A(_273_),
    .B(_269_),
    .C(_209_),
    .Y(_274_)
);

FILL FILL254250x90150 (
);

FILL FILL_1__11395_ (
);

FILL FILL_0__10388_ (
);

AND2X2 _10673_ (
    .A(_3936_),
    .B(_3935_),
    .Y(_3978_[12])
);

NAND3X1 _10253_ (
    .A(_3511_),
    .B(_3526_),
    .C(_3527_),
    .Y(_3531_)
);

FILL FILL_3__11302_ (
);

FILL FILL_2__9781_ (
);

FILL FILL_2__9361_ (
);

FILL FILL_2__13187_ (
);

FILL FILL_0__6715_ (
);

OR2X2 _8821_ (
    .A(_2241_),
    .B(_2246_),
    .Y(_2248_)
);

INVX1 _8401_ (
    .A(_1834_),
    .Y(_1840_)
);

FILL FILL254250x57750 (
);

FILL FILL_0__9187_ (
);

OAI21X1 _11878_ (
    .A(_4921_),
    .B(_4996_),
    .C(_4925_),
    .Y(_4997_)
);

NOR2X1 _11458_ (
    .A(_4643_),
    .B(_4642_),
    .Y(_4644_)
);

AOI22X1 _11038_ (
    .A(_4072_),
    .B(_4143_),
    .C(_4146_),
    .D(_4142_),
    .Y(_4237_)
);

FILL FILL_3__12927_ (
);

FILL FILL_1__13121_ (
);

FILL FILL_0__12954_ (
);

FILL FILL_0__12534_ (
);

FILL FILL_0__12114_ (
);

AOI21X1 _9606_ (
    .A(gnd),
    .B(_2957_),
    .C(_2959_),
    .Y(_2960_)
);

FILL FILL_1__8563_ (
);

FILL FILL_1__8143_ (
);

FILL FILL253950x108150 (
);

FILL FILL_3__8489_ (
);

FILL FILL_3__8069_ (
);

FILL FILL_3__9010_ (
);

FILL FILL_0__13319_ (
);

FILL FILL_2__6486_ (
);

FILL FILL_1__9768_ (
);

FILL FILL_1__9348_ (
);

FILL FILL_3__12680_ (
);

FILL FILL_3__12260_ (
);

FILL FILL_2__11673_ (
);

FILL FILL_2__11253_ (
);

FILL FILL_1__10666_ (
);

FILL FILL_1__10246_ (
);

FILL FILL_0__7673_ (
);

FILL FILL254550x201750 (
);

FILL FILL_2__8632_ (
);

FILL FILL_2__8212_ (
);

FILL FILL_0__10600_ (
);

FILL FILL_3__13045_ (
);

FILL FILL_2__12878_ (
);

FILL FILL_2__12458_ (
);

FILL FILL_2__12038_ (
);

FILL FILL_0__13072_ (
);

FILL FILL_0__8878_ (
);

FILL FILL_0__8458_ (
);

DFFPOSX1 _10729_ (
    .D(\X[4] [6]),
    .CLK(clk_bF$buf3),
    .Q(\X[5] [6])
);

FILL FILL_0__8038_ (
);

NOR2X1 _10309_ (
    .A(_3320_),
    .B(_3509_),
    .Y(_3586_)
);

FILL FILL_1__12812_ (
);

FILL FILL_2__9417_ (
);

FILL FILL_0__11805_ (
);

FILL FILL_1__7834_ (
);

FILL FILL_1__7414_ (
);

NAND2X1 _6484_ (
    .A(gnd),
    .B(Xin[4]),
    .Y(_85_)
);

FILL FILL_3__8701_ (
);

NOR2X1 _10482_ (
    .A(_3755_),
    .B(_3754_),
    .Y(_3756_)
);

FILL FILL_0__10197_ (
);

AOI22X1 _10062_ (
    .A(gnd),
    .B(\X[4] [2]),
    .C(gnd),
    .D(\X[4] [3]),
    .Y(_3342_)
);

FILL FILL_1__8619_ (
);

FILL FILL_3__11531_ (
);

FILL FILL_2__10944_ (
);

FILL FILL_2__9590_ (
);

FILL FILL_2__10524_ (
);

FILL FILL_2__9170_ (
);

FILL FILL_2__10104_ (
);

AOI22X1 _7689_ (
    .A(_1039_),
    .B(_1205_),
    .C(_1131_),
    .D(_1127_),
    .Y(_1206_)
);

NOR2X1 _7269_ (
    .A(_1580_),
    .B(_1579_),
    .Y(_1581_)
);

FILL FILL_0__6944_ (
);

FILL FILL_0__6524_ (
);

OAI21X1 _8630_ (
    .A(_2013_),
    .B(_2065_),
    .C(_2001_),
    .Y(_2066_)
);

NAND2X1 _8210_ (
    .A(_1648_),
    .B(_1651_),
    .Y(_1652_)
);

AOI22X1 _11687_ (
    .A(\X[7] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[7] [4]),
    .Y(_4809_)
);

FILL FILL_3__7093_ (
);

AND2X2 _11267_ (
    .A(\X[5]_5_bF$buf0 ),
    .B(gnd),
    .Y(_4463_)
);

FILL FILL_2__7903_ (
);

FILL FILL_3__12316_ (
);

FILL FILL_2__11729_ (
);

FILL FILL_0__12763_ (
);

FILL FILL_2__11309_ (
);

FILL FILL_0__12343_ (
);

FILL FILL_0__7729_ (
);

DFFPOSX1 _9835_ (
    .D(_3181_[5]),
    .CLK(clk_bF$buf38),
    .Q(\Y[4] [5])
);

FILL FILL_0__7309_ (
);

AOI21X1 _9415_ (
    .A(_2752_),
    .B(_2751_),
    .C(_2694_),
    .Y(_2772_)
);

FILL FILL_1__8792_ (
);

FILL FILL_1__8372_ (
);

FILL FILL_0__13128_ (
);

BUFX2 _13413_ (
    .A(_6377_[5]),
    .Y(Yout[5])
);

FILL FILL_1__9997_ (
);

FILL FILL_1__9577_ (
);

FILL FILL_1__9157_ (
);

FILL FILL_2__11482_ (
);

FILL FILL_2__11062_ (
);

FILL FILL_1__10895_ (
);

FILL FILL_1__10475_ (
);

FILL FILL_1__10055_ (
);

FILL FILL_0__7482_ (
);

FILL FILL_0__7062_ (
);

FILL FILL_3__10802_ (
);

FILL FILL_2__8861_ (
);

FILL FILL_2__8441_ (
);

FILL FILL_3__13274_ (
);

FILL FILL_2__8021_ (
);

FILL FILL_2__12687_ (
);

FILL FILL_2__12267_ (
);

OAI21X1 _7901_ (
    .A(_1381_),
    .B(_1406_),
    .C(_1405_),
    .Y(_1413_)
);

FILL FILL_0__8687_ (
);

FILL FILL_3__6784_ (
);

FILL FILL_0__8267_ (
);

NAND2X1 _10958_ (
    .A(_4136_),
    .B(_4132_),
    .Y(_4158_)
);

OAI21X1 _10538_ (
    .A(_3804_),
    .B(_3803_),
    .C(_3809_),
    .Y(_3810_)
);

OAI21X1 _10118_ (
    .A(_3324_),
    .B(_3396_),
    .C(_3365_),
    .Y(_3397_)
);

FILL FILL_1__12621_ (
);

FILL FILL_1__12201_ (
);

FILL FILL_2__9646_ (
);

FILL FILL_2__9226_ (
);

FILL FILL_1__7643_ (
);

FILL FILL_3__7569_ (
);

FILL FILL_1__13406_ (
);

FILL FILL_3__8930_ (
);

FILL FILL_0__12819_ (
);

FILL FILL_3__10399_ (
);

AOI21X1 _10291_ (
    .A(_3485_),
    .B(_3555_),
    .C(_3567_),
    .Y(_3568_)
);

FILL FILL_1__8848_ (
);

FILL FILL_3__11760_ (
);

FILL FILL_1__8428_ (
);

FILL FILL_1__8008_ (
);

FILL FILL_2__10333_ (
);

NOR2X1 _7498_ (
    .A(_1010_),
    .B(_1012_),
    .Y(_1017_)
);

AND2X2 _7078_ (
    .A(_663_),
    .B(_662_),
    .Y(_790_[4])
);

FILL FILL_3__9715_ (
);

FILL FILL_0__6753_ (
);

NAND2X1 _11496_ (
    .A(_4642_),
    .B(_4654_),
    .Y(_4679_)
);

OAI21X1 _11076_ (
    .A(_4192_),
    .B(_4189_),
    .C(_4274_),
    .Y(_4275_)
);

FILL FILL_2__7712_ (
);

FILL FILL_3__12545_ (
);

FILL FILL_3__12125_ (
);

FILL FILL_2__11958_ (
);

FILL FILL_0__12992_ (
);

FILL FILL_2__11538_ (
);

FILL FILL_0__12572_ (
);

FILL FILL_2__11118_ (
);

FILL FILL_0__12152_ (
);

FILL FILL_0__7958_ (
);

FILL FILL_0__7538_ (
);

OAI21X1 _9644_ (
    .A(_2954_),
    .B(_2967_),
    .C(_2971_),
    .Y(_2997_)
);

FILL FILL_0__7118_ (
);

AOI21X1 _9224_ (
    .A(_2583_),
    .B(_2582_),
    .C(_2581_),
    .Y(_2584_)
);

FILL FILL_1__8181_ (
);

FILL FILL_2__8917_ (
);

NOR2X1 _13222_ (
    .A(\u_fir_pe7.rYin [5]),
    .B(\u_fir_pe7.mul [5]),
    .Y(_6247_)
);

FILL FILL_1__6914_ (
);

FILL FILL_1__9386_ (
);

FILL FILL_2__11291_ (
);

FILL FILL_1__10284_ (
);

FILL FILL_0__7291_ (
);

FILL FILL_3__10611_ (
);

FILL FILL_2__8670_ (
);

FILL FILL_2__8250_ (
);

OAI21X1 _6769_ (
    .A(_366_),
    .B(_363_),
    .C(_299_),
    .Y(_367_)
);

FILL FILL_2__12076_ (
);

OAI21X1 _7710_ (
    .A(_1226_),
    .B(_1225_),
    .C(_1224_),
    .Y(_1227_)
);

FILL FILL_1__11489_ (
);

FILL FILL_1__11069_ (
);

FILL FILL_0__8496_ (
);

NAND2X1 _10767_ (
    .A(gnd),
    .B(\X[5] [1]),
    .Y(_4716_)
);

OAI21X1 _10347_ (
    .A(_3623_),
    .B(_3622_),
    .C(_3621_),
    .Y(_3624_)
);

FILL FILL_1__12850_ (
);

FILL FILL_1__12430_ (
);

FILL FILL_1__12010_ (
);

FILL FILL_2__10809_ (
);

FILL FILL_2__9455_ (
);

FILL FILL_0__11843_ (
);

FILL FILL_2__9035_ (
);

FILL FILL_0__11423_ (
);

FILL FILL_0__11003_ (
);

FILL FILL_0__6809_ (
);

NOR2X1 _8915_ (
    .A(\u_fir_pe2.rYin [12]),
    .B(\u_fir_pe2.mul [12]),
    .Y(_2339_)
);

FILL FILL_1__7872_ (
);

FILL FILL_1__7452_ (
);

FILL FILL_1__7032_ (
);

FILL FILL_3__7798_ (
);

FILL FILL_1__13215_ (
);

NAND3X1 _12913_ (
    .A(_5948_),
    .B(_5949_),
    .C(_5950_),
    .Y(_5951_)
);

FILL FILL_0__12628_ (
);

FILL FILL_0__12208_ (
);

FILL FILL_1__8657_ (
);

FILL FILL_1__8237_ (
);

FILL FILL_2__10982_ (
);

FILL FILL_2__10562_ (
);

FILL FILL_2__10142_ (
);

FILL FILL_3__9944_ (
);

FILL FILL_3__9104_ (
);

FILL FILL_0__6982_ (
);

FILL FILL_0__6562_ (
);

FILL FILL_2__7941_ (
);

FILL FILL_3__12774_ (
);

FILL FILL_2__7521_ (
);

FILL FILL_3__12354_ (
);

FILL FILL_2__7101_ (
);

FILL FILL_2__11767_ (
);

FILL FILL_2__11347_ (
);

FILL FILL_0__12381_ (
);

FILL FILL_0__7767_ (
);

DFFPOSX1 _9873_ (
    .D(_3185_[3]),
    .CLK(clk_bF$buf42),
    .Q(\u_fir_pe3.mul [3])
);

FILL FILL_0__7347_ (
);

OAI21X1 _9453_ (
    .A(_2416_),
    .B(_2807_),
    .C(_2809_),
    .Y(_2810_)
);

INVX1 _9033_ (
    .A(_2395_),
    .Y(_2396_)
);

FILL FILL_1__11701_ (
);

FILL FILL_2__8726_ (
);

FILL FILL_2__8306_ (
);

FILL FILL_3__13139_ (
);

FILL FILL_0__13166_ (
);

NAND2X1 _13031_ (
    .A(_6048_),
    .B(_6045_),
    .Y(_6067_)
);

FILL FILL_1__6723_ (
);

FILL FILL_1__9195_ (
);

FILL FILL_1__12906_ (
);

FILL FILL_0__9913_ (
);

FILL FILL_1__10093_ (
);

FILL FILL_1__7928_ (
);

FILL FILL_1__7508_ (
);

FILL FILL_3__10000_ (
);

NOR2X1 _6998_ (
    .A(_560_),
    .B(_583_),
    .Y(_591_)
);

INVX1 _6578_ (
    .A(_96_),
    .Y(_178_)
);

FILL FILL_1__11298_ (
);

NAND2X1 _10996_ (
    .A(\X[5] [0]),
    .B(gnd),
    .Y(_4195_)
);

NAND2X1 _10576_ (
    .A(_3841_),
    .B(_3842_),
    .Y(_3978_[3])
);

NAND2X1 _10156_ (
    .A(_3346_),
    .B(_3430_),
    .Y(_3435_)
);

FILL FILL_2__9684_ (
);

FILL FILL_2__10618_ (
);

FILL FILL_2__9264_ (
);

FILL FILL_0__11652_ (
);

FILL FILL_0__11232_ (
);

FILL FILL_0__6618_ (
);

INVX1 _8724_ (
    .A(_2120_),
    .Y(_2158_)
);

NAND2X1 _8304_ (
    .A(_1743_),
    .B(_1735_),
    .Y(_1744_)
);

FILL FILL_1__7681_ (
);

FILL FILL_1__7261_ (
);

FILL FILL_3__7187_ (
);

FILL FILL_1__13024_ (
);

FILL FILL_0__12857_ (
);

NAND3X1 _12722_ (
    .A(_5715_),
    .B(_5756_),
    .C(_5761_),
    .Y(_5762_)
);

FILL FILL_0__12437_ (
);

FILL FILL_0__12017_ (
);

NAND2X1 _12302_ (
    .A(_5412_),
    .B(_5411_),
    .Y(_5578_[15])
);

NOR2X1 _9929_ (
    .A(_3211_),
    .B(_3210_),
    .Y(_3982_[3])
);

NOR2X1 _9509_ (
    .A(_2864_),
    .B(_2807_),
    .Y(_2865_)
);

FILL FILL_1__8886_ (
);

FILL FILL_1__8466_ (
);

FILL FILL_1__8046_ (
);

FILL FILL_2__10791_ (
);

FILL FILL_2__10371_ (
);

FILL FILL_3__9753_ (
);

FILL FILL_3__9333_ (
);

FILL FILL_0__6791_ (
);

FILL FILL_2__6389_ (
);

FILL FILL_2__7750_ (
);

FILL FILL_2__7330_ (
);

FILL FILL_2__11996_ (
);

FILL FILL_2__11576_ (
);

FILL FILL_2__11156_ (
);

FILL FILL_0__12190_ (
);

FILL FILL_1__10989_ (
);

FILL FILL_1__10569_ (
);

FILL FILL_1__10149_ (
);

FILL FILL_0__7996_ (
);

FILL FILL_0__7576_ (
);

NOR2X1 _9682_ (
    .A(_3030_),
    .B(_3029_),
    .Y(_3181_[1])
);

FILL FILL_0__7156_ (
);

AOI22X1 _9262_ (
    .A(gnd),
    .B(\X[3] [7]),
    .C(\X[3] [3]),
    .D(gnd),
    .Y(_2621_)
);

FILL FILL_1__11930_ (
);

FILL FILL_1__11510_ (
);

FILL FILL_2__8535_ (
);

FILL FILL_0__10923_ (
);

FILL FILL_0__10503_ (
);

FILL FILL_0__13395_ (
);

NOR2X1 _13260_ (
    .A(_6272_),
    .B(_6271_),
    .Y(_6284_)
);

FILL FILL_1__6952_ (
);

FILL FILL_1__6532_ (
);

FILL FILL_2__13302_ (
);

FILL FILL_3__6878_ (
);

FILL FILL_3__6458_ (
);

FILL FILL_1__12715_ (
);

FILL FILL_0__9722_ (
);

FILL FILL_0__9302_ (
);

FILL FILL_0__11708_ (
);

FILL FILL_1__7737_ (
);

FILL FILL_1__7317_ (
);

INVX2 _6387_ (
    .A(gnd),
    .Y(_778_)
);

NAND2X1 _10385_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3661_)
);

FILL FILL_3__11854_ (
);

FILL FILL_2__6601_ (
);

FILL FILL_3__11014_ (
);

FILL FILL_2__10847_ (
);

FILL FILL_2__9493_ (
);

FILL FILL_0__11881_ (
);

FILL FILL_2__10427_ (
);

FILL FILL_2__9073_ (
);

FILL FILL_0__11461_ (
);

FILL FILL_2__10007_ (
);

FILL FILL_0__11041_ (
);

FILL FILL_3__9809_ (
);

FILL FILL_0__6847_ (
);

DFFPOSX1 _8953_ (
    .D(_2383_[0]),
    .CLK(clk_bF$buf56),
    .Q(\Y[3] [0])
);

FILL FILL_0__6427_ (
);

AND2X2 _8533_ (
    .A(_1961_),
    .B(_1966_),
    .Y(_1971_)
);

DFFPOSX1 _8113_ (
    .D(\Y[1] [13]),
    .CLK(clk_bF$buf32),
    .Q(\u_fir_pe1.rYin [13])
);

FILL FILL_1__7490_ (
);

FILL FILL_1__7070_ (
);

FILL FILL_2__7806_ (
);

FILL FILL_3__12639_ (
);

FILL FILL_1__13253_ (
);

AOI22X1 _12951_ (
    .A(_5821_),
    .B(_5987_),
    .C(_5913_),
    .D(_5909_),
    .Y(_5988_)
);

FILL FILL_0__12666_ (
);

FILL FILL_0__12246_ (
);

NOR2X1 _12531_ (
    .A(_6362_),
    .B(_6361_),
    .Y(_6363_)
);

NAND3X1 _12111_ (
    .A(_5208_),
    .B(_5212_),
    .C(_5215_),
    .Y(_5228_)
);

INVX1 _9738_ (
    .A(\u_fir_pe3.rYin [8]),
    .Y(_3081_)
);

NAND3X1 _9318_ (
    .A(_2672_),
    .B(_2673_),
    .C(_2674_),
    .Y(_2677_)
);

FILL FILL_1__8695_ (
);

FILL FILL_1__8275_ (
);

FILL FILL_2__10180_ (
);

FILL FILL_3__9562_ (
);

INVX1 _13316_ (
    .A(\u_fir_pe7.mul [14]),
    .Y(_6340_)
);

FILL FILL_1_CLKBUF1_insert40 (
);

FILL FILL_1_CLKBUF1_insert41 (
);

FILL FILL_1_CLKBUF1_insert42 (
);

FILL FILL_1_CLKBUF1_insert43 (
);

FILL FILL_1_CLKBUF1_insert44 (
);

FILL FILL_1_CLKBUF1_insert45 (
);

FILL FILL_1_CLKBUF1_insert46 (
);

FILL FILL_1_CLKBUF1_insert47 (
);

FILL FILL_1_CLKBUF1_insert48 (
);

FILL FILL_1_CLKBUF1_insert49 (
);

FILL FILL_2__11385_ (
);

FILL FILL_1__10798_ (
);

FILL FILL_1__10378_ (
);

FILL FILL_0__7385_ (
);

AOI21X1 _9491_ (
    .A(_2832_),
    .B(_2828_),
    .C(_2773_),
    .Y(_2847_)
);

NAND2X1 _9071_ (
    .A(gnd),
    .B(\X[3] [2]),
    .Y(_2433_)
);

FILL FILL_3__10705_ (
);

FILL FILL_2__8764_ (
);

FILL FILL_2__8344_ (
);

FILL FILL_0__10312_ (
);

OAI21X1 _7804_ (
    .A(_871_),
    .B(_1102_),
    .C(_1276_),
    .Y(_1319_)
);

FILL FILL_1__6761_ (
);

FILL FILL_2__13111_ (
);

FILL FILL_3__6687_ (
);

FILL FILL_1__12944_ (
);

FILL FILL_1__12524_ (
);

FILL FILL_1__12104_ (
);

FILL FILL_2__9969_ (
);

FILL FILL_0__9951_ (
);

FILL FILL_2__9549_ (
);

FILL FILL_0__9531_ (
);

FILL FILL_0__11937_ (
);

FILL FILL_2__9129_ (
);

FILL FILL_0__9111_ (
);

INVX1 _11802_ (
    .A(_4921_),
    .Y(_4922_)
);

FILL FILL_0__11517_ (
);

FILL FILL_1__7966_ (
);

FILL FILL_1__7546_ (
);

FILL FILL_1__7126_ (
);

FILL FILL_1__13309_ (
);

FILL FILL_3__8413_ (
);

OAI21X1 _10194_ (
    .A(_3472_),
    .B(_3468_),
    .C(_3384_),
    .Y(_3473_)
);

FILL FILL_2__6830_ (
);

FILL FILL_2__6410_ (
);

FILL FILL_3__11243_ (
);

FILL FILL_2__10656_ (
);

FILL FILL_0__11690_ (
);

FILL FILL_2__10236_ (
);

FILL FILL_0__11270_ (
);

FILL FILL_0__6656_ (
);

NAND2X1 _8762_ (
    .A(_2193_),
    .B(_2194_),
    .Y(_2195_)
);

AOI22X1 _8342_ (
    .A(_1705_),
    .B(_1700_),
    .C(_1777_),
    .D(_1781_),
    .Y(_1782_)
);

AND2X2 _11399_ (
    .A(_4588_),
    .B(_4587_),
    .Y(_4592_)
);

FILL FILL_3__12868_ (
);

FILL FILL_2__7615_ (
);

FILL FILL_3__12448_ (
);

FILL FILL_3__12028_ (
);

FILL FILL_1__13062_ (
);

FILL FILL_0__12895_ (
);

NOR2X1 _12760_ (
    .A(_5792_),
    .B(_5794_),
    .Y(_5799_)
);

FILL FILL_0__12055_ (
);

AND2X2 _12340_ (
    .A(_5445_),
    .B(_5444_),
    .Y(_5572_[4])
);

FILL FILL_2__12802_ (
);

NAND3X1 _9967_ (
    .A(_3216_),
    .B(_3233_),
    .C(_3236_),
    .Y(_3249_)
);

NAND3X1 _9547_ (
    .A(_2886_),
    .B(_2892_),
    .C(_2850_),
    .Y(_2902_)
);

INVX1 _9127_ (
    .A(_2475_),
    .Y(_2488_)
);

FILL FILL_0__8802_ (
);

FILL FILL_3__9371_ (
);

NAND3X1 _13125_ (
    .A(_6140_),
    .B(_6157_),
    .C(_6156_),
    .Y(_6159_)
);

FILL FILL_1__6817_ (
);

FILL FILL_1__9289_ (
);

FILL FILL_2__11194_ (
);

FILL FILL_1__10187_ (
);

FILL FILL_0__7194_ (
);

FILL FILL_2__8573_ (
);

FILL FILL_0__10961_ (
);

FILL FILL_2__8153_ (
);

FILL FILL_0__10541_ (
);

FILL FILL_0__10121_ (
);

FILL FILL_2__12399_ (
);

NAND2X1 _7613_ (
    .A(_1122_),
    .B(_1130_),
    .Y(_1131_)
);

FILL FILL_1__6990_ (
);

FILL FILL_1__6570_ (
);

FILL FILL_0__8399_ (
);

FILL FILL_1__12753_ (
);

FILL FILL_1__12333_ (
);

FILL FILL_0__9760_ (
);

FILL FILL_2__9778_ (
);

FILL FILL_2__9358_ (
);

FILL FILL_0__9340_ (
);

FILL FILL_0__11746_ (
);

DFFPOSX1 _11611_ (
    .D(\Y[5] [3]),
    .CLK(clk_bF$buf39),
    .Q(\u_fir_pe5.rYin [3])
);

FILL FILL_0__11326_ (
);

NOR2X1 _8818_ (
    .A(\u_fir_pe2.rYin [3]),
    .B(\u_fir_pe2.mul [3]),
    .Y(_2245_)
);

FILL FILL_1__7775_ (
);

FILL FILL_1__7355_ (
);

FILL FILL_1__13118_ (
);

FILL FILL_3__8642_ (
);

AOI21X1 _12816_ (
    .A(_5763_),
    .B(_5761_),
    .C(_5854_),
    .Y(_5855_)
);

FILL FILL_3__11472_ (
);

FILL FILL_2__10885_ (
);

FILL FILL_2__10465_ (
);

FILL FILL_2__10045_ (
);

FILL FILL_1__9921_ (
);

FILL FILL_1__9501_ (
);

FILL FILL_3__9427_ (
);

FILL FILL_0__6885_ (
);

DFFPOSX1 _8991_ (
    .D(\Y[2] [14]),
    .CLK(clk_bF$buf0),
    .Q(\u_fir_pe2.rYin [14])
);

FILL FILL_0__6465_ (
);

NAND2X1 _8571_ (
    .A(_2007_),
    .B(_2003_),
    .Y(_2008_)
);

NAND2X1 _8151_ (
    .A(gnd),
    .B(\X[2] [2]),
    .Y(_1594_)
);

FILL FILL_2__7844_ (
);

FILL FILL_2__7424_ (
);

FILL FILL_2__7004_ (
);

FILL FILL_1__13291_ (
);

FILL FILL_0__12284_ (
);

FILL FILL_2__12611_ (
);

NAND2X1 _9776_ (
    .A(_3119_),
    .B(_3114_),
    .Y(_3120_)
);

OAI21X1 _9356_ (
    .A(_2631_),
    .B(_2639_),
    .C(_2638_),
    .Y(_2714_)
);

FILL FILL_2__8629_ (
);

FILL FILL_0__8611_ (
);

FILL FILL_2__8209_ (
);

FILL FILL_3__9180_ (
);

FILL FILL_0__13069_ (
);

DFFPOSX1 _13354_ (
    .D(\X[6] [0]),
    .CLK(clk_bF$buf2),
    .Q(\X[7] [0])
);

FILL FILL_1__6626_ (
);

FILL FILL_1__9098_ (
);

FILL FILL_1__12809_ (
);

FILL FILL_0__9816_ (
);

FILL FILL_3__10323_ (
);

FILL FILL_2__8382_ (
);

FILL FILL_0__10770_ (
);

FILL FILL_0__10350_ (
);

AOI21X1 _7842_ (
    .A(_1353_),
    .B(_1254_),
    .C(_1355_),
    .Y(_1356_)
);

NAND2X1 _7422_ (
    .A(\X[1] [2]),
    .B(gnd),
    .Y(_942_)
);

NOR2X1 _7002_ (
    .A(_235_),
    .B(_462_),
    .Y(_595_)
);

NAND3X1 _10899_ (
    .A(_4097_),
    .B(_4098_),
    .C(_4099_),
    .Y(_4100_)
);

NOR2X1 _10479_ (
    .A(_3262_),
    .B(_3650_),
    .Y(_3753_)
);

NAND3X1 _10059_ (
    .A(_3327_),
    .B(_3336_),
    .C(_3338_),
    .Y(_3339_)
);

FILL FILL_3__11948_ (
);

FILL FILL_1__12982_ (
);

FILL FILL_1__12562_ (
);

FILL FILL_3__11108_ (
);

FILL FILL_1__12142_ (
);

FILL FILL_0__11975_ (
);

FILL FILL_2__9587_ (
);

FILL FILL_2__9167_ (
);

INVX1 _11840_ (
    .A(_4878_),
    .Y(_4960_)
);

FILL FILL_0__11555_ (
);

INVX1 _11420_ (
    .A(_4606_),
    .Y(_4612_)
);

FILL FILL_0__11135_ (
);

AND2X2 _11000_ (
    .A(_4130_),
    .B(_4134_),
    .Y(_4199_)
);

NAND3X1 _8627_ (
    .A(_2061_),
    .B(_2058_),
    .C(_2062_),
    .Y(_2063_)
);

NAND2X1 _8207_ (
    .A(_1603_),
    .B(_1608_),
    .Y(_1649_)
);

FILL FILL_1__7584_ (
);

FILL FILL_1__7164_ (
);

FILL FILL_3__8871_ (
);

AND2X2 _12625_ (
    .A(vdd),
    .B(\X[6] [3]),
    .Y(_5666_)
);

FILL FILL_3__8031_ (
);

AOI21X1 _12205_ (
    .A(_5197_),
    .B(_5189_),
    .C(_5267_),
    .Y(_5320_)
);

FILL FILL_1__8789_ (
);

FILL FILL_1__8369_ (
);

FILL FILL_2__10694_ (
);

FILL FILL_2__10274_ (
);

FILL FILL_1__9730_ (
);

FILL FILL_1__9310_ (
);

FILL FILL_3__9656_ (
);

FILL FILL_0__6694_ (
);

NAND2X1 _8380_ (
    .A(\X[2] [2]),
    .B(gnd),
    .Y(_1819_)
);

FILL FILL_2__7653_ (
);

FILL FILL_3__12066_ (
);

FILL FILL_2__11899_ (
);

FILL FILL_2__11479_ (
);

FILL FILL_2__11059_ (
);

FILL FILL_0__12093_ (
);

FILL FILL_2__12840_ (
);

FILL FILL_2__12420_ (
);

FILL FILL_0__7899_ (
);

FILL FILL_2__12000_ (
);

FILL FILL_0__7479_ (
);

AOI21X1 _9585_ (
    .A(_2878_),
    .B(_2882_),
    .C(_2852_),
    .Y(_2940_)
);

FILL FILL_0__7059_ (
);

OR2X2 _9165_ (
    .A(_2524_),
    .B(_2522_),
    .Y(_2525_)
);

FILL FILL_1__11833_ (
);

FILL FILL_1__11413_ (
);

FILL FILL_0__8840_ (
);

FILL FILL_2__8858_ (
);

FILL FILL_0__8420_ (
);

FILL FILL_2__8438_ (
);

FILL FILL_0__10826_ (
);

FILL FILL_0__10406_ (
);

FILL FILL_0__8000_ (
);

FILL FILL_2__8018_ (
);

FILL FILL_0__13298_ (
);

OAI21X1 _13163_ (
    .A(_6163_),
    .B(_6188_),
    .C(_6187_),
    .Y(_6195_)
);

FILL FILL_1__6855_ (
);

FILL FILL_1__6435_ (
);

FILL FILL_2__13205_ (
);

FILL FILL_1__12618_ (
);

FILL FILL_0__9625_ (
);

FILL FILL_3__7722_ (
);

FILL FILL_0__9205_ (
);

FILL FILL_3__7302_ (
);

FILL FILL_3__10972_ (
);

FILL FILL_3__10552_ (
);

FILL FILL_2__8191_ (
);

BUFX2 BUFX2_insert10 (
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf1 )
);

BUFX2 BUFX2_insert11 (
    .A(\X[5] [5]),
    .Y(\X[5]_5_bF$buf0 )
);

FILL FILL_3__8507_ (
);

NAND3X1 _7651_ (
    .A(_1166_),
    .B(_1167_),
    .C(_1168_),
    .Y(_1169_)
);

DFFPOSX1 _7231_ (
    .D(Yin[8]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.rYin [8])
);

NAND2X1 _10288_ (
    .A(_3565_),
    .B(_3564_),
    .Y(_3566_)
);

FILL FILL_2__6924_ (
);

FILL FILL_2__6504_ (
);

FILL FILL_1__12791_ (
);

FILL FILL_3__11337_ (
);

FILL FILL_1__12371_ (
);

FILL FILL_2__9396_ (
);

FILL FILL_0__11784_ (
);

FILL FILL_0__11364_ (
);

OAI21X1 _8856_ (
    .A(_2277_),
    .B(_2278_),
    .C(_2274_),
    .Y(_2279_)
);

INVX1 _8436_ (
    .A(_1729_),
    .Y(_1875_)
);

INVX1 _8016_ (
    .A(_1519_),
    .Y(_1520_)
);

FILL FILL_1__7393_ (
);

FILL FILL_2__7709_ (
);

FILL FILL_1__13156_ (
);

FILL FILL_0__12989_ (
);

NAND2X1 _12854_ (
    .A(_5885_),
    .B(_5886_),
    .Y(_5892_)
);

FILL FILL_0__12569_ (
);

FILL FILL_3__8260_ (
);

FILL FILL_0__12149_ (
);

NAND2X1 _12434_ (
    .A(_5537_),
    .B(_5531_),
    .Y(_5538_)
);

NAND3X1 _12014_ (
    .A(_5104_),
    .B(_5122_),
    .C(_5118_),
    .Y(_5132_)
);

FILL FILL_1__8598_ (
);

FILL FILL_1__8178_ (
);

FILL FILL_3__11090_ (
);

FILL FILL_2__10083_ (
);

FILL FILL_3__9045_ (
);

INVX1 _13219_ (
    .A(\u_fir_pe7.rYin [5]),
    .Y(_6244_)
);

FILL FILL_2__7882_ (
);

FILL FILL_2__7462_ (
);

FILL FILL_3__12295_ (
);

FILL FILL_2__7042_ (
);

FILL FILL_2__11288_ (
);

NOR3X1 _6922_ (
    .A(_305_),
    .B(_473_),
    .C(_416_),
    .Y(_517_)
);

OAI21X1 _6502_ (
    .A(_98_),
    .B(_99_),
    .C(_84_),
    .Y(_103_)
);

FILL FILL_0__7288_ (
);

NAND3X1 _9394_ (
    .A(_2706_),
    .B(_2737_),
    .C(_2742_),
    .Y(_2752_)
);

FILL FILL_1__11642_ (
);

FILL FILL_1__11222_ (
);

FILL FILL_2__8667_ (
);

FILL FILL_2__8247_ (
);

FILL FILL_0__10635_ (
);

NAND2X1 _10920_ (
    .A(_4116_),
    .B(_4118_),
    .Y(_4120_)
);

FILL FILL_0__10215_ (
);

AOI21X1 _10500_ (
    .A(_3745_),
    .B(_3747_),
    .C(_3773_),
    .Y(_3774_)
);

DFFPOSX1 _13392_ (
    .D(_6375_[14]),
    .CLK(clk_bF$buf24),
    .Q(\u_fir_pe7.mul [14])
);

NAND2X1 _7707_ (
    .A(_1188_),
    .B(_1191_),
    .Y(_1224_)
);

FILL FILL_1__6664_ (
);

FILL FILL_2__13014_ (
);

FILL FILL254250x172950 (
);

FILL FILL_1__12847_ (
);

FILL FILL_1__12427_ (
);

FILL FILL_1__12007_ (
);

FILL FILL_3__7951_ (
);

FILL FILL_0__9434_ (
);

FILL FILL_0__9014_ (
);

NAND3X1 _11705_ (
    .A(_4814_),
    .B(_4826_),
    .C(_4822_),
    .Y(_4827_)
);

FILL FILL_3__7111_ (
);

FILL FILL_1__7869_ (
);

FILL FILL_3__10781_ (
);

FILL FILL_1__7449_ (
);

FILL FILL_1__7029_ (
);

FILL FILL_1__8810_ (
);

FILL FILL_3__8736_ (
);

NAND2X1 _7880_ (
    .A(_1364_),
    .B(_1392_),
    .Y(_1393_)
);

NAND3X1 _7460_ (
    .A(_933_),
    .B(_974_),
    .C(_979_),
    .Y(_980_)
);

NAND2X1 _7040_ (
    .A(_630_),
    .B(_629_),
    .Y(_796_[15])
);

AOI21X1 _10097_ (
    .A(_3289_),
    .B(_3293_),
    .C(_3257_),
    .Y(_3377_)
);

FILL FILL_2__6733_ (
);

FILL FILL_3__11566_ (
);

FILL FILL_1__12180_ (
);

FILL FILL_2__10979_ (
);

FILL FILL_2__10559_ (
);

FILL FILL_2__10139_ (
);

FILL FILL_0__11173_ (
);

FILL FILL_2__11920_ (
);

FILL FILL_2__11500_ (
);

FILL FILL_0__6979_ (
);

FILL FILL_0__6559_ (
);

AOI21X1 _8665_ (
    .A(_2049_),
    .B(_2052_),
    .C(_2100_),
    .Y(_2101_)
);

NAND3X1 _8245_ (
    .A(gnd),
    .B(\X[2] [3]),
    .C(_1677_),
    .Y(_1686_)
);

FILL FILL_1__10913_ (
);

FILL FILL_0__7920_ (
);

FILL FILL_2__7938_ (
);

FILL FILL_2__7518_ (
);

FILL FILL_0__7500_ (
);

FILL FILL_0__12798_ (
);

NAND3X1 _12663_ (
    .A(_5702_),
    .B(_5703_),
    .C(_5701_),
    .Y(_5704_)
);

FILL FILL_0__12378_ (
);

OAI21X1 _12243_ (
    .A(_5355_),
    .B(_5356_),
    .C(_5308_),
    .Y(_5357_)
);

FILL FILL_2__12705_ (
);

FILL FILL_0__8705_ (
);

FILL FILL_3__9694_ (
);

FILL FILL_3__9274_ (
);

NAND2X1 _13028_ (
    .A(_6061_),
    .B(_6055_),
    .Y(_6064_)
);

FILL FILL_2__7691_ (
);

FILL FILL_2__7271_ (
);

FILL FILL_2__11097_ (
);

AOI21X1 _6731_ (
    .A(_328_),
    .B(_326_),
    .C(_324_),
    .Y(_329_)
);

FILL FILL_0__7097_ (
);

FILL FILL_3__10837_ (
);

FILL FILL_1__11871_ (
);

FILL FILL_3__10417_ (
);

FILL FILL_1__11451_ (
);

FILL FILL_1__11031_ (
);

FILL FILL_2__8896_ (
);

FILL FILL_2__8476_ (
);

FILL FILL_0__10864_ (
);

FILL FILL_0__10444_ (
);

FILL FILL_2__8056_ (
);

FILL FILL_0__10024_ (
);

NAND2X1 _7936_ (
    .A(_1440_),
    .B(_1443_),
    .Y(_1587_[2])
);

NAND2X1 _7516_ (
    .A(_1029_),
    .B(_1034_),
    .Y(_1035_)
);

FILL FILL_1__6893_ (
);

FILL FILL_1__6473_ (
);

FILL FILL_2__13243_ (
);

FILL FILL_3__6399_ (
);

FILL FILL_1__12656_ (
);

FILL FILL_1__12236_ (
);

FILL FILL_0__9663_ (
);

FILL FILL_0__9243_ (
);

NAND3X1 _11934_ (
    .A(_5006_),
    .B(_5048_),
    .C(_5049_),
    .Y(_5053_)
);

FILL FILL_0__11649_ (
);

FILL FILL_3__7340_ (
);

NOR2X1 _11514_ (
    .A(\u_fir_pe5.rYin [9]),
    .B(\u_fir_pe5.mul [9]),
    .Y(_4698_)
);

FILL FILL_0__11229_ (
);

FILL FILL_1__7678_ (
);

FILL FILL_1__7258_ (
);

FILL FILL_3__10170_ (
);

AOI21X1 _12719_ (
    .A(_5753_),
    .B(_5754_),
    .C(_5752_),
    .Y(_5759_)
);

FILL FILL_1_BUFX2_insert70 (
);

FILL FILL_1_BUFX2_insert71 (
);

FILL FILL_1_BUFX2_insert72 (
);

FILL FILL_1_BUFX2_insert73 (
);

FILL FILL_1_BUFX2_insert74 (
);

FILL FILL_1_BUFX2_insert75 (
);

FILL FILL_1_BUFX2_insert76 (
);

FILL FILL_1_BUFX2_insert77 (
);

FILL FILL_1_BUFX2_insert78 (
);

FILL FILL_1_BUFX2_insert79 (
);

FILL FILL_2__6962_ (
);

FILL FILL_3__11795_ (
);

FILL FILL_2__6542_ (
);

FILL FILL_2__10788_ (
);

FILL FILL_2__10368_ (
);

FILL FILL_1__9824_ (
);

FILL FILL_1__9404_ (
);

FILL FILL_0_CLKBUF1_insert50 (
);

FILL FILL_0_CLKBUF1_insert51 (
);

FILL FILL_0_CLKBUF1_insert52 (
);

FILL FILL_0_CLKBUF1_insert53 (
);

FILL FILL_0_CLKBUF1_insert54 (
);

FILL FILL_0__6788_ (
);

FILL FILL_0_CLKBUF1_insert55 (
);

INVX1 _8894_ (
    .A(\u_fir_pe2.rYin [10]),
    .Y(_2318_)
);

NAND2X1 _8474_ (
    .A(\X[2] [3]),
    .B(vdd),
    .Y(_1912_)
);

FILL FILL_0_CLKBUF1_insert56 (
);

FILL FILL_0_CLKBUF1_insert57 (
);

INVX1 _8054_ (
    .A(\u_fir_pe1.mul [14]),
    .Y(_1558_)
);

FILL FILL_0_CLKBUF1_insert58 (
);

FILL FILL_0_CLKBUF1_insert59 (
);

FILL FILL_1__10302_ (
);

FILL FILL_2__7747_ (
);

FILL FILL_2__7327_ (
);

FILL FILL_1__13194_ (
);

NAND3X1 _12892_ (
    .A(_5928_),
    .B(_5929_),
    .C(_5927_),
    .Y(_5930_)
);

FILL FILL_0__12187_ (
);

DFFPOSX1 _12472_ (
    .D(_5572_[11]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[11])
);

NOR2X1 _12052_ (
    .A(_5100_),
    .B(_5103_),
    .Y(_5169_)
);

FILL FILL_2__12934_ (
);

NAND2X1 _9679_ (
    .A(_3022_),
    .B(_3027_),
    .Y(_3028_)
);

AND2X2 _9259_ (
    .A(\X[3] [3]),
    .B(gnd),
    .Y(_2618_)
);

FILL FILL_1__11927_ (
);

FILL FILL_1__11507_ (
);

FILL FILL_0__8934_ (
);

FILL FILL_0__8514_ (
);

FILL FILL_3__6611_ (
);

NAND3X1 _13257_ (
    .A(_6280_),
    .B(_6277_),
    .C(_6240_),
    .Y(_6281_)
);

FILL FILL_1__6949_ (
);

FILL FILL_1__6529_ (
);

FILL FILL_2__7080_ (
);

FILL FILL_0__9719_ (
);

FILL FILL_3__7816_ (
);

OAI21X1 _6960_ (
    .A(_504_),
    .B(_507_),
    .C(_552_),
    .Y(_555_)
);

INVX1 _6540_ (
    .A(_139_),
    .Y(_140_)
);

FILL FILL_3__10646_ (
);

FILL FILL_1__11680_ (
);

FILL FILL_1__11260_ (
);

FILL FILL_2__8285_ (
);

FILL FILL_0__10673_ (
);

FILL FILL_0__10253_ (
);

OAI22X1 _7745_ (
    .A(_1214_),
    .B(_1102_),
    .C(_822_),
    .D(_1213_),
    .Y(_1261_)
);

NAND2X1 _7325_ (
    .A(_829_),
    .B(_844_),
    .Y(_847_)
);

FILL FILL_2__13052_ (
);

FILL FILL_1__12885_ (
);

FILL FILL_1__12045_ (
);

FILL FILL_0__9892_ (
);

FILL FILL_0__9472_ (
);

FILL FILL_0__11878_ (
);

FILL FILL_0__9052_ (
);

AND2X2 _11743_ (
    .A(_4859_),
    .B(_4863_),
    .Y(_4864_)
);

FILL FILL_0__11458_ (
);

FILL FILL_0__11038_ (
);

AND2X2 _11323_ (
    .A(_4508_),
    .B(_4504_),
    .Y(_4518_)
);

FILL FILL_1__7487_ (
);

FILL FILL_1__7067_ (
);

AOI21X1 _12948_ (
    .A(_5910_),
    .B(_5984_),
    .C(_5983_),
    .Y(_5985_)
);

FILL FILL_3__8354_ (
);

NAND2X1 _12528_ (
    .A(_6359_),
    .B(_6339_),
    .Y(_6360_)
);

INVX1 _12108_ (
    .A(_5146_),
    .Y(_5225_)
);

FILL FILL_2__6771_ (
);

FILL FILL_3__11184_ (
);

FILL FILL_2__10597_ (
);

FILL FILL_2__10177_ (
);

FILL FILL_1__9633_ (
);

FILL FILL_1__9213_ (
);

FILL FILL_3__9979_ (
);

FILL FILL_3__9139_ (
);

FILL FILL_0__6597_ (
);

OAI21X1 _8283_ (
    .A(_1722_),
    .B(_1723_),
    .C(_1721_),
    .Y(_1724_)
);

FILL FILL_1__10951_ (
);

FILL FILL_1__10531_ (
);

FILL FILL_1__10111_ (
);

FILL FILL_2__7976_ (
);

FILL FILL_2__7556_ (
);

FILL FILL_3__12389_ (
);

FILL FILL_2__7136_ (
);

AND2X2 _12281_ (
    .A(_5390_),
    .B(_5387_),
    .Y(_5394_)
);

FILL FILL_2__12743_ (
);

FILL FILL_2__12323_ (
);

NAND2X1 _9488_ (
    .A(_2833_),
    .B(_2840_),
    .Y(_2844_)
);

INVX1 _9068_ (
    .A(_2429_),
    .Y(_2430_)
);

FILL FILL_1__11736_ (
);

FILL FILL_1__11316_ (
);

FILL FILL_0__8743_ (
);

FILL FILL_3__6840_ (
);

FILL FILL_0__8323_ (
);

FILL FILL_0__10309_ (
);

FILL FILL254550x118950 (
);

OAI21X1 _13066_ (
    .A(_5653_),
    .B(_5884_),
    .C(_6058_),
    .Y(_6101_)
);

FILL FILL_2__9702_ (
);

FILL FILL_1__6758_ (
);

FILL FILL_2__13108_ (
);

FILL FILL_0__9948_ (
);

FILL FILL_0__9528_ (
);

FILL FILL_3__7625_ (
);

FILL FILL_0__9108_ (
);

FILL FILL_3__10035_ (
);

FILL FILL_0__10482_ (
);

FILL FILL_0__10062_ (
);

FILL FILL_1__8904_ (
);

OAI21X1 _7974_ (
    .A(_1470_),
    .B(_1471_),
    .C(_1475_),
    .Y(_1477_)
);

AOI21X1 _7554_ (
    .A(_981_),
    .B(_979_),
    .C(_1072_),
    .Y(_1073_)
);

NAND2X1 _7134_ (
    .A(_717_),
    .B(_716_),
    .Y(_790_[9])
);

FILL FILL_2__13281_ (
);

FILL FILL_2__6827_ (
);

FILL FILL_2__6407_ (
);

FILL FILL_1__12694_ (
);

FILL FILL_1__12274_ (
);

FILL FILL_0__9281_ (
);

FILL FILL_2__9299_ (
);

NOR2X1 _11972_ (
    .A(_5088_),
    .B(_5089_),
    .Y(_5090_)
);

FILL FILL_0__11687_ (
);

INVX1 _11552_ (
    .A(\u_fir_pe5.rYin [13]),
    .Y(_4736_)
);

FILL FILL_0__11267_ (
);

AOI21X1 _11132_ (
    .A(_4329_),
    .B(_4328_),
    .C(_4327_),
    .Y(_4330_)
);

NAND2X1 _8759_ (
    .A(_2191_),
    .B(_2190_),
    .Y(_2192_)
);

OAI21X1 _8339_ (
    .A(_1774_),
    .B(_1775_),
    .C(_1732_),
    .Y(_1779_)
);

FILL FILL_1__7296_ (
);

INVX1 _9700_ (
    .A(\u_fir_pe3.rYin [4]),
    .Y(_3046_)
);

FILL FILL_1__13059_ (
);

FILL FILL_3__8583_ (
);

NAND3X1 _12757_ (
    .A(_5722_),
    .B(_5791_),
    .C(_5726_),
    .Y(_5796_)
);

OAI21X1 _12337_ (
    .A(_5433_),
    .B(_5429_),
    .C(_5442_),
    .Y(_5443_)
);

FILL FILL_0__13413_ (
);

FILL FILL_2__6580_ (
);

FILL FILL_1__9442_ (
);

FILL FILL_1__9022_ (
);

FILL FILL_3__9788_ (
);

FILL FILL_3__9368_ (
);

DFFPOSX1 _8092_ (
    .D(\X[1] [0]),
    .CLK(clk_bF$buf10),
    .Q(\X[2] [0])
);

FILL FILL_1__10340_ (
);

FILL FILL_2__7785_ (
);

FILL FILL_2__7365_ (
);

NAND3X1 _12090_ (
    .A(_5125_),
    .B(_5131_),
    .C(_5206_),
    .Y(_5207_)
);

NAND3X1 _6825_ (
    .A(_419_),
    .B(_420_),
    .C(_421_),
    .Y(_422_)
);

OAI21X1 _6405_ (
    .A(_4_),
    .B(_7_),
    .C(_0_),
    .Y(_8_)
);

FILL FILL_2__12972_ (
);

FILL FILL_2__12552_ (
);

FILL FILL_2__12132_ (
);

AOI21X1 _9297_ (
    .A(_2543_),
    .B(_2562_),
    .C(_2655_),
    .Y(_2656_)
);

FILL FILL_1__11965_ (
);

FILL FILL_1__11545_ (
);

FILL FILL_1__11125_ (
);

FILL FILL_0__8552_ (
);

FILL FILL_0__10958_ (
);

FILL FILL_0__8132_ (
);

FILL FILL_0__10538_ (
);

NAND3X1 _10823_ (
    .A(_4019_),
    .B(_4024_),
    .C(_4022_),
    .Y(_4025_)
);

NAND3X1 _10403_ (
    .A(_3676_),
    .B(_3678_),
    .C(_3677_),
    .Y(_3679_)
);

FILL FILL_0__10118_ (
);

NAND2X1 _13295_ (
    .A(_6314_),
    .B(_6307_),
    .Y(_6318_)
);

FILL FILL_2__9931_ (
);

FILL FILL_2__9511_ (
);

FILL FILL_1__6987_ (
);

FILL FILL_1__6567_ (
);

FILL FILL_2__13337_ (
);

FILL FILL_0__9757_ (
);

FILL FILL_0__9337_ (
);

DFFPOSX1 _11608_ (
    .D(\Y[5] [0]),
    .CLK(clk_bF$buf40),
    .Q(\u_fir_pe5.rYin [0])
);

FILL FILL_3__10264_ (
);

FILL FILL_0__10291_ (
);

FILL FILL_1__8713_ (
);

FILL FILL_3__8219_ (
);

AOI21X1 _7783_ (
    .A(_1292_),
    .B(_1298_),
    .C(_1256_),
    .Y(_1299_)
);

AND2X2 _7363_ (
    .A(vdd),
    .B(\X[1] [3]),
    .Y(_884_)
);

FILL FILL_2__13090_ (
);

FILL FILL_3__11889_ (
);

FILL FILL_2__6636_ (
);

FILL FILL_3__11049_ (
);

FILL FILL_1__12083_ (
);

FILL FILL_0__9090_ (
);

NAND3X1 _11781_ (
    .A(_4898_),
    .B(_4901_),
    .C(_4850_),
    .Y(_4902_)
);

FILL FILL_0__11496_ (
);

FILL FILL_0__11076_ (
);

OR2X2 _11361_ (
    .A(_4554_),
    .B(_4550_),
    .Y(_4555_)
);

FILL FILL_1__9918_ (
);

FILL FILL_3__12410_ (
);

FILL FILL_2__11823_ (
);

FILL FILL_2__11403_ (
);

DFFPOSX1 _8988_ (
    .D(\Y[2] [11]),
    .CLK(clk_bF$buf7),
    .Q(\u_fir_pe2.rYin [11])
);

NAND2X1 _8568_ (
    .A(_1995_),
    .B(_2004_),
    .Y(_2005_)
);

INVX1 _8148_ (
    .A(_2379_),
    .Y(_2380_)
);

FILL FILL_1__10816_ (
);

FILL FILL_0__7823_ (
);

FILL FILL_0__7403_ (
);

FILL FILL_1__13288_ (
);

AOI21X1 _12986_ (
    .A(_5879_),
    .B(_5944_),
    .C(_6022_),
    .Y(_6023_)
);

INVX1 _12566_ (
    .A(_5607_),
    .Y(_5608_)
);

OAI21X1 _12146_ (
    .A(_4856_),
    .B(_5101_),
    .C(_5255_),
    .Y(_5262_)
);

FILL FILL_2__12608_ (
);

FILL FILL_0__13222_ (
);

FILL FILL_0__8608_ (
);

FILL FILL_3__6705_ (
);

FILL FILL_1__9671_ (
);

FILL FILL_1__9251_ (
);

FILL FILL_3__9597_ (
);

FILL FILL_2__7594_ (
);

FILL FILL_2__7174_ (
);

INVX1 _6634_ (
    .A(gnd),
    .Y(_233_)
);

FILL FILL_2__12781_ (
);

FILL FILL_2__12361_ (
);

FILL FILL_1__11774_ (
);

FILL FILL_1__11354_ (
);

FILL FILL_0__8781_ (
);

FILL FILL_2__8799_ (
);

FILL FILL_2__8379_ (
);

FILL FILL_0__8361_ (
);

FILL FILL_0__10767_ (
);

NAND2X1 _10632_ (
    .A(_3892_),
    .B(_3895_),
    .Y(_3978_[8])
);

FILL FILL_0__10347_ (
);

AOI21X1 _10212_ (
    .A(_3454_),
    .B(_3455_),
    .C(_3412_),
    .Y(_3490_)
);

FILL FILL_2__9740_ (
);

FILL FILL_2__9320_ (
);

NOR3X1 _7839_ (
    .A(_1299_),
    .B(_1301_),
    .C(_1349_),
    .Y(_1353_)
);

AND2X2 _7419_ (
    .A(gnd),
    .B(\X[1] [6]),
    .Y(_939_)
);

FILL FILL_1__6796_ (
);

FILL FILL_2__13146_ (
);

FILL FILL_1__12979_ (
);

FILL FILL_1__12559_ (
);

FILL FILL_1__12139_ (
);

FILL FILL_0__9986_ (
);

FILL FILL_0__9566_ (
);

FILL FILL_3__7663_ (
);

FILL FILL_0__9146_ (
);

NAND3X1 _11837_ (
    .A(_4944_),
    .B(_4948_),
    .C(_4950_),
    .Y(_4957_)
);

NOR3X1 _11417_ (
    .A(_4608_),
    .B(_4576_),
    .C(_4594_),
    .Y(_4609_)
);

FILL FILL_0__12913_ (
);

FILL FILL_3__10493_ (
);

FILL FILL254250x104550 (
);

FILL FILL_1__8942_ (
);

FILL FILL_1__8522_ (
);

FILL FILL_3__8448_ (
);

NAND2X1 _7592_ (
    .A(_1103_),
    .B(_1104_),
    .Y(_1110_)
);

NAND2X1 _7172_ (
    .A(_755_),
    .B(_749_),
    .Y(_756_)
);

FILL FILL_2__6865_ (
);

FILL FILL253950x43350 (
);

FILL FILL_2__6445_ (
);

FILL FILL_3__11278_ (
);

DFFPOSX1 _11590_ (
    .D(_4775_[6]),
    .CLK(clk_bF$buf48),
    .Q(\Y[6] [6])
);

OAI21X1 _11170_ (
    .A(_4286_),
    .B(_4366_),
    .C(_4349_),
    .Y(_4367_)
);

FILL FILL_1__9727_ (
);

FILL FILL_1__9307_ (
);

FILL FILL_2__11212_ (
);

INVX1 _8797_ (
    .A(\u_fir_pe2.rYin [1]),
    .Y(_2226_)
);

NAND2X1 _8377_ (
    .A(_1812_),
    .B(_1815_),
    .Y(_1816_)
);

FILL FILL_1__10625_ (
);

FILL FILL_1__10205_ (
);

FILL FILL_0__7632_ (
);

FILL FILL_1__13097_ (
);

NOR2X1 _12795_ (
    .A(_5820_),
    .B(_5833_),
    .Y(_5834_)
);

NAND2X1 _12375_ (
    .A(_5457_),
    .B(_5469_),
    .Y(_5478_)
);

FILL FILL_3__13004_ (
);

FILL FILL_2__12837_ (
);

FILL FILL_2__12417_ (
);

FILL FILL_0__13031_ (
);

FILL FILL_0__8837_ (
);

FILL FILL_3__6934_ (
);

FILL FILL_0__8417_ (
);

FILL FILL_1__9480_ (
);

FILL FILL_1__9060_ (
);

FILL FILL_3__7719_ (
);

OAI21X1 _6863_ (
    .A(_438_),
    .B(_440_),
    .C(_431_),
    .Y(_459_)
);

NAND3X1 _6443_ (
    .A(_32_),
    .B(_44_),
    .C(_40_),
    .Y(_45_)
);

FILL FILL_2__12590_ (
);

FILL FILL_2__12170_ (
);

FILL FILL_1__11583_ (
);

FILL FILL_3__10129_ (
);

FILL FILL_1__11163_ (
);

FILL FILL_0__8590_ (
);

FILL FILL_0__10996_ (
);

FILL FILL_2__8188_ (
);

FILL FILL_0__8170_ (
);

FILL FILL_0__10576_ (
);

NAND3X1 _10861_ (
    .A(_4061_),
    .B(_4056_),
    .C(_4058_),
    .Y(_4062_)
);

OAI21X1 _10441_ (
    .A(_3661_),
    .B(_3714_),
    .C(_3715_),
    .Y(_3716_)
);

FILL FILL_0__10156_ (
);

NAND3X1 _10021_ (
    .A(_3289_),
    .B(_3293_),
    .C(_3295_),
    .Y(_3302_)
);

FILL FILL_3__11910_ (
);

FILL FILL_2__10903_ (
);

OAI21X1 _7648_ (
    .A(_932_),
    .B(_1165_),
    .C(_1079_),
    .Y(_1166_)
);

DFFPOSX1 _7228_ (
    .D(Yin[5]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [5])
);

FILL FILL_0__6903_ (
);

FILL FILL_1__12788_ (
);

FILL FILL_1__12368_ (
);

FILL FILL_0__9795_ (
);

FILL FILL_3__7892_ (
);

FILL FILL_0__9375_ (
);

AOI22X1 _11646_ (
    .A(\X[7] [0]),
    .B(vdd),
    .C(\X[7] [1]),
    .D(gnd),
    .Y(_5532_)
);

FILL FILL_3__7052_ (
);

INVX1 _11226_ (
    .A(_4368_),
    .Y(_4423_)
);

FILL FILL_0__12722_ (
);

FILL FILL_0__12302_ (
);

FILL FILL_1__8751_ (
);

FILL FILL_1__8331_ (
);

FILL FILL_3__8677_ (
);

FILL FILL_2__6674_ (
);

FILL FILL_1__9956_ (
);

FILL FILL_1__9536_ (
);

FILL FILL_1__9116_ (
);

FILL FILL_2__11861_ (
);

FILL FILL_2__11441_ (
);

FILL FILL_2__11021_ (
);

INVX1 _8186_ (
    .A(_1627_),
    .Y(_1628_)
);

FILL FILL_1__10854_ (
);

FILL FILL_1__10434_ (
);

FILL FILL_1__10014_ (
);

FILL FILL_0__7861_ (
);

FILL FILL_2__7879_ (
);

FILL FILL_2__7459_ (
);

FILL FILL_0__7441_ (
);

FILL FILL_0__7021_ (
);

FILL FILL_2__7039_ (
);

NOR3X1 _12184_ (
    .A(_5087_),
    .B(_5255_),
    .C(_5198_),
    .Y(_5299_)
);

FILL FILL_2__8820_ (
);

FILL FILL_2__8400_ (
);

FILL FILL_3__13233_ (
);

AOI21X1 _6919_ (
    .A(_460_),
    .B(_494_),
    .C(_513_),
    .Y(_514_)
);

FILL FILL_2__12646_ (
);

FILL FILL_2__12226_ (
);

FILL FILL_0__13260_ (
);

FILL FILL_1__11219_ (
);

FILL FILL_0__8646_ (
);

FILL FILL_0__8226_ (
);

NAND2X1 _10917_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf1 ),
    .Y(_4117_)
);

DFFPOSX1 _13389_ (
    .D(_6375_[11]),
    .CLK(clk_bF$buf40),
    .Q(\u_fir_pe7.mul [11])
);

FILL FILL_2__9605_ (
);

FILL FILL_1__7602_ (
);

FILL FILL_3__7948_ (
);

NAND3X1 _6672_ (
    .A(_224_),
    .B(_266_),
    .C(_267_),
    .Y(_271_)
);

FILL FILL_3__10778_ (
);

FILL FILL_3__10358_ (
);

FILL FILL_1__11392_ (
);

FILL FILL_0__10385_ (
);

NOR2X1 _10670_ (
    .A(_3933_),
    .B(_3932_),
    .Y(_3934_)
);

NAND3X1 _10250_ (
    .A(_3526_),
    .B(_3527_),
    .C(_3525_),
    .Y(_3528_)
);

FILL FILL_1__8807_ (
);

OAI21X1 _7877_ (
    .A(_1102_),
    .B(_1389_),
    .C(_1368_),
    .Y(_1390_)
);

AOI21X1 _7457_ (
    .A(_971_),
    .B(_972_),
    .C(_970_),
    .Y(_977_)
);

NAND2X1 _7037_ (
    .A(_628_),
    .B(_622_),
    .Y(_796_[14])
);

FILL FILL_2__13184_ (
);

FILL FILL_0__6712_ (
);

FILL FILL_1__12597_ (
);

FILL FILL_1__12177_ (
);

FILL FILL_0__9184_ (
);

NAND2X1 _11875_ (
    .A(\X[7] [1]),
    .B(gnd),
    .Y(_4994_)
);

FILL FILL_3__7281_ (
);

INVX1 _11455_ (
    .A(\u_fir_pe5.mul [4]),
    .Y(_4641_)
);

INVX1 _11035_ (
    .A(_4233_),
    .Y(_4234_)
);

FILL FILL_2__11917_ (
);

FILL FILL_0__12951_ (
);

FILL FILL_0__12531_ (
);

FILL FILL_0__12111_ (
);

FILL FILL_0__7917_ (
);

NOR2X1 _9603_ (
    .A(_2864_),
    .B(_2917_),
    .Y(_2957_)
);

FILL FILL_1__8560_ (
);

FILL FILL_1__8140_ (
);

FILL FILL_3__8066_ (
);

FILL FILL_0__13316_ (
);

FILL FILL_2__6483_ (
);

FILL FILL_1__9765_ (
);

FILL FILL_1__9345_ (
);

FILL FILL_2__11670_ (
);

FILL FILL_2__11250_ (
);

FILL FILL_1__10663_ (
);

FILL FILL_1__10243_ (
);

FILL FILL_0__7670_ (
);

FILL FILL_2__7688_ (
);

FILL FILL_2__7268_ (
);

NAND3X1 _6728_ (
    .A(vdd),
    .B(Xin[6]),
    .C(_325_),
    .Y(_326_)
);

FILL FILL_2__12875_ (
);

FILL FILL_2__12455_ (
);

FILL FILL_2__12035_ (
);

FILL FILL_1__11868_ (
);

FILL FILL_1__11448_ (
);

FILL FILL_1__11028_ (
);

FILL FILL_0__8875_ (
);

FILL FILL_0__8455_ (
);

FILL FILL_3__6552_ (
);

FILL FILL_0__8035_ (
);

DFFPOSX1 _10726_ (
    .D(\X[4] [3]),
    .CLK(clk_bF$buf25),
    .Q(\X[5] [3])
);

AND2X2 _10306_ (
    .A(_3582_),
    .B(_3579_),
    .Y(_3583_)
);

NAND2X1 _13198_ (
    .A(_6222_),
    .B(_6225_),
    .Y(_6369_[2])
);

FILL FILL_2__9414_ (
);

FILL FILL_0__11802_ (
);

FILL FILL_1__7831_ (
);

FILL FILL_1__7411_ (
);

FILL FILL_3__7757_ (
);

FILL FILL_3__7337_ (
);

AND2X2 _6481_ (
    .A(_77_),
    .B(_81_),
    .Y(_82_)
);

FILL FILL_3__10587_ (
);

FILL FILL_0__10194_ (
);

FILL FILL_1__8616_ (
);

FILL FILL_2__10941_ (
);

FILL FILL_2__10521_ (
);

FILL FILL_2__10101_ (
);

AOI21X1 _7686_ (
    .A(_1128_),
    .B(_1202_),
    .C(_1201_),
    .Y(_1203_)
);

NAND2X1 _7266_ (
    .A(_1577_),
    .B(_1557_),
    .Y(_1578_)
);

FILL FILL_0__6941_ (
);

FILL FILL_2__6959_ (
);

FILL FILL_2__6539_ (
);

FILL FILL_0__6521_ (
);

NAND2X1 _11684_ (
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4806_)
);

FILL FILL_0__11399_ (
);

AND2X2 _11264_ (
    .A(_4458_),
    .B(_4401_),
    .Y(_4460_)
);

FILL FILL_2__7900_ (
);

FILL FILL_3__12733_ (
);

FILL FILL_2__11726_ (
);

FILL FILL_0__12760_ (
);

FILL FILL_2__11306_ (
);

FILL FILL_0__12340_ (
);

FILL FILL_0__7726_ (
);

DFFPOSX1 _9832_ (
    .D(_3181_[2]),
    .CLK(clk_bF$buf55),
    .Q(\Y[4] [2])
);

FILL FILL_0__7306_ (
);

NAND2X1 _9412_ (
    .A(_2765_),
    .B(_2769_),
    .Y(_3187_[8])
);

AOI21X1 _12889_ (
    .A(_5838_),
    .B(_5840_),
    .C(_5926_),
    .Y(_5927_)
);

FILL FILL_3__8295_ (
);

DFFPOSX1 _12469_ (
    .D(_5572_[8]),
    .CLK(clk_bF$buf23),
    .Q(_6377_[8])
);

AOI21X1 _12049_ (
    .A(_5131_),
    .B(_5132_),
    .C(_5099_),
    .Y(_5166_)
);

FILL FILL_0__13125_ (
);

BUFX2 _13410_ (
    .A(_6377_[2]),
    .Y(Yout[2])
);

FILL FILL_1__9994_ (
);

FILL FILL_1__9574_ (
);

FILL FILL_1__9154_ (
);

FILL FILL_1__10892_ (
);

FILL FILL_1__10472_ (
);

FILL FILL_1__10052_ (
);

FILL FILL_2__7497_ (
);

FILL FILL_2__7077_ (
);

NAND2X1 _6957_ (
    .A(_548_),
    .B(_551_),
    .Y(_552_)
);

AOI21X1 _6537_ (
    .A(_91_),
    .B(_95_),
    .C(_84_),
    .Y(_137_)
);

FILL FILL_2__12684_ (
);

FILL FILL_2__12264_ (
);

FILL FILL_1__11677_ (
);

FILL FILL_1__11257_ (
);

FILL FILL_0__8684_ (
);

FILL FILL_3__6781_ (
);

FILL FILL_0__8264_ (
);

AOI22X1 _10955_ (
    .A(gnd),
    .B(\X[5]_5_bF$buf1 ),
    .C(_4144_),
    .D(_4146_),
    .Y(_4155_)
);

OR2X2 _10535_ (
    .A(_3805_),
    .B(_3806_),
    .Y(_3807_)
);

NOR2X1 _10115_ (
    .A(_3392_),
    .B(_3394_),
    .Y(_3984_[6])
);

FILL FILL_2__9643_ (
);

FILL FILL_2__9223_ (
);

FILL FILL_1__6699_ (
);

FILL FILL_2__13049_ (
);

FILL FILL_1__7640_ (
);

FILL FILL_0__9889_ (
);

FILL FILL_3__7986_ (
);

FILL FILL_0__9469_ (
);

FILL FILL_3__7566_ (
);

FILL FILL_0__9049_ (
);

FILL FILL_3__7146_ (
);

FILL FILL_1__13403_ (
);

FILL FILL_0__12816_ (
);

FILL FILL_1__8845_ (
);

FILL FILL_1__8425_ (
);

FILL FILL_1__8005_ (
);

FILL FILL_2__10330_ (
);

NAND3X1 _7495_ (
    .A(_940_),
    .B(_1009_),
    .C(_944_),
    .Y(_1014_)
);

OAI21X1 _7075_ (
    .A(_651_),
    .B(_647_),
    .C(_660_),
    .Y(_661_)
);

FILL FILL_0__6750_ (
);

FILL FILL_2__6768_ (
);

INVX1 _11493_ (
    .A(\u_fir_pe5.mul [8]),
    .Y(_4676_)
);

NAND3X1 _11073_ (
    .A(_4120_),
    .B(_4259_),
    .C(_4264_),
    .Y(_4272_)
);

FILL FILL_3__12962_ (
);

FILL FILL_3__12122_ (
);

FILL FILL_2__11955_ (
);

FILL FILL_2__11535_ (
);

FILL FILL_2__11115_ (
);

FILL FILL_1__10948_ (
);

FILL FILL_1__10528_ (
);

FILL FILL_1__10108_ (
);

FILL FILL_0__7955_ (
);

FILL FILL_0__7535_ (
);

OR2X2 _9641_ (
    .A(_2992_),
    .B(_2985_),
    .Y(_2994_)
);

FILL FILL_0__7115_ (
);

OAI21X1 _9221_ (
    .A(_2503_),
    .B(_2580_),
    .C(_2497_),
    .Y(_2581_)
);

NAND2X1 _12698_ (
    .A(_5666_),
    .B(_5737_),
    .Y(_5738_)
);

NAND2X1 _12278_ (
    .A(_5387_),
    .B(_5390_),
    .Y(_5391_)
);

FILL FILL_2__8914_ (
);

FILL FILL_3__13327_ (
);

FILL FILL_1__6911_ (
);

FILL FILL_3__6417_ (
);

FILL FILL_1__9383_ (
);

FILL FILL_1__10281_ (
);

FILL FILL_3__13080_ (
);

NAND3X1 _6766_ (
    .A(_303_),
    .B(_360_),
    .C(_361_),
    .Y(_364_)
);

FILL FILL_2__12073_ (
);

FILL FILL_1__11486_ (
);

FILL FILL_1__11066_ (
);

FILL FILL_0__8493_ (
);

FILL FILL_0__10899_ (
);

FILL FILL_0__10479_ (
);

AND2X2 _10764_ (
    .A(\X[5] [1]),
    .B(vdd),
    .Y(_4685_)
);

FILL FILL_0__8073_ (
);

AOI21X1 _10344_ (
    .A(_3541_),
    .B(_3543_),
    .C(_3620_),
    .Y(_3621_)
);

FILL FILL_0__10059_ (
);

FILL FILL_2__10806_ (
);

FILL FILL_2__9452_ (
);

FILL FILL_0__11840_ (
);

FILL FILL_2__9032_ (
);

FILL FILL_0__11420_ (
);

FILL FILL_0__11000_ (
);

FILL FILL_2__13278_ (
);

FILL FILL_0__6806_ (
);

INVX1 _8912_ (
    .A(\u_fir_pe2.rYin [12]),
    .Y(_2336_)
);

FILL FILL_0__9698_ (
);

FILL FILL_0__9278_ (
);

INVX2 _11969_ (
    .A(gnd),
    .Y(_5087_)
);

FILL FILL_3__7375_ (
);

OR2X2 _11549_ (
    .A(_4726_),
    .B(_4731_),
    .Y(_4733_)
);

INVX1 _11129_ (
    .A(_4307_),
    .Y(_4327_)
);

FILL FILL_1__13212_ (
);

OAI21X1 _12910_ (
    .A(_5714_),
    .B(_5947_),
    .C(_5861_),
    .Y(_5948_)
);

FILL FILL_0__12625_ (
);

FILL FILL_0__12205_ (
);

FILL FILL_1__8654_ (
);

FILL FILL_1__8234_ (
);

FILL FILL_3__9521_ (
);

FILL FILL_2__6997_ (
);

FILL FILL_2__6577_ (
);

FILL FILL_1__9439_ (
);

FILL FILL_1__9019_ (
);

FILL FILL_3__12351_ (
);

FILL FILL_2__11764_ (
);

FILL FILL_2__11344_ (
);

DFFPOSX1 _8089_ (
    .D(_1587_[13]),
    .CLK(clk_bF$buf3),
    .Q(\Y[2] [13])
);

FILL FILL_1__10337_ (
);

FILL FILL_0__7764_ (
);

DFFPOSX1 _9870_ (
    .D(_3182_[0]),
    .CLK(clk_bF$buf28),
    .Q(\u_fir_pe3.mul [0])
);

FILL FILL_0__7344_ (
);

NAND2X1 _9450_ (
    .A(\X[3]_5_bF$buf3 ),
    .B(vdd),
    .Y(_2807_)
);

NAND2X1 _9030_ (
    .A(gnd),
    .B(\X[3] [0]),
    .Y(_2393_)
);

NAND3X1 _12087_ (
    .A(_5201_),
    .B(_5202_),
    .C(_5203_),
    .Y(_5204_)
);

FILL FILL_2__8723_ (
);

FILL FILL_2__8303_ (
);

FILL FILL_2__12969_ (
);

FILL FILL_2__12549_ (
);

FILL FILL_2__12129_ (
);

FILL FILL_0__13163_ (
);

FILL FILL_1__6720_ (
);

FILL FILL_0__8549_ (
);

FILL FILL_3__6646_ (
);

FILL FILL_1__9192_ (
);

FILL FILL_1__12903_ (
);

FILL FILL_2__9928_ (
);

FILL FILL_0__9910_ (
);

FILL FILL_2__9508_ (
);

FILL FILL_1__10090_ (
);

FILL FILL_1__7925_ (
);

FILL FILL_1__7505_ (
);

INVX1 _6995_ (
    .A(_585_),
    .Y(_589_)
);

NAND3X1 _6575_ (
    .A(_162_),
    .B(_166_),
    .C(_168_),
    .Y(_175_)
);

FILL FILL_1__11295_ (
);

INVX1 _10993_ (
    .A(_4187_),
    .Y(_4192_)
);

NOR2X1 _10573_ (
    .A(_3839_),
    .B(_3838_),
    .Y(_3840_)
);

FILL FILL_0__10288_ (
);

OAI21X1 _10153_ (
    .A(_3277_),
    .B(_3262_),
    .C(_3346_),
    .Y(_3432_)
);

FILL FILL_3__11202_ (
);

FILL FILL_2__9681_ (
);

FILL FILL_2__10615_ (
);

FILL FILL_2__9261_ (
);

FILL FILL_2__13087_ (
);

FILL FILL_0__6615_ (
);

OAI21X1 _8721_ (
    .A(_1899_),
    .B(_2073_),
    .C(_2117_),
    .Y(_2155_)
);

NAND3X1 _8301_ (
    .A(_1740_),
    .B(_1734_),
    .C(_1737_),
    .Y(_1741_)
);

FILL FILL_0__9087_ (
);

NAND3X1 _11778_ (
    .A(_4894_),
    .B(_4888_),
    .C(_4892_),
    .Y(_4899_)
);

NOR2X1 _11358_ (
    .A(_4129_),
    .B(_4290_),
    .Y(_4552_)
);

FILL FILL_3__12827_ (
);

FILL FILL_1__13021_ (
);

FILL FILL_0__12854_ (
);

FILL FILL_0__12434_ (
);

FILL FILL_0__12014_ (
);

NAND3X1 _9926_ (
    .A(_3208_),
    .B(_3974_),
    .C(_3207_),
    .Y(_3209_)
);

NOR2X1 _9506_ (
    .A(_2797_),
    .B(_2794_),
    .Y(_2862_)
);

FILL FILL_1__8883_ (
);

FILL FILL_1__8463_ (
);

FILL FILL_1__8043_ (
);

FILL FILL_3__8389_ (
);

FILL FILL_3__9750_ (
);

FILL FILL_0__13219_ (
);

FILL FILL_2__6386_ (
);

FILL FILL_1__9668_ (
);

FILL FILL_1__9248_ (
);

FILL FILL_3__12580_ (
);

FILL FILL_2__11993_ (
);

FILL FILL_2__11573_ (
);

FILL FILL_2__11153_ (
);

FILL FILL_1__10986_ (
);

FILL FILL_1__10566_ (
);

FILL FILL_1__10146_ (
);

FILL FILL_0__7993_ (
);

FILL FILL_0__7573_ (
);

FILL FILL_0__7153_ (
);

FILL FILL_2__8952_ (
);

FILL FILL_2__8532_ (
);

FILL FILL_0__10920_ (
);

FILL FILL_0__10500_ (
);

FILL FILL_2__12778_ (
);

FILL FILL_2__12358_ (
);

FILL FILL_0__8778_ (
);

FILL FILL_3__6875_ (
);

FILL FILL_0__8358_ (
);

NOR2X1 _10629_ (
    .A(_3881_),
    .B(_3880_),
    .Y(_3893_)
);

AOI21X1 _10209_ (
    .A(_3469_),
    .B(_3471_),
    .C(_3486_),
    .Y(_3487_)
);

FILL FILL_1__12712_ (
);

FILL FILL_2__9737_ (
);

FILL FILL_2__9317_ (
);

FILL FILL_0__11705_ (
);

FILL FILL_1__7734_ (
);

FILL FILL_1__7314_ (
);

AOI22X1 _6384_ (
    .A(Xin[0]),
    .B(vdd),
    .C(Xin[1]),
    .D(gnd),
    .Y(_750_)
);

FILL FILL_3__8601_ (
);

AND2X2 _10382_ (
    .A(_3654_),
    .B(_3657_),
    .Y(_3658_)
);

FILL FILL_0__10097_ (
);

FILL FILL_1__8939_ (
);

FILL FILL_3__11851_ (
);

FILL FILL_1__8519_ (
);

FILL FILL_3__11431_ (
);

FILL FILL_2__10844_ (
);

FILL FILL_2__9490_ (
);

FILL FILL_2__10424_ (
);

FILL FILL_2__9070_ (
);

FILL FILL_2__10004_ (
);

OAI21X1 _7589_ (
    .A(_1105_),
    .B(_1106_),
    .C(_1101_),
    .Y(_1107_)
);

NOR2X1 _7169_ (
    .A(_751_),
    .B(_752_),
    .Y(_753_)
);

FILL FILL_0__6844_ (
);

NOR2X1 _8950_ (
    .A(_2371_),
    .B(_2314_),
    .Y(_2386_[1])
);

FILL FILL_0__6424_ (
);

NAND2X1 _8530_ (
    .A(_1967_),
    .B(_1891_),
    .Y(_1968_)
);

DFFPOSX1 _8110_ (
    .D(\Y[1] [10]),
    .CLK(clk_bF$buf54),
    .Q(\u_fir_pe1.rYin [10])
);

DFFPOSX1 _11587_ (
    .D(_4775_[3]),
    .CLK(clk_bF$buf48),
    .Q(\Y[6] [3])
);

INVX1 _11167_ (
    .A(_4357_),
    .Y(_4364_)
);

FILL FILL_2__7803_ (
);

FILL FILL_3__12216_ (
);

FILL FILL_1__13250_ (
);

FILL FILL_0__12663_ (
);

FILL FILL_2__11209_ (
);

FILL FILL_0__12243_ (
);

FILL FILL_0__7629_ (
);

NOR2X1 _9735_ (
    .A(_3075_),
    .B(_3074_),
    .Y(_3078_)
);

OAI21X1 _9315_ (
    .A(_2660_),
    .B(_2664_),
    .C(_2667_),
    .Y(_2674_)
);

FILL FILL_1__8692_ (
);

FILL FILL_1__8272_ (
);

FILL FILL_0__13028_ (
);

AND2X2 _13313_ (
    .A(_6336_),
    .B(_6335_),
    .Y(_6369_[13])
);

FILL FILL_1_CLKBUF1_insert12 (
);

FILL FILL_1_CLKBUF1_insert13 (
);

FILL FILL_1_CLKBUF1_insert14 (
);

FILL FILL_1__9897_ (
);

FILL FILL_1__9477_ (
);

FILL FILL_1_CLKBUF1_insert15 (
);

FILL FILL_1__9057_ (
);

FILL FILL_1_CLKBUF1_insert16 (
);

FILL FILL_1_CLKBUF1_insert17 (
);

FILL FILL_1_CLKBUF1_insert18 (
);

FILL FILL254550x36150 (
);

FILL FILL_1_CLKBUF1_insert19 (
);

FILL FILL_2__11382_ (
);

FILL FILL_1__10795_ (
);

FILL FILL_1__10375_ (
);

FILL FILL_0__7382_ (
);

FILL FILL_2__8761_ (
);

FILL FILL_2__8341_ (
);

FILL FILL_3__13174_ (
);

FILL FILL_2__12587_ (
);

FILL FILL_2__12167_ (
);

OAI22X1 _7801_ (
    .A(_1214_),
    .B(_1259_),
    .C(_1315_),
    .D(_1314_),
    .Y(_1316_)
);

FILL FILL254250x43350 (
);

FILL FILL_0__8587_ (
);

FILL FILL_0__8167_ (
);

INVX2 _10858_ (
    .A(\X[5]_5_bF$buf1 ),
    .Y(_4059_)
);

NAND2X1 _10438_ (
    .A(_3519_),
    .B(_3593_),
    .Y(_3713_)
);

NAND3X1 _10018_ (
    .A(_3214_),
    .B(_3294_),
    .C(_3298_),
    .Y(_3299_)
);

FILL FILL_1__12941_ (
);

FILL FILL_1__12521_ (
);

FILL FILL_1__12101_ (
);

FILL FILL_2__9966_ (
);

FILL FILL_0__11934_ (
);

FILL FILL_2__9546_ (
);

FILL FILL_2__9126_ (
);

FILL FILL_0__11514_ (
);

FILL FILL_1__7963_ (
);

FILL FILL_1__7543_ (
);

FILL FILL_1__7123_ (
);

FILL FILL_1__13306_ (
);

FILL FILL_3__8830_ (
);

FILL FILL_0__12719_ (
);

FILL FILL_3__10299_ (
);

NAND3X1 _10191_ (
    .A(_3397_),
    .B(_3465_),
    .C(_3466_),
    .Y(_3470_)
);

FILL FILL_1__8748_ (
);

FILL FILL_3__11660_ (
);

FILL FILL_1__8328_ (
);

FILL FILL_2__10653_ (
);

FILL FILL_2__10233_ (
);

NAND3X1 _7398_ (
    .A(_918_),
    .B(_851_),
    .C(_854_),
    .Y(_919_)
);

FILL FILL_3__9615_ (
);

FILL FILL_0__6653_ (
);

NAND2X1 _11396_ (
    .A(_4587_),
    .B(_4588_),
    .Y(_4589_)
);

FILL FILL_2__7612_ (
);

FILL FILL_3__12445_ (
);

FILL FILL_2__11858_ (
);

FILL FILL_0__12892_ (
);

FILL FILL_2__11438_ (
);

FILL FILL_2__11018_ (
);

FILL FILL_0__12052_ (
);

FILL FILL_0__7858_ (
);

NAND2X1 _9964_ (
    .A(_3242_),
    .B(_3245_),
    .Y(_3246_)
);

FILL FILL_0__7438_ (
);

OAI21X1 _9544_ (
    .A(_2899_),
    .B(_2767_),
    .C(_2849_),
    .Y(_2900_)
);

FILL FILL_0__7018_ (
);

NAND3X1 _9124_ (
    .A(gnd),
    .B(\X[3] [2]),
    .C(_2484_),
    .Y(_2485_)
);

FILL FILL_2__8817_ (
);

FILL FILL_0__13257_ (
);

NAND2X1 _13122_ (
    .A(_6142_),
    .B(_6155_),
    .Y(_6156_)
);

FILL FILL_1__6814_ (
);

FILL FILL_1__9286_ (
);

FILL FILL_2__11191_ (
);

FILL FILL_1__10184_ (
);

FILL FILL_0__7191_ (
);

FILL FILL_3__10931_ (
);

FILL FILL_3__10511_ (
);

FILL FILL_2__8570_ (
);

FILL FILL_2__8150_ (
);

NAND3X1 _6669_ (
    .A(_266_),
    .B(_267_),
    .C(_265_),
    .Y(_268_)
);

FILL FILL_2__12396_ (
);

AND2X2 _7610_ (
    .A(vdd),
    .B(\X[1] [6]),
    .Y(_1128_)
);

FILL FILL_1__11389_ (
);

FILL FILL_0__8396_ (
);

FILL FILL_3__6493_ (
);

INVX1 _10667_ (
    .A(\u_fir_pe4.mul [12]),
    .Y(_3931_)
);

AOI21X1 _10247_ (
    .A(_3434_),
    .B(_3437_),
    .C(_3443_),
    .Y(_3525_)
);

FILL FILL_3__11716_ (
);

FILL FILL_1__12750_ (
);

FILL FILL_1__12330_ (
);

FILL FILL_2__9775_ (
);

FILL FILL_2__9355_ (
);

FILL FILL_0__11743_ (
);

FILL FILL_0__11323_ (
);

FILL FILL_0__6709_ (
);

INVX1 _8815_ (
    .A(\u_fir_pe2.rYin [3]),
    .Y(_2242_)
);

FILL FILL_1__7772_ (
);

FILL FILL_1__7352_ (
);

FILL FILL_3__7698_ (
);

FILL FILL_3__7278_ (
);

FILL FILL_1__13115_ (
);

FILL FILL_0__12948_ (
);

AOI21X1 _12813_ (
    .A(_5851_),
    .B(_5850_),
    .C(_5849_),
    .Y(_5852_)
);

FILL FILL_0__12528_ (
);

FILL FILL_0__12108_ (
);

FILL FILL_1__8557_ (
);

FILL FILL_1__8137_ (
);

FILL FILL_2__10882_ (
);

FILL FILL_2__10462_ (
);

FILL FILL_2__10042_ (
);

FILL FILL_0__6882_ (
);

FILL FILL_0__6462_ (
);

FILL FILL_2__7841_ (
);

FILL FILL_3__12674_ (
);

FILL FILL_2__7421_ (
);

FILL FILL_2__7001_ (
);

FILL FILL_2__11667_ (
);

FILL FILL_2__11247_ (
);

FILL FILL_0__12281_ (
);

FILL FILL_0__7667_ (
);

NOR2X1 _9773_ (
    .A(_3115_),
    .B(_3116_),
    .Y(_3117_)
);

OAI21X1 _9353_ (
    .A(_2406_),
    .B(_2710_),
    .C(_2416_),
    .Y(_2711_)
);

FILL FILL_2__8626_ (
);

FILL FILL_2__8206_ (
);

FILL FILL_3__13039_ (
);

FILL FILL_0__13066_ (
);

DFFPOSX1 _13351_ (
    .D(_6369_[13]),
    .CLK(clk_bF$buf9),
    .Q(\Y[7] [13])
);

FILL FILL_1__6623_ (
);

FILL FILL_3__6969_ (
);

FILL FILL_1__9095_ (
);

FILL FILL_1__12806_ (
);

FILL FILL_0__9813_ (
);

FILL FILL_1__7828_ (
);

FILL FILL_1__7408_ (
);

FILL FILL_3__10320_ (
);

NAND3X1 _6898_ (
    .A(_423_),
    .B(_426_),
    .C(_493_),
    .Y(_494_)
);

NAND2X1 _6478_ (
    .A(gnd),
    .B(Xin_5_bF$buf1),
    .Y(_79_)
);

FILL FILL_1__11198_ (
);

INVX1 _10896_ (
    .A(_4011_),
    .Y(_4097_)
);

OAI21X1 _10476_ (
    .A(_3718_),
    .B(_3712_),
    .C(_3722_),
    .Y(_3750_)
);

NAND3X1 _10056_ (
    .A(gnd),
    .B(\X[4] [6]),
    .C(_3333_),
    .Y(_3336_)
);

FILL FILL_3__11945_ (
);

FILL FILL_3__11525_ (
);

FILL FILL_2__10938_ (
);

FILL FILL_0__11972_ (
);

FILL FILL_2__9584_ (
);

FILL FILL_2__10518_ (
);

FILL FILL_2__9164_ (
);

FILL FILL_0__11552_ (
);

FILL FILL_0__11132_ (
);

FILL FILL_0__6938_ (
);

FILL FILL_0__6518_ (
);

OAI22X1 _8624_ (
    .A(_1609_),
    .B(_2056_),
    .C(_2057_),
    .D(_2059_),
    .Y(_2060_)
);

NAND3X1 _8204_ (
    .A(_1622_),
    .B(_1645_),
    .C(_1644_),
    .Y(_1646_)
);

FILL FILL_1__7581_ (
);

FILL FILL_1__7161_ (
);

FILL FILL_3__7087_ (
);

FILL FILL_0__12757_ (
);

OAI22X1 _12622_ (
    .A(_6310_),
    .B(_5662_),
    .C(_5612_),
    .D(_5617_),
    .Y(_5663_)
);

FILL FILL_0__12337_ (
);

NAND3X1 _12202_ (
    .A(_5311_),
    .B(_5316_),
    .C(_5315_),
    .Y(_5317_)
);

NOR2X1 _9829_ (
    .A(_3170_),
    .B(_3177_),
    .Y(_3184_[2])
);

AOI21X1 _9409_ (
    .A(_2680_),
    .B(_2595_),
    .C(_2766_),
    .Y(_2767_)
);

FILL FILL_1__8786_ (
);

FILL FILL_1__8366_ (
);

FILL FILL_2__10691_ (
);

FILL FILL_2__10271_ (
);

FILL FILL_3__9233_ (
);

BUFX2 _13407_ (
    .A(_6377_[13]),
    .Y(Yout[13])
);

FILL FILL_0__6691_ (
);

FILL FILL_2__7650_ (
);

FILL FILL_3__12063_ (
);

FILL FILL_2__11896_ (
);

FILL FILL_2__11476_ (
);

FILL FILL_2__11056_ (
);

FILL FILL_0__12090_ (
);

FILL FILL_1__10889_ (
);

FILL FILL_1__10469_ (
);

FILL FILL_1__10049_ (
);

FILL FILL_0__7896_ (
);

FILL FILL_0__7476_ (
);

NAND3X1 _9582_ (
    .A(_2934_),
    .B(_2936_),
    .C(_2935_),
    .Y(_2937_)
);

FILL FILL_0__7056_ (
);

AND2X2 _9162_ (
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2522_)
);

FILL FILL_1__11830_ (
);

FILL FILL_1__11410_ (
);

FILL FILL_2__8855_ (
);

FILL FILL_2__8435_ (
);

FILL FILL_0__10823_ (
);

FILL FILL_3__13268_ (
);

FILL FILL_0__10403_ (
);

FILL FILL_2__8015_ (
);

FILL FILL_0__13295_ (
);

NAND2X1 _13160_ (
    .A(_6192_),
    .B(_6189_),
    .Y(_6375_[13])
);

FILL FILL_1__6852_ (
);

FILL FILL_1__6432_ (
);

FILL FILL_2__13202_ (
);

FILL FILL_1__12615_ (
);

FILL FILL254550x86550 (
);

FILL FILL_0__9622_ (
);

FILL FILL_0__9202_ (
);

FILL FILL_1__7637_ (
);

FILL FILL_3__8924_ (
);

FILL FILL_3__8504_ (
);

OAI21X1 _10285_ (
    .A(_3390_),
    .B(_3480_),
    .C(_3476_),
    .Y(_3563_)
);

FILL FILL_2__6921_ (
);

FILL FILL_2__6501_ (
);

FILL FILL_2__9393_ (
);

FILL FILL_0__11781_ (
);

FILL FILL_2__10327_ (
);

FILL FILL_0__11361_ (
);

FILL FILL_3__9709_ (
);

FILL FILL_0__6747_ (
);

INVX1 _8853_ (
    .A(\u_fir_pe2.mul [7]),
    .Y(_2276_)
);

NAND3X1 _8433_ (
    .A(_1816_),
    .B(_1857_),
    .C(_1862_),
    .Y(_1872_)
);

AOI21X1 _8013_ (
    .A(_1511_),
    .B(_1489_),
    .C(_1509_),
    .Y(_1516_)
);

FILL FILL_1__7390_ (
);

FILL FILL_2__7706_ (
);

FILL FILL_3__12539_ (
);

FILL FILL_1__13153_ (
);

FILL FILL_0__12986_ (
);

OAI21X1 _12851_ (
    .A(_5887_),
    .B(_5888_),
    .C(_5883_),
    .Y(_5889_)
);

FILL FILL_0__12566_ (
);

FILL FILL_0__12146_ (
);

NOR2X1 _12431_ (
    .A(_5533_),
    .B(_5534_),
    .Y(_5535_)
);

INVX1 _12011_ (
    .A(_5042_),
    .Y(_5129_)
);

OR2X2 _9638_ (
    .A(_2963_),
    .B(_2989_),
    .Y(_2991_)
);

NAND3X1 _9218_ (
    .A(_2575_),
    .B(_2576_),
    .C(_2577_),
    .Y(_2578_)
);

FILL FILL_1__8595_ (
);

FILL FILL_1__8175_ (
);

FILL FILL_2__10080_ (
);

FILL FILL_3__9462_ (
);

OR2X2 _13216_ (
    .A(_6240_),
    .B(_6238_),
    .Y(_6242_)
);

FILL FILL_1__6908_ (
);

FILL FILL_3__12292_ (
);

FILL FILL_2__11285_ (
);

FILL FILL_1__10698_ (
);

FILL FILL_1__10278_ (
);

FILL FILL_0__7285_ (
);

INVX1 _9391_ (
    .A(_2662_),
    .Y(_2749_)
);

FILL FILL_2__8664_ (
);

FILL FILL_2__8244_ (
);

FILL FILL_0__10632_ (
);

FILL FILL_0__10212_ (
);

NAND2X1 _7704_ (
    .A(_1212_),
    .B(_1219_),
    .Y(_1221_)
);

FILL FILL_1__6661_ (
);

FILL FILL_2__13011_ (
);

FILL FILL_3__6587_ (
);

FILL FILL_1__12844_ (
);

FILL FILL_1__12424_ (
);

FILL FILL_1__12004_ (
);

FILL FILL_0__9431_ (
);

FILL FILL_2__9449_ (
);

FILL FILL_0__11837_ (
);

FILL FILL_2__9029_ (
);

FILL FILL_0__9011_ (
);

NAND2X1 _11702_ (
    .A(vdd),
    .B(\X[7] [2]),
    .Y(_4824_)
);

FILL FILL_0__11417_ (
);

AOI21X1 _8909_ (
    .A(_2329_),
    .B(_2320_),
    .C(_2327_),
    .Y(_2332_)
);

FILL FILL_1__7866_ (
);

FILL FILL_1__7446_ (
);

FILL FILL_1__7026_ (
);

FILL FILL_1__13209_ (
);

AOI21X1 _12907_ (
    .A(_5944_),
    .B(_5943_),
    .C(_5879_),
    .Y(_5945_)
);

NAND3X1 _10094_ (
    .A(_3360_),
    .B(_3364_),
    .C(_3367_),
    .Y(_3374_)
);

FILL FILL_3__11983_ (
);

FILL FILL_2__6730_ (
);

FILL FILL_3__11143_ (
);

FILL FILL_2__10976_ (
);

FILL FILL_2__10556_ (
);

FILL FILL_2__10136_ (
);

FILL FILL_0__11170_ (
);

FILL FILL_0__6976_ (
);

FILL FILL_0__6556_ (
);

AOI21X1 _8662_ (
    .A(_2025_),
    .B(_2031_),
    .C(_2097_),
    .Y(_2098_)
);

INVX1 _8242_ (
    .A(gnd),
    .Y(_1683_)
);

FILL FILL_1__10910_ (
);

NOR2X1 _11299_ (
    .A(_4490_),
    .B(_4494_),
    .Y(_4495_)
);

FILL FILL_2__7935_ (
);

FILL FILL_3__12768_ (
);

FILL FILL_2__7515_ (
);

FILL FILL_0__12795_ (
);

NAND3X1 _12660_ (
    .A(_5700_),
    .B(_5633_),
    .C(_5636_),
    .Y(_5701_)
);

FILL FILL_0__12375_ (
);

NAND3X1 _12240_ (
    .A(_5346_),
    .B(_5353_),
    .C(_5352_),
    .Y(_5354_)
);

FILL FILL_2__12702_ (
);

DFFPOSX1 _9867_ (
    .D(\Y[3] [13]),
    .CLK(clk_bF$buf12),
    .Q(\u_fir_pe3.rYin [13])
);

OAI21X1 _9447_ (
    .A(_2724_),
    .B(_2803_),
    .C(_2802_),
    .Y(_2804_)
);

INVX1 _9027_ (
    .A(_3178_),
    .Y(_3179_)
);

FILL FILL_0__8702_ (
);

FILL FILL_3__9691_ (
);

NAND3X1 _13025_ (
    .A(_6059_),
    .B(_6060_),
    .C(_6058_),
    .Y(_6061_)
);

FILL FILL_1__6717_ (
);

FILL FILL_1__9189_ (
);

FILL FILL_0__9907_ (
);

FILL FILL_2__11094_ (
);

FILL FILL_1__10087_ (
);

FILL FILL_0__7094_ (
);

FILL FILL_3__10414_ (
);

FILL FILL_2__8893_ (
);

FILL FILL_2__8473_ (
);

FILL FILL_0__10861_ (
);

FILL FILL_0__10441_ (
);

FILL FILL_2__8053_ (
);

FILL FILL_0__10021_ (
);

FILL FILL_2__12299_ (
);

INVX1 _7933_ (
    .A(_1437_),
    .Y(_1441_)
);

INVX1 _7513_ (
    .A(\X[1] [7]),
    .Y(_1032_)
);

FILL FILL_1__6890_ (
);

FILL FILL_1__6470_ (
);

FILL FILL_2__13240_ (
);

FILL FILL_0__8299_ (
);

FILL FILL_1__12653_ (
);

FILL FILL_1__12233_ (
);

FILL FILL_0__9660_ (
);

FILL FILL_2__9678_ (
);

FILL FILL_0__9240_ (
);

FILL FILL_2__9258_ (
);

NAND3X1 _11931_ (
    .A(_5048_),
    .B(_5049_),
    .C(_5047_),
    .Y(_5050_)
);

FILL FILL_0__11646_ (
);

INVX1 _11511_ (
    .A(_4690_),
    .Y(_4694_)
);

FILL FILL_0__11226_ (
);

OAI21X1 _8718_ (
    .A(_2105_),
    .B(_2146_),
    .C(_2145_),
    .Y(_2152_)
);

FILL FILL_1__7675_ (
);

FILL FILL_1__7255_ (
);

FILL FILL_1__13018_ (
);

FILL FILL_3__8542_ (
);

NAND3X1 _12716_ (
    .A(_5751_),
    .B(_5717_),
    .C(_5755_),
    .Y(_5756_)
);

FILL FILL_3__11372_ (
);

FILL FILL_2__10785_ (
);

FILL FILL_2__10365_ (
);

FILL FILL_1__9821_ (
);

FILL FILL_1__9401_ (
);

FILL FILL_0_CLKBUF1_insert20 (
);

FILL FILL_3__9327_ (
);

FILL FILL_0_CLKBUF1_insert21 (
);

FILL FILL_0_CLKBUF1_insert22 (
);

FILL FILL_0_CLKBUF1_insert23 (
);

FILL FILL_0_CLKBUF1_insert24 (
);

FILL FILL_0__6785_ (
);

INVX1 _8891_ (
    .A(_2313_),
    .Y(_2315_)
);

FILL FILL_0_CLKBUF1_insert25 (
);

NAND2X1 _8471_ (
    .A(_1904_),
    .B(_1908_),
    .Y(_1909_)
);

FILL FILL_0_CLKBUF1_insert26 (
);

FILL FILL_0_CLKBUF1_insert27 (
);

AND2X2 _8051_ (
    .A(_1554_),
    .B(_1553_),
    .Y(_1587_[13])
);

FILL FILL_0_CLKBUF1_insert28 (
);

FILL FILL_0_CLKBUF1_insert29 (
);

FILL FILL_3__12997_ (
);

FILL FILL_2__7744_ (
);

FILL FILL_2__7324_ (
);

FILL FILL_3__12157_ (
);

FILL FILL_1__13191_ (
);

FILL FILL_0__12184_ (
);

FILL FILL_2__12931_ (
);

NOR2X1 _9676_ (
    .A(_3023_),
    .B(_3024_),
    .Y(_3025_)
);

OAI21X1 _9256_ (
    .A(_2564_),
    .B(_2614_),
    .C(_2558_),
    .Y(_2615_)
);

FILL FILL_1__11924_ (
);

FILL FILL_1__11504_ (
);

FILL FILL_0__8931_ (
);

FILL FILL_2__8949_ (
);

FILL FILL_2__8529_ (
);

FILL FILL_0__8511_ (
);

FILL FILL_0__10917_ (
);

FILL FILL_3__9080_ (
);

AND2X2 _13254_ (
    .A(_6256_),
    .B(_6266_),
    .Y(_6277_)
);

FILL FILL_1__6946_ (
);

FILL FILL_1__6526_ (
);

FILL FILL_1__12709_ (
);

FILL FILL_0__9716_ (
);

FILL FILL_3__7813_ (
);

FILL FILL_2__8282_ (
);

FILL FILL_0__10670_ (
);

FILL FILL_0__10250_ (
);

OAI21X1 _7742_ (
    .A(_1224_),
    .B(_1226_),
    .C(_1220_),
    .Y(_1258_)
);

NAND2X1 _7322_ (
    .A(_841_),
    .B(_837_),
    .Y(_844_)
);

OAI21X1 _10799_ (
    .A(_4763_),
    .B(_4000_),
    .C(_4001_),
    .Y(_4002_)
);

NOR2X1 _10379_ (
    .A(_3203_),
    .B(_3650_),
    .Y(_3655_)
);

FILL FILL_1__12882_ (
);

FILL FILL_3__11008_ (
);

FILL FILL_1__12042_ (
);

FILL FILL_2__9487_ (
);

FILL FILL_0__11875_ (
);

FILL FILL_2__9067_ (
);

NAND2X1 _11740_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf2 ),
    .Y(_4861_)
);

FILL FILL_0__11455_ (
);

FILL FILL_0__11035_ (
);

INVX1 _11320_ (
    .A(_4514_),
    .Y(_4515_)
);

NOR2X1 _8947_ (
    .A(\u_fir_pe2.rYin [0]),
    .B(\u_fir_pe2.mul [0]),
    .Y(_2370_)
);

NAND3X1 _8527_ (
    .A(_1895_),
    .B(_1956_),
    .C(_1951_),
    .Y(_1965_)
);

DFFPOSX1 _8107_ (
    .D(\Y[1] [7]),
    .CLK(clk_bF$buf32),
    .Q(\u_fir_pe1.rYin [7])
);

FILL FILL_1__7484_ (
);

FILL FILL_1__7064_ (
);

FILL FILL_1__13247_ (
);

FILL FILL_3__8771_ (
);

OAI22X1 _12945_ (
    .A(_5833_),
    .B(_5980_),
    .C(_5903_),
    .D(_5981_),
    .Y(_5982_)
);

INVX1 _12525_ (
    .A(\X[6] [2]),
    .Y(_6349_)
);

AOI21X1 _12105_ (
    .A(_5212_),
    .B(_5208_),
    .C(_5167_),
    .Y(_5222_)
);

FILL FILL_1__8689_ (
);

FILL FILL_1__8269_ (
);

FILL FILL_2__10594_ (
);

FILL FILL_2__10174_ (
);

FILL FILL_1__9630_ (
);

FILL FILL_1__9210_ (
);

FILL FILL_3__9976_ (
);

FILL FILL_3__9556_ (
);

FILL FILL_0__6594_ (
);

INVX1 _8280_ (
    .A(_1661_),
    .Y(_1721_)
);

FILL FILL_2__7973_ (
);

FILL FILL_2__7553_ (
);

FILL FILL_3__12386_ (
);

FILL FILL_2__7133_ (
);

FILL FILL_2__11799_ (
);

FILL FILL_2__11379_ (
);

FILL FILL_2__12740_ (
);

FILL FILL_2__12320_ (
);

FILL FILL_0__7799_ (
);

FILL FILL_0__7379_ (
);

OR2X2 _9485_ (
    .A(_2771_),
    .B(_2841_),
    .Y(_2842_)
);

AND2X2 _9065_ (
    .A(gnd),
    .B(\X[3] [2]),
    .Y(_2427_)
);

FILL FILL_1__11733_ (
);

FILL FILL_1__11313_ (
);

FILL FILL_0__8740_ (
);

FILL FILL_2__8758_ (
);

FILL FILL_0__8320_ (
);

FILL FILL_2__8338_ (
);

FILL FILL_0__10306_ (
);

FILL FILL_0__13198_ (
);

OAI22X1 _13063_ (
    .A(_5996_),
    .B(_6041_),
    .C(_6097_),
    .D(_6096_),
    .Y(_6098_)
);

FILL FILL_1__6755_ (
);

FILL FILL_2__13105_ (
);

FILL FILL_1__12938_ (
);

FILL FILL_1__12518_ (
);

FILL FILL_0__9945_ (
);

FILL FILL_0__9525_ (
);

FILL FILL_0__9105_ (
);

FILL FILL_3__10872_ (
);

FILL FILL_3__10452_ (
);

FILL FILL_3__10032_ (
);

FILL FILL_1__8901_ (
);

NAND2X1 _7971_ (
    .A(_1474_),
    .B(_1469_),
    .Y(_1475_)
);

AOI21X1 _7551_ (
    .A(_1069_),
    .B(_1068_),
    .C(_1067_),
    .Y(_1070_)
);

INVX1 _7131_ (
    .A(_714_),
    .Y(_715_)
);

NAND3X1 _10188_ (
    .A(_3465_),
    .B(_3466_),
    .C(_3464_),
    .Y(_3467_)
);

FILL FILL_2__6824_ (
);

FILL FILL_3__11657_ (
);

FILL FILL_2__6404_ (
);

FILL FILL_1__12691_ (
);

FILL FILL_3__11237_ (
);

FILL FILL_1__12271_ (
);

FILL FILL_2__9296_ (
);

FILL FILL_0__11684_ (
);

FILL FILL_0__11264_ (
);

FILL FILL254550x172950 (
);

NOR2X1 _8756_ (
    .A(_1829_),
    .B(_2056_),
    .Y(_2189_)
);

OAI21X1 _8336_ (
    .A(_1774_),
    .B(_1775_),
    .C(_1773_),
    .Y(_1776_)
);

FILL FILL_1__7293_ (
);

FILL FILL_2__7609_ (
);

FILL FILL_1__13056_ (
);

FILL FILL_0__12889_ (
);

AND2X2 _12754_ (
    .A(_5724_),
    .B(_5728_),
    .Y(_5793_)
);

FILL FILL_3__8160_ (
);

FILL FILL_0__12049_ (
);

NOR2X1 _12334_ (
    .A(\u_fir_pe6.rYin [4]),
    .B(\u_fir_pe6.mul [4]),
    .Y(_5440_)
);

FILL FILL_0__13410_ (
);

FILL FILL_1__8498_ (
);

FILL FILL_3__9785_ (
);

INVX1 _13119_ (
    .A(_6150_),
    .Y(_6153_)
);

FILL FILL_2__7782_ (
);

FILL FILL_2__7362_ (
);

FILL FILL_2__11188_ (
);

OAI21X1 _6822_ (
    .A(_25_),
    .B(_416_),
    .C(_418_),
    .Y(_419_)
);

INVX1 _6402_ (
    .A(_4_),
    .Y(_5_)
);

FILL FILL_0__7188_ (
);

AOI21X1 _9294_ (
    .A(_2652_),
    .B(_2651_),
    .C(_2650_),
    .Y(_2653_)
);

FILL FILL_1__11962_ (
);

FILL FILL_3__10508_ (
);

FILL FILL_1__11542_ (
);

FILL FILL_1__11122_ (
);

FILL FILL_2__8567_ (
);

FILL FILL_0__10955_ (
);

FILL FILL_2__8147_ (
);

FILL FILL_0__10535_ (
);

NAND2X1 _10820_ (
    .A(_4020_),
    .B(_4021_),
    .Y(_4022_)
);

NAND2X1 _10400_ (
    .A(_3657_),
    .B(_3654_),
    .Y(_3676_)
);

FILL FILL_0__10115_ (
);

AND2X2 _13292_ (
    .A(_6311_),
    .B(_6314_),
    .Y(_6316_)
);

OAI21X1 _7607_ (
    .A(_886_),
    .B(_941_),
    .C(_1124_),
    .Y(_1125_)
);

FILL FILL_1__6984_ (
);

FILL FILL_1__6564_ (
);

FILL FILL_2__13334_ (
);

FILL FILL_1__12747_ (
);

FILL FILL_1__12327_ (
);

FILL FILL_0__9754_ (
);

FILL FILL_0__9334_ (
);

FILL FILL_3__7431_ (
);

DFFPOSX1 _11605_ (
    .D(\X[5]_5_bF$buf2 ),
    .CLK(clk_bF$buf11),
    .Q(\X[6] [5])
);

FILL FILL_3__7011_ (
);

FILL FILL_1__7769_ (
);

FILL FILL_3__10681_ (
);

FILL FILL_1__7349_ (
);

FILL FILL_1__8710_ (
);

FILL FILL_3__8636_ (
);

FILL FILL_3__8216_ (
);

AND2X2 _7780_ (
    .A(_1284_),
    .B(_1288_),
    .Y(_1296_)
);

OAI22X1 _7360_ (
    .A(_1528_),
    .B(_880_),
    .C(_830_),
    .D(_835_),
    .Y(_881_)
);

FILL FILL_3__11886_ (
);

FILL FILL_2__6633_ (
);

FILL FILL_3__11466_ (
);

FILL FILL_1__12080_ (
);

FILL FILL_2__10879_ (
);

FILL FILL_2__10459_ (
);

FILL FILL_2__10039_ (
);

FILL FILL_0__11493_ (
);

FILL FILL_0__11073_ (
);

FILL FILL_1__9915_ (
);

FILL FILL_2__11820_ (
);

FILL FILL_0__6879_ (
);

FILL FILL_2__11400_ (
);

DFFPOSX1 _8985_ (
    .D(\Y[2] [8]),
    .CLK(clk_bF$buf12),
    .Q(\u_fir_pe2.rYin [8])
);

FILL FILL_0__6459_ (
);

AND2X2 _8565_ (
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_2002_)
);

NOR2X1 _8145_ (
    .A(_2374_),
    .B(_2354_),
    .Y(_2377_)
);

FILL FILL_1__10813_ (
);

FILL FILL_2__7838_ (
);

FILL FILL_0__7820_ (
);

FILL FILL_0__7400_ (
);

FILL FILL_2__7418_ (
);

FILL FILL_1__13285_ (
);

OAI21X1 _12983_ (
    .A(_6019_),
    .B(_6018_),
    .C(_6017_),
    .Y(_6020_)
);

FILL FILL_0__12698_ (
);

FILL FILL_0__12278_ (
);

NOR2X1 _12563_ (
    .A(_5603_),
    .B(_5604_),
    .Y(_5605_)
);

AND2X2 _12143_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5259_)
);

FILL FILL_2__12605_ (
);

FILL FILL_0__8605_ (
);

FILL FILL_3__9174_ (
);

DFFPOSX1 _13348_ (
    .D(_6369_[10]),
    .CLK(clk_bF$buf48),
    .Q(\Y[7] [10])
);

FILL FILL_2__7591_ (
);

FILL FILL_2__7171_ (
);

FILL FILL_3__7907_ (
);

AOI22X1 _6631_ (
    .A(gnd),
    .B(Xin[7]),
    .C(Xin[3]),
    .D(gnd),
    .Y(_230_)
);

FILL FILL_1__11771_ (
);

FILL FILL_1__11351_ (
);

FILL FILL_2__8796_ (
);

FILL FILL_2__8376_ (
);

FILL FILL_0__10764_ (
);

FILL FILL_0__10344_ (
);

NAND3X1 _7836_ (
    .A(_1308_),
    .B(_1350_),
    .C(_1309_),
    .Y(_1351_)
);

NAND2X1 _7416_ (
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_936_)
);

FILL FILL_1__6793_ (
);

FILL FILL_2__13143_ (
);

FILL FILL_1__12976_ (
);

FILL FILL_1__12556_ (
);

FILL FILL_1__12136_ (
);

FILL FILL_0__9983_ (
);

FILL FILL_0__9563_ (
);

FILL FILL_0__11969_ (
);

FILL FILL_3__7660_ (
);

FILL FILL_0__9143_ (
);

NAND3X1 _11834_ (
    .A(_4949_),
    .B(_4934_),
    .C(_4953_),
    .Y(_4954_)
);

FILL FILL_0__11549_ (
);

NAND2X1 _11414_ (
    .A(_4605_),
    .B(_4604_),
    .Y(_4606_)
);

FILL FILL_0__11129_ (
);

FILL FILL_0__12910_ (
);

FILL FILL_1__7998_ (
);

FILL FILL_1__7578_ (
);

FILL FILL_1__7158_ (
);

FILL FILL_3__10070_ (
);

FILL FILL_3__8865_ (
);

FILL FILL_3__8445_ (
);

NAND3X1 _12619_ (
    .A(_5649_),
    .B(_5657_),
    .C(_5659_),
    .Y(_5660_)
);

FILL FILL_3__8025_ (
);

FILL FILL_2__6862_ (
);

FILL FILL_2__6442_ (
);

FILL FILL_2__10688_ (
);

FILL FILL_2__10268_ (
);

FILL FILL_1__9724_ (
);

FILL FILL_1__9304_ (
);

FILL FILL_0__6688_ (
);

NAND2X1 _8794_ (
    .A(_2224_),
    .B(_2223_),
    .Y(_2390_[15])
);

AOI21X1 _8374_ (
    .A(_1741_),
    .B(_1737_),
    .C(_1806_),
    .Y(_1813_)
);

FILL FILL_1__10622_ (
);

FILL FILL_1__10202_ (
);

FILL FILL_2__7647_ (
);

FILL FILL_1__13094_ (
);

AOI22X1 _12792_ (
    .A(_5666_),
    .B(_5737_),
    .C(_5740_),
    .D(_5736_),
    .Y(_5831_)
);

FILL FILL_0__12087_ (
);

NOR2X1 _12372_ (
    .A(\u_fir_pe6.rYin [8]),
    .B(\u_fir_pe6.mul [8]),
    .Y(_5475_)
);

FILL FILL_3__13001_ (
);

FILL FILL_2__12834_ (
);

FILL FILL_2__12414_ (
);

NAND3X1 _9999_ (
    .A(gnd),
    .B(\X[4] [3]),
    .C(_3271_),
    .Y(_3280_)
);

INVX1 _9579_ (
    .A(_2906_),
    .Y(_2934_)
);

INVX1 _9159_ (
    .A(_2516_),
    .Y(_2520_)
);

FILL FILL_1__11827_ (
);

FILL FILL_1__11407_ (
);

FILL FILL_0__8834_ (
);

FILL FILL_0__8414_ (
);

FILL FILL_3__6511_ (
);

NAND2X1 _13157_ (
    .A(_6168_),
    .B(_6167_),
    .Y(_6190_)
);

FILL FILL_1__6849_ (
);

FILL FILL_1__6429_ (
);

FILL FILL_0__9619_ (
);

AOI21X1 _6860_ (
    .A(_441_),
    .B(_437_),
    .C(_382_),
    .Y(_456_)
);

NAND2X1 _6440_ (
    .A(vdd),
    .B(Xin[2]),
    .Y(_42_)
);

FILL FILL_3__10966_ (
);

FILL FILL_3__10546_ (
);

FILL FILL_1__11580_ (
);

FILL FILL_3__10126_ (
);

FILL FILL_1__11160_ (
);

FILL FILL_0__10993_ (
);

FILL FILL_2__8185_ (
);

FILL FILL_0__10573_ (
);

FILL FILL_0__10153_ (
);

FILL FILL_2__10900_ (
);

AOI21X1 _7645_ (
    .A(_1162_),
    .B(_1161_),
    .C(_1097_),
    .Y(_1163_)
);

DFFPOSX1 _7225_ (
    .D(Yin[2]),
    .CLK(clk_bF$buf20),
    .Q(\u_fir_pe0.rYin [2])
);

FILL FILL_0__6900_ (
);

FILL FILL_2__6918_ (
);

FILL FILL_1__12785_ (
);

FILL FILL_1__12365_ (
);

FILL FILL_0__9792_ (
);

FILL FILL_0__9372_ (
);

FILL FILL_0__11778_ (
);

NOR2X1 _11643_ (
    .A(_5471_),
    .B(_5492_),
    .Y(_5502_)
);

FILL FILL_0__11358_ (
);

AOI21X1 _11223_ (
    .A(_4410_),
    .B(_4408_),
    .C(_4380_),
    .Y(_4420_)
);

FILL FILL_1__7387_ (
);

OAI21X1 _12848_ (
    .A(_5804_),
    .B(_5809_),
    .C(_5808_),
    .Y(_5886_)
);

FILL FILL_3__8254_ (
);

OAI21X1 _12428_ (
    .A(_5524_),
    .B(_5525_),
    .C(_5529_),
    .Y(_5531_)
);

OAI21X1 _12008_ (
    .A(_5117_),
    .B(_5111_),
    .C(_5119_),
    .Y(_5126_)
);

FILL FILL_2__6671_ (
);

FILL FILL_3__11084_ (
);

FILL FILL_2__10497_ (
);

FILL FILL_2__10077_ (
);

FILL FILL_1__9953_ (
);

FILL FILL_1__9533_ (
);

FILL FILL_1__9113_ (
);

FILL FILL_3__9039_ (
);

FILL FILL_0__6497_ (
);

NAND2X1 _8183_ (
    .A(vdd),
    .B(\X[2] [1]),
    .Y(_1625_)
);

FILL FILL_1__10851_ (
);

FILL FILL_1__10431_ (
);

FILL FILL_1__10011_ (
);

FILL FILL_2__7876_ (
);

FILL FILL_2__7456_ (
);

FILL FILL_2__7036_ (
);

AOI21X1 _12181_ (
    .A(_5242_),
    .B(_5276_),
    .C(_5295_),
    .Y(_5296_)
);

FILL FILL_3__13230_ (
);

NAND3X1 _6916_ (
    .A(_495_),
    .B(_501_),
    .C(_459_),
    .Y(_511_)
);

FILL FILL_2__12643_ (
);

FILL FILL_2__12223_ (
);

OAI21X1 _9388_ (
    .A(_2732_),
    .B(_2736_),
    .C(_2739_),
    .Y(_2746_)
);

FILL FILL_1__11216_ (
);

FILL FILL_0__8643_ (
);

FILL FILL_3__6740_ (
);

FILL FILL_0__8223_ (
);

FILL FILL_0__10629_ (
);

OAI21X1 _10914_ (
    .A(_4113_),
    .B(_4114_),
    .C(_4112_),
    .Y(_4115_)
);

FILL FILL_0__10209_ (
);

DFFPOSX1 _13386_ (
    .D(_6375_[8]),
    .CLK(clk_bF$buf24),
    .Q(\u_fir_pe7.mul [8])
);

FILL FILL_2__9602_ (
);

FILL FILL_1__6658_ (
);

FILL FILL_2__13008_ (
);

FILL FILL_0__9428_ (
);

FILL FILL_3__7525_ (
);

FILL FILL_3__7105_ (
);

FILL FILL_3__10355_ (
);

FILL FILL_0__10382_ (
);

FILL FILL_1__8804_ (
);

NOR2X1 _7874_ (
    .A(_1383_),
    .B(_1387_),
    .Y(_1593_[12])
);

NAND3X1 _7454_ (
    .A(_969_),
    .B(_935_),
    .C(_973_),
    .Y(_974_)
);

INVX1 _7034_ (
    .A(_616_),
    .Y(_626_)
);

FILL FILL_2__13181_ (
);

FILL FILL_2__6727_ (
);

FILL FILL_1__12594_ (
);

FILL FILL_1__12174_ (
);

FILL FILL_2__9199_ (
);

FILL FILL_0__9181_ (
);

OAI21X1 _11872_ (
    .A(_4918_),
    .B(_4990_),
    .C(_4959_),
    .Y(_4991_)
);

OR2X2 _11452_ (
    .A(_4632_),
    .B(_4637_),
    .Y(_4639_)
);

FILL FILL_0__11167_ (
);

INVX1 _11032_ (
    .A(_4225_),
    .Y(_4231_)
);

FILL FILL_3__12921_ (
);

FILL FILL_2__11914_ (
);

NAND3X1 _8659_ (
    .A(_2090_),
    .B(_2091_),
    .C(_2094_),
    .Y(_2095_)
);

INVX1 _8239_ (
    .A(_1679_),
    .Y(_1680_)
);

FILL FILL_1__7196_ (
);

FILL FILL_1__10907_ (
);

FILL FILL_0__7914_ (
);

INVX1 _9600_ (
    .A(_2953_),
    .Y(_2954_)
);

FILL FILL_3__8483_ (
);

NAND3X1 _12657_ (
    .A(_5633_),
    .B(_5696_),
    .C(_5697_),
    .Y(_5698_)
);

AOI21X1 _12237_ (
    .A(gnd),
    .B(_5348_),
    .C(_5350_),
    .Y(_5351_)
);

FILL FILL_0__13313_ (
);

FILL FILL_2__6480_ (
);

FILL FILL_1__9762_ (
);

FILL FILL_1__9342_ (
);

FILL FILL_3__9268_ (
);

FILL FILL_1__10660_ (
);

FILL FILL_1__10240_ (
);

FILL FILL_2__7685_ (
);

FILL FILL_2__7265_ (
);

FILL FILL_3__12098_ (
);

OAI21X1 _6725_ (
    .A(_240_),
    .B(_248_),
    .C(_247_),
    .Y(_323_)
);

FILL FILL_2__12872_ (
);

FILL FILL_2__12452_ (
);

FILL FILL_2__12032_ (
);

NAND3X1 _9197_ (
    .A(_2547_),
    .B(_2554_),
    .C(_2556_),
    .Y(_2557_)
);

FILL FILL_1__11865_ (
);

FILL FILL_1__11445_ (
);

FILL FILL_1__11025_ (
);

FILL FILL_0__8872_ (
);

FILL FILL_0__8452_ (
);

FILL FILL_0__10858_ (
);

FILL FILL_0__10438_ (
);

DFFPOSX1 _10723_ (
    .D(\X[4] [0]),
    .CLK(clk_bF$buf35),
    .Q(\X[5] [0])
);

FILL FILL_0__8032_ (
);

INVX1 _10303_ (
    .A(_3574_),
    .Y(_3580_)
);

FILL FILL_0__10018_ (
);

INVX1 _13195_ (
    .A(_6219_),
    .Y(_6223_)
);

FILL FILL_2__9411_ (
);

FILL FILL_1__6887_ (
);

FILL FILL_1__6467_ (
);

FILL FILL_2__13237_ (
);

FILL FILL_0__9657_ (
);

FILL FILL_3__7754_ (
);

FILL FILL_0__9237_ (
);

AOI21X1 _11928_ (
    .A(_4934_),
    .B(_4953_),
    .C(_5046_),
    .Y(_5047_)
);

NAND2X1 _11508_ (
    .A(_4690_),
    .B(_4691_),
    .Y(_4692_)
);

FILL FILL_0__10191_ (
);

FILL FILL_1__8613_ (
);

FILL FILL_3__8539_ (
);

OAI22X1 _7683_ (
    .A(_1051_),
    .B(_1198_),
    .C(_1121_),
    .D(_1199_),
    .Y(_1200_)
);

INVX1 _7263_ (
    .A(\X[1] [2]),
    .Y(_1567_)
);

FILL FILL_3__9900_ (
);

FILL FILL_2__6956_ (
);

FILL FILL_2__6536_ (
);

INVX1 _11681_ (
    .A(_4803_),
    .Y(_4804_)
);

FILL FILL_0__11396_ (
);

OAI21X1 _11261_ (
    .A(_4404_),
    .B(_4456_),
    .C(_4392_),
    .Y(_4457_)
);

FILL FILL_1__9818_ (
);

FILL FILL_3__12310_ (
);

FILL FILL_2__11723_ (
);

FILL FILL_2__11303_ (
);

NAND2X1 _8888_ (
    .A(_2311_),
    .B(_2310_),
    .Y(_2384_[9])
);

OR2X2 _8468_ (
    .A(_1901_),
    .B(_1900_),
    .Y(_1906_)
);

NOR2X1 _8048_ (
    .A(_1551_),
    .B(_1550_),
    .Y(_1552_)
);

FILL FILL_0__7723_ (
);

FILL FILL_0__7303_ (
);

FILL FILL_1__13188_ (
);

AOI21X1 _12886_ (
    .A(_5923_),
    .B(_5922_),
    .C(_5921_),
    .Y(_5924_)
);

FILL FILL254550x104550 (
);

DFFPOSX1 _12466_ (
    .D(_5572_[5]),
    .CLK(clk_bF$buf22),
    .Q(_6377_[5])
);

AOI21X1 _12046_ (
    .A(_5143_),
    .B(_5142_),
    .C(_5085_),
    .Y(_5163_)
);

FILL FILL253950x183750 (
);

FILL FILL_2__12928_ (
);

FILL FILL_0__13122_ (
);

FILL FILL_0__8928_ (
);

FILL FILL_0__8508_ (
);

FILL FILL_3__6605_ (
);

FILL FILL_1__9991_ (
);

FILL FILL_1__9571_ (
);

FILL FILL_1__9151_ (
);

FILL FILL_3__9497_ (
);

FILL FILL_2__7494_ (
);

FILL FILL_2__7074_ (
);

AOI21X1 _6954_ (
    .A(_487_),
    .B(_491_),
    .C(_461_),
    .Y(_549_)
);

OR2X2 _6534_ (
    .A(_133_),
    .B(_131_),
    .Y(_134_)
);

FILL FILL_2__12681_ (
);

FILL FILL_2__12261_ (
);

FILL FILL_1__11674_ (
);

FILL FILL_1__11254_ (
);

FILL FILL_2__8699_ (
);

FILL FILL_0__8681_ (
);

FILL FILL_0__8261_ (
);

FILL FILL_2__8279_ (
);

FILL FILL_0__10667_ (
);

NAND3X1 _10952_ (
    .A(_4140_),
    .B(_4151_),
    .C(_4147_),
    .Y(_4152_)
);

OAI21X1 _10532_ (
    .A(_3772_),
    .B(_3797_),
    .C(_3796_),
    .Y(_3804_)
);

FILL FILL_0__10247_ (
);

AOI21X1 _10112_ (
    .A(_3308_),
    .B(_3314_),
    .C(_3391_),
    .Y(_3392_)
);

FILL FILL_2__9640_ (
);

FILL FILL_2__9220_ (
);

INVX1 _7739_ (
    .A(_1254_),
    .Y(_1255_)
);

NAND3X1 _7319_ (
    .A(_830_),
    .B(_838_),
    .C(_840_),
    .Y(_841_)
);

FILL FILL_1__6696_ (
);

FILL FILL_2__13046_ (
);

FILL FILL_1__12879_ (
);

FILL FILL_1__12459_ (
);

FILL FILL_1__12039_ (
);

FILL FILL_0__9886_ (
);

FILL FILL_3__7983_ (
);

FILL FILL_0__9466_ (
);

FILL FILL_0__9046_ (
);

OAI21X1 _11737_ (
    .A(_5560_),
    .B(_4856_),
    .C(_4857_),
    .Y(_4858_)
);

OAI22X1 _11317_ (
    .A(_4218_),
    .B(_4220_),
    .C(_4304_),
    .D(_4129_),
    .Y(_4512_)
);

FILL FILL_1__13400_ (
);

FILL FILL_0__12813_ (
);

FILL FILL_3__10393_ (
);

FILL FILL_1__8842_ (
);

FILL FILL_1__8422_ (
);

FILL FILL_1__8002_ (
);

AND2X2 _7492_ (
    .A(_942_),
    .B(_946_),
    .Y(_1011_)
);

NOR2X1 _7072_ (
    .A(\u_fir_pe0.rYin [4]),
    .B(\u_fir_pe0.mul [4]),
    .Y(_658_)
);

FILL FILL_2__6765_ (
);

FILL FILL_3__11178_ (
);

NAND2X1 _11490_ (
    .A(_4672_),
    .B(_4671_),
    .Y(_4673_)
);

AOI21X1 _11070_ (
    .A(_4268_),
    .B(_4267_),
    .C(_4266_),
    .Y(_4269_)
);

FILL FILL_1__9627_ (
);

FILL FILL_1__9207_ (
);

FILL FILL_2__11952_ (
);

FILL FILL_2__11532_ (
);

FILL FILL_2__11112_ (
);

AOI21X1 _8697_ (
    .A(_2009_),
    .B(_2001_),
    .C(_2079_),
    .Y(_2132_)
);

NAND3X1 _8277_ (
    .A(_1647_),
    .B(_1711_),
    .C(_1712_),
    .Y(_1718_)
);

FILL FILL_1__10945_ (
);

FILL FILL_1__10525_ (
);

FILL FILL_1__10105_ (
);

FILL FILL_0__7952_ (
);

FILL FILL_0__7532_ (
);

FILL FILL_0__7112_ (
);

NAND2X1 _12695_ (
    .A(gnd),
    .B(\X[6]_5_bF$buf3 ),
    .Y(_5735_)
);

OAI21X1 _12275_ (
    .A(_5345_),
    .B(_5358_),
    .C(_5362_),
    .Y(_5388_)
);

FILL FILL_2__8911_ (
);

FILL FILL_3__13324_ (
);

FILL FILL_2__12737_ (
);

FILL FILL_2__12317_ (
);

FILL FILL_0__8737_ (
);

FILL FILL_3__6834_ (
);

FILL FILL_0__8317_ (
);

FILL FILL_1__9380_ (
);

FILL FILL_3__7619_ (
);

NAND3X1 _6763_ (
    .A(_315_),
    .B(_346_),
    .C(_351_),
    .Y(_361_)
);

FILL FILL_2__12070_ (
);

FILL FILL_3__10449_ (
);

FILL FILL_1__11483_ (
);

FILL FILL_1__11063_ (
);

FILL FILL_0__8490_ (
);

FILL FILL_0__10896_ (
);

FILL FILL_0__10476_ (
);

DFFPOSX1 _10761_ (
    .D(_3984_[14]),
    .CLK(clk_bF$buf38),
    .Q(\u_fir_pe4.mul [14])
);

FILL FILL_0__8070_ (
);

OAI21X1 _10341_ (
    .A(_3617_),
    .B(_3616_),
    .C(_3615_),
    .Y(_3618_)
);

FILL FILL_0__10056_ (
);

FILL FILL_3__11810_ (
);

FILL FILL_2__10803_ (
);

NOR2X1 _7968_ (
    .A(_1470_),
    .B(_1471_),
    .Y(_1472_)
);

AND2X2 _7548_ (
    .A(_1018_),
    .B(_1015_),
    .Y(_1067_)
);

AND2X2 _7128_ (
    .A(\u_fir_pe0.rYin [9]),
    .B(\u_fir_pe0.mul [9]),
    .Y(_712_)
);

FILL FILL_2__13275_ (
);

FILL FILL_0__6803_ (
);

FILL FILL_1__12688_ (
);

FILL FILL_1__12268_ (
);

FILL FILL_0__9695_ (
);

FILL FILL_0__9275_ (
);

AOI21X1 _11966_ (
    .A(_5048_),
    .B(_5049_),
    .C(_5006_),
    .Y(_5084_)
);

FILL FILL_3__7372_ (
);

NOR2X1 _11546_ (
    .A(\u_fir_pe5.rYin [12]),
    .B(\u_fir_pe5.mul [12]),
    .Y(_4730_)
);

NAND3X1 _11126_ (
    .A(_4309_),
    .B(_4311_),
    .C(_4313_),
    .Y(_4324_)
);

FILL FILL_0__12622_ (
);

FILL FILL_0__12202_ (
);

FILL FILL_1__8651_ (
);

FILL FILL_1__8231_ (
);

FILL FILL_3__8577_ (
);

FILL FILL_3__8157_ (
);

FILL FILL_0__13407_ (
);

FILL FILL_2__6994_ (
);

FILL FILL_2__6574_ (
);

FILL FILL_1__9436_ (
);

FILL FILL_1__9016_ (
);

FILL FILL_2__11761_ (
);

FILL FILL_2__11341_ (
);

DFFPOSX1 _8086_ (
    .D(_1587_[10]),
    .CLK(clk_bF$buf10),
    .Q(\Y[2] [10])
);

FILL FILL_1__10334_ (
);

FILL FILL_0__7761_ (
);

FILL FILL_2__7779_ (
);

FILL FILL_0__7341_ (
);

FILL FILL_2__7359_ (
);

OAI21X1 _12084_ (
    .A(_4807_),
    .B(_5198_),
    .C(_5200_),
    .Y(_5201_)
);

FILL FILL_2__8720_ (
);

FILL FILL_2__8300_ (
);

NAND2X1 _6819_ (
    .A(Xin_5_bF$buf3),
    .B(gnd),
    .Y(_416_)
);

FILL FILL_2__12966_ (
);

FILL FILL_2__12546_ (
);

FILL FILL_2__12126_ (
);

FILL FILL_0__13160_ (
);

FILL FILL_1__11959_ (
);

FILL FILL_1__11539_ (
);

FILL FILL_1__11119_ (
);

FILL FILL_0__8546_ (
);

INVX1 _10817_ (
    .A(_4018_),
    .Y(_4019_)
);

FILL FILL_1__12900_ (
);

NOR2X1 _13289_ (
    .A(\u_fir_pe7.rYin [11]),
    .B(\u_fir_pe7.mul [11]),
    .Y(_6313_)
);

FILL FILL_2__9925_ (
);

FILL FILL_2__9505_ (
);

FILL FILL_1__7922_ (
);

FILL FILL_1__7502_ (
);

FILL FILL_3__7848_ (
);

FILL FILL_3__7008_ (
);

AOI21X1 _6992_ (
    .A(_557_),
    .B(_559_),
    .C(_585_),
    .Y(_586_)
);

NAND3X1 _6572_ (
    .A(_167_),
    .B(_152_),
    .C(_171_),
    .Y(_172_)
);

FILL FILL_3__10678_ (
);

FILL FILL_1__11292_ (
);

OAI21X1 _10990_ (
    .A(_4114_),
    .B(_4112_),
    .C(_4105_),
    .Y(_4190_)
);

INVX1 _10570_ (
    .A(\u_fir_pe4.mul [3]),
    .Y(_3837_)
);

FILL FILL_0__10285_ (
);

NAND2X1 _10150_ (
    .A(gnd),
    .B(\X[4] [4]),
    .Y(_3429_)
);

FILL FILL_1__8707_ (
);

FILL FILL_2__10612_ (
);

INVX1 _7777_ (
    .A(_1257_),
    .Y(_1293_)
);

NAND3X1 _7357_ (
    .A(_867_),
    .B(_875_),
    .C(_877_),
    .Y(_878_)
);

FILL FILL_2__13084_ (
);

FILL FILL_0__6612_ (
);

FILL FILL_1__12077_ (
);

FILL FILL_0__9084_ (
);

NAND3X1 _11775_ (
    .A(_4883_),
    .B(_4887_),
    .C(_4889_),
    .Y(_4896_)
);

FILL FILL_3__7181_ (
);

INVX1 _11355_ (
    .A(_4511_),
    .Y(_4549_)
);

FILL FILL_3__12824_ (
);

FILL FILL_3__12404_ (
);

FILL FILL_2__11817_ (
);

FILL FILL_0__12851_ (
);

FILL FILL_0__12431_ (
);

FILL FILL_0__12011_ (
);

FILL FILL_1__7099_ (
);

FILL FILL_0__7817_ (
);

NAND2X1 _9923_ (
    .A(_3202_),
    .B(_3205_),
    .Y(_3206_)
);

NAND2X1 _9503_ (
    .A(gnd),
    .B(_2789_),
    .Y(_2859_)
);

FILL FILL_1__8880_ (
);

FILL FILL_1__8460_ (
);

FILL FILL_1__8040_ (
);

FILL FILL_0__13216_ (
);

FILL FILL_2__6383_ (
);

FILL FILL_1__9665_ (
);

FILL FILL_1__9245_ (
);

FILL FILL_2__11990_ (
);

FILL FILL_2__11570_ (
);

FILL FILL_2__11150_ (
);

FILL FILL_1__10983_ (
);

FILL FILL_1__10563_ (
);

FILL FILL_1__10143_ (
);

FILL FILL_0__7990_ (
);

FILL FILL_2__7588_ (
);

FILL FILL_0__7570_ (
);

FILL FILL_2__7168_ (
);

FILL FILL_0__7150_ (
);

AND2X2 _6628_ (
    .A(Xin[3]),
    .B(gnd),
    .Y(_227_)
);

FILL FILL_2__12775_ (
);

FILL FILL_2__12355_ (
);

FILL FILL_1__11768_ (
);

FILL FILL_1__11348_ (
);

FILL FILL_0__8775_ (
);

FILL FILL_0__8355_ (
);

FILL FILL_3__6452_ (
);

NAND3X1 _10626_ (
    .A(_3889_),
    .B(_3886_),
    .C(_3849_),
    .Y(_3890_)
);

AOI21X1 _10206_ (
    .A(_3395_),
    .B(_3473_),
    .C(_3481_),
    .Y(_3484_)
);

NAND3X1 _13098_ (
    .A(_6090_),
    .B(_6132_),
    .C(_6091_),
    .Y(_6133_)
);

FILL FILL_2__9734_ (
);

FILL FILL_2__9314_ (
);

FILL FILL_0__11702_ (
);

FILL FILL_1__7731_ (
);

FILL FILL_1__7311_ (
);

NOR2X1 _6381_ (
    .A(_689_),
    .B(_710_),
    .Y(_720_)
);

FILL FILL_0__12907_ (
);

FILL FILL_3__10487_ (
);

FILL FILL_3__10067_ (
);

FILL FILL_0__10094_ (
);

FILL FILL_1__8936_ (
);

FILL FILL_1__8516_ (
);

FILL FILL_2__10841_ (
);

FILL FILL_2__10421_ (
);

FILL FILL_2__10001_ (
);

OAI21X1 _7586_ (
    .A(_1022_),
    .B(_1027_),
    .C(_1026_),
    .Y(_1104_)
);

OAI21X1 _7166_ (
    .A(_742_),
    .B(_743_),
    .C(_747_),
    .Y(_749_)
);

FILL FILL_3__9803_ (
);

FILL FILL_2__6859_ (
);

FILL FILL_0__6841_ (
);

FILL FILL_0__6421_ (
);

FILL FILL_2__6439_ (
);

DFFPOSX1 _11584_ (
    .D(_4774_[0]),
    .CLK(clk_bF$buf40),
    .Q(\Y[6] [0])
);

FILL FILL_0__11299_ (
);

AND2X2 _11164_ (
    .A(_4352_),
    .B(_4357_),
    .Y(_4362_)
);

FILL FILL_2__7800_ (
);

FILL FILL_0__12660_ (
);

FILL FILL_2__11206_ (
);

FILL FILL_0__12240_ (
);

FILL FILL_1__10619_ (
);

FILL FILL_0__7626_ (
);

NOR2X1 _9732_ (
    .A(\u_fir_pe3.rYin [7]),
    .B(\u_fir_pe3.mul [7]),
    .Y(_3075_)
);

AOI21X1 _9312_ (
    .A(_2670_),
    .B(_2665_),
    .C(_2526_),
    .Y(_2671_)
);

INVX1 _12789_ (
    .A(_5827_),
    .Y(_5828_)
);

FILL FILL_3__8195_ (
);

INVX1 _12369_ (
    .A(\u_fir_pe6.rYin [8]),
    .Y(_5472_)
);

FILL FILL_0__13025_ (
);

NOR2X1 _13310_ (
    .A(_6333_),
    .B(_6332_),
    .Y(_6334_)
);

FILL FILL_3__6928_ (
);

FILL FILL_3__6508_ (
);

FILL FILL_1__9894_ (
);

FILL FILL_1__9474_ (
);

FILL FILL_1__9054_ (
);

FILL FILL_1__10792_ (
);

FILL FILL_1__10372_ (
);

FILL FILL_2__7397_ (
);

FILL FILL_3__13171_ (
);

NAND2X1 _6857_ (
    .A(_442_),
    .B(_449_),
    .Y(_453_)
);

INVX1 _6437_ (
    .A(_38_),
    .Y(_39_)
);

FILL FILL_2__12584_ (
);

FILL FILL_2__12164_ (
);

FILL FILL_1__11997_ (
);

FILL FILL_1__11577_ (
);

FILL FILL_1__11157_ (
);

FILL FILL_0__8584_ (
);

FILL FILL_3__6681_ (
);

FILL FILL_0__8164_ (
);

INVX1 _10855_ (
    .A(_4055_),
    .Y(_4056_)
);

OAI21X1 _10435_ (
    .A(_3262_),
    .B(_3493_),
    .C(_3667_),
    .Y(_3710_)
);

AOI21X1 _10015_ (
    .A(_3291_),
    .B(_3292_),
    .C(_3290_),
    .Y(_3296_)
);

FILL FILL_3__11904_ (
);

FILL FILL_2__9963_ (
);

FILL FILL_0__11931_ (
);

FILL FILL_2__9543_ (
);

FILL FILL_2__9123_ (
);

FILL FILL_0__11511_ (
);

FILL FILL_1__6599_ (
);

FILL FILL_1__7960_ (
);

FILL FILL_1__7540_ (
);

FILL FILL_1__7120_ (
);

FILL FILL_0__9789_ (
);

FILL FILL_0__9369_ (
);

FILL FILL_3__7466_ (
);

FILL FILL_3__7046_ (
);

FILL FILL_1__13303_ (
);

FILL FILL_0__12716_ (
);

FILL FILL_3__10296_ (
);

FILL FILL_1__8745_ (
);

FILL FILL_1__8325_ (
);

FILL FILL_2__10650_ (
);

FILL FILL_2__10230_ (
);

NAND3X1 _7395_ (
    .A(_851_),
    .B(_914_),
    .C(_915_),
    .Y(_916_)
);

FILL FILL254550x57750 (
);

FILL FILL_0__6650_ (
);

FILL FILL_2__6668_ (
);

NAND2X1 _11393_ (
    .A(_4584_),
    .B(_4585_),
    .Y(_4586_)
);

FILL FILL_3__12862_ (
);

FILL FILL_3__12022_ (
);

FILL FILL_2__11855_ (
);

FILL FILL_2__11435_ (
);

FILL FILL_2__11015_ (
);

FILL FILL_1__10848_ (
);

FILL FILL_1__10428_ (
);

FILL FILL_1__10008_ (
);

FILL FILL_0__7855_ (
);

NAND2X1 _9961_ (
    .A(_3197_),
    .B(_3202_),
    .Y(_3243_)
);

FILL FILL_0__7435_ (
);

INVX1 _9541_ (
    .A(_2896_),
    .Y(_2897_)
);

FILL FILL_0__7015_ (
);

NAND3X1 _9121_ (
    .A(_2477_),
    .B(_2481_),
    .C(_2479_),
    .Y(_2482_)
);

NAND3X1 _12598_ (
    .A(_5607_),
    .B(_5624_),
    .C(_5627_),
    .Y(_5640_)
);

NAND3X1 _12178_ (
    .A(_5277_),
    .B(_5283_),
    .C(_5241_),
    .Y(_5293_)
);

FILL FILL_2__8814_ (
);

FILL FILL_0__13254_ (
);

FILL FILL_1__6811_ (
);

FILL FILL_1__9283_ (
);

FILL FILL253950x115350 (
);

FILL FILL_1__10181_ (
);

AOI21X1 _6666_ (
    .A(_152_),
    .B(_171_),
    .C(_264_),
    .Y(_265_)
);

FILL FILL_2__12393_ (
);

FILL FILL_1__11386_ (
);

FILL FILL_0__8393_ (
);

FILL FILL_0__10799_ (
);

FILL FILL_0__10379_ (
);

NAND2X1 _10664_ (
    .A(_3923_),
    .B(_3916_),
    .Y(_3927_)
);

NAND2X1 _10244_ (
    .A(_3513_),
    .B(_3521_),
    .Y(_3522_)
);

FILL FILL_2__9772_ (
);

FILL FILL_2__10706_ (
);

FILL FILL_2__9352_ (
);

FILL FILL_0__11740_ (
);

FILL FILL_0__11320_ (
);

FILL FILL_2__13178_ (
);

FILL FILL_0__6706_ (
);

NAND2X1 _8812_ (
    .A(_2239_),
    .B(_2238_),
    .Y(_2240_)
);

FILL FILL_0__9598_ (
);

FILL FILL_3__7695_ (
);

FILL FILL_0__9178_ (
);

NOR2X1 _11869_ (
    .A(_4986_),
    .B(_4988_),
    .Y(_5578_[6])
);

NOR2X1 _11449_ (
    .A(\u_fir_pe5.rYin [3]),
    .B(\u_fir_pe5.mul [3]),
    .Y(_4636_)
);

NAND2X1 _11029_ (
    .A(_4226_),
    .B(_4227_),
    .Y(_4228_)
);

FILL FILL_3__12918_ (
);

FILL FILL_1__13112_ (
);

FILL FILL_0__12945_ (
);

AND2X2 _12810_ (
    .A(_5800_),
    .B(_5797_),
    .Y(_5849_)
);

FILL FILL_0__12525_ (
);

FILL FILL_0__12105_ (
);

FILL FILL_1__8554_ (
);

FILL FILL_1__8134_ (
);

FILL FILL_3__9421_ (
);

FILL FILL_2__6897_ (
);

FILL FILL_2__6477_ (
);

FILL FILL_1__9759_ (
);

FILL FILL_1__9339_ (
);

FILL FILL_3__12251_ (
);

FILL FILL_2__11664_ (
);

FILL FILL_2__11244_ (
);

FILL FILL_1__10657_ (
);

FILL FILL_1__10237_ (
);

FILL FILL_0__7664_ (
);

INVX1 _9770_ (
    .A(_3113_),
    .Y(_3114_)
);

OAI21X1 _9350_ (
    .A(_2629_),
    .B(_2707_),
    .C(_2651_),
    .Y(_2708_)
);

FILL FILL_2__8623_ (
);

FILL FILL_2__8203_ (
);

FILL FILL_3__13036_ (
);

FILL FILL_2__12869_ (
);

FILL FILL_2__12449_ (
);

FILL FILL_2__12029_ (
);

FILL FILL_0__13063_ (
);

FILL FILL_1__6620_ (
);

FILL FILL_0__8869_ (
);

FILL FILL_0__8449_ (
);

FILL FILL_3__6546_ (
);

FILL FILL_0__8029_ (
);

FILL FILL_1__9092_ (
);

FILL FILL_1__12803_ (
);

FILL FILL_2__9828_ (
);

FILL FILL_0__9810_ (
);

FILL FILL_2__9408_ (
);

FILL FILL_1__7825_ (
);

FILL FILL_1__7405_ (
);

NAND3X1 _6895_ (
    .A(_488_),
    .B(_490_),
    .C(_489_),
    .Y(_491_)
);

OAI21X1 _6475_ (
    .A(_778_),
    .B(_74_),
    .C(_75_),
    .Y(_76_)
);

FILL FILL_1__11195_ (
);

AOI21X1 _10893_ (
    .A(_4085_),
    .B(_4081_),
    .C(_4067_),
    .Y(_4094_)
);

AOI21X1 _10473_ (
    .A(_3744_),
    .B(_3645_),
    .C(_3746_),
    .Y(_3747_)
);

FILL FILL_0__10188_ (
);

NAND2X1 _10053_ (
    .A(\X[4] [2]),
    .B(gnd),
    .Y(_3333_)
);

FILL FILL_2__10935_ (
);

FILL FILL_2__9581_ (
);

FILL FILL_2__10515_ (
);

FILL FILL_2__9161_ (
);

FILL FILL_0__6935_ (
);

FILL FILL_0__6515_ (
);

NOR3X1 _8621_ (
    .A(_1899_),
    .B(_1726_),
    .C(_1915_),
    .Y(_2057_)
);

NAND3X1 _8201_ (
    .A(_1623_),
    .B(_1639_),
    .C(_1642_),
    .Y(_1643_)
);

NAND2X1 _11678_ (
    .A(_5563_),
    .B(_4800_),
    .Y(_4801_)
);

NAND3X1 _11258_ (
    .A(_4452_),
    .B(_4449_),
    .C(_4453_),
    .Y(_4454_)
);

FILL FILL_0__12754_ (
);

FILL FILL_0__12334_ (
);

AOI21X1 _9826_ (
    .A(\X[3] [0]),
    .B(vdd),
    .C(_3091_),
    .Y(_3168_)
);

NAND2X1 _9406_ (
    .A(_2763_),
    .B(_2758_),
    .Y(_2764_)
);

FILL FILL_1__8783_ (
);

FILL FILL_1__8363_ (
);

FILL FILL253050x198150 (
);

FILL FILL_3__9650_ (
);

FILL FILL_0__13119_ (
);

BUFX2 _13404_ (
    .A(_6377_[10]),
    .Y(Yout[10])
);

FILL FILL_1__9988_ (
);

FILL FILL_1__9568_ (
);

FILL FILL_1__9148_ (
);

FILL FILL_2__11893_ (
);

FILL FILL_2__11473_ (
);

FILL FILL_2__11053_ (
);

FILL FILL_1__10886_ (
);

FILL FILL_1__10466_ (
);

FILL FILL_1__10046_ (
);

FILL FILL_0__7893_ (
);

FILL FILL_0__7473_ (
);

FILL FILL_0__7053_ (
);

FILL FILL_2__8852_ (
);

FILL FILL_2__8432_ (
);

FILL FILL_0__10820_ (
);

FILL FILL_3__13265_ (
);

FILL FILL_0__10400_ (
);

FILL FILL_2__8012_ (
);

FILL FILL_2__12678_ (
);

FILL FILL_2__12258_ (
);

FILL FILL_0__13292_ (
);

FILL FILL_0__8678_ (
);

FILL FILL_3__6775_ (
);

FILL FILL_0__8258_ (
);

NAND2X1 _10949_ (
    .A(gnd),
    .B(\X[5] [4]),
    .Y(_4149_)
);

NAND2X1 _10529_ (
    .A(_3801_),
    .B(_3798_),
    .Y(_3984_[13])
);

OAI21X1 _10109_ (
    .A(_3387_),
    .B(_3388_),
    .C(_3386_),
    .Y(_3389_)
);

FILL FILL_1__12612_ (
);

FILL FILL_2__9637_ (
);

FILL FILL_2__9217_ (
);

FILL FILL_1__7634_ (
);

FILL FILL_3__8921_ (
);

NAND3X1 _10282_ (
    .A(_3557_),
    .B(_3558_),
    .C(_3559_),
    .Y(_3560_)
);

FILL FILL_1__8839_ (
);

FILL FILL_3__11751_ (
);

FILL FILL_1__8419_ (
);

FILL FILL_3__11331_ (
);

FILL FILL_2__9390_ (
);

FILL FILL_2__10324_ (
);

INVX1 _7489_ (
    .A(_1007_),
    .Y(_1008_)
);

INVX1 _7069_ (
    .A(\u_fir_pe0.rYin [4]),
    .Y(_655_)
);

FILL FILL_0__6744_ (
);

AND2X2 _8850_ (
    .A(_2273_),
    .B(_2272_),
    .Y(_2384_[6])
);

INVX1 _8430_ (
    .A(_1771_),
    .Y(_1869_)
);

OAI21X1 _8010_ (
    .A(_1509_),
    .B(_1510_),
    .C(_1508_),
    .Y(_1514_)
);

OAI21X1 _11487_ (
    .A(_4668_),
    .B(_4669_),
    .C(_4665_),
    .Y(_4670_)
);

INVX1 _11067_ (
    .A(_4120_),
    .Y(_4266_)
);

FILL FILL_3__12956_ (
);

FILL FILL_2__7703_ (
);

FILL FILL_3__12536_ (
);

FILL FILL_3__12116_ (
);

FILL FILL_1__13150_ (
);

FILL FILL_2__11949_ (
);

FILL FILL_0__12983_ (
);

FILL FILL_2__11529_ (
);

FILL FILL_0__12563_ (
);

FILL FILL_2__11109_ (
);

FILL FILL_0__12143_ (
);

FILL FILL_0__7949_ (
);

FILL FILL_0__7529_ (
);

OAI22X1 _9635_ (
    .A(_2535_),
    .B(_2853_),
    .C(_2696_),
    .D(_2626_),
    .Y(_2988_)
);

FILL FILL_0__7109_ (
);

AND2X2 _9215_ (
    .A(_2525_),
    .B(_2526_),
    .Y(_2575_)
);

FILL FILL_1__8592_ (
);

FILL FILL_1__8172_ (
);

FILL FILL_2__8908_ (
);

INVX1 _13213_ (
    .A(_6229_),
    .Y(_6239_)
);

FILL FILL_1__6905_ (
);

FILL FILL_1__9797_ (
);

FILL FILL_1__9377_ (
);

FILL FILL_2__11282_ (
);

FILL FILL_1__10695_ (
);

FILL FILL_1__10275_ (
);

FILL FILL_0__7282_ (
);

FILL FILL_3__10602_ (
);

FILL FILL_2__8661_ (
);

FILL FILL_2__8241_ (
);

FILL FILL_2__12067_ (
);

NAND2X1 _7701_ (
    .A(_1203_),
    .B(_1206_),
    .Y(_1218_)
);

FILL FILL_0__8487_ (
);

DFFPOSX1 _10758_ (
    .D(_3984_[11]),
    .CLK(clk_bF$buf7),
    .Q(\u_fir_pe4.mul [11])
);

FILL FILL_0__8067_ (
);

NAND2X1 _10338_ (
    .A(_3579_),
    .B(_3582_),
    .Y(_3615_)
);

FILL FILL_1__12841_ (
);

FILL FILL_1__12421_ (
);

FILL FILL_1__12001_ (
);

FILL FILL_2__9446_ (
);

FILL FILL_0__11834_ (
);

FILL FILL_2__9026_ (
);

FILL FILL_0__11414_ (
);

NOR2X1 _8906_ (
    .A(_2329_),
    .B(_2326_),
    .Y(_2330_)
);

FILL FILL_1__7863_ (
);

FILL FILL_1__7443_ (
);

FILL FILL_1__7023_ (
);

FILL FILL_3__7789_ (
);

FILL FILL_1__13206_ (
);

AOI21X1 _12904_ (
    .A(_5936_),
    .B(_5941_),
    .C(_5880_),
    .Y(_5942_)
);

FILL FILL_0__12619_ (
);

FILL FILL_3__8310_ (
);

NAND3X1 _10091_ (
    .A(_3324_),
    .B(_3365_),
    .C(_3370_),
    .Y(_3371_)
);

FILL FILL_3__11980_ (
);

FILL FILL_1__8648_ (
);

FILL FILL_1__8228_ (
);

FILL FILL_3__11560_ (
);

FILL FILL_2__10973_ (
);

FILL FILL_2__10553_ (
);

FILL FILL_2__10133_ (
);

NOR2X1 _7298_ (
    .A(_820_),
    .B(_819_),
    .Y(_1591_[3])
);

FILL FILL_3__9935_ (
);

FILL FILL_3__9515_ (
);

FILL FILL_0__6973_ (
);

FILL FILL_0__6553_ (
);

AOI21X1 _11296_ (
    .A(_4440_),
    .B(_4443_),
    .C(_4491_),
    .Y(_4492_)
);

FILL FILL_2__7932_ (
);

FILL FILL_3__12765_ (
);

FILL FILL_2__7512_ (
);

FILL FILL_3__12345_ (
);

FILL FILL_2__11758_ (
);

FILL FILL_0__12792_ (
);

FILL FILL_2__11338_ (
);

FILL FILL_0__12372_ (
);

FILL FILL_0__7758_ (
);

DFFPOSX1 _9864_ (
    .D(\Y[3] [10]),
    .CLK(clk_bF$buf17),
    .Q(\u_fir_pe3.rYin [10])
);

FILL FILL_0__7338_ (
);

NAND2X1 _9444_ (
    .A(gnd),
    .B(\X[3] [7]),
    .Y(_2801_)
);

NAND2X1 _9024_ (
    .A(_3111_),
    .B(_3175_),
    .Y(_3176_)
);

FILL FILL_2__8717_ (
);

FILL FILL_0__13157_ (
);

NAND2X1 _13022_ (
    .A(_6056_),
    .B(_6057_),
    .Y(_6058_)
);

FILL FILL_1__6714_ (
);

FILL FILL_1__9186_ (
);

FILL FILL_0__9904_ (
);

FILL FILL_2__11091_ (
);

FILL FILL_1__10084_ (
);

FILL FILL_0__7091_ (
);

FILL FILL_1__7919_ (
);

FILL FILL_3__10831_ (
);

FILL FILL_2__8890_ (
);

FILL FILL_2__8470_ (
);

FILL FILL_2__8050_ (
);

OR2X2 _6989_ (
    .A(_581_),
    .B(_579_),
    .Y(_583_)
);

AOI21X1 _6569_ (
    .A(_163_),
    .B(_165_),
    .C(_156_),
    .Y(_169_)
);

FILL FILL_2__12296_ (
);

AND2X2 _7930_ (
    .A(\u_fir_pe1.rYin [2]),
    .B(\u_fir_pe1.mul [2]),
    .Y(_1438_)
);

NAND3X1 _7510_ (
    .A(_1023_),
    .B(_1028_),
    .C(_1026_),
    .Y(_1029_)
);

FILL FILL_1__11289_ (
);

FILL FILL_0__8296_ (
);

NAND3X1 _10987_ (
    .A(_4180_),
    .B(_4181_),
    .C(_4186_),
    .Y(_4187_)
);

FILL FILL_3__6393_ (
);

NAND2X1 _10567_ (
    .A(_3831_),
    .B(_3834_),
    .Y(_3978_[2])
);

NAND2X1 _10147_ (
    .A(_3420_),
    .B(_3425_),
    .Y(_3426_)
);

FILL FILL_1__12650_ (
);

FILL FILL_1__12230_ (
);

FILL FILL_2__9675_ (
);

FILL FILL_2__10609_ (
);

FILL FILL_2__9255_ (
);

FILL FILL_0__11643_ (
);

FILL FILL_0__11223_ (
);

FILL FILL_0__6609_ (
);

NAND2X1 _8715_ (
    .A(_2148_),
    .B(_2149_),
    .Y(_2390_[11])
);

FILL FILL_1__7672_ (
);

FILL FILL_1__13015_ (
);

FILL FILL_0__12848_ (
);

OAI21X1 _12713_ (
    .A(_5748_),
    .B(_5749_),
    .C(_5734_),
    .Y(_5753_)
);

FILL FILL_0__12428_ (
);

FILL FILL_0__12008_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1__8877_ (
);

FILL FILL_1__8457_ (
);

FILL FILL_1__8037_ (
);

FILL FILL_2__10782_ (
);

FILL FILL_2__10362_ (
);

FILL FILL_3__9744_ (
);

FILL FILL_0__6782_ (
);

FILL FILL_2__7741_ (
);

FILL FILL_3__12574_ (
);

FILL FILL_2__7321_ (
);

FILL FILL_2__11987_ (
);

FILL FILL_2__11567_ (
);

FILL FILL_2__11147_ (
);

FILL FILL_0__12181_ (
);

FILL FILL_0__7987_ (
);

FILL FILL_0__7567_ (
);

AND2X2 _9673_ (
    .A(\u_fir_pe3.rYin [0]),
    .B(\u_fir_pe3.mul [0]),
    .Y(_3022_)
);

FILL FILL_0__7147_ (
);

OAI21X1 _9253_ (
    .A(_2610_),
    .B(_2611_),
    .C(_2601_),
    .Y(_2612_)
);

FILL FILL_1__11921_ (
);

FILL FILL_1__11501_ (
);

FILL FILL_2__8946_ (
);

FILL FILL_2__8526_ (
);

FILL FILL_0__10914_ (
);

OAI21X1 _13251_ (
    .A(_6244_),
    .B(_6245_),
    .C(_6273_),
    .Y(_6274_)
);

FILL FILL_1__6943_ (
);

FILL FILL_1__6523_ (
);

FILL FILL_3__6869_ (
);

FILL FILL_3__6449_ (
);

FILL FILL_1__12706_ (
);

FILL FILL_0__9713_ (
);

FILL FILL_1__7728_ (
);

FILL FILL_1__7308_ (
);

FILL FILL_3__10220_ (
);

AND2X2 _6798_ (
    .A(_394_),
    .B(_391_),
    .Y(_395_)
);

NAND2X1 _6378_ (
    .A(Xin[0]),
    .B(gnd),
    .Y(_689_)
);

FILL FILL_1__11098_ (
);

NAND3X1 _10796_ (
    .A(_4773_),
    .B(_3998_),
    .C(_3994_),
    .Y(_3999_)
);

OAI22X1 _10376_ (
    .A(_3605_),
    .B(_3493_),
    .C(_3213_),
    .D(_3604_),
    .Y(_3652_)
);

FILL FILL_3__11845_ (
);

FILL FILL_3__11425_ (
);

FILL FILL_3__11005_ (
);

FILL FILL_2__10838_ (
);

FILL FILL_2__9484_ (
);

FILL FILL_0__11872_ (
);

FILL FILL_2__10418_ (
);

FILL FILL_2__9064_ (
);

FILL FILL_0__11452_ (
);

FILL FILL_0__11032_ (
);

FILL FILL_0__6838_ (
);

NAND3X1 _8944_ (
    .A(_2361_),
    .B(_2367_),
    .C(_2362_),
    .Y(_2368_)
);

FILL FILL_0__6418_ (
);

AOI21X1 _8524_ (
    .A(_1872_),
    .B(_1871_),
    .C(_1803_),
    .Y(_1962_)
);

DFFPOSX1 _8104_ (
    .D(\Y[1] [4]),
    .CLK(clk_bF$buf52),
    .Q(\u_fir_pe1.rYin [4])
);

FILL FILL_1__7481_ (
);

FILL FILL_1__7061_ (
);

FILL FILL_1__13244_ (
);

NOR2X1 _12942_ (
    .A(_5977_),
    .B(_5978_),
    .Y(_5979_)
);

FILL FILL_0__12657_ (
);

FILL FILL_0__12237_ (
);

NOR2X1 _12522_ (
    .A(_6268_),
    .B(_6310_),
    .Y(_6319_)
);

NAND3X1 _12102_ (
    .A(_5165_),
    .B(_5213_),
    .C(_5218_),
    .Y(_5219_)
);

INVX1 _9729_ (
    .A(\u_fir_pe3.rYin [7]),
    .Y(_3072_)
);

NAND3X1 _9309_ (
    .A(_2662_),
    .B(_2661_),
    .C(_2663_),
    .Y(_2668_)
);

FILL FILL_1__8686_ (
);

FILL FILL_1__8266_ (
);

FILL FILL_2__10591_ (
);

FILL FILL_2__10171_ (
);

FILL FILL_3__9133_ (
);

INVX1 _13307_ (
    .A(\u_fir_pe7.mul [13]),
    .Y(_6331_)
);

FILL FILL_0__6591_ (
);

FILL FILL_2__7970_ (
);

FILL FILL_2__7550_ (
);

FILL FILL_2__7130_ (
);

FILL FILL_2__11796_ (
);

FILL FILL_2__11376_ (
);

FILL FILL_1__10789_ (
);

FILL FILL_1__10369_ (
);

FILL FILL_0__7796_ (
);

FILL FILL_0__7376_ (
);

AOI21X1 _9482_ (
    .A(_2827_),
    .B(_2822_),
    .C(_2774_),
    .Y(_2839_)
);

NAND2X1 _9062_ (
    .A(vdd),
    .B(\X[3] [3]),
    .Y(_2424_)
);

FILL FILL_1__11730_ (
);

FILL FILL_1__11310_ (
);

FILL FILL_2__8755_ (
);

FILL FILL_2__8335_ (
);

FILL FILL_0__10303_ (
);

FILL FILL_0__13195_ (
);

NAND2X1 _13060_ (
    .A(_6063_),
    .B(_6066_),
    .Y(_6095_)
);

FILL FILL_1__6752_ (
);

FILL FILL_2__13102_ (
);

FILL FILL_1__12935_ (
);

FILL FILL_0__9942_ (
);

FILL FILL_0__9522_ (
);

FILL FILL_0__11928_ (
);

FILL FILL_0__9102_ (
);

FILL FILL_0__11508_ (
);

FILL FILL_1__7957_ (
);

FILL FILL_1__7537_ (
);

FILL FILL_1__7117_ (
);

FILL FILL_3__8404_ (
);

AOI21X1 _10185_ (
    .A(_3372_),
    .B(_3370_),
    .C(_3463_),
    .Y(_3464_)
);

FILL FILL_2__6821_ (
);

FILL FILL_2__6401_ (
);

FILL FILL_3__11234_ (
);

FILL FILL_2__10647_ (
);

FILL FILL_2__9293_ (
);

FILL FILL_0__11681_ (
);

FILL FILL_2__10227_ (
);

FILL FILL_0__11261_ (
);

FILL FILL_0__6647_ (
);

INVX1 _8753_ (
    .A(_2160_),
    .Y(_2186_)
);

AOI21X1 _8333_ (
    .A(_1676_),
    .B(_1694_),
    .C(_1772_),
    .Y(_1773_)
);

FILL FILL_1__7290_ (
);

FILL FILL_3__12859_ (
);

FILL FILL_2__7606_ (
);

FILL FILL_3__12439_ (
);

FILL FILL_1__13053_ (
);

FILL FILL_0__12886_ (
);

INVX1 _12751_ (
    .A(_5789_),
    .Y(_5790_)
);

FILL FILL_0__12046_ (
);

INVX1 _12331_ (
    .A(\u_fir_pe6.rYin [4]),
    .Y(_5437_)
);

NAND3X1 _9958_ (
    .A(_3216_),
    .B(_3239_),
    .C(_3238_),
    .Y(_3240_)
);

NAND2X1 _9538_ (
    .A(_2886_),
    .B(_2892_),
    .Y(_2894_)
);

NAND2X1 _9118_ (
    .A(_2427_),
    .B(_2478_),
    .Y(_2479_)
);

FILL FILL_1__8495_ (
);

FILL FILL_1__8075_ (
);

FILL FILL_3__9362_ (
);

NAND2X1 _13116_ (
    .A(_6144_),
    .B(_6148_),
    .Y(_6150_)
);

FILL FILL_1__6808_ (
);

FILL FILL_3__12192_ (
);

FILL FILL_2__11185_ (
);

FILL FILL_1__10598_ (
);

FILL FILL_1__10178_ (
);

FILL FILL_0__7185_ (
);

AND2X2 _9291_ (
    .A(_2628_),
    .B(_2623_),
    .Y(_2650_)
);

FILL FILL_3__10925_ (
);

FILL FILL_2__8564_ (
);

FILL FILL_0__10952_ (
);

FILL FILL_2__8144_ (
);

FILL FILL_0__10532_ (
);

FILL FILL_0__10112_ (
);

NAND2X1 _7604_ (
    .A(vdd),
    .B(\X[1]_5_bF$buf3 ),
    .Y(_1122_)
);

FILL FILL_1__6981_ (
);

FILL FILL_1__6561_ (
);

FILL FILL_2__13331_ (
);

FILL FILL_3__6487_ (
);

FILL FILL_1__12744_ (
);

FILL FILL_1__12324_ (
);

FILL FILL_2__9769_ (
);

FILL FILL_0__9751_ (
);

FILL FILL_2__9349_ (
);

FILL FILL_0__9331_ (
);

FILL FILL_0__11737_ (
);

DFFPOSX1 _11602_ (
    .D(\X[5] [2]),
    .CLK(clk_bF$buf5),
    .Q(\X[6] [2])
);

FILL FILL_0__11317_ (
);

OAI21X1 _8809_ (
    .A(_2235_),
    .B(_2236_),
    .C(_2234_),
    .Y(_2237_)
);

FILL FILL_1__7766_ (
);

FILL FILL_1__7346_ (
);

FILL FILL_1__13109_ (
);

FILL FILL_3__8633_ (
);

NAND3X1 _12807_ (
    .A(_5817_),
    .B(_5836_),
    .C(_5830_),
    .Y(_5846_)
);

FILL FILL254250x216150 (
);

FILL FILL_2__6630_ (
);

FILL FILL_2__10876_ (
);

FILL FILL_2__10456_ (
);

FILL FILL_0__11490_ (
);

FILL FILL_2__10036_ (
);

FILL FILL_0__11070_ (
);

FILL FILL_1__9912_ (
);

FILL FILL_3__9418_ (
);

FILL FILL_0__6876_ (
);

DFFPOSX1 _8982_ (
    .D(\Y[2] [5]),
    .CLK(clk_bF$buf0),
    .Q(\u_fir_pe2.rYin [5])
);

FILL FILL_0__6456_ (
);

AND2X2 _8562_ (
    .A(vdd),
    .B(\X[2] [7]),
    .Y(_1999_)
);

NOR2X1 _8142_ (
    .A(_2364_),
    .B(_2372_),
    .Y(_2374_)
);

FILL FILL_1__10810_ (
);

NAND2X1 _11199_ (
    .A(_4386_),
    .B(_4395_),
    .Y(_4396_)
);

FILL FILL_2__7835_ (
);

FILL FILL_2__7415_ (
);

FILL FILL_1__13282_ (
);

INVX1 _12980_ (
    .A(_5962_),
    .Y(_6017_)
);

FILL FILL_0__12695_ (
);

FILL FILL_0__12275_ (
);

NOR2X1 _12560_ (
    .A(_5602_),
    .B(_5601_),
    .Y(_6373_[3])
);

NOR2X1 _12140_ (
    .A(_5255_),
    .B(_5198_),
    .Y(_5256_)
);

FILL FILL_2__12602_ (
);

AOI21X1 _9767_ (
    .A(_3105_),
    .B(_3083_),
    .C(_3103_),
    .Y(_3110_)
);

NAND3X1 _9347_ (
    .A(_2702_),
    .B(_2704_),
    .C(_2703_),
    .Y(_2705_)
);

FILL FILL254550x72150 (
);

FILL FILL_0__8602_ (
);

FILL FILL_3__9591_ (
);

DFFPOSX1 _13345_ (
    .D(_6369_[7]),
    .CLK(clk_bF$buf22),
    .Q(\Y[7] [7])
);

FILL FILL_1__6617_ (
);

FILL FILL_1__9089_ (
);

FILL FILL_0__9807_ (
);

FILL FILL_3__10314_ (
);

FILL FILL_2__8793_ (
);

FILL FILL_2__8373_ (
);

FILL FILL_0__10341_ (
);

FILL FILL_2__12199_ (
);

NAND3X1 _7833_ (
    .A(_1339_),
    .B(_1343_),
    .C(_1347_),
    .Y(_1348_)
);

NAND2X1 _7413_ (
    .A(_932_),
    .B(_931_),
    .Y(_933_)
);

FILL FILL_1__6790_ (
);

FILL FILL_2__13140_ (
);

FILL FILL_0__8199_ (
);

FILL FILL_3__11939_ (
);

FILL FILL_1__12973_ (
);

FILL FILL_1__12553_ (
);

FILL FILL_1__12133_ (
);

FILL FILL_0__9980_ (
);

FILL FILL_2__9998_ (
);

FILL FILL_2__9578_ (
);

FILL FILL_0__11966_ (
);

FILL FILL_0__9560_ (
);

FILL FILL_0__9140_ (
);

FILL FILL_2__9158_ (
);

AOI21X1 _11831_ (
    .A(_4945_),
    .B(_4947_),
    .C(_4938_),
    .Y(_4951_)
);

FILL FILL_0__11546_ (
);

AND2X2 _11411_ (
    .A(_4581_),
    .B(_4580_),
    .Y(_4603_)
);

FILL FILL_0__11126_ (
);

OAI21X1 _8618_ (
    .A(_1980_),
    .B(_1984_),
    .C(_1982_),
    .Y(_2054_)
);

FILL FILL_1__7995_ (
);

FILL FILL_1__7575_ (
);

FILL FILL_1__7155_ (
);

FILL FILL_3__8862_ (
);

NAND3X1 _12616_ (
    .A(gnd),
    .B(\X[6]_5_bF$buf3 ),
    .C(_5654_),
    .Y(_5657_)
);

FILL FILL_3__11692_ (
);

FILL FILL_3__11272_ (
);

FILL FILL_2__10685_ (
);

FILL FILL_2__10265_ (
);

FILL FILL254550x150 (
);

FILL FILL_1__9721_ (
);

FILL FILL_1__9301_ (
);

FILL FILL_0__6685_ (
);

NAND2X1 _8791_ (
    .A(_2222_),
    .B(_2216_),
    .Y(_2390_[14])
);

NAND2X1 _8371_ (
    .A(_1807_),
    .B(_1809_),
    .Y(_1810_)
);

FILL FILL_3__12897_ (
);

FILL FILL_2__7644_ (
);

FILL FILL_3__12057_ (
);

FILL FILL_1__13091_ (
);

FILL FILL_0__12084_ (
);

FILL FILL_2__12831_ (
);

FILL FILL_2__12411_ (
);

INVX1 _9996_ (
    .A(gnd),
    .Y(_3277_)
);

NAND2X1 _9576_ (
    .A(_2923_),
    .B(_2926_),
    .Y(_2931_)
);

NAND3X1 _9156_ (
    .A(_2511_),
    .B(_2516_),
    .C(_2458_),
    .Y(_2517_)
);

FILL FILL_1__11824_ (
);

FILL FILL_1__11404_ (
);

FILL FILL_2__8849_ (
);

FILL FILL_0__8831_ (
);

FILL FILL_0__8411_ (
);

FILL FILL_2__8429_ (
);

FILL FILL_0__10817_ (
);

FILL FILL_2__8009_ (
);

FILL FILL_0__13289_ (
);

NAND2X1 _13154_ (
    .A(_6185_),
    .B(_6186_),
    .Y(_6187_)
);

FILL FILL_1__6846_ (
);

FILL FILL_1__6426_ (
);

FILL FILL_1__12609_ (
);

FILL FILL_0__9616_ (
);

FILL FILL_3__7713_ (
);

FILL FILL_3__10543_ (
);

FILL FILL_0__10990_ (
);

FILL FILL_2__8182_ (
);

FILL FILL_0__10570_ (
);

FILL FILL_0__10150_ (
);

AOI21X1 _7642_ (
    .A(_1154_),
    .B(_1159_),
    .C(_1098_),
    .Y(_1160_)
);

DFFPOSX1 _7222_ (
    .D(Xin[7]),
    .CLK(clk_bF$buf34),
    .Q(\X[1] [7])
);

OAI21X1 _10699_ (
    .A(_3950_),
    .B(_3953_),
    .C(_3960_),
    .Y(_3963_)
);

OAI21X1 _10279_ (
    .A(_3323_),
    .B(_3556_),
    .C(_3470_),
    .Y(_3557_)
);

FILL FILL_2__6915_ (
);

FILL FILL_1__12782_ (
);

FILL FILL_3__11328_ (
);

FILL FILL_1__12362_ (
);

FILL FILL_2__9387_ (
);

FILL FILL_0__11775_ (
);

NAND2X1 _11640_ (
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_5471_)
);

FILL FILL_0__11355_ (
);

INVX1 _11220_ (
    .A(_4339_),
    .Y(_4417_)
);

NOR2X1 _8847_ (
    .A(_2270_),
    .B(_2269_),
    .Y(_2271_)
);

OAI21X1 _8427_ (
    .A(_1852_),
    .B(_1856_),
    .C(_1859_),
    .Y(_1866_)
);

NOR2X1 _8007_ (
    .A(_1510_),
    .B(_1509_),
    .Y(_1511_)
);

FILL FILL_1__7384_ (
);

FILL FILL_1__13147_ (
);

FILL FILL_3__8671_ (
);

NAND2X1 _12845_ (
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5883_)
);

FILL FILL_3__8251_ (
);

NAND2X1 _12425_ (
    .A(_5528_),
    .B(_5523_),
    .Y(_5529_)
);

AOI21X1 _12005_ (
    .A(_5118_),
    .B(_5122_),
    .C(_5104_),
    .Y(_5123_)
);

FILL FILL_1__8589_ (
);

FILL FILL_1__8169_ (
);

FILL FILL_2__10494_ (
);

FILL FILL_2__10074_ (
);

FILL FILL_1__9950_ (
);

FILL FILL_1__9530_ (
);

FILL FILL_1__9110_ (
);

FILL FILL_3__9456_ (
);

FILL FILL_3__9036_ (
);

FILL FILL_0__6494_ (
);

NOR2X1 _8180_ (
    .A(_1621_),
    .B(_1620_),
    .Y(_1622_)
);

FILL FILL_2__7873_ (
);

FILL FILL_2__7453_ (
);

FILL FILL_3__12286_ (
);

FILL FILL_2__7033_ (
);

FILL FILL_2__11699_ (
);

FILL FILL_2__11279_ (
);

OAI21X1 _6913_ (
    .A(_508_),
    .B(_376_),
    .C(_458_),
    .Y(_509_)
);

FILL FILL_2__12640_ (
);

FILL FILL_2__12220_ (
);

FILL FILL_0__7699_ (
);

FILL FILL_0__7279_ (
);

AOI21X1 _9385_ (
    .A(_2742_),
    .B(_2737_),
    .C(_2706_),
    .Y(_2743_)
);

FILL FILL_1__11213_ (
);

FILL FILL_2__8658_ (
);

FILL FILL_0__8640_ (
);

FILL FILL_2__8238_ (
);

FILL FILL_0__8220_ (
);

FILL FILL_0__10626_ (
);

INVX1 _10911_ (
    .A(_4052_),
    .Y(_4112_)
);

FILL FILL_0__10206_ (
);

FILL FILL_0__13098_ (
);

DFFPOSX1 _13383_ (
    .D(_6375_[5]),
    .CLK(clk_bF$buf48),
    .Q(\u_fir_pe7.mul [5])
);

FILL FILL_1__6655_ (
);

FILL FILL_2__13005_ (
);

FILL FILL_1__12838_ (
);

FILL FILL_1__12418_ (
);

FILL FILL_3__7942_ (
);

FILL FILL_0__9425_ (
);

FILL FILL_3__7102_ (
);

FILL FILL_3__10772_ (
);

FILL FILL_1__8801_ (
);

FILL FILL_3__8727_ (
);

OAI21X1 _7871_ (
    .A(_1173_),
    .B(_1384_),
    .C(_1356_),
    .Y(_1385_)
);

OAI21X1 _7451_ (
    .A(_966_),
    .B(_967_),
    .C(_952_),
    .Y(_971_)
);

INVX1 _7031_ (
    .A(_582_),
    .Y(_623_)
);

AOI21X1 _10088_ (
    .A(_3362_),
    .B(_3363_),
    .C(_3361_),
    .Y(_3368_)
);

FILL FILL_2__6724_ (
);

FILL FILL_1__12591_ (
);

FILL FILL_1__12171_ (
);

FILL FILL_2__9196_ (
);

FILL FILL_0__11164_ (
);

FILL FILL_2__11911_ (
);

AOI21X1 _8656_ (
    .A(_1989_),
    .B(_2019_),
    .C(_2022_),
    .Y(_2092_)
);

NAND2X1 _8236_ (
    .A(vdd),
    .B(\X[2] [2]),
    .Y(_1677_)
);

FILL FILL_1__7193_ (
);

FILL FILL_1__10904_ (
);

FILL FILL_0__7911_ (
);

FILL FILL_2__7929_ (
);

FILL FILL_2__7509_ (
);

FILL FILL_0__12789_ (
);

FILL FILL_3__8480_ (
);

NAND3X1 _12654_ (
    .A(_5632_),
    .B(_5690_),
    .C(_5694_),
    .Y(_5695_)
);

FILL FILL_0__12369_ (
);

FILL FILL_3__8060_ (
);

NOR2X1 _12234_ (
    .A(_5255_),
    .B(_5308_),
    .Y(_5348_)
);

FILL FILL_0__13310_ (
);

FILL FILL_1__8398_ (
);

FILL FILL_3__9685_ (
);

OAI22X1 _13019_ (
    .A(_5910_),
    .B(_5991_),
    .C(_6053_),
    .D(_6054_),
    .Y(_6055_)
);

FILL FILL_2__7682_ (
);

FILL FILL_2__7262_ (
);

FILL FILL_2__11088_ (
);

OAI21X1 _6722_ (
    .A(_15_),
    .B(_319_),
    .C(_25_),
    .Y(_320_)
);

FILL FILL_0__7088_ (
);

NAND3X1 _9194_ (
    .A(gnd),
    .B(\X[3] [4]),
    .C(_2544_),
    .Y(_2554_)
);

FILL FILL_3__10828_ (
);

FILL FILL_1__11862_ (
);

FILL FILL_3__10408_ (
);

FILL FILL_1__11442_ (
);

FILL FILL_1__11022_ (
);

FILL FILL_2__8887_ (
);

FILL FILL_2__8467_ (
);

FILL FILL_0__10855_ (
);

FILL FILL_0__10435_ (
);

DFFPOSX1 _10720_ (
    .D(_3978_[13]),
    .CLK(clk_bF$buf57),
    .Q(\Y[5] [13])
);

FILL FILL_2__8047_ (
);

INVX1 _10300_ (
    .A(_3576_),
    .Y(_3577_)
);

FILL FILL_0__10015_ (
);

AND2X2 _13192_ (
    .A(\u_fir_pe7.rYin [2]),
    .B(\u_fir_pe7.mul [2]),
    .Y(_6220_)
);

NOR2X1 _7927_ (
    .A(_1428_),
    .B(_1433_),
    .Y(_1436_)
);

NAND2X1 _7507_ (
    .A(_1024_),
    .B(_1025_),
    .Y(_1026_)
);

FILL FILL_1__6884_ (
);

FILL FILL_1__6464_ (
);

FILL FILL_2__13234_ (
);

FILL FILL_1__12647_ (
);

FILL FILL_1__12227_ (
);

FILL FILL_0__9654_ (
);

AOI21X1 _11925_ (
    .A(_5043_),
    .B(_5042_),
    .C(_5041_),
    .Y(_5044_)
);

FILL FILL_0__9234_ (
);

FILL FILL_3__7331_ (
);

OAI21X1 _11505_ (
    .A(_4677_),
    .B(_4678_),
    .C(_4688_),
    .Y(_4689_)
);

FILL FILL_1__7669_ (
);

FILL FILL_3__10161_ (
);

FILL FILL_1__8610_ (
);

NOR2X1 _7680_ (
    .A(_1195_),
    .B(_1196_),
    .Y(_1197_)
);

NOR2X1 _7260_ (
    .A(_1486_),
    .B(_1528_),
    .Y(_1537_)
);

FILL FILL_2__6953_ (
);

FILL FILL_3__11786_ (
);

FILL FILL_2__6533_ (
);

FILL FILL_3__11366_ (
);

FILL FILL_2__10779_ (
);

FILL FILL_2__10359_ (
);

FILL FILL_0__11393_ (
);

FILL FILL_1__9815_ (
);

FILL FILL_2__11720_ (
);

FILL FILL_2__11300_ (
);

FILL FILL_0__6779_ (
);

INVX1 _8885_ (
    .A(_2308_),
    .Y(_2309_)
);

AND2X2 _8465_ (
    .A(_1901_),
    .B(_1900_),
    .Y(_1903_)
);

INVX1 _8045_ (
    .A(\u_fir_pe1.mul [13]),
    .Y(_1549_)
);

FILL FILL_2__7738_ (
);

FILL FILL_0__7720_ (
);

FILL FILL_0__7300_ (
);

FILL FILL_2__7318_ (
);

FILL FILL_1__13185_ (
);

INVX1 _12883_ (
    .A(_5901_),
    .Y(_5921_)
);

FILL FILL_0__12598_ (
);

FILL FILL_0__12178_ (
);

DFFPOSX1 _12463_ (
    .D(_5572_[2]),
    .CLK(clk_bF$buf2),
    .Q(_6377_[2])
);

NAND2X1 _12043_ (
    .A(_5156_),
    .B(_5160_),
    .Y(_5578_[8])
);

FILL FILL_2__12925_ (
);

FILL FILL_1__11918_ (
);

FILL FILL_0__8925_ (
);

FILL FILL_0__8505_ (
);

FILL FILL_3__6602_ (
);

FILL FILL_3__9074_ (
);

NOR2X1 _13248_ (
    .A(_6269_),
    .B(_6270_),
    .Y(_6271_)
);

FILL FILL_2__7491_ (
);

FILL FILL_2__7071_ (
);

FILL FILL_3__7807_ (
);

NAND3X1 _6951_ (
    .A(_543_),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

AND2X2 _6531_ (
    .A(Xin[0]),
    .B(gnd),
    .Y(_131_)
);

FILL FILL_3__10637_ (
);

FILL FILL_1__11671_ (
);

FILL FILL_1__11251_ (
);

FILL FILL_2__8696_ (
);

FILL FILL_2__8276_ (
);

FILL FILL_0__10664_ (
);

FILL FILL_0__10244_ (
);

NAND2X1 _7736_ (
    .A(_1251_),
    .B(_1094_),
    .Y(_1252_)
);

NAND3X1 _7316_ (
    .A(vdd),
    .B(\X[1] [2]),
    .C(_828_),
    .Y(_838_)
);

FILL FILL_1__6693_ (
);

FILL FILL_2__13043_ (
);

FILL FILL_1__12876_ (
);

FILL FILL_1__12456_ (
);

FILL FILL_1__12036_ (
);

FILL FILL_0__9463_ (
);

FILL FILL_0__11869_ (
);

FILL FILL_3__7560_ (
);

FILL FILL_0__9043_ (
);

NAND2X1 _11734_ (
    .A(_5482_),
    .B(_4854_),
    .Y(_4855_)
);

FILL FILL_0__11449_ (
);

FILL FILL_3__7140_ (
);

FILL FILL_0__11029_ (
);

NAND2X1 _11314_ (
    .A(_4504_),
    .B(_4508_),
    .Y(_4509_)
);

FILL FILL_0__12810_ (
);

FILL FILL_1__7898_ (
);

FILL FILL_1__7478_ (
);

FILL FILL_3__10390_ (
);

FILL FILL_1__7058_ (
);

OAI21X1 _12939_ (
    .A(_5901_),
    .B(_5975_),
    .C(_5922_),
    .Y(_5976_)
);

FILL FILL_3__8345_ (
);

INVX1 _12519_ (
    .A(_6279_),
    .Y(_6289_)
);

FILL FILL_2__6762_ (
);

FILL FILL_3__11175_ (
);

FILL FILL_2__10588_ (
);

FILL FILL_2__10168_ (
);

FILL FILL_1__9624_ (
);

FILL FILL_1__9204_ (
);

FILL FILL_0__6588_ (
);

NAND3X1 _8694_ (
    .A(_2123_),
    .B(_2128_),
    .C(_2127_),
    .Y(_2129_)
);

INVX1 _8274_ (
    .A(_1614_),
    .Y(_1715_)
);

FILL FILL_1__10942_ (
);

FILL FILL_1__10522_ (
);

FILL FILL_1__10102_ (
);

FILL FILL_2__7967_ (
);

FILL FILL_2__7547_ (
);

FILL FILL_2__7127_ (
);

NAND2X1 _12692_ (
    .A(vdd),
    .B(\X[6] [3]),
    .Y(_5732_)
);

OR2X2 _12272_ (
    .A(_5383_),
    .B(_5376_),
    .Y(_5385_)
);

FILL FILL_2__12734_ (
);

FILL FILL_2__12314_ (
);

NOR2X1 _9899_ (
    .A(_3968_),
    .B(_3948_),
    .Y(_3971_)
);

OAI21X1 _9479_ (
    .A(_2826_),
    .B(_2825_),
    .C(_2776_),
    .Y(_2836_)
);

NAND2X1 _9059_ (
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2421_)
);

FILL FILL_1__11727_ (
);

FILL FILL_1__11307_ (
);

FILL FILL_0__8734_ (
);

FILL FILL_0__8314_ (
);

NOR2X1 _13057_ (
    .A(_6072_),
    .B(_6077_),
    .Y(_6092_)
);

FILL FILL_1__6749_ (
);

FILL FILL_0__9939_ (
);

FILL FILL_0__9519_ (
);

INVX1 _6760_ (
    .A(_271_),
    .Y(_358_)
);

FILL FILL_3__10866_ (
);

FILL FILL_1__11480_ (
);

FILL FILL_3__10026_ (
);

FILL FILL_1__11060_ (
);

FILL FILL_0__10893_ (
);

FILL FILL_0__10473_ (
);

FILL FILL_0__10053_ (
);

FILL FILL_2__10800_ (
);

OAI21X1 _7965_ (
    .A(_1462_),
    .B(_1463_),
    .C(_1467_),
    .Y(_1469_)
);

NAND3X1 _7545_ (
    .A(_1035_),
    .B(_1054_),
    .C(_1048_),
    .Y(_1064_)
);

INVX1 _7125_ (
    .A(_692_),
    .Y(_708_)
);

FILL FILL_2__13272_ (
);

FILL FILL_2__6818_ (
);

FILL FILL_0__6800_ (
);

FILL FILL_1__12685_ (
);

FILL FILL_1__12265_ (
);

FILL FILL_0__9692_ (
);

FILL FILL_0__9272_ (
);

AOI21X1 _11963_ (
    .A(_5063_),
    .B(_5065_),
    .C(_5080_),
    .Y(_5081_)
);

FILL FILL_0__11678_ (
);

INVX1 _11543_ (
    .A(\u_fir_pe5.rYin [12]),
    .Y(_4727_)
);

FILL FILL_0__11258_ (
);

OAI21X1 _11123_ (
    .A(_4320_),
    .B(_4314_),
    .C(_4308_),
    .Y(_4321_)
);

FILL FILL_1__7287_ (
);

FILL FILL_3__8574_ (
);

AOI21X1 _12748_ (
    .A(_5751_),
    .B(_5755_),
    .C(_5717_),
    .Y(_5787_)
);

NAND2X1 _12328_ (
    .A(_5434_),
    .B(_5429_),
    .Y(_5435_)
);

FILL FILL_0__13404_ (
);

FILL FILL_2__6991_ (
);

FILL FILL_2__6571_ (
);

FILL FILL_2__10397_ (
);

FILL FILL_1__9433_ (
);

FILL FILL_1__9013_ (
);

FILL FILL_3__9779_ (
);

FILL FILL_3__9359_ (
);

FILL FILL_0__6397_ (
);

DFFPOSX1 _8083_ (
    .D(_1587_[7]),
    .CLK(clk_bF$buf44),
    .Q(\Y[2] [7])
);

FILL FILL_1__10331_ (
);

FILL FILL_2__7776_ (
);

FILL FILL_2__7356_ (
);

NAND2X1 _12081_ (
    .A(\X[7]_5_bF$buf0 ),
    .B(gnd),
    .Y(_5198_)
);

FILL FILL_3__13130_ (
);

OAI21X1 _6816_ (
    .A(_333_),
    .B(_412_),
    .C(_411_),
    .Y(_413_)
);

FILL FILL_2__12963_ (
);

FILL FILL_2__12543_ (
);

FILL FILL_2__12123_ (
);

OAI21X1 _9288_ (
    .A(_2639_),
    .B(_2646_),
    .C(_2631_),
    .Y(_2647_)
);

FILL FILL_1__11956_ (
);

FILL FILL_1__11536_ (
);

FILL FILL_1__11116_ (
);

FILL FILL253950x201750 (
);

FILL FILL_0__8543_ (
);

FILL FILL_0__10949_ (
);

FILL FILL_3__6640_ (
);

FILL FILL_0__10529_ (
);

NAND2X1 _10814_ (
    .A(vdd),
    .B(\X[5] [1]),
    .Y(_4016_)
);

FILL FILL_0__10109_ (
);

AND2X2 _13286_ (
    .A(_6308_),
    .B(_6309_),
    .Y(_6369_[10])
);

FILL FILL_2__9922_ (
);

FILL FILL_2__9502_ (
);

FILL FILL_1__6978_ (
);

FILL FILL_1__6558_ (
);

FILL FILL_2__13328_ (
);

FILL FILL_0__9748_ (
);

FILL FILL_0__9328_ (
);

FILL FILL_3__7425_ (
);

FILL FILL_3__10255_ (
);

FILL FILL_0__10282_ (
);

FILL FILL_1__8704_ (
);

NAND2X1 _7774_ (
    .A(_1288_),
    .B(_1284_),
    .Y(_1290_)
);

NAND3X1 _7354_ (
    .A(gnd),
    .B(\X[1]_5_bF$buf0 ),
    .C(_872_),
    .Y(_875_)
);

FILL FILL_2__13081_ (
);

FILL FILL_2__6627_ (
);

FILL FILL_1__12074_ (
);

FILL FILL_2__9099_ (
);

FILL FILL_0__9081_ (
);

NAND3X1 _11772_ (
    .A(_4808_),
    .B(_4888_),
    .C(_4892_),
    .Y(_4893_)
);

FILL FILL_0__11487_ (
);

FILL FILL_0__11067_ (
);

OAI21X1 _11352_ (
    .A(_4290_),
    .B(_4464_),
    .C(_4508_),
    .Y(_4546_)
);

FILL FILL_1__9909_ (
);

FILL FILL_2__11814_ (
);

DFFPOSX1 _8979_ (
    .D(\Y[2] [2]),
    .CLK(clk_bF$buf12),
    .Q(\u_fir_pe2.rYin [2])
);

AOI22X1 _8559_ (
    .A(vdd),
    .B(\X[2]_5_bF$buf0 ),
    .C(gnd),
    .D(\X[2] [6]),
    .Y(_1996_)
);

NOR2X1 _8139_ (
    .A(_2344_),
    .B(_2334_),
    .Y(_2354_)
);

FILL FILL_1__7096_ (
);

FILL FILL_1__10807_ (
);

FILL FILL_0__7814_ (
);

INVX2 _9920_ (
    .A(\X[4] [3]),
    .Y(_3203_)
);

INVX1 _9500_ (
    .A(_2855_),
    .Y(_2856_)
);

FILL FILL_1__13279_ (
);

AOI21X1 _12977_ (
    .A(_6004_),
    .B(_6002_),
    .C(_5974_),
    .Y(_6014_)
);

NAND3X1 _12557_ (
    .A(_5599_),
    .B(_6365_),
    .C(_5598_),
    .Y(_5600_)
);

NOR2X1 _12137_ (
    .A(_5188_),
    .B(_5185_),
    .Y(_5253_)
);

FILL FILL_0__13213_ (
);

FILL FILL_2__6380_ (
);

FILL FILL254250x111750 (
);

FILL FILL_1__9662_ (
);

FILL FILL_1__9242_ (
);

FILL FILL_3__9168_ (
);

FILL FILL_1__10980_ (
);

FILL FILL_1__10560_ (
);

FILL FILL_1__10140_ (
);

FILL FILL_2__7585_ (
);

FILL FILL_2__7165_ (
);

OAI21X1 _6625_ (
    .A(_173_),
    .B(_223_),
    .C(_167_),
    .Y(_224_)
);

FILL FILL_2__12772_ (
);

FILL FILL_2__12352_ (
);

NOR2X1 _9097_ (
    .A(_2412_),
    .B(_2449_),
    .Y(_2458_)
);

FILL FILL_1__11765_ (
);

FILL FILL_1__11345_ (
);

FILL FILL_0__8772_ (
);

FILL FILL_0__8352_ (
);

FILL FILL_0__10338_ (
);

AND2X2 _10623_ (
    .A(_3865_),
    .B(_3875_),
    .Y(_3886_)
);

OAI21X1 _10203_ (
    .A(_3480_),
    .B(_3481_),
    .C(_3479_),
    .Y(_3482_)
);

NAND3X1 _13095_ (
    .A(_6121_),
    .B(_6125_),
    .C(_6129_),
    .Y(_6130_)
);

FILL FILL_2__9731_ (
);

FILL FILL_2__9311_ (
);

FILL FILL_1__6787_ (
);

FILL FILL_2__13137_ (
);

FILL FILL_0__9977_ (
);

FILL FILL_0__9557_ (
);

FILL FILL_3__7654_ (
);

FILL FILL_0__9137_ (
);

NAND3X1 _11828_ (
    .A(_4938_),
    .B(_4945_),
    .C(_4947_),
    .Y(_4948_)
);

AOI21X1 _11408_ (
    .A(_4542_),
    .B(_4544_),
    .C(_4599_),
    .Y(_4600_)
);

FILL FILL_0__12904_ (
);

FILL FILL_3__10484_ (
);

FILL FILL_0__10091_ (
);

FILL FILL_1__8933_ (
);

FILL FILL_1__8513_ (
);

FILL FILL_3__8439_ (
);

FILL FILL_3__8019_ (
);

NAND2X1 _7583_ (
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_1101_)
);

NAND2X1 _7163_ (
    .A(_746_),
    .B(_741_),
    .Y(_747_)
);

FILL FILL_3__9800_ (
);

FILL FILL_2__6856_ (
);

FILL FILL_2__6436_ (
);

FILL FILL_3__11269_ (
);

NOR2X1 _11581_ (
    .A(_4762_),
    .B(_4705_),
    .Y(_4777_[1])
);

FILL FILL_0__11296_ (
);

NAND2X1 _11161_ (
    .A(_4358_),
    .B(_4282_),
    .Y(_4359_)
);

FILL FILL_1__9718_ (
);

FILL FILL_3__12630_ (
);

FILL FILL_3__12210_ (
);

FILL FILL_2__11203_ (
);

INVX1 _8788_ (
    .A(_2210_),
    .Y(_2220_)
);

INVX1 _8368_ (
    .A(_1806_),
    .Y(_1807_)
);

FILL FILL_1__10616_ (
);

FILL FILL_0__7623_ (
);

FILL FILL_1__13088_ (
);

INVX1 _12786_ (
    .A(_5819_),
    .Y(_5825_)
);

FILL FILL_3__8192_ (
);

NOR2X1 _12366_ (
    .A(_5466_),
    .B(_5465_),
    .Y(_5469_)
);

FILL FILL_3__13415_ (
);

FILL FILL_2__12828_ (
);

FILL FILL_2__12408_ (
);

FILL FILL_0__13022_ (
);

FILL FILL_0__8828_ (
);

FILL FILL_3__6925_ (
);

FILL FILL_0__8408_ (
);

FILL FILL_1__9891_ (
);

FILL FILL_1__9471_ (
);

FILL FILL_1__9051_ (
);

FILL FILL_3__9397_ (
);

FILL FILL_2__7394_ (
);

OR2X2 _6854_ (
    .A(_380_),
    .B(_450_),
    .Y(_451_)
);

AND2X2 _6434_ (
    .A(gnd),
    .B(Xin[2]),
    .Y(_36_)
);

FILL FILL_2__12581_ (
);

FILL FILL_2__12161_ (
);

FILL FILL_1__11994_ (
);

FILL FILL_1__11574_ (
);

FILL FILL_1__11154_ (
);

FILL FILL_0__8581_ (
);

FILL FILL_2__8599_ (
);

FILL FILL_0__10987_ (
);

FILL FILL_0__8161_ (
);

FILL FILL_2__8179_ (
);

FILL FILL_0__10567_ (
);

NOR3X1 _10852_ (
    .A(_4038_),
    .B(_4005_),
    .C(_4050_),
    .Y(_4053_)
);

OAI22X1 _10432_ (
    .A(_3605_),
    .B(_3650_),
    .C(_3706_),
    .D(_3705_),
    .Y(_3707_)
);

FILL FILL_0__10147_ (
);

NAND3X1 _10012_ (
    .A(_3290_),
    .B(_3292_),
    .C(_3291_),
    .Y(_3293_)
);

FILL FILL_2__9960_ (
);

FILL FILL_2__9540_ (
);

FILL FILL_2__9120_ (
);

NAND3X1 _7639_ (
    .A(_1150_),
    .B(_1151_),
    .C(_1152_),
    .Y(_1157_)
);

DFFPOSX1 _7219_ (
    .D(Xin[4]),
    .CLK(clk_bF$buf41),
    .Q(\X[1] [4])
);

FILL FILL_1__6596_ (
);

FILL FILL_1__12779_ (
);

FILL FILL_1__12359_ (
);

FILL FILL_0__9786_ (
);

FILL FILL_3__7883_ (
);

FILL FILL_0__9366_ (
);

DFFPOSX1 _11637_ (
    .D(_4781_[13]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [13])
);

FILL FILL_3__7043_ (
);

AOI21X1 _11217_ (
    .A(_4400_),
    .B(_4407_),
    .C(_4382_),
    .Y(_4414_)
);

FILL FILL_1__13300_ (
);

FILL FILL_0__12713_ (
);

FILL FILL_1__8742_ (
);

FILL FILL_1__8322_ (
);

FILL FILL_3__8668_ (
);

NAND3X1 _7392_ (
    .A(_850_),
    .B(_908_),
    .C(_912_),
    .Y(_913_)
);

FILL FILL_2__6665_ (
);

NAND2X1 _11390_ (
    .A(_4582_),
    .B(_4581_),
    .Y(_4583_)
);

FILL FILL_1__9947_ (
);

FILL FILL_1__9527_ (
);

FILL FILL_1__9107_ (
);

FILL FILL_2__11852_ (
);

FILL FILL_2__11432_ (
);

FILL FILL_2__11012_ (
);

AOI21X1 _8597_ (
    .A(_2024_),
    .B(_2020_),
    .C(_1979_),
    .Y(_2034_)
);

NAND2X1 _8177_ (
    .A(\X[2] [4]),
    .B(vdd),
    .Y(_1619_)
);

FILL FILL_1__10845_ (
);

FILL FILL_1__10425_ (
);

FILL FILL_1__10005_ (
);

FILL FILL_0__7852_ (
);

FILL FILL_0__7432_ (
);

FILL FILL_0__7012_ (
);

NAND2X1 _12595_ (
    .A(_5633_),
    .B(_5636_),
    .Y(_5637_)
);

OAI21X1 _12175_ (
    .A(_5290_),
    .B(_5158_),
    .C(_5240_),
    .Y(_5291_)
);

FILL FILL_2__8811_ (
);

FILL FILL_3__13224_ (
);

FILL FILL_2__12637_ (
);

FILL FILL_2__12217_ (
);

FILL FILL_0__13251_ (
);

FILL FILL_0__8637_ (
);

FILL FILL_0__8217_ (
);

NAND3X1 _10908_ (
    .A(_4038_),
    .B(_4102_),
    .C(_4103_),
    .Y(_4109_)
);

FILL FILL_1__9280_ (
);

FILL FILL_3__7519_ (
);

AOI21X1 _6663_ (
    .A(_261_),
    .B(_260_),
    .C(_259_),
    .Y(_262_)
);

FILL FILL_2__12390_ (
);

FILL FILL_3__10769_ (
);

FILL FILL_3__10349_ (
);

FILL FILL_1__11383_ (
);

FILL FILL_0__8390_ (
);

FILL FILL_0__10796_ (
);

FILL FILL_0__10376_ (
);

AND2X2 _10661_ (
    .A(_3920_),
    .B(_3923_),
    .Y(_3925_)
);

AND2X2 _10241_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3519_)
);

FILL FILL_3__11710_ (
);

FILL FILL_2__10703_ (
);

NAND2X1 _7868_ (
    .A(_1379_),
    .B(_1381_),
    .Y(_1382_)
);

OAI21X1 _7448_ (
    .A(_966_),
    .B(_967_),
    .C(_965_),
    .Y(_968_)
);

NAND2X1 _7028_ (
    .A(_618_),
    .B(_617_),
    .Y(_620_)
);

FILL FILL_2__13175_ (
);

FILL FILL_0__6703_ (
);

FILL FILL_1__12588_ (
);

FILL FILL_1__12168_ (
);

FILL FILL_0__9595_ (
);

FILL FILL_0__9175_ (
);

AOI21X1 _11866_ (
    .A(_4902_),
    .B(_4908_),
    .C(_4985_),
    .Y(_4986_)
);

FILL FILL_3__7272_ (
);

INVX1 _11446_ (
    .A(\u_fir_pe5.rYin [3]),
    .Y(_4633_)
);

NAND2X1 _11026_ (
    .A(gnd),
    .B(\X[5] [6]),
    .Y(_4225_)
);

FILL FILL_2__11908_ (
);

FILL FILL_0__12942_ (
);

FILL FILL_0__12522_ (
);

FILL FILL_0__12102_ (
);

FILL FILL_0__7908_ (
);

FILL FILL_1__8551_ (
);

FILL FILL_3__8897_ (
);

FILL FILL_0__13307_ (
);

FILL FILL_2__6894_ (
);

FILL FILL_2__6474_ (
);

FILL FILL_1__9756_ (
);

FILL FILL_1__9336_ (
);

FILL FILL_2__11661_ (
);

FILL FILL_2__11241_ (
);

FILL FILL_1__10654_ (
);

FILL FILL_1__10234_ (
);

FILL FILL_2__7679_ (
);

FILL FILL_0__7661_ (
);

FILL FILL_2__7259_ (
);

FILL FILL_2__8620_ (
);

FILL FILL_2__8200_ (
);

OAI21X1 _6719_ (
    .A(_238_),
    .B(_316_),
    .C(_260_),
    .Y(_317_)
);

FILL FILL_2__12866_ (
);

FILL FILL_2__12446_ (
);

FILL FILL_2__12026_ (
);

FILL FILL_0__13060_ (
);

FILL FILL_1__11859_ (
);

FILL FILL_1__11439_ (
);

FILL FILL_1__11019_ (
);

FILL FILL_0__8866_ (
);

FILL FILL_3__6963_ (
);

FILL FILL_0__8446_ (
);

FILL FILL_3__6543_ (
);

DFFPOSX1 _10717_ (
    .D(_3978_[10]),
    .CLK(clk_bF$buf18),
    .Q(\Y[5] [10])
);

FILL FILL_0__8026_ (
);

FILL FILL_1__12800_ (
);

NOR2X1 _13189_ (
    .A(_6210_),
    .B(_6215_),
    .Y(_6218_)
);

FILL FILL_2__9825_ (
);

FILL FILL_2__9405_ (
);

FILL FILL_1__7822_ (
);

FILL FILL_1__7402_ (
);

FILL FILL_3__7748_ (
);

FILL FILL_3__7328_ (
);

NAND2X1 _6892_ (
    .A(_469_),
    .B(_466_),
    .Y(_488_)
);

NAND2X1 _6472_ (
    .A(_700_),
    .B(_72_),
    .Y(_73_)
);

FILL FILL_3__10578_ (
);

FILL FILL_1__11192_ (
);

NAND3X1 _10890_ (
    .A(_4086_),
    .B(_4090_),
    .C(_4054_),
    .Y(_4091_)
);

NOR3X1 _10470_ (
    .A(_3690_),
    .B(_3692_),
    .C(_3740_),
    .Y(_3744_)
);

FILL FILL_0__10185_ (
);

AND2X2 _10050_ (
    .A(gnd),
    .B(\X[4] [6]),
    .Y(_3330_)
);

FILL FILL_1__8607_ (
);

FILL FILL_2__10932_ (
);

FILL FILL_2__10512_ (
);

OAI21X1 _7677_ (
    .A(_1119_),
    .B(_1193_),
    .C(_1140_),
    .Y(_1194_)
);

INVX1 _7257_ (
    .A(_1497_),
    .Y(_1507_)
);

FILL FILL_0__6932_ (
);

FILL FILL_0__6512_ (
);

FILL FILL_1__12397_ (
);

NAND2X1 _11675_ (
    .A(_4795_),
    .B(_4791_),
    .Y(_4798_)
);

FILL FILL_3__7081_ (
);

OAI22X1 _11255_ (
    .A(_4000_),
    .B(_4447_),
    .C(_4448_),
    .D(_4450_),
    .Y(_4451_)
);

FILL FILL_3__12724_ (
);

FILL FILL_3__12304_ (
);

FILL FILL_2__11717_ (
);

FILL FILL_0__12751_ (
);

FILL FILL_0__12331_ (
);

FILL FILL_0__7717_ (
);

NAND2X1 _9823_ (
    .A(_3165_),
    .B(_3166_),
    .Y(_3181_[15])
);

NAND3X1 _9403_ (
    .A(_2691_),
    .B(_2755_),
    .C(_2756_),
    .Y(_2761_)
);

FILL FILL_1__8780_ (
);

FILL FILL_1__8360_ (
);

FILL FILL_3__8286_ (
);

BUFX2 _13401_ (
    .A(_6376_[7]),
    .Y(Xout[7])
);

FILL FILL_0__13116_ (
);

FILL FILL_1__9985_ (
);

FILL FILL_1__9565_ (
);

FILL FILL_1__9145_ (
);

FILL FILL_2__11890_ (
);

FILL FILL_2__11470_ (
);

FILL FILL_2__11050_ (
);

FILL FILL_1__10883_ (
);

FILL FILL_1__10463_ (
);

FILL FILL_1__10043_ (
);

FILL FILL_0__7890_ (
);

FILL FILL_0__7470_ (
);

FILL FILL_2__7488_ (
);

FILL FILL_0__7050_ (
);

FILL FILL_2__7068_ (
);

INVX1 _6948_ (
    .A(_515_),
    .Y(_543_)
);

INVX1 _6528_ (
    .A(_125_),
    .Y(_129_)
);

FILL FILL_2__12675_ (
);

FILL FILL_2__12255_ (
);

FILL FILL_1__11668_ (
);

FILL FILL_1__11248_ (
);

FILL FILL_0__8675_ (
);

FILL FILL_0__8255_ (
);

INVX1 _10946_ (
    .A(_4145_),
    .Y(_4146_)
);

NAND2X1 _10526_ (
    .A(_3777_),
    .B(_3776_),
    .Y(_3799_)
);

AOI21X1 _10106_ (
    .A(_3214_),
    .B(_3298_),
    .C(_3385_),
    .Y(_3386_)
);

FILL FILL_2__9634_ (
);

FILL FILL_2__9214_ (
);

FILL FILL_1__7631_ (
);

FILL FILL_3__7977_ (
);

FILL FILL_3__7137_ (
);

FILL FILL_0__12807_ (
);

FILL FILL_1__8836_ (
);

FILL FILL_1__8416_ (
);

FILL FILL_2__10321_ (
);

AOI21X1 _7486_ (
    .A(_969_),
    .B(_973_),
    .C(_935_),
    .Y(_1005_)
);

NAND2X1 _7066_ (
    .A(_652_),
    .B(_647_),
    .Y(_653_)
);

FILL FILL_0__6741_ (
);

FILL FILL_2__6759_ (
);

INVX1 _11484_ (
    .A(\u_fir_pe5.mul [7]),
    .Y(_4667_)
);

FILL FILL_0__11199_ (
);

NAND3X1 _11064_ (
    .A(_4207_),
    .B(_4248_),
    .C(_4253_),
    .Y(_4263_)
);

FILL FILL_3__12953_ (
);

FILL FILL_2__7700_ (
);

FILL FILL_3__12113_ (
);

FILL FILL_2__11946_ (
);

FILL FILL_0__12980_ (
);

FILL FILL_2__11526_ (
);

FILL FILL_0__12560_ (
);

FILL FILL_2__11106_ (
);

FILL FILL_0__12140_ (
);

FILL FILL_1__10939_ (
);

FILL FILL_1__10519_ (
);

FILL FILL_0__7946_ (
);

FILL FILL_0__7526_ (
);

INVX1 _9632_ (
    .A(_2984_),
    .Y(_2985_)
);

FILL FILL_0__7106_ (
);

AOI21X1 _9212_ (
    .A(_2562_),
    .B(_2558_),
    .C(_2543_),
    .Y(_2572_)
);

NAND2X1 _12689_ (
    .A(_5728_),
    .B(_5720_),
    .Y(_5729_)
);

OR2X2 _12269_ (
    .A(_5354_),
    .B(_5380_),
    .Y(_5382_)
);

FILL FILL_2__8905_ (
);

FILL FILL_3__13318_ (
);

NOR2X1 _13210_ (
    .A(_6234_),
    .B(_6235_),
    .Y(_6236_)
);

FILL FILL_1__6902_ (
);

FILL FILL_3__6408_ (
);

FILL FILL_1__9794_ (
);

FILL FILL_1__9374_ (
);

FILL FILL_1__10692_ (
);

FILL FILL_1__10272_ (
);

FILL FILL_2__7297_ (
);

FILL FILL_3__13071_ (
);

OAI21X1 _6757_ (
    .A(_341_),
    .B(_345_),
    .C(_348_),
    .Y(_355_)
);

FILL FILL_2__12064_ (
);

FILL FILL_1__11897_ (
);

FILL FILL_1__11477_ (
);

FILL FILL_1__11057_ (
);

FILL FILL_0__8484_ (
);

FILL FILL_3__6581_ (
);

DFFPOSX1 _10755_ (
    .D(_3984_[8]),
    .CLK(clk_bF$buf21),
    .Q(\u_fir_pe4.mul [8])
);

FILL FILL_0__8064_ (
);

NAND2X1 _10335_ (
    .A(_3603_),
    .B(_3610_),
    .Y(_3612_)
);

FILL FILL_3__11804_ (
);

FILL FILL_2__9443_ (
);

FILL FILL_0__11831_ (
);

FILL FILL_2__9023_ (
);

FILL FILL_0__11411_ (
);

FILL FILL_1__6499_ (
);

FILL FILL_2__13269_ (
);

AND2X2 _8903_ (
    .A(\u_fir_pe2.rYin [11]),
    .B(\u_fir_pe2.mul [11]),
    .Y(_2327_)
);

FILL FILL_1__7860_ (
);

FILL FILL_1__7440_ (
);

FILL FILL_1__7020_ (
);

FILL FILL_0__9689_ (
);

FILL FILL_0__9269_ (
);

FILL FILL_3__7366_ (
);

FILL FILL_1__13203_ (
);

NAND3X1 _12901_ (
    .A(_5932_),
    .B(_5933_),
    .C(_5934_),
    .Y(_5939_)
);

FILL FILL_0__12616_ (
);

FILL FILL_3__10196_ (
);

FILL FILL_1__8645_ (
);

FILL FILL_1__8225_ (
);

FILL FILL_2__10970_ (
);

FILL FILL_2__10550_ (
);

FILL FILL_2__10130_ (
);

NAND3X1 _7295_ (
    .A(_817_),
    .B(_1583_),
    .C(_816_),
    .Y(_818_)
);

FILL FILL_3__9512_ (
);

FILL FILL_2__6988_ (
);

FILL FILL_0__6970_ (
);

FILL FILL_0__6550_ (
);

FILL FILL_2__6568_ (
);

AOI21X1 _11293_ (
    .A(_4416_),
    .B(_4422_),
    .C(_4488_),
    .Y(_4489_)
);

FILL FILL_2__11755_ (
);

FILL FILL_2__11335_ (
);

FILL FILL_1__10328_ (
);

FILL FILL_0__7755_ (
);

DFFPOSX1 _9861_ (
    .D(\Y[3] [7]),
    .CLK(clk_bF$buf47),
    .Q(\u_fir_pe3.rYin [7])
);

FILL FILL_0__7335_ (
);

NAND2X1 _9441_ (
    .A(_2797_),
    .B(_2794_),
    .Y(_2798_)
);

INVX1 _9021_ (
    .A(_3172_),
    .Y(_3173_)
);

DFFPOSX1 _12498_ (
    .D(\Y[7] [13]),
    .CLK(clk_bF$buf11),
    .Q(\u_fir_pe6.rYin [13])
);

OAI21X1 _12078_ (
    .A(_5115_),
    .B(_5194_),
    .C(_5193_),
    .Y(_5195_)
);

FILL FILL_2__8714_ (
);

FILL FILL_0__13154_ (
);

FILL FILL_1__6711_ (
);

FILL FILL_3__6637_ (
);

FILL FILL_1__9183_ (
);

FILL FILL_0__9901_ (
);

FILL FILL_2__9919_ (
);

FILL FILL_1__10081_ (
);

FILL FILL_1__7916_ (
);

NAND3X1 _6986_ (
    .A(_561_),
    .B(_578_),
    .C(_577_),
    .Y(_580_)
);

NAND3X1 _6566_ (
    .A(_156_),
    .B(_163_),
    .C(_165_),
    .Y(_166_)
);

FILL FILL_2__12293_ (
);

FILL FILL_1__11286_ (
);

FILL FILL_0__8293_ (
);

FILL FILL_0__10699_ (
);

AOI21X1 _10984_ (
    .A(_4171_),
    .B(_4170_),
    .C(_4121_),
    .Y(_4184_)
);

INVX1 _10564_ (
    .A(_3828_),
    .Y(_3832_)
);

FILL FILL_0__10279_ (
);

INVX1 _10144_ (
    .A(\X[4] [7]),
    .Y(_3423_)
);

FILL FILL_2__9672_ (
);

FILL FILL_2__10606_ (
);

FILL FILL_2__9252_ (
);

FILL FILL_0__11640_ (
);

FILL FILL_0__11220_ (
);

FILL FILL_2__13078_ (
);

FILL FILL_0__6606_ (
);

INVX1 _8712_ (
    .A(_2146_),
    .Y(_2147_)
);

FILL FILL_0__9498_ (
);

FILL FILL_3__7595_ (
);

FILL FILL_0__9078_ (
);

AOI21X1 _11769_ (
    .A(_4885_),
    .B(_4886_),
    .C(_4884_),
    .Y(_4890_)
);

OAI21X1 _11349_ (
    .A(_4496_),
    .B(_4537_),
    .C(_4536_),
    .Y(_4543_)
);

FILL FILL_3__12818_ (
);

FILL FILL_1__13012_ (
);

FILL FILL_0__12845_ (
);

OAI21X1 _12710_ (
    .A(_5748_),
    .B(_5749_),
    .C(_5747_),
    .Y(_5750_)
);

FILL FILL_0__12425_ (
);

FILL FILL_0__12005_ (
);

OAI21X1 _9917_ (
    .A(_3192_),
    .B(_3195_),
    .C(_3189_),
    .Y(_3200_)
);

FILL FILL_1__8874_ (
);

FILL FILL_1__8454_ (
);

FILL FILL_1__8034_ (
);

FILL FILL_3__9741_ (
);

FILL FILL_2__6797_ (
);

FILL FILL_1__9659_ (
);

FILL FILL_1__9239_ (
);

FILL FILL_3__12571_ (
);

FILL FILL_3__12151_ (
);

FILL FILL_2__11984_ (
);

FILL FILL_2__11564_ (
);

FILL FILL_2__11144_ (
);

FILL FILL_1__10977_ (
);

FILL FILL_1__10557_ (
);

FILL FILL_1__10137_ (
);

FILL FILL_0__7984_ (
);

FILL FILL_0__7564_ (
);

OAI21X1 _9670_ (
    .A(_2958_),
    .B(_3008_),
    .C(_2986_),
    .Y(_3021_)
);

FILL FILL_0__7144_ (
);

NAND3X1 _9250_ (
    .A(_2602_),
    .B(_2608_),
    .C(_2607_),
    .Y(_2609_)
);

FILL FILL_2__8943_ (
);

FILL FILL_2__8523_ (
);

FILL FILL_0__10911_ (
);

FILL FILL_2__12769_ (
);

FILL FILL_2__12349_ (
);

FILL FILL253350x198150 (
);

FILL FILL_1__6940_ (
);

FILL FILL_1__6520_ (
);

FILL FILL_0__8769_ (
);

FILL FILL_3__6866_ (
);

FILL FILL_0__8349_ (
);

FILL FILL_1__12703_ (
);

FILL FILL_2__9728_ (
);

FILL FILL_0__9710_ (
);

FILL FILL_2__9308_ (
);

FILL FILL_1__7725_ (
);

FILL FILL_1__7305_ (
);

INVX1 _6795_ (
    .A(_386_),
    .Y(_392_)
);

FILL FILL254550x43350 (
);

FILL FILL_1__11095_ (
);

NAND3X1 _10793_ (
    .A(_3985_),
    .B(_3990_),
    .C(_3988_),
    .Y(_3996_)
);

OAI21X1 _10373_ (
    .A(_3615_),
    .B(_3617_),
    .C(_3611_),
    .Y(_3649_)
);

FILL FILL_0__10088_ (
);

FILL FILL_3__11422_ (
);

FILL FILL_2__10835_ (
);

FILL FILL_2__9481_ (
);

FILL FILL_2__10415_ (
);

FILL FILL_2__9061_ (
);

FILL FILL_0__6835_ (
);

OR2X2 _8941_ (
    .A(\u_fir_pe2.rYin [15]),
    .B(\u_fir_pe2.mul [15]),
    .Y(_2365_)
);

FILL FILL_0__6415_ (
);

OAI21X1 _8521_ (
    .A(_1950_),
    .B(_1946_),
    .C(_1953_),
    .Y(_1959_)
);

DFFPOSX1 _8101_ (
    .D(\Y[1] [1]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.rYin [1])
);

FILL FILL254250x50550 (
);

NAND2X1 _11998_ (
    .A(_5107_),
    .B(_5115_),
    .Y(_5116_)
);

NOR2X1 _11578_ (
    .A(\u_fir_pe5.rYin [0]),
    .B(\u_fir_pe5.mul [0]),
    .Y(_4761_)
);

NAND3X1 _11158_ (
    .A(_4286_),
    .B(_4347_),
    .C(_4342_),
    .Y(_4356_)
);

FILL FILL_3__12207_ (
);

FILL FILL_1__13241_ (
);

FILL FILL_0__12654_ (
);

FILL FILL_0__12234_ (
);

OR2X2 _9726_ (
    .A(_3063_),
    .B(_3068_),
    .Y(_3070_)
);

OAI21X1 _9306_ (
    .A(_2664_),
    .B(_2660_),
    .C(_2600_),
    .Y(_2665_)
);

FILL FILL_1__8683_ (
);

FILL FILL_1__8263_ (
);

FILL FILL_3__9970_ (
);

FILL FILL_3__9550_ (
);

FILL FILL_3__9130_ (
);

FILL FILL_0__13019_ (
);

AND2X2 _13304_ (
    .A(_6327_),
    .B(_6326_),
    .Y(_6369_[12])
);

FILL FILL_1__9888_ (
);

FILL FILL_1__9468_ (
);

FILL FILL_1__9048_ (
);

FILL FILL_3__12380_ (
);

FILL FILL_2__11793_ (
);

FILL FILL_2__11373_ (
);

FILL FILL_1__10786_ (
);

FILL FILL_1__10366_ (
);

FILL FILL_0__7793_ (
);

FILL FILL_0__7373_ (
);

FILL FILL_2__8752_ (
);

FILL FILL_2__8332_ (
);

FILL FILL_3__13165_ (
);

FILL FILL_0__10300_ (
);

FILL FILL_2__12998_ (
);

FILL FILL_2__12578_ (
);

FILL FILL_2__12158_ (
);

FILL FILL_0__13192_ (
);

FILL FILL_0__8578_ (
);

FILL FILL_3__6675_ (
);

FILL FILL_0__8158_ (
);

OAI21X1 _10849_ (
    .A(_4038_),
    .B(_4050_),
    .C(_4044_),
    .Y(_4051_)
);

NAND2X1 _10429_ (
    .A(_3672_),
    .B(_3675_),
    .Y(_3704_)
);

NAND2X1 _10009_ (
    .A(_3269_),
    .B(_3265_),
    .Y(_3290_)
);

FILL FILL_1__12932_ (
);

FILL FILL_2__9957_ (
);

FILL FILL_2__9537_ (
);

FILL FILL_0__11925_ (
);

FILL FILL_2__9117_ (
);

FILL FILL_0__11505_ (
);

FILL FILL_1__7954_ (
);

FILL FILL_1__7534_ (
);

FILL FILL_1__7114_ (
);

FILL FILL_3__8821_ (
);

AOI21X1 _10182_ (
    .A(_3460_),
    .B(_3459_),
    .C(_3458_),
    .Y(_3461_)
);

FILL FILL_1__8739_ (
);

FILL FILL_1__8319_ (
);

FILL FILL_3__11651_ (
);

FILL FILL_2__10644_ (
);

FILL FILL_2__9290_ (
);

FILL FILL_2__10224_ (
);

OAI21X1 _7389_ (
    .A(_905_),
    .B(_906_),
    .C(_866_),
    .Y(_910_)
);

FILL FILL_3__9606_ (
);

FILL FILL_0__6644_ (
);

NOR2X1 _8750_ (
    .A(_2183_),
    .B(_2182_),
    .Y(_2184_)
);

NAND3X1 _8330_ (
    .A(_1767_),
    .B(_1769_),
    .C(_1768_),
    .Y(_1770_)
);

NOR2X1 _11387_ (
    .A(_4220_),
    .B(_4447_),
    .Y(_4580_)
);

FILL FILL_2__7603_ (
);

FILL FILL_1__13050_ (
);

FILL FILL_2__11849_ (
);

FILL FILL_0__12883_ (
);

FILL FILL_2__11429_ (
);

FILL FILL_2__11009_ (
);

FILL FILL_0__12043_ (
);

FILL FILL_0__7849_ (
);

NAND3X1 _9955_ (
    .A(_3217_),
    .B(_3233_),
    .C(_3236_),
    .Y(_3237_)
);

FILL FILL_0__7429_ (
);

NAND2X1 _9535_ (
    .A(_2889_),
    .B(_2890_),
    .Y(_2891_)
);

FILL FILL_0__7009_ (
);

NAND2X1 _9115_ (
    .A(vdd),
    .B(\X[3] [4]),
    .Y(_2476_)
);

FILL FILL_1__8492_ (
);

FILL FILL_1__8072_ (
);

FILL FILL_2__8808_ (
);

FILL FILL_0__13248_ (
);

NOR2X1 _13113_ (
    .A(_6146_),
    .B(_6145_),
    .Y(_6147_)
);

FILL FILL_1__6805_ (
);

FILL FILL_1__9697_ (
);

FILL FILL_1__9277_ (
);

FILL FILL_2__11182_ (
);

FILL FILL_1__10595_ (
);

FILL FILL_1__10175_ (
);

FILL FILL_0__7182_ (
);

FILL FILL_3__10922_ (
);

FILL FILL_3__10502_ (
);

FILL FILL_2__8561_ (
);

FILL FILL_2__8141_ (
);

FILL FILL_3__13394_ (
);

FILL FILL_2__12387_ (
);

OAI21X1 _7601_ (
    .A(_1115_),
    .B(_1118_),
    .C(_1117_),
    .Y(_1119_)
);

FILL FILL_0__8387_ (
);

FILL FILL_3__6484_ (
);

NOR2X1 _10658_ (
    .A(\u_fir_pe4.rYin [11]),
    .B(\u_fir_pe4.mul [11]),
    .Y(_3922_)
);

OAI21X1 _10238_ (
    .A(_3277_),
    .B(_3332_),
    .C(_3515_),
    .Y(_3516_)
);

FILL FILL_3__11707_ (
);

FILL FILL_1__12741_ (
);

FILL FILL_1__12321_ (
);

FILL FILL_2__9766_ (
);

FILL FILL_2__9346_ (
);

FILL FILL_0__11734_ (
);

FILL FILL_0__11314_ (
);

OAI21X1 _8806_ (
    .A(_2226_),
    .B(_2227_),
    .C(_2231_),
    .Y(_2234_)
);

FILL FILL_1__7763_ (
);

FILL FILL_1__7343_ (
);

FILL FILL_3__7689_ (
);

FILL FILL_1__13106_ (
);

FILL FILL_0__12939_ (
);

INVX1 _12804_ (
    .A(_5746_),
    .Y(_5843_)
);

FILL FILL_0__12519_ (
);

FILL FILL_3__8210_ (
);

FILL FILL_3__11880_ (
);

FILL FILL_1__8548_ (
);

FILL FILL_3__11040_ (
);

FILL FILL_2__10873_ (
);

FILL FILL_2__10453_ (
);

FILL FILL_2__10033_ (
);

NOR2X1 _7198_ (
    .A(_779_),
    .B(_786_),
    .Y(_793_[2])
);

FILL FILL_0__6873_ (
);

FILL FILL_0__6453_ (
);

AND2X2 _11196_ (
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4393_)
);

FILL FILL_2__7832_ (
);

FILL FILL_3__12665_ (
);

FILL FILL_2__7412_ (
);

FILL FILL_3__12245_ (
);

FILL FILL_2__11658_ (
);

FILL FILL_0__12692_ (
);

FILL FILL_2__11238_ (
);

FILL FILL_0__12272_ (
);

FILL FILL_0__7658_ (
);

OAI21X1 _9764_ (
    .A(_3103_),
    .B(_3104_),
    .C(_3102_),
    .Y(_3108_)
);

INVX1 _9344_ (
    .A(_2695_),
    .Y(_2702_)
);

FILL FILL_2__8617_ (
);

FILL FILL_0__13057_ (
);

DFFPOSX1 _13342_ (
    .D(_6369_[4]),
    .CLK(clk_bF$buf46),
    .Q(\Y[7] [4])
);

FILL FILL_1__6614_ (
);

FILL FILL_1__9086_ (
);

FILL FILL_0__9804_ (
);

FILL FILL_3__7901_ (
);

FILL FILL_1__7819_ (
);

FILL FILL254250x237750 (
);

FILL FILL_2__8790_ (
);

FILL FILL_2__8370_ (
);

NAND2X1 _6889_ (
    .A(_482_),
    .B(_476_),
    .Y(_485_)
);

NAND2X1 _6469_ (
    .A(Xin[0]),
    .B(gnd),
    .Y(_70_)
);

FILL FILL_2__12196_ (
);

NAND2X1 _7830_ (
    .A(_1344_),
    .B(_1311_),
    .Y(_1345_)
);

OAI21X1 _7410_ (
    .A(_1507_),
    .B(_929_),
    .C(_874_),
    .Y(_930_)
);

FILL FILL_1__11189_ (
);

FILL FILL_0__8196_ (
);

OAI21X1 _10887_ (
    .A(_4083_),
    .B(_4084_),
    .C(_4069_),
    .Y(_4088_)
);

NAND3X1 _10467_ (
    .A(_3699_),
    .B(_3741_),
    .C(_3700_),
    .Y(_3742_)
);

NAND2X1 _10047_ (
    .A(\X[4] [1]),
    .B(vdd),
    .Y(_3327_)
);

FILL FILL_1__12970_ (
);

FILL FILL_3__11516_ (
);

FILL FILL_1__12550_ (
);

FILL FILL_1__12130_ (
);

FILL FILL_2__9995_ (
);

FILL FILL_2__10929_ (
);

FILL FILL_2__9575_ (
);

FILL FILL_0__11963_ (
);

FILL FILL_2__10509_ (
);

FILL FILL_2__9155_ (
);

FILL FILL_0__11543_ (
);

FILL FILL_0__11123_ (
);

FILL FILL_0__6929_ (
);

FILL FILL_0__6509_ (
);

AOI21X1 _8615_ (
    .A(_1966_),
    .B(_2036_),
    .C(_2050_),
    .Y(_2051_)
);

FILL FILL_1__7992_ (
);

FILL FILL_1__7572_ (
);

FILL FILL_1__7152_ (
);

FILL FILL_3__7078_ (
);

FILL FILL_1__13335_ (
);

FILL FILL254550x93750 (
);

FILL FILL_0__12748_ (
);

NAND2X1 _12613_ (
    .A(\X[6] [1]),
    .B(gnd),
    .Y(_5654_)
);

FILL FILL_0__12328_ (
);

FILL FILL_1__8777_ (
);

FILL FILL_1__8357_ (
);

FILL FILL_2__10682_ (
);

FILL FILL_2__10262_ (
);

FILL FILL_3__9224_ (
);

FILL FILL_0__6682_ (
);

FILL FILL_3__12894_ (
);

FILL FILL_2__7641_ (
);

FILL FILL_2__11887_ (
);

FILL FILL_2__11467_ (
);

FILL FILL_2__11047_ (
);

FILL FILL_0__12081_ (
);

FILL FILL_0__7887_ (
);

INVX1 _9993_ (
    .A(_3273_),
    .Y(_3274_)
);

FILL FILL_0__7467_ (
);

NAND2X1 _9573_ (
    .A(_2927_),
    .B(_2907_),
    .Y(_2928_)
);

FILL FILL_0__7047_ (
);

NAND3X1 _9153_ (
    .A(_2445_),
    .B(_2502_),
    .C(_2506_),
    .Y(_2514_)
);

FILL FILL_1__11821_ (
);

FILL FILL_1__11401_ (
);

FILL FILL_2__8846_ (
);

FILL FILL_2__8426_ (
);

FILL FILL_0__10814_ (
);

FILL FILL_3__13259_ (
);

FILL FILL_2__8006_ (
);

FILL FILL_0__13286_ (
);

NAND3X1 _13151_ (
    .A(_6157_),
    .B(_6159_),
    .C(_6183_),
    .Y(_6184_)
);

FILL FILL_1__6843_ (
);

FILL FILL_1__6423_ (
);

FILL FILL_1__12606_ (
);

FILL FILL_0__9613_ (
);

FILL FILL_3__10960_ (
);

FILL FILL_1__7628_ (
);

FILL FILL_3__10120_ (
);

AOI21X1 _6698_ (
    .A(_207_),
    .B(_285_),
    .C(_293_),
    .Y(_296_)
);

FILL FILL_3__8915_ (
);

NAND2X1 _10696_ (
    .A(_3957_),
    .B(_3959_),
    .Y(_3960_)
);

AOI21X1 _10276_ (
    .A(_3553_),
    .B(_3552_),
    .C(_3488_),
    .Y(_3554_)
);

FILL FILL_2__6912_ (
);

FILL FILL_3__11745_ (
);

FILL FILL_2__9384_ (
);

FILL FILL_0__11772_ (
);

FILL FILL_2__10318_ (
);

FILL FILL_0__11352_ (
);

FILL FILL_0__6738_ (
);

INVX1 _8844_ (
    .A(\u_fir_pe2.mul [6]),
    .Y(_2268_)
);

AOI21X1 _8424_ (
    .A(_1862_),
    .B(_1857_),
    .C(_1816_),
    .Y(_1863_)
);

OAI21X1 _8004_ (
    .A(_1506_),
    .B(_1503_),
    .C(_1505_),
    .Y(_1508_)
);

FILL FILL_1__7381_ (
);

FILL FILL_1__13144_ (
);

FILL FILL_0__12977_ (
);

INVX1 _12842_ (
    .A(_5879_),
    .Y(_5880_)
);

FILL FILL_0__12557_ (
);

FILL FILL_0__12137_ (
);

NOR2X1 _12422_ (
    .A(_5524_),
    .B(_5525_),
    .Y(_5526_)
);

NAND3X1 _12002_ (
    .A(_5112_),
    .B(_5116_),
    .C(_5114_),
    .Y(_5120_)
);

NOR2X1 _9629_ (
    .A(_2951_),
    .B(_2974_),
    .Y(_2982_)
);

INVX1 _9209_ (
    .A(_2487_),
    .Y(_2569_)
);

FILL FILL_1__8586_ (
);

FILL FILL_1__8166_ (
);

FILL FILL_2__10491_ (
);

FILL FILL_2__10071_ (
);

FILL FILL_3__9453_ (
);

NAND2X1 _13207_ (
    .A(_6232_),
    .B(_6233_),
    .Y(_6369_[3])
);

FILL FILL_0__6491_ (
);

FILL FILL_2__7870_ (
);

FILL FILL_2__7450_ (
);

FILL FILL_2__7030_ (
);

FILL FILL_2__11696_ (
);

FILL FILL_2__11276_ (
);

INVX1 _6910_ (
    .A(_505_),
    .Y(_506_)
);

FILL FILL_1__10689_ (
);

FILL FILL_1__10269_ (
);

FILL FILL_0__7696_ (
);

FILL FILL_0__7276_ (
);

NAND3X1 _9382_ (
    .A(_2733_),
    .B(_2734_),
    .C(_2735_),
    .Y(_2740_)
);

FILL FILL_1__11210_ (
);

FILL FILL_2__8655_ (
);

FILL FILL_2__8235_ (
);

FILL FILL_0__10623_ (
);

FILL FILL_0__10203_ (
);

FILL FILL_0__13095_ (
);

DFFPOSX1 _13380_ (
    .D(_6372_[2]),
    .CLK(clk_bF$buf27),
    .Q(\u_fir_pe7.mul [2])
);

FILL FILL_1__6652_ (
);

FILL FILL_3__6998_ (
);

FILL FILL_2__13002_ (
);

FILL FILL_3__6578_ (
);

FILL FILL_1__12835_ (
);

FILL FILL_1__12415_ (
);

FILL FILL_0__9422_ (
);

FILL FILL_0__11828_ (
);

FILL FILL_0__11408_ (
);

FILL FILL_1__7857_ (
);

FILL FILL_1__7437_ (
);

FILL FILL_1__7017_ (
);

FILL FILL_3__8304_ (
);

NAND3X1 _10085_ (
    .A(_3360_),
    .B(_3326_),
    .C(_3364_),
    .Y(_3365_)
);

FILL FILL_3__11974_ (
);

FILL FILL_2__6721_ (
);

FILL FILL_3__11134_ (
);

FILL FILL_2__10967_ (
);

FILL FILL_2__10547_ (
);

FILL FILL_2__9193_ (
);

FILL FILL_0__11581_ (
);

FILL FILL_2__10127_ (
);

FILL FILL_0__11161_ (
);

FILL FILL_3__9929_ (
);

FILL FILL_0__6967_ (
);

FILL FILL_0__6547_ (
);

NAND3X1 _8653_ (
    .A(_2054_),
    .B(_2088_),
    .C(_2086_),
    .Y(_2089_)
);

NAND3X1 _8233_ (
    .A(\X[2] [1]),
    .B(vdd),
    .C(_1673_),
    .Y(_1674_)
);

FILL FILL_1__7190_ (
);

FILL FILL_1__10901_ (
);

FILL FILL_2__7926_ (
);

FILL FILL_3__12759_ (
);

FILL FILL_2__7506_ (
);

FILL FILL_0__12786_ (
);

OAI21X1 _12651_ (
    .A(_5687_),
    .B(_5688_),
    .C(_5648_),
    .Y(_5692_)
);

FILL FILL_0__12366_ (
);

INVX1 _12231_ (
    .A(_5344_),
    .Y(_5345_)
);

DFFPOSX1 _9858_ (
    .D(\Y[3] [4]),
    .CLK(clk_bF$buf47),
    .Q(\u_fir_pe3.rYin [4])
);

AOI22X1 _9438_ (
    .A(gnd),
    .B(\X[3] [6]),
    .C(gnd),
    .D(\X[3] [7]),
    .Y(_2795_)
);

INVX2 _9018_ (
    .A(gnd),
    .Y(_3169_)
);

FILL FILL_1__8395_ (
);

FILL FILL254550x216150 (
);

NAND2X1 _13016_ (
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_6052_)
);

FILL FILL_1__6708_ (
);

FILL FILL_3__12092_ (
);

FILL FILL_2__11085_ (
);

FILL FILL_1__10498_ (
);

FILL FILL_1__10078_ (
);

FILL FILL_0__7085_ (
);

AOI22X1 _9191_ (
    .A(gnd),
    .B(\X[3] [3]),
    .C(gnd),
    .D(\X[3] [4]),
    .Y(_2551_)
);

FILL FILL_2__8884_ (
);

FILL FILL_2__8464_ (
);

FILL FILL_0__10852_ (
);

FILL FILL_0__10432_ (
);

FILL FILL_2__8044_ (
);

FILL FILL_0__10012_ (
);

NOR2X1 _7924_ (
    .A(_1432_),
    .B(_1431_),
    .Y(_1433_)
);

INVX1 _7504_ (
    .A(_1022_),
    .Y(_1023_)
);

FILL FILL_1__6881_ (
);

FILL FILL_1__6461_ (
);

FILL FILL_2__13231_ (
);

FILL FILL_1__12644_ (
);

FILL FILL_1__12224_ (
);

FILL FILL_0__9651_ (
);

FILL FILL_2__9669_ (
);

FILL FILL_2__9249_ (
);

FILL FILL_0__9231_ (
);

AND2X2 _11922_ (
    .A(_5019_),
    .B(_5014_),
    .Y(_5041_)
);

AND2X2 _11502_ (
    .A(_4644_),
    .B(_4654_),
    .Y(_4686_)
);

FILL FILL_0__11217_ (
);

OAI21X1 _8709_ (
    .A(_2090_),
    .B(_2143_),
    .C(_2086_),
    .Y(_2144_)
);

FILL FILL_1__7666_ (
);

FILL FILL_1__13009_ (
);

FILL FILL_3__8533_ (
);

INVX1 _12707_ (
    .A(_5734_),
    .Y(_5747_)
);

FILL FILL_2__6950_ (
);

FILL FILL_2__6530_ (
);

FILL FILL_3__11363_ (
);

FILL FILL_2__10776_ (
);

FILL FILL_2__10356_ (
);

FILL FILL_0__11390_ (
);

FILL FILL_1__9812_ (
);

FILL FILL_3__9318_ (
);

FILL FILL_0__6776_ (
);

AND2X2 _8882_ (
    .A(\u_fir_pe2.rYin [9]),
    .B(\u_fir_pe2.mul [9]),
    .Y(_2306_)
);

NOR2X1 _8462_ (
    .A(_2364_),
    .B(_1899_),
    .Y(_1900_)
);

AND2X2 _8042_ (
    .A(_1545_),
    .B(_1544_),
    .Y(_1587_[12])
);

OR2X2 _11099_ (
    .A(_4292_),
    .B(_4291_),
    .Y(_4297_)
);

FILL FILL_3__12988_ (
);

FILL FILL_2__7735_ (
);

FILL FILL_2__7315_ (
);

FILL FILL_3__12148_ (
);

FILL FILL_1__13182_ (
);

NAND3X1 _12880_ (
    .A(_5903_),
    .B(_5905_),
    .C(_5907_),
    .Y(_5918_)
);

FILL FILL_0__12595_ (
);

FILL FILL_0__12175_ (
);

NOR2X1 _12460_ (
    .A(_5561_),
    .B(_5568_),
    .Y(_5575_[2])
);

AOI21X1 _12040_ (
    .A(_5071_),
    .B(_4986_),
    .C(_5157_),
    .Y(_5158_)
);

FILL FILL_2__12922_ (
);

NAND3X1 _9667_ (
    .A(_3017_),
    .B(_3018_),
    .C(_3016_),
    .Y(_3019_)
);

OAI21X1 _9247_ (
    .A(_2530_),
    .B(_2605_),
    .C(_2534_),
    .Y(_2606_)
);

FILL FILL_1__11915_ (
);

FILL FILL_0__8922_ (
);

FILL FILL_0__8502_ (
);

FILL FILL_0__10908_ (
);

FILL FILL_3__9491_ (
);

FILL FILL_3__9071_ (
);

NAND2X1 _13245_ (
    .A(_6264_),
    .B(_6267_),
    .Y(_6369_[7])
);

FILL FILL_1__6937_ (
);

FILL FILL_1__6517_ (
);

FILL FILL_0__9707_ (
);

FILL FILL_3__7804_ (
);

FILL FILL_3__10214_ (
);

FILL FILL_2__8693_ (
);

FILL FILL_2__8273_ (
);

FILL FILL_0__10661_ (
);

FILL FILL_0__10241_ (
);

FILL FILL_2__12099_ (
);

NAND2X1 _7733_ (
    .A(_1249_),
    .B(_1248_),
    .Y(_1593_[9])
);

AOI22X1 _7313_ (
    .A(vdd),
    .B(\X[1] [1]),
    .C(vdd),
    .D(\X[1] [2]),
    .Y(_835_)
);

FILL FILL_1__6690_ (
);

FILL FILL_2__13040_ (
);

FILL FILL_3__11839_ (
);

FILL FILL_1__12873_ (
);

FILL FILL_1__12453_ (
);

FILL FILL_1__12033_ (
);

FILL FILL_2__9898_ (
);

FILL FILL_0__9460_ (
);

FILL FILL_2__9478_ (
);

FILL FILL_0__11866_ (
);

FILL FILL_2__9058_ (
);

FILL FILL_0__9040_ (
);

NAND2X1 _11731_ (
    .A(\X[7] [0]),
    .B(gnd),
    .Y(_4852_)
);

FILL FILL_0__11446_ (
);

FILL FILL_0__11026_ (
);

NAND2X1 _11311_ (
    .A(gnd),
    .B(_4459_),
    .Y(_4506_)
);

INVX1 _8938_ (
    .A(_2356_),
    .Y(_2361_)
);

NAND3X1 _8518_ (
    .A(_1954_),
    .B(_1955_),
    .C(_1953_),
    .Y(_1956_)
);

FILL FILL_1__7895_ (
);

FILL FILL_1__7475_ (
);

FILL FILL_1__7055_ (
);

FILL FILL_1__13238_ (
);

FILL FILL_3__8762_ (
);

NAND3X1 _12936_ (
    .A(_5971_),
    .B(_5967_),
    .C(_5972_),
    .Y(_5973_)
);

DFFPOSX1 _12516_ (
    .D(_5578_[15]),
    .CLK(clk_bF$buf49),
    .Q(\u_fir_pe6.mul [15])
);

FILL FILL_2__10585_ (
);

FILL FILL_2__10165_ (
);

FILL FILL_1__9621_ (
);

FILL FILL_1__9201_ (
);

FILL FILL_3__9547_ (
);

FILL FILL_0__6585_ (
);

OAI21X1 _8691_ (
    .A(_2125_),
    .B(_2124_),
    .C(_2118_),
    .Y(_2126_)
);

NAND3X1 _8271_ (
    .A(_1620_),
    .B(_1707_),
    .C(_1708_),
    .Y(_1712_)
);

FILL FILL_2__7964_ (
);

FILL FILL_2__7544_ (
);

FILL FILL_2__7124_ (
);

FILL FILL_2__12731_ (
);

FILL FILL_2__12311_ (
);

NOR2X1 _9896_ (
    .A(_3958_),
    .B(_3966_),
    .Y(_3968_)
);

NAND3X1 _9476_ (
    .A(_2773_),
    .B(_2828_),
    .C(_2832_),
    .Y(_2833_)
);

AOI22X1 _9056_ (
    .A(\X[3] [0]),
    .B(gnd),
    .C(gnd),
    .D(\X[3] [4]),
    .Y(_2418_)
);

FILL FILL_1__11724_ (
);

FILL FILL_1__11304_ (
);

FILL FILL_0__8731_ (
);

FILL FILL_2__8749_ (
);

FILL FILL_0__8311_ (
);

FILL FILL_2__8329_ (
);

FILL FILL_0__13189_ (
);

NOR2X1 _13054_ (
    .A(_6086_),
    .B(_6089_),
    .Y(_6375_[10])
);

FILL FILL_1__6746_ (
);

FILL FILL_1__12929_ (
);

FILL FILL_0__9936_ (
);

FILL FILL_0__9516_ (
);

FILL FILL_3__10863_ (
);

FILL FILL_3__10443_ (
);

FILL FILL_0__10890_ (
);

FILL FILL_0__10470_ (
);

FILL FILL_0__10050_ (
);

NAND2X1 _7962_ (
    .A(_1466_),
    .B(_1461_),
    .Y(_1467_)
);

INVX1 _7542_ (
    .A(_964_),
    .Y(_1061_)
);

INVX1 _7122_ (
    .A(_703_),
    .Y(_706_)
);

NOR2X1 _10599_ (
    .A(_3861_),
    .B(_3862_),
    .Y(_3863_)
);

AND2X2 _10179_ (
    .A(_3409_),
    .B(_3406_),
    .Y(_3458_)
);

FILL FILL_2__6815_ (
);

FILL FILL_3__11648_ (
);

FILL FILL_1__12682_ (
);

FILL FILL_3__11228_ (
);

FILL FILL_1__12262_ (
);

FILL FILL_2__9287_ (
);

AOI21X1 _11960_ (
    .A(_4989_),
    .B(_5067_),
    .C(_5075_),
    .Y(_5078_)
);

FILL FILL_0__11675_ (
);

AOI21X1 _11540_ (
    .A(_4720_),
    .B(_4711_),
    .C(_4718_),
    .Y(_4723_)
);

FILL FILL_0__11255_ (
);

NAND2X1 _11120_ (
    .A(gnd),
    .B(\X[5] [6]),
    .Y(_4318_)
);

NAND3X1 _8747_ (
    .A(_1971_),
    .B(_2044_),
    .C(_2150_),
    .Y(_2181_)
);

NAND2X1 _8327_ (
    .A(_1745_),
    .B(_1741_),
    .Y(_1767_)
);

FILL FILL_1__7284_ (
);

FILL FILL_1__13047_ (
);

AOI21X1 _12745_ (
    .A(_5773_),
    .B(_5781_),
    .C(_5784_),
    .Y(_5785_)
);

FILL FILL_3__8151_ (
);

NOR2X1 _12325_ (
    .A(_5430_),
    .B(_5431_),
    .Y(_5432_)
);

FILL FILL_0__13401_ (
);

FILL FILL_1__8489_ (
);

FILL FILL_1__8069_ (
);

FILL FILL_2__10394_ (
);

FILL FILL_1__9430_ (
);

FILL FILL_1__9010_ (
);

FILL FILL_3__9776_ (
);

FILL FILL_0__6394_ (
);

DFFPOSX1 _8080_ (
    .D(_1587_[4]),
    .CLK(clk_bF$buf44),
    .Q(\Y[2] [4])
);

FILL FILL_2__7773_ (
);

FILL FILL_2__7353_ (
);

FILL FILL_3__12186_ (
);

FILL FILL_2__11179_ (
);

NAND2X1 _6813_ (
    .A(vdd),
    .B(Xin[7]),
    .Y(_410_)
);

FILL FILL_2__12960_ (
);

FILL FILL_2__12540_ (
);

FILL FILL_2__12120_ (
);

FILL FILL_0__7599_ (
);

FILL FILL_0__7179_ (
);

NAND3X1 _9285_ (
    .A(_2637_),
    .B(_2640_),
    .C(_2638_),
    .Y(_2644_)
);

FILL FILL_1__11953_ (
);

FILL FILL_1__11533_ (
);

FILL FILL_1__11113_ (
);

FILL FILL_2__8558_ (
);

FILL FILL_0__8540_ (
);

FILL FILL_0__10946_ (
);

FILL FILL_2__8138_ (
);

FILL FILL_0__10526_ (
);

NOR2X1 _10811_ (
    .A(_4012_),
    .B(_4011_),
    .Y(_4013_)
);

FILL FILL_0__10106_ (
);

NOR2X1 _13283_ (
    .A(_6306_),
    .B(_6305_),
    .Y(_6307_)
);

FILL FILL_1__6975_ (
);

FILL FILL_1__6555_ (
);

FILL FILL_2__13325_ (
);

FILL FILL_1__12738_ (
);

FILL FILL_1__12318_ (
);

FILL FILL_0__9745_ (
);

FILL FILL_3__7842_ (
);

FILL FILL_0__9325_ (
);

FILL FILL_3__7422_ (
);

FILL FILL_3__7002_ (
);

FILL FILL_3__10672_ (
);

FILL FILL_1__8701_ (
);

FILL FILL_3__8627_ (
);

NAND3X1 _7771_ (
    .A(_1204_),
    .B(_1280_),
    .C(_1212_),
    .Y(_1287_)
);

NAND2X1 _7351_ (
    .A(\X[1] [1]),
    .B(gnd),
    .Y(_872_)
);

FILL FILL_2__6624_ (
);

FILL FILL_3__11457_ (
);

FILL FILL_1__12071_ (
);

FILL FILL_2__9096_ (
);

FILL FILL_0__11484_ (
);

FILL FILL_0__11064_ (
);

FILL FILL_1__9906_ (
);

FILL FILL_2__11811_ (
);

DFFPOSX1 _8976_ (
    .D(\X[2] [7]),
    .CLK(clk_bF$buf14),
    .Q(\X[3] [7])
);

AND2X2 _8556_ (
    .A(_1726_),
    .B(_1915_),
    .Y(_1993_)
);

NAND2X1 _8136_ (
    .A(gnd),
    .B(\X[2] [1]),
    .Y(_2325_)
);

FILL FILL_1__7093_ (
);

FILL FILL_1__10804_ (
);

FILL FILL_0__7811_ (
);

FILL FILL_2__7829_ (
);

FILL FILL_2__7409_ (
);

FILL FILL_1__13276_ (
);

INVX1 _12974_ (
    .A(_5933_),
    .Y(_6011_)
);

FILL FILL_0__12689_ (
);

FILL FILL_3__8380_ (
);

FILL FILL_0__12269_ (
);

NAND2X1 _12554_ (
    .A(_5593_),
    .B(_5596_),
    .Y(_5597_)
);

NAND2X1 _12134_ (
    .A(gnd),
    .B(_5180_),
    .Y(_5250_)
);

FILL FILL_0__13210_ (
);

FILL FILL_1__8298_ (
);

FILL FILL_3__9165_ (
);

DFFPOSX1 _13339_ (
    .D(_6369_[1]),
    .CLK(clk_bF$buf27),
    .Q(\Y[7] [1])
);

FILL FILL_2__7582_ (
);

FILL FILL_2__7162_ (
);

OAI21X1 _6622_ (
    .A(_219_),
    .B(_220_),
    .C(_210_),
    .Y(_221_)
);

AOI21X1 _9094_ (
    .A(_2452_),
    .B(_2455_),
    .C(_2446_),
    .Y(_2456_)
);

FILL FILL_1__11762_ (
);

FILL FILL_3__10308_ (
);

FILL FILL_1__11342_ (
);

FILL FILL_2__8787_ (
);

FILL FILL_2__8367_ (
);

FILL FILL_0__10335_ (
);

OAI21X1 _10620_ (
    .A(_3853_),
    .B(_3854_),
    .C(_3882_),
    .Y(_3883_)
);

NOR2X1 _10200_ (
    .A(_3395_),
    .B(_3392_),
    .Y(_3479_)
);

NAND2X1 _13092_ (
    .A(_6126_),
    .B(_6093_),
    .Y(_6127_)
);

NAND2X1 _7827_ (
    .A(_1336_),
    .B(_1333_),
    .Y(_1342_)
);

AND2X2 _7407_ (
    .A(_927_),
    .B(_923_),
    .Y(_1593_[5])
);

FILL FILL_1__6784_ (
);

FILL FILL_2__13134_ (
);

FILL FILL_1__12967_ (
);

FILL FILL_1__12547_ (
);

FILL FILL_1__12127_ (
);

FILL FILL_0__9974_ (
);

FILL FILL_0__9554_ (
);

FILL FILL_0__9134_ (
);

NAND3X1 _11825_ (
    .A(vdd),
    .B(\X[7] [4]),
    .C(_4935_),
    .Y(_4945_)
);

NAND3X1 _11405_ (
    .A(_4569_),
    .B(_4597_),
    .C(_4596_),
    .Y(_4598_)
);

FILL FILL_0__12901_ (
);

FILL FILL_1__7989_ (
);

FILL FILL_1__7569_ (
);

FILL FILL_1__7149_ (
);

FILL FILL_3__10061_ (
);

FILL FILL_1__8930_ (
);

FILL FILL_1__8510_ (
);

FILL FILL_3__8856_ (
);

FILL FILL_3__8016_ (
);

INVX1 _7580_ (
    .A(_1097_),
    .Y(_1098_)
);

NOR2X1 _7160_ (
    .A(_742_),
    .B(_743_),
    .Y(_744_)
);

FILL FILL_2__6853_ (
);

FILL FILL_3__11686_ (
);

FILL FILL_2__6433_ (
);

FILL FILL_2__10679_ (
);

FILL FILL_2__10259_ (
);

FILL FILL_0__11293_ (
);

FILL FILL_1__9715_ (
);

FILL FILL_2__11200_ (
);

FILL FILL_0__6679_ (
);

INVX1 _8785_ (
    .A(_2176_),
    .Y(_2217_)
);

NAND2X1 _8365_ (
    .A(\X[2] [0]),
    .B(gnd),
    .Y(_1804_)
);

FILL FILL_1__10613_ (
);

FILL FILL_0__7620_ (
);

FILL FILL_2__7638_ (
);

FILL FILL_1__13085_ (
);

NAND2X1 _12783_ (
    .A(_5820_),
    .B(_5821_),
    .Y(_5822_)
);

FILL FILL_0__12078_ (
);

NOR2X1 _12363_ (
    .A(\u_fir_pe6.rYin [7]),
    .B(\u_fir_pe6.mul [7]),
    .Y(_5466_)
);

FILL FILL_2__12825_ (
);

FILL FILL_2__12405_ (
);

FILL FILL_1__11818_ (
);

FILL FILL_0__8825_ (
);

FILL FILL_0__8405_ (
);

FILL FILL_3__6502_ (
);

FILL FILL_3__9394_ (
);

NAND2X1 _13148_ (
    .A(_6173_),
    .B(_6180_),
    .Y(_6181_)
);

FILL FILL_2__7391_ (
);

AOI21X1 _6851_ (
    .A(_436_),
    .B(_431_),
    .C(_383_),
    .Y(_448_)
);

NAND2X1 _6431_ (
    .A(gnd),
    .B(Xin[3]),
    .Y(_33_)
);

FILL FILL_3__10957_ (
);

FILL FILL_1__11991_ (
);

FILL FILL_3__10537_ (
);

FILL FILL_1__11571_ (
);

FILL FILL_3__10117_ (
);

FILL FILL_1__11151_ (
);

FILL FILL_2__8596_ (
);

FILL FILL_0__10984_ (
);

FILL FILL_2__8176_ (
);

FILL FILL_0__10564_ (
);

FILL FILL_0__10144_ (
);

OAI21X1 _7636_ (
    .A(_1153_),
    .B(_1149_),
    .C(_1100_),
    .Y(_1154_)
);

DFFPOSX1 _7216_ (
    .D(Xin[1]),
    .CLK(clk_bF$buf41),
    .Q(\X[1] [1])
);

FILL FILL_1__6593_ (
);

FILL FILL_2__6909_ (
);

FILL FILL_1__12776_ (
);

FILL FILL_1__12356_ (
);

FILL FILL_0__9783_ (
);

FILL FILL_0__9363_ (
);

FILL FILL_0__11769_ (
);

FILL FILL_3__7460_ (
);

DFFPOSX1 _11634_ (
    .D(_4781_[10]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.mul [10])
);

FILL FILL_0__11349_ (
);

NAND3X1 _11214_ (
    .A(_4380_),
    .B(_4408_),
    .C(_4410_),
    .Y(_4411_)
);

FILL FILL_0__12710_ (
);

FILL FILL_1__7798_ (
);

FILL FILL_1__7378_ (
);

FILL FILL_3__10290_ (
);

INVX1 _12839_ (
    .A(_5861_),
    .Y(_5877_)
);

FILL FILL_3__8245_ (
);

OAI21X1 _12419_ (
    .A(_5521_),
    .B(_5504_),
    .C(_5520_),
    .Y(_5523_)
);

FILL FILL_2__6662_ (
);

FILL FILL_3__11075_ (
);

FILL FILL_2__10488_ (
);

FILL FILL_2__10068_ (
);

FILL FILL_1__9944_ (
);

FILL FILL_1__9524_ (
);

FILL FILL_1__9104_ (
);

FILL FILL_0__6488_ (
);

NAND3X1 _8594_ (
    .A(_1977_),
    .B(_2025_),
    .C(_2030_),
    .Y(_2031_)
);

AOI21X1 _8174_ (
    .A(_1613_),
    .B(_1614_),
    .C(_2380_),
    .Y(_1617_)
);

FILL FILL_1__10842_ (
);

FILL FILL_1__10422_ (
);

FILL FILL_1__10002_ (
);

FILL FILL_2__7867_ (
);

FILL FILL_2__7447_ (
);

FILL FILL_2__7027_ (
);

NAND2X1 _12592_ (
    .A(_5588_),
    .B(_5593_),
    .Y(_5634_)
);

INVX1 _12172_ (
    .A(_5287_),
    .Y(_5288_)
);

NAND2X1 _6907_ (
    .A(_495_),
    .B(_501_),
    .Y(_503_)
);

FILL FILL_2__12634_ (
);

FILL FILL_2__12214_ (
);

INVX1 _9799_ (
    .A(\u_fir_pe3.mul [13]),
    .Y(_3143_)
);

OAI21X1 _9379_ (
    .A(_2732_),
    .B(_2736_),
    .C(_2708_),
    .Y(_2737_)
);

FILL FILL_1__11207_ (
);

FILL FILL_0__8634_ (
);

FILL FILL_3__6731_ (
);

FILL FILL_0__8214_ (
);

INVX1 _10905_ (
    .A(_4005_),
    .Y(_4106_)
);

DFFPOSX1 _13377_ (
    .D(\Y[6] [15]),
    .CLK(clk_bF$buf26),
    .Q(\u_fir_pe7.rYin [15])
);

FILL FILL_1__6649_ (
);

FILL FILL_3__7936_ (
);

FILL FILL_0__9419_ (
);

FILL FILL_3__7516_ (
);

AND2X2 _6660_ (
    .A(_237_),
    .B(_232_),
    .Y(_259_)
);

FILL FILL_1__11380_ (
);

FILL FILL_0__10793_ (
);

FILL FILL_0__10373_ (
);

FILL FILL_2__10700_ (
);

OAI21X1 _7865_ (
    .A(_1376_),
    .B(_1378_),
    .C(_1357_),
    .Y(_1379_)
);

INVX1 _7445_ (
    .A(_952_),
    .Y(_965_)
);

OAI21X1 _7025_ (
    .A(_594_),
    .B(_601_),
    .C(_600_),
    .Y(_617_)
);

FILL FILL_2__13172_ (
);

FILL FILL_2__6718_ (
);

FILL FILL_0__6700_ (
);

FILL FILL_1__12585_ (
);

FILL FILL_1__12165_ (
);

FILL FILL_0__11998_ (
);

FILL FILL_0__9592_ (
);

FILL FILL_0__9172_ (
);

OAI21X1 _11863_ (
    .A(_4981_),
    .B(_4982_),
    .C(_4980_),
    .Y(_4983_)
);

FILL FILL_0__11578_ (
);

NAND2X1 _11443_ (
    .A(_4630_),
    .B(_4629_),
    .Y(_4631_)
);

FILL FILL_0__11158_ (
);

NAND3X1 _11023_ (
    .A(_4210_),
    .B(_4219_),
    .C(_4221_),
    .Y(_4222_)
);

FILL FILL_3__12912_ (
);

FILL FILL_2__11905_ (
);

FILL FILL_1__7187_ (
);

FILL FILL_0__7905_ (
);

FILL FILL_3__8474_ (
);

OAI21X1 _12648_ (
    .A(_5687_),
    .B(_5688_),
    .C(_5686_),
    .Y(_5689_)
);

AND2X2 _12228_ (
    .A(_5324_),
    .B(_5319_),
    .Y(_5342_)
);

FILL FILL_0__13304_ (
);

FILL FILL_2__6891_ (
);

FILL FILL_2__6471_ (
);

FILL FILL_2__10297_ (
);

FILL FILL_1__9753_ (
);

FILL FILL_1__9333_ (
);

FILL FILL_3__9259_ (
);

FILL FILL_1__10651_ (
);

FILL FILL_1__10231_ (
);

FILL FILL_2__7676_ (
);

FILL FILL_2__7256_ (
);

FILL FILL_3__12089_ (
);

FILL FILL_3__13030_ (
);

NAND3X1 _6716_ (
    .A(_311_),
    .B(_313_),
    .C(_312_),
    .Y(_314_)
);

FILL FILL_2__12863_ (
);

FILL FILL_2__12443_ (
);

FILL FILL_2__12023_ (
);

INVX1 _9188_ (
    .A(_2547_),
    .Y(_2548_)
);

FILL FILL_1__11856_ (
);

FILL FILL_1__11436_ (
);

FILL FILL_1__11016_ (
);

FILL FILL_0__8863_ (
);

FILL FILL_3__6960_ (
);

FILL FILL_0__8443_ (
);

FILL FILL_0__10849_ (
);

FILL FILL_0__10429_ (
);

DFFPOSX1 _10714_ (
    .D(_3978_[7]),
    .CLK(clk_bF$buf18),
    .Q(\Y[5] [7])
);

FILL FILL_0__8023_ (
);

FILL FILL_0__10009_ (
);

FILL FILL254550x111750 (
);

NOR2X1 _13186_ (
    .A(_6214_),
    .B(_6213_),
    .Y(_6215_)
);

FILL FILL_2__9822_ (
);

FILL FILL_2__9402_ (
);

FILL FILL_1__6878_ (
);

FILL FILL_1__6458_ (
);

FILL FILL_2__13228_ (
);

FILL FILL_0__9648_ (
);

FILL FILL_3__7745_ (
);

FILL FILL_0__9228_ (
);

OAI21X1 _11919_ (
    .A(_5030_),
    .B(_5037_),
    .C(_5022_),
    .Y(_5038_)
);

FILL FILL_3__10155_ (
);

FILL FILL_0__10182_ (
);

FILL FILL_1__8604_ (
);

NAND3X1 _7674_ (
    .A(_1189_),
    .B(_1185_),
    .C(_1190_),
    .Y(_1191_)
);

DFFPOSX1 _7254_ (
    .D(_796_[15]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.mul [15])
);

FILL FILL_2__6947_ (
);

FILL FILL_2__6527_ (
);

FILL FILL_1__12394_ (
);

NAND3X1 _11672_ (
    .A(_4792_),
    .B(_4794_),
    .C(_4793_),
    .Y(_4795_)
);

FILL FILL_0__11387_ (
);

NOR3X1 _11252_ (
    .A(_4290_),
    .B(_4117_),
    .C(_4306_),
    .Y(_4448_)
);

FILL FILL_1__9809_ (
);

FILL FILL_3__12301_ (
);

FILL FILL_2__11714_ (
);

INVX1 _8879_ (
    .A(_2286_),
    .Y(_2302_)
);

OAI21X1 _8459_ (
    .A(_1816_),
    .B(_1896_),
    .C(_1865_),
    .Y(_1897_)
);

NOR2X1 _8039_ (
    .A(_1542_),
    .B(_1541_),
    .Y(_1543_)
);

FILL FILL_0__7714_ (
);

INVX1 _9820_ (
    .A(_3163_),
    .Y(_3164_)
);

OAI21X1 _9400_ (
    .A(_2757_),
    .B(_2754_),
    .C(_2690_),
    .Y(_2758_)
);

FILL FILL_1__13179_ (
);

OAI21X1 _12877_ (
    .A(_5914_),
    .B(_5908_),
    .C(_5902_),
    .Y(_5915_)
);

AOI21X1 _12457_ (
    .A(\X[7] [0]),
    .B(gnd),
    .C(_5482_),
    .Y(_5559_)
);

NAND2X1 _12037_ (
    .A(_5154_),
    .B(_5149_),
    .Y(_5155_)
);

FILL FILL_2__12919_ (
);

FILL FILL_0__13113_ (
);

FILL FILL_0__8919_ (
);

FILL FILL_1__9982_ (
);

FILL FILL_1__9562_ (
);

FILL FILL_1__9142_ (
);

FILL FILL_3__9488_ (
);

FILL FILL_1__10880_ (
);

FILL FILL_1__10460_ (
);

FILL FILL_1__10040_ (
);

FILL FILL_2__7485_ (
);

FILL FILL_2__7065_ (
);

NAND2X1 _6945_ (
    .A(_532_),
    .B(_535_),
    .Y(_540_)
);

NAND3X1 _6525_ (
    .A(_120_),
    .B(_125_),
    .C(_67_),
    .Y(_126_)
);

FILL FILL_2__12672_ (
);

FILL FILL_2__12252_ (
);

FILL FILL_1__11665_ (
);

FILL FILL_1__11245_ (
);

FILL FILL_0__8672_ (
);

FILL FILL_0__8252_ (
);

FILL FILL_0__10658_ (
);

AND2X2 _10943_ (
    .A(vdd),
    .B(\X[5] [4]),
    .Y(_4143_)
);

NAND2X1 _10523_ (
    .A(_3794_),
    .B(_3795_),
    .Y(_3796_)
);

FILL FILL_0__10238_ (
);

AOI21X1 _10103_ (
    .A(_3306_),
    .B(_3305_),
    .C(_3242_),
    .Y(_3383_)
);

FILL FILL_2__9631_ (
);

FILL FILL_2__9211_ (
);

FILL FILL_1__6687_ (
);

FILL FILL_2__13037_ (
);

FILL FILL_0__9457_ (
);

FILL FILL_3__7554_ (
);

FILL FILL_0__9037_ (
);

NOR2X1 _11728_ (
    .A(_4803_),
    .B(_4840_),
    .Y(_4849_)
);

AOI22X1 _11308_ (
    .A(\X[5]_5_bF$buf0 ),
    .B(gnd),
    .C(_4462_),
    .D(_4463_),
    .Y(_4503_)
);

FILL FILL_0__12804_ (
);

FILL FILL_3__10384_ (
);

FILL FILL_1__8833_ (
);

FILL FILL_1__8413_ (
);

FILL FILL_3__8339_ (
);

AOI21X1 _7483_ (
    .A(_991_),
    .B(_999_),
    .C(_1002_),
    .Y(_1003_)
);

NOR2X1 _7063_ (
    .A(_648_),
    .B(_649_),
    .Y(_650_)
);

FILL FILL_3__9700_ (
);

FILL FILL_2__6756_ (
);

FILL FILL_3__11169_ (
);

AND2X2 _11481_ (
    .A(_4664_),
    .B(_4663_),
    .Y(_4775_[6])
);

FILL FILL_0__11196_ (
);

INVX1 _11061_ (
    .A(_4162_),
    .Y(_4260_)
);

FILL FILL_1__9618_ (
);

FILL FILL_3__12530_ (
);

FILL FILL_2__11943_ (
);

FILL FILL_2__11523_ (
);

FILL FILL_2__11103_ (
);

NAND3X1 _8688_ (
    .A(_2119_),
    .B(_2122_),
    .C(_2076_),
    .Y(_2123_)
);

NAND3X1 _8268_ (
    .A(_1706_),
    .B(_1707_),
    .C(_1708_),
    .Y(_1709_)
);

FILL FILL_1__10936_ (
);

FILL FILL_1__10516_ (
);

FILL FILL_0__7943_ (
);

FILL FILL_0__7523_ (
);

FILL FILL_0__7103_ (
);

NAND3X1 _12686_ (
    .A(_5725_),
    .B(_5719_),
    .C(_5722_),
    .Y(_5726_)
);

OAI22X1 _12266_ (
    .A(_4926_),
    .B(_5244_),
    .C(_5087_),
    .D(_5017_),
    .Y(_5379_)
);

FILL FILL_2__8902_ (
);

FILL FILL_2__12728_ (
);

FILL FILL_2__12308_ (
);

FILL FILL_0__8728_ (
);

FILL FILL_3__6825_ (
);

FILL FILL_0__8308_ (
);

FILL FILL_1__9791_ (
);

FILL FILL_1__9371_ (
);

FILL FILL_2__7294_ (
);

FILL FILL254250x187350 (
);

AOI21X1 _6754_ (
    .A(_351_),
    .B(_346_),
    .C(_315_),
    .Y(_352_)
);

FILL FILL_2__12061_ (
);

FILL FILL_1__11894_ (
);

FILL FILL_1__11474_ (
);

FILL FILL_1__11054_ (
);

FILL FILL_2__8499_ (
);

FILL FILL_0__8481_ (
);

FILL FILL_0__10887_ (
);

FILL FILL_0__10467_ (
);

FILL FILL_0__8061_ (
);

DFFPOSX1 _10752_ (
    .D(_3984_[5]),
    .CLK(clk_bF$buf21),
    .Q(\u_fir_pe4.mul [5])
);

NAND2X1 _10332_ (
    .A(_3594_),
    .B(_3597_),
    .Y(_3609_)
);

FILL FILL_0__10047_ (
);

FILL FILL_3__11801_ (
);

FILL FILL_2__9440_ (
);

FILL FILL_2__9020_ (
);

NOR2X1 _7959_ (
    .A(_1462_),
    .B(_1463_),
    .Y(_1464_)
);

OAI21X1 _7539_ (
    .A(_1047_),
    .B(_1042_),
    .C(_1049_),
    .Y(_1058_)
);

NAND2X1 _7119_ (
    .A(_699_),
    .B(_702_),
    .Y(_703_)
);

FILL FILL_1__6496_ (
);

FILL FILL_2__13266_ (
);

OAI21X1 _8900_ (
    .A(_2320_),
    .B(_2321_),
    .C(_2316_),
    .Y(_2324_)
);

FILL FILL_1__12679_ (
);

FILL FILL_1__12259_ (
);

FILL FILL_0__9686_ (
);

FILL FILL_3__7783_ (
);

FILL FILL_0__9266_ (
);

OAI21X1 _11957_ (
    .A(_5074_),
    .B(_5075_),
    .C(_5073_),
    .Y(_5076_)
);

FILL FILL_3__7363_ (
);

NOR2X1 _11537_ (
    .A(_4720_),
    .B(_4717_),
    .Y(_4721_)
);

INVX1 _11117_ (
    .A(_4309_),
    .Y(_4315_)
);

FILL FILL_1__13200_ (
);

FILL FILL_0__12613_ (
);

FILL FILL_1__8642_ (
);

FILL FILL_1__8222_ (
);

FILL FILL_3__8568_ (
);

NAND2X1 _7292_ (
    .A(_811_),
    .B(_814_),
    .Y(_815_)
);

FILL FILL_2__6985_ (
);

FILL FILL_2__6565_ (
);

FILL FILL_3__11398_ (
);

NAND3X1 _11290_ (
    .A(_4481_),
    .B(_4482_),
    .C(_4485_),
    .Y(_4486_)
);

FILL FILL_1__9427_ (
);

FILL FILL_2__11752_ (
);

FILL FILL_2__11332_ (
);

AOI21X1 _8497_ (
    .A(_1930_),
    .B(_1934_),
    .C(_1916_),
    .Y(_1935_)
);

DFFPOSX1 _8077_ (
    .D(_1587_[1]),
    .CLK(clk_bF$buf45),
    .Q(\Y[2] [1])
);

FILL FILL_1__10325_ (
);

FILL FILL_0__7752_ (
);

FILL FILL_0__7332_ (
);

DFFPOSX1 _12495_ (
    .D(\Y[7] [10]),
    .CLK(clk_bF$buf39),
    .Q(\u_fir_pe6.rYin [10])
);

NAND2X1 _12075_ (
    .A(vdd),
    .B(\X[7] [7]),
    .Y(_5192_)
);

FILL FILL_2__8711_ (
);

FILL FILL_3__13124_ (
);

FILL FILL_2__12957_ (
);

FILL FILL_2__12537_ (
);

FILL FILL_2__12117_ (
);

FILL FILL_0__13151_ (
);

FILL FILL_0__8537_ (
);

NAND2X1 _10808_ (
    .A(\X[5] [4]),
    .B(vdd),
    .Y(_4010_)
);

FILL FILL_1__9180_ (
);

FILL FILL_2__9916_ (
);

FILL FILL_1__7913_ (
);

FILL FILL_3__7839_ (
);

NAND2X1 _6983_ (
    .A(_563_),
    .B(_576_),
    .Y(_577_)
);

NAND3X1 _6563_ (
    .A(vdd),
    .B(Xin[4]),
    .C(_153_),
    .Y(_163_)
);

FILL FILL_2__12290_ (
);

FILL FILL_3__10249_ (
);

FILL FILL_1__11283_ (
);

FILL FILL_0__8290_ (
);

FILL FILL_0__10696_ (
);

NAND3X1 _10981_ (
    .A(_4175_),
    .B(_4176_),
    .C(_4177_),
    .Y(_4181_)
);

AND2X2 _10561_ (
    .A(\u_fir_pe4.rYin [2]),
    .B(\u_fir_pe4.mul [2]),
    .Y(_3829_)
);

FILL FILL_0__10276_ (
);

NAND3X1 _10141_ (
    .A(_3414_),
    .B(_3419_),
    .C(_3417_),
    .Y(_3420_)
);

FILL FILL_2__10603_ (
);

NAND3X1 _7768_ (
    .A(_1267_),
    .B(_1283_),
    .C(_1281_),
    .Y(_1284_)
);

AND2X2 _7348_ (
    .A(gnd),
    .B(\X[1]_5_bF$buf1 ),
    .Y(_869_)
);

FILL FILL_2__13075_ (
);

FILL FILL_0__6603_ (
);

FILL FILL_1__12068_ (
);

FILL FILL_0__9495_ (
);

FILL FILL_0__9075_ (
);

NAND3X1 _11766_ (
    .A(_4884_),
    .B(_4886_),
    .C(_4885_),
    .Y(_4887_)
);

FILL FILL_3__7172_ (
);

NAND2X1 _11346_ (
    .A(_4539_),
    .B(_4540_),
    .Y(_4781_[11])
);

FILL FILL_2__11808_ (
);

FILL FILL_0__12842_ (
);

FILL FILL_0__12422_ (
);

FILL FILL_0__12002_ (
);

FILL FILL_0__7808_ (
);

NAND3X1 _9914_ (
    .A(_3928_),
    .B(_3196_),
    .C(_3194_),
    .Y(_3197_)
);

FILL FILL_1__8871_ (
);

FILL FILL_1__8451_ (
);

FILL FILL_1__8031_ (
);

FILL FILL_3__8797_ (
);

FILL FILL_0__13207_ (
);

FILL FILL_2__6794_ (
);

FILL FILL_1__9656_ (
);

FILL FILL_1__9236_ (
);

FILL FILL_2__11981_ (
);

FILL FILL_2__11561_ (
);

FILL FILL_2__11141_ (
);

FILL FILL_1__10974_ (
);

FILL FILL_1__10554_ (
);

FILL FILL_1__10134_ (
);

FILL FILL_2__7999_ (
);

FILL FILL_0__7981_ (
);

FILL FILL_0__7561_ (
);

FILL FILL_2__7579_ (
);

FILL FILL_0__7141_ (
);

FILL FILL_2__7159_ (
);

FILL FILL_2__8940_ (
);

FILL FILL_2__8520_ (
);

NAND3X1 _6619_ (
    .A(_211_),
    .B(_217_),
    .C(_216_),
    .Y(_218_)
);

FILL FILL_2__12766_ (
);

FILL FILL_2__12346_ (
);

FILL FILL_1__11759_ (
);

FILL FILL_1__11339_ (
);

FILL FILL_0__8766_ (
);

FILL FILL_0__8346_ (
);

FILL FILL_3__6443_ (
);

NOR2X1 _10617_ (
    .A(_3878_),
    .B(_3879_),
    .Y(_3880_)
);

FILL FILL_1__12700_ (
);

NAND2X1 _13089_ (
    .A(_6118_),
    .B(_6115_),
    .Y(_6124_)
);

FILL FILL_2__9725_ (
);

FILL FILL_2__9305_ (
);

FILL FILL_1__7722_ (
);

FILL FILL_1__7302_ (
);

INVX1 _6792_ (
    .A(_388_),
    .Y(_389_)
);

FILL FILL_3__10898_ (
);

FILL FILL_3__10478_ (
);

FILL FILL_3__10058_ (
);

FILL FILL_1__11092_ (
);

OAI21X1 _10790_ (
    .A(_3989_),
    .B(_3992_),
    .C(_3985_),
    .Y(_3993_)
);

INVX1 _10370_ (
    .A(_3645_),
    .Y(_3646_)
);

FILL FILL_0__10085_ (
);

FILL FILL_1__8927_ (
);

FILL FILL_1__8507_ (
);

FILL FILL_2__10832_ (
);

FILL FILL_2__10412_ (
);

OAI21X1 _7997_ (
    .A(_1489_),
    .B(_1490_),
    .C(_1500_),
    .Y(_1501_)
);

INVX1 _7577_ (
    .A(_1079_),
    .Y(_1095_)
);

OAI21X1 _7157_ (
    .A(_739_),
    .B(_722_),
    .C(_738_),
    .Y(_741_)
);

FILL FILL_0__6832_ (
);

FILL FILL_0__6412_ (
);

FILL FILL_1__12297_ (
);

AND2X2 _11995_ (
    .A(vdd),
    .B(\X[7] [6]),
    .Y(_5113_)
);

NAND3X1 _11575_ (
    .A(_4752_),
    .B(_4758_),
    .C(_4753_),
    .Y(_4759_)
);

AOI21X1 _11155_ (
    .A(_4263_),
    .B(_4262_),
    .C(_4194_),
    .Y(_4353_)
);

FILL FILL_3__12624_ (
);

FILL FILL_0__12651_ (
);

FILL FILL_0__12231_ (
);

FILL FILL_0__7617_ (
);

NOR2X1 _9723_ (
    .A(\u_fir_pe3.rYin [6]),
    .B(\u_fir_pe3.mul [6]),
    .Y(_3067_)
);

NAND3X1 _9303_ (
    .A(_2615_),
    .B(_2657_),
    .C(_2658_),
    .Y(_2662_)
);

FILL FILL_1__8680_ (
);

FILL FILL_1__8260_ (
);

FILL FILL_3__8186_ (
);

FILL FILL_3__13409_ (
);

FILL FILL_0__13016_ (
);

NOR2X1 _13301_ (
    .A(_6324_),
    .B(_6323_),
    .Y(_6325_)
);

FILL FILL_3__6919_ (
);

FILL FILL_1__9465_ (
);

FILL FILL_1__9045_ (
);

FILL FILL_2__11790_ (
);

FILL FILL_2__11370_ (
);

FILL FILL_1__10783_ (
);

FILL FILL_1__10363_ (
);

FILL FILL_0__7790_ (
);

FILL FILL_2__7388_ (
);

FILL FILL_0__7370_ (
);

OAI21X1 _6848_ (
    .A(_435_),
    .B(_434_),
    .C(_385_),
    .Y(_445_)
);

NAND2X1 _6428_ (
    .A(Xin[0]),
    .B(vdd),
    .Y(_30_)
);

FILL FILL_2__12995_ (
);

FILL FILL_2__12575_ (
);

FILL FILL_2__12155_ (
);

FILL FILL_1__11988_ (
);

FILL FILL_1__11568_ (
);

FILL FILL_1__11148_ (
);

FILL FILL_0__8575_ (
);

FILL FILL_3__6672_ (
);

FILL FILL_0__8155_ (
);

AOI21X1 _10846_ (
    .A(_4025_),
    .B(_4029_),
    .C(_4017_),
    .Y(_4048_)
);

NOR2X1 _10426_ (
    .A(_3681_),
    .B(_3686_),
    .Y(_3701_)
);

AOI22X1 _10006_ (
    .A(vdd),
    .B(\X[4] [4]),
    .C(_3276_),
    .D(_3278_),
    .Y(_3287_)
);

FILL FILL_2__9954_ (
);

FILL FILL_2__9534_ (
);

FILL FILL_0__11922_ (
);

FILL FILL_2__9114_ (
);

FILL FILL_0__11502_ (
);

FILL FILL_1__7951_ (
);

FILL FILL_1__7531_ (
);

FILL FILL_1__7111_ (
);

FILL FILL_3__7877_ (
);

FILL FILL_3__7457_ (
);

FILL FILL_3__7037_ (
);

FILL FILL_0__12707_ (
);

FILL FILL_1__8736_ (
);

FILL FILL_1__8316_ (
);

FILL FILL_2__10641_ (
);

FILL FILL_2__10221_ (
);

OAI21X1 _7386_ (
    .A(_905_),
    .B(_906_),
    .C(_904_),
    .Y(_907_)
);

FILL FILL_0__6641_ (
);

FILL FILL_2__6659_ (
);

FILL FILL_0__11099_ (
);

INVX1 _11384_ (
    .A(_4551_),
    .Y(_4577_)
);

FILL FILL_3__12853_ (
);

FILL FILL_2__7600_ (
);

FILL FILL_3__12013_ (
);

FILL FILL_2__11846_ (
);

FILL FILL_0__12880_ (
);

FILL FILL_2__11426_ (
);

FILL FILL_0__12460_ (
);

FILL FILL_2__11006_ (
);

FILL FILL_0__12040_ (
);

FILL FILL_1__10839_ (
);

FILL FILL_1__10419_ (
);

FILL FILL_0__7846_ (
);

INVX1 _9952_ (
    .A(_3220_),
    .Y(_3234_)
);

FILL FILL_0__7426_ (
);

NAND2X1 _9532_ (
    .A(_2884_),
    .B(_2852_),
    .Y(_2888_)
);

FILL FILL_0__7006_ (
);

AND2X2 _9112_ (
    .A(_2468_),
    .B(_2472_),
    .Y(_2473_)
);

NAND3X1 _12589_ (
    .A(_5607_),
    .B(_5630_),
    .C(_5629_),
    .Y(_5631_)
);

NAND2X1 _12169_ (
    .A(_5277_),
    .B(_5283_),
    .Y(_5285_)
);

FILL FILL_2__8805_ (
);

FILL FILL_3__13218_ (
);

FILL FILL_0__13245_ (
);

NOR2X1 _13110_ (
    .A(_5653_),
    .B(_6041_),
    .Y(_6144_)
);

FILL FILL_1__6802_ (
);

FILL FILL_1__9694_ (
);

FILL FILL_1__9274_ (
);

FILL FILL_1__10592_ (
);

FILL FILL_1__10172_ (
);

FILL FILL_2__7197_ (
);

OAI21X1 _6657_ (
    .A(_248_),
    .B(_255_),
    .C(_240_),
    .Y(_256_)
);

FILL FILL_2__12384_ (
);

FILL FILL_1__11797_ (
);

FILL FILL_1__11377_ (
);

FILL FILL_0__8384_ (
);

AND2X2 _10655_ (
    .A(_3917_),
    .B(_3918_),
    .Y(_3978_[10])
);

NAND2X1 _10235_ (
    .A(gnd),
    .B(\X[4]_5_bF$buf2 ),
    .Y(_3513_)
);

FILL FILL_2__9763_ (
);

FILL FILL_2__9343_ (
);

FILL FILL_0__11731_ (
);

FILL FILL_0__11311_ (
);

FILL FILL_1__6399_ (
);

FILL FILL_2__13169_ (
);

INVX1 _8803_ (
    .A(_2231_),
    .Y(_2232_)
);

FILL FILL_1__7760_ (
);

FILL FILL_1__7340_ (
);

FILL FILL_0__9589_ (
);

FILL FILL_0__9169_ (
);

FILL FILL_1__13103_ (
);

FILL FILL_0__12936_ (
);

OAI21X1 _12801_ (
    .A(_5829_),
    .B(_5824_),
    .C(_5831_),
    .Y(_5840_)
);

FILL FILL_3__10096_ (
);

FILL FILL_1__8545_ (
);

FILL FILL_2__10870_ (
);

FILL FILL_2__10450_ (
);

FILL FILL_2__10030_ (
);

AOI21X1 _7195_ (
    .A(Xin[0]),
    .B(gnd),
    .C(_700_),
    .Y(_777_)
);

FILL FILL_3__9412_ (
);

FILL FILL_2__6888_ (
);

FILL FILL_0__6870_ (
);

FILL FILL_0__6450_ (
);

FILL FILL_2__6468_ (
);

AND2X2 _11193_ (
    .A(vdd),
    .B(\X[5] [7]),
    .Y(_4390_)
);

FILL FILL_3__12242_ (
);

FILL FILL_2__11655_ (
);

FILL FILL_2__11235_ (
);

FILL FILL_1__10648_ (
);

FILL FILL_1__10228_ (
);

CLKBUF1 CLKBUF1_insert90 (
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert91 (
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert92 (
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert93 (
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert94 (
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

FILL FILL_0__7655_ (
);

NOR2X1 _9761_ (
    .A(_3104_),
    .B(_3103_),
    .Y(_3105_)
);

CLKBUF1 CLKBUF1_insert95 (
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

NOR2X1 _9341_ (
    .A(_2697_),
    .B(_2698_),
    .Y(_2699_)
);

CLKBUF1 CLKBUF1_insert96 (
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

AOI21X1 _12398_ (
    .A(_5496_),
    .B(_5474_),
    .C(_5494_),
    .Y(_5501_)
);

FILL FILL_2__8614_ (
);

FILL FILL_3__13027_ (
);

FILL FILL_0__13054_ (
);

FILL FILL_1__6611_ (
);

FILL FILL_3__6537_ (
);

FILL FILL_1__9083_ (
);

FILL FILL_2__9819_ (
);

FILL FILL_0__9801_ (
);

FILL FILL_1__7816_ (
);

NAND3X1 _6886_ (
    .A(_480_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

NOR2X1 _6466_ (
    .A(_21_),
    .B(_58_),
    .Y(_67_)
);

FILL FILL_2__12193_ (
);

FILL FILL_1__11186_ (
);

FILL FILL_0__8193_ (
);

FILL FILL_0__10599_ (
);

OAI21X1 _10884_ (
    .A(_4083_),
    .B(_4084_),
    .C(_4082_),
    .Y(_4085_)
);

NAND3X1 _10464_ (
    .A(_3730_),
    .B(_3734_),
    .C(_3738_),
    .Y(_3739_)
);

FILL FILL_0__10179_ (
);

NAND2X1 _10044_ (
    .A(_3323_),
    .B(_3322_),
    .Y(_3324_)
);

FILL FILL253650x198150 (
);

FILL FILL_2__9992_ (
);

FILL FILL_2__10926_ (
);

FILL FILL_2__9572_ (
);

FILL FILL_0__11960_ (
);

FILL FILL_2__10506_ (
);

FILL FILL_2__9152_ (
);

FILL FILL_0__11540_ (
);

FILL FILL_0__11120_ (
);

FILL FILL_2__13398_ (
);

FILL FILL_0__6926_ (
);

FILL FILL_0__6506_ (
);

NOR2X1 _8612_ (
    .A(_1967_),
    .B(_2047_),
    .Y(_2048_)
);

FILL FILL_0__9398_ (
);

FILL FILL_3__7495_ (
);

INVX1 _11669_ (
    .A(_5522_),
    .Y(_4792_)
);

OAI21X1 _11249_ (
    .A(_4371_),
    .B(_4375_),
    .C(_4373_),
    .Y(_4445_)
);

FILL FILL_3__12718_ (
);

FILL FILL_1__13332_ (
);

FILL FILL_0__12745_ (
);

AND2X2 _12610_ (
    .A(gnd),
    .B(\X[6]_5_bF$buf1 ),
    .Y(_5651_)
);

FILL FILL_0__12325_ (
);

NAND2X1 _9817_ (
    .A(\u_fir_pe3.rYin [15]),
    .B(\u_fir_pe3.mul [15]),
    .Y(_3160_)
);

FILL FILL_1__8774_ (
);

FILL FILL_1__8354_ (
);

FILL FILL_3__9641_ (
);

FILL FILL_2__6697_ (
);

FILL FILL_1__9979_ (
);

FILL FILL_1__9559_ (
);

FILL FILL_1__9139_ (
);

FILL FILL_2__11884_ (
);

FILL FILL_2__11464_ (
);

FILL FILL_2__11044_ (
);

FILL FILL_1__10877_ (
);

FILL FILL_1__10457_ (
);

FILL FILL_1__10037_ (
);

FILL FILL_0__7884_ (
);

NAND2X1 _9990_ (
    .A(gnd),
    .B(\X[4] [2]),
    .Y(_3271_)
);

FILL FILL_0__7464_ (
);

INVX1 _9570_ (
    .A(_2922_),
    .Y(_2925_)
);

FILL FILL_0__7044_ (
);

NAND3X1 _9150_ (
    .A(_2507_),
    .B(_2510_),
    .C(_2459_),
    .Y(_2511_)
);

FILL FILL_2__8843_ (
);

FILL FILL_2__8423_ (
);

FILL FILL_0__10811_ (
);

FILL FILL_2__8003_ (
);

FILL FILL_2__12669_ (
);

FILL FILL_2__12249_ (
);

FILL FILL_0__13283_ (
);

FILL FILL_1__6840_ (
);

FILL FILL_1__6420_ (
);

FILL FILL_0__8669_ (
);

FILL FILL_3__6766_ (
);

FILL FILL_0__8249_ (
);

FILL FILL_1__12603_ (
);

FILL FILL_0__9610_ (
);

FILL FILL_2__9628_ (
);

FILL FILL_2__9208_ (
);

FILL FILL_1__7625_ (
);

OAI21X1 _6695_ (
    .A(_292_),
    .B(_293_),
    .C(_291_),
    .Y(_294_)
);

NAND2X1 _10693_ (
    .A(_3952_),
    .B(_3946_),
    .Y(_3956_)
);

AOI21X1 _10273_ (
    .A(_3545_),
    .B(_3550_),
    .C(_3489_),
    .Y(_3551_)
);

FILL FILL_3__11742_ (
);

FILL FILL_3__11322_ (
);

FILL FILL_2__9381_ (
);

FILL FILL_2__10315_ (
);

FILL FILL_0__6735_ (
);

AND2X2 _8841_ (
    .A(_2265_),
    .B(_2264_),
    .Y(_2384_[5])
);

NAND3X1 _8421_ (
    .A(_1854_),
    .B(_1853_),
    .C(_1855_),
    .Y(_1860_)
);

NAND2X1 _8001_ (
    .A(_1501_),
    .B(_1504_),
    .Y(_1587_[8])
);

INVX1 _11898_ (
    .A(\X[7] [7]),
    .Y(_5017_)
);

NOR2X1 _11478_ (
    .A(_4661_),
    .B(_4660_),
    .Y(_4662_)
);

OAI21X1 _11058_ (
    .A(_4243_),
    .B(_4247_),
    .C(_4250_),
    .Y(_4257_)
);

FILL FILL_3__12947_ (
);

FILL FILL_3__12527_ (
);

FILL FILL_3__12107_ (
);

FILL FILL_1__13141_ (
);

FILL FILL_0__12974_ (
);

FILL FILL_0__12554_ (
);

FILL FILL_0__12134_ (
);

INVX1 _9626_ (
    .A(_2976_),
    .Y(_2980_)
);

NAND3X1 _9206_ (
    .A(_2553_),
    .B(_2557_),
    .C(_2559_),
    .Y(_2566_)
);

FILL FILL_1__8583_ (
);

FILL FILL_1__8163_ (
);

FILL FILL_3__9030_ (
);

NOR2X1 _13204_ (
    .A(_6230_),
    .B(_6229_),
    .Y(_6231_)
);

FILL FILL_1__9788_ (
);

FILL FILL_1__9368_ (
);

FILL FILL_3__12280_ (
);

FILL FILL_2__11693_ (
);

FILL FILL_2__11273_ (
);

FILL FILL_1__10686_ (
);

FILL FILL_1__10266_ (
);

FILL FILL_0__7693_ (
);

FILL FILL_0__7273_ (
);

FILL FILL_2__8652_ (
);

FILL FILL_2__8232_ (
);

FILL FILL_0__10620_ (
);

FILL FILL_3__13065_ (
);

FILL FILL_0__10200_ (
);

FILL FILL_2__12898_ (
);

FILL FILL_2__12058_ (
);

FILL FILL_0__13092_ (
);

FILL FILL_0__8898_ (
);

FILL FILL_3__6995_ (
);

FILL FILL_0__8478_ (
);

DFFPOSX1 _10749_ (
    .D(_3981_[2]),
    .CLK(clk_bF$buf3),
    .Q(\u_fir_pe4.mul [2])
);

FILL FILL_0__8058_ (
);

OAI21X1 _10329_ (
    .A(_3605_),
    .B(_3507_),
    .C(_3320_),
    .Y(_3606_)
);

FILL FILL_1__12832_ (
);

FILL FILL_1__12412_ (
);

FILL FILL_2__9437_ (
);

FILL FILL_0__11825_ (
);

FILL FILL_2__9017_ (
);

FILL FILL_0__11405_ (
);

FILL FILL_1__7854_ (
);

FILL FILL_1__7434_ (
);

FILL FILL_1__7014_ (
);

FILL FILL_3__8721_ (
);

FILL FILL_3__8301_ (
);

OAI21X1 _10082_ (
    .A(_3357_),
    .B(_3358_),
    .C(_3343_),
    .Y(_3362_)
);

FILL FILL_1__8639_ (
);

FILL FILL_1__8219_ (
);

FILL FILL_3__11551_ (
);

FILL FILL_2__10964_ (
);

FILL FILL_2__10544_ (
);

FILL FILL_2__9190_ (
);

FILL FILL_2__10124_ (
);

INVX2 _7289_ (
    .A(\X[1] [3]),
    .Y(_812_)
);

FILL FILL_3__9926_ (
);

FILL FILL_3__9506_ (
);

FILL FILL_0__6964_ (
);

FILL FILL_0__6544_ (
);

NAND3X1 _8650_ (
    .A(_2081_),
    .B(_2085_),
    .C(_2055_),
    .Y(_2086_)
);

NAND3X1 _8230_ (
    .A(_1670_),
    .B(_1665_),
    .C(_1667_),
    .Y(_1671_)
);

AOI21X1 _11287_ (
    .A(_4380_),
    .B(_4410_),
    .C(_4413_),
    .Y(_4483_)
);

FILL FILL_2__7923_ (
);

FILL FILL_2__7503_ (
);

FILL FILL_3__12336_ (
);

FILL FILL_2__11749_ (
);

FILL FILL_0__12783_ (
);

FILL FILL_2__11329_ (
);

FILL FILL_0__12363_ (
);

FILL FILL_0__7749_ (
);

DFFPOSX1 _9855_ (
    .D(\Y[3] [1]),
    .CLK(clk_bF$buf56),
    .Q(\u_fir_pe3.rYin [1])
);

FILL FILL_0__7329_ (
);

NAND2X1 _9435_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2792_)
);

AOI22X1 _9015_ (
    .A(\X[3] [0]),
    .B(gnd),
    .C(\X[3] [1]),
    .D(vdd),
    .Y(_3141_)
);

FILL FILL_1__8392_ (
);

FILL FILL_2__8708_ (
);

FILL FILL_0__13148_ (
);

AND2X2 _13013_ (
    .A(_6045_),
    .B(_6048_),
    .Y(_6049_)
);

FILL FILL_1__6705_ (
);

FILL FILL_1__9597_ (
);

FILL FILL_1__9177_ (
);

FILL FILL_2__11082_ (
);

FILL FILL_1__10495_ (
);

FILL FILL_1__10075_ (
);

FILL FILL_0__7082_ (
);

FILL FILL_3__10822_ (
);

FILL FILL_2__8881_ (
);

FILL FILL_2__8461_ (
);

FILL FILL_3__13294_ (
);

FILL FILL_2__8041_ (
);

FILL FILL_2__12287_ (
);

INVX1 _7921_ (
    .A(\u_fir_pe1.mul [1]),
    .Y(_1430_)
);

AOI21X1 _7501_ (
    .A(_959_),
    .B(_963_),
    .C(_952_),
    .Y(_1020_)
);

FILL FILL_0__8287_ (
);

AOI21X1 _10978_ (
    .A(_4177_),
    .B(_4176_),
    .C(_4175_),
    .Y(_4178_)
);

FILL FILL_3__6384_ (
);

NOR2X1 _10558_ (
    .A(_3819_),
    .B(_3824_),
    .Y(_3827_)
);

NAND2X1 _10138_ (
    .A(_3415_),
    .B(_3416_),
    .Y(_3417_)
);

FILL FILL_1__12641_ (
);

FILL FILL_1__12221_ (
);

FILL FILL_2__9666_ (
);

FILL FILL_2__9246_ (
);

FILL FILL_0__11214_ (
);

NAND2X1 _8706_ (
    .A(_2136_),
    .B(_2140_),
    .Y(_2141_)
);

FILL FILL_1__7663_ (
);

FILL FILL_1__13006_ (
);

FILL FILL_3__8950_ (
);

FILL FILL_0__12839_ (
);

NAND3X1 _12704_ (
    .A(vdd),
    .B(\X[6] [3]),
    .C(_5743_),
    .Y(_5744_)
);

FILL FILL_0__12419_ (
);

FILL FILL254550x237750 (
);

FILL FILL_1__8868_ (
);

FILL FILL_3__11780_ (
);

FILL FILL_1__8448_ (
);

FILL FILL_1__8028_ (
);

FILL FILL_2__10773_ (
);

FILL FILL_2__10353_ (
);

INVX1 _7098_ (
    .A(\u_fir_pe0.rYin [7]),
    .Y(_681_)
);

FILL FILL_3__9735_ (
);

FILL FILL_0__6773_ (
);

AND2X2 _11096_ (
    .A(_4292_),
    .B(_4291_),
    .Y(_4294_)
);

FILL FILL_2__7732_ (
);

FILL FILL_3__12565_ (
);

FILL FILL_2__7312_ (
);

FILL FILL_2__11978_ (
);

FILL FILL_2__11558_ (
);

FILL FILL_0__12592_ (
);

FILL FILL_2__11138_ (
);

FILL FILL_0__12172_ (
);

FILL FILL_0__7978_ (
);

FILL FILL_0__7558_ (
);

NAND2X1 _9664_ (
    .A(_3015_),
    .B(_2979_),
    .Y(_3016_)
);

FILL FILL_0__7138_ (
);

NAND2X1 _9244_ (
    .A(\X[3] [1]),
    .B(gnd),
    .Y(_2603_)
);

FILL FILL_1__11912_ (
);

FILL FILL_2__8937_ (
);

FILL FILL_2__8517_ (
);

FILL FILL_0__10905_ (
);

INVX1 _13242_ (
    .A(_6259_),
    .Y(_6265_)
);

FILL FILL_1__6934_ (
);

FILL FILL_1__6514_ (
);

FILL FILL_0__9704_ (
);

FILL FILL_1__7719_ (
);

FILL FILL_3__10631_ (
);

FILL FILL_3__10211_ (
);

FILL FILL_2__8690_ (
);

FILL FILL_2__8270_ (
);

NAND2X1 _6789_ (
    .A(Xin[2]),
    .B(gnd),
    .Y(_386_)
);

FILL FILL_2__12096_ (
);

AND2X2 _7730_ (
    .A(_1246_),
    .B(_1239_),
    .Y(_1247_)
);

AND2X2 _7310_ (
    .A(vdd),
    .B(\X[1] [1]),
    .Y(_832_)
);

FILL FILL_1__11089_ (
);

INVX1 _10787_ (
    .A(_3989_),
    .Y(_3990_)
);

NAND2X1 _10367_ (
    .A(_3642_),
    .B(_3485_),
    .Y(_3643_)
);

FILL FILL_3__11836_ (
);

FILL FILL_1__12870_ (
);

FILL FILL_3__11416_ (
);

FILL FILL_1__12450_ (
);

FILL FILL_1__12030_ (
);

FILL FILL_2__10829_ (
);

FILL FILL_2__9895_ (
);

FILL FILL_2__9475_ (
);

FILL FILL_0__11863_ (
);

FILL FILL_2__10409_ (
);

FILL FILL_2__9055_ (
);

FILL FILL_0__11443_ (
);

FILL FILL_0__11023_ (
);

FILL FILL_0__6829_ (
);

AND2X2 _8935_ (
    .A(_2352_),
    .B(_2358_),
    .Y(_2359_)
);

FILL FILL_0__6409_ (
);

AOI21X1 _8515_ (
    .A(_1864_),
    .B(_1866_),
    .C(_1952_),
    .Y(_1953_)
);

FILL FILL_1__7892_ (
);

FILL FILL_1__7472_ (
);

FILL FILL_1__7052_ (
);

FILL FILL_3__7398_ (
);

FILL FILL_3_BUFX2_insert71 (
);

FILL FILL_1__13235_ (
);

FILL FILL_3_BUFX2_insert73 (
);

FILL FILL_3_BUFX2_insert74 (
);

FILL FILL_3_BUFX2_insert76 (
);

OAI21X1 _12933_ (
    .A(_5969_),
    .B(_5968_),
    .C(_5965_),
    .Y(_5970_)
);

FILL FILL_3_BUFX2_insert78 (
);

FILL FILL_0__12648_ (
);

FILL FILL_0__12228_ (
);

DFFPOSX1 _12513_ (
    .D(_5578_[12]),
    .CLK(clk_bF$buf46),
    .Q(\u_fir_pe6.mul [12])
);

FILL FILL_1__8677_ (
);

FILL FILL_1__8257_ (
);

FILL FILL_2__10582_ (
);

FILL FILL_2__10162_ (
);

FILL FILL_3__9964_ (
);

FILL FILL_3__9124_ (
);

FILL FILL_0__6582_ (
);

FILL FILL_2__7961_ (
);

FILL FILL_3__12794_ (
);

FILL FILL_2__7541_ (
);

FILL FILL_2__7121_ (
);

FILL FILL_2__11787_ (
);

FILL FILL_2__11367_ (
);

FILL FILL_0__7787_ (
);

NOR2X1 _9893_ (
    .A(_3938_),
    .B(_3928_),
    .Y(_3948_)
);

FILL FILL_0__7367_ (
);

INVX1 _9473_ (
    .A(_2822_),
    .Y(_2830_)
);

NAND2X1 _9053_ (
    .A(\X[3] [0]),
    .B(gnd),
    .Y(_2415_)
);

FILL FILL_1__11721_ (
);

FILL FILL_1__11301_ (
);

FILL FILL_2__8746_ (
);

FILL FILL_2__8326_ (
);

FILL FILL_3__13159_ (
);

FILL FILL_0__13186_ (
);

NAND2X1 _13051_ (
    .A(_5956_),
    .B(_6029_),
    .Y(_6087_)
);

FILL FILL_1__6743_ (
);

FILL FILL_1__12926_ (
);

FILL FILL_0__9933_ (
);

FILL FILL_0__11919_ (
);

FILL FILL_0__9513_ (
);

FILL FILL_3__7610_ (
);

FILL FILL_1__7948_ (
);

FILL FILL_1__7528_ (
);

FILL FILL_1__7108_ (
);

AOI21X1 _6598_ (
    .A(_26_),
    .B(_110_),
    .C(_197_),
    .Y(_198_)
);

FILL FILL_3__8815_ (
);

OAI21X1 _10596_ (
    .A(_3853_),
    .B(_3854_),
    .C(_3858_),
    .Y(_3860_)
);

NAND3X1 _10176_ (
    .A(_3426_),
    .B(_3445_),
    .C(_3439_),
    .Y(_3455_)
);

FILL FILL_2__6812_ (
);

FILL FILL_2__10638_ (
);

FILL FILL_2__9284_ (
);

FILL FILL_0__11672_ (
);

FILL FILL_2__10218_ (
);

FILL FILL_0__11252_ (
);

FILL FILL_0__6638_ (
);

OR2X2 _8744_ (
    .A(_2177_),
    .B(_2154_),
    .Y(_2178_)
);

AOI22X1 _8324_ (
    .A(gnd),
    .B(\X[2]_5_bF$buf3 ),
    .C(_1753_),
    .D(_1755_),
    .Y(_1764_)
);

FILL FILL_1__7281_ (
);

FILL FILL_1__13044_ (
);

FILL FILL_0__12877_ (
);

NAND2X1 _12742_ (
    .A(_5781_),
    .B(_5773_),
    .Y(_5782_)
);

FILL FILL_0__12457_ (
);

FILL FILL_0__12037_ (
);

AOI21X1 _12322_ (
    .A(_5422_),
    .B(_5427_),
    .C(_5423_),
    .Y(_5429_)
);

NAND3X1 _9949_ (
    .A(gnd),
    .B(\X[4] [1]),
    .C(_3230_),
    .Y(_3231_)
);

NAND3X1 _9529_ (
    .A(_2814_),
    .B(_2817_),
    .C(_2884_),
    .Y(_2885_)
);

NAND2X1 _9109_ (
    .A(gnd),
    .B(\X[3]_5_bF$buf1 ),
    .Y(_2470_)
);

FILL FILL_1__8486_ (
);

FILL FILL_1__8066_ (
);

FILL FILL_2__10391_ (
);

FILL FILL_3__9353_ (
);

OAI21X1 _13107_ (
    .A(_6109_),
    .B(_6103_),
    .C(_6113_),
    .Y(_6141_)
);

FILL FILL_0__6391_ (
);

FILL FILL254250x223350 (
);

FILL FILL_2__7770_ (
);

FILL FILL_2__7350_ (
);

FILL FILL_3__12183_ (
);

FILL FILL_2__11176_ (
);

NAND2X1 _6810_ (
    .A(_406_),
    .B(_403_),
    .Y(_407_)
);

FILL FILL_1__10589_ (
);

FILL FILL_1__10169_ (
);

FILL FILL_0__7596_ (
);

FILL FILL_0__7176_ (
);

AOI21X1 _9282_ (
    .A(_2638_),
    .B(_2640_),
    .C(_2637_),
    .Y(_2641_)
);

FILL FILL_3__10916_ (
);

FILL FILL_1__11950_ (
);

FILL FILL_1__11530_ (
);

FILL FILL_1__11110_ (
);

FILL FILL_2__8555_ (
);

FILL FILL_0__10943_ (
);

FILL FILL_2__8135_ (
);

FILL FILL_0__10523_ (
);

FILL FILL_0__10103_ (
);

INVX1 _13280_ (
    .A(\u_fir_pe7.mul [10]),
    .Y(_6304_)
);

FILL FILL_1__6972_ (
);

FILL FILL_1__6552_ (
);

FILL FILL_2__13322_ (
);

FILL FILL_3__6478_ (
);

FILL FILL_1__12735_ (
);

FILL FILL_1__12315_ (
);

FILL FILL_0__9742_ (
);

FILL FILL_0__9322_ (
);

FILL FILL_0__11728_ (
);

FILL FILL_0__11308_ (
);

FILL FILL_1__7757_ (
);

FILL FILL_1__7337_ (
);

FILL FILL_3__8624_ (
);

FILL FILL_2__6621_ (
);

FILL FILL_3__11034_ (
);

FILL FILL_2__10867_ (
);

FILL FILL_2__10447_ (
);

FILL FILL_2__9093_ (
);

FILL FILL_0__11481_ (
);

FILL FILL_2__10027_ (
);

FILL FILL_0__11061_ (
);

FILL FILL_1__9903_ (
);

FILL FILL_3__9829_ (
);

FILL FILL_0__6867_ (
);

DFFPOSX1 _8973_ (
    .D(\X[2] [4]),
    .CLK(clk_bF$buf28),
    .Q(\X[3] [4])
);

FILL FILL_0__6447_ (
);

AOI21X1 _8553_ (
    .A(_1933_),
    .B(_1932_),
    .C(_1917_),
    .Y(_1990_)
);

AND2X2 _8133_ (
    .A(\X[2] [1]),
    .B(vdd),
    .Y(_2294_)
);

FILL FILL_1__7090_ (
);

FILL FILL_1__10801_ (
);

FILL FILL_2__7826_ (
);

FILL FILL_3__12659_ (
);

FILL FILL_2__7406_ (
);

FILL FILL_1__13273_ (
);

AOI21X1 _12971_ (
    .A(_5994_),
    .B(_6001_),
    .C(_5976_),
    .Y(_6008_)
);

FILL FILL_0__12686_ (
);

FILL FILL_0__12266_ (
);

INVX2 _12551_ (
    .A(\X[6] [3]),
    .Y(_5594_)
);

INVX1 _12131_ (
    .A(_5246_),
    .Y(_5247_)
);

OAI21X1 _9758_ (
    .A(_3100_),
    .B(_3097_),
    .C(_3099_),
    .Y(_3102_)
);

INVX2 _9338_ (
    .A(gnd),
    .Y(_2696_)
);

FILL FILL_1__8295_ (
);

FILL FILL_3__9582_ (
);

NOR2X1 _13336_ (
    .A(_6299_),
    .B(_6363_),
    .Y(_6358_)
);

FILL FILL_1__6608_ (
);

FILL FILL253350x61350 (
);

FILL FILL_1__10398_ (
);

INVX1 _9091_ (
    .A(_2436_),
    .Y(_2453_)
);

FILL FILL_3__10305_ (
);

FILL FILL_2__8784_ (
);

FILL FILL_2__8364_ (
);

FILL FILL_0__10332_ (
);

NAND3X1 _7824_ (
    .A(_1312_),
    .B(_1338_),
    .C(_1334_),
    .Y(_1339_)
);

INVX1 _7404_ (
    .A(_917_),
    .Y(_925_)
);

FILL FILL_1__6781_ (
);

FILL FILL_2__13131_ (
);

FILL FILL_1__12964_ (
);

FILL FILL_1__12544_ (
);

FILL FILL_1__12124_ (
);

FILL FILL_2__9989_ (
);

FILL FILL_0__9971_ (
);

FILL FILL_0__9551_ (
);

FILL FILL_2__9569_ (
);

FILL FILL_0__11957_ (
);

FILL FILL_0__9131_ (
);

FILL FILL_2__9149_ (
);

AOI22X1 _11822_ (
    .A(gnd),
    .B(\X[7] [3]),
    .C(vdd),
    .D(\X[7] [4]),
    .Y(_4942_)
);

FILL FILL_0__11537_ (
);

OAI21X1 _11402_ (
    .A(_4576_),
    .B(_4571_),
    .C(_4594_),
    .Y(_4595_)
);

FILL FILL_0__11117_ (
);

NAND2X1 _8609_ (
    .A(_2044_),
    .B(_1974_),
    .Y(_2046_)
);

FILL FILL_1__7986_ (
);

FILL FILL_1__7566_ (
);

FILL FILL_1__7146_ (
);

FILL FILL_1__13329_ (
);

FILL FILL_3__8433_ (
);

OAI21X1 _12607_ (
    .A(_5608_),
    .B(_5642_),
    .C(_5624_),
    .Y(_5648_)
);

FILL FILL_2__6850_ (
);

FILL FILL_3__11683_ (
);

FILL FILL_2__6430_ (
);

FILL FILL_3__11263_ (
);

FILL FILL_2__10676_ (
);

FILL FILL_2__10256_ (
);

FILL FILL_0__11290_ (
);

FILL FILL_1__9712_ (
);

FILL FILL_3__9218_ (
);

FILL FILL_0__6676_ (
);

NAND2X1 _8782_ (
    .A(_2212_),
    .B(_2211_),
    .Y(_2214_)
);

INVX1 _8362_ (
    .A(_1796_),
    .Y(_1801_)
);

FILL FILL_1__10610_ (
);

FILL FILL_3__12888_ (
);

FILL FILL_2__7635_ (
);

FILL FILL_3__12048_ (
);

FILL FILL_1__13082_ (
);

NAND2X1 _12780_ (
    .A(gnd),
    .B(\X[6] [6]),
    .Y(_5819_)
);

FILL FILL_0__12075_ (
);

INVX1 _12360_ (
    .A(\u_fir_pe6.rYin [7]),
    .Y(_5463_)
);

FILL FILL_2__12822_ (
);

FILL FILL_2__12402_ (
);

NAND3X1 _9987_ (
    .A(\X[4] [1]),
    .B(gnd),
    .C(_3267_),
    .Y(_3268_)
);

AOI21X1 _9567_ (
    .A(_2873_),
    .B(_2916_),
    .C(_2919_),
    .Y(_2922_)
);

NAND3X1 _9147_ (
    .A(_2503_),
    .B(_2497_),
    .C(_2501_),
    .Y(_2508_)
);

FILL FILL_1__11815_ (
);

FILL FILL_0__8822_ (
);

FILL FILL_0__8402_ (
);

FILL FILL_0__10808_ (
);

NAND2X1 _13145_ (
    .A(_6177_),
    .B(_6151_),
    .Y(_6178_)
);

FILL FILL_1__6837_ (
);

FILL FILL_1__6417_ (
);

FILL FILL_0__9607_ (
);

FILL FILL_3__7704_ (
);

FILL FILL_3__10534_ (
);

FILL FILL_2__8593_ (
);

FILL FILL_0__10981_ (
);

FILL FILL_2__8173_ (
);

FILL FILL_0__10561_ (
);

FILL FILL_0__10141_ (
);

NAND3X1 _7633_ (
    .A(_1146_),
    .B(_1147_),
    .C(_1114_),
    .Y(_1151_)
);

DFFPOSX1 _7213_ (
    .D(_790_[14]),
    .CLK(clk_bF$buf25),
    .Q(\Y[1] [14])
);

FILL FILL_1__6590_ (
);

FILL FILL_2__6906_ (
);

FILL FILL_1__12773_ (
);

FILL FILL_1__12353_ (
);

FILL FILL_0__9780_ (
);

FILL FILL_2__9798_ (
);

FILL FILL_2__9378_ (
);

FILL FILL_0__9360_ (
);

FILL FILL_0__11766_ (
);

DFFPOSX1 _11631_ (
    .D(_4781_[7]),
    .CLK(clk_bF$buf31),
    .Q(\u_fir_pe5.mul [7])
);

FILL FILL_0__11346_ (
);

NAND3X1 _11211_ (
    .A(_4400_),
    .B(_4407_),
    .C(_4382_),
    .Y(_4408_)
);

NOR2X1 _8838_ (
    .A(_2262_),
    .B(_2261_),
    .Y(_2263_)
);

OAI21X1 _8418_ (
    .A(_1852_),
    .B(_1856_),
    .C(_1818_),
    .Y(_1857_)
);

FILL FILL_1__7795_ (
);

FILL FILL_1__7375_ (
);

FILL FILL_1__13138_ (
);

FILL FILL_3__8662_ (
);

NAND3X1 _12836_ (
    .A(_5864_),
    .B(_5867_),
    .C(_5783_),
    .Y(_5874_)
);

FILL FILL_3__8242_ (
);

NOR2X1 _12416_ (
    .A(_5518_),
    .B(_5519_),
    .Y(_5572_[11])
);

FILL FILL_3__11492_ (
);

FILL FILL_2__10485_ (
);

FILL FILL_2__10065_ (
);

FILL FILL_1__9941_ (
);

FILL FILL_1__9521_ (
);

FILL FILL_1__9101_ (
);

FILL FILL_3__9447_ (
);

FILL FILL_0__6485_ (
);

INVX1 _8591_ (
    .A(_2020_),
    .Y(_2028_)
);

NAND3X1 _8171_ (
    .A(_2376_),
    .B(_1608_),
    .C(_1611_),
    .Y(_1614_)
);

FILL FILL_2__7864_ (
);

FILL FILL_2__7444_ (
);

FILL FILL_3__12277_ (
);

FILL FILL_2__7024_ (
);

NAND2X1 _6904_ (
    .A(_498_),
    .B(_499_),
    .Y(_500_)
);

FILL FILL_2__12631_ (
);

FILL FILL_2__12211_ (
);

AND2X2 _9796_ (
    .A(_3139_),
    .B(_3138_),
    .Y(_3181_[12])
);

NAND3X1 _9376_ (
    .A(_2714_),
    .B(_2729_),
    .C(_2730_),
    .Y(_2734_)
);

FILL FILL_1__11204_ (
);

FILL FILL_2__8649_ (
);

FILL FILL_0__8631_ (
);

FILL FILL_2__8229_ (
);

FILL FILL_0__8211_ (
);

FILL FILL_0__10617_ (
);

NAND3X1 _10902_ (
    .A(_4011_),
    .B(_4098_),
    .C(_4099_),
    .Y(_4103_)
);

FILL FILL_0__13089_ (
);

DFFPOSX1 _13374_ (
    .D(\Y[6] [12]),
    .CLK(clk_bF$buf50),
    .Q(\u_fir_pe7.rYin [12])
);

FILL FILL_1__6646_ (
);

FILL FILL_2__13416_ (
);

FILL FILL_1__12829_ (
);

FILL FILL_1__12409_ (
);

FILL FILL_3__7933_ (
);

FILL FILL_0__9416_ (
);

FILL FILL_3__10763_ (
);

FILL FILL_0__10790_ (
);

FILL FILL_0__10370_ (
);

FILL FILL_3__8718_ (
);

AOI21X1 _7862_ (
    .A(_1374_),
    .B(_1375_),
    .C(_1358_),
    .Y(_1376_)
);

NAND3X1 _7442_ (
    .A(vdd),
    .B(\X[1] [3]),
    .C(_961_),
    .Y(_962_)
);

NAND3X1 _7022_ (
    .A(_582_),
    .B(_584_),
    .C(_612_),
    .Y(_614_)
);

NAND2X1 _10499_ (
    .A(_3770_),
    .B(_3772_),
    .Y(_3773_)
);

OAI21X1 _10079_ (
    .A(_3357_),
    .B(_3358_),
    .C(_3356_),
    .Y(_3359_)
);

FILL FILL_2__6715_ (
);

FILL FILL_1__12582_ (
);

FILL FILL_3__11128_ (
);

FILL FILL_1__12162_ (
);

FILL FILL_0__11995_ (
);

FILL FILL_2__9187_ (
);

AOI21X1 _11860_ (
    .A(_4808_),
    .B(_4892_),
    .C(_4979_),
    .Y(_4980_)
);

FILL FILL_0__11575_ (
);

OAI21X1 _11440_ (
    .A(_4626_),
    .B(_4627_),
    .C(_4625_),
    .Y(_4628_)
);

FILL FILL_0__11155_ (
);

OAI21X1 _11020_ (
    .A(_4000_),
    .B(_4218_),
    .C(_4213_),
    .Y(_4219_)
);

FILL FILL_2__11902_ (
);

NAND2X1 _8647_ (
    .A(_2079_),
    .B(_2066_),
    .Y(_2083_)
);

INVX2 _8227_ (
    .A(\X[2]_5_bF$buf2 ),
    .Y(_1668_)
);

FILL FILL_1__7184_ (
);

FILL FILL_0__7902_ (
);

FILL FILL_3__8891_ (
);

AOI21X1 _12645_ (
    .A(_5607_),
    .B(_5627_),
    .C(_5641_),
    .Y(_5686_)
);

FILL FILL_3__8051_ (
);

NAND3X1 _12225_ (
    .A(_5236_),
    .B(_5338_),
    .C(_5079_),
    .Y(_5339_)
);

FILL FILL_0__13301_ (
);

FILL FILL_1__8389_ (
);

FILL FILL_2__10294_ (
);

FILL FILL_1__9750_ (
);

FILL FILL_1__9330_ (
);

FILL FILL_3__9676_ (
);

FILL FILL_2__7673_ (
);

FILL FILL_2__11499_ (
);

FILL FILL_2__11079_ (
);

INVX1 _6713_ (
    .A(_304_),
    .Y(_311_)
);

FILL FILL_2__12860_ (
);

FILL FILL_2__12440_ (
);

FILL FILL_2__12020_ (
);

FILL FILL_0__7499_ (
);

FILL FILL_0__7079_ (
);

AOI22X1 _9185_ (
    .A(gnd),
    .B(\X[3] [2]),
    .C(gnd),
    .D(\X[3] [3]),
    .Y(_2545_)
);

FILL FILL_1__11853_ (
);

FILL FILL_1__11433_ (
);

FILL FILL_1__11013_ (
);

FILL FILL_0__8860_ (
);

FILL FILL_2__8878_ (
);

FILL FILL_2__8458_ (
);

FILL FILL_0__8440_ (
);

FILL FILL_0__10846_ (
);

FILL FILL_0__10426_ (
);

DFFPOSX1 _10711_ (
    .D(_3978_[4]),
    .CLK(clk_bF$buf35),
    .Q(\Y[5] [4])
);

FILL FILL_2__8038_ (
);

FILL FILL_0__8020_ (
);

FILL FILL_0__10006_ (
);

INVX1 _13183_ (
    .A(\u_fir_pe7.mul [1]),
    .Y(_6212_)
);

INVX1 _7918_ (
    .A(_821_),
    .Y(_1588_[0])
);

FILL FILL_1__6875_ (
);

FILL FILL_1__6455_ (
);

FILL FILL_2__13225_ (
);

FILL FILL_1__12638_ (
);

FILL FILL_1__12218_ (
);

FILL FILL_0__9645_ (
);

NAND3X1 _11916_ (
    .A(_5028_),
    .B(_5031_),
    .C(_5029_),
    .Y(_5035_)
);

FILL FILL_0__9225_ (
);

FILL FILL_3__7322_ (
);

FILL FILL_3__10992_ (
);

FILL FILL_3__10572_ (
);

FILL FILL_3__10152_ (
);

FILL FILL_1__8601_ (
);

OAI21X1 _7671_ (
    .A(_1187_),
    .B(_1186_),
    .C(_1183_),
    .Y(_1188_)
);

DFFPOSX1 _7251_ (
    .D(_796_[12]),
    .CLK(clk_bF$buf34),
    .Q(\u_fir_pe0.mul [12])
);

FILL FILL_2__6944_ (
);

FILL FILL_3__11777_ (
);

FILL FILL_2__6524_ (
);

FILL FILL_3__11357_ (
);

FILL FILL_1__12391_ (
);

FILL FILL_0__11384_ (
);

FILL FILL_1__9806_ (
);

FILL FILL_2__11711_ (
);

INVX1 _8876_ (
    .A(_2297_),
    .Y(_2300_)
);

OAI21X1 _8456_ (
    .A(_1804_),
    .B(_1814_),
    .C(_1810_),
    .Y(_1894_)
);

INVX1 _8036_ (
    .A(\u_fir_pe1.mul [12]),
    .Y(_1540_)
);

FILL FILL_1__10704_ (
);

FILL FILL_0__7711_ (
);

FILL FILL_2__7729_ (
);

FILL FILL_2__7309_ (
);

FILL FILL_1__13176_ (
);

NAND2X1 _12874_ (
    .A(vdd),
    .B(\X[6] [6]),
    .Y(_5912_)
);

FILL FILL_0__12589_ (
);

FILL FILL_3__8280_ (
);

FILL FILL_0__12169_ (
);

NAND2X1 _12454_ (
    .A(_5556_),
    .B(_5557_),
    .Y(_5572_[15])
);

NAND3X1 _12034_ (
    .A(_5082_),
    .B(_5146_),
    .C(_5147_),
    .Y(_5152_)
);

FILL FILL_2__12916_ (
);

FILL FILL_0__13110_ (
);

FILL FILL_1__8198_ (
);

FILL FILL_1__11909_ (
);

FILL FILL_0__8916_ (
);

FILL FILL_3__9065_ (
);

NOR2X1 _13239_ (
    .A(_6260_),
    .B(_6261_),
    .Y(_6262_)
);

FILL FILL_2__7482_ (
);

FILL FILL_2__7062_ (
);

NAND2X1 _6942_ (
    .A(_536_),
    .B(_516_),
    .Y(_537_)
);

NAND3X1 _6522_ (
    .A(_54_),
    .B(_111_),
    .C(_115_),
    .Y(_123_)
);

FILL FILL_3__10628_ (
);

FILL FILL_1__11662_ (
);

FILL FILL_1__11242_ (
);

FILL FILL_2__8687_ (
);

FILL FILL_2__8267_ (
);

FILL FILL_0__10655_ (
);

OAI22X1 _10940_ (
    .A(_4027_),
    .B(_4138_),
    .C(_4070_),
    .D(_4139_),
    .Y(_4140_)
);

FILL FILL_0__10235_ (
);

NAND3X1 _10520_ (
    .A(_3766_),
    .B(_3768_),
    .C(_3792_),
    .Y(_3793_)
);

NAND3X1 _10100_ (
    .A(_3324_),
    .B(_3373_),
    .C(_3374_),
    .Y(_3380_)
);

AOI21X1 _7727_ (
    .A(_1243_),
    .B(_1242_),
    .C(_1235_),
    .Y(_1244_)
);

OAI22X1 _7307_ (
    .A(_827_),
    .B(_828_),
    .C(_797_),
    .D(_801_),
    .Y(_829_)
);

FILL FILL_1__6684_ (
);

FILL FILL_2__13034_ (
);

FILL FILL_1__12867_ (
);

FILL FILL_1__12447_ (
);

FILL FILL_1__12027_ (
);

FILL FILL_3__7971_ (
);

FILL FILL_0__9454_ (
);

FILL FILL_3__7551_ (
);

FILL FILL_0__9034_ (
);

AOI21X1 _11725_ (
    .A(_4843_),
    .B(_4846_),
    .C(_4837_),
    .Y(_4847_)
);

FILL FILL_3__7131_ (
);

NAND2X1 _11305_ (
    .A(_4453_),
    .B(_4454_),
    .Y(_4500_)
);

FILL FILL_0__12801_ (
);

FILL FILL_1__7889_ (
);

FILL FILL_1__7469_ (
);

FILL FILL_1__7049_ (
);

FILL FILL_1__8830_ (
);

FILL FILL_1__8410_ (
);

FILL FILL_3__8756_ (
);

FILL FILL_3__8336_ (
);

NAND2X1 _7480_ (
    .A(_999_),
    .B(_991_),
    .Y(_1000_)
);

AOI21X1 _7060_ (
    .A(_640_),
    .B(_645_),
    .C(_641_),
    .Y(_647_)
);

FILL FILL_2__6753_ (
);

FILL FILL_2__10999_ (
);

FILL FILL_2__10579_ (
);

FILL FILL_2__10159_ (
);

FILL FILL_0__11193_ (
);

FILL FILL_1__9615_ (
);

FILL FILL_2__11940_ (
);

FILL FILL_2__11520_ (
);

FILL FILL_0__6999_ (
);

FILL FILL_2__11100_ (
);

FILL FILL_0__6579_ (
);

NAND2X1 _8685_ (
    .A(gnd),
    .B(\X[2] [7]),
    .Y(_2120_)
);

INVX1 _8265_ (
    .A(_1620_),
    .Y(_1706_)
);

FILL FILL_1__10933_ (
);

FILL FILL_1__10513_ (
);

FILL FILL_0__7940_ (
);

FILL FILL_2__7958_ (
);

FILL FILL_0__7520_ (
);

FILL FILL_2__7538_ (
);

FILL FILL_2__7118_ (
);

FILL FILL_0__7100_ (
);

INVX2 _12683_ (
    .A(\X[6] [6]),
    .Y(_5723_)
);

FILL FILL_0__12398_ (
);

INVX1 _12263_ (
    .A(_5375_),
    .Y(_5376_)
);

FILL FILL_2__12725_ (
);

FILL FILL_2__12305_ (
);

FILL FILL_1__11718_ (
);

FILL FILL_0__8725_ (
);

FILL FILL_0__8305_ (
);

FILL FILL_3__6402_ (
);

FILL FILL_3__9294_ (
);

NOR2X1 _13048_ (
    .A(_6081_),
    .B(_6083_),
    .Y(_6084_)
);

FILL FILL_2__7291_ (
);

NAND3X1 _6751_ (
    .A(_342_),
    .B(_343_),
    .C(_344_),
    .Y(_349_)
);

FILL FILL_3__10857_ (
);

FILL FILL_1__11891_ (
);

FILL FILL_1__11471_ (
);

FILL FILL_3__10017_ (
);

FILL FILL_1__11051_ (
);

FILL FILL_2__8496_ (
);

FILL FILL_0__10884_ (
);

FILL FILL_0__10464_ (
);

FILL FILL_0__10044_ (
);

OAI21X1 _7956_ (
    .A(_1452_),
    .B(_1453_),
    .C(_1459_),
    .Y(_1461_)
);

AOI21X1 _7536_ (
    .A(_1048_),
    .B(_1054_),
    .C(_1035_),
    .Y(_1055_)
);

AOI21X1 _7116_ (
    .A(_695_),
    .B(_698_),
    .C(_697_),
    .Y(_699_)
);

FILL FILL_1__6493_ (
);

FILL FILL_2__13263_ (
);

FILL FILL_2__6809_ (
);

FILL FILL_1__12676_ (
);

FILL FILL_1__12256_ (
);

FILL FILL_0__9683_ (
);

FILL FILL_3__7780_ (
);

FILL FILL_0__9263_ (
);

NOR2X1 _11954_ (
    .A(_4989_),
    .B(_4986_),
    .Y(_5073_)
);

FILL FILL_0__11669_ (
);

AND2X2 _11534_ (
    .A(\u_fir_pe5.rYin [11]),
    .B(\u_fir_pe5.mul [11]),
    .Y(_4718_)
);

FILL FILL_0__11249_ (
);

AND2X2 _11114_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf3 ),
    .Y(_4312_)
);

FILL FILL_0__12610_ (
);

FILL FILL_1__7698_ (
);

FILL FILL_1__7278_ (
);

FILL FILL_3__10190_ (
);

AOI21X1 _12739_ (
    .A(_5761_),
    .B(_5756_),
    .C(_5763_),
    .Y(_5779_)
);

NOR2X1 _12319_ (
    .A(_5424_),
    .B(_5423_),
    .Y(_5427_)
);

FILL FILL_2__6982_ (
);

FILL FILL_2__6562_ (
);

FILL FILL_2__10388_ (
);

FILL FILL_1__9424_ (
);

FILL FILL_0__6388_ (
);

NAND3X1 _8494_ (
    .A(_1924_),
    .B(_1928_),
    .C(_1926_),
    .Y(_1932_)
);

NOR2X1 _8074_ (
    .A(_1517_),
    .B(_1581_),
    .Y(_1576_)
);

FILL FILL_1__10322_ (
);

FILL FILL_2__7767_ (
);

FILL FILL_2__7347_ (
);

DFFPOSX1 _12492_ (
    .D(\Y[7] [7]),
    .CLK(clk_bF$buf22),
    .Q(\u_fir_pe6.rYin [7])
);

NAND2X1 _12072_ (
    .A(_5188_),
    .B(_5185_),
    .Y(_5189_)
);

FILL FILL_3__13121_ (
);

AOI22X1 _6807_ (
    .A(gnd),
    .B(Xin[6]),
    .C(vdd),
    .D(Xin[7]),
    .Y(_404_)
);

FILL FILL_2__12954_ (
);

FILL FILL_2__12534_ (
);

FILL FILL_2__12114_ (
);

NAND2X1 _9699_ (
    .A(_3044_),
    .B(_3045_),
    .Y(_3181_[3])
);

NAND2X1 _9279_ (
    .A(_2549_),
    .B(_2633_),
    .Y(_2638_)
);

FILL FILL_1__11947_ (
);

FILL FILL_1__11527_ (
);

FILL FILL_1__11107_ (
);

FILL FILL_0__8534_ (
);

FILL FILL_3__6631_ (
);

AOI21X1 _10805_ (
    .A(_4004_),
    .B(_4005_),
    .C(_4771_),
    .Y(_4008_)
);

AOI21X1 _13277_ (
    .A(_6282_),
    .B(_6297_),
    .C(_6300_),
    .Y(_6301_)
);

FILL FILL_2__9913_ (
);

FILL FILL_1__6969_ (
);

FILL FILL_1__6549_ (
);

FILL FILL_2__13319_ (
);

FILL FILL_1__7910_ (
);

FILL FILL_0__9739_ (
);

FILL FILL_0__9319_ (
);

FILL FILL_3__7416_ (
);

INVX1 _6980_ (
    .A(_571_),
    .Y(_574_)
);

AOI22X1 _6560_ (
    .A(gnd),
    .B(Xin[3]),
    .C(vdd),
    .D(Xin[4]),
    .Y(_160_)
);

FILL FILL_3__10666_ (
);

FILL FILL_3__10246_ (
);

FILL FILL_1__11280_ (
);

FILL FILL_0__10693_ (
);

FILL FILL_0__10273_ (
);

FILL FILL_2__10600_ (
);

NAND2X1 _7765_ (
    .A(_1280_),
    .B(_1269_),
    .Y(_1281_)
);

OAI21X1 _7345_ (
    .A(_826_),
    .B(_860_),
    .C(_842_),
    .Y(_866_)
);

FILL FILL_2__13072_ (
);

FILL FILL_2__6618_ (
);

FILL FILL_0__6600_ (
);

FILL FILL_1__12065_ (
);

FILL FILL_0__9492_ (
);

FILL FILL_0__11898_ (
);

FILL FILL_0__9072_ (
);

NAND2X1 _11763_ (
    .A(_4863_),
    .B(_4859_),
    .Y(_4884_)
);

FILL FILL_0__11478_ (
);

FILL FILL_0__11058_ (
);

INVX1 _11343_ (
    .A(_4537_),
    .Y(_4538_)
);

FILL FILL_2__11805_ (
);

FILL FILL_1__7087_ (
);

FILL FILL_0__7805_ (
);

NAND3X1 _9911_ (
    .A(_3189_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3194_)
);

NAND3X1 _12968_ (
    .A(_5974_),
    .B(_6002_),
    .C(_6004_),
    .Y(_6005_)
);

FILL FILL_3__8374_ (
);

OAI21X1 _12548_ (
    .A(_5583_),
    .B(_5586_),
    .C(_5580_),
    .Y(_5591_)
);

INVX2 _12128_ (
    .A(gnd),
    .Y(_5244_)
);

FILL FILL_0__13204_ (
);

FILL FILL_2__6791_ (
);

FILL FILL_2__10197_ (
);

FILL FILL_1__9653_ (
);

FILL FILL_1__9233_ (
);

FILL FILL_3__9999_ (
);

FILL FILL_3__9159_ (
);

FILL FILL_1__10971_ (
);

FILL FILL_1__10551_ (
);

FILL FILL_1__10131_ (
);

FILL FILL_2__7996_ (
);

FILL FILL_2__7576_ (
);

FILL FILL_2__7156_ (
);

OAI21X1 _6616_ (
    .A(_139_),
    .B(_214_),
    .C(_143_),
    .Y(_215_)
);

FILL FILL_2__12763_ (
);

FILL FILL_2__12343_ (
);

OAI21X1 _9088_ (
    .A(_3172_),
    .B(_2409_),
    .C(_2412_),
    .Y(_2450_)
);

FILL FILL_1__11756_ (
);

FILL FILL_1__11336_ (
);

FILL FILL_0__8763_ (
);

FILL FILL_3__6860_ (
);

FILL FILL_0__8343_ (
);

FILL FILL_0__10329_ (
);

NAND2X1 _10614_ (
    .A(_3873_),
    .B(_3876_),
    .Y(_3978_[7])
);

NAND3X1 _13086_ (
    .A(_6094_),
    .B(_6120_),
    .C(_6116_),
    .Y(_6121_)
);

FILL FILL_2__9722_ (
);

FILL FILL_2__9302_ (
);

FILL FILL_1__6778_ (
);

FILL FILL_2__13128_ (
);

FILL FILL_0__9968_ (
);

FILL FILL_0__9548_ (
);

FILL FILL_3__7645_ (
);

FILL FILL_0__9128_ (
);

INVX1 _11819_ (
    .A(_4938_),
    .Y(_4939_)
);

FILL FILL_3__10475_ (
);

FILL FILL_0__10082_ (
);

FILL FILL_1__8924_ (
);

FILL FILL_1__8504_ (
);

AND2X2 _7994_ (
    .A(_1456_),
    .B(_1466_),
    .Y(_1498_)
);

NAND3X1 _7574_ (
    .A(_1082_),
    .B(_1085_),
    .C(_1001_),
    .Y(_1092_)
);

NOR2X1 _7154_ (
    .A(_736_),
    .B(_737_),
    .Y(_790_[11])
);

FILL FILL_2__6847_ (
);

FILL FILL_2__6427_ (
);

FILL FILL_1__12294_ (
);

OAI21X1 _11992_ (
    .A(_4871_),
    .B(_4926_),
    .C(_5109_),
    .Y(_5110_)
);

OR2X2 _11572_ (
    .A(\u_fir_pe5.rYin [15]),
    .B(\u_fir_pe5.mul [15]),
    .Y(_4756_)
);

FILL FILL_0__11287_ (
);

OAI21X1 _11152_ (
    .A(_4341_),
    .B(_4337_),
    .C(_4344_),
    .Y(_4350_)
);

FILL FILL_1__9709_ (
);

FILL FILL_3__12621_ (
);

FILL FILL_3__12201_ (
);

OAI21X1 _8779_ (
    .A(_2188_),
    .B(_2195_),
    .C(_2194_),
    .Y(_2211_)
);

OAI21X1 _8359_ (
    .A(_1723_),
    .B(_1721_),
    .C(_1714_),
    .Y(_1799_)
);

FILL FILL_1__10607_ (
);

FILL FILL_0__7614_ (
);

INVX1 _9720_ (
    .A(\u_fir_pe3.rYin [6]),
    .Y(_3064_)
);

NAND3X1 _9300_ (
    .A(_2657_),
    .B(_2658_),
    .C(_2656_),
    .Y(_2659_)
);

FILL FILL_1__13079_ (
);

NAND3X1 _12777_ (
    .A(_5804_),
    .B(_5813_),
    .C(_5815_),
    .Y(_5816_)
);

OR2X2 _12357_ (
    .A(_5454_),
    .B(_5459_),
    .Y(_5461_)
);

FILL FILL_2__12819_ (
);

FILL FILL_0__13013_ (
);

FILL FILL_0__8819_ (
);

FILL FILL_1__9462_ (
);

FILL FILL_1__9042_ (
);

FILL FILL_3__9388_ (
);

FILL FILL_1__10780_ (
);

FILL FILL_1__10360_ (
);

FILL FILL_2__7385_ (
);

NAND3X1 _6845_ (
    .A(_382_),
    .B(_437_),
    .C(_441_),
    .Y(_442_)
);

AOI22X1 _6425_ (
    .A(Xin[0]),
    .B(gnd),
    .C(gnd),
    .D(Xin[4]),
    .Y(_27_)
);

FILL FILL_2__12992_ (
);

FILL FILL_2__12572_ (
);

FILL FILL_2__12152_ (
);

FILL FILL_1__11985_ (
);

FILL FILL_1__11565_ (
);

FILL FILL_1__11145_ (
);

FILL FILL_0__8572_ (
);

FILL FILL_0__10978_ (
);

FILL FILL_0__8152_ (
);

FILL FILL_0__10558_ (
);

OR2X2 _10843_ (
    .A(_4044_),
    .B(_4043_),
    .Y(_4045_)
);

NOR2X1 _10423_ (
    .A(_3695_),
    .B(_3698_),
    .Y(_3984_[10])
);

FILL FILL_0__10138_ (
);

NAND3X1 _10003_ (
    .A(_3272_),
    .B(_3283_),
    .C(_3279_),
    .Y(_3284_)
);

FILL FILL_2__9951_ (
);

FILL FILL_2__9531_ (
);

FILL FILL_2__9111_ (
);

FILL FILL_1__6587_ (
);

FILL FILL_0__9777_ (
);

FILL FILL_3__7874_ (
);

FILL FILL_0__9357_ (
);

DFFPOSX1 _11628_ (
    .D(_4780_[4]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.mul [4])
);

NAND2X1 _11208_ (
    .A(_4388_),
    .B(_4398_),
    .Y(_4405_)
);

FILL FILL_0__12704_ (
);

FILL FILL254550x187350 (
);

FILL FILL_3__10284_ (
);

FILL FILL_1__8733_ (
);

FILL FILL_1__8313_ (
);

FILL FILL_3__8659_ (
);

AOI21X1 _7383_ (
    .A(_825_),
    .B(_845_),
    .C(_859_),
    .Y(_904_)
);

FILL FILL_3__9600_ (
);

FILL FILL_2__6656_ (
);

FILL FILL_3__11069_ (
);

NOR2X1 _11381_ (
    .A(_4574_),
    .B(_4573_),
    .Y(_4575_)
);

FILL FILL_0__11096_ (
);

FILL FILL_1__9938_ (
);

FILL FILL_1__9518_ (
);

FILL FILL_3__12430_ (
);

FILL FILL_2__11843_ (
);

FILL FILL_2__11423_ (
);

FILL FILL_2__11003_ (
);

NAND3X1 _8588_ (
    .A(_2020_),
    .B(_2024_),
    .C(_1979_),
    .Y(_2025_)
);

OAI21X1 _8168_ (
    .A(_2372_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1611_)
);

FILL FILL_1__10836_ (
);

FILL FILL_1__10416_ (
);

FILL FILL_0__7843_ (
);

FILL FILL_0__7423_ (
);

FILL FILL_0__7003_ (
);

NAND3X1 _12586_ (
    .A(_5608_),
    .B(_5624_),
    .C(_5627_),
    .Y(_5628_)
);

NAND2X1 _12166_ (
    .A(_5280_),
    .B(_5281_),
    .Y(_5282_)
);

FILL FILL_2__8802_ (
);

FILL FILL_3__13215_ (
);

FILL FILL_2__12628_ (
);

FILL FILL_2__12208_ (
);

FILL FILL_0__13242_ (
);

FILL FILL_0__8628_ (
);

FILL FILL_3__6725_ (
);

FILL FILL_0__8208_ (
);

FILL FILL_1__9691_ (
);

FILL FILL_1__9271_ (
);

FILL FILL_2__7194_ (
);

NAND3X1 _6654_ (
    .A(_246_),
    .B(_249_),
    .C(_247_),
    .Y(_253_)
);

FILL FILL_2__12381_ (
);

FILL FILL_1__11794_ (
);

FILL FILL_1__11374_ (
);

FILL FILL_0__8381_ (
);

FILL FILL_2__8399_ (
);

FILL FILL_0__10787_ (
);

NOR2X1 _10652_ (
    .A(_3915_),
    .B(_3914_),
    .Y(_3916_)
);

FILL FILL_0__10367_ (
);

OAI21X1 _10232_ (
    .A(_3506_),
    .B(_3509_),
    .C(_3508_),
    .Y(_3510_)
);

FILL FILL_3__11701_ (
);

FILL FILL_2__9760_ (
);

FILL FILL_2__9340_ (
);

NAND2X1 _7859_ (
    .A(_1369_),
    .B(_1372_),
    .Y(_1373_)
);

NAND3X1 _7439_ (
    .A(_954_),
    .B(_958_),
    .C(_956_),
    .Y(_959_)
);

AND2X2 _7019_ (
    .A(_608_),
    .B(_605_),
    .Y(_612_)
);

FILL FILL_1__6396_ (
);

FILL FILL_2__13166_ (
);

FILL FILL_1__12999_ (
);

NOR2X1 _8800_ (
    .A(\u_fir_pe2.rYin [1]),
    .B(\u_fir_pe2.mul [1]),
    .Y(_2229_)
);

FILL FILL_1__12579_ (
);

FILL FILL_1__12159_ (
);

FILL FILL_0__9586_ (
);

FILL FILL_0__9166_ (
);

AOI21X1 _11857_ (
    .A(_4900_),
    .B(_4899_),
    .C(_4836_),
    .Y(_4977_)
);

FILL FILL_3__7263_ (
);

OAI21X1 _11437_ (
    .A(_4617_),
    .B(_4618_),
    .C(_4622_),
    .Y(_4625_)
);

INVX1 _11017_ (
    .A(_4215_),
    .Y(_4216_)
);

FILL FILL_1__13100_ (
);

FILL FILL_0__12933_ (
);

FILL FILL_3__10093_ (
);

FILL FILL_1__8542_ (
);

NAND2X1 _7192_ (
    .A(_774_),
    .B(_775_),
    .Y(_790_[15])
);

FILL FILL_2__6885_ (
);

FILL FILL_2__6465_ (
);

FILL FILL_3__11298_ (
);

AOI22X1 _11190_ (
    .A(vdd),
    .B(\X[5]_5_bF$buf3 ),
    .C(gnd),
    .D(\X[5] [6]),
    .Y(_4387_)
);

FILL FILL_1__9747_ (
);

FILL FILL_1__9327_ (
);

FILL FILL_2__11652_ (
);

FILL FILL_2__11232_ (
);

AND2X2 _8397_ (
    .A(gnd),
    .B(\X[2]_5_bF$buf3 ),
    .Y(_1836_)
);

FILL FILL_1__10645_ (
);

FILL FILL_1__10225_ (
);

CLKBUF1 CLKBUF1_insert60 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert61 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert62 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert63 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert64 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf5)
);

FILL FILL_0__7652_ (
);

CLKBUF1 CLKBUF1_insert65 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert66 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert67 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert68 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert69 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf0)
);

OAI21X1 _12395_ (
    .A(_5494_),
    .B(_5495_),
    .C(_5493_),
    .Y(_5499_)
);

FILL FILL_2__8611_ (
);

FILL FILL_2__12857_ (
);

FILL FILL_2__12437_ (
);

FILL FILL_2__12017_ (
);

FILL FILL_0__13051_ (
);

FILL FILL_0__8857_ (
);

FILL FILL_3__6954_ (
);

FILL FILL_0__8437_ (
);

DFFPOSX1 _10708_ (
    .D(_3978_[1]),
    .CLK(clk_bF$buf6),
    .Q(\Y[5] [1])
);

FILL FILL_0__8017_ (
);

FILL FILL_1__9080_ (
);

FILL FILL_2__9816_ (
);

FILL FILL_1__7813_ (
);

FILL FILL_3__7739_ (
);

NAND2X1 _6883_ (
    .A(_477_),
    .B(_478_),
    .Y(_479_)
);

AOI21X1 _6463_ (
    .A(_61_),
    .B(_64_),
    .C(_55_),
    .Y(_65_)
);

FILL FILL_2__12190_ (
);

FILL FILL_3__10569_ (
);

FILL FILL_1__11183_ (
);

FILL FILL_0__8190_ (
);

FILL FILL_0__10596_ (
);

INVX1 _10881_ (
    .A(_4069_),
    .Y(_4082_)
);

NAND2X1 _10461_ (
    .A(_3735_),
    .B(_3702_),
    .Y(_3736_)
);

FILL FILL_0__10176_ (
);

OAI21X1 _10041_ (
    .A(_3898_),
    .B(_3320_),
    .C(_3265_),
    .Y(_3321_)
);

FILL FILL_3__11930_ (
);

FILL FILL_3__11510_ (
);

FILL FILL_2__10923_ (
);

FILL FILL_2__10503_ (
);

NAND2X1 _7668_ (
    .A(gnd),
    .B(_1184_),
    .Y(_1185_)
);

DFFPOSX1 _7248_ (
    .D(_796_[9]),
    .CLK(clk_bF$buf41),
    .Q(\u_fir_pe0.mul [9])
);

FILL FILL_2__13395_ (
);

FILL FILL_0__6923_ (
);

FILL FILL_0__6503_ (
);

FILL FILL_1__12388_ (
);

FILL FILL_0__9395_ (
);

FILL FILL_3__7492_ (
);

NOR2X1 _11666_ (
    .A(_5513_),
    .B(_4784_),
    .Y(_4789_)
);

FILL FILL_3__7072_ (
);

AOI21X1 _11246_ (
    .A(_4357_),
    .B(_4427_),
    .C(_4441_),
    .Y(_4442_)
);

FILL FILL_3__12715_ (
);

FILL FILL_2__11708_ (
);

FILL FILL_0__12742_ (
);

FILL FILL_0__12322_ (
);

FILL FILL_0__7708_ (
);

NOR2X1 _9814_ (
    .A(_3157_),
    .B(_3156_),
    .Y(_3181_[14])
);

FILL FILL_1__8771_ (
);

FILL FILL_1__8351_ (
);

FILL FILL_3__8697_ (
);

FILL FILL_3__8277_ (
);

FILL FILL_0__13107_ (
);

FILL FILL_2__6694_ (
);

FILL FILL_1__9976_ (
);

FILL FILL_1__9556_ (
);

FILL FILL_1__9136_ (
);

FILL FILL_2__11881_ (
);

FILL FILL_2__11461_ (
);

FILL FILL_2__11041_ (
);

FILL FILL_1__10874_ (
);

FILL FILL_1__10454_ (
);

FILL FILL_1__10034_ (
);

FILL FILL_2__7899_ (
);

FILL FILL_0__7881_ (
);

FILL FILL_2__7479_ (
);

FILL FILL_0__7461_ (
);

FILL FILL_2__7059_ (
);

FILL FILL_0__7041_ (
);

FILL FILL_2__8840_ (
);

FILL FILL_2__8420_ (
);

FILL FILL_2__8000_ (
);

INVX1 _6939_ (
    .A(_531_),
    .Y(_534_)
);

NAND3X1 _6519_ (
    .A(_116_),
    .B(_119_),
    .C(_68_),
    .Y(_120_)
);

FILL FILL_2__12666_ (
);

FILL FILL_2__12246_ (
);

FILL FILL_0__13280_ (
);

FILL FILL_1__11659_ (
);

FILL FILL_1__11239_ (
);

FILL FILL_0__8666_ (
);

FILL FILL_0__8246_ (
);

AND2X2 _10937_ (
    .A(_4132_),
    .B(_4136_),
    .Y(_4137_)
);

NAND2X1 _10517_ (
    .A(_3782_),
    .B(_3789_),
    .Y(_3790_)
);

FILL FILL_1__12600_ (
);

FILL FILL253950x79350 (
);

FILL FILL_2__9625_ (
);

FILL FILL_2__9205_ (
);

FILL FILL_1__7622_ (
);

FILL FILL_3__7968_ (
);

FILL FILL_3__7128_ (
);

NOR2X1 _6692_ (
    .A(_207_),
    .B(_204_),
    .Y(_291_)
);

FILL FILL_3__10798_ (
);

NOR2X1 _10690_ (
    .A(_3952_),
    .B(_3946_),
    .Y(_3954_)
);

NAND3X1 _10270_ (
    .A(_3541_),
    .B(_3542_),
    .C(_3543_),
    .Y(_3548_)
);

FILL FILL_1__8827_ (
);

FILL FILL_1__8407_ (
);

FILL FILL_2__10312_ (
);

NAND3X1 _7897_ (
    .A(_1381_),
    .B(_1409_),
    .C(_1408_),
    .Y(_1410_)
);

AOI21X1 _7477_ (
    .A(_979_),
    .B(_974_),
    .C(_981_),
    .Y(_997_)
);

NOR2X1 _7057_ (
    .A(_642_),
    .B(_641_),
    .Y(_645_)
);

FILL FILL_0__6732_ (
);

FILL FILL_1__12197_ (
);

NAND3X1 _11895_ (
    .A(_5008_),
    .B(_5013_),
    .C(_5011_),
    .Y(_5014_)
);

INVX1 _11475_ (
    .A(\u_fir_pe5.mul [6]),
    .Y(_4659_)
);

AOI21X1 _11055_ (
    .A(_4253_),
    .B(_4248_),
    .C(_4207_),
    .Y(_4254_)
);

FILL FILL_3__12944_ (
);

FILL FILL_2__11937_ (
);

FILL FILL_0__12971_ (
);

FILL FILL_2__11517_ (
);

FILL FILL_0__12551_ (
);

FILL FILL_0__12131_ (
);

FILL FILL_0__7937_ (
);

FILL FILL_0__7517_ (
);

AOI21X1 _9623_ (
    .A(_2948_),
    .B(_2950_),
    .C(_2976_),
    .Y(_2977_)
);

NAND3X1 _9203_ (
    .A(_2558_),
    .B(_2543_),
    .C(_2562_),
    .Y(_2563_)
);

FILL FILL_1__8580_ (
);

FILL FILL_1__8160_ (
);

FILL FILL_3__13309_ (
);

FILL FILL_0__13336_ (
);

INVX1 _13201_ (
    .A(\u_fir_pe7.mul [3]),
    .Y(_6228_)
);

FILL FILL_3__6819_ (
);

FILL FILL_1__9785_ (
);

FILL FILL_1__9365_ (
);

FILL FILL_2__11690_ (
);

FILL FILL_2__11270_ (
);

FILL FILL_1__10683_ (
);

FILL FILL_1__10263_ (
);

FILL FILL_0__7690_ (
);

FILL FILL_0__7270_ (
);

FILL FILL_2__7288_ (
);

FILL FILL_3__13062_ (
);

OAI21X1 _6748_ (
    .A(_341_),
    .B(_345_),
    .C(_317_),
    .Y(_346_)
);

FILL FILL_2__12895_ (
);

FILL FILL_2__12055_ (
);

FILL FILL_1__11888_ (
);

FILL FILL_1__11468_ (
);

FILL FILL_1__11048_ (
);

FILL FILL_0__8895_ (
);

FILL FILL_0__8475_ (
);

FILL FILL_3__6572_ (
);

DFFPOSX1 _10746_ (
    .D(\Y[4] [15]),
    .CLK(clk_bF$buf45),
    .Q(\u_fir_pe4.rYin [15])
);

FILL FILL_0__8055_ (
);

NAND3X1 _10326_ (
    .A(_3588_),
    .B(_3595_),
    .C(_3602_),
    .Y(_3603_)
);

FILL FILL_2__9434_ (
);

FILL FILL_0__11822_ (
);

FILL FILL_2__9014_ (
);

FILL FILL_0__11402_ (
);

FILL FILL_1__7851_ (
);

FILL FILL_1__7431_ (
);

FILL FILL_1__7011_ (
);

FILL FILL_3__7357_ (
);

FILL FILL_0__12607_ (
);

FILL FILL_3__10187_ (
);

FILL FILL_1__8636_ (
);

FILL FILL_1__8216_ (
);

FILL FILL_2__10961_ (
);

FILL FILL_2__10541_ (
);

FILL FILL_2__10121_ (
);

OAI21X1 _7286_ (
    .A(_801_),
    .B(_804_),
    .C(_798_),
    .Y(_809_)
);

FILL FILL_2__6979_ (
);

FILL FILL_0__6961_ (
);

FILL FILL_0__6541_ (
);

FILL FILL_2__6559_ (
);

NAND3X1 _11284_ (
    .A(_4445_),
    .B(_4479_),
    .C(_4477_),
    .Y(_4480_)
);

FILL FILL_2__7920_ (
);

FILL FILL_3__12753_ (
);

FILL FILL_2__7500_ (
);

FILL FILL_2__11746_ (
);

FILL FILL_0__12780_ (
);

FILL FILL_2__11326_ (
);

FILL FILL_0__12360_ (
);

FILL FILL_1__10319_ (
);

FILL FILL_0__7746_ (
);

DFFPOSX1 _9852_ (
    .D(\X[3] [6]),
    .CLK(clk_bF$buf42),
    .Q(\X[4] [6])
);

FILL FILL_0__7326_ (
);

NOR2X1 _9432_ (
    .A(_2523_),
    .B(_2712_),
    .Y(_2789_)
);

NOR2X1 _9012_ (
    .A(_3080_),
    .B(_3101_),
    .Y(_3111_)
);

DFFPOSX1 _12489_ (
    .D(\Y[7] [4]),
    .CLK(clk_bF$buf8),
    .Q(\u_fir_pe6.rYin [4])
);

AOI22X1 _12069_ (
    .A(gnd),
    .B(\X[7] [6]),
    .C(vdd),
    .D(\X[7] [7]),
    .Y(_5186_)
);

FILL FILL_2__8705_ (
);

FILL FILL_0__13145_ (
);

NOR2X1 _13010_ (
    .A(_5594_),
    .B(_6041_),
    .Y(_6046_)
);

FILL FILL_1__6702_ (
);

FILL FILL_3__6628_ (
);

FILL FILL_1__9594_ (
);

FILL FILL_1__9174_ (
);

FILL FILL_1__10492_ (
);

FILL FILL_1__10072_ (
);

FILL FILL_2__7097_ (
);

FILL FILL_1__7907_ (
);

NAND2X1 _6977_ (
    .A(_565_),
    .B(_569_),
    .Y(_571_)
);

INVX1 _6557_ (
    .A(_156_),
    .Y(_157_)
);

FILL FILL_2__12284_ (
);

FILL FILL_1__11697_ (
);

FILL FILL_1__11277_ (
);

FILL FILL_0__8284_ (
);

OAI21X1 _10975_ (
    .A(_4097_),
    .B(_4174_),
    .C(_4091_),
    .Y(_4175_)
);

NOR2X1 _10555_ (
    .A(_3823_),
    .B(_3822_),
    .Y(_3824_)
);

INVX1 _10135_ (
    .A(_3413_),
    .Y(_3414_)
);

FILL FILL_2__9663_ (
);

FILL FILL_2__9243_ (
);

FILL FILL_0__11211_ (
);

FILL FILL_2__13069_ (
);

NAND2X1 _8703_ (
    .A(_2134_),
    .B(_2110_),
    .Y(_2138_)
);

FILL FILL_1__7660_ (
);

FILL FILL_0__9489_ (
);

FILL FILL_3__7586_ (
);

FILL FILL_0__9069_ (
);

FILL FILL_3__7166_ (
);

FILL FILL_3__12809_ (
);

FILL FILL_1__13003_ (
);

FILL FILL_0__12836_ (
);

NAND3X1 _12701_ (
    .A(_5736_),
    .B(_5740_),
    .C(_5738_),
    .Y(_5741_)
);

FILL FILL_0__12416_ (
);

OR2X2 _9908_ (
    .A(_3919_),
    .B(_3190_),
    .Y(_3191_)
);

FILL FILL_1__8865_ (
);

FILL FILL_1__8445_ (
);

FILL FILL_1__8025_ (
);

FILL FILL_2__10770_ (
);

FILL FILL_2__10350_ (
);

OR2X2 _7095_ (
    .A(_672_),
    .B(_677_),
    .Y(_679_)
);

FILL FILL254550x50550 (
);

FILL FILL_3__9312_ (
);

FILL FILL253950x198150 (
);

FILL FILL_2__6788_ (
);

FILL FILL_0__6770_ (
);

NOR2X1 _11093_ (
    .A(_4755_),
    .B(_4290_),
    .Y(_4291_)
);

FILL FILL_3__12982_ (
);

FILL FILL_3__12562_ (
);

FILL FILL_3__12142_ (
);

FILL FILL_2__11975_ (
);

FILL FILL_2__11555_ (
);

FILL FILL_2__11135_ (
);

FILL FILL_1__10968_ (
);

FILL FILL_1__10548_ (
);

FILL FILL_1__10128_ (
);

FILL FILL_0__7975_ (
);

FILL FILL_0__7555_ (
);

OAI21X1 _9661_ (
    .A(_3007_),
    .B(_3006_),
    .C(_3012_),
    .Y(_3013_)
);

FILL FILL_0__7135_ (
);

OAI21X1 _9241_ (
    .A(_2527_),
    .B(_2599_),
    .C(_2568_),
    .Y(_2600_)
);

NAND3X1 _12298_ (
    .A(_5408_),
    .B(_5409_),
    .C(_5407_),
    .Y(_5410_)
);

FILL FILL_2__8934_ (
);

FILL FILL_2__8514_ (
);

FILL FILL_0__10902_ (
);

FILL FILL_1__6931_ (
);

FILL FILL_1__6511_ (
);

FILL FILL_3__6437_ (
);

FILL FILL_0__9701_ (
);

FILL FILL_2__9719_ (
);

FILL FILL_1__7716_ (
);

OAI21X1 _6786_ (
    .A(_304_),
    .B(_308_),
    .C(_313_),
    .Y(_383_)
);

FILL FILL_2__12093_ (
);

FILL FILL_1__11086_ (
);

FILL FILL_0__10499_ (
);

NAND2X1 _10784_ (
    .A(vdd),
    .B(\X[5] [0]),
    .Y(_3987_)
);

NAND2X1 _10364_ (
    .A(_3640_),
    .B(_3639_),
    .Y(_3984_[9])
);

FILL FILL_0__10079_ (
);

FILL FILL_3__11413_ (
);

FILL FILL_2__10826_ (
);

FILL FILL_2__9892_ (
);

FILL FILL_2__9472_ (
);

FILL FILL_0__11860_ (
);

FILL FILL_2__10406_ (
);

FILL FILL_2__9052_ (
);

FILL FILL_0__11440_ (
);

FILL FILL_0__11020_ (
);

FILL FILL_2__13298_ (
);

FILL FILL_0__6826_ (
);

NOR2X1 _8932_ (
    .A(_2353_),
    .B(_2355_),
    .Y(_2356_)
);

FILL FILL_0__6406_ (
);

AOI21X1 _8512_ (
    .A(_1949_),
    .B(_1948_),
    .C(_1947_),
    .Y(_1950_)
);

FILL FILL_0__9298_ (
);

NAND2X1 _11989_ (
    .A(gnd),
    .B(\X[7]_5_bF$buf3 ),
    .Y(_5107_)
);

INVX1 _11569_ (
    .A(_4747_),
    .Y(_4752_)
);

NAND3X1 _11149_ (
    .A(_4345_),
    .B(_4346_),
    .C(_4344_),
    .Y(_4347_)
);

FILL FILL_1__13232_ (
);

NAND2X1 _12930_ (
    .A(gnd),
    .B(_5966_),
    .Y(_5967_)
);

FILL FILL_0__12645_ (
);

FILL FILL_0__12225_ (
);

DFFPOSX1 _12510_ (
    .D(_5578_[9]),
    .CLK(clk_bF$buf22),
    .Q(\u_fir_pe6.mul [9])
);

OR2X2 _9717_ (
    .A(_3055_),
    .B(_3060_),
    .Y(_3062_)
);

FILL FILL_1__8674_ (
);

FILL FILL_1__8254_ (
);

FILL FILL_3__9961_ (
);

FILL FILL_3__9541_ (
);

FILL FILL_3__9121_ (
);

FILL FILL_2__6597_ (
);

FILL FILL_1__9459_ (
);

FILL FILL_1__9039_ (
);

FILL FILL_3__12371_ (
);

FILL FILL_2__11784_ (
);

FILL FILL_2__11364_ (
);

FILL FILL_1__10777_ (
);

FILL FILL_1__10357_ (
);

FILL FILL_0__7784_ (
);

NAND2X1 _9890_ (
    .A(gnd),
    .B(\X[4] [1]),
    .Y(_3919_)
);

FILL FILL_0__7364_ (
);

OAI21X1 _9470_ (
    .A(_2826_),
    .B(_2825_),
    .C(_2824_),
    .Y(_2827_)
);

INVX1 _9050_ (
    .A(_2412_),
    .Y(_2413_)
);

FILL FILL_2__8743_ (
);

FILL FILL_2__8323_ (
);

FILL FILL_3__13156_ (
);

FILL FILL_2__12989_ (
);

FILL FILL_2__12569_ (
);

FILL FILL_2__12149_ (
);

FILL FILL_0__13183_ (
);

FILL FILL_1__6740_ (
);

FILL FILL_0__8569_ (
);

FILL FILL_3__6666_ (
);

FILL FILL_0__8149_ (
);

FILL FILL_1__12923_ (
);

FILL FILL_0__9930_ (
);

FILL FILL_2__9948_ (
);

FILL FILL_2__9528_ (
);

FILL FILL_0__11916_ (
);

FILL FILL_0__9510_ (
);

FILL FILL_2__9108_ (
);

FILL FILL252750x248550 (
);

FILL FILL_1__7945_ (
);

FILL FILL_1__7525_ (
);

FILL FILL_1__7105_ (
);

AOI21X1 _6595_ (
    .A(_118_),
    .B(_117_),
    .C(_54_),
    .Y(_195_)
);

FILL FILL_3__8812_ (
);

NAND2X1 _10593_ (
    .A(_3857_),
    .B(_3852_),
    .Y(_3858_)
);

INVX1 _10173_ (
    .A(_3355_),
    .Y(_3452_)
);

FILL FILL_3__11642_ (
);

FILL FILL_3__11222_ (
);

FILL FILL_2__10635_ (
);

FILL FILL_2__9281_ (
);

FILL FILL_2__10215_ (
);

FILL FILL_0__6635_ (
);

INVX1 _8741_ (
    .A(_2174_),
    .Y(_2175_)
);

NAND3X1 _8321_ (
    .A(_1749_),
    .B(_1760_),
    .C(_1756_),
    .Y(_1761_)
);

NAND2X1 _11798_ (
    .A(_4917_),
    .B(_4916_),
    .Y(_4918_)
);

NAND3X1 _11378_ (
    .A(_4362_),
    .B(_4435_),
    .C(_4541_),
    .Y(_4572_)
);

FILL FILL_3__12007_ (
);

FILL FILL254250x7350 (
);

FILL FILL_1__13041_ (
);

FILL FILL_0__12874_ (
);

FILL FILL_0__12454_ (
);

FILL FILL_0__12034_ (
);

NAND3X1 _9946_ (
    .A(_3222_),
    .B(_3227_),
    .C(_3225_),
    .Y(_3228_)
);

NAND3X1 _9526_ (
    .A(_2879_),
    .B(_2881_),
    .C(_2880_),
    .Y(_2882_)
);

OAI21X1 _9106_ (
    .A(_3169_),
    .B(_2465_),
    .C(_2466_),
    .Y(_2467_)
);

FILL FILL_1__8483_ (
);

FILL FILL_1__8063_ (
);

FILL FILL_3__9770_ (
);

FILL FILL_0__13239_ (
);

AOI21X1 _13104_ (
    .A(_6135_),
    .B(_6036_),
    .C(_6137_),
    .Y(_6138_)
);

FILL FILL_1__9688_ (
);

FILL FILL_1__9268_ (
);

FILL FILL_2__11173_ (
);

FILL FILL_1__10586_ (
);

FILL FILL_1__10166_ (
);

FILL FILL_0__7593_ (
);

FILL FILL_0__7173_ (
);

FILL FILL_2__8552_ (
);

FILL FILL_0__10940_ (
);

FILL FILL_2__8132_ (
);

FILL FILL_0__10520_ (
);

FILL FILL_0__10100_ (
);

FILL FILL_2__12798_ (
);

FILL FILL_2__12378_ (
);

FILL FILL_0__8798_ (
);

FILL FILL_3__6895_ (
);

FILL FILL_0__8378_ (
);

INVX1 _10649_ (
    .A(\u_fir_pe4.mul [10]),
    .Y(_3913_)
);

INVX1 _10229_ (
    .A(vdd),
    .Y(_3507_)
);

FILL FILL_1__12732_ (
);

FILL FILL_1__12312_ (
);

FILL FILL_2__9757_ (
);

FILL FILL_2__9337_ (
);

FILL FILL_0__11725_ (
);

FILL FILL_0__11305_ (
);

FILL FILL_1__7754_ (
);

FILL FILL_1__7334_ (
);

FILL FILL_3__8201_ (
);

FILL FILL_3__11871_ (
);

FILL FILL_1__8539_ (
);

FILL FILL_3__11451_ (
);

FILL FILL_3__11031_ (
);

FILL FILL254250x244950 (
);

FILL FILL_2__10864_ (
);

FILL FILL_2__10444_ (
);

FILL FILL_2__9090_ (
);

FILL FILL_2__10024_ (
);

FILL FILL_1__9900_ (
);

INVX1 _7189_ (
    .A(_772_),
    .Y(_773_)
);

FILL FILL_0__6864_ (
);

DFFPOSX1 _8970_ (
    .D(\X[2] [1]),
    .CLK(clk_bF$buf28),
    .Q(\X[3] [1])
);

FILL FILL_0__6444_ (
);

INVX1 _8550_ (
    .A(_1984_),
    .Y(_1987_)
);

DFFPOSX1 _8130_ (
    .D(_1593_[14]),
    .CLK(clk_bF$buf13),
    .Q(\u_fir_pe1.mul [14])
);

AND2X2 _11187_ (
    .A(_4117_),
    .B(_4306_),
    .Y(_4384_)
);

FILL FILL_2__7823_ (
);

FILL FILL_3__12656_ (
);

FILL FILL_2__7403_ (
);

FILL FILL_3__12236_ (
);

FILL FILL_1__13270_ (
);

FILL FILL_2__11649_ (
);

FILL FILL_0__12683_ (
);

FILL FILL_2__11229_ (
);

FILL FILL_0__12263_ (
);

FILL FILL_0__7649_ (
);

NAND2X1 _9755_ (
    .A(_3095_),
    .B(_3098_),
    .Y(_3181_[8])
);

AOI21X1 _9335_ (
    .A(_2657_),
    .B(_2658_),
    .C(_2615_),
    .Y(_2693_)
);

FILL FILL_1__8292_ (
);

FILL FILL_2__8608_ (
);

FILL FILL_0__13048_ (
);

NOR2X1 _13333_ (
    .A(_6355_),
    .B(_6210_),
    .Y(_6368_[0])
);

FILL FILL_1__6605_ (
);

FILL FILL_1__9497_ (
);

FILL FILL_1__9077_ (
);

FILL FILL_1__10395_ (
);

FILL FILL_2__8781_ (
);

FILL FILL_2__8361_ (
);

FILL FILL_3__13194_ (
);

FILL FILL_2__12187_ (
);

AOI21X1 _7821_ (
    .A(_1267_),
    .B(_1283_),
    .C(_1335_),
    .Y(_1336_)
);

NAND3X1 _7401_ (
    .A(_920_),
    .B(_921_),
    .C(_919_),
    .Y(_922_)
);

FILL FILL_0__8187_ (
);

NAND3X1 _10878_ (
    .A(vdd),
    .B(\X[5] [2]),
    .C(_4078_),
    .Y(_4079_)
);

NAND2X1 _10458_ (
    .A(_3727_),
    .B(_3724_),
    .Y(_3733_)
);

AND2X2 _10038_ (
    .A(_3318_),
    .B(_3314_),
    .Y(_3984_[5])
);

FILL FILL_1__12961_ (
);

FILL FILL_3__11507_ (
);

FILL FILL_1__12541_ (
);

FILL FILL_1__12121_ (
);

FILL FILL_2__9986_ (
);

FILL FILL_2__9566_ (
);

FILL FILL_0__11954_ (
);

FILL FILL_2__9146_ (
);

FILL FILL_0__11534_ (
);

FILL FILL_0__11114_ (
);

OAI21X1 _8606_ (
    .A(_2041_),
    .B(_2042_),
    .C(_2038_),
    .Y(_2043_)
);

FILL FILL_1__7983_ (
);

FILL FILL_1__7563_ (
);

FILL FILL_1__7143_ (
);

FILL FILL_3__7069_ (
);

FILL FILL_1__13326_ (
);

FILL FILL_3__8850_ (
);

FILL FILL_0__12739_ (
);

FILL FILL_3__8430_ (
);

NAND2X1 _12604_ (
    .A(_5645_),
    .B(_5639_),
    .Y(_6374_[4])
);

FILL FILL_0__12319_ (
);

FILL FILL_3__8010_ (
);

FILL FILL_1__8768_ (
);

FILL FILL_1__8348_ (
);

FILL FILL_2__10673_ (
);

FILL FILL_2__10253_ (
);

FILL FILL_3__9635_ (
);

FILL FILL_3__9215_ (
);

FILL FILL_0__6673_ (
);

FILL FILL_2__7632_ (
);

FILL FILL_2__11878_ (
);

FILL FILL_2__11458_ (
);

FILL FILL_2__11038_ (
);

FILL FILL_0__12072_ (
);

FILL FILL_0__7878_ (
);

NAND3X1 _9984_ (
    .A(_3264_),
    .B(_3259_),
    .C(_3261_),
    .Y(_3265_)
);

FILL FILL_0__7458_ (
);

OAI21X1 _9564_ (
    .A(_2864_),
    .B(_2917_),
    .C(_2918_),
    .Y(_2919_)
);

FILL FILL_0__7038_ (
);

NAND3X1 _9144_ (
    .A(_2492_),
    .B(_2496_),
    .C(_2498_),
    .Y(_2505_)
);

FILL FILL_1__11812_ (
);

FILL FILL_2__8837_ (
);

FILL FILL_2__8417_ (
);

FILL FILL_0__10805_ (
);

FILL FILL_0__13277_ (
);

NAND2X1 _13142_ (
    .A(_6146_),
    .B(_6174_),
    .Y(_6175_)
);

FILL FILL_1__6834_ (
);

FILL FILL_1__6414_ (
);

FILL FILL_0__9604_ (
);

FILL FILL_3__10951_ (
);

FILL FILL_1__7619_ (
);

FILL FILL_3__10111_ (
);

FILL FILL_2__8590_ (
);

FILL FILL_2__8170_ (
);

NAND3X1 _6689_ (
    .A(_188_),
    .B(_286_),
    .C(_287_),
    .Y(_288_)
);

FILL FILL_3__8906_ (
);

NAND3X1 _7630_ (
    .A(_1146_),
    .B(_1147_),
    .C(_1145_),
    .Y(_1148_)
);

DFFPOSX1 _7210_ (
    .D(_790_[11]),
    .CLK(clk_bF$buf54),
    .Q(\Y[1] [11])
);

NOR2X1 _10687_ (
    .A(\u_fir_pe4.rYin [14]),
    .B(\u_fir_pe4.mul [14]),
    .Y(_3951_)
);

OAI21X1 _10267_ (
    .A(_3544_),
    .B(_3540_),
    .C(_3491_),
    .Y(_3545_)
);

FILL FILL_2__6903_ (
);

FILL FILL_3__11736_ (
);

FILL FILL_1__12770_ (
);

FILL FILL_1__12350_ (
);

FILL FILL_2__9795_ (
);

FILL FILL_2__9375_ (
);

FILL FILL_0__11763_ (
);

FILL FILL_2__10309_ (
);

FILL FILL_0__11343_ (
);

FILL FILL_0__6729_ (
);

INVX1 _8835_ (
    .A(\u_fir_pe2.mul [5]),
    .Y(_2260_)
);

NAND3X1 _8415_ (
    .A(_1833_),
    .B(_1847_),
    .C(_1850_),
    .Y(_1854_)
);

FILL FILL_1__7792_ (
);

FILL FILL_1__7372_ (
);

FILL FILL_3__7298_ (
);

FILL FILL_1__13135_ (
);

FILL FILL_0__12968_ (
);

INVX1 _12833_ (
    .A(_5867_),
    .Y(_5872_)
);

FILL FILL_0__12548_ (
);

FILL FILL_0__12128_ (
);

NOR2X1 _12413_ (
    .A(_5516_),
    .B(_5515_),
    .Y(_5517_)
);

FILL FILL_1__8577_ (
);

FILL FILL_1__8157_ (
);

FILL FILL_2__10482_ (
);

FILL FILL_2__10062_ (
);

FILL FILL254250x79350 (
);

FILL FILL_0__6482_ (
);

FILL FILL_2__7861_ (
);

FILL FILL_3__12694_ (
);

FILL FILL_2__7441_ (
);

FILL FILL_2__7021_ (
);

FILL FILL_2__11687_ (
);

FILL FILL_2__11267_ (
);

NAND2X1 _6901_ (
    .A(_493_),
    .B(_461_),
    .Y(_497_)
);

FILL FILL_0__7687_ (
);

NOR2X1 _9793_ (
    .A(_3136_),
    .B(_3135_),
    .Y(_3137_)
);

FILL FILL_0__7267_ (
);

NAND3X1 _9373_ (
    .A(_2729_),
    .B(_2730_),
    .C(_2728_),
    .Y(_2731_)
);

FILL FILL_1__11201_ (
);

FILL FILL_2__8646_ (
);

FILL FILL_2__8226_ (
);

FILL FILL_0__10614_ (
);

FILL FILL_0__13086_ (
);

DFFPOSX1 _13371_ (
    .D(\Y[6] [9]),
    .CLK(clk_bF$buf5),
    .Q(\u_fir_pe7.rYin [9])
);

FILL FILL_1__6643_ (
);

FILL FILL_2__13413_ (
);

FILL FILL_3__6989_ (
);

FILL FILL_1__12826_ (
);

FILL FILL_1__12406_ (
);

FILL FILL_0__9413_ (
);

FILL FILL_0__11819_ (
);

FILL FILL_3__7510_ (
);

FILL FILL254550x223350 (
);

FILL FILL_1__7848_ (
);

FILL FILL_1__7428_ (
);

FILL FILL_3__10340_ (
);

FILL FILL_1__7008_ (
);

AOI22X1 _6498_ (
    .A(gnd),
    .B(Xin[4]),
    .C(_88_),
    .D(_90_),
    .Y(_99_)
);

OAI21X1 _10496_ (
    .A(_3767_),
    .B(_3769_),
    .C(_3748_),
    .Y(_3770_)
);

INVX1 _10076_ (
    .A(_3343_),
    .Y(_3356_)
);

FILL FILL_3__11965_ (
);

FILL FILL_2__6712_ (
);

FILL FILL_3__11545_ (
);

FILL FILL_3__11125_ (
);

FILL FILL_2__10958_ (
);

FILL FILL_0__11992_ (
);

FILL FILL_2__10538_ (
);

FILL FILL_2__9184_ (
);

FILL FILL_0__11572_ (
);

FILL FILL_2__10118_ (
);

FILL FILL_0__11152_ (
);

FILL FILL_0__6958_ (
);

FILL FILL_0__6538_ (
);

NAND3X1 _8644_ (
    .A(_2001_),
    .B(_2079_),
    .C(_2009_),
    .Y(_2080_)
);

INVX1 _8224_ (
    .A(_1664_),
    .Y(_1665_)
);

FILL FILL_1__7181_ (
);

FILL FILL_2__7917_ (
);

FILL FILL_0__12777_ (
);

NAND3X1 _12642_ (
    .A(_5674_),
    .B(_5670_),
    .C(_5676_),
    .Y(_5683_)
);

FILL FILL_0__12357_ (
);

OAI21X1 _12222_ (
    .A(_5286_),
    .B(_5289_),
    .C(_5334_),
    .Y(_5337_)
);

DFFPOSX1 _9849_ (
    .D(\X[3] [3]),
    .CLK(clk_bF$buf15),
    .Q(\X[4] [3])
);

AND2X2 _9429_ (
    .A(_2785_),
    .B(_2782_),
    .Y(_2786_)
);

NAND2X1 _9009_ (
    .A(\X[3] [0]),
    .B(vdd),
    .Y(_3080_)
);

FILL FILL_1__8386_ (
);

FILL FILL_2__10291_ (
);

FILL FILL_3__9253_ (
);

OAI22X1 _13007_ (
    .A(_5996_),
    .B(_5884_),
    .C(_5604_),
    .D(_5995_),
    .Y(_6043_)
);

FILL FILL_2__7670_ (
);

FILL FILL_3__12083_ (
);

FILL FILL_2__11496_ (
);

FILL FILL_2__11076_ (
);

NOR2X1 _6710_ (
    .A(_306_),
    .B(_307_),
    .Y(_308_)
);

FILL FILL_1__10489_ (
);

FILL FILL_1__10069_ (
);

FILL FILL_0__7496_ (
);

FILL FILL_0__7076_ (
);

NAND3X1 _9182_ (
    .A(_2530_),
    .B(_2539_),
    .C(_2541_),
    .Y(_2542_)
);

FILL FILL_1__11850_ (
);

FILL FILL_1__11430_ (
);

FILL FILL_1__11010_ (
);

FILL FILL_2__8875_ (
);

FILL FILL_2__8455_ (
);

FILL FILL_0__10843_ (
);

FILL FILL_0__10423_ (
);

FILL FILL_2__8035_ (
);

FILL FILL_0__10003_ (
);

INVX1 _13180_ (
    .A(_5603_),
    .Y(_6370_[0])
);

OAI21X1 _7915_ (
    .A(_1413_),
    .B(_1412_),
    .C(_1424_),
    .Y(_1426_)
);

FILL FILL_1__6872_ (
);

FILL FILL_1__6452_ (
);

FILL FILL_2__13222_ (
);

FILL FILL_3__6378_ (
);

FILL FILL_1__12635_ (
);

FILL FILL_1__12215_ (
);

FILL FILL_0__9642_ (
);

FILL FILL_0__9222_ (
);

AOI21X1 _11913_ (
    .A(_5029_),
    .B(_5031_),
    .C(_5028_),
    .Y(_5032_)
);

FILL FILL_0__11208_ (
);

FILL FILL_1__7657_ (
);

FILL FILL_3__8524_ (
);

FILL FILL_2__6941_ (
);

FILL FILL_2__6521_ (
);

FILL FILL_3__11354_ (
);

FILL FILL_2__10767_ (
);

FILL FILL_2__10347_ (
);

FILL FILL_0__11381_ (
);

FILL FILL_1__9803_ (
);

FILL FILL_3__9729_ (
);

FILL FILL_3__9309_ (
);

FILL FILL_0__6767_ (
);

NAND2X1 _8873_ (
    .A(_2293_),
    .B(_2296_),
    .Y(_2297_)
);

NAND2X1 _8453_ (
    .A(_1890_),
    .B(_1889_),
    .Y(_1891_)
);

NAND2X1 _8033_ (
    .A(_1532_),
    .B(_1525_),
    .Y(_1536_)
);

FILL FILL_1__10701_ (
);

FILL FILL_3__12979_ (
);

FILL FILL_2__7726_ (
);

FILL FILL_2__7306_ (
);

FILL FILL_1__13173_ (
);

INVX1 _12871_ (
    .A(_5903_),
    .Y(_5909_)
);

FILL FILL_0__12586_ (
);

FILL FILL_0__12166_ (
);

INVX1 _12451_ (
    .A(_5554_),
    .Y(_5555_)
);

OAI21X1 _12031_ (
    .A(_5148_),
    .B(_5145_),
    .C(_5081_),
    .Y(_5149_)
);

FILL FILL_2__12913_ (
);

OR2X2 _9658_ (
    .A(_3008_),
    .B(_3009_),
    .Y(_3010_)
);

NOR2X1 _9238_ (
    .A(_2595_),
    .B(_2597_),
    .Y(_3187_[6])
);

FILL FILL_1__8195_ (
);

FILL FILL_1__11906_ (
);

FILL FILL_0__8913_ (
);

FILL FILL_3__9482_ (
);

OAI21X1 _13236_ (
    .A(_6252_),
    .B(_6253_),
    .C(_6257_),
    .Y(_6259_)
);

FILL FILL_1__6928_ (
);

FILL FILL_1__6508_ (
);

FILL FILL_1__10298_ (
);

FILL FILL_3__10205_ (
);

FILL FILL_2__8684_ (
);

FILL FILL_2__8264_ (
);

FILL FILL_0__10652_ (
);

FILL FILL_3__13097_ (
);

FILL FILL_0__10232_ (
);

AOI21X1 _7724_ (
    .A(_1097_),
    .B(_1162_),
    .C(_1240_),
    .Y(_1241_)
);

INVX1 _7304_ (
    .A(_825_),
    .Y(_826_)
);

FILL FILL_1__6681_ (
);

FILL FILL_2__13031_ (
);

FILL FILL_1__12864_ (
);

FILL FILL_1__12444_ (
);

FILL FILL_1__12024_ (
);

FILL FILL_2__9889_ (
);

FILL FILL_2__9469_ (
);

FILL FILL_0__9451_ (
);

FILL FILL_0__11857_ (
);

FILL FILL_0__9031_ (
);

FILL FILL_2__9049_ (
);

INVX1 _11722_ (
    .A(_4827_),
    .Y(_4844_)
);

FILL FILL_0__11437_ (
);

NAND2X1 _11302_ (
    .A(_4490_),
    .B(_4494_),
    .Y(_4497_)
);

FILL FILL_0__11017_ (
);

OAI21X1 _8929_ (
    .A(_2345_),
    .B(_2346_),
    .C(_2350_),
    .Y(_2352_)
);

AND2X2 _8509_ (
    .A(_1908_),
    .B(_1904_),
    .Y(_1947_)
);

FILL FILL_1__7886_ (
);

FILL FILL_1__7466_ (
);

FILL FILL_1__7046_ (
);

FILL FILL_1__13229_ (
);

FILL FILL_3__8753_ (
);

OAI21X1 _12927_ (
    .A(_5894_),
    .B(_5963_),
    .C(_5933_),
    .Y(_5964_)
);

DFFPOSX1 _12507_ (
    .D(_5578_[6]),
    .CLK(clk_bF$buf29),
    .Q(\u_fir_pe6.mul [6])
);

FILL FILL_2__6750_ (
);

FILL FILL_3__11163_ (
);

FILL FILL_2__10996_ (
);

FILL FILL_2__10576_ (
);

FILL FILL_2__10156_ (
);

FILL FILL_0__11190_ (
);

FILL FILL_1__9612_ (
);

FILL FILL_3__9538_ (
);

FILL FILL_0__6996_ (
);

FILL FILL_0__6576_ (
);

NAND3X1 _8682_ (
    .A(_2114_),
    .B(_2115_),
    .C(_2116_),
    .Y(_2117_)
);

AOI21X1 _8262_ (
    .A(_1694_),
    .B(_1690_),
    .C(_1676_),
    .Y(_1703_)
);

FILL FILL_1__10930_ (
);

FILL FILL_1__10510_ (
);

FILL FILL_2__7955_ (
);

FILL FILL_2__7535_ (
);

FILL FILL_2__7115_ (
);

AND2X2 _12680_ (
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5720_)
);

FILL FILL_0__12395_ (
);

NOR2X1 _12260_ (
    .A(_5342_),
    .B(_5365_),
    .Y(_5373_)
);

FILL FILL_2__12722_ (
);

FILL FILL_2__12302_ (
);

AND2X2 _9887_ (
    .A(\X[4] [1]),
    .B(gnd),
    .Y(_3888_)
);

AOI21X1 _9467_ (
    .A(_2744_),
    .B(_2746_),
    .C(_2823_),
    .Y(_2824_)
);

NAND2X1 _9047_ (
    .A(_3172_),
    .B(_2409_),
    .Y(_2410_)
);

FILL FILL_1__11715_ (
);

FILL FILL_0__8722_ (
);

FILL FILL_0__8302_ (
);

AOI21X1 _13045_ (
    .A(_6074_),
    .B(_6080_),
    .C(_6038_),
    .Y(_6081_)
);

FILL FILL_1__6737_ (
);

FILL FILL_0__9927_ (
);

FILL FILL_0__9507_ (
);

FILL FILL_3__7604_ (
);

FILL FILL_3__10434_ (
);

FILL FILL_2__8493_ (
);

FILL FILL_0__10881_ (
);

FILL FILL_0__10461_ (
);

FILL FILL_2__8073_ (
);

FILL FILL_0__10041_ (
);

NAND2X1 _7953_ (
    .A(_1456_),
    .B(_1458_),
    .Y(_1459_)
);

NOR2X1 _7533_ (
    .A(_1038_),
    .B(_1051_),
    .Y(_1052_)
);

NAND2X1 _7113_ (
    .A(_675_),
    .B(_687_),
    .Y(_696_)
);

FILL FILL_1__6490_ (
);

FILL FILL_2__13260_ (
);

FILL FILL_2__6806_ (
);

FILL FILL_1__12673_ (
);

FILL FILL_3__11219_ (
);

FILL FILL_1__12253_ (
);

FILL FILL_0__9680_ (
);

FILL FILL_2__9698_ (
);

FILL FILL_2__9278_ (
);

FILL FILL_0__9260_ (
);

NAND3X1 _11951_ (
    .A(_4970_),
    .B(_5068_),
    .C(_5069_),
    .Y(_5070_)
);

FILL FILL_0__11666_ (
);

OAI21X1 _11531_ (
    .A(_4711_),
    .B(_4712_),
    .C(_4707_),
    .Y(_4715_)
);

FILL FILL_0__11246_ (
);

NAND2X1 _11111_ (
    .A(gnd),
    .B(\X[5] [7]),
    .Y(_4309_)
);

NAND3X1 _8738_ (
    .A(_2156_),
    .B(_2166_),
    .C(_2169_),
    .Y(_2172_)
);

NAND2X1 _8318_ (
    .A(gnd),
    .B(\X[2] [4]),
    .Y(_1758_)
);

FILL FILL_1__7695_ (
);

FILL FILL_1__7275_ (
);

FILL FILL_1__13038_ (
);

INVX1 _12736_ (
    .A(_5685_),
    .Y(_5776_)
);

FILL FILL_3__8142_ (
);

NOR2X1 _12316_ (
    .A(\u_fir_pe6.rYin [2]),
    .B(\u_fir_pe6.mul [2]),
    .Y(_5424_)
);

FILL FILL_3__11392_ (
);

FILL FILL_2__10385_ (
);

FILL FILL_1__9421_ (
);

FILL FILL_3__9347_ (
);

FILL FILL_0__6385_ (
);

AOI21X1 _8491_ (
    .A(_1926_),
    .B(_1928_),
    .C(_1924_),
    .Y(_1929_)
);

NOR2X1 _8071_ (
    .A(_1573_),
    .B(_1428_),
    .Y(_1586_[0])
);

FILL FILL_2__7764_ (
);

FILL FILL_3__12597_ (
);

FILL FILL_2__7344_ (
);

FILL FILL_3__12177_ (
);

NAND2X1 _6804_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_401_)
);

FILL FILL_2__12951_ (
);

FILL FILL_2__12531_ (
);

FILL FILL_2__12111_ (
);

NOR2X1 _9696_ (
    .A(_3042_),
    .B(_3041_),
    .Y(_3043_)
);

OAI21X1 _9276_ (
    .A(_2480_),
    .B(_2465_),
    .C(_2549_),
    .Y(_2635_)
);

FILL FILL_1__11944_ (
);

FILL FILL_1__11524_ (
);

FILL FILL_1__11104_ (
);

FILL FILL_0__8951_ (
);

FILL FILL_2__8549_ (
);

FILL FILL_0__8531_ (
);

FILL FILL_0__10937_ (
);

FILL FILL_0__10517_ (
);

NAND3X1 _10802_ (
    .A(_4767_),
    .B(_3999_),
    .C(_4002_),
    .Y(_4005_)
);

NOR2X1 _13274_ (
    .A(_6294_),
    .B(_6288_),
    .Y(_6297_)
);

FILL FILL_2__9910_ (
);

FILL FILL_1__6966_ (
);

FILL FILL_1__6546_ (
);

FILL FILL_2__13316_ (
);

FILL FILL_1__12729_ (
);

FILL FILL_1__12309_ (
);

FILL FILL_0__9736_ (
);

FILL FILL_3__7833_ (
);

FILL FILL_0__9316_ (
);

FILL FILL_3__10663_ (
);

FILL FILL_0__10690_ (
);

FILL FILL_0__10270_ (
);

FILL FILL_3__8618_ (
);

AOI21X1 _7762_ (
    .A(vdd),
    .B(\X[1] [6]),
    .C(_1209_),
    .Y(_1278_)
);

NAND2X1 _7342_ (
    .A(_863_),
    .B(_857_),
    .Y(_1592_[4])
);

NAND3X1 _10399_ (
    .A(_3658_),
    .B(_3674_),
    .C(_3672_),
    .Y(_3675_)
);

FILL FILL_2__6615_ (
);

FILL FILL_3__11448_ (
);

FILL FILL_1__12062_ (
);

FILL FILL_0__11895_ (
);

FILL FILL_2__9087_ (
);

AOI22X1 _11760_ (
    .A(gnd),
    .B(\X[7] [4]),
    .C(_4870_),
    .D(_4872_),
    .Y(_4881_)
);

FILL FILL_0__11475_ (
);

FILL FILL_0__11055_ (
);

OAI21X1 _11340_ (
    .A(_4481_),
    .B(_4534_),
    .C(_4477_),
    .Y(_4535_)
);

FILL FILL_2__11802_ (
);

DFFPOSX1 _8967_ (
    .D(_2384_[14]),
    .CLK(clk_bF$buf36),
    .Q(\Y[3] [14])
);

AOI21X1 _8547_ (
    .A(\X[2] [3]),
    .B(gnd),
    .C(_1981_),
    .Y(_1984_)
);

DFFPOSX1 _8127_ (
    .D(_1593_[11]),
    .CLK(clk_bF$buf32),
    .Q(\u_fir_pe1.mul [11])
);

FILL FILL_1__7084_ (
);

FILL FILL_0__7802_ (
);

FILL FILL_1__13267_ (
);

FILL FILL_3__8791_ (
);

NAND3X1 _12965_ (
    .A(_5994_),
    .B(_6001_),
    .C(_5976_),
    .Y(_6002_)
);

FILL FILL_3__8371_ (
);

NAND3X1 _12545_ (
    .A(_6319_),
    .B(_5587_),
    .C(_5585_),
    .Y(_5588_)
);

OAI21X1 _12125_ (
    .A(_5220_),
    .B(_5222_),
    .C(_5213_),
    .Y(_5241_)
);

FILL FILL_0__13201_ (
);

FILL FILL_1__8289_ (
);

FILL FILL_2__10194_ (
);

FILL FILL_1__9650_ (
);

FILL FILL_1__9230_ (
);

FILL FILL_3__9996_ (
);

FILL FILL_3__9576_ (
);

FILL FILL_3__9156_ (
);

FILL FILL_2__7993_ (
);

FILL FILL_2__7573_ (
);

FILL FILL_2__7153_ (
);

FILL FILL_2__11399_ (
);

NAND2X1 _6613_ (
    .A(Xin[1]),
    .B(gnd),
    .Y(_212_)
);

FILL FILL_2__12760_ (
);

FILL FILL_2__12340_ (
);

FILL FILL_0__7399_ (
);

NAND2X1 _9085_ (
    .A(_2440_),
    .B(_2443_),
    .Y(_2447_)
);

FILL FILL_1__11753_ (
);

FILL FILL_1__11333_ (
);

FILL FILL_0__8760_ (
);

FILL FILL_2__8778_ (
);

FILL FILL_0__8340_ (
);

FILL FILL_2__8358_ (
);

FILL FILL_0__10326_ (
);

INVX1 _10611_ (
    .A(_3868_),
    .Y(_3874_)
);

AOI21X1 _13083_ (
    .A(_6049_),
    .B(_6065_),
    .C(_6117_),
    .Y(_6118_)
);

AND2X2 _7818_ (
    .A(_1332_),
    .B(_1329_),
    .Y(_1333_)
);

FILL FILL_1__6775_ (
);

FILL FILL_2__13125_ (
);

FILL FILL_1__12958_ (
);

FILL FILL_1__12538_ (
);

FILL FILL_1__12118_ (
);

FILL FILL_0__9965_ (
);

FILL FILL_0__9545_ (
);

FILL FILL_0__9125_ (
);

AOI22X1 _11816_ (
    .A(gnd),
    .B(\X[7] [2]),
    .C(vdd),
    .D(\X[7] [3]),
    .Y(_4936_)
);

FILL FILL_3__10892_ (
);

FILL FILL_3__10052_ (
);

FILL FILL_1__8921_ (
);

FILL FILL_1__8501_ (
);

FILL FILL_3__8847_ (
);

FILL FILL_3__8007_ (
);

OAI21X1 _7991_ (
    .A(_1478_),
    .B(_1479_),
    .C(_1493_),
    .Y(_1494_)
);

INVX1 _7571_ (
    .A(_1085_),
    .Y(_1090_)
);

NOR2X1 _7151_ (
    .A(_734_),
    .B(_733_),
    .Y(_735_)
);

FILL FILL_2__6844_ (
);

FILL FILL_3__11677_ (
);

FILL FILL_2__6424_ (
);

FILL FILL_1__12291_ (
);

FILL FILL_0__11284_ (
);

FILL FILL_1__9706_ (
);

NAND3X1 _8776_ (
    .A(_2176_),
    .B(_2178_),
    .C(_2206_),
    .Y(_2208_)
);

NAND3X1 _8356_ (
    .A(_1789_),
    .B(_1790_),
    .C(_1795_),
    .Y(_1796_)
);

FILL FILL_1__10604_ (
);

FILL FILL_0__7611_ (
);

FILL FILL_2__7629_ (
);

FILL FILL_1__13076_ (
);

OAI21X1 _12774_ (
    .A(_5594_),
    .B(_5812_),
    .C(_5807_),
    .Y(_5813_)
);

FILL FILL_0__12069_ (
);

NOR2X1 _12354_ (
    .A(\u_fir_pe6.rYin [6]),
    .B(\u_fir_pe6.mul [6]),
    .Y(_5458_)
);

FILL FILL_2__12816_ (
);

FILL FILL_0__13010_ (
);

FILL FILL_1__11809_ (
);

FILL FILL_0__8816_ (
);

OAI21X1 _13139_ (
    .A(_5884_),
    .B(_6171_),
    .C(_6150_),
    .Y(_6172_)
);

FILL FILL_2__7382_ (
);

INVX1 _6842_ (
    .A(_431_),
    .Y(_439_)
);

NAND2X1 _6422_ (
    .A(Xin[0]),
    .B(gnd),
    .Y(_24_)
);

FILL FILL_3__10948_ (
);

FILL FILL_1__11982_ (
);

FILL FILL_3__10528_ (
);

FILL FILL_1__11562_ (
);

FILL FILL_1__11142_ (
);

FILL FILL_2__8587_ (
);

FILL FILL_0__10975_ (
);

FILL FILL_2__8167_ (
);

FILL FILL_0__10555_ (
);

OR2X2 _10840_ (
    .A(_4041_),
    .B(_4040_),
    .Y(_4042_)
);

NAND2X1 _10420_ (
    .A(_3565_),
    .B(_3638_),
    .Y(_3696_)
);

FILL FILL_0__10135_ (
);

NAND2X1 _10000_ (
    .A(gnd),
    .B(\X[4] [3]),
    .Y(_3281_)
);

AOI21X1 _7627_ (
    .A(_1056_),
    .B(_1058_),
    .C(_1144_),
    .Y(_1145_)
);

DFFPOSX1 _7207_ (
    .D(_790_[8]),
    .CLK(clk_bF$buf16),
    .Q(\Y[1] [8])
);

FILL FILL_1__6584_ (
);

FILL FILL_1__12767_ (
);

FILL FILL_1__12347_ (
);

FILL FILL_0__9774_ (
);

FILL FILL_0__9354_ (
);

FILL FILL_3__7451_ (
);

DFFPOSX1 _11625_ (
    .D(_4777_[1]),
    .CLK(clk_bF$buf50),
    .Q(\u_fir_pe5.mul [1])
);

INVX1 _11205_ (
    .A(\X[5] [4]),
    .Y(_4402_)
);

FILL FILL_0__12701_ (
);

FILL FILL_1__7789_ (
);

FILL FILL_1__7369_ (
);

FILL FILL_3__10281_ (
);

FILL FILL_1__8730_ (
);

FILL FILL_1__8310_ (
);

FILL FILL_3__8236_ (
);

NAND3X1 _7380_ (
    .A(_892_),
    .B(_888_),
    .C(_894_),
    .Y(_901_)
);

FILL FILL_2__6653_ (
);

FILL FILL_3__11486_ (
);

FILL FILL_3__11066_ (
);

FILL FILL_2__10899_ (
);

FILL FILL_2__10479_ (
);

FILL FILL_2__10059_ (
);

FILL FILL_0__11093_ (
);

FILL FILL_1__9935_ (
);

FILL FILL_1__9515_ (
);

FILL FILL_2__11840_ (
);

FILL FILL_2__11420_ (
);

FILL FILL_0__6899_ (
);

FILL FILL_2__11000_ (
);

FILL FILL_0__6479_ (
);

AOI21X1 _8585_ (
    .A(_1937_),
    .B(_1943_),
    .C(_2018_),
    .Y(_2022_)
);

NAND3X1 _8165_ (
    .A(_2382_),
    .B(_1607_),
    .C(_1603_),
    .Y(_1608_)
);

FILL FILL_1__10833_ (
);

FILL FILL_1__10413_ (
);

FILL FILL_2__7858_ (
);

FILL FILL_0__7840_ (
);

FILL FILL_0__7420_ (
);

FILL FILL_2__7438_ (
);

FILL FILL_0__7000_ (
);

FILL FILL_2__7018_ (
);

FILL FILL_0__12298_ (
);

INVX1 _12583_ (
    .A(_5611_),
    .Y(_5625_)
);

NAND2X1 _12163_ (
    .A(_5275_),
    .B(_5243_),
    .Y(_5279_)
);

FILL FILL_2__12625_ (
);

FILL FILL_2__12205_ (
);

FILL FILL_0__8625_ (
);

FILL FILL_3__6722_ (
);

FILL FILL_0__8205_ (
);

FILL FILL_3__9194_ (
);

DFFPOSX1 _13368_ (
    .D(\Y[6] [6]),
    .CLK(clk_bF$buf48),
    .Q(\u_fir_pe7.rYin [6])
);

FILL FILL_2__7191_ (
);

FILL FILL_3__7927_ (
);

AOI21X1 _6651_ (
    .A(_247_),
    .B(_249_),
    .C(_246_),
    .Y(_250_)
);

FILL FILL_1__11791_ (
);

FILL FILL_1__11371_ (
);

FILL FILL_2__8396_ (
);

FILL FILL_0__10784_ (
);

FILL FILL_0__10364_ (
);

NOR2X1 _7856_ (
    .A(_1362_),
    .B(_1366_),
    .Y(_1370_)
);

NAND2X1 _7436_ (
    .A(_884_),
    .B(_955_),
    .Y(_956_)
);

NAND2X1 _7016_ (
    .A(_605_),
    .B(_608_),
    .Y(_609_)
);

FILL FILL_1__6393_ (
);

FILL FILL_2__13163_ (
);

FILL FILL_2__6709_ (
);

FILL FILL_1__12996_ (
);

FILL FILL_1__12576_ (
);

FILL FILL_1__12156_ (
);

FILL FILL_0__11989_ (
);

FILL FILL_0__9583_ (
);

FILL FILL_3__7680_ (
);

FILL FILL_0__9163_ (
);

NAND3X1 _11854_ (
    .A(_4918_),
    .B(_4967_),
    .C(_4968_),
    .Y(_4974_)
);

FILL FILL_0__11569_ (
);

INVX1 _11434_ (
    .A(_4622_),
    .Y(_4623_)
);

FILL FILL_0__11149_ (
);

AND2X2 _11014_ (
    .A(vdd),
    .B(\X[5] [7]),
    .Y(_4213_)
);

FILL FILL_3__12903_ (
);

FILL FILL_0__12930_ (
);

FILL FILL_1__7598_ (
);

FILL FILL_1__7178_ (
);

FILL FILL_3__8465_ (
);

NAND3X1 _12639_ (
    .A(_5675_),
    .B(_5661_),
    .C(_5679_),
    .Y(_5680_)
);

FILL FILL_3__8045_ (
);

NAND2X1 _12219_ (
    .A(_5330_),
    .B(_5333_),
    .Y(_5334_)
);

FILL FILL_2__6882_ (
);

FILL FILL_2__6462_ (
);

FILL FILL_2__10288_ (
);

FILL FILL_1__9744_ (
);

FILL FILL_1__9324_ (
);

OAI21X1 _8394_ (
    .A(_1750_),
    .B(_1754_),
    .C(_1753_),
    .Y(_1833_)
);

FILL FILL_1__10642_ (
);

FILL FILL_1__10222_ (
);

CLKBUF1 CLKBUF1_insert30 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert31 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert32 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert33 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert34 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf35)
);

FILL FILL_2__7667_ (
);

CLKBUF1 CLKBUF1_insert35 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert36 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert37 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert38 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert39 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf30)
);

NOR2X1 _12392_ (
    .A(_5495_),
    .B(_5494_),
    .Y(_5496_)
);

FILL FILL_3__13021_ (
);

INVX2 _6707_ (
    .A(gnd),
    .Y(_305_)
);

FILL FILL_2__12854_ (
);

FILL FILL_2__12434_ (
);

FILL FILL_2__12014_ (
);

OAI21X1 _9599_ (
    .A(_2921_),
    .B(_2915_),
    .C(_2925_),
    .Y(_2953_)
);

NAND3X1 _9179_ (
    .A(gnd),
    .B(\X[3] [6]),
    .C(_2536_),
    .Y(_2539_)
);

FILL FILL_1__11847_ (
);

FILL FILL_1__11427_ (
);

FILL FILL_1__11007_ (
);

FILL FILL_0__8854_ (
);

FILL FILL_0__8434_ (
);

NOR2X1 _10705_ (
    .A(_3908_),
    .B(_3972_),
    .Y(_3967_)
);

FILL FILL_0__8014_ (
);

OAI21X1 _13177_ (
    .A(_6195_),
    .B(_6194_),
    .C(_6206_),
    .Y(_6208_)
);

FILL FILL_2__9813_ (
);

FILL FILL_1__6869_ (
);

FILL FILL_1__6449_ (
);

FILL FILL_2__13219_ (
);

FILL FILL_1__7810_ (
);

FILL FILL_0__9639_ (
);

FILL FILL_0__9219_ (
);

FILL FILL_3__7316_ (
);

OAI22X1 _6880_ (
    .A(_331_),
    .B(_412_),
    .C(_474_),
    .D(_475_),
    .Y(_476_)
);

INVX1 _6460_ (
    .A(_45_),
    .Y(_62_)
);

FILL FILL_3__10986_ (
);

FILL FILL_3__10146_ (
);

FILL FILL_1__11180_ (
);

FILL FILL_0__10593_ (
);

FILL FILL_0__10173_ (
);

FILL FILL_2__10920_ (
);

FILL FILL_2__10500_ (
);

OAI21X1 _7665_ (
    .A(_1112_),
    .B(_1181_),
    .C(_1151_),
    .Y(_1182_)
);

DFFPOSX1 _7245_ (
    .D(_796_[6]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.mul [6])
);

FILL FILL_2__6938_ (
);

FILL FILL_0__6920_ (
);

FILL FILL_0__6500_ (
);

FILL FILL_2__6518_ (
);

FILL FILL_1__12385_ (
);

FILL FILL_0__9392_ (
);

FILL FILL_0__11798_ (
);

AOI22X1 _11663_ (
    .A(gnd),
    .B(\X[7] [0]),
    .C(vdd),
    .D(\X[7] [1]),
    .Y(_4786_)
);

FILL FILL_0__11378_ (
);

NOR2X1 _11243_ (
    .A(_4358_),
    .B(_4438_),
    .Y(_4439_)
);

FILL FILL_2__11705_ (
);

FILL FILL_0__7705_ (
);

NOR2X1 _9811_ (
    .A(_3154_),
    .B(_3153_),
    .Y(_3155_)
);

FILL FILL_3__8694_ (
);

AND2X2 _12868_ (
    .A(vdd),
    .B(\X[6]_5_bF$buf0 ),
    .Y(_5906_)
);

NAND2X1 _12448_ (
    .A(\u_fir_pe6.rYin [15]),
    .B(\u_fir_pe6.mul [15]),
    .Y(_5551_)
);

NAND3X1 _12028_ (
    .A(_5085_),
    .B(_5142_),
    .C(_5143_),
    .Y(_5146_)
);

FILL FILL_0__13104_ (
);

FILL FILL_2__6691_ (
);

FILL FILL_2__10097_ (
);

FILL FILL_1__9973_ (
);

FILL FILL_1__9553_ (
);

FILL FILL_1__9133_ (
);

FILL FILL_1__10871_ (
);

FILL FILL_1__10451_ (
);

FILL FILL_1__10031_ (
);

FILL FILL_2__7896_ (
);

FILL FILL_2__7476_ (
);

FILL FILL_2__7056_ (
);

FILL FILL_3__13250_ (
);

AOI21X1 _6936_ (
    .A(_482_),
    .B(_525_),
    .C(_528_),
    .Y(_531_)
);

NAND3X1 _6516_ (
    .A(_112_),
    .B(_106_),
    .C(_110_),
    .Y(_117_)
);

FILL FILL_2__12663_ (
);

FILL FILL_2__12243_ (
);

FILL FILL_1__11656_ (
);

FILL FILL_1__11236_ (
);

FILL FILL_0__8663_ (
);

FILL FILL_3__6760_ (
);

FILL FILL_0__8243_ (
);

FILL FILL_0__10649_ (
);

NAND2X1 _10934_ (
    .A(vdd),
    .B(\X[5] [6]),
    .Y(_4134_)
);

NAND2X1 _10514_ (
    .A(_3786_),
    .B(_3760_),
    .Y(_3787_)
);

FILL FILL_0__10229_ (
);

FILL FILL_2__9622_ (
);

FILL FILL_2__9202_ (
);

FILL FILL_1__6678_ (
);

FILL FILL_2__13028_ (
);

FILL FILL_0__9448_ (
);

FILL FILL_3__7545_ (
);

FILL FILL_0__9028_ (
);

OAI21X1 _11719_ (
    .A(_5563_),
    .B(_4800_),
    .C(_4803_),
    .Y(_4841_)
);

FILL FILL_3__10375_ (
);

FILL FILL_1__8824_ (
);

FILL FILL_1__8404_ (
);

OAI21X1 _7894_ (
    .A(_1388_),
    .B(_1383_),
    .C(_1406_),
    .Y(_1407_)
);

INVX1 _7474_ (
    .A(_903_),
    .Y(_994_)
);

NOR2X1 _7054_ (
    .A(\u_fir_pe0.rYin [2]),
    .B(\u_fir_pe0.mul [2]),
    .Y(_642_)
);

FILL FILL_2__6747_ (
);

FILL FILL_1__12194_ (
);

NAND2X1 _11892_ (
    .A(_5009_),
    .B(_5010_),
    .Y(_5011_)
);

AND2X2 _11472_ (
    .A(_4656_),
    .B(_4655_),
    .Y(_4775_[5])
);

FILL FILL_0__11187_ (
);

NAND3X1 _11052_ (
    .A(_4245_),
    .B(_4244_),
    .C(_4246_),
    .Y(_4251_)
);

FILL FILL_1__9609_ (
);

FILL FILL_3__12521_ (
);

FILL FILL_3__12101_ (
);

FILL FILL_2__11934_ (
);

FILL FILL_2__11514_ (
);

NOR2X1 _8679_ (
    .A(_2011_),
    .B(_2056_),
    .Y(_2114_)
);

NAND3X1 _8259_ (
    .A(_1695_),
    .B(_1699_),
    .C(_1663_),
    .Y(_1700_)
);

FILL FILL_1__10927_ (
);

FILL FILL_1__10507_ (
);

FILL FILL_0__7934_ (
);

FILL FILL_0__7514_ (
);

OR2X2 _9620_ (
    .A(_2972_),
    .B(_2970_),
    .Y(_2974_)
);

AOI21X1 _9200_ (
    .A(_2554_),
    .B(_2556_),
    .C(_2547_),
    .Y(_2560_)
);

FILL FILL_1__13399_ (
);

OAI21X1 _12677_ (
    .A(_5681_),
    .B(_5716_),
    .C(_5675_),
    .Y(_5717_)
);

INVX1 _12257_ (
    .A(_5367_),
    .Y(_5371_)
);

FILL FILL_2__12719_ (
);

FILL FILL_0__13333_ (
);

FILL FILL_0__8719_ (
);

FILL FILL_3__6816_ (
);

FILL FILL_1__9782_ (
);

FILL FILL_1__9362_ (
);

FILL FILL_3__9288_ (
);

FILL FILL_1__10680_ (
);

FILL FILL_1__10260_ (
);

FILL FILL_2__7285_ (
);

NAND3X1 _6745_ (
    .A(_323_),
    .B(_338_),
    .C(_339_),
    .Y(_343_)
);

FILL FILL_2__12892_ (
);

FILL FILL_2__12052_ (
);

FILL FILL_1__11885_ (
);

FILL FILL_1__11465_ (
);

FILL FILL_1__11045_ (
);

FILL FILL_0__8892_ (
);

FILL FILL_0__8472_ (
);

FILL FILL_0__10878_ (
);

FILL FILL_0__10458_ (
);

DFFPOSX1 _10743_ (
    .D(\Y[4] [12]),
    .CLK(clk_bF$buf43),
    .Q(\u_fir_pe4.rYin [12])
);

FILL FILL_0__8052_ (
);

NAND2X1 _10323_ (
    .A(gnd),
    .B(\X[4] [7]),
    .Y(_3600_)
);

FILL FILL_0__10038_ (
);

FILL FILL253950x10950 (
);

FILL FILL_2__9431_ (
);

FILL FILL_2__9011_ (
);

FILL FILL_1__6487_ (
);

FILL FILL_2__13257_ (
);

FILL FILL_0__9677_ (
);

FILL FILL_3__7774_ (
);

FILL FILL_0__9257_ (
);

OAI21X1 _11948_ (
    .A(_5066_),
    .B(_5062_),
    .C(_4978_),
    .Y(_5067_)
);

NOR2X1 _11528_ (
    .A(\u_fir_pe5.rYin [10]),
    .B(\u_fir_pe5.mul [10]),
    .Y(_4712_)
);

NAND2X1 _11108_ (
    .A(\X[5] [4]),
    .B(gnd),
    .Y(_4306_)
);

FILL FILL_0__12604_ (
);

FILL FILL_1__8633_ (
);

FILL FILL_1__8213_ (
);

FILL FILL_3__8559_ (
);

NAND3X1 _7283_ (
    .A(_1537_),
    .B(_805_),
    .C(_803_),
    .Y(_806_)
);

FILL FILL_3__9920_ (
);

FILL FILL_2__6976_ (
);

FILL FILL_2__6556_ (
);

FILL FILL_3__11389_ (
);

NAND3X1 _11281_ (
    .A(_4472_),
    .B(_4476_),
    .C(_4446_),
    .Y(_4477_)
);

FILL FILL_1__9418_ (
);

FILL FILL_3__12750_ (
);

FILL FILL_3__12330_ (
);

FILL FILL_2__11743_ (
);

FILL FILL_2__11323_ (
);

NAND2X1 _8488_ (
    .A(_1921_),
    .B(_1925_),
    .Y(_1926_)
);

OAI21X1 _8068_ (
    .A(_1559_),
    .B(_1562_),
    .C(_1569_),
    .Y(_1572_)
);

FILL FILL_1__10316_ (
);

FILL FILL_0__7743_ (
);

FILL FILL_0__7323_ (
);

DFFPOSX1 _12486_ (
    .D(\Y[7] [1]),
    .CLK(clk_bF$buf27),
    .Q(\u_fir_pe6.rYin [1])
);

NAND2X1 _12066_ (
    .A(gnd),
    .B(\X[7] [6]),
    .Y(_5183_)
);

FILL FILL_2__8702_ (
);

FILL FILL_3__13115_ (
);

FILL FILL_2__12948_ (
);

FILL FILL_2__12528_ (
);

FILL FILL_2__12108_ (
);

FILL FILL_0__13142_ (
);

FILL FILL_0__8948_ (
);

FILL FILL_0__8528_ (
);

FILL FILL_1__9591_ (
);

FILL FILL_1__9171_ (
);

FILL FILL_3__9097_ (
);

FILL FILL_2__9907_ (
);

FILL FILL_2__7094_ (
);

FILL FILL_1__7904_ (
);

NOR2X1 _6974_ (
    .A(_567_),
    .B(_566_),
    .Y(_568_)
);

AOI22X1 _6554_ (
    .A(gnd),
    .B(Xin[2]),
    .C(vdd),
    .D(Xin[3]),
    .Y(_154_)
);

FILL FILL_2__12281_ (
);

FILL FILL_1__11694_ (
);

FILL FILL_1__11274_ (
);

FILL FILL253650x237750 (
);

FILL FILL_2__8299_ (
);

FILL FILL_0__8281_ (
);

FILL FILL_0__10687_ (
);

NAND3X1 _10972_ (
    .A(_4169_),
    .B(_4170_),
    .C(_4171_),
    .Y(_4172_)
);

INVX1 _10552_ (
    .A(\u_fir_pe4.mul [1]),
    .Y(_3821_)
);

FILL FILL_0__10267_ (
);

AOI21X1 _10132_ (
    .A(_3350_),
    .B(_3354_),
    .C(_3343_),
    .Y(_3411_)
);

FILL FILL_2__9660_ (
);

FILL FILL_2__9240_ (
);

AND2X2 _7759_ (
    .A(\X[1]_5_bF$buf1 ),
    .B(gnd),
    .Y(_1275_)
);

OAI21X1 _7339_ (
    .A(_860_),
    .B(_859_),
    .C(_826_),
    .Y(_861_)
);

FILL FILL_2__13066_ (
);

FILL FILL_1__12899_ (
);

NAND2X1 _8700_ (
    .A(_2134_),
    .B(_2133_),
    .Y(_2135_)
);

FILL FILL_1__12059_ (
);

FILL FILL_0__9486_ (
);

FILL FILL_0__9066_ (
);

NAND3X1 _11757_ (
    .A(_4866_),
    .B(_4877_),
    .C(_4873_),
    .Y(_4878_)
);

FILL FILL_3__7163_ (
);

NAND2X1 _11337_ (
    .A(_4527_),
    .B(_4531_),
    .Y(_4532_)
);

FILL FILL_1__13000_ (
);

FILL FILL_0__12833_ (
);

FILL FILL_0__12413_ (
);

NAND2X1 _9905_ (
    .A(vdd),
    .B(\X[4] [2]),
    .Y(_3188_)
);

FILL FILL_1__8862_ (
);

FILL FILL_1__8442_ (
);

FILL FILL_1__8022_ (
);

FILL FILL_3__8788_ (
);

NOR2X1 _7092_ (
    .A(\u_fir_pe0.rYin [6]),
    .B(\u_fir_pe0.mul [6]),
    .Y(_676_)
);

FILL FILL_2__6785_ (
);

OAI21X1 _11090_ (
    .A(_4207_),
    .B(_4287_),
    .C(_4256_),
    .Y(_4288_)
);

FILL FILL_1__9647_ (
);

FILL FILL_1__9227_ (
);

FILL FILL_2__11972_ (
);

FILL FILL_2__11552_ (
);

FILL FILL_2__11132_ (
);

NAND2X1 _8297_ (
    .A(_1735_),
    .B(_1736_),
    .Y(_1737_)
);

FILL FILL_1__10965_ (
);

FILL FILL_1__10545_ (
);

FILL FILL_1__10125_ (
);

FILL FILL_0__7972_ (
);

FILL FILL_0__7552_ (
);

FILL FILL_0__7132_ (
);

NAND2X1 _12295_ (
    .A(_5406_),
    .B(_5370_),
    .Y(_5407_)
);

FILL FILL_2__8931_ (
);

FILL FILL_2__8511_ (
);

FILL FILL_2__12757_ (
);

FILL FILL_2__12337_ (
);

FILL FILL_0__8757_ (
);

FILL FILL_3__6854_ (
);

FILL FILL_0__8337_ (
);

FILL FILL_3__6434_ (
);

NOR2X1 _10608_ (
    .A(_3869_),
    .B(_3870_),
    .Y(_3871_)
);

FILL FILL_2__9716_ (
);

FILL FILL_1__7713_ (
);

FILL FILL_3__7639_ (
);

AOI21X1 _6783_ (
    .A(_297_),
    .B(_367_),
    .C(_379_),
    .Y(_380_)
);

FILL FILL_2__12090_ (
);

FILL FILL_3__10889_ (
);

FILL FILL_3__10469_ (
);

FILL FILL_1__11083_ (
);

FILL FILL_0__10496_ (
);

INVX1 _10781_ (
    .A(_4772_),
    .Y(_4773_)
);

AND2X2 _10361_ (
    .A(_3637_),
    .B(_3630_),
    .Y(_3638_)
);

FILL FILL_0__10076_ (
);

FILL FILL_1__8918_ (
);

FILL FILL_3__11830_ (
);

FILL FILL_2__10823_ (
);

FILL FILL_2__10403_ (
);

NAND2X1 _7988_ (
    .A(_1454_),
    .B(_1466_),
    .Y(_1491_)
);

OAI21X1 _7568_ (
    .A(_1004_),
    .B(_1001_),
    .C(_1086_),
    .Y(_1087_)
);

OAI21X1 _7148_ (
    .A(_724_),
    .B(_725_),
    .C(_729_),
    .Y(_732_)
);

FILL FILL_2__13295_ (
);

FILL FILL_0__6823_ (
);

FILL FILL_0__6403_ (
);

FILL FILL_1__12288_ (
);

FILL FILL_0__9295_ (
);

OAI21X1 _11986_ (
    .A(_5100_),
    .B(_5103_),
    .C(_5102_),
    .Y(_5104_)
);

FILL FILL_3__7392_ (
);

AND2X2 _11566_ (
    .A(_4743_),
    .B(_4749_),
    .Y(_4750_)
);

AOI21X1 _11146_ (
    .A(_4255_),
    .B(_4257_),
    .C(_4343_),
    .Y(_4344_)
);

FILL FILL_3__12615_ (
);

FILL FILL_3_BUFX2_insert10 (
);

FILL FILL_0__12642_ (
);

FILL FILL_0__12222_ (
);

FILL FILL_0__7608_ (
);

NOR2X1 _9714_ (
    .A(\u_fir_pe3.rYin [5]),
    .B(\u_fir_pe3.mul [5]),
    .Y(_3059_)
);

FILL FILL_1__8671_ (
);

FILL FILL_1__8251_ (
);

FILL FILL_3__8177_ (
);

FILL FILL_0__13007_ (
);

FILL FILL_2__6594_ (
);

FILL FILL_1__9456_ (
);

FILL FILL_1__9036_ (
);

FILL FILL_2__11781_ (
);

FILL FILL_2__11361_ (
);

FILL FILL_1__10774_ (
);

FILL FILL_1__10354_ (
);

FILL FILL_2__7799_ (
);

FILL FILL_0__7781_ (
);

FILL FILL_2__7379_ (
);

FILL FILL_0__7361_ (
);

FILL FILL_2__8740_ (
);

FILL FILL_2__8320_ (
);

OAI21X1 _6839_ (
    .A(_435_),
    .B(_434_),
    .C(_433_),
    .Y(_436_)
);

INVX1 _6419_ (
    .A(_21_),
    .Y(_22_)
);

FILL FILL_2__12986_ (
);

FILL FILL_2__12566_ (
);

FILL FILL_2__12146_ (
);

FILL FILL_0__13180_ (
);

FILL FILL_1__11979_ (
);

FILL FILL_1__11559_ (
);

FILL FILL_1__11139_ (
);

FILL FILL_0__8566_ (
);

FILL FILL_3__6663_ (
);

FILL FILL_0__8146_ (
);

INVX1 _10837_ (
    .A(_4038_),
    .Y(_4039_)
);

NOR2X1 _10417_ (
    .A(_3690_),
    .B(_3692_),
    .Y(_3693_)
);

FILL FILL_1__12920_ (
);

FILL FILL_2__9945_ (
);

FILL FILL_0__11913_ (
);

FILL FILL_2__9525_ (
);

FILL FILL_2__9105_ (
);

FILL FILL_1__7942_ (
);

FILL FILL_1__7522_ (
);

FILL FILL_1__7102_ (
);

FILL FILL_3__7868_ (
);

FILL FILL_3__7028_ (
);

NAND3X1 _6592_ (
    .A(_136_),
    .B(_185_),
    .C(_186_),
    .Y(_192_)
);

FILL FILL_3__10698_ (
);

NOR2X1 _10590_ (
    .A(_3853_),
    .B(_3854_),
    .Y(_3855_)
);

OAI21X1 _10170_ (
    .A(_3438_),
    .B(_3433_),
    .C(_3440_),
    .Y(_3449_)
);

FILL FILL_1__8727_ (
);

FILL FILL_1__8307_ (
);

FILL FILL_2__10632_ (
);

FILL FILL_2__10212_ (
);

NAND2X1 _7797_ (
    .A(_1265_),
    .B(_1266_),
    .Y(_1312_)
);

NAND3X1 _7377_ (
    .A(_893_),
    .B(_879_),
    .C(_897_),
    .Y(_898_)
);

FILL FILL_0__6632_ (
);

FILL FILL_1__12097_ (
);

OAI21X1 _11795_ (
    .A(_5492_),
    .B(_4914_),
    .C(_4859_),
    .Y(_4915_)
);

OR2X2 _11375_ (
    .A(_4568_),
    .B(_4545_),
    .Y(_4569_)
);

FILL FILL_3__12844_ (
);

FILL FILL_3__12424_ (
);

FILL FILL_3__12004_ (
);

FILL FILL_2__11837_ (
);

FILL FILL_0__12871_ (
);

FILL FILL_2__11417_ (
);

FILL FILL_0__12451_ (
);

FILL FILL_0__12031_ (
);

FILL FILL_0__7837_ (
);

NAND2X1 _9943_ (
    .A(_3223_),
    .B(_3224_),
    .Y(_3225_)
);

FILL FILL_0__7417_ (
);

NAND2X1 _9523_ (
    .A(_2860_),
    .B(_2857_),
    .Y(_2879_)
);

NAND2X1 _9103_ (
    .A(_3091_),
    .B(_2463_),
    .Y(_2464_)
);

FILL FILL_1__8480_ (
);

FILL FILL_1__8060_ (
);

FILL FILL_3__13209_ (
);

FILL FILL_0__13236_ (
);

NOR3X1 _13101_ (
    .A(_6081_),
    .B(_6083_),
    .C(_6131_),
    .Y(_6135_)
);

FILL FILL_1__9685_ (
);

FILL FILL_1__9265_ (
);

FILL FILL253950x216150 (
);

FILL FILL_2__11170_ (
);

FILL FILL_1__10583_ (
);

FILL FILL_1__10163_ (
);

FILL FILL_0__7590_ (
);

FILL FILL_2__7188_ (
);

FILL FILL_0__7170_ (
);

NAND2X1 _6648_ (
    .A(_158_),
    .B(_242_),
    .Y(_247_)
);

FILL FILL_2__12795_ (
);

FILL FILL_2__12375_ (
);

FILL FILL_1__11788_ (
);

FILL FILL_1__11368_ (
);

FILL FILL_0__8795_ (
);

FILL FILL_0__8375_ (
);

AOI21X1 _10646_ (
    .A(_3891_),
    .B(_3906_),
    .C(_3909_),
    .Y(_3910_)
);

AOI21X1 _10226_ (
    .A(_3444_),
    .B(_3441_),
    .C(_3427_),
    .Y(_3504_)
);

FILL FILL_2__9754_ (
);

FILL FILL_2__9334_ (
);

FILL FILL_0__11722_ (
);

FILL FILL_0__11302_ (
);

FILL FILL_1__7751_ (
);

FILL FILL_1__7331_ (
);

FILL FILL_3__7257_ (
);

FILL FILL_0__12927_ (
);

FILL FILL_3__10087_ (
);

FILL FILL_1__8536_ (
);

FILL FILL_2__10861_ (
);

FILL FILL_2__10441_ (
);

FILL FILL_2__10021_ (
);

NAND2X1 _7186_ (
    .A(\u_fir_pe0.rYin [15]),
    .B(\u_fir_pe0.mul [15]),
    .Y(_769_)
);

FILL FILL_3__9403_ (
);

FILL FILL_2__6879_ (
);

FILL FILL_0__6861_ (
);

FILL FILL_0__6441_ (
);

FILL FILL_2__6459_ (
);

AOI21X1 _11184_ (
    .A(_4324_),
    .B(_4323_),
    .C(_4308_),
    .Y(_4381_)
);

FILL FILL_2__7820_ (
);

FILL FILL_2__7400_ (
);

FILL FILL254250x126150 (
);

FILL FILL_2__11646_ (
);

FILL FILL_0__12680_ (
);

FILL FILL_2__11226_ (
);

FILL FILL_0__12260_ (
);

FILL FILL_1__10639_ (
);

FILL FILL_1__10219_ (
);

FILL FILL_0__7646_ (
);

NOR2X1 _9752_ (
    .A(_3084_),
    .B(_3083_),
    .Y(_3096_)
);

AOI21X1 _9332_ (
    .A(_2672_),
    .B(_2674_),
    .C(_2689_),
    .Y(_2690_)
);

OAI21X1 _12389_ (
    .A(_5491_),
    .B(_5488_),
    .C(_5490_),
    .Y(_5493_)
);

FILL FILL_2__8605_ (
);

FILL FILL_0__13045_ (
);

OAI21X1 _13330_ (
    .A(_6341_),
    .B(_6344_),
    .C(_6351_),
    .Y(_6354_)
);

FILL FILL_1__6602_ (
);

FILL FILL_3__6528_ (
);

FILL FILL_1__9494_ (
);

FILL FILL_1__9074_ (
);

FILL FILL_1__10392_ (
);

FILL FILL_1__7807_ (
);

FILL FILL_3__13191_ (
);

NAND2X1 _6877_ (
    .A(gnd),
    .B(Xin[6]),
    .Y(_473_)
);

OAI21X1 _6457_ (
    .A(_781_),
    .B(_18_),
    .C(_21_),
    .Y(_59_)
);

FILL FILL_2__12184_ (
);

FILL FILL_1__11177_ (
);

FILL FILL_0__8184_ (
);

NAND3X1 _10875_ (
    .A(_4071_),
    .B(_4075_),
    .C(_4073_),
    .Y(_4076_)
);

NAND3X1 _10455_ (
    .A(_3703_),
    .B(_3729_),
    .C(_3725_),
    .Y(_3730_)
);

INVX1 _10035_ (
    .A(_3308_),
    .Y(_3316_)
);

FILL FILL_3__11924_ (
);

FILL FILL_2__9983_ (
);

FILL FILL_2__10917_ (
);

FILL FILL_2__9563_ (
);

FILL FILL_0__11951_ (
);

FILL FILL_2__9143_ (
);

FILL FILL_0__11531_ (
);

FILL FILL_0__11111_ (
);

FILL FILL_0__6917_ (
);

NAND3X1 _8603_ (
    .A(_2020_),
    .B(_2024_),
    .C(_2027_),
    .Y(_2040_)
);

FILL FILL_1__7980_ (
);

FILL FILL_1__7560_ (
);

FILL FILL_1__7140_ (
);

FILL FILL_0__9389_ (
);

FILL FILL_3__7486_ (
);

FILL FILL_3__12709_ (
);

FILL FILL_1__13323_ (
);

FILL FILL_0__12736_ (
);

OAI21X1 _12601_ (
    .A(_5642_),
    .B(_5641_),
    .C(_5608_),
    .Y(_5643_)
);

FILL FILL_0__12316_ (
);

INVX1 _9808_ (
    .A(\u_fir_pe3.mul [14]),
    .Y(_3152_)
);

FILL FILL_1__8765_ (
);

FILL FILL_1__8345_ (
);

FILL FILL_2__10670_ (
);

FILL FILL_2__10250_ (
);

FILL FILL_3__9632_ (
);

FILL FILL_2__6688_ (
);

FILL FILL_0__6670_ (
);

FILL FILL_3__12042_ (
);

FILL FILL_2__11875_ (
);

FILL FILL_2__11455_ (
);

FILL FILL_2__11035_ (
);

FILL FILL_1__10868_ (
);

FILL FILL_1__10448_ (
);

FILL FILL_1__10028_ (
);

FILL FILL_0__7875_ (
);

INVX2 _9981_ (
    .A(\X[4]_5_bF$buf2 ),
    .Y(_3262_)
);

FILL FILL_0__7455_ (
);

NAND2X1 _9561_ (
    .A(_2722_),
    .B(_2796_),
    .Y(_2916_)
);

FILL FILL_0__7035_ (
);

NAND3X1 _9141_ (
    .A(_2417_),
    .B(_2497_),
    .C(_2501_),
    .Y(_2502_)
);

AOI21X1 _12198_ (
    .A(_5264_),
    .B(_5307_),
    .C(_5310_),
    .Y(_5313_)
);

FILL FILL_2__8834_ (
);

FILL FILL_2__8414_ (
);

FILL FILL_0__10802_ (
);

FILL FILL_0__13274_ (
);

FILL FILL_1__6831_ (
);

FILL FILL_1__6411_ (
);

FILL FILL_3__6757_ (
);

FILL FILL_2__9619_ (
);

FILL FILL_0__9601_ (
);

FILL FILL_1__7616_ (
);

OAI21X1 _6686_ (
    .A(_284_),
    .B(_280_),
    .C(_196_),
    .Y(_285_)
);

INVX1 _10684_ (
    .A(\u_fir_pe4.rYin [14]),
    .Y(_3947_)
);

FILL FILL_0__10399_ (
);

NAND3X1 _10264_ (
    .A(_3537_),
    .B(_3538_),
    .C(_3505_),
    .Y(_3542_)
);

FILL FILL_2__6900_ (
);

FILL FILL_3__11313_ (
);

FILL FILL_2__9792_ (
);

FILL FILL_2__9372_ (
);

FILL FILL_0__11760_ (
);

FILL FILL_2__10306_ (
);

FILL FILL_0__11340_ (
);

FILL FILL_2__13198_ (
);

FILL FILL_0__6726_ (
);

AND2X2 _8832_ (
    .A(_2257_),
    .B(_2256_),
    .Y(_2384_[4])
);

NAND3X1 _8412_ (
    .A(_1847_),
    .B(_1846_),
    .C(_1850_),
    .Y(_1851_)
);

FILL FILL_0__9198_ (
);

INVX1 _11889_ (
    .A(_5007_),
    .Y(_5008_)
);

NOR2X1 _11469_ (
    .A(_4653_),
    .B(_4652_),
    .Y(_4654_)
);

OAI21X1 _11049_ (
    .A(_4243_),
    .B(_4247_),
    .C(_4209_),
    .Y(_4248_)
);

FILL FILL_3__12938_ (
);

FILL FILL_1__13132_ (
);

FILL FILL_0__12965_ (
);

OAI21X1 _12830_ (
    .A(_5786_),
    .B(_5783_),
    .C(_5868_),
    .Y(_5869_)
);

FILL FILL_0__12545_ (
);

FILL FILL_0__12125_ (
);

OAI21X1 _12410_ (
    .A(_5506_),
    .B(_5507_),
    .C(_5511_),
    .Y(_5514_)
);

NAND3X1 _9617_ (
    .A(_2952_),
    .B(_2969_),
    .C(_2968_),
    .Y(_2971_)
);

FILL FILL_1__8574_ (
);

FILL FILL_1__8154_ (
);

FILL FILL_3__9021_ (
);

FILL FILL_2__6497_ (
);

FILL FILL_1__9779_ (
);

FILL FILL_1__9359_ (
);

FILL FILL_3__12691_ (
);

FILL FILL_3__12271_ (
);

FILL FILL_2__11684_ (
);

FILL FILL_2__11264_ (
);

FILL FILL_1__10677_ (
);

FILL FILL_1__10257_ (
);

FILL FILL_0__7684_ (
);

INVX1 _9790_ (
    .A(\u_fir_pe3.mul [12]),
    .Y(_3134_)
);

FILL FILL_0__7264_ (
);

AOI21X1 _9370_ (
    .A(_2637_),
    .B(_2640_),
    .C(_2646_),
    .Y(_2728_)
);

FILL FILL_2__8643_ (
);

FILL FILL_2__8223_ (
);

FILL FILL_0__10611_ (
);

FILL FILL_3__13056_ (
);

FILL FILL_2__12889_ (
);

FILL FILL_2__12049_ (
);

FILL FILL_0__13083_ (
);

FILL FILL_1__6640_ (
);

FILL FILL_2__13410_ (
);

FILL FILL_0__8889_ (
);

FILL FILL_0__8469_ (
);

FILL FILL_0__8049_ (
);

FILL FILL_1__12823_ (
);

FILL FILL_1__12403_ (
);

FILL FILL_2__9428_ (
);

FILL FILL_0__9410_ (
);

FILL FILL_0__11816_ (
);

FILL FILL253350x158550 (
);

FILL FILL_1__7845_ (
);

FILL FILL_1__7425_ (
);

FILL FILL_1__7005_ (
);

NAND3X1 _6495_ (
    .A(_84_),
    .B(_95_),
    .C(_91_),
    .Y(_96_)
);

FILL FILL_3__8712_ (
);

AOI21X1 _10493_ (
    .A(_3765_),
    .B(_3766_),
    .C(_3749_),
    .Y(_3767_)
);

NAND3X1 _10073_ (
    .A(gnd),
    .B(\X[4] [3]),
    .C(_3352_),
    .Y(_3353_)
);

FILL FILL_3__11542_ (
);

FILL FILL_2__10955_ (
);

FILL FILL_2__10535_ (
);

FILL FILL_2__9181_ (
);

FILL FILL_2__10115_ (
);

FILL FILL_0__6955_ (
);

FILL FILL_0__6535_ (
);

AND2X2 _8641_ (
    .A(_2070_),
    .B(_2076_),
    .Y(_2077_)
);

NOR3X1 _8221_ (
    .A(_1647_),
    .B(_1614_),
    .C(_1659_),
    .Y(_1662_)
);

AOI22X1 _11698_ (
    .A(gnd),
    .B(\X[7] [1]),
    .C(vdd),
    .D(\X[7] [2]),
    .Y(_4820_)
);

NAND2X1 _11278_ (
    .A(_4470_),
    .B(_4457_),
    .Y(_4474_)
);

FILL FILL_2__7914_ (
);

FILL FILL_3__12327_ (
);

FILL FILL_0__12774_ (
);

FILL FILL_0__12354_ (
);

DFFPOSX1 _9846_ (
    .D(\X[3] [0]),
    .CLK(clk_bF$buf15),
    .Q(\X[4] [0])
);

INVX1 _9426_ (
    .A(_2777_),
    .Y(_2783_)
);

DFFPOSX1 _9006_ (
    .D(_2390_[13]),
    .CLK(clk_bF$buf28),
    .Q(\u_fir_pe2.mul [13])
);

FILL FILL_1__8383_ (
);

FILL FILL254250x10950 (
);

FILL FILL_3__9670_ (
);

FILL FILL_3__9250_ (
);

FILL FILL_0__13139_ (
);

OAI21X1 _13004_ (
    .A(_6006_),
    .B(_6008_),
    .C(_6002_),
    .Y(_6040_)
);

FILL FILL254550x244950 (
);

FILL FILL_1__9588_ (
);

FILL FILL_1__9168_ (
);

FILL FILL_2__11493_ (
);

FILL FILL_2__11073_ (
);

FILL FILL_1__10486_ (
);

FILL FILL_1__10066_ (
);

FILL FILL_0__7493_ (
);

FILL FILL_0__7073_ (
);

FILL FILL_3__10813_ (
);

FILL FILL_2__8872_ (
);

FILL FILL_2__8452_ (
);

FILL FILL_0__10840_ (
);

FILL FILL_3__13285_ (
);

FILL FILL_0__10420_ (
);

FILL FILL_2__8032_ (
);

FILL FILL_0__10000_ (
);

FILL FILL_2__12698_ (
);

FILL FILL_2__12278_ (
);

INVX1 _7912_ (
    .A(_1418_),
    .Y(_1424_)
);

FILL FILL_0__8698_ (
);

FILL FILL_3__6795_ (
);

FILL FILL_0__8278_ (
);

AND2X2 _10969_ (
    .A(_4119_),
    .B(_4120_),
    .Y(_4169_)
);

INVX1 _10549_ (
    .A(_3212_),
    .Y(_3979_[0])
);

NOR2X1 _10129_ (
    .A(_3401_),
    .B(_3403_),
    .Y(_3408_)
);

FILL FILL_1__12632_ (
);

FILL FILL_1__12212_ (
);

FILL FILL_2__9657_ (
);

NAND2X1 _11910_ (
    .A(_4940_),
    .B(_5024_),
    .Y(_5029_)
);

FILL FILL_2__9237_ (
);

FILL FILL_0__11205_ (
);

FILL FILL_1__7654_ (
);

FILL FILL_1__13417_ (
);

FILL FILL_3__8941_ (
);

FILL FILL_1__8859_ (
);

FILL FILL_3__11771_ (
);

FILL FILL_1__8439_ (
);

FILL FILL_1__8019_ (
);

FILL FILL_2__10764_ (
);

FILL FILL_2__10344_ (
);

FILL FILL_1__9800_ (
);

INVX1 _7089_ (
    .A(\u_fir_pe0.rYin [6]),
    .Y(_673_)
);

FILL FILL_3__9726_ (
);

FILL FILL_0__6764_ (
);

AOI21X1 _8870_ (
    .A(_2289_),
    .B(_2292_),
    .C(_2291_),
    .Y(_2293_)
);

AND2X2 _8450_ (
    .A(_1888_),
    .B(_1884_),
    .Y(_2390_[7])
);

AND2X2 _8030_ (
    .A(_1529_),
    .B(_1532_),
    .Y(_1534_)
);

OAI21X1 _11087_ (
    .A(_4195_),
    .B(_4205_),
    .C(_4201_),
    .Y(_4285_)
);

FILL FILL_2__7723_ (
);

FILL FILL_3__12556_ (
);

FILL FILL_2__7303_ (
);

FILL FILL_1__13170_ (
);

FILL FILL_2__11969_ (
);

FILL FILL_2__11549_ (
);

FILL FILL_0__12583_ (
);

FILL FILL_2__11129_ (
);

FILL FILL_0__12163_ (
);

FILL FILL_2__12910_ (
);

FILL FILL_0__7969_ (
);

FILL FILL_0__7549_ (
);

OAI21X1 _9655_ (
    .A(_2975_),
    .B(_3000_),
    .C(_2999_),
    .Y(_3007_)
);

FILL FILL_0__7129_ (
);

AOI21X1 _9235_ (
    .A(_2511_),
    .B(_2517_),
    .C(_2594_),
    .Y(_2595_)
);

FILL FILL_1__8192_ (
);

FILL FILL_1__11903_ (
);

FILL FILL_0__8910_ (
);

FILL FILL_2__8928_ (
);

FILL FILL_2__8508_ (
);

NAND2X1 _13233_ (
    .A(_6256_),
    .B(_6251_),
    .Y(_6257_)
);

FILL FILL_1__6925_ (
);

FILL FILL_1__6505_ (
);

FILL FILL_1__9397_ (
);

FILL FILL_1__10295_ (
);

FILL FILL_3__10622_ (
);

FILL FILL_2__8681_ (
);

FILL FILL_2__8261_ (
);

FILL FILL_2__12087_ (
);

OAI21X1 _7721_ (
    .A(_1237_),
    .B(_1236_),
    .C(_1235_),
    .Y(_1238_)
);

NOR2X1 _7301_ (
    .A(_821_),
    .B(_822_),
    .Y(_823_)
);

NAND2X1 _10778_ (
    .A(_4705_),
    .B(_4769_),
    .Y(_4770_)
);

AOI21X1 _10358_ (
    .A(_3634_),
    .B(_3633_),
    .C(_3626_),
    .Y(_3635_)
);

FILL FILL_3__11827_ (
);

FILL FILL_1__12861_ (
);

FILL FILL_3__11407_ (
);

FILL FILL_1__12441_ (
);

FILL FILL_1__12021_ (
);

FILL FILL_2__9886_ (
);

FILL FILL_2__9466_ (
);

FILL FILL_0__11854_ (
);

FILL FILL_2__9046_ (
);

FILL FILL_0__11434_ (
);

FILL FILL_0__11014_ (
);

NAND2X1 _8926_ (
    .A(_2349_),
    .B(_2343_),
    .Y(_2350_)
);

NAND3X1 _8506_ (
    .A(_1916_),
    .B(_1934_),
    .C(_1930_),
    .Y(_1944_)
);

FILL FILL_1__7883_ (
);

FILL FILL_1__7463_ (
);

FILL FILL_1__7043_ (
);

FILL FILL_1__13226_ (
);

OAI21X1 _12924_ (
    .A(_5880_),
    .B(_5960_),
    .C(_5943_),
    .Y(_5961_)
);

FILL FILL_0__12639_ (
);

FILL FILL_3__8330_ (
);

FILL FILL_0__12219_ (
);

DFFPOSX1 _12504_ (
    .D(_5576_[3]),
    .CLK(clk_bF$buf8),
    .Q(\u_fir_pe6.mul [3])
);

FILL FILL_1__8668_ (
);

FILL FILL_1__8248_ (
);

FILL FILL_3__11580_ (
);

FILL FILL_3__11160_ (
);

FILL FILL_2__10993_ (
);

FILL FILL_2__10573_ (
);

FILL FILL_2__10153_ (
);

FILL FILL_3__9955_ (
);

FILL FILL_3__9115_ (
);

FILL FILL_0__6993_ (
);

FILL FILL_0__6573_ (
);

FILL FILL_2__7952_ (
);

FILL FILL_3__12785_ (
);

FILL FILL_2__7532_ (
);

FILL FILL_3__12365_ (
);

FILL FILL_2__7112_ (
);

FILL FILL_2__11778_ (
);

FILL FILL_2__11358_ (
);

FILL FILL_0__12392_ (
);

FILL FILL_0__7778_ (
);

DFFPOSX1 _9884_ (
    .D(_3187_[14]),
    .CLK(clk_bF$buf56),
    .Q(\u_fir_pe3.mul [14])
);

FILL FILL_0__7358_ (
);

OAI21X1 _9464_ (
    .A(_2820_),
    .B(_2819_),
    .C(_2818_),
    .Y(_2821_)
);

NAND2X1 _9044_ (
    .A(_2404_),
    .B(_2400_),
    .Y(_2407_)
);

FILL FILL_1__11712_ (
);

FILL FILL_2__8737_ (
);

FILL FILL_2__8317_ (
);

FILL FILL_0__10705_ (
);

FILL FILL_0__13177_ (
);

AND2X2 _13042_ (
    .A(_6066_),
    .B(_6070_),
    .Y(_6078_)
);

FILL FILL_1__6734_ (
);

FILL FILL_1__12917_ (
);

FILL FILL_0__9924_ (
);

FILL FILL_0__9504_ (
);

FILL FILL_3__7601_ (
);

FILL FILL_1__7939_ (
);

FILL FILL_1__7519_ (
);

FILL FILL_3__10011_ (
);

FILL FILL254250x230550 (
);

FILL FILL_2__8490_ (
);

FILL FILL_2__8070_ (
);

AOI21X1 _6589_ (
    .A(_101_),
    .B(_105_),
    .C(_69_),
    .Y(_189_)
);

FILL FILL_3__8806_ (
);

NOR2X1 _7950_ (
    .A(_1455_),
    .B(_1454_),
    .Y(_1456_)
);

AOI22X1 _7530_ (
    .A(_884_),
    .B(_955_),
    .C(_958_),
    .D(_954_),
    .Y(_1049_)
);

NOR2X1 _7110_ (
    .A(\u_fir_pe0.rYin [8]),
    .B(\u_fir_pe0.mul [8]),
    .Y(_693_)
);

OAI21X1 _10587_ (
    .A(_3843_),
    .B(_3844_),
    .C(_3850_),
    .Y(_3852_)
);

AOI21X1 _10167_ (
    .A(_3439_),
    .B(_3445_),
    .C(_3426_),
    .Y(_3446_)
);

FILL FILL_2__6803_ (
);

FILL FILL_1__12670_ (
);

FILL FILL_1__12250_ (
);

FILL FILL_2__9695_ (
);

FILL FILL_2__10629_ (
);

FILL FILL_2__9275_ (
);

FILL FILL_0__11663_ (
);

FILL FILL_2__10209_ (
);

FILL FILL_0__11243_ (
);

FILL FILL_0__6629_ (
);

OAI21X1 _8735_ (
    .A(_2167_),
    .B(_2168_),
    .C(_2120_),
    .Y(_2169_)
);

INVX1 _8315_ (
    .A(_1754_),
    .Y(_1755_)
);

FILL FILL_1__7692_ (
);

FILL FILL_1__7272_ (
);

FILL FILL_3__7198_ (
);

FILL FILL_1__13035_ (
);

FILL FILL_0__12868_ (
);

OAI21X1 _12733_ (
    .A(_5772_),
    .B(_5767_),
    .C(_5695_),
    .Y(_5773_)
);

FILL FILL_0__12448_ (
);

FILL FILL_0__12028_ (
);

NOR2X1 _12313_ (
    .A(_5421_),
    .B(_5420_),
    .Y(_5572_[1])
);

FILL FILL_1__8897_ (
);

FILL FILL_1__8477_ (
);

FILL FILL_1__8057_ (
);

FILL FILL_2__10382_ (
);

FILL FILL_3__9344_ (
);

FILL FILL_0__6382_ (
);

FILL FILL_2__7761_ (
);

FILL FILL_2__7341_ (
);

FILL FILL_2__11167_ (
);

NOR2X1 _6801_ (
    .A(_132_),
    .B(_321_),
    .Y(_398_)
);

FILL FILL_0__7587_ (
);

INVX1 _9693_ (
    .A(\u_fir_pe3.mul [3]),
    .Y(_3040_)
);

FILL FILL_0__7167_ (
);

NAND2X1 _9273_ (
    .A(gnd),
    .B(\X[3] [4]),
    .Y(_2632_)
);

FILL FILL_3__10907_ (
);

FILL FILL_1__11941_ (
);

FILL FILL_1__11521_ (
);

FILL FILL_1__11101_ (
);

FILL FILL_2__8546_ (
);

FILL FILL_0__10934_ (
);

FILL FILL_0__10514_ (
);

OR2X2 _13271_ (
    .A(_6290_),
    .B(_6294_),
    .Y(_6295_)
);

FILL FILL_1__6963_ (
);

FILL FILL_1__6543_ (
);

FILL FILL_2__13313_ (
);

FILL FILL_3__6469_ (
);

FILL FILL_1__12726_ (
);

FILL FILL_1__12306_ (
);

FILL FILL_0__9733_ (
);

FILL FILL_0__9313_ (
);

FILL FILL_0__11719_ (
);

FILL FILL_1__7748_ (
);

FILL FILL_1__7328_ (
);

FILL FILL_3__10240_ (
);

INVX1 _6398_ (
    .A(_0_),
    .Y(_1_)
);

NAND2X1 _10396_ (
    .A(_3671_),
    .B(_3660_),
    .Y(_3672_)
);

FILL FILL_3__11865_ (
);

FILL FILL_2__6612_ (
);

FILL FILL_3__11025_ (
);

FILL FILL_2__10858_ (
);

FILL FILL_0__11892_ (
);

FILL FILL_2__10438_ (
);

FILL FILL_2__9084_ (
);

FILL FILL_0__11472_ (
);

FILL FILL_2__10018_ (
);

FILL FILL_0__11052_ (
);

FILL FILL_0__6858_ (
);

DFFPOSX1 _8964_ (
    .D(_2384_[11]),
    .CLK(clk_bF$buf47),
    .Q(\Y[3] [11])
);

FILL FILL_0__6438_ (
);

NOR2X1 _8544_ (
    .A(_1912_),
    .B(_1915_),
    .Y(_1981_)
);

DFFPOSX1 _8124_ (
    .D(_1593_[8]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.mul [8])
);

FILL FILL_1__7081_ (
);

FILL FILL_2__7817_ (
);

FILL FILL_1__13264_ (
);

NAND2X1 _12962_ (
    .A(_5982_),
    .B(_5992_),
    .Y(_5999_)
);

FILL FILL_0__12677_ (
);

FILL FILL_0__12257_ (
);

NAND3X1 _12542_ (
    .A(_5580_),
    .B(_5584_),
    .C(_5582_),
    .Y(_5585_)
);

AOI21X1 _12122_ (
    .A(_5223_),
    .B(_5219_),
    .C(_5164_),
    .Y(_5238_)
);

NAND3X1 _9749_ (
    .A(_3092_),
    .B(_3089_),
    .C(_3052_),
    .Y(_3093_)
);

AOI21X1 _9329_ (
    .A(_2598_),
    .B(_2676_),
    .C(_2684_),
    .Y(_2687_)
);

FILL FILL_1__8286_ (
);

FILL FILL_2__10191_ (
);

FILL FILL_3__9573_ (
);

NAND2X1 _13327_ (
    .A(_6348_),
    .B(_6350_),
    .Y(_6351_)
);

FILL FILL_2__7990_ (
);

FILL FILL_2__7570_ (
);

FILL FILL_2__7150_ (
);

FILL FILL_2__11396_ (
);

OAI21X1 _6610_ (
    .A(_136_),
    .B(_208_),
    .C(_177_),
    .Y(_209_)
);

FILL FILL_1__10389_ (
);

FILL FILL_0__7396_ (
);

AOI22X1 _9082_ (
    .A(_2400_),
    .B(_2405_),
    .C(_2440_),
    .D(_2443_),
    .Y(_2444_)
);

FILL FILL_1__11750_ (
);

FILL FILL_1__11330_ (
);

FILL FILL_2__8775_ (
);

FILL FILL_2__8355_ (
);

FILL FILL_0__10323_ (
);

AND2X2 _13080_ (
    .A(_6114_),
    .B(_6111_),
    .Y(_6115_)
);

AND2X2 _7815_ (
    .A(_1320_),
    .B(_1316_),
    .Y(_1330_)
);

FILL FILL_1__6772_ (
);

FILL FILL_2__13122_ (
);

FILL FILL_3__6698_ (
);

FILL FILL_1__12955_ (
);

FILL FILL_1__12535_ (
);

FILL FILL_1__12115_ (
);

FILL FILL_0__9962_ (
);

FILL FILL_0__9542_ (
);

FILL FILL_0__11948_ (
);

FILL FILL_0__9122_ (
);

NAND3X1 _11813_ (
    .A(_4921_),
    .B(_4930_),
    .C(_4932_),
    .Y(_4933_)
);

FILL FILL_0__11528_ (
);

FILL FILL_0__11108_ (
);

FILL FILL_1__7977_ (
);

FILL FILL_1__7557_ (
);

FILL FILL_1__7137_ (
);

FILL FILL_3__8424_ (
);

FILL FILL_2__6841_ (
);

FILL FILL_2__6421_ (
);

FILL FILL_3__11254_ (
);

FILL FILL_2__10667_ (
);

FILL FILL_2__10247_ (
);

FILL FILL_0__11281_ (
);

FILL FILL_1__9703_ (
);

FILL FILL_3__9209_ (
);

FILL FILL_0__6667_ (
);

AND2X2 _8773_ (
    .A(_2202_),
    .B(_2199_),
    .Y(_2206_)
);

AOI21X1 _8353_ (
    .A(_1780_),
    .B(_1779_),
    .C(_1730_),
    .Y(_1793_)
);

FILL FILL_1__10601_ (
);

FILL FILL_3__12879_ (
);

FILL FILL_2__7626_ (
);

FILL FILL_3__12459_ (
);

FILL FILL_3__12039_ (
);

FILL FILL_1__13073_ (
);

INVX1 _12771_ (
    .A(_5809_),
    .Y(_5810_)
);

FILL FILL_0__12066_ (
);

INVX1 _12351_ (
    .A(\u_fir_pe6.rYin [6]),
    .Y(_5455_)
);

FILL FILL_3__13400_ (
);

FILL FILL_2__12813_ (
);

INVX1 _9978_ (
    .A(_3258_),
    .Y(_3259_)
);

OAI21X1 _9558_ (
    .A(_2465_),
    .B(_2696_),
    .C(_2870_),
    .Y(_2913_)
);

AOI21X1 _9138_ (
    .A(_2494_),
    .B(_2495_),
    .C(_2493_),
    .Y(_2499_)
);

FILL FILL_1__11806_ (
);

FILL FILL_0__8813_ (
);

FILL FILL_3__6910_ (
);

NOR2X1 _13136_ (
    .A(_6165_),
    .B(_6169_),
    .Y(_6375_[12])
);

FILL FILL_1__6828_ (
);

FILL FILL_1__6408_ (
);

FILL FILL_1__10198_ (
);

FILL FILL_3__10105_ (
);

FILL FILL_2__8584_ (
);

FILL FILL_0__10972_ (
);

FILL FILL_2__8164_ (
);

FILL FILL_0__10552_ (
);

FILL FILL_0__10132_ (
);

AOI21X1 _7624_ (
    .A(_1141_),
    .B(_1140_),
    .C(_1139_),
    .Y(_1142_)
);

DFFPOSX1 _7204_ (
    .D(_790_[5]),
    .CLK(clk_bF$buf32),
    .Q(\Y[1] [5])
);

FILL FILL_1__6581_ (
);

FILL FILL_1__12764_ (
);

FILL FILL_1__12344_ (
);

FILL FILL_2__9789_ (
);

FILL FILL_0__9771_ (
);

FILL FILL_2__9369_ (
);

FILL FILL_0__9351_ (
);

FILL FILL_0__11757_ (
);

DFFPOSX1 _11622_ (
    .D(\Y[5] [14]),
    .CLK(clk_bF$buf18),
    .Q(\u_fir_pe5.rYin [14])
);

FILL FILL_0__11337_ (
);

NAND2X1 _11202_ (
    .A(_4398_),
    .B(_4394_),
    .Y(_4399_)
);

OAI21X1 _8829_ (
    .A(_2245_),
    .B(_2241_),
    .C(_2254_),
    .Y(_2255_)
);

NAND2X1 _8409_ (
    .A(gnd),
    .B(\X[2]_5_bF$buf0 ),
    .Y(_1848_)
);

FILL FILL_1__7786_ (
);

FILL FILL_1__7366_ (
);

FILL FILL_1__13129_ (
);

FILL FILL_3__8653_ (
);

NAND3X1 _12827_ (
    .A(_5714_),
    .B(_5853_),
    .C(_5858_),
    .Y(_5866_)
);

NAND2X1 _12407_ (
    .A(_5510_),
    .B(_5505_),
    .Y(_5511_)
);

FILL FILL_2__6650_ (
);

FILL FILL_3__11483_ (
);

FILL FILL_2__10896_ (
);

FILL FILL_2__10476_ (
);

FILL FILL_2__10056_ (
);

FILL FILL_0__11090_ (
);

FILL FILL_1__9932_ (
);

FILL FILL_1__9512_ (
);

FILL FILL_3__9438_ (
);

FILL FILL_0__6896_ (
);

FILL FILL_0__6476_ (
);

NAND3X1 _8582_ (
    .A(_1937_),
    .B(_1943_),
    .C(_2018_),
    .Y(_2019_)
);

NAND3X1 _8162_ (
    .A(_1594_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1605_)
);

FILL FILL_1__10830_ (
);

FILL FILL_1__10410_ (
);

FILL FILL_2__7855_ (
);

FILL FILL_2__7435_ (
);

FILL FILL_3__12268_ (
);

FILL FILL_2__7015_ (
);

NAND3X1 _12580_ (
    .A(vdd),
    .B(\X[6] [1]),
    .C(_5621_),
    .Y(_5622_)
);

FILL FILL_0__12295_ (
);

NAND3X1 _12160_ (
    .A(_5205_),
    .B(_5208_),
    .C(_5275_),
    .Y(_5276_)
);

FILL FILL_2__12622_ (
);

FILL FILL_2__12202_ (
);

NAND2X1 _9787_ (
    .A(_3126_),
    .B(_3119_),
    .Y(_3130_)
);

NAND2X1 _9367_ (
    .A(_2716_),
    .B(_2724_),
    .Y(_2725_)
);

FILL FILL_0__8622_ (
);

FILL FILL_0__8202_ (
);

FILL FILL_0__10608_ (
);

FILL FILL_3__9191_ (
);

DFFPOSX1 _13365_ (
    .D(\Y[6] [3]),
    .CLK(clk_bF$buf48),
    .Q(\u_fir_pe7.rYin [3])
);

FILL FILL_1__6637_ (
);

FILL FILL_2__13407_ (
);

FILL FILL_0__9827_ (
);

FILL FILL_3__7924_ (
);

FILL FILL_0__9407_ (
);

FILL FILL_3__10334_ (
);

FILL FILL_2__8393_ (
);

FILL FILL_0__10781_ (
);

FILL FILL_0__10361_ (
);

OR2X2 _7853_ (
    .A(_1366_),
    .B(_1362_),
    .Y(_1367_)
);

NAND2X1 _7433_ (
    .A(gnd),
    .B(\X[1]_5_bF$buf3 ),
    .Y(_953_)
);

OAI21X1 _7013_ (
    .A(_563_),
    .B(_576_),
    .C(_580_),
    .Y(_606_)
);

FILL FILL_1__6390_ (
);

FILL FILL_2__13160_ (
);

FILL FILL_3__11959_ (
);

FILL FILL_2__6706_ (
);

FILL FILL_1__12993_ (
);

FILL FILL_1__12573_ (
);

FILL FILL_3__11119_ (
);

FILL FILL_1__12153_ (
);

FILL FILL_0__11986_ (
);

FILL FILL_0__9580_ (
);

FILL FILL_2__9598_ (
);

FILL FILL_2__9178_ (
);

FILL FILL_0__9160_ (
);

AOI21X1 _11851_ (
    .A(_4883_),
    .B(_4887_),
    .C(_4851_),
    .Y(_4971_)
);

FILL FILL_0__11566_ (
);

NOR2X1 _11431_ (
    .A(\u_fir_pe5.rYin [1]),
    .B(\u_fir_pe5.mul [1]),
    .Y(_4620_)
);

FILL FILL_0__11146_ (
);

NAND2X1 _11011_ (
    .A(\X[5] [2]),
    .B(gnd),
    .Y(_4210_)
);

OAI21X1 _8638_ (
    .A(_1668_),
    .B(_1913_),
    .C(_2067_),
    .Y(_2074_)
);

OAI21X1 _8218_ (
    .A(_1647_),
    .B(_1659_),
    .C(_1653_),
    .Y(_1660_)
);

FILL FILL_1__7595_ (
);

FILL FILL_1__7175_ (
);

FILL FILL_3__8882_ (
);

AOI21X1 _12636_ (
    .A(_5671_),
    .B(_5673_),
    .C(_5664_),
    .Y(_5677_)
);

FILL FILL_3__8042_ (
);

AOI21X1 _12216_ (
    .A(_5269_),
    .B(_5273_),
    .C(_5243_),
    .Y(_5331_)
);

FILL FILL_2__10285_ (
);

FILL FILL_1__9741_ (
);

FILL FILL_1__9321_ (
);

FILL FILL_3__9667_ (
);

OAI21X1 _8391_ (
    .A(_2372_),
    .B(_1829_),
    .C(_1821_),
    .Y(_1830_)
);

FILL FILL_2__7664_ (
);

FILL FILL_3__12077_ (
);

AOI21X1 _6704_ (
    .A(_266_),
    .B(_267_),
    .C(_224_),
    .Y(_302_)
);

FILL FILL_2__12851_ (
);

FILL FILL_2__12431_ (
);

FILL FILL_2__12011_ (
);

AOI21X1 _9596_ (
    .A(_2947_),
    .B(_2848_),
    .C(_2949_),
    .Y(_2950_)
);

NAND2X1 _9176_ (
    .A(\X[3] [2]),
    .B(gnd),
    .Y(_2536_)
);

FILL FILL_1__11844_ (
);

FILL FILL_1__11424_ (
);

FILL FILL_1__11004_ (
);

FILL FILL_0__8851_ (
);

FILL FILL_2__8869_ (
);

FILL FILL_0__8431_ (
);

FILL FILL_2__8449_ (
);

FILL FILL_0__10837_ (
);

NOR2X1 _10702_ (
    .A(_3964_),
    .B(_3819_),
    .Y(_3977_[0])
);

FILL FILL_0__10417_ (
);

FILL FILL_0__8011_ (
);

FILL FILL_2__8029_ (
);

INVX1 _13174_ (
    .A(_6200_),
    .Y(_6206_)
);

FILL FILL_2__9810_ (
);

NOR3X1 _7909_ (
    .A(_1420_),
    .B(_1388_),
    .C(_1406_),
    .Y(_1421_)
);

FILL FILL_1__6866_ (
);

FILL FILL_1__6446_ (
);

FILL FILL_2__13216_ (
);

FILL FILL_1__12629_ (
);

FILL FILL_1__12209_ (
);

FILL FILL_0__9636_ (
);

FILL FILL_3__7733_ (
);

FILL FILL_0__9216_ (
);

OAI21X1 _11907_ (
    .A(_4871_),
    .B(_4856_),
    .C(_4940_),
    .Y(_5026_)
);

FILL FILL_3__7313_ (
);

FILL FILL_3__10983_ (
);

FILL FILL_3__10563_ (
);

FILL FILL_0__10590_ (
);

FILL FILL_0__10170_ (
);

FILL FILL_3__8518_ (
);

OAI21X1 _7662_ (
    .A(_1098_),
    .B(_1178_),
    .C(_1161_),
    .Y(_1179_)
);

DFFPOSX1 _7242_ (
    .D(_794_[3]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.mul [3])
);

NAND2X1 _10299_ (
    .A(gnd),
    .B(_3575_),
    .Y(_3576_)
);

FILL FILL_2__6935_ (
);

FILL FILL_2__6515_ (
);

FILL FILL_3__11348_ (
);

FILL FILL_1__12382_ (
);

FILL FILL_0__11795_ (
);

INVX1 _11660_ (
    .A(_4782_),
    .Y(_4783_)
);

FILL FILL_0__11375_ (
);

NAND2X1 _11240_ (
    .A(_4435_),
    .B(_4365_),
    .Y(_4437_)
);

FILL FILL_2__11702_ (
);

NAND2X1 _8867_ (
    .A(_2269_),
    .B(_2281_),
    .Y(_2290_)
);

AOI21X1 _8447_ (
    .A(_1881_),
    .B(_1880_),
    .C(_1782_),
    .Y(_1886_)
);

NOR2X1 _8027_ (
    .A(\u_fir_pe1.rYin [11]),
    .B(\u_fir_pe1.mul [11]),
    .Y(_1531_)
);

FILL FILL_0__7702_ (
);

FILL FILL_1__13167_ (
);

NAND2X1 _12865_ (
    .A(gnd),
    .B(\X[6] [7]),
    .Y(_5903_)
);

FILL FILL_3__8271_ (
);

NOR2X1 _12445_ (
    .A(_5548_),
    .B(_5547_),
    .Y(_5572_[14])
);

NAND3X1 _12025_ (
    .A(_5097_),
    .B(_5128_),
    .C(_5133_),
    .Y(_5143_)
);

FILL FILL_2__12907_ (
);

FILL FILL_0__13101_ (
);

FILL FILL_1__8189_ (
);

FILL FILL_0__8907_ (
);

FILL FILL_2__10094_ (
);

FILL FILL_1__9970_ (
);

FILL FILL_1__9550_ (
);

FILL FILL_1__9130_ (
);

FILL FILL_3__9896_ (
);

FILL FILL_3__9056_ (
);

FILL FILL_2__7893_ (
);

FILL FILL_2__7473_ (
);

FILL FILL_2__7053_ (
);

FILL FILL_2__11299_ (
);

OAI21X1 _6933_ (
    .A(_473_),
    .B(_526_),
    .C(_527_),
    .Y(_528_)
);

NAND3X1 _6513_ (
    .A(_101_),
    .B(_105_),
    .C(_107_),
    .Y(_114_)
);

FILL FILL_2__12660_ (
);

FILL FILL_2__12240_ (
);

FILL FILL_0__7299_ (
);

FILL FILL_1__11653_ (
);

FILL FILL_1__11233_ (
);

FILL FILL_2__8678_ (
);

FILL FILL_0__8660_ (
);

FILL FILL_0__8240_ (
);

FILL FILL_2__8258_ (
);

FILL FILL_0__10646_ (
);

OAI21X1 _10931_ (
    .A(_4763_),
    .B(_4129_),
    .C(_4130_),
    .Y(_4131_)
);

NAND2X1 _10511_ (
    .A(_3755_),
    .B(_3783_),
    .Y(_3784_)
);

FILL FILL_0__10226_ (
);

INVX1 _7718_ (
    .A(_1180_),
    .Y(_1235_)
);

FILL FILL_1__6675_ (
);

FILL FILL_2__13025_ (
);

FILL FILL_1__12858_ (
);

FILL FILL_1__12438_ (
);

FILL FILL_1__12018_ (
);

FILL FILL_0_BUFX2_insert0 (
);

FILL FILL_0_BUFX2_insert1 (
);

FILL FILL_0_BUFX2_insert2 (
);

FILL FILL_3__7962_ (
);

FILL FILL_0_BUFX2_insert3 (
);

FILL FILL_0__9445_ (
);

FILL FILL_0_BUFX2_insert4 (
);

FILL FILL_3__7542_ (
);

FILL FILL_0_BUFX2_insert5 (
);

FILL FILL_0__9025_ (
);

NAND2X1 _11716_ (
    .A(_4831_),
    .B(_4834_),
    .Y(_4838_)
);

FILL FILL_3__7122_ (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_1__8821_ (
);

FILL FILL_1__8401_ (
);

FILL FILL_3__8747_ (
);

AND2X2 _7891_ (
    .A(_1400_),
    .B(_1399_),
    .Y(_1404_)
);

OAI21X1 _7471_ (
    .A(_990_),
    .B(_985_),
    .C(_913_),
    .Y(_991_)
);

NOR2X1 _7051_ (
    .A(_639_),
    .B(_638_),
    .Y(_790_[1])
);

FILL FILL_2__6744_ (
);

FILL FILL_3__11577_ (
);

FILL FILL_1__12191_ (
);

FILL FILL_0__11184_ (
);

FILL FILL_1__9606_ (
);

FILL FILL_2__11931_ (
);

FILL FILL_2__11511_ (
);

NOR3X1 _8676_ (
    .A(_1899_),
    .B(_2067_),
    .C(_2010_),
    .Y(_2111_)
);

OAI21X1 _8256_ (
    .A(_1692_),
    .B(_1693_),
    .C(_1678_),
    .Y(_1697_)
);

FILL FILL_1__10924_ (
);

FILL FILL_1__10504_ (
);

FILL FILL_0__7931_ (
);

FILL FILL_2__7949_ (
);

FILL FILL_0__7511_ (
);

FILL FILL_2__7529_ (
);

FILL FILL_2__7109_ (
);

FILL FILL_1__13396_ (
);

NAND2X1 _12674_ (
    .A(_5710_),
    .B(_5712_),
    .Y(_5714_)
);

FILL FILL_0__12389_ (
);

AOI21X1 _12254_ (
    .A(_5339_),
    .B(_5341_),
    .C(_5367_),
    .Y(_5368_)
);

FILL FILL_3__13303_ (
);

FILL FILL_2__12716_ (
);

FILL FILL_0__13330_ (
);

FILL FILL_1__11709_ (
);

FILL FILL_0__8716_ (
);

FILL FILL_3__9285_ (
);

INVX1 _13039_ (
    .A(_6039_),
    .Y(_6075_)
);

FILL FILL_2__7282_ (
);

NAND3X1 _6742_ (
    .A(_338_),
    .B(_339_),
    .C(_337_),
    .Y(_340_)
);

FILL FILL_3__10848_ (
);

FILL FILL_1__11882_ (
);

FILL FILL_3__10428_ (
);

FILL FILL_1__11462_ (
);

FILL FILL_3__10008_ (
);

FILL FILL_1__11042_ (
);

FILL FILL_2__8487_ (
);

FILL FILL_0__10875_ (
);

DFFPOSX1 _10740_ (
    .D(\Y[4] [9]),
    .CLK(clk_bF$buf55),
    .Q(\u_fir_pe4.rYin [9])
);

FILL FILL_0__10455_ (
);

FILL FILL_2__8067_ (
);

AOI22X1 _10320_ (
    .A(_3430_),
    .B(_3596_),
    .C(_3522_),
    .D(_3518_),
    .Y(_3597_)
);

FILL FILL_0__10035_ (
);

INVX1 _7947_ (
    .A(\u_fir_pe1.mul [4]),
    .Y(_1453_)
);

INVX1 _7527_ (
    .A(_1045_),
    .Y(_1046_)
);

INVX1 _7107_ (
    .A(\u_fir_pe0.rYin [8]),
    .Y(_690_)
);

FILL FILL_1__6484_ (
);

FILL FILL_2__13254_ (
);

FILL FILL_1__12667_ (
);

FILL FILL_1__12247_ (
);

FILL FILL_0__9674_ (
);

FILL FILL_0__9254_ (
);

NAND3X1 _11945_ (
    .A(_4991_),
    .B(_5059_),
    .C(_5060_),
    .Y(_5064_)
);

FILL FILL_3__7351_ (
);

INVX1 _11525_ (
    .A(\u_fir_pe5.rYin [10]),
    .Y(_4709_)
);

NAND2X1 _11105_ (
    .A(\X[5] [3]),
    .B(vdd),
    .Y(_4303_)
);

FILL FILL_0__12601_ (
);

FILL FILL_1__7689_ (
);

FILL FILL_1__7269_ (
);

FILL FILL_3__10181_ (
);

FILL FILL_1__8630_ (
);

FILL FILL_1__8210_ (
);

FILL FILL_3__8136_ (
);

NAND3X1 _7280_ (
    .A(_798_),
    .B(_802_),
    .C(_800_),
    .Y(_803_)
);

FILL FILL_2__6973_ (
);

FILL FILL_2__6553_ (
);

FILL FILL_2__10799_ (
);

FILL FILL_2__10379_ (
);

FILL FILL_1__9415_ (
);

FILL FILL_2__11740_ (
);

FILL FILL_0__6799_ (
);

FILL FILL_2__11320_ (
);

FILL FILL_0__6379_ (
);

AOI21X1 _8485_ (
    .A(_1922_),
    .B(_1920_),
    .C(_1918_),
    .Y(_1923_)
);

NAND2X1 _8065_ (
    .A(_1566_),
    .B(_1568_),
    .Y(_1569_)
);

FILL FILL_1__10313_ (
);

FILL FILL_2__7758_ (
);

FILL FILL_0__7740_ (
);

FILL FILL_2__7338_ (
);

FILL FILL_0__7320_ (
);

DFFPOSX1 _12483_ (
    .D(\X[7] [6]),
    .CLK(clk_bF$buf37),
    .Q(_6376_[6])
);

FILL FILL_0__12198_ (
);

NOR2X1 _12063_ (
    .A(_4914_),
    .B(_5103_),
    .Y(_5180_)
);

FILL FILL_2__12945_ (
);

FILL FILL_2__12525_ (
);

FILL FILL_2__12105_ (
);

FILL FILL_1__11938_ (
);

FILL FILL_1__11518_ (
);

FILL FILL_0__8945_ (
);

FILL FILL_0__8525_ (
);

FILL FILL_3__6622_ (
);

NOR2X1 _13268_ (
    .A(\u_fir_pe7.rYin [9]),
    .B(\u_fir_pe7.mul [9]),
    .Y(_6292_)
);

FILL FILL_2__9904_ (
);

FILL FILL_2__7091_ (
);

FILL FILL_1__7901_ (
);

FILL FILL_3__7407_ (
);

NOR2X1 _6971_ (
    .A(_74_),
    .B(_462_),
    .Y(_565_)
);

NAND3X1 _6551_ (
    .A(_139_),
    .B(_148_),
    .C(_150_),
    .Y(_151_)
);

FILL FILL_3__10657_ (
);

FILL FILL_1__11691_ (
);

FILL FILL_1__11271_ (
);

FILL FILL_2__8296_ (
);

FILL FILL_0__10684_ (
);

FILL FILL_0__10264_ (
);

AND2X2 _7756_ (
    .A(_1270_),
    .B(_1213_),
    .Y(_1272_)
);

NAND3X1 _7336_ (
    .A(_825_),
    .B(_842_),
    .C(_845_),
    .Y(_858_)
);

FILL FILL_2__13063_ (
);

FILL FILL_2__6609_ (
);

FILL FILL_1__12896_ (
);

FILL FILL_1__12056_ (
);

FILL FILL_0__9483_ (
);

FILL FILL_0__11889_ (
);

FILL FILL_3__7580_ (
);

FILL FILL_0__9063_ (
);

NAND2X1 _11754_ (
    .A(vdd),
    .B(\X[7] [3]),
    .Y(_4875_)
);

FILL FILL_0__11469_ (
);

FILL FILL_0__11049_ (
);

NAND2X1 _11334_ (
    .A(_4525_),
    .B(_4501_),
    .Y(_4529_)
);

FILL FILL_3__12803_ (
);

FILL FILL_0__12830_ (
);

FILL FILL_0__12410_ (
);

FILL FILL_1__7498_ (
);

FILL FILL_1__7078_ (
);

INVX1 _9902_ (
    .A(_3973_),
    .Y(_3974_)
);

INVX1 _12959_ (
    .A(\X[6] [4]),
    .Y(_5996_)
);

FILL FILL_3__8365_ (
);

OR2X2 _12539_ (
    .A(_6310_),
    .B(_5581_),
    .Y(_5582_)
);

NAND2X1 _12119_ (
    .A(_5224_),
    .B(_5231_),
    .Y(_5235_)
);

FILL FILL_2__6782_ (
);

FILL FILL_3__11195_ (
);

FILL FILL_2__10188_ (
);

FILL FILL_1__9644_ (
);

FILL FILL_1__9224_ (
);

INVX1 _8294_ (
    .A(_1733_),
    .Y(_1734_)
);

FILL FILL_1__10962_ (
);

FILL FILL_1__10542_ (
);

FILL FILL_1__10122_ (
);

FILL FILL_2__7987_ (
);

FILL FILL_2__7567_ (
);

FILL FILL_2__7147_ (
);

OAI21X1 _12292_ (
    .A(_5398_),
    .B(_5397_),
    .C(_5403_),
    .Y(_5404_)
);

NOR2X1 _6607_ (
    .A(_204_),
    .B(_206_),
    .Y(_796_[6])
);

FILL FILL_2__12754_ (
);

FILL FILL_2__12334_ (
);

OAI22X1 _9499_ (
    .A(_2808_),
    .B(_2696_),
    .C(_2416_),
    .D(_2807_),
    .Y(_2855_)
);

NAND2X1 _9079_ (
    .A(_2423_),
    .B(_2438_),
    .Y(_2441_)
);

FILL FILL_1__11747_ (
);

FILL FILL_1__11327_ (
);

FILL FILL_0__8754_ (
);

FILL FILL_3__6851_ (
);

FILL FILL_0__8334_ (
);

OAI21X1 _10605_ (
    .A(_3861_),
    .B(_3862_),
    .C(_3866_),
    .Y(_3868_)
);

FILL FILL_0_BUFX2_insert80 (
);

FILL FILL_0_BUFX2_insert81 (
);

FILL FILL_0_BUFX2_insert82 (
);

FILL FILL_0_BUFX2_insert83 (
);

FILL FILL_0_BUFX2_insert84 (
);

FILL FILL_0_BUFX2_insert85 (
);

FILL FILL_0_BUFX2_insert86 (
);

FILL FILL_0_BUFX2_insert87 (
);

AND2X2 _13077_ (
    .A(_6102_),
    .B(_6098_),
    .Y(_6112_)
);

FILL FILL_0_BUFX2_insert88 (
);

FILL FILL_0_BUFX2_insert89 (
);

FILL FILL_2__9713_ (
);

FILL FILL_1__6769_ (
);

FILL FILL_2__13119_ (
);

FILL FILL_1__7710_ (
);

FILL FILL_0__9959_ (
);

FILL FILL_0__9539_ (
);

FILL FILL_3__7636_ (
);

FILL FILL_0__9119_ (
);

NAND2X1 _6780_ (
    .A(_377_),
    .B(_376_),
    .Y(_378_)
);

FILL FILL_3__10046_ (
);

FILL FILL_1__11080_ (
);

FILL FILL_0__10493_ (
);

FILL FILL_0__10073_ (
);

FILL FILL_1__8915_ (
);

FILL FILL_2__10820_ (
);

FILL FILL_2__10400_ (
);

INVX1 _7985_ (
    .A(\u_fir_pe1.mul [8]),
    .Y(_1488_)
);

NAND3X1 _7565_ (
    .A(_932_),
    .B(_1071_),
    .C(_1076_),
    .Y(_1084_)
);

NAND2X1 _7145_ (
    .A(_728_),
    .B(_723_),
    .Y(_729_)
);

FILL FILL_2__13292_ (
);

FILL FILL_0__6820_ (
);

FILL FILL_2__6838_ (
);

FILL FILL_0__6400_ (
);

FILL FILL_2__6418_ (
);

FILL FILL_1__12285_ (
);

FILL FILL253650x43350 (
);

FILL FILL_0__9292_ (
);

INVX1 _11983_ (
    .A(gnd),
    .Y(_5101_)
);

FILL FILL_0__11698_ (
);

NOR2X1 _11563_ (
    .A(_4744_),
    .B(_4746_),
    .Y(_4747_)
);

FILL FILL_0__11278_ (
);

AOI21X1 _11143_ (
    .A(_4340_),
    .B(_4339_),
    .C(_4338_),
    .Y(_4341_)
);

FILL FILL_0__7605_ (
);

INVX1 _9711_ (
    .A(\u_fir_pe3.rYin [5]),
    .Y(_3056_)
);

FILL FILL_3__8594_ (
);

AND2X2 _12768_ (
    .A(gnd),
    .B(\X[6] [7]),
    .Y(_5807_)
);

OR2X2 _12348_ (
    .A(_5446_),
    .B(_5451_),
    .Y(_5453_)
);

FILL FILL_0__13004_ (
);

FILL FILL_2__6591_ (
);

FILL FILL254550x194550 (
);

FILL FILL_1__9453_ (
);

FILL FILL_1__9033_ (
);

FILL FILL_3__9379_ (
);

FILL FILL_1__10771_ (
);

FILL FILL_1__10351_ (
);

FILL FILL_2__7796_ (
);

FILL FILL_2__7376_ (
);

FILL FILL_3__13150_ (
);

AOI21X1 _6836_ (
    .A(_353_),
    .B(_355_),
    .C(_432_),
    .Y(_433_)
);

NAND2X1 _6416_ (
    .A(_781_),
    .B(_18_),
    .Y(_19_)
);

FILL FILL_2__12983_ (
);

FILL FILL_2__12563_ (
);

FILL FILL_2__12143_ (
);

FILL FILL_1__11976_ (
);

FILL FILL_1__11556_ (
);

FILL FILL_1__11136_ (
);

FILL FILL_0__8563_ (
);

FILL FILL_0__10969_ (
);

FILL FILL_0__8143_ (
);

FILL FILL_0__10549_ (
);

NAND3X1 _10834_ (
    .A(_4025_),
    .B(_4029_),
    .C(_4031_),
    .Y(_4036_)
);

AOI21X1 _10414_ (
    .A(_3683_),
    .B(_3689_),
    .C(_3647_),
    .Y(_3690_)
);

FILL FILL_0__10129_ (
);

FILL FILL_2__9942_ (
);

FILL FILL_0__11910_ (
);

FILL FILL_2__9522_ (
);

FILL FILL_2__9102_ (
);

FILL FILL_1__6998_ (
);

FILL FILL_1__6578_ (
);

FILL FILL_0__9768_ (
);

FILL FILL_0__9348_ (
);

DFFPOSX1 _11619_ (
    .D(\Y[5] [11]),
    .CLK(clk_bF$buf35),
    .Q(\u_fir_pe5.rYin [11])
);

FILL FILL_3__10275_ (
);

FILL FILL_2_BUFX2_insert0 (
);

FILL FILL_2_BUFX2_insert1 (
);

FILL FILL_2_BUFX2_insert2 (
);

FILL FILL_2_BUFX2_insert3 (
);

FILL FILL_2_BUFX2_insert4 (
);

FILL FILL_2_BUFX2_insert5 (
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_1__8724_ (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_1__8304_ (
);

FILL FILL_2_BUFX2_insert9 (
);

NAND2X1 _7794_ (
    .A(_1302_),
    .B(_1306_),
    .Y(_1309_)
);

AOI21X1 _7374_ (
    .A(_889_),
    .B(_891_),
    .C(_882_),
    .Y(_895_)
);

FILL FILL_2__6647_ (
);

FILL FILL_1__12094_ (
);

AND2X2 _11792_ (
    .A(_4912_),
    .B(_4908_),
    .Y(_5578_[5])
);

FILL FILL_0__11087_ (
);

INVX1 _11372_ (
    .A(_4565_),
    .Y(_4566_)
);

FILL FILL_1__9929_ (
);

FILL FILL_1__9509_ (
);

FILL FILL_3__12421_ (
);

FILL FILL_2__11834_ (
);

FILL FILL_2__11414_ (
);

DFFPOSX1 _8999_ (
    .D(_2390_[6]),
    .CLK(clk_bF$buf51),
    .Q(\u_fir_pe2.mul [6])
);

NAND3X1 _8579_ (
    .A(_2013_),
    .B(_2014_),
    .C(_2015_),
    .Y(_2016_)
);

OAI21X1 _8159_ (
    .A(_1598_),
    .B(_1601_),
    .C(_1594_),
    .Y(_1602_)
);

FILL FILL_1__10827_ (
);

FILL FILL_1__10407_ (
);

FILL FILL_0__7834_ (
);

INVX1 _9940_ (
    .A(_3221_),
    .Y(_3222_)
);

FILL FILL_0__7414_ (
);

NAND2X1 _9520_ (
    .A(_2873_),
    .B(_2867_),
    .Y(_2876_)
);

NAND2X1 _9100_ (
    .A(\X[3] [0]),
    .B(vdd),
    .Y(_2461_)
);

FILL FILL_1__13299_ (
);

NOR2X1 _12997_ (
    .A(_5952_),
    .B(_6032_),
    .Y(_6033_)
);

NAND3X1 _12577_ (
    .A(_5613_),
    .B(_5618_),
    .C(_5616_),
    .Y(_5619_)
);

NAND3X1 _12157_ (
    .A(_5270_),
    .B(_5272_),
    .C(_5271_),
    .Y(_5273_)
);

FILL FILL_3__13206_ (
);

FILL FILL_2__12619_ (
);

FILL FILL_0__13233_ (
);

FILL FILL_0__8619_ (
);

FILL FILL_3__6716_ (
);

FILL FILL_1__9682_ (
);

FILL FILL_1__9262_ (
);

FILL FILL_1__10580_ (
);

FILL FILL_1__10160_ (
);

FILL FILL_2__7185_ (
);

OAI21X1 _6645_ (
    .A(_89_),
    .B(_74_),
    .C(_158_),
    .Y(_244_)
);

FILL FILL_2__12792_ (
);

FILL FILL_2__12372_ (
);

FILL FILL_1__11785_ (
);

FILL FILL_1__11365_ (
);

FILL FILL_0__8792_ (
);

FILL FILL_0__8372_ (
);

FILL FILL_0__10778_ (
);

FILL FILL_0__10358_ (
);

NOR2X1 _10643_ (
    .A(_3903_),
    .B(_3897_),
    .Y(_3906_)
);

NAND2X1 _10223_ (
    .A(_3494_),
    .B(_3495_),
    .Y(_3501_)
);

FILL FILL_2__9751_ (
);

FILL FILL_2__9331_ (
);

FILL FILL_1__6387_ (
);

FILL FILL_2__13157_ (
);

FILL FILL_0__9997_ (
);

FILL FILL_0__9577_ (
);

FILL FILL_3__7674_ (
);

FILL FILL_0__9157_ (
);

NAND3X1 _11848_ (
    .A(_4954_),
    .B(_4958_),
    .C(_4961_),
    .Y(_4968_)
);

INVX1 _11428_ (
    .A(\u_fir_pe5.rYin [1]),
    .Y(_4617_)
);

NAND2X1 _11008_ (
    .A(_4203_),
    .B(_4206_),
    .Y(_4207_)
);

FILL FILL_0__12924_ (
);

FILL FILL_1__8533_ (
);

FILL FILL_3__8459_ (
);

NOR2X1 _7183_ (
    .A(_766_),
    .B(_765_),
    .Y(_790_[14])
);

FILL FILL253950x237750 (
);

FILL FILL_3__9820_ (
);

FILL FILL_2__6876_ (
);

FILL FILL_2__6456_ (
);

FILL FILL_3__11289_ (
);

INVX1 _11181_ (
    .A(_4375_),
    .Y(_4378_)
);

FILL FILL_1__9738_ (
);

FILL FILL_1__9318_ (
);

FILL FILL_3__12650_ (
);

FILL FILL_2__11643_ (
);

FILL FILL_2__11223_ (
);

INVX1 _8388_ (
    .A(vdd),
    .Y(_1827_)
);

FILL FILL_1__10636_ (
);

FILL FILL_1__10216_ (
);

FILL FILL_0__7643_ (
);

NAND2X1 _12386_ (
    .A(_5486_),
    .B(_5489_),
    .Y(_5572_[8])
);

FILL FILL_2__8602_ (
);

FILL FILL_2__12848_ (
);

FILL FILL_2__12428_ (
);

FILL FILL_2__12008_ (
);

FILL FILL_0__13042_ (
);

FILL FILL_0__8848_ (
);

FILL FILL_3__6945_ (
);

FILL FILL_0__8428_ (
);

FILL FILL_0__8008_ (
);

FILL FILL_1__9491_ (
);

FILL FILL_1__9071_ (
);

FILL FILL_2__9807_ (
);

FILL FILL_1__7804_ (
);

FILL FILL254250x180150 (
);

AND2X2 _6874_ (
    .A(_466_),
    .B(_469_),
    .Y(_470_)
);

NAND2X1 _6454_ (
    .A(_49_),
    .B(_52_),
    .Y(_56_)
);

FILL FILL_2__12181_ (
);

FILL FILL_1__11174_ (
);

FILL FILL_2__8199_ (
);

FILL FILL_0__8181_ (
);

FILL FILL_0__10587_ (
);

NAND2X1 _10872_ (
    .A(_4021_),
    .B(_4072_),
    .Y(_4073_)
);

AOI21X1 _10452_ (
    .A(_3658_),
    .B(_3674_),
    .C(_3726_),
    .Y(_3727_)
);

FILL FILL_0__10167_ (
);

NAND3X1 _10032_ (
    .A(_3311_),
    .B(_3312_),
    .C(_3310_),
    .Y(_3313_)
);

FILL FILL_3__11921_ (
);

FILL FILL_3__11501_ (
);

FILL FILL_2__10914_ (
);

FILL FILL_2__9980_ (
);

FILL FILL_2__9560_ (
);

FILL FILL_2__9140_ (
);

INVX1 _7659_ (
    .A(_1169_),
    .Y(_1176_)
);

DFFPOSX1 _7239_ (
    .D(_791_[0]),
    .CLK(clk_bF$buf16),
    .Q(\u_fir_pe0.mul [0])
);

FILL FILL_0__6914_ (
);

FILL FILL_1__12799_ (
);

INVX1 _8600_ (
    .A(_1958_),
    .Y(_2037_)
);

FILL FILL_1__12379_ (
);

FILL FILL_0__9386_ (
);

FILL FILL_3__7483_ (
);

NAND2X1 _11657_ (
    .A(gnd),
    .B(\X[7] [3]),
    .Y(_5569_)
);

FILL FILL_3__7063_ (
);

OAI21X1 _11237_ (
    .A(_4432_),
    .B(_4433_),
    .C(_4429_),
    .Y(_4434_)
);

FILL FILL_3__12706_ (
);

FILL FILL_1__13320_ (
);

FILL FILL253950x86550 (
);

FILL FILL_0__12733_ (
);

FILL FILL_0__12313_ (
);

AND2X2 _9805_ (
    .A(_3148_),
    .B(_3147_),
    .Y(_3181_[13])
);

FILL FILL_1__8762_ (
);

FILL FILL_1__8342_ (
);

FILL FILL_3__8688_ (
);

FILL FILL_2__6685_ (
);

FILL FILL_1__9967_ (
);

FILL FILL_1__9547_ (
);

FILL FILL_1__9127_ (
);

FILL FILL_2__11872_ (
);

FILL FILL_2__11452_ (
);

FILL FILL_2__11032_ (
);

NAND3X1 _8197_ (
    .A(_1626_),
    .B(_1638_),
    .C(_1634_),
    .Y(_1639_)
);

FILL FILL_1__10865_ (
);

FILL FILL_1__10445_ (
);

FILL FILL_1__10025_ (
);

FILL FILL_0__7872_ (
);

FILL FILL_0__7452_ (
);

FILL FILL_0__7032_ (
);

OAI21X1 _12195_ (
    .A(_5255_),
    .B(_5308_),
    .C(_5309_),
    .Y(_5310_)
);

FILL FILL_2__8831_ (
);

FILL FILL_2__8411_ (
);

FILL FILL_3__13244_ (
);

FILL FILL_2__12657_ (
);

FILL FILL_2__12237_ (
);

FILL FILL_0__13271_ (
);

FILL FILL_0__8657_ (
);

FILL FILL_0__8237_ (
);

NAND2X1 _10928_ (
    .A(_4126_),
    .B(_4127_),
    .Y(_4128_)
);

OAI21X1 _10508_ (
    .A(_3493_),
    .B(_3780_),
    .C(_3759_),
    .Y(_3781_)
);

FILL FILL_2__9616_ (
);

FILL FILL_1__7613_ (
);

FILL FILL_3__7959_ (
);

NAND3X1 _6683_ (
    .A(_209_),
    .B(_277_),
    .C(_278_),
    .Y(_282_)
);

FILL FILL_3__8900_ (
);

FILL FILL_3__10789_ (
);

FILL FILL_3__10369_ (
);

FILL FILL_0__10396_ (
);

OR2X2 _10681_ (
    .A(_3937_),
    .B(_3943_),
    .Y(_3945_)
);

NAND3X1 _10261_ (
    .A(_3537_),
    .B(_3538_),
    .C(_3536_),
    .Y(_3539_)
);

FILL FILL_1__8818_ (
);

FILL FILL_2__10303_ (
);

NAND2X1 _7888_ (
    .A(_1399_),
    .B(_1400_),
    .Y(_1401_)
);

NAND3X1 _7468_ (
    .A(_981_),
    .B(_974_),
    .C(_979_),
    .Y(_988_)
);

NAND2X1 _7048_ (
    .A(_631_),
    .B(_636_),
    .Y(_637_)
);

FILL FILL_2__13195_ (
);

FILL FILL_0__6723_ (
);

FILL FILL_1__12188_ (
);

FILL FILL_0__9195_ (
);

AOI21X1 _11886_ (
    .A(_4944_),
    .B(_4948_),
    .C(_4937_),
    .Y(_5005_)
);

FILL FILL_3__7292_ (
);

INVX1 _11466_ (
    .A(\u_fir_pe5.mul [5]),
    .Y(_4651_)
);

NAND3X1 _11046_ (
    .A(_4224_),
    .B(_4238_),
    .C(_4241_),
    .Y(_4245_)
);

FILL FILL_2__11928_ (
);

FILL FILL_0__12962_ (
);

FILL FILL_2__11508_ (
);

FILL FILL_0__12542_ (
);

FILL FILL_0__12122_ (
);

FILL FILL_0__7928_ (
);

FILL FILL_0__7508_ (
);

NAND2X1 _9614_ (
    .A(_2954_),
    .B(_2967_),
    .Y(_2968_)
);

FILL FILL253050x230550 (
);

FILL FILL_1__8571_ (
);

FILL FILL_1__8151_ (
);

FILL FILL_0__13327_ (
);

FILL FILL_2__6494_ (
);

FILL FILL_1__9776_ (
);

FILL FILL_1__9356_ (
);

FILL FILL_2__11681_ (
);

FILL FILL_2__11261_ (
);

FILL FILL_1__10674_ (
);

FILL FILL_1__10254_ (
);

FILL FILL_2__7699_ (
);

FILL FILL_0__7681_ (
);

FILL FILL_0__7261_ (
);

FILL FILL_2__7279_ (
);

FILL FILL_2__8640_ (
);

FILL FILL_2__8220_ (
);

AOI21X1 _6739_ (
    .A(_246_),
    .B(_249_),
    .C(_255_),
    .Y(_337_)
);

FILL FILL_2__12886_ (
);

FILL FILL_2__12046_ (
);

FILL FILL_0__13080_ (
);

FILL FILL_1__11879_ (
);

FILL FILL_1__11459_ (
);

FILL FILL_1__11039_ (
);

FILL FILL_0__8886_ (
);

FILL FILL_0__8466_ (
);

FILL FILL_3__6563_ (
);

DFFPOSX1 _10737_ (
    .D(\Y[4] [6]),
    .CLK(clk_bF$buf7),
    .Q(\u_fir_pe4.rYin [6])
);

FILL FILL_0__8046_ (
);

AOI21X1 _10317_ (
    .A(_3519_),
    .B(_3593_),
    .C(_3592_),
    .Y(_3594_)
);

FILL FILL_1__12820_ (
);

FILL FILL_1__12400_ (
);

FILL FILL_2__9425_ (
);

FILL FILL_0__11813_ (
);

FILL FILL_1__7842_ (
);

FILL FILL_1__7422_ (
);

FILL FILL_1__7002_ (
);

FILL FILL_3__7348_ (
);

NAND2X1 _6492_ (
    .A(vdd),
    .B(Xin[3]),
    .Y(_93_)
);

FILL FILL_3__10598_ (
);

NAND2X1 _10490_ (
    .A(_3760_),
    .B(_3763_),
    .Y(_3764_)
);

NAND3X1 _10070_ (
    .A(_3345_),
    .B(_3349_),
    .C(_3347_),
    .Y(_3350_)
);

FILL FILL_1__8627_ (
);

FILL FILL_1__8207_ (
);

FILL FILL_2__10952_ (
);

FILL FILL_2__10532_ (
);

FILL FILL_2__10112_ (
);

INVX1 _7697_ (
    .A(\X[1] [4]),
    .Y(_1214_)
);

OR2X2 _7277_ (
    .A(_1528_),
    .B(_799_),
    .Y(_800_)
);

FILL FILL_0__6952_ (
);

FILL FILL_0__6532_ (
);

AND2X2 _11695_ (
    .A(vdd),
    .B(\X[7] [1]),
    .Y(_4817_)
);

NAND3X1 _11275_ (
    .A(_4392_),
    .B(_4470_),
    .C(_4400_),
    .Y(_4471_)
);

FILL FILL_2__7911_ (
);

FILL FILL_3__12744_ (
);

FILL FILL_2__11737_ (
);

FILL FILL_0__12771_ (
);

FILL FILL_2__11317_ (
);

FILL FILL_0__12351_ (
);

FILL FILL_0__7737_ (
);

DFFPOSX1 _9843_ (
    .D(_3181_[13]),
    .CLK(clk_bF$buf12),
    .Q(\Y[4] [13])
);

FILL FILL_0__7317_ (
);

INVX1 _9423_ (
    .A(_2779_),
    .Y(_2780_)
);

DFFPOSX1 _9003_ (
    .D(_2390_[10]),
    .CLK(clk_bF$buf51),
    .Q(\u_fir_pe2.mul [10])
);

FILL FILL_1__8380_ (
);

FILL FILL_0__13136_ (
);

INVX1 _13001_ (
    .A(_6036_),
    .Y(_6037_)
);

FILL FILL_1__9585_ (
);

FILL FILL_1__9165_ (
);

FILL FILL_2__11490_ (
);

FILL FILL_2__11070_ (
);

FILL FILL_1__10483_ (
);

FILL FILL_1__10063_ (
);

FILL FILL254550x126150 (
);

FILL FILL_0__7490_ (
);

FILL FILL_2__7088_ (
);

FILL FILL_0__7070_ (
);

OAI21X1 _6968_ (
    .A(_530_),
    .B(_524_),
    .C(_534_),
    .Y(_562_)
);

NAND3X1 _6548_ (
    .A(gnd),
    .B(Xin[6]),
    .C(_145_),
    .Y(_148_)
);

FILL FILL_2__12695_ (
);

FILL FILL_2__12275_ (
);

FILL FILL_1__11688_ (
);

FILL FILL_1__11268_ (
);

FILL FILL_0__8695_ (
);

FILL FILL_3__6792_ (
);

FILL FILL_0__8275_ (
);

AOI21X1 _10966_ (
    .A(_4156_),
    .B(_4152_),
    .C(_4137_),
    .Y(_4166_)
);

OAI21X1 _10546_ (
    .A(_3804_),
    .B(_3803_),
    .C(_3815_),
    .Y(_3817_)
);

NAND3X1 _10126_ (
    .A(_3331_),
    .B(_3400_),
    .C(_3335_),
    .Y(_3405_)
);

FILL FILL_2__9654_ (
);

FILL FILL_2__9234_ (
);

FILL FILL_0__11202_ (
);

FILL FILL_1__7651_ (
);

FILL FILL_3__7997_ (
);

FILL FILL_3__7577_ (
);

FILL FILL_3__7157_ (
);

FILL FILL_1__13414_ (
);

FILL FILL_0__12827_ (
);

FILL FILL_0__12407_ (
);

FILL FILL_1__8856_ (
);

FILL FILL_1__8436_ (
);

FILL FILL_1__8016_ (
);

FILL FILL_2__10341_ (
);

OR2X2 _7086_ (
    .A(_664_),
    .B(_669_),
    .Y(_671_)
);

FILL FILL_3__9303_ (
);

FILL FILL_2__6779_ (
);

FILL FILL_0__6761_ (
);

NAND2X1 _11084_ (
    .A(_4281_),
    .B(_4280_),
    .Y(_4282_)
);

FILL FILL_3__12973_ (
);

FILL FILL_2__7720_ (
);

FILL FILL_2__7300_ (
);

FILL FILL_3__12133_ (
);

FILL FILL_2__11966_ (
);

FILL FILL_2__11546_ (
);

FILL FILL_0__12580_ (
);

FILL FILL_2__11126_ (
);

FILL FILL_0__12160_ (
);

FILL FILL_1__10959_ (
);

FILL FILL_1__10539_ (
);

FILL FILL_1__10119_ (
);

FILL FILL_0__7966_ (
);

FILL FILL_0__7546_ (
);

NAND2X1 _9652_ (
    .A(_3004_),
    .B(_3001_),
    .Y(_3187_[13])
);

FILL FILL_0__7126_ (
);

OAI21X1 _9232_ (
    .A(_2590_),
    .B(_2591_),
    .C(_2589_),
    .Y(_2592_)
);

FILL FILL_1__11900_ (
);

OR2X2 _12289_ (
    .A(_5399_),
    .B(_5400_),
    .Y(_5401_)
);

FILL FILL_2__8925_ (
);

FILL FILL_2__8505_ (
);

NOR2X1 _13230_ (
    .A(_6252_),
    .B(_6253_),
    .Y(_6254_)
);

FILL FILL_1__6922_ (
);

FILL FILL_1__6502_ (
);

FILL FILL_3__6428_ (
);

FILL FILL_1__9394_ (
);

FILL FILL_1__10292_ (
);

FILL FILL_1__7707_ (
);

FILL FILL_3__13091_ (
);

OAI21X1 _6777_ (
    .A(_202_),
    .B(_292_),
    .C(_288_),
    .Y(_375_)
);

FILL FILL_2__12084_ (
);

FILL FILL_1__11497_ (
);

FILL FILL_1__11077_ (
);

INVX1 _10775_ (
    .A(_4766_),
    .Y(_4767_)
);

AOI21X1 _10355_ (
    .A(_3488_),
    .B(_3553_),
    .C(_3631_),
    .Y(_3632_)
);

FILL FILL_2__10817_ (
);

FILL FILL_2__9463_ (
);

FILL FILL_0__11851_ (
);

FILL FILL_2__9043_ (
);

FILL FILL_0__11431_ (
);

FILL FILL_0__11011_ (
);

FILL FILL_2__13289_ (
);

FILL FILL_0__6817_ (
);

NOR2X1 _8923_ (
    .A(_2345_),
    .B(_2346_),
    .Y(_2347_)
);

INVX1 _8503_ (
    .A(_1854_),
    .Y(_1941_)
);

FILL FILL_1__7880_ (
);

FILL FILL_1__7460_ (
);

FILL FILL_1__7040_ (
);

FILL FILL_0__9289_ (
);

FILL FILL_1__13223_ (
);

INVX1 _12921_ (
    .A(_5951_),
    .Y(_5958_)
);

FILL FILL_0__12636_ (
);

FILL FILL_0__12216_ (
);

DFFPOSX1 _12501_ (
    .D(_5573_[0]),
    .CLK(clk_bF$buf49),
    .Q(\u_fir_pe6.mul [0])
);

OR2X2 _9708_ (
    .A(_3052_),
    .B(_3050_),
    .Y(_3054_)
);

FILL FILL_1__8665_ (
);

FILL FILL_1__8245_ (
);

FILL FILL_2__10990_ (
);

FILL FILL_2__10570_ (
);

FILL FILL_2__10150_ (
);

FILL FILL_3__9952_ (
);

FILL FILL_3__9532_ (
);

FILL FILL_0__6990_ (
);

FILL FILL_0__6570_ (
);

FILL FILL_2__6588_ (
);

FILL FILL_3__12362_ (
);

FILL FILL_2__11775_ (
);

FILL FILL_2__11355_ (
);

FILL FILL_1__10768_ (
);

FILL FILL_1__10348_ (
);

FILL FILL_0__7775_ (
);

DFFPOSX1 _9881_ (
    .D(_3187_[11]),
    .CLK(clk_bF$buf4),
    .Q(\u_fir_pe3.mul [11])
);

FILL FILL_0__7355_ (
);

NAND2X1 _9461_ (
    .A(_2782_),
    .B(_2785_),
    .Y(_2818_)
);

NAND3X1 _9041_ (
    .A(_2401_),
    .B(_2403_),
    .C(_2402_),
    .Y(_2404_)
);

AOI21X1 _12098_ (
    .A(_5135_),
    .B(_5137_),
    .C(_5214_),
    .Y(_5215_)
);

FILL FILL_2__8734_ (
);

FILL FILL_2__8314_ (
);

FILL FILL_0__10702_ (
);

FILL FILL_3__13147_ (
);

FILL FILL_0__13174_ (
);

FILL FILL_1__6731_ (
);

FILL FILL_3__6657_ (
);

FILL FILL_1__12914_ (
);

FILL FILL_0__9921_ (
);

FILL FILL_2__9939_ (
);

FILL FILL_2__9519_ (
);

FILL FILL_0__9501_ (
);

FILL FILL_0__11907_ (
);

FILL FILL_1__7936_ (
);

FILL FILL_1__7516_ (
);

NAND3X1 _6586_ (
    .A(_172_),
    .B(_176_),
    .C(_179_),
    .Y(_186_)
);

FILL FILL_0__10299_ (
);

NAND2X1 _10584_ (
    .A(_3847_),
    .B(_3849_),
    .Y(_3850_)
);

NOR2X1 _10164_ (
    .A(_3429_),
    .B(_3442_),
    .Y(_3443_)
);

FILL FILL_2__6800_ (
);

FILL FILL_3__11213_ (
);

FILL FILL_2__9692_ (
);

FILL FILL_2__10626_ (
);

FILL FILL_2__9272_ (
);

FILL FILL_0__11660_ (
);

FILL FILL_2__10206_ (
);

FILL FILL_0__11240_ (
);

FILL FILL_2__13098_ (
);

FILL FILL_0__6626_ (
);

NAND3X1 _8732_ (
    .A(_2158_),
    .B(_2165_),
    .C(_2164_),
    .Y(_2166_)
);

AND2X2 _8312_ (
    .A(vdd),
    .B(\X[2] [4]),
    .Y(_1752_)
);

FILL FILL_0__9098_ (
);

INVX1 _11789_ (
    .A(_4902_),
    .Y(_4910_)
);

NAND3X1 _11369_ (
    .A(_4547_),
    .B(_4557_),
    .C(_4560_),
    .Y(_4563_)
);

FILL FILL_3__12838_ (
);

FILL FILL_1__13032_ (
);

FILL FILL253650x158550 (
);

FILL FILL_0__12865_ (
);

NAND3X1 _12730_ (
    .A(_5763_),
    .B(_5756_),
    .C(_5761_),
    .Y(_5770_)
);

FILL FILL_0__12445_ (
);

FILL FILL_0__12025_ (
);

NAND2X1 _12310_ (
    .A(_5413_),
    .B(_5418_),
    .Y(_5419_)
);

NAND2X1 _9937_ (
    .A(gnd),
    .B(\X[4] [1]),
    .Y(_3219_)
);

NAND3X1 _9517_ (
    .A(_2871_),
    .B(_2872_),
    .C(_2870_),
    .Y(_2873_)
);

FILL FILL_1__8894_ (
);

FILL FILL_1__8474_ (
);

FILL FILL_1__8054_ (
);

FILL FILL253950x18150 (
);

FILL FILL_3__9761_ (
);

FILL FILL_2__6397_ (
);

FILL FILL_1__9679_ (
);

FILL FILL_1__9259_ (
);

FILL FILL_3__12591_ (
);

FILL FILL_2__11164_ (
);

FILL FILL_1__10997_ (
);

FILL FILL_1__10577_ (
);

FILL FILL_1__10157_ (
);

FILL FILL_0__7584_ (
);

NAND2X1 _9690_ (
    .A(_3034_),
    .B(_3037_),
    .Y(_3181_[2])
);

FILL FILL_0__7164_ (
);

NAND2X1 _9270_ (
    .A(_2623_),
    .B(_2628_),
    .Y(_2629_)
);

FILL FILL_2__8543_ (
);

FILL FILL_0__10931_ (
);

FILL FILL_0__10511_ (
);

FILL FILL_2__12789_ (
);

FILL FILL_2__12369_ (
);

FILL FILL_1__6960_ (
);

FILL FILL_1__6540_ (
);

FILL FILL_0__8789_ (
);

FILL FILL_2__13310_ (
);

FILL FILL_3__6886_ (
);

FILL FILL_0__8369_ (
);

FILL FILL_1__12723_ (
);

FILL FILL_1__12303_ (
);

FILL FILL_0__9730_ (
);

FILL FILL_2__9748_ (
);

FILL FILL_0__9310_ (
);

FILL FILL_2__9328_ (
);

FILL FILL_0__11716_ (
);

FILL FILL_1__7745_ (
);

FILL FILL_1__7325_ (
);

NAND2X1 _6395_ (
    .A(gnd),
    .B(Xin[3]),
    .Y(_787_)
);

FILL FILL_3__8612_ (
);

AOI21X1 _10393_ (
    .A(gnd),
    .B(\X[4] [6]),
    .C(_3600_),
    .Y(_3669_)
);

FILL FILL_3__11862_ (
);

FILL FILL_3__11442_ (
);

FILL FILL_2__10855_ (
);

FILL FILL_2__10435_ (
);

FILL FILL_2__9081_ (
);

FILL FILL_2__10015_ (
);

FILL FILL_0__6855_ (
);

DFFPOSX1 _8961_ (
    .D(_2384_[8]),
    .CLK(clk_bF$buf0),
    .Q(\Y[3] [8])
);

FILL FILL_0__6435_ (
);

AOI21X1 _8541_ (
    .A(_1943_),
    .B(_1944_),
    .C(_1911_),
    .Y(_1978_)
);

DFFPOSX1 _8121_ (
    .D(_1593_[5]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.mul [5])
);

DFFPOSX1 _11598_ (
    .D(_4775_[14]),
    .CLK(clk_bF$buf6),
    .Q(\Y[6] [14])
);

AOI21X1 _11178_ (
    .A(\X[5] [3]),
    .B(gnd),
    .C(_4372_),
    .Y(_4375_)
);

FILL FILL_2__7814_ (
);

FILL FILL_3__12227_ (
);

FILL FILL_1__13261_ (
);

FILL FILL_0__12674_ (
);

FILL FILL_0__12254_ (
);

AND2X2 _9746_ (
    .A(_3068_),
    .B(_3078_),
    .Y(_3089_)
);

OAI21X1 _9326_ (
    .A(_2683_),
    .B(_2684_),
    .C(_2682_),
    .Y(_2685_)
);

FILL FILL_1__8283_ (
);

FILL FILL_3__9990_ (
);

FILL FILL_3__9150_ (
);

FILL FILL_0__13039_ (
);

NAND2X1 _13324_ (
    .A(_6343_),
    .B(_6337_),
    .Y(_6347_)
);

FILL FILL_1__9488_ (
);

FILL FILL_1__9068_ (
);

FILL FILL_2__11393_ (
);

FILL FILL_1__10386_ (
);

FILL FILL_0__7393_ (
);

FILL FILL_2__8772_ (
);

FILL FILL_2__8352_ (
);

FILL FILL_3__13185_ (
);

FILL FILL_0__10320_ (
);

FILL FILL_2__12598_ (
);

FILL FILL_2__12178_ (
);

INVX1 _7812_ (
    .A(_1326_),
    .Y(_1327_)
);

FILL FILL_0__8598_ (
);

FILL FILL_0__8178_ (
);

NAND2X1 _10869_ (
    .A(gnd),
    .B(\X[5] [4]),
    .Y(_4070_)
);

AND2X2 _10449_ (
    .A(_3723_),
    .B(_3720_),
    .Y(_3724_)
);

NAND3X1 _10029_ (
    .A(_3309_),
    .B(_3242_),
    .C(_3245_),
    .Y(_3310_)
);

FILL FILL_1__12952_ (
);

FILL FILL_1__12532_ (
);

FILL FILL_1__12112_ (
);

FILL FILL_2__9977_ (
);

FILL FILL_2__9557_ (
);

FILL FILL_0__11945_ (
);

FILL FILL_2__9137_ (
);

NAND3X1 _11810_ (
    .A(gnd),
    .B(\X[7] [6]),
    .C(_4927_),
    .Y(_4930_)
);

FILL FILL_0__11525_ (
);

FILL FILL_0__11105_ (
);

FILL FILL_1__7974_ (
);

FILL FILL_1__7554_ (
);

FILL FILL_1__7134_ (
);

FILL FILL_1__13317_ (
);

FILL FILL_3__8841_ (
);

FILL FILL_3__8421_ (
);

FILL FILL_3__8001_ (
);

FILL FILL_1__8759_ (
);

FILL FILL_1__8339_ (
);

FILL FILL_2__10664_ (
);

FILL FILL_2__10244_ (
);

FILL FILL_1__9700_ (
);

FILL FILL_3__9626_ (
);

FILL FILL_0__6664_ (
);

NAND2X1 _8770_ (
    .A(_2199_),
    .B(_2202_),
    .Y(_2203_)
);

NAND3X1 _8350_ (
    .A(_1784_),
    .B(_1785_),
    .C(_1786_),
    .Y(_1790_)
);

FILL FILL_2__7623_ (
);

FILL FILL_3__12456_ (
);

FILL FILL_1__13070_ (
);

FILL FILL_2__11869_ (
);

FILL FILL_2__11449_ (
);

FILL FILL_2__11029_ (
);

FILL FILL_0__12063_ (
);

FILL FILL_2__12810_ (
);

FILL FILL_0__7869_ (
);

NOR3X1 _9975_ (
    .A(_3241_),
    .B(_3208_),
    .C(_3253_),
    .Y(_3256_)
);

FILL FILL_0__7449_ (
);

OAI22X1 _9555_ (
    .A(_2808_),
    .B(_2853_),
    .C(_2909_),
    .D(_2908_),
    .Y(_2910_)
);

FILL FILL_0__7029_ (
);

NAND3X1 _9135_ (
    .A(_2493_),
    .B(_2495_),
    .C(_2494_),
    .Y(_2496_)
);

FILL FILL_1__11803_ (
);

FILL FILL_0__8810_ (
);

FILL FILL_2__8828_ (
);

FILL FILL_2__8408_ (
);

FILL FILL_0__13268_ (
);

OAI21X1 _13133_ (
    .A(_5955_),
    .B(_6166_),
    .C(_6138_),
    .Y(_6167_)
);

FILL FILL_1__6825_ (
);

FILL FILL_1__6405_ (
);

FILL FILL_1__9297_ (
);

FILL FILL254250x86550 (
);

FILL FILL_1__10195_ (
);

FILL FILL_3__10942_ (
);

FILL FILL_3__10102_ (
);

FILL FILL_2__8581_ (
);

FILL FILL_2__8161_ (
);

INVX1 _7621_ (
    .A(_1119_),
    .Y(_1139_)
);

DFFPOSX1 _7201_ (
    .D(_790_[2]),
    .CLK(clk_bF$buf52),
    .Q(\Y[1] [2])
);

NOR2X1 _10678_ (
    .A(\u_fir_pe4.rYin [13]),
    .B(\u_fir_pe4.mul [13]),
    .Y(_3942_)
);

AOI21X1 _10258_ (
    .A(_3447_),
    .B(_3449_),
    .C(_3535_),
    .Y(_3536_)
);

FILL FILL_3__11727_ (
);

FILL FILL_1__12761_ (
);

FILL FILL_3__11307_ (
);

FILL FILL_1__12341_ (
);

FILL FILL_2__9786_ (
);

FILL FILL_2__9366_ (
);

FILL FILL_0__11754_ (
);

FILL FILL_0__11334_ (
);

NOR2X1 _8826_ (
    .A(\u_fir_pe2.rYin [4]),
    .B(\u_fir_pe2.mul [4]),
    .Y(_2252_)
);

OAI21X1 _8406_ (
    .A(_1844_),
    .B(_1839_),
    .C(_1833_),
    .Y(_1845_)
);

FILL FILL_1__7783_ (
);

FILL FILL_1__7363_ (
);

FILL FILL_3__7289_ (
);

FILL FILL_1__13126_ (
);

FILL FILL_0__12959_ (
);

AOI21X1 _12824_ (
    .A(_5862_),
    .B(_5861_),
    .C(_5860_),
    .Y(_5863_)
);

FILL FILL_3__8230_ (
);

FILL FILL_0__12539_ (
);

NOR2X1 _12404_ (
    .A(_5506_),
    .B(_5507_),
    .Y(_5508_)
);

FILL FILL_0__12119_ (
);

FILL FILL254550x230550 (
);

FILL FILL_1__8568_ (
);

FILL FILL_1__8148_ (
);

FILL FILL_3__11060_ (
);

FILL FILL_2__10893_ (
);

FILL FILL_2__10473_ (
);

FILL FILL_2__10053_ (
);

FILL FILL_3__9015_ (
);

FILL FILL_0__6893_ (
);

FILL FILL_0__6473_ (
);

FILL FILL_2__7852_ (
);

FILL FILL_3__12685_ (
);

FILL FILL_2__7432_ (
);

FILL FILL_2__7012_ (
);

FILL FILL_2__11678_ (
);

FILL FILL_2__11258_ (
);

FILL FILL_0__12292_ (
);

FILL FILL_0__7678_ (
);

AND2X2 _9784_ (
    .A(_3123_),
    .B(_3126_),
    .Y(_3128_)
);

FILL FILL_0__7258_ (
);

AND2X2 _9364_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2722_)
);

FILL FILL_2__8637_ (
);

FILL FILL_2__8217_ (
);

FILL FILL_0__10605_ (
);

FILL FILL_0__13077_ (
);

DFFPOSX1 _13362_ (
    .D(\Y[6] [0]),
    .CLK(clk_bF$buf40),
    .Q(\u_fir_pe7.rYin [0])
);

FILL FILL_1__6634_ (
);

FILL FILL_2__13404_ (
);

FILL FILL_1__12817_ (
);

FILL FILL_0__9824_ (
);

FILL FILL_0__9404_ (
);

FILL FILL_3__7501_ (
);

FILL FILL_1__7839_ (
);

FILL FILL_1__7419_ (
);

FILL FILL_3__10331_ (
);

FILL FILL_2__8390_ (
);

OAI21X1 _6489_ (
    .A(_89_),
    .B(_15_),
    .C(_83_),
    .Y(_90_)
);

NOR2X1 _7850_ (
    .A(_941_),
    .B(_1102_),
    .Y(_1364_)
);

NAND2X1 _7430_ (
    .A(vdd),
    .B(\X[1] [3]),
    .Y(_950_)
);

OR2X2 _7010_ (
    .A(_601_),
    .B(_594_),
    .Y(_603_)
);

NOR2X1 _10487_ (
    .A(_3753_),
    .B(_3757_),
    .Y(_3761_)
);

NAND2X1 _10067_ (
    .A(_3275_),
    .B(_3346_),
    .Y(_3347_)
);

FILL FILL_3__11956_ (
);

FILL FILL_2__6703_ (
);

FILL FILL_1__12990_ (
);

FILL FILL_3__11536_ (
);

FILL FILL_1__12570_ (
);

FILL FILL_1__12150_ (
);

FILL FILL_2__10949_ (
);

FILL FILL_2__9595_ (
);

FILL FILL_0__11983_ (
);

FILL FILL_2__10529_ (
);

FILL FILL_2__9175_ (
);

FILL FILL_0__11563_ (
);

FILL FILL_2__10109_ (
);

FILL FILL_0__11143_ (
);

FILL FILL_0__6949_ (
);

FILL FILL_0__6529_ (
);

AND2X2 _8635_ (
    .A(vdd),
    .B(\X[2] [6]),
    .Y(_2071_)
);

AOI21X1 _8215_ (
    .A(_1634_),
    .B(_1638_),
    .C(_1626_),
    .Y(_1657_)
);

FILL FILL_1__7592_ (
);

FILL FILL_1__7172_ (
);

FILL FILL_3__7098_ (
);

FILL FILL_2__7908_ (
);

FILL FILL_0__12768_ (
);

NAND3X1 _12633_ (
    .A(_5664_),
    .B(_5671_),
    .C(_5673_),
    .Y(_5674_)
);

FILL FILL_0__12348_ (
);

NAND3X1 _12213_ (
    .A(_5325_),
    .B(_5327_),
    .C(_5326_),
    .Y(_5328_)
);

FILL FILL_1__8797_ (
);

FILL FILL_1__8377_ (
);

FILL FILL_2__10282_ (
);

FILL FILL_3__9244_ (
);

FILL FILL_2__7661_ (
);

FILL FILL_3__12074_ (
);

FILL FILL_2__11487_ (
);

FILL FILL_2__11067_ (
);

AOI21X1 _6701_ (
    .A(_281_),
    .B(_283_),
    .C(_298_),
    .Y(_299_)
);

FILL FILL_0__7487_ (
);

NOR3X1 _9593_ (
    .A(_2893_),
    .B(_2895_),
    .C(_2943_),
    .Y(_2947_)
);

FILL FILL_0__7067_ (
);

AND2X2 _9173_ (
    .A(gnd),
    .B(\X[3] [6]),
    .Y(_2533_)
);

FILL FILL_3__10807_ (
);

FILL FILL_1__11841_ (
);

FILL FILL_1__11421_ (
);

FILL FILL_1__11001_ (
);

FILL FILL_2__8866_ (
);

FILL FILL_2__8446_ (
);

FILL FILL_0__10834_ (
);

FILL FILL_3__13279_ (
);

FILL FILL_0__10414_ (
);

FILL FILL_2__8026_ (
);

NOR3X1 _13171_ (
    .A(_6202_),
    .B(_6170_),
    .C(_6188_),
    .Y(_6203_)
);

NAND2X1 _7906_ (
    .A(_1417_),
    .B(_1416_),
    .Y(_1418_)
);

FILL FILL_1__6863_ (
);

FILL FILL_1__6443_ (
);

FILL FILL_2__13213_ (
);

FILL FILL_1__12626_ (
);

FILL FILL_1__12206_ (
);

FILL FILL_0__9633_ (
);

FILL FILL_3__7730_ (
);

FILL FILL_0__9213_ (
);

NAND2X1 _11904_ (
    .A(gnd),
    .B(\X[7] [4]),
    .Y(_5023_)
);

FILL FILL_1__7648_ (
);

FILL FILL_3__8935_ (
);

FILL FILL_3__8515_ (
);

OAI21X1 _10296_ (
    .A(_3503_),
    .B(_3572_),
    .C(_3542_),
    .Y(_3573_)
);

FILL FILL_2__6932_ (
);

FILL FILL_2__6512_ (
);

FILL FILL_0__11792_ (
);

FILL FILL_2__10338_ (
);

FILL FILL_0__11372_ (
);

FILL FILL_0__6758_ (
);

NOR2X1 _8864_ (
    .A(\u_fir_pe2.rYin [8]),
    .B(\u_fir_pe2.mul [8]),
    .Y(_2287_)
);

AND2X2 _8444_ (
    .A(_1879_),
    .B(_1882_),
    .Y(_1883_)
);

AND2X2 _8024_ (
    .A(_1526_),
    .B(_1527_),
    .Y(_1587_[10])
);

FILL FILL_2__7717_ (
);

FILL FILL_1__13164_ (
);

FILL FILL_0__12997_ (
);

NAND2X1 _12862_ (
    .A(\X[6] [4]),
    .B(gnd),
    .Y(_5900_)
);

FILL FILL_0__12577_ (
);

FILL FILL_0__12157_ (
);

NOR2X1 _12442_ (
    .A(_5545_),
    .B(_5544_),
    .Y(_5546_)
);

INVX1 _12022_ (
    .A(_5053_),
    .Y(_5140_)
);

FILL FILL_2__12904_ (
);

NAND2X1 _9649_ (
    .A(_2980_),
    .B(_2979_),
    .Y(_3002_)
);

AOI21X1 _9229_ (
    .A(_2417_),
    .B(_2501_),
    .C(_2588_),
    .Y(_2589_)
);

FILL FILL_1__8186_ (
);

FILL FILL_0__8904_ (
);

FILL FILL_2__10091_ (
);

FILL FILL_3__9473_ (
);

OAI21X1 _13227_ (
    .A(_6244_),
    .B(_6245_),
    .C(_6249_),
    .Y(_6251_)
);

FILL FILL_1__6919_ (
);

FILL FILL_2__7890_ (
);

FILL FILL_2__7470_ (
);

FILL FILL_2__7050_ (
);

FILL FILL_2__11296_ (
);

NAND2X1 _6930_ (
    .A(_331_),
    .B(_405_),
    .Y(_525_)
);

NAND3X1 _6510_ (
    .A(_26_),
    .B(_106_),
    .C(_110_),
    .Y(_111_)
);

FILL FILL_1__10289_ (
);

FILL FILL_0__7296_ (
);

FILL FILL_1__11650_ (
);

FILL FILL_1__11230_ (
);

FILL FILL_2__8675_ (
);

FILL FILL_2__8255_ (
);

FILL FILL_0__10643_ (
);

FILL FILL_0__10223_ (
);

AOI21X1 _7715_ (
    .A(_1222_),
    .B(_1220_),
    .C(_1192_),
    .Y(_1232_)
);

FILL FILL_1__6672_ (
);

FILL FILL_2__13022_ (
);

FILL FILL_3__6598_ (
);

FILL FILL_1__12855_ (
);

FILL FILL_1__12435_ (
);

FILL FILL_1__12015_ (
);

FILL FILL_0__9442_ (
);

FILL FILL_0__11848_ (
);

FILL FILL_0__9022_ (
);

AOI22X1 _11713_ (
    .A(_4791_),
    .B(_4796_),
    .C(_4831_),
    .D(_4834_),
    .Y(_4835_)
);

FILL FILL_0__11428_ (
);

FILL FILL_0__11008_ (
);

FILL FILL_1__7877_ (
);

FILL FILL_1__7457_ (
);

FILL FILL_1__7037_ (
);

AND2X2 _12918_ (
    .A(_5946_),
    .B(_5951_),
    .Y(_5956_)
);

FILL FILL_3__11994_ (
);

FILL FILL_2__6741_ (
);

FILL FILL_3__11154_ (
);

FILL FILL_2__10987_ (
);

FILL FILL_2__10567_ (
);

FILL FILL_2__10147_ (
);

FILL FILL_0__11181_ (
);

FILL FILL_1__9603_ (
);

FILL FILL_3__9109_ (
);

FILL FILL_0__6987_ (
);

FILL FILL_0__6567_ (
);

AOI21X1 _8673_ (
    .A(_2054_),
    .B(_2088_),
    .C(_2107_),
    .Y(_2108_)
);

OAI21X1 _8253_ (
    .A(_1692_),
    .B(_1693_),
    .C(_1691_),
    .Y(_1694_)
);

FILL FILL_1__10921_ (
);

FILL FILL_1__10501_ (
);

FILL FILL_2__7946_ (
);

FILL FILL_3__12779_ (
);

FILL FILL_2__7526_ (
);

FILL FILL_2__7106_ (
);

NAND2X1 _12671_ (
    .A(gnd),
    .B(\X[6]_5_bF$buf2 ),
    .Y(_5711_)
);

FILL FILL_0__12386_ (
);

OR2X2 _12251_ (
    .A(_5363_),
    .B(_5361_),
    .Y(_5365_)
);

FILL FILL_3__13300_ (
);

FILL FILL_2__12713_ (
);

DFFPOSX1 _9878_ (
    .D(_3187_[8]),
    .CLK(clk_bF$buf4),
    .Q(\u_fir_pe3.mul [8])
);

NAND2X1 _9458_ (
    .A(_2806_),
    .B(_2813_),
    .Y(_2815_)
);

INVX1 _9038_ (
    .A(_3131_),
    .Y(_2401_)
);

FILL FILL_1__11706_ (
);

FILL FILL_0__8713_ (
);

FILL FILL_3__6810_ (
);

NAND2X1 _13036_ (
    .A(_6070_),
    .B(_6066_),
    .Y(_6072_)
);

FILL FILL_1__6728_ (
);

FILL FILL_0__9918_ (
);

FILL FILL_1__10098_ (
);

FILL FILL_3__10425_ (
);

FILL FILL_2__8484_ (
);

FILL FILL_0__10872_ (
);

FILL FILL_0__10452_ (
);

FILL FILL_2__8064_ (
);

FILL FILL_0__10032_ (
);

OR2X2 _7944_ (
    .A(_1444_),
    .B(_1449_),
    .Y(_1451_)
);

INVX1 _7524_ (
    .A(_1037_),
    .Y(_1043_)
);

NOR2X1 _7104_ (
    .A(_684_),
    .B(_683_),
    .Y(_687_)
);

FILL FILL_1__6481_ (
);

FILL FILL_2__13251_ (
);

FILL FILL_1__12664_ (
);

FILL FILL_1__12244_ (
);

FILL FILL_0__9671_ (
);

FILL FILL_2__9689_ (
);

FILL FILL_0__9251_ (
);

FILL FILL_2__9269_ (
);

NAND3X1 _11942_ (
    .A(_5059_),
    .B(_5060_),
    .C(_5058_),
    .Y(_5061_)
);

FILL FILL_0__11657_ (
);

INVX1 _11522_ (
    .A(_4704_),
    .Y(_4706_)
);

FILL FILL_0__11237_ (
);

NAND2X1 _11102_ (
    .A(_4295_),
    .B(_4299_),
    .Y(_4300_)
);

AOI21X1 _8729_ (
    .A(gnd),
    .B(_2160_),
    .C(_2162_),
    .Y(_2163_)
);

OAI22X1 _8309_ (
    .A(_1636_),
    .B(_1747_),
    .C(_1679_),
    .D(_1748_),
    .Y(_1749_)
);

FILL FILL_1__7686_ (
);

FILL FILL_1__7266_ (
);

FILL FILL_1__13029_ (
);

FILL FILL_3__8553_ (
);

AOI22X1 _12727_ (
    .A(_5690_),
    .B(_5685_),
    .C(_5762_),
    .D(_5766_),
    .Y(_5767_)
);

FILL FILL_3__8133_ (
);

NOR2X1 _12307_ (
    .A(_5414_),
    .B(_5415_),
    .Y(_5416_)
);

FILL FILL_2__6970_ (
);

FILL FILL_2__6550_ (
);

FILL FILL_3__11383_ (
);

FILL FILL_2__10796_ (
);

FILL FILL_2__10376_ (
);

FILL FILL_1__9412_ (
);

FILL FILL_3__9338_ (
);

FILL FILL_0__6796_ (
);

NAND3X1 _8482_ (
    .A(gnd),
    .B(\X[2] [6]),
    .C(_1919_),
    .Y(_1920_)
);

NAND2X1 _8062_ (
    .A(_1561_),
    .B(_1555_),
    .Y(_1565_)
);

FILL FILL_1__10310_ (
);

FILL FILL_2__7755_ (
);

FILL FILL_2__7335_ (
);

FILL FILL_3__12168_ (
);

FILL FILL_0__12195_ (
);

DFFPOSX1 _12480_ (
    .D(\X[7] [3]),
    .CLK(clk_bF$buf29),
    .Q(_6376_[3])
);

AND2X2 _12060_ (
    .A(_5176_),
    .B(_5173_),
    .Y(_5177_)
);

FILL FILL_2__12942_ (
);

FILL FILL_2__12522_ (
);

FILL FILL_2__12102_ (
);

INVX1 _9687_ (
    .A(_3031_),
    .Y(_3035_)
);

INVX1 _9267_ (
    .A(\X[3] [7]),
    .Y(_2626_)
);

FILL FILL_1__11935_ (
);

FILL FILL_1__11515_ (
);

FILL FILL_0__8942_ (
);

FILL FILL_0__8522_ (
);

FILL FILL_0__10928_ (
);

FILL FILL_0__10508_ (
);

FILL FILL_3__9091_ (
);

INVX1 _13265_ (
    .A(_6284_),
    .Y(_6288_)
);

FILL FILL_2__9901_ (
);

FILL FILL_1__6957_ (
);

FILL FILL_1__6537_ (
);

FILL FILL_2__13307_ (
);

FILL FILL_0__9727_ (
);

FILL FILL_3__7824_ (
);

FILL FILL_0__9307_ (
);

FILL FILL_3__10654_ (
);

FILL FILL_2__8293_ (
);

FILL FILL_0__10681_ (
);

FILL FILL_0__10261_ (
);

FILL FILL254250x18150 (
);

FILL FILL_3__8609_ (
);

OAI21X1 _7753_ (
    .A(_1216_),
    .B(_1268_),
    .C(_1204_),
    .Y(_1269_)
);

NAND2X1 _7333_ (
    .A(_851_),
    .B(_854_),
    .Y(_855_)
);

FILL FILL_2__13060_ (
);

FILL FILL_2__6606_ (
);

FILL FILL_1__12893_ (
);

FILL FILL_1__12053_ (
);

FILL FILL_0__9480_ (
);

FILL FILL_2__9498_ (
);

FILL FILL_0__11886_ (
);

FILL FILL_0__9060_ (
);

FILL FILL_2__9078_ (
);

OAI21X1 _11751_ (
    .A(_4871_),
    .B(_4797_),
    .C(_4865_),
    .Y(_4872_)
);

FILL FILL_0__11466_ (
);

FILL FILL_0__11046_ (
);

NAND2X1 _11331_ (
    .A(_4525_),
    .B(_4524_),
    .Y(_4526_)
);

FILL FILL_3__12800_ (
);

DFFPOSX1 _8958_ (
    .D(_2384_[5]),
    .CLK(clk_bF$buf47),
    .Q(\Y[3] [5])
);

AOI21X1 _8538_ (
    .A(_1955_),
    .B(_1954_),
    .C(_1897_),
    .Y(_1975_)
);

DFFPOSX1 _8118_ (
    .D(_1590_[2]),
    .CLK(clk_bF$buf19),
    .Q(\u_fir_pe1.mul [2])
);

FILL FILL_1__7495_ (
);

FILL FILL_1__7075_ (
);

FILL FILL_1__13258_ (
);

FILL FILL_3__8782_ (
);

NAND2X1 _12956_ (
    .A(_5992_),
    .B(_5988_),
    .Y(_5993_)
);

NAND2X1 _12536_ (
    .A(gnd),
    .B(\X[6] [2]),
    .Y(_5579_)
);

OR2X2 _12116_ (
    .A(_5162_),
    .B(_5232_),
    .Y(_5233_)
);

FILL FILL_2__10185_ (
);

FILL FILL_1__9641_ (
);

FILL FILL_1__9221_ (
);

FILL FILL_3__9987_ (
);

FILL FILL_3__9567_ (
);

AOI21X1 _8291_ (
    .A(_1685_),
    .B(_1689_),
    .C(_1678_),
    .Y(_1731_)
);

FILL FILL_1_CLKBUF1_insert90 (
);

FILL FILL_1_CLKBUF1_insert91 (
);

FILL FILL_1_CLKBUF1_insert92 (
);

FILL FILL_1_CLKBUF1_insert93 (
);

FILL FILL_1_CLKBUF1_insert94 (
);

FILL FILL_2__7984_ (
);

FILL FILL_1_CLKBUF1_insert95 (
);

FILL FILL_2__7564_ (
);

FILL FILL_3__12397_ (
);

FILL FILL_1_CLKBUF1_insert96 (
);

FILL FILL_2__7144_ (
);

AOI21X1 _6604_ (
    .A(_120_),
    .B(_126_),
    .C(_203_),
    .Y(_204_)
);

FILL FILL_2__12751_ (
);

FILL FILL_2__12331_ (
);

OAI21X1 _9496_ (
    .A(_2818_),
    .B(_2820_),
    .C(_2814_),
    .Y(_2852_)
);

NAND2X1 _9076_ (
    .A(_2435_),
    .B(_2431_),
    .Y(_2438_)
);

FILL FILL_1__11744_ (
);

FILL FILL_1__11324_ (
);

FILL FILL_2__8769_ (
);

FILL FILL_0__8751_ (
);

FILL FILL_0__8331_ (
);

FILL FILL_2__8349_ (
);

FILL FILL_0__10317_ (
);

NAND2X1 _10602_ (
    .A(_3865_),
    .B(_3860_),
    .Y(_3866_)
);

INVX1 _13074_ (
    .A(_6108_),
    .Y(_6109_)
);

FILL FILL_2__9710_ (
);

OAI22X1 _7809_ (
    .A(_1030_),
    .B(_1032_),
    .C(_1116_),
    .D(_941_),
    .Y(_1324_)
);

FILL FILL_1__6766_ (
);

FILL FILL_2__13116_ (
);

FILL FILL_1__12949_ (
);

FILL FILL_1__12529_ (
);

FILL FILL_1__12109_ (
);

FILL FILL_0__9956_ (
);

FILL FILL_0__9536_ (
);

FILL FILL_0__9116_ (
);

NAND2X1 _11807_ (
    .A(\X[7] [2]),
    .B(gnd),
    .Y(_4927_)
);

FILL FILL_3__10883_ (
);

FILL FILL_3__10463_ (
);

FILL FILL_3__10043_ (
);

FILL FILL_0__10490_ (
);

FILL FILL_0__10070_ (
);

FILL FILL_1__8912_ (
);

FILL FILL_3__8838_ (
);

NAND2X1 _7982_ (
    .A(_1484_),
    .B(_1483_),
    .Y(_1485_)
);

AOI21X1 _7562_ (
    .A(_1080_),
    .B(_1079_),
    .C(_1078_),
    .Y(_1081_)
);

NOR2X1 _7142_ (
    .A(_724_),
    .B(_725_),
    .Y(_726_)
);

OAI21X1 _10199_ (
    .A(_3395_),
    .B(_3392_),
    .C(_3477_),
    .Y(_3478_)
);

FILL FILL_2__6835_ (
);

FILL FILL_3__11668_ (
);

FILL FILL_2__6415_ (
);

FILL FILL_3__11248_ (
);

FILL FILL_1__12282_ (
);

AOI21X1 _11980_ (
    .A(_5038_),
    .B(_5035_),
    .C(_5021_),
    .Y(_5098_)
);

FILL FILL_0__11695_ (
);

OAI21X1 _11560_ (
    .A(_4736_),
    .B(_4737_),
    .C(_4741_),
    .Y(_4743_)
);

FILL FILL_0__11275_ (
);

AND2X2 _11140_ (
    .A(_4299_),
    .B(_4295_),
    .Y(_4338_)
);

OAI21X1 _8767_ (
    .A(_2157_),
    .B(_2170_),
    .C(_2174_),
    .Y(_2200_)
);

AOI21X1 _8347_ (
    .A(_1786_),
    .B(_1785_),
    .C(_1784_),
    .Y(_1787_)
);

FILL FILL_0__7602_ (
);

FILL FILL_1__13067_ (
);

NAND2X1 _12765_ (
    .A(\X[6] [2]),
    .B(gnd),
    .Y(_5804_)
);

FILL FILL_3__8171_ (
);

NOR2X1 _12345_ (
    .A(\u_fir_pe6.rYin [5]),
    .B(\u_fir_pe6.mul [5]),
    .Y(_5450_)
);

FILL FILL_2__12807_ (
);

FILL FILL_0__13001_ (
);

FILL FILL_0__8807_ (
);

FILL FILL_3__6904_ (
);

FILL FILL_1__9450_ (
);

FILL FILL_1__9030_ (
);

FILL FILL_3__9796_ (
);

FILL FILL_2__7793_ (
);

FILL FILL_2__7373_ (
);

FILL FILL_2__11199_ (
);

OAI21X1 _6833_ (
    .A(_429_),
    .B(_428_),
    .C(_427_),
    .Y(_430_)
);

NAND2X1 _6413_ (
    .A(_13_),
    .B(_9_),
    .Y(_16_)
);

FILL FILL_2__12980_ (
);

FILL FILL_2__12560_ (
);

FILL FILL_2__12140_ (
);

FILL FILL_1__11973_ (
);

FILL FILL_3__10519_ (
);

FILL FILL_1__11553_ (
);

FILL FILL_1__11133_ (
);

FILL FILL_2__8578_ (
);

FILL FILL_0__8560_ (
);

FILL FILL_0__10966_ (
);

FILL FILL_0__8140_ (
);

FILL FILL_2__8158_ (
);

FILL FILL_0__10546_ (
);

NAND2X1 _10831_ (
    .A(_4031_),
    .B(_4032_),
    .Y(_4033_)
);

AND2X2 _10411_ (
    .A(_3675_),
    .B(_3679_),
    .Y(_3687_)
);

FILL FILL_0__10126_ (
);

NAND3X1 _7618_ (
    .A(_1121_),
    .B(_1123_),
    .C(_1125_),
    .Y(_1136_)
);

FILL FILL_1__6995_ (
);

FILL FILL_1__6575_ (
);

FILL FILL_1__12758_ (
);

FILL FILL_1__12338_ (
);

FILL FILL_0__9765_ (
);

FILL FILL_0__9345_ (
);

FILL FILL_3__7442_ (
);

DFFPOSX1 _11616_ (
    .D(\Y[5] [8]),
    .CLK(clk_bF$buf30),
    .Q(\u_fir_pe5.rYin [8])
);

FILL FILL_3__7022_ (
);

FILL FILL_3__10692_ (
);

FILL FILL_3__10272_ (
);

FILL FILL_1__8721_ (
);

FILL FILL_1__8301_ (
);

FILL FILL_3__8647_ (
);

FILL FILL_3__8227_ (
);

NOR2X1 _7791_ (
    .A(_1302_),
    .B(_1306_),
    .Y(_1307_)
);

NAND3X1 _7371_ (
    .A(_882_),
    .B(_889_),
    .C(_891_),
    .Y(_892_)
);

FILL FILL_3__11897_ (
);

FILL FILL_2__6644_ (
);

FILL FILL_3__11477_ (
);

FILL FILL_1__12091_ (
);

FILL FILL_0__11084_ (
);

FILL FILL_1__9926_ (
);

FILL FILL_1__9506_ (
);

FILL FILL_2__11831_ (
);

FILL FILL_2__11411_ (
);

DFFPOSX1 _8996_ (
    .D(_2388_[3]),
    .CLK(clk_bF$buf0),
    .Q(\u_fir_pe2.mul [3])
);

OAI21X1 _8576_ (
    .A(_1619_),
    .B(_2010_),
    .C(_2012_),
    .Y(_2013_)
);

INVX1 _8156_ (
    .A(_1598_),
    .Y(_1599_)
);

FILL FILL_1__10824_ (
);

FILL FILL_1__10404_ (
);

FILL FILL_2__7849_ (
);

FILL FILL_0__7831_ (
);

FILL FILL_0__7411_ (
);

FILL FILL_2__7429_ (
);

FILL FILL_2__7009_ (
);

FILL FILL_1__13296_ (
);

NAND2X1 _12994_ (
    .A(_6029_),
    .B(_5959_),
    .Y(_6031_)
);

FILL FILL_0__12289_ (
);

NAND2X1 _12574_ (
    .A(_5614_),
    .B(_5615_),
    .Y(_5616_)
);

NAND2X1 _12154_ (
    .A(_5251_),
    .B(_5248_),
    .Y(_5270_)
);

FILL FILL_2__12616_ (
);

FILL FILL_0__13230_ (
);

FILL FILL_0__8616_ (
);

FILL FILL_3__9185_ (
);

DFFPOSX1 _13359_ (
    .D(\X[6]_5_bF$buf3 ),
    .CLK(clk_bF$buf37),
    .Q(\X[7] [5])
);

FILL FILL_2__7182_ (
);

FILL FILL_3__7918_ (
);

NAND2X1 _6642_ (
    .A(gnd),
    .B(Xin[4]),
    .Y(_241_)
);

FILL FILL_1__11782_ (
);

FILL FILL_1__11362_ (
);

FILL FILL_2__8387_ (
);

FILL FILL_0__10775_ (
);

OR2X2 _10640_ (
    .A(_3899_),
    .B(_3903_),
    .Y(_3904_)
);

FILL FILL_0__10355_ (
);

OAI21X1 _10220_ (
    .A(_3496_),
    .B(_3497_),
    .C(_3492_),
    .Y(_3498_)
);

INVX1 _7847_ (
    .A(_1323_),
    .Y(_1361_)
);

NAND2X1 _7427_ (
    .A(_946_),
    .B(_938_),
    .Y(_947_)
);

OR2X2 _7007_ (
    .A(_572_),
    .B(_598_),
    .Y(_600_)
);

FILL FILL_1__6384_ (
);

FILL FILL_2__13154_ (
);

FILL FILL_1__12987_ (
);

FILL FILL_1__12567_ (
);

FILL FILL_1__12147_ (
);

FILL FILL_0__9994_ (
);

FILL FILL_0__9574_ (
);

FILL FILL_3__7671_ (
);

FILL FILL_0__9154_ (
);

NAND3X1 _11845_ (
    .A(_4918_),
    .B(_4959_),
    .C(_4964_),
    .Y(_4965_)
);

NAND2X1 _11425_ (
    .A(_4615_),
    .B(_4614_),
    .Y(_4781_[15])
);

AOI21X1 _11005_ (
    .A(_4132_),
    .B(_4128_),
    .C(_4197_),
    .Y(_4204_)
);

FILL FILL_0__12921_ (
);

FILL FILL_1__7589_ (
);

FILL FILL_1__7169_ (
);

FILL FILL_3__10081_ (
);

FILL FILL_1__8950_ (
);

FILL FILL_1__8530_ (
);

FILL FILL_3__8876_ (
);

FILL FILL_3__8456_ (
);

FILL FILL_3__8036_ (
);

NOR2X1 _7180_ (
    .A(_763_),
    .B(_762_),
    .Y(_764_)
);

FILL FILL_2__6873_ (
);

FILL FILL_2__6453_ (
);

FILL FILL_2__10699_ (
);

FILL FILL_2__10279_ (
);

FILL FILL_1__9735_ (
);

FILL FILL_1__9315_ (
);

FILL FILL_2__11640_ (
);

FILL FILL_2__11220_ (
);

FILL FILL_0__6699_ (
);

AOI22X1 _8385_ (
    .A(vdd),
    .B(\X[2] [7]),
    .C(\X[2] [3]),
    .D(vdd),
    .Y(_1824_)
);

FILL FILL_1__10633_ (
);

FILL FILL_1__10213_ (
);

FILL FILL_2__7658_ (
);

FILL FILL_0__7640_ (
);

FILL FILL_0__12098_ (
);

NOR2X1 _12383_ (
    .A(_5475_),
    .B(_5474_),
    .Y(_5487_)
);

FILL FILL_3__13012_ (
);

FILL FILL_2__12845_ (
);

FILL FILL_2__12425_ (
);

FILL FILL_2__12005_ (
);

FILL FILL_1__11838_ (
);

FILL FILL_1__11418_ (
);

FILL FILL_0__8845_ (
);

FILL FILL_0__8425_ (
);

FILL FILL_3__6522_ (
);

FILL FILL_0__8005_ (
);

NAND2X1 _13168_ (
    .A(_6199_),
    .B(_6198_),
    .Y(_6200_)
);

FILL FILL_2__9804_ (
);

FILL FILL_1__7801_ (
);

FILL FILL_3__7307_ (
);

NOR2X1 _6871_ (
    .A(_15_),
    .B(_462_),
    .Y(_467_)
);

AOI22X1 _6451_ (
    .A(_9_),
    .B(_14_),
    .C(_49_),
    .D(_52_),
    .Y(_53_)
);

FILL FILL_3__10977_ (
);

FILL FILL_3__10137_ (
);

FILL FILL_1__11171_ (
);

FILL FILL_2__8196_ (
);

FILL FILL_0__10584_ (
);

FILL FILL_0__10164_ (
);

FILL FILL_2__10911_ (
);

AND2X2 _7656_ (
    .A(_1164_),
    .B(_1169_),
    .Y(_1174_)
);

DFFPOSX1 _7236_ (
    .D(Yin[13]),
    .CLK(clk_bF$buf33),
    .Q(\u_fir_pe0.rYin [13])
);

FILL FILL_2__6929_ (
);

FILL FILL_0__6911_ (
);

FILL FILL_2__6509_ (
);

FILL FILL_1__12796_ (
);

FILL FILL_1__12376_ (
);

FILL FILL_0__9383_ (
);

FILL FILL_0__11789_ (
);

NOR2X1 _11654_ (
    .A(_5565_),
    .B(_5564_),
    .Y(_5566_)
);

FILL FILL_0__11369_ (
);

NAND3X1 _11234_ (
    .A(_4411_),
    .B(_4415_),
    .C(_4418_),
    .Y(_4431_)
);

FILL FILL_0__12730_ (
);

FILL FILL_0__12310_ (
);

FILL FILL_1__7398_ (
);

NOR2X1 _9802_ (
    .A(_3145_),
    .B(_3144_),
    .Y(_3146_)
);

NAND2X1 _12859_ (
    .A(\X[6] [3]),
    .B(gnd),
    .Y(_5897_)
);

INVX1 _12439_ (
    .A(\u_fir_pe6.mul [14]),
    .Y(_5543_)
);

OAI21X1 _12019_ (
    .A(_5123_),
    .B(_5127_),
    .C(_5130_),
    .Y(_5137_)
);

FILL FILL_2__6682_ (
);

FILL FILL_3__11095_ (
);

FILL FILL_2__10088_ (
);

FILL FILL_1__9964_ (
);

FILL FILL_1__9544_ (
);

FILL FILL_1__9124_ (
);

NAND2X1 _8194_ (
    .A(gnd),
    .B(\X[2] [2]),
    .Y(_1636_)
);

FILL FILL_1__10862_ (
);

FILL FILL_1__10442_ (
);

FILL FILL_1__10022_ (
);

FILL FILL_2__7887_ (
);

FILL FILL_2__7467_ (
);

FILL FILL_2__7047_ (
);

NAND2X1 _12192_ (
    .A(_5113_),
    .B(_5187_),
    .Y(_5307_)
);

FILL FILL_3__13241_ (
);

OAI21X1 _6927_ (
    .A(_74_),
    .B(_305_),
    .C(_479_),
    .Y(_522_)
);

AOI21X1 _6507_ (
    .A(_103_),
    .B(_104_),
    .C(_102_),
    .Y(_108_)
);

FILL FILL_2__12654_ (
);

FILL FILL_2__12234_ (
);

AOI21X1 _9399_ (
    .A(_2756_),
    .B(_2755_),
    .C(_2691_),
    .Y(_2757_)
);

FILL FILL_1__11647_ (
);

FILL FILL_1__11227_ (
);

FILL FILL_0__8654_ (
);

FILL FILL_3__6751_ (
);

FILL FILL_0__8234_ (
);

INVX1 _10925_ (
    .A(_4124_),
    .Y(_4125_)
);

NOR2X1 _10505_ (
    .A(_3774_),
    .B(_3778_),
    .Y(_3984_[12])
);

BUFX2 _13397_ (
    .A(_6376_[3]),
    .Y(Xout[3])
);

FILL FILL_2__9613_ (
);

FILL FILL_1__6669_ (
);

FILL FILL_2__13019_ (
);

FILL FILL_1__7610_ (
);

FILL FILL_0__9439_ (
);

FILL FILL_3__7536_ (
);

FILL FILL_0__9019_ (
);

NAND3X1 _6680_ (
    .A(_277_),
    .B(_278_),
    .C(_276_),
    .Y(_279_)
);

FILL FILL_3__10366_ (
);

FILL FILL_0__10393_ (
);

FILL FILL_1__8815_ (
);

FILL FILL_2__10300_ (
);

NAND2X1 _7885_ (
    .A(_1396_),
    .B(_1397_),
    .Y(_1398_)
);

AOI22X1 _7465_ (
    .A(_908_),
    .B(_903_),
    .C(_980_),
    .D(_984_),
    .Y(_985_)
);

NOR2X1 _7045_ (
    .A(_632_),
    .B(_633_),
    .Y(_634_)
);

FILL FILL_2__13192_ (
);

FILL FILL_0__6720_ (
);

FILL FILL_2__6738_ (
);

FILL FILL_1__12185_ (
);

FILL FILL_0__9192_ (
);

NOR2X1 _11883_ (
    .A(_4995_),
    .B(_4997_),
    .Y(_5002_)
);

AND2X2 _11463_ (
    .A(_4648_),
    .B(_4647_),
    .Y(_4775_[4])
);

FILL FILL_0__11178_ (
);

NAND3X1 _11043_ (
    .A(_4238_),
    .B(_4237_),
    .C(_4241_),
    .Y(_4242_)
);

FILL FILL_3__12932_ (
);

FILL FILL_2__11925_ (
);

FILL FILL_2__11505_ (
);

FILL FILL_1__10918_ (
);

FILL FILL_0__7925_ (
);

FILL FILL_0__7505_ (
);

INVX1 _9611_ (
    .A(_2962_),
    .Y(_2965_)
);

FILL FILL_3__8494_ (
);

OAI21X1 _12668_ (
    .A(_5707_),
    .B(_5708_),
    .C(_5706_),
    .Y(_5709_)
);

NAND3X1 _12248_ (
    .A(_5343_),
    .B(_5360_),
    .C(_5359_),
    .Y(_5362_)
);

FILL FILL_0__13324_ (
);

FILL FILL_2__6491_ (
);

FILL FILL_3__6807_ (
);

FILL FILL_1__9773_ (
);

FILL FILL_1__9353_ (
);

FILL FILL_3__9279_ (
);

FILL FILL_1__10671_ (
);

FILL FILL_1__10251_ (
);

FILL FILL_2__7696_ (
);

FILL FILL_2__7276_ (
);

NAND2X1 _6736_ (
    .A(_325_),
    .B(_333_),
    .Y(_334_)
);

FILL FILL_2__12883_ (
);

FILL FILL_2__12043_ (
);

FILL FILL_1__11876_ (
);

FILL FILL_1__11456_ (
);

FILL FILL_1__11036_ (
);

FILL FILL_0__8883_ (
);

FILL FILL_3__6980_ (
);

FILL FILL_0__8463_ (
);

FILL FILL_0__10869_ (
);

FILL FILL_0__10449_ (
);

DFFPOSX1 _10734_ (
    .D(\Y[4] [3]),
    .CLK(clk_bF$buf55),
    .Q(\u_fir_pe4.rYin [3])
);

FILL FILL_0__8043_ (
);

OAI22X1 _10314_ (
    .A(_3442_),
    .B(_3589_),
    .C(_3512_),
    .D(_3590_),
    .Y(_3591_)
);

FILL FILL_0__10029_ (
);

FILL FILL_2__9422_ (
);

FILL FILL_0__11810_ (
);

FILL FILL_1__6898_ (
);

FILL FILL_1__6478_ (
);

FILL FILL_2__13248_ (
);

FILL FILL_3_CLKBUF1_insert41 (
);

FILL FILL_3_CLKBUF1_insert43 (
);

FILL FILL_3_CLKBUF1_insert45 (
);

FILL FILL_3_CLKBUF1_insert47 (
);

FILL FILL_3_CLKBUF1_insert49 (
);

FILL FILL_0__9668_ (
);

FILL FILL_3__7765_ (
);

FILL FILL_0__9248_ (
);

AOI21X1 _11939_ (
    .A(_4966_),
    .B(_4964_),
    .C(_5057_),
    .Y(_5058_)
);

NAND2X1 _11519_ (
    .A(_4702_),
    .B(_4701_),
    .Y(_4775_[9])
);

FILL FILL_1__8624_ (
);

FILL FILL_1__8204_ (
);

NAND2X1 _7694_ (
    .A(_1210_),
    .B(_1206_),
    .Y(_1211_)
);

NAND2X1 _7274_ (
    .A(gnd),
    .B(\X[1] [2]),
    .Y(_797_)
);

FILL FILL_3__9911_ (
);

FILL FILL_2__6967_ (
);

FILL FILL_2__6547_ (
);

OAI22X1 _11692_ (
    .A(_4812_),
    .B(_4813_),
    .C(_4782_),
    .D(_4786_),
    .Y(_4814_)
);

AND2X2 _11272_ (
    .A(_4461_),
    .B(_4467_),
    .Y(_4468_)
);

FILL FILL_1__9829_ (
);

FILL FILL_1__9409_ (
);

FILL FILL_3__12741_ (
);

FILL FILL_3__12321_ (
);

FILL FILL_2__11734_ (
);

FILL FILL_2__11314_ (
);

NAND2X1 _8899_ (
    .A(_2322_),
    .B(_2317_),
    .Y(_2323_)
);

OAI21X1 _8479_ (
    .A(_1834_),
    .B(_1842_),
    .C(_1841_),
    .Y(_1917_)
);

NOR2X1 _8059_ (
    .A(_1561_),
    .B(_1555_),
    .Y(_1563_)
);

FILL FILL_1__10307_ (
);

FILL FILL_0__7734_ (
);

DFFPOSX1 _9840_ (
    .D(_3181_[10]),
    .CLK(clk_bF$buf26),
    .Q(\Y[4] [10])
);

FILL FILL_0__7314_ (
);

NAND2X1 _9420_ (
    .A(\X[3] [2]),
    .B(gnd),
    .Y(_2777_)
);

FILL FILL_1__13199_ (
);

DFFPOSX1 _9000_ (
    .D(_2390_[7]),
    .CLK(clk_bF$buf51),
    .Q(\u_fir_pe2.mul [7])
);

AOI21X1 _12897_ (
    .A(_5934_),
    .B(_5933_),
    .C(_5932_),
    .Y(_5935_)
);

DFFPOSX1 _12477_ (
    .D(\X[7] [0]),
    .CLK(clk_bF$buf29),
    .Q(_6376_[0])
);

INVX1 _12057_ (
    .A(_5168_),
    .Y(_5174_)
);

FILL FILL_3__13106_ (
);

FILL FILL_2__12939_ (
);

FILL FILL_2__12519_ (
);

FILL FILL_0__13133_ (
);

FILL FILL_0__8939_ (
);

FILL FILL_0__8519_ (
);

FILL FILL_3__6616_ (
);

FILL FILL_1__9582_ (
);

FILL FILL_1__9162_ (
);

FILL FILL_1__10480_ (
);

FILL FILL_1__10060_ (
);

FILL FILL_2__7085_ (
);

AOI21X1 _6965_ (
    .A(_556_),
    .B(_457_),
    .C(_558_),
    .Y(_559_)
);

NAND2X1 _6545_ (
    .A(Xin[2]),
    .B(gnd),
    .Y(_145_)
);

FILL FILL_2__12692_ (
);

FILL FILL_2__12272_ (
);

FILL FILL_1__11685_ (
);

FILL FILL_1__11265_ (
);

FILL FILL_0__8692_ (
);

FILL FILL_0__8272_ (
);

FILL FILL_0__10678_ (
);

INVX1 _10963_ (
    .A(_4081_),
    .Y(_4163_)
);

INVX1 _10543_ (
    .A(_3809_),
    .Y(_3815_)
);

FILL FILL_0__10258_ (
);

AND2X2 _10123_ (
    .A(_3333_),
    .B(_3337_),
    .Y(_3402_)
);

FILL FILL_2__9651_ (
);

FILL FILL_2__9231_ (
);

FILL FILL_2__13057_ (
);

FILL FILL_0__9897_ (
);

FILL FILL_3__7994_ (
);

FILL FILL_0__9477_ (
);

FILL FILL_0__9057_ (
);

AND2X2 _11748_ (
    .A(vdd),
    .B(\X[7] [3]),
    .Y(_4869_)
);

AOI21X1 _11328_ (
    .A(_4400_),
    .B(_4392_),
    .C(_4470_),
    .Y(_4523_)
);

FILL FILL_1__13411_ (
);

FILL FILL_0__12824_ (
);

FILL FILL_0__12404_ (
);

FILL FILL254550x180150 (
);

FILL FILL_1__8853_ (
);

FILL FILL_1__8433_ (
);

FILL FILL_1__8013_ (
);

FILL FILL_3__8779_ (
);

NOR2X1 _7083_ (
    .A(\u_fir_pe0.rYin [5]),
    .B(\u_fir_pe0.mul [5]),
    .Y(_668_)
);

FILL FILL_3__9720_ (
);

FILL FILL_3__9300_ (
);

FILL FILL_2__6776_ (
);

FILL FILL_3__11189_ (
);

FILL FILL254550x147750 (
);

AND2X2 _11081_ (
    .A(_4279_),
    .B(_4275_),
    .Y(_4781_[7])
);

FILL FILL_1__9638_ (
);

FILL FILL_1__9218_ (
);

FILL FILL_2__11963_ (
);

FILL FILL_2__11543_ (
);

FILL FILL_2__11123_ (
);

OR2X2 _8288_ (
    .A(_1727_),
    .B(_1725_),
    .Y(_1728_)
);

FILL FILL_1__10956_ (
);

FILL FILL_1__10536_ (
);

FILL FILL_1__10116_ (
);

FILL FILL_0__7963_ (
);

FILL FILL_0__7543_ (
);

FILL FILL_0__7123_ (
);

OAI21X1 _12286_ (
    .A(_5366_),
    .B(_5391_),
    .C(_5390_),
    .Y(_5398_)
);

FILL FILL_2__8922_ (
);

FILL FILL_2__8502_ (
);

FILL FILL_3__13335_ (
);

FILL FILL_2__12748_ (
);

FILL FILL_2__12328_ (
);

FILL FILL_0__8748_ (
);

FILL FILL_3__6845_ (
);

FILL FILL_0__8328_ (
);

FILL FILL_3__6425_ (
);

FILL FILL_1__9391_ (
);

FILL FILL_2__9707_ (
);

FILL FILL_1__7704_ (
);

NAND3X1 _6774_ (
    .A(_369_),
    .B(_370_),
    .C(_371_),
    .Y(_372_)
);

FILL FILL_2__12081_ (
);

FILL FILL_1__11494_ (
);

FILL FILL_1__11074_ (
);

FILL FILL_0__10487_ (
);

INVX2 _10772_ (
    .A(vdd),
    .Y(_4763_)
);

OAI21X1 _10352_ (
    .A(_3628_),
    .B(_3627_),
    .C(_3626_),
    .Y(_3629_)
);

FILL FILL_0__10067_ (
);

FILL FILL_1__8909_ (
);

FILL FILL_3__11821_ (
);

FILL FILL_3__11401_ (
);

FILL FILL_2__10814_ (
);

FILL FILL_2__9460_ (
);

FILL FILL_2__9040_ (
);

OAI21X1 _7979_ (
    .A(_1480_),
    .B(_1481_),
    .C(_1477_),
    .Y(_1482_)
);

INVX1 _7559_ (
    .A(_932_),
    .Y(_1078_)
);

INVX1 _7139_ (
    .A(_722_),
    .Y(_723_)
);

FILL FILL_2__13286_ (
);

FILL FILL_0__6814_ (
);

OAI21X1 _8920_ (
    .A(_2336_),
    .B(_2337_),
    .C(_2341_),
    .Y(_2343_)
);

FILL FILL_1__12699_ (
);

OAI21X1 _8500_ (
    .A(_1929_),
    .B(_1923_),
    .C(_1931_),
    .Y(_1938_)
);

FILL FILL_1__12279_ (
);

FILL FILL_0__9286_ (
);

NAND2X1 _11977_ (
    .A(_5088_),
    .B(_5089_),
    .Y(_5095_)
);

FILL FILL_3__7383_ (
);

NAND2X1 _11557_ (
    .A(_4740_),
    .B(_4734_),
    .Y(_4741_)
);

NAND3X1 _11137_ (
    .A(_4307_),
    .B(_4325_),
    .C(_4321_),
    .Y(_4335_)
);

FILL FILL_3__12606_ (
);

FILL FILL_1__13220_ (
);

FILL FILL_0__12633_ (
);

FILL FILL_0__12213_ (
);

INVX1 _9705_ (
    .A(_3041_),
    .Y(_3051_)
);

FILL FILL_1__8662_ (
);

FILL FILL_1__8242_ (
);

FILL FILL_3__8588_ (
);

FILL FILL_3__8168_ (
);

FILL FILL_2__6585_ (
);

FILL FILL_1__9447_ (
);

FILL FILL_1__9027_ (
);

FILL FILL_2__11772_ (
);

FILL FILL_2__11352_ (
);

DFFPOSX1 _8097_ (
    .D(\X[1]_5_bF$buf1 ),
    .CLK(clk_bF$buf7),
    .Q(\X[2] [5])
);

FILL FILL_1__10765_ (
);

FILL FILL_1__10345_ (
);

FILL FILL_0__7772_ (
);

FILL FILL_0__7352_ (
);

OAI21X1 _12095_ (
    .A(_5211_),
    .B(_5210_),
    .C(_5209_),
    .Y(_5212_)
);

FILL FILL_2__8731_ (
);

FILL FILL_2__8311_ (
);

FILL FILL253350x230550 (
);

FILL FILL_2__12977_ (
);

FILL FILL_2__12557_ (
);

FILL FILL_2__12137_ (
);

FILL FILL_0__13171_ (
);

FILL FILL_0__8557_ (
);

FILL FILL_0__8137_ (
);

NAND3X1 _10828_ (
    .A(_4017_),
    .B(_4029_),
    .C(_4025_),
    .Y(_4030_)
);

INVX1 _10408_ (
    .A(_3648_),
    .Y(_3684_)
);

FILL FILL_1__12911_ (
);

FILL FILL_2__9936_ (
);

FILL FILL_0__11904_ (
);

FILL FILL_2__9516_ (
);

FILL FILL_1__7933_ (
);

FILL FILL_1__7513_ (
);

FILL FILL_3__7859_ (
);

FILL FILL_3__7019_ (
);

NAND3X1 _6583_ (
    .A(_136_),
    .B(_177_),
    .C(_182_),
    .Y(_183_)
);

FILL FILL_3__10689_ (
);

FILL FILL_0__10296_ (
);

NOR2X1 _10581_ (
    .A(_3846_),
    .B(_3845_),
    .Y(_3847_)
);

AOI22X1 _10161_ (
    .A(_3275_),
    .B(_3346_),
    .C(_3349_),
    .D(_3345_),
    .Y(_3440_)
);

FILL FILL_1__8718_ (
);

FILL FILL_3__11210_ (
);

FILL FILL_2__10623_ (
);

FILL FILL_2__10203_ (
);

AOI21X1 _7788_ (
    .A(_1252_),
    .B(_1255_),
    .C(_1303_),
    .Y(_1304_)
);

NAND3X1 _7368_ (
    .A(vdd),
    .B(\X[1] [3]),
    .C(_880_),
    .Y(_889_)
);

FILL FILL_2__13095_ (
);

FILL FILL_0__6623_ (
);

FILL FILL_1__12088_ (
);

FILL FILL_0__9095_ (
);

NAND3X1 _11786_ (
    .A(_4905_),
    .B(_4906_),
    .C(_4904_),
    .Y(_4907_)
);

FILL FILL_3__7192_ (
);

OAI21X1 _11366_ (
    .A(_4558_),
    .B(_4559_),
    .C(_4511_),
    .Y(_4560_)
);

FILL FILL_3__12835_ (
);

FILL FILL_3__12415_ (
);

FILL FILL_2__11828_ (
);

FILL FILL_0__12862_ (
);

FILL FILL_2__11408_ (
);

FILL FILL_0__12442_ (
);

FILL FILL_0__12022_ (
);

FILL FILL_0__7828_ (
);

NOR2X1 _9934_ (
    .A(_3215_),
    .B(_3214_),
    .Y(_3216_)
);

FILL FILL_0__7408_ (
);

NAND2X1 _9514_ (
    .A(_2868_),
    .B(_2869_),
    .Y(_2870_)
);

FILL FILL_1__8891_ (
);

FILL FILL_1__8471_ (
);

FILL FILL_1__8051_ (
);

FILL FILL_3__8397_ (
);

FILL FILL_0__13227_ (
);

FILL FILL_2__6394_ (
);

FILL FILL_1__9676_ (
);

FILL FILL_1__9256_ (
);

FILL FILL_2__11581_ (
);

FILL FILL_2__11161_ (
);

FILL FILL_1__10994_ (
);

FILL FILL_1__10574_ (
);

FILL FILL_1__10154_ (
);

FILL FILL_2__7599_ (
);

FILL FILL_0__7581_ (
);

FILL FILL_2__7179_ (
);

FILL FILL_0__7161_ (
);

FILL FILL_3__10901_ (
);

FILL FILL_2__8540_ (
);

FILL FILL254250x133350 (
);

NAND2X1 _6639_ (
    .A(_232_),
    .B(_237_),
    .Y(_238_)
);

FILL FILL_2__12786_ (
);

FILL FILL_2__12366_ (
);

FILL FILL_1__11779_ (
);

FILL FILL_1__11359_ (
);

FILL FILL_0__8786_ (
);

FILL FILL_0__8366_ (
);

FILL FILL_3__6463_ (
);

NOR2X1 _10637_ (
    .A(\u_fir_pe4.rYin [9]),
    .B(\u_fir_pe4.mul [9]),
    .Y(_3901_)
);

OAI21X1 _10217_ (
    .A(_3413_),
    .B(_3418_),
    .C(_3417_),
    .Y(_3495_)
);

FILL FILL_1__12720_ (
);

FILL FILL_1__12300_ (
);

FILL FILL_2__9745_ (
);

FILL FILL253950x72150 (
);

FILL FILL_2__9325_ (
);

FILL FILL_0__11713_ (
);

FILL FILL_1__7742_ (
);

FILL FILL_1__7322_ (
);

NOR2X1 _6392_ (
    .A(_783_),
    .B(_782_),
    .Y(_784_)
);

FILL FILL_0__12918_ (
);

FILL FILL_3__10078_ (
);

AND2X2 _10390_ (
    .A(\X[4]_5_bF$buf0 ),
    .B(vdd),
    .Y(_3666_)
);

FILL FILL_1__8947_ (
);

FILL FILL_1__8527_ (
);

FILL FILL_2__10852_ (
);

FILL FILL_2__10432_ (
);

FILL FILL_2__10012_ (
);

NAND2X1 _7597_ (
    .A(\X[1] [3]),
    .B(gnd),
    .Y(_1115_)
);

INVX1 _7177_ (
    .A(\u_fir_pe0.mul [14]),
    .Y(_761_)
);

FILL FILL_3__9814_ (
);

FILL FILL_0__6852_ (
);

FILL FILL_0__6432_ (
);

DFFPOSX1 _11595_ (
    .D(_4775_[11]),
    .CLK(clk_bF$buf35),
    .Q(\Y[6] [11])
);

NOR2X1 _11175_ (
    .A(_4303_),
    .B(_4306_),
    .Y(_4372_)
);

FILL FILL_2__7811_ (
);

FILL FILL_0__12671_ (
);

FILL FILL_2__11217_ (
);

FILL FILL_0__12251_ (
);

FILL FILL_0__7637_ (
);

OAI21X1 _9743_ (
    .A(_3056_),
    .B(_3057_),
    .C(_3085_),
    .Y(_3086_)
);

NOR2X1 _9323_ (
    .A(_2598_),
    .B(_2595_),
    .Y(_2682_)
);

FILL FILL_1__8280_ (
);

FILL FILL_0__13036_ (
);

NOR2X1 _13321_ (
    .A(_6343_),
    .B(_6337_),
    .Y(_6345_)
);

FILL FILL_3__6939_ (
);

FILL FILL_3__6519_ (
);

FILL FILL_1__9485_ (
);

FILL FILL_1__9065_ (
);

FILL FILL_2__11390_ (
);

FILL FILL_1__10383_ (
);

FILL FILL_0__7390_ (
);

FILL FILL_3__13182_ (
);

OAI22X1 _6868_ (
    .A(_417_),
    .B(_305_),
    .C(_25_),
    .D(_416_),
    .Y(_464_)
);

NAND2X1 _6448_ (
    .A(_32_),
    .B(_47_),
    .Y(_50_)
);

FILL FILL_2__12595_ (
);

FILL FILL_2__12175_ (
);

FILL FILL_1__11168_ (
);

FILL FILL_0__8595_ (
);

FILL FILL_3__6692_ (
);

FILL FILL_0__8175_ (
);

AND2X2 _10866_ (
    .A(_4062_),
    .B(_4066_),
    .Y(_4067_)
);

AND2X2 _10446_ (
    .A(_3711_),
    .B(_3707_),
    .Y(_3721_)
);

NAND3X1 _10026_ (
    .A(_3242_),
    .B(_3305_),
    .C(_3306_),
    .Y(_3307_)
);

FILL FILL_3__11915_ (
);

FILL FILL_2__10908_ (
);

FILL FILL_2__9974_ (
);

FILL FILL_2__9554_ (
);

FILL FILL_0__11942_ (
);

FILL FILL_2__9134_ (
);

FILL FILL_0__11522_ (
);

FILL FILL_0__11102_ (
);

FILL FILL_0__6908_ (
);

FILL FILL_1__7971_ (
);

FILL FILL_1__7551_ (
);

FILL FILL_1__7131_ (
);

FILL FILL_3__7477_ (
);

FILL FILL_3__7057_ (
);

FILL FILL_1__13314_ (
);

FILL FILL_0__12727_ (
);

FILL FILL_0__12307_ (
);

FILL FILL_1__8756_ (
);

FILL FILL_1__8336_ (
);

FILL FILL_2__10661_ (
);

FILL FILL_2__10241_ (
);

FILL FILL_0__6661_ (
);

FILL FILL_2__6679_ (
);

FILL FILL_3__12873_ (
);

FILL FILL_2__7620_ (
);

FILL FILL_3__12033_ (
);

FILL FILL_2__11866_ (
);

FILL FILL_2__11446_ (
);

FILL FILL_2__11026_ (
);

FILL FILL_0__12060_ (
);

FILL FILL_1__10859_ (
);

FILL FILL_1__10439_ (
);

FILL FILL_1__10019_ (
);

FILL FILL_0__7866_ (
);

OAI21X1 _9972_ (
    .A(_3241_),
    .B(_3253_),
    .C(_3247_),
    .Y(_3254_)
);

FILL FILL_0__7446_ (
);

NAND2X1 _9552_ (
    .A(_2875_),
    .B(_2878_),
    .Y(_2907_)
);

FILL FILL_0__7026_ (
);

NAND2X1 _9132_ (
    .A(_2472_),
    .B(_2468_),
    .Y(_2493_)
);

FILL FILL_1__11800_ (
);

OAI21X1 _12189_ (
    .A(_4856_),
    .B(_5087_),
    .C(_5261_),
    .Y(_5304_)
);

FILL FILL_2__8825_ (
);

FILL FILL_2__8405_ (
);

FILL FILL_0__13265_ (
);

NAND2X1 _13130_ (
    .A(_6161_),
    .B(_6163_),
    .Y(_6164_)
);

FILL FILL_1__6822_ (
);

FILL FILL_1__6402_ (
);

FILL FILL_1__9294_ (
);

FILL FILL_2_CLKBUF1_insert50 (
);

FILL FILL_2_CLKBUF1_insert51 (
);

FILL FILL_2_CLKBUF1_insert52 (
);

FILL FILL_2_CLKBUF1_insert53 (
);

FILL FILL_2_CLKBUF1_insert54 (
);

FILL FILL_2_CLKBUF1_insert55 (
);

FILL FILL_2_CLKBUF1_insert56 (
);

FILL FILL_2_CLKBUF1_insert57 (
);

FILL FILL_2_CLKBUF1_insert58 (
);

FILL FILL_2_CLKBUF1_insert59 (
);

FILL FILL_1__10192_ (
);

FILL FILL_1__7607_ (
);

AOI21X1 _6677_ (
    .A(_184_),
    .B(_182_),
    .C(_275_),
    .Y(_276_)
);

FILL FILL_1__11397_ (
);

INVX1 _10675_ (
    .A(\u_fir_pe4.rYin [13]),
    .Y(_3939_)
);

AOI21X1 _10255_ (
    .A(_3532_),
    .B(_3531_),
    .C(_3530_),
    .Y(_3533_)
);

FILL FILL_3__11304_ (
);

FILL FILL_2__9783_ (
);

FILL FILL_2__9363_ (
);

FILL FILL_0__11751_ (
);

FILL FILL_0__11331_ (
);

FILL FILL_2__13189_ (
);

FILL FILL_0__6717_ (
);

INVX1 _8823_ (
    .A(\u_fir_pe2.rYin [4]),
    .Y(_2249_)
);

AOI22X1 _8403_ (
    .A(vdd),
    .B(\X[2] [4]),
    .C(gnd),
    .D(\X[2]_5_bF$buf3 ),
    .Y(_1842_)
);

FILL FILL_1__7780_ (
);

FILL FILL_1__7360_ (
);

FILL FILL_0__9189_ (
);

FILL FILL_3__12929_ (
);

FILL FILL_1__13123_ (
);

FILL FILL_0__12956_ (
);

INVX1 _12821_ (
    .A(_5714_),
    .Y(_5860_)
);

FILL FILL_0__12536_ (
);

FILL FILL_0__12116_ (
);

INVX1 _12401_ (
    .A(_5504_),
    .Y(_5505_)
);

NAND2X1 _9608_ (
    .A(_2956_),
    .B(_2960_),
    .Y(_2962_)
);

FILL FILL_1__8565_ (
);

FILL FILL_1__8145_ (
);

FILL FILL_2__10890_ (
);

FILL FILL_2__10470_ (
);

FILL FILL_2__10050_ (
);

FILL FILL_3__9432_ (
);

FILL FILL_3__9012_ (
);

FILL FILL_0__6890_ (
);

FILL FILL_0__6470_ (
);

FILL FILL_2__6488_ (
);

FILL FILL_3__12682_ (
);

FILL FILL_3__12262_ (
);

FILL FILL_2__11675_ (
);

FILL FILL_2__11255_ (
);

FILL FILL_1__10668_ (
);

FILL FILL_1__10248_ (
);

FILL FILL254550x10950 (
);

FILL FILL_0__7675_ (
);

NOR2X1 _9781_ (
    .A(\u_fir_pe3.rYin [11]),
    .B(\u_fir_pe3.mul [11]),
    .Y(_3125_)
);

FILL FILL_0__7255_ (
);

OAI21X1 _9361_ (
    .A(_2480_),
    .B(_2535_),
    .C(_2718_),
    .Y(_2719_)
);

FILL FILL253950x158550 (
);

FILL FILL_2__8634_ (
);

FILL FILL_2__8214_ (
);

FILL FILL_0__10602_ (
);

FILL FILL_3__13047_ (
);

FILL FILL_0__13074_ (
);

FILL FILL_1__6631_ (
);

FILL FILL_2__13401_ (
);

FILL FILL_3__6557_ (
);

FILL FILL_1__12814_ (
);

FILL FILL_0__9821_ (
);

FILL FILL_2__9419_ (
);

FILL FILL_0__9401_ (
);

FILL FILL_0__11807_ (
);

FILL FILL_1__7836_ (
);

FILL FILL_1__7416_ (
);

AND2X2 _6486_ (
    .A(vdd),
    .B(Xin[3]),
    .Y(_87_)
);

FILL FILL_3__8703_ (
);

OR2X2 _10484_ (
    .A(_3757_),
    .B(_3753_),
    .Y(_3758_)
);

FILL FILL_0__10199_ (
);

NAND2X1 _10064_ (
    .A(vdd),
    .B(\X[4]_5_bF$buf3 ),
    .Y(_3344_)
);

FILL FILL_2__6700_ (
);

FILL FILL_2__10946_ (
);

FILL FILL_0__11980_ (
);

FILL FILL_2__9592_ (
);

FILL FILL_2__10526_ (
);

FILL FILL_2__9172_ (
);

FILL FILL_0__11560_ (
);

FILL FILL_2__10106_ (
);

FILL FILL_0__11140_ (
);

FILL FILL_0__6946_ (
);

FILL FILL_0__6526_ (
);

NOR2X1 _8632_ (
    .A(_2067_),
    .B(_2010_),
    .Y(_2068_)
);

OR2X2 _8212_ (
    .A(_1653_),
    .B(_1652_),
    .Y(_1654_)
);

endmodule
