magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect 13 71 57 79
rect -7 39 57 71
rect -7 30 37 39
<< nwell >>
rect -6 77 57 136
<< ntransistor >>
rect 9 7 11 27
rect 19 7 21 27
rect 29 7 31 27
rect 39 7 41 27
<< ptransistor >>
rect 9 83 11 123
rect 19 83 21 123
rect 29 83 31 123
rect 39 83 41 123
<< ndiffusion >>
rect 8 7 9 27
rect 11 7 12 27
rect 18 7 19 27
rect 21 7 22 27
rect 28 7 29 27
rect 31 7 32 27
rect 38 7 39 27
rect 41 7 42 27
<< pdiffusion >>
rect 8 83 9 123
rect 11 83 12 123
rect 18 83 19 123
rect 21 83 22 123
rect 28 83 29 123
rect 31 83 32 123
rect 38 83 39 123
rect 41 83 42 123
<< ndcontact >>
rect 2 7 8 27
rect 12 7 18 27
rect 22 7 28 27
rect 32 7 38 27
rect 42 7 48 27
<< pdcontact >>
rect 2 83 8 123
rect 12 83 18 123
rect 22 83 28 123
rect 32 83 38 123
rect 42 83 48 123
<< psubstratepcontact >>
rect -3 -3 53 3
<< nsubstratencontact >>
rect -3 127 53 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 39 123 41 125
rect 9 82 11 83
rect 19 82 21 83
rect 29 82 31 83
rect 39 82 41 83
rect 9 80 41 82
rect 9 64 11 80
rect 9 58 12 64
rect 9 31 11 58
rect 9 29 41 31
rect 9 27 11 29
rect 19 27 21 29
rect 29 27 31 29
rect 39 27 41 29
rect 9 5 11 7
rect 19 5 21 7
rect 29 5 31 7
rect 39 5 41 7
<< polycontact >>
rect 12 58 18 64
<< metal1 >>
rect -3 133 53 134
rect -3 126 53 127
rect 2 123 8 126
rect 22 123 28 126
rect 42 123 48 126
rect 12 80 18 83
rect 32 80 36 83
rect 12 77 36 80
rect 32 58 36 77
rect 32 34 36 51
rect 12 30 36 34
rect 12 27 16 30
rect 32 27 36 30
rect 2 4 8 7
rect 22 4 28 7
rect 42 4 48 7
rect -3 3 53 4
rect -3 -4 53 -3
<< m2contact >>
rect 12 51 19 58
rect 32 51 39 58
<< metal2 >>
rect 33 58 37 67
rect 13 43 17 51
<< m1p >>
rect -3 126 53 134
rect -3 -4 53 4
<< m2p >>
rect 33 59 37 67
rect 13 43 17 50
<< labels >>
rlabel metal2 15 44 15 44 1 A
port 1 n signal input
rlabel metal2 35 65 35 65 1 Y
port 2 n signal output
rlabel metal1 -3 126 53 134 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -3 -4 53 4 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 50 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
