magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -56 -56 84 404
<< genericcontact >>
rect 11 325 17 331
rect 11 297 17 303
rect 11 269 17 275
rect 11 241 17 247
rect 11 213 17 219
rect 11 185 17 191
rect 11 157 17 163
rect 11 129 17 135
rect 11 101 17 107
rect 11 73 17 79
rect 11 45 17 51
rect 11 17 17 23
<< metal1 >>
rect 4 4 24 344
<< end >>
