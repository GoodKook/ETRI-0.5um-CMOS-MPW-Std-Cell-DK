magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -60 -60 330 330
<< psubstratepdiff >>
rect 85 85 185 185
<< metal1 >>
rect 85 85 185 185
use ntap_ring_pdiode_CDNS_7230122529128  ntap_ring_pdiode_CDNS_7230122529128_0
timestamp 1569140870
transform 1 0 0 0 1 0
box 0 0 270 270
use ptap_CDNS_7230122529127  ptap_CDNS_7230122529127_0
timestamp 1569140870
transform 1 0 82 0 1 82
box 4 4 102 102
<< end >>
