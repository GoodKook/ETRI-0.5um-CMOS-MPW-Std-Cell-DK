magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -17 71 57 79
rect -17 39 67 71
rect -7 30 67 39
<< nwell >>
rect -6 77 57 136
rect 6 73 39 77
<< ntransistor >>
rect 9 11 11 21
rect 19 11 21 31
rect 24 11 26 31
rect 34 11 36 31
rect 39 11 41 31
<< ptransistor >>
rect 9 99 11 119
rect 19 79 21 119
rect 24 79 26 119
rect 34 83 36 123
rect 39 83 41 123
<< ndiffusion >>
rect 12 29 19 31
rect 8 11 9 21
rect 11 13 12 21
rect 18 13 19 29
rect 11 11 19 13
rect 21 11 24 31
rect 26 27 34 31
rect 26 11 27 27
rect 33 11 34 27
rect 36 11 39 31
rect 41 11 42 31
<< pdiffusion >>
rect 8 99 9 119
rect 11 99 12 119
rect 18 85 19 119
rect 14 79 19 85
rect 21 79 24 119
rect 26 87 27 119
rect 33 87 34 123
rect 26 83 34 87
rect 36 83 39 123
rect 41 83 42 123
rect 26 79 29 83
<< ndcontact >>
rect 2 11 8 21
rect 12 13 18 29
rect 27 11 33 27
rect 42 11 48 31
<< pdcontact >>
rect 2 99 8 119
rect 12 85 18 119
rect 27 87 33 123
rect 42 83 48 123
<< psubstratepcontact >>
rect -3 -3 53 3
<< nsubstratencontact >>
rect -3 127 53 133
<< polysilicon >>
rect 9 124 26 126
rect 9 119 11 124
rect 19 119 21 121
rect 24 119 26 124
rect 34 123 36 125
rect 39 123 41 125
rect 9 98 11 99
rect 4 96 11 98
rect 4 51 6 96
rect 19 72 21 79
rect 24 77 26 79
rect 34 72 36 83
rect 13 70 21 72
rect 26 70 36 72
rect 13 64 15 70
rect 26 64 28 70
rect 4 24 6 45
rect 13 34 15 58
rect 13 32 21 34
rect 19 31 21 32
rect 24 31 26 58
rect 34 31 36 33
rect 39 31 41 83
rect 4 22 11 24
rect 9 21 11 22
rect 9 6 11 11
rect 19 9 21 11
rect 24 9 26 11
rect 34 6 36 11
rect 39 9 41 11
rect 9 4 36 6
<< polycontact >>
rect 12 58 18 64
rect 22 58 28 64
rect 2 45 8 51
rect 41 58 47 64
<< metal1 >>
rect -3 133 53 134
rect -3 126 53 127
rect 12 119 18 126
rect 42 123 48 126
rect 2 82 5 99
rect 33 87 34 88
rect 27 85 34 87
rect 2 79 28 82
rect 24 64 28 79
rect 31 58 34 85
rect 22 35 26 58
rect 2 32 26 35
rect 2 21 5 32
rect 31 29 34 51
rect 27 27 34 29
rect 12 4 16 13
rect 33 26 34 27
rect 42 4 46 11
rect -3 3 53 4
rect -3 -4 53 -3
<< m2contact >>
rect 2 51 9 58
rect 12 51 19 58
rect 31 51 38 58
rect 41 51 48 58
<< metal2 >>
rect 3 58 7 67
rect 33 58 37 67
rect 13 43 17 51
rect 43 43 47 51
<< m1p >>
rect -3 126 53 134
rect -3 -4 53 4
<< m2p >>
rect 3 59 7 67
rect 33 59 37 67
rect 13 43 17 50
rect 43 43 47 50
<< labels >>
rlabel metal2 45 45 45 45 1 A
port 1 n signal input
rlabel metal2 15 45 15 45 1 B
port 2 n signal input
rlabel metal2 5 65 5 65 1 S
port 3 n signal input
rlabel metal2 35 66 35 66 5 Y
port 4 n signal output
rlabel metal1 -3 126 53 134 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -3 -4 53 4 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 50 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
