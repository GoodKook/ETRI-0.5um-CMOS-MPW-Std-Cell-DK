magic
tech scmos
magscale 1 6
timestamp 1727178736
<< error_s >>
rect 12 18732 18408 18768
rect 12 17952 18408 17988
rect 12 17172 18408 17208
rect 12 16392 18408 16428
rect 12 15612 18408 15648
rect 12 14832 18408 14868
rect 12 14052 18408 14088
rect 12 13272 18408 13308
rect 12 12492 18408 12528
rect 12 11712 18408 11748
rect 12 10932 18408 10968
rect 12 10152 18408 10188
rect 12 9372 18408 9408
rect 12 8592 18408 8628
rect 12 7812 18408 7848
rect 12 7032 18408 7068
rect 12 6252 18408 6288
rect 12 5472 18408 5508
rect 12 4692 18408 4728
rect 12 3912 18408 3948
rect 12 3132 18408 3168
rect 12 2352 18408 2388
rect 12 1572 18408 1608
rect 12 792 18408 828
rect 12 12 18408 48
<< nwell >>
rect 17791 18648 18001 18672
rect 6600 11253 6645 11268
<< metal1 >>
rect -189 18726 90 18774
rect -189 17214 -9 18726
rect 6861 18411 6999 18429
rect 7641 18411 7959 18429
rect 16821 18411 17079 18429
rect 11739 18369 11781 18399
rect 11691 18360 11781 18369
rect 11691 18351 11769 18360
rect 11691 18261 11709 18351
rect 12081 18369 12120 18381
rect 17700 18369 17739 18381
rect 12081 18339 12129 18369
rect 12111 18261 12129 18339
rect 17691 18339 17739 18369
rect 13761 18309 13800 18321
rect 13761 18291 13842 18309
rect 13761 18279 13800 18291
rect 17691 18261 17709 18339
rect 11691 18231 11739 18261
rect 11700 18219 11739 18231
rect 12111 18231 12159 18261
rect 12120 18219 12159 18231
rect 14160 18249 14199 18261
rect 14151 18231 14199 18249
rect 14160 18219 14199 18231
rect 17691 18231 17739 18261
rect 17700 18219 17739 18231
rect 15561 18171 15759 18189
rect 18429 17994 18609 18774
rect 18330 17946 18609 17994
rect 8583 17811 8679 17829
rect 6441 17751 6579 17769
rect 8421 17751 8559 17769
rect 12861 17751 13059 17769
rect 621 17709 660 17721
rect 11100 17709 11139 17721
rect 621 17679 669 17709
rect 651 17601 669 17679
rect 11091 17679 11139 17709
rect 15921 17709 15960 17721
rect 16860 17709 16899 17721
rect 15921 17679 15969 17709
rect 11091 17601 11109 17679
rect 15951 17601 15969 17679
rect 621 17571 669 17601
rect 621 17559 660 17571
rect 8961 17571 9039 17589
rect 11040 17598 11109 17601
rect 11061 17571 11109 17598
rect 11061 17559 11100 17571
rect 15921 17571 15969 17601
rect 16851 17679 16899 17709
rect 16851 17601 16869 17679
rect 16851 17571 16899 17601
rect 15921 17559 15960 17571
rect 16860 17559 16899 17571
rect 7761 17511 7959 17529
rect 12561 17511 12699 17529
rect 16341 17511 16539 17529
rect -189 17166 90 17214
rect -189 15654 -9 17166
rect 1161 16851 1299 16869
rect 6801 16851 6879 16869
rect 9021 16851 9159 16869
rect 14661 16851 14739 16869
rect 6639 16809 6681 16839
rect 1581 16791 1749 16809
rect 6639 16800 6729 16809
rect 6651 16791 6729 16800
rect 1581 16671 1659 16689
rect 1731 16641 1749 16791
rect 6711 16689 6729 16791
rect 13161 16791 13329 16809
rect 13311 16701 13329 16791
rect 14481 16791 14649 16809
rect 14631 16701 14649 16791
rect 16440 16749 16479 16761
rect 15981 16731 16122 16749
rect 16431 16731 16479 16749
rect 16440 16719 16479 16731
rect 6711 16671 6819 16689
rect 13311 16671 13359 16701
rect 13320 16659 13359 16671
rect 14631 16671 14679 16701
rect 14640 16659 14679 16671
rect 1680 16638 1749 16641
rect 1701 16611 1749 16638
rect 1701 16599 1740 16611
rect 3321 16611 3459 16629
rect 10383 16611 10479 16629
rect 15441 16611 15579 16629
rect 15621 16611 15699 16629
rect 4941 16551 5139 16569
rect 5781 16491 5919 16509
rect 18429 16434 18609 17946
rect 18330 16386 18609 16434
rect 3231 16029 3249 16179
rect 7800 16149 7839 16161
rect 7791 16119 7839 16149
rect 8121 16149 8160 16161
rect 8121 16119 8169 16149
rect 8541 16149 8580 16161
rect 8880 16149 8919 16161
rect 8541 16119 8589 16149
rect 7791 16041 7809 16119
rect 8151 16041 8169 16119
rect 8571 16041 8589 16119
rect 3231 16011 3399 16029
rect 4551 16011 4659 16029
rect 7791 16011 7839 16041
rect 7800 15999 7839 16011
rect 8121 16011 8169 16041
rect 8121 15999 8160 16011
rect 8541 16011 8589 16041
rect 8871 16119 8919 16149
rect 9561 16149 9600 16161
rect 10140 16149 10179 16161
rect 9561 16119 9609 16149
rect 8871 16041 8889 16119
rect 9591 16041 9609 16119
rect 8871 16011 8919 16041
rect 8541 15999 8580 16011
rect 8880 15999 8919 16011
rect 9561 16011 9609 16041
rect 10131 16119 10179 16149
rect 10941 16149 10980 16161
rect 10941 16119 10989 16149
rect 13101 16149 13140 16161
rect 13101 16119 13149 16149
rect 10131 16041 10149 16119
rect 10971 16041 10989 16119
rect 13131 16041 13149 16119
rect 16791 16131 16899 16149
rect 16791 16041 16809 16131
rect 10131 16011 10179 16041
rect 9561 15999 9600 16011
rect 10140 15999 10179 16011
rect 10941 16011 10989 16041
rect 10941 15999 10980 16011
rect 12741 16011 12819 16029
rect 13101 16011 13149 16041
rect 13101 15999 13140 16011
rect 16761 16011 16809 16041
rect 16761 15999 16800 16011
rect 3381 15951 3459 15969
rect 5961 15951 6159 15969
rect 7161 15951 7539 15969
rect 9621 15951 9819 15969
rect 9981 15951 10119 15969
rect 14121 15951 14319 15969
rect 7701 15891 7899 15909
rect -189 15606 90 15654
rect -189 14094 -9 15606
rect 12501 15531 12579 15549
rect 11991 15291 12159 15309
rect 5040 15249 5079 15261
rect 5031 15219 5079 15249
rect 7341 15249 7380 15261
rect 7341 15219 7389 15249
rect 7821 15231 7929 15249
rect 5031 15141 5049 15219
rect 7371 15141 7389 15219
rect 7911 15141 7929 15231
rect 9621 15231 9699 15249
rect 10581 15231 10659 15249
rect 11001 15249 11040 15261
rect 11001 15219 11049 15249
rect 11031 15141 11049 15219
rect 11991 15141 12009 15291
rect 15171 15291 15339 15309
rect 12540 15249 12579 15261
rect 3501 15111 3579 15129
rect 5031 15111 5079 15141
rect 5040 15099 5079 15111
rect 7371 15111 7419 15141
rect 7380 15099 7419 15111
rect 7911 15111 7959 15141
rect 7920 15099 7959 15111
rect 8241 15111 8319 15129
rect 11001 15111 11049 15141
rect 11001 15099 11040 15111
rect 11961 15111 12009 15141
rect 12531 15219 12579 15249
rect 13920 15249 13959 15261
rect 13911 15219 13959 15249
rect 14301 15249 14340 15261
rect 14301 15219 14349 15249
rect 12531 15141 12549 15219
rect 13911 15141 13929 15219
rect 14331 15141 14349 15219
rect 15171 15141 15189 15291
rect 15621 15249 15660 15261
rect 16140 15249 16179 15261
rect 15621 15219 15669 15249
rect 12531 15111 12579 15141
rect 11961 15099 12000 15111
rect 12540 15099 12579 15111
rect 13911 15111 13959 15141
rect 13920 15099 13959 15111
rect 14331 15111 14379 15141
rect 14340 15099 14379 15111
rect 15141 15111 15189 15141
rect 15141 15099 15180 15111
rect 4221 15051 4659 15069
rect 9681 15051 9759 15069
rect 15651 15069 15669 15219
rect 16131 15219 16179 15249
rect 16131 15129 16149 15219
rect 16041 15111 16149 15129
rect 15651 15051 15759 15069
rect 18429 14874 18609 16386
rect 18330 14826 18609 14874
rect 17181 14751 17259 14769
rect 6321 14631 6399 14649
rect 7881 14631 8019 14649
rect 12231 14631 12459 14649
rect 8241 14589 8280 14601
rect 8400 14589 8439 14601
rect 8241 14559 8289 14589
rect 8271 14481 8289 14559
rect 7731 14451 7839 14469
rect 8241 14451 8289 14481
rect 8391 14559 8439 14589
rect 10080 14589 10119 14601
rect 9201 14571 9309 14589
rect 8241 14439 8280 14451
rect 2781 14391 3039 14409
rect 6861 14391 6999 14409
rect 8391 14418 8409 14559
rect 9291 14469 9309 14571
rect 10071 14559 10119 14589
rect 10821 14589 10860 14601
rect 10821 14559 10869 14589
rect 9291 14451 9369 14469
rect 9351 14421 9369 14451
rect 9351 14391 9399 14421
rect 9360 14379 9399 14391
rect 10071 14409 10089 14559
rect 10851 14481 10869 14559
rect 10821 14451 10869 14481
rect 12231 14481 12249 14631
rect 13941 14631 14079 14649
rect 15831 14631 15999 14649
rect 13041 14589 13080 14601
rect 13560 14589 13599 14601
rect 13041 14559 13089 14589
rect 13071 14481 13089 14559
rect 13551 14559 13599 14589
rect 13980 14589 14019 14601
rect 13971 14559 14019 14589
rect 14481 14589 14520 14601
rect 14481 14559 14529 14589
rect 15420 14589 15459 14601
rect 14781 14571 14889 14589
rect 13551 14481 13569 14559
rect 13971 14481 13989 14559
rect 14511 14481 14529 14559
rect 12231 14451 12279 14481
rect 10821 14439 10860 14451
rect 12240 14439 12279 14451
rect 13041 14451 13089 14481
rect 13041 14439 13080 14451
rect 13521 14451 13569 14481
rect 13521 14439 13560 14451
rect 13941 14451 13989 14481
rect 13941 14439 13980 14451
rect 14481 14451 14529 14481
rect 14871 14481 14889 14571
rect 15411 14559 15459 14589
rect 15411 14481 15429 14559
rect 15831 14481 15849 14631
rect 16320 14589 16359 14601
rect 14871 14451 14919 14481
rect 14481 14439 14520 14451
rect 14880 14439 14919 14451
rect 15411 14451 15459 14481
rect 15420 14439 15459 14451
rect 15801 14451 15849 14481
rect 16311 14559 16359 14589
rect 17601 14571 17829 14589
rect 16311 14481 16329 14559
rect 18180 14529 18219 14541
rect 18138 14511 18219 14529
rect 18180 14499 18219 14511
rect 16311 14451 16359 14481
rect 15801 14439 15840 14451
rect 16320 14439 16359 14451
rect 17601 14451 17679 14469
rect 9981 14391 10089 14409
rect 15201 14391 15339 14409
rect 17061 14391 17259 14409
rect 13461 14271 13539 14289
rect -189 14046 90 14094
rect -189 12534 -9 14046
rect 15561 13971 15759 13989
rect 14001 13851 14199 13869
rect 1221 13731 1419 13749
rect 8700 13749 8739 13761
rect 8691 13719 8739 13749
rect 15120 13749 15159 13761
rect 15111 13719 15159 13749
rect 3921 13689 3960 13701
rect 3921 13659 3969 13689
rect 7341 13689 7380 13701
rect 8340 13689 8379 13701
rect 7341 13659 7389 13689
rect 2838 13611 2979 13629
rect 1839 13569 1881 13599
rect 3951 13581 3969 13659
rect 7371 13629 7389 13659
rect 8331 13659 8379 13689
rect 8691 13689 8709 13719
rect 8631 13671 8709 13689
rect 7800 13629 7839 13641
rect 7371 13611 7482 13629
rect 7791 13611 7839 13629
rect 7800 13599 7839 13611
rect 8331 13581 8349 13659
rect 1839 13560 1959 13569
rect 1851 13551 1959 13560
rect 2481 13569 2520 13581
rect 2481 13551 2529 13569
rect 3951 13551 3999 13581
rect 2481 13539 2520 13551
rect 3960 13539 3999 13551
rect 4281 13551 4359 13569
rect 8301 13551 8349 13581
rect 8631 13581 8649 13671
rect 14061 13689 14100 13701
rect 14061 13659 14109 13689
rect 10041 13629 10080 13641
rect 10440 13629 10479 13641
rect 10041 13611 10089 13629
rect 10398 13611 10479 13629
rect 10041 13599 10080 13611
rect 10440 13599 10479 13611
rect 8631 13551 8679 13581
rect 8301 13539 8340 13551
rect 8640 13539 8679 13551
rect 10551 13521 10569 13659
rect 14091 13581 14109 13659
rect 14241 13629 14280 13641
rect 14241 13611 14289 13629
rect 14598 13611 14709 13629
rect 14241 13599 14280 13611
rect 14061 13551 14109 13581
rect 14691 13581 14709 13611
rect 15111 13581 15129 13719
rect 15180 13689 15219 13701
rect 14691 13551 14739 13581
rect 14061 13539 14100 13551
rect 14700 13539 14739 13551
rect 15081 13551 15129 13581
rect 15171 13659 15219 13689
rect 16461 13671 16569 13689
rect 15171 13581 15189 13659
rect 15171 13551 15219 13581
rect 15081 13539 15120 13551
rect 15180 13539 15219 13551
rect 16551 13569 16569 13671
rect 16941 13671 17109 13689
rect 17091 13629 17109 13671
rect 17091 13611 17202 13629
rect 17991 13581 18009 13719
rect 16551 13551 16629 13569
rect 17511 13551 17679 13569
rect 5121 13491 5319 13509
rect 6021 13491 6159 13509
rect 10521 13491 10569 13521
rect 16611 13521 16629 13551
rect 17961 13551 18009 13581
rect 17961 13539 18000 13551
rect 16611 13491 16659 13521
rect 10521 13479 10560 13491
rect 16620 13479 16659 13491
rect 18429 13314 18609 14826
rect 18330 13266 18609 13314
rect 3741 13191 3819 13209
rect 1341 13029 1380 13041
rect 1341 12999 1389 13029
rect 7401 13029 7440 13041
rect 7401 12999 7449 13029
rect 7911 13011 8019 13029
rect 13191 13011 13299 13029
rect 1371 12909 1389 12999
rect 4680 12969 4719 12981
rect 4671 12951 4719 12969
rect 4680 12939 4719 12951
rect 1371 12891 1449 12909
rect 2751 12891 2859 12909
rect 1431 12861 1449 12891
rect 4320 12918 4380 12921
rect 4341 12909 4380 12918
rect 7431 12909 7449 12999
rect 7521 12969 7560 12981
rect 7521 12951 7602 12969
rect 7521 12939 7560 12951
rect 13191 12909 13209 13011
rect 13791 13029 13809 13119
rect 14061 13071 14319 13089
rect 15681 13071 15879 13089
rect 13701 13011 13809 13029
rect 14181 13011 14289 13029
rect 4341 12891 4389 12909
rect 7431 12891 7509 12909
rect 13071 12891 13209 12909
rect 14271 12921 14289 13011
rect 14931 13011 15039 13029
rect 14931 12921 14949 13011
rect 15381 13011 15489 13029
rect 14271 12891 14319 12921
rect 4341 12879 4380 12891
rect 1431 12831 1479 12861
rect 1440 12819 1479 12831
rect 4311 12849 4329 12876
rect 7491 12861 7509 12891
rect 14280 12879 14319 12891
rect 14901 12891 14949 12921
rect 15471 12921 15489 13011
rect 16101 13029 16140 13041
rect 16101 12999 16149 13029
rect 16581 13011 16659 13029
rect 17100 13029 17139 13041
rect 17091 12999 17139 13029
rect 17481 13029 17520 13041
rect 17481 12999 17529 13029
rect 16131 12921 16149 12999
rect 15471 12891 15519 12921
rect 14901 12879 14940 12891
rect 15480 12879 15519 12891
rect 16101 12891 16149 12921
rect 17091 12909 17109 12999
rect 17511 12909 17529 12999
rect 17091 12891 17169 12909
rect 16101 12879 16140 12891
rect 17151 12861 17169 12891
rect 17451 12891 17529 12909
rect 17451 12861 17469 12891
rect 4101 12831 4329 12849
rect 6081 12831 6339 12849
rect 7491 12831 7539 12861
rect 7500 12819 7539 12831
rect 13581 12831 13779 12849
rect 14001 12831 14259 12849
rect 17151 12831 17199 12861
rect 17160 12819 17199 12831
rect 17421 12831 17469 12861
rect 17421 12819 17460 12831
rect -189 12486 90 12534
rect -189 10974 -9 12486
rect 8001 12279 8019 12321
rect 621 12171 819 12189
rect 5361 12171 5559 12189
rect 5901 12171 6039 12189
rect 7101 12171 7179 12189
rect 12261 12171 12459 12189
rect 12981 12171 13239 12189
rect 15621 12171 15879 12189
rect 17121 12171 17259 12189
rect 17781 12171 17979 12189
rect 18051 12171 18219 12189
rect 2640 12129 2679 12141
rect 2631 12111 2679 12129
rect 2640 12099 2679 12111
rect 4740 12129 4779 12141
rect 4731 12099 4779 12129
rect 5001 12129 5040 12141
rect 5580 12129 5619 12141
rect 5001 12099 5049 12129
rect 3240 12069 3279 12081
rect 3198 12051 3279 12069
rect 3240 12039 3279 12051
rect 4731 12021 4749 12099
rect 1401 11991 1539 12009
rect 4731 11991 4779 12021
rect 4740 11979 4779 11991
rect 5031 12009 5049 12099
rect 5571 12099 5619 12129
rect 5940 12129 5979 12141
rect 5931 12099 5979 12129
rect 6291 12111 6399 12129
rect 5571 12021 5589 12099
rect 5031 11991 5199 12009
rect 5541 11991 5589 12021
rect 5541 11979 5580 11991
rect 5931 11961 5949 12099
rect 6291 12021 6309 12111
rect 8361 12129 8400 12141
rect 8820 12129 8859 12141
rect 8361 12099 8409 12129
rect 8391 12021 8409 12099
rect 6261 11991 6309 12021
rect 6261 11979 6300 11991
rect 8361 11991 8409 12021
rect 8811 12099 8859 12129
rect 12741 12129 12780 12141
rect 12741 12099 12789 12129
rect 13881 12129 13920 12141
rect 15300 12129 15339 12141
rect 13881 12099 13929 12129
rect 8811 12021 8829 12099
rect 8811 11991 8859 12021
rect 8361 11979 8400 11991
rect 8820 11979 8859 11991
rect 12771 11961 12789 12099
rect 5901 11931 5949 11961
rect 5901 11919 5940 11931
rect 7041 11931 7119 11949
rect 13521 11931 13659 11949
rect 13911 11898 13929 12099
rect 15291 12099 15339 12129
rect 16221 12129 16260 12141
rect 18051 12129 18069 12171
rect 16221 12099 16281 12129
rect 15291 12069 15309 12099
rect 16239 12081 16281 12099
rect 17991 12111 18069 12129
rect 16620 12069 16659 12081
rect 15138 12051 15309 12069
rect 16578 12051 16659 12069
rect 15291 12021 15309 12051
rect 16620 12039 16659 12051
rect 17991 12021 18009 12111
rect 14781 12009 14820 12021
rect 14781 11991 14829 12009
rect 15291 11991 15339 12021
rect 14781 11979 14820 11991
rect 15300 11979 15339 11991
rect 16041 11991 16269 12009
rect 17991 11991 18039 12021
rect 18000 11979 18039 11991
rect 18429 11754 18609 13266
rect 18330 11706 18609 11754
rect 7881 11631 7959 11649
rect 7941 11571 8139 11589
rect 17061 11571 17139 11589
rect 4521 11511 4629 11529
rect 2280 11469 2319 11481
rect 2271 11439 2319 11469
rect 2601 11451 2679 11469
rect 3660 11469 3699 11481
rect 3651 11439 3699 11469
rect 2271 11361 2289 11439
rect 3651 11361 3669 11439
rect 4071 11361 4089 11439
rect 4611 11361 4629 11511
rect 5760 11529 5799 11541
rect 4881 11511 4989 11529
rect 4971 11361 4989 11511
rect 5751 11499 5799 11529
rect 14901 11511 14979 11529
rect 15021 11511 15099 11529
rect 17421 11511 17619 11529
rect 5751 11361 5769 11499
rect 5820 11469 5859 11481
rect 2271 11331 2319 11361
rect 2280 11319 2319 11331
rect 3651 11331 3699 11361
rect 3660 11319 3699 11331
rect 4071 11331 4119 11361
rect 4080 11319 4119 11331
rect 4611 11331 4659 11361
rect 4620 11319 4659 11331
rect 4941 11331 4989 11361
rect 4941 11319 4980 11331
rect 5721 11331 5769 11361
rect 5811 11439 5859 11469
rect 6231 11451 6399 11469
rect 5811 11361 5829 11439
rect 6231 11361 6249 11451
rect 8400 11469 8439 11481
rect 8391 11439 8439 11469
rect 11961 11469 12000 11481
rect 11961 11439 12009 11469
rect 17061 11451 17169 11469
rect 5811 11331 5859 11361
rect 5721 11319 5760 11331
rect 5820 11319 5859 11331
rect 6201 11331 6249 11361
rect 6201 11319 6240 11331
rect 2781 11271 2919 11289
rect 5181 11271 5259 11289
rect 6261 11271 6399 11289
rect 8391 11298 8409 11439
rect 11991 11358 12009 11439
rect 17151 11361 17169 11451
rect 17481 11469 17520 11481
rect 17481 11439 17529 11469
rect 17841 11469 17880 11481
rect 17841 11439 17889 11469
rect 17511 11361 17529 11439
rect 17871 11361 17889 11439
rect 17151 11331 17199 11361
rect 17160 11319 17199 11331
rect 17511 11331 17559 11361
rect 17520 11319 17559 11331
rect 17841 11331 17889 11361
rect 17841 11319 17880 11331
rect 9201 11271 9399 11289
rect 16881 11271 17259 11289
rect 17421 11271 17619 11289
rect -189 10926 90 10974
rect -189 9414 -9 10926
rect 8061 10851 8139 10869
rect 5601 10731 5799 10749
rect 4701 10671 4959 10689
rect 201 10611 399 10629
rect 1521 10611 1779 10629
rect 5751 10611 5859 10629
rect 4860 10569 4899 10581
rect 4851 10539 4899 10569
rect 5751 10569 5769 10611
rect 8421 10611 8559 10629
rect 16461 10611 16599 10629
rect 16971 10611 17139 10629
rect 6120 10569 6159 10581
rect 5691 10560 5769 10569
rect 5679 10551 5769 10560
rect 4851 10461 4869 10539
rect 5679 10518 5721 10551
rect 6111 10539 6159 10569
rect 11361 10551 11439 10569
rect 13380 10569 13419 10581
rect 13371 10539 13419 10569
rect 15960 10569 15999 10581
rect 15951 10539 15999 10569
rect 6111 10461 6129 10539
rect 13371 10461 13389 10539
rect 4851 10431 4899 10461
rect 4860 10419 4899 10431
rect 6111 10431 6159 10461
rect 6120 10419 6159 10431
rect 13341 10431 13389 10461
rect 15951 10461 15969 10539
rect 16971 10461 16989 10611
rect 17931 10551 18039 10569
rect 17931 10461 17949 10551
rect 15951 10431 15999 10461
rect 13341 10419 13380 10431
rect 15960 10419 15999 10431
rect 16941 10431 16989 10461
rect 16941 10419 16980 10431
rect 17901 10431 17949 10461
rect 17901 10419 17940 10431
rect 6801 10371 7059 10389
rect 18429 10194 18609 11706
rect 18330 10146 18609 10194
rect 7521 10071 7659 10089
rect 9111 9981 9129 10059
rect 7080 9969 7119 9981
rect 7071 9939 7119 9969
rect 1821 9909 1860 9921
rect 1920 9909 1959 9921
rect 1821 9879 1869 9909
rect 1851 9801 1869 9879
rect 1821 9771 1869 9801
rect 1911 9879 1959 9909
rect 2301 9909 2340 9921
rect 4620 9909 4659 9921
rect 2301 9879 2349 9909
rect 1821 9759 1860 9771
rect 1911 9741 1929 9879
rect 2331 9801 2349 9879
rect 2301 9771 2349 9801
rect 4611 9879 4659 9909
rect 4881 9909 4920 9921
rect 4881 9879 4929 9909
rect 5841 9909 5880 9921
rect 5841 9879 5889 9909
rect 4611 9801 4629 9879
rect 4611 9771 4659 9801
rect 2301 9759 2340 9771
rect 4620 9759 4659 9771
rect 1401 9711 1539 9729
rect 3621 9711 3819 9729
rect 4911 9729 4929 9879
rect 5871 9801 5889 9879
rect 5841 9771 5889 9801
rect 7071 9789 7089 9939
rect 7140 9909 7179 9921
rect 7011 9771 7089 9789
rect 7131 9879 7179 9909
rect 7941 9909 7980 9921
rect 7941 9879 7989 9909
rect 8661 9909 8700 9921
rect 10080 9909 10119 9921
rect 8661 9879 8709 9909
rect 7131 9801 7149 9879
rect 7971 9801 7989 9879
rect 8691 9849 8709 9879
rect 10071 9879 10119 9909
rect 12201 9909 12240 9921
rect 12201 9879 12249 9909
rect 8691 9831 8769 9849
rect 7131 9771 7179 9801
rect 5841 9759 5880 9771
rect 7011 9741 7029 9771
rect 7140 9759 7179 9771
rect 7941 9771 7989 9801
rect 8751 9801 8769 9831
rect 10071 9801 10089 9879
rect 12231 9801 12249 9879
rect 14511 9891 14619 9909
rect 14511 9801 14529 9891
rect 8751 9771 8799 9801
rect 7941 9759 7980 9771
rect 8760 9759 8799 9771
rect 10071 9771 10119 9801
rect 10080 9759 10119 9771
rect 12201 9771 12249 9801
rect 13200 9789 13239 9801
rect 12201 9759 12240 9771
rect 13191 9759 13239 9789
rect 14481 9771 14529 9801
rect 14481 9759 14520 9771
rect 15471 9789 15489 9939
rect 16641 9909 16680 9921
rect 16641 9879 16689 9909
rect 16671 9801 16689 9879
rect 17901 9891 18009 9909
rect 15321 9771 15489 9789
rect 16641 9771 16689 9801
rect 17991 9789 18009 9891
rect 17991 9771 18069 9789
rect 16641 9759 16680 9771
rect 4911 9711 5079 9729
rect 7041 9711 7239 9729
rect 7521 9711 7659 9729
rect 11661 9711 11979 9729
rect 13191 9678 13209 9759
rect 13281 9711 13359 9729
rect 14841 9711 15039 9729
rect 18051 9729 18069 9771
rect 18051 9720 18129 9729
rect 18051 9711 18141 9720
rect 18099 9678 18141 9711
rect 16941 9591 17019 9609
rect -189 9366 90 9414
rect -189 7854 -9 9366
rect 6321 9291 6459 9309
rect 861 9051 1179 9069
rect 5001 9051 5139 9069
rect 5841 9051 6099 9069
rect 8181 9051 8259 9069
rect 8481 9051 8679 9069
rect 3261 9009 3300 9021
rect 3261 8979 3309 9009
rect 3291 8901 3309 8979
rect 4071 8991 4239 9009
rect 4071 8901 4089 8991
rect 5481 8991 5559 9009
rect 5901 9009 5940 9021
rect 6480 9009 6519 9021
rect 5901 8979 5949 9009
rect 2421 8871 2559 8889
rect 3261 8871 3309 8901
rect 3261 8859 3300 8871
rect 4041 8871 4089 8901
rect 4041 8859 4080 8871
rect 5931 8841 5949 8979
rect 6471 8979 6519 9009
rect 7680 9009 7719 9021
rect 7671 8979 7719 9009
rect 9120 9009 9159 9021
rect 9111 8979 9159 9009
rect 9480 9009 9519 9021
rect 9471 8979 9519 9009
rect 9861 9009 9900 9021
rect 12000 9009 12039 9021
rect 9861 8979 9909 9009
rect 6471 8901 6489 8979
rect 6471 8871 6519 8901
rect 6480 8859 6519 8871
rect 6741 8811 6999 8829
rect 7671 8829 7689 8979
rect 7671 8811 7779 8829
rect 9111 8838 9129 8979
rect 9471 8901 9489 8979
rect 9891 8901 9909 8979
rect 9471 8871 9519 8901
rect 9480 8859 9519 8871
rect 9861 8871 9909 8901
rect 11991 8979 12039 9009
rect 12321 8991 12489 9009
rect 11991 8901 12009 8979
rect 12471 8901 12489 8991
rect 12861 9009 12900 9021
rect 15960 9009 15999 9021
rect 12861 8979 12909 9009
rect 12891 8901 12909 8979
rect 15951 8979 15999 9009
rect 16920 9009 16959 9021
rect 16911 8979 16959 9009
rect 15951 8901 15969 8979
rect 11991 8871 12039 8901
rect 9861 8859 9900 8871
rect 12000 8859 12039 8871
rect 12471 8871 12519 8901
rect 12480 8859 12519 8871
rect 12891 8871 12939 8901
rect 12900 8859 12939 8871
rect 14841 8871 14919 8889
rect 15951 8871 15999 8901
rect 15960 8859 15999 8871
rect 16911 8889 16929 8979
rect 16821 8871 16929 8889
rect 15501 8811 15639 8829
rect 17481 8751 17619 8769
rect 18429 8634 18609 10146
rect 18330 8586 18609 8634
rect 4941 8451 5139 8469
rect 16611 8421 16629 8499
rect 17019 8481 17061 8499
rect 17001 8460 17061 8481
rect 17001 8451 17049 8460
rect 17001 8439 17040 8451
rect 4461 8391 4539 8409
rect 4611 8391 4779 8409
rect 2880 8349 2919 8361
rect 2871 8319 2919 8349
rect 2871 8241 2889 8319
rect 2871 8211 2919 8241
rect 2880 8199 2919 8211
rect 1281 8151 1599 8169
rect 2661 8151 2859 8169
rect 4611 8178 4629 8391
rect 5781 8391 5979 8409
rect 7401 8391 7599 8409
rect 16101 8391 16299 8409
rect 16581 8391 16629 8421
rect 16581 8379 16620 8391
rect 4971 8331 5139 8349
rect 4971 8241 4989 8331
rect 6300 8349 6339 8361
rect 6291 8340 6339 8349
rect 6279 8319 6339 8340
rect 6720 8349 6759 8361
rect 6711 8319 6759 8349
rect 7431 8331 7539 8349
rect 6279 8298 6321 8319
rect 4941 8211 4989 8241
rect 6711 8241 6729 8319
rect 7431 8241 7449 8331
rect 8340 8349 8379 8361
rect 8331 8319 8379 8349
rect 9141 8349 9180 8361
rect 9840 8349 9879 8361
rect 9141 8319 9189 8349
rect 7779 8241 7821 8259
rect 8331 8241 8349 8319
rect 9171 8241 9189 8319
rect 9831 8319 9879 8349
rect 15300 8349 15339 8361
rect 15291 8319 15339 8349
rect 15681 8349 15720 8361
rect 15681 8319 15729 8349
rect 16041 8349 16080 8361
rect 16041 8319 16089 8349
rect 16131 8340 16239 8349
rect 9321 8289 9360 8301
rect 9720 8289 9759 8301
rect 9321 8271 9402 8289
rect 9711 8271 9759 8289
rect 9321 8259 9360 8271
rect 9720 8259 9759 8271
rect 6711 8211 6759 8241
rect 4941 8199 4980 8211
rect 6720 8199 6759 8211
rect 7401 8211 7449 8241
rect 7401 8199 7440 8211
rect 7761 8220 7821 8241
rect 7761 8211 7809 8220
rect 7761 8199 7800 8211
rect 8301 8211 8349 8241
rect 8301 8199 8340 8211
rect 9141 8211 9189 8241
rect 9831 8241 9849 8319
rect 15291 8301 15309 8319
rect 15240 8298 15309 8301
rect 15261 8271 15309 8298
rect 15261 8259 15300 8271
rect 15711 8241 15729 8319
rect 16071 8241 16089 8319
rect 16119 8331 16239 8340
rect 16119 8301 16161 8331
rect 16671 8241 16689 8439
rect 17301 8391 17439 8409
rect 17721 8391 17829 8409
rect 16980 8349 17019 8361
rect 9831 8211 9879 8241
rect 9141 8199 9180 8211
rect 9840 8199 9879 8211
rect 15321 8229 15360 8241
rect 15321 8220 15369 8229
rect 15321 8199 15381 8220
rect 15711 8211 15759 8241
rect 15720 8199 15759 8211
rect 16041 8211 16089 8241
rect 16041 8199 16080 8211
rect 16641 8211 16689 8241
rect 16971 8319 17019 8349
rect 17421 8349 17460 8361
rect 17421 8319 17469 8349
rect 16971 8241 16989 8319
rect 17451 8241 17469 8319
rect 17811 8241 17829 8391
rect 16971 8211 17019 8241
rect 16641 8199 16680 8211
rect 16980 8199 17019 8211
rect 17421 8211 17469 8241
rect 17421 8199 17460 8211
rect 17781 8211 17829 8241
rect 17781 8199 17820 8211
rect 15339 8181 15381 8199
rect 6561 8151 6639 8169
rect 7461 8151 7599 8169
rect 7881 8151 7959 8169
rect 15981 8151 16119 8169
rect 2841 8031 2919 8049
rect -189 7806 90 7854
rect -189 6294 -9 7806
rect 5901 7611 6099 7629
rect 3321 7551 3519 7569
rect 4101 7491 4299 7509
rect 5943 7491 6159 7509
rect 8121 7491 8559 7509
rect 11001 7491 11199 7509
rect 13161 7491 13269 7509
rect 501 7449 540 7461
rect 3060 7449 3099 7461
rect 501 7419 549 7449
rect 531 7341 549 7419
rect 3051 7419 3099 7449
rect 3681 7449 3720 7461
rect 3681 7440 3729 7449
rect 3681 7419 3741 7440
rect 8280 7449 8319 7461
rect 7281 7431 7389 7449
rect 531 7311 579 7341
rect 540 7299 579 7311
rect 3051 7269 3069 7419
rect 3699 7398 3741 7419
rect 3771 7341 3789 7419
rect 7371 7341 7389 7431
rect 8271 7419 8319 7449
rect 8781 7449 8820 7461
rect 8781 7419 8829 7449
rect 9321 7449 9360 7461
rect 9321 7419 9369 7449
rect 10101 7449 10140 7461
rect 10101 7419 10149 7449
rect 3771 7311 3819 7341
rect 3780 7299 3819 7311
rect 7371 7311 7419 7341
rect 7380 7299 7419 7311
rect 8271 7329 8289 7419
rect 8811 7341 8829 7419
rect 8181 7311 8289 7329
rect 8781 7311 8829 7341
rect 9351 7341 9369 7419
rect 10131 7341 10149 7419
rect 13251 7341 13269 7491
rect 17931 7491 18039 7509
rect 14061 7449 14100 7461
rect 14061 7419 14109 7449
rect 14481 7449 14520 7461
rect 14481 7419 14529 7449
rect 15321 7449 15360 7461
rect 15321 7419 15369 7449
rect 17061 7449 17100 7461
rect 17061 7419 17109 7449
rect 9351 7311 9399 7341
rect 8781 7299 8820 7311
rect 9360 7299 9399 7311
rect 10131 7311 10179 7341
rect 10140 7299 10179 7311
rect 13221 7311 13269 7341
rect 14091 7329 14109 7419
rect 14511 7341 14529 7419
rect 14091 7311 14199 7329
rect 13221 7299 13260 7311
rect 14481 7311 14529 7341
rect 15351 7341 15369 7419
rect 17091 7341 17109 7419
rect 17511 7431 17619 7449
rect 17511 7341 17529 7431
rect 17931 7341 17949 7491
rect 15351 7311 15399 7341
rect 14481 7299 14520 7311
rect 15360 7299 15399 7311
rect 17091 7311 17139 7341
rect 17100 7299 17139 7311
rect 17481 7311 17529 7341
rect 17481 7299 17520 7311
rect 17901 7311 17949 7341
rect 17901 7299 17940 7311
rect 2961 7251 3069 7269
rect 8181 7251 8439 7269
rect 18429 7074 18609 8586
rect 18330 7026 18609 7074
rect 15261 6951 15339 6969
rect 5061 6891 5199 6909
rect 7221 6831 7359 6849
rect 180 6789 219 6801
rect 171 6759 219 6789
rect 1521 6789 1560 6801
rect 3360 6789 3399 6801
rect 1521 6759 1569 6789
rect 171 6669 189 6759
rect 600 6729 639 6741
rect 591 6699 639 6729
rect 591 6681 609 6699
rect 171 6651 249 6669
rect 231 6621 249 6651
rect 561 6651 609 6681
rect 1551 6681 1569 6759
rect 3351 6759 3399 6789
rect 5121 6789 5160 6801
rect 5121 6759 5169 6789
rect 6120 6789 6159 6801
rect 6111 6759 6159 6789
rect 1551 6651 1599 6681
rect 561 6639 600 6651
rect 1560 6639 1599 6651
rect 2541 6651 2619 6669
rect 3351 6669 3369 6759
rect 5151 6681 5169 6759
rect 3291 6651 3369 6669
rect 231 6615 300 6621
rect 231 6591 279 6615
rect 240 6579 279 6591
rect 3291 6609 3309 6651
rect 4701 6651 4839 6669
rect 5151 6651 5199 6681
rect 5160 6639 5199 6651
rect 5631 6669 5649 6759
rect 5571 6651 5649 6669
rect 6111 6681 6129 6759
rect 6531 6681 6549 6819
rect 7161 6789 7200 6801
rect 7161 6759 7209 6789
rect 8121 6789 8160 6801
rect 8121 6759 8169 6789
rect 9681 6789 9720 6801
rect 9681 6759 9729 6789
rect 12081 6789 12120 6801
rect 12180 6789 12219 6801
rect 12081 6759 12129 6789
rect 6111 6651 6159 6681
rect 3141 6591 3309 6609
rect 5571 6609 5589 6651
rect 6120 6639 6159 6651
rect 6531 6651 6579 6681
rect 6540 6639 6579 6651
rect 7191 6669 7209 6759
rect 8151 6678 8169 6759
rect 9711 6681 9729 6759
rect 7191 6651 7299 6669
rect 9681 6651 9729 6681
rect 11631 6669 11649 6759
rect 12111 6681 12129 6759
rect 11631 6651 11709 6669
rect 9681 6639 9720 6651
rect 5481 6591 5679 6609
rect 11691 6609 11709 6651
rect 12081 6651 12129 6681
rect 12171 6759 12219 6789
rect 14601 6771 14679 6789
rect 15201 6771 15369 6789
rect 12171 6681 12189 6759
rect 15351 6681 15369 6771
rect 12171 6651 12219 6681
rect 12081 6639 12120 6651
rect 12180 6639 12219 6651
rect 15351 6651 15399 6681
rect 15360 6639 15399 6651
rect 11691 6591 11799 6609
rect 16041 6531 16239 6549
rect 5961 6471 6219 6489
rect -189 6246 90 6294
rect -189 4734 -9 6246
rect 4761 6051 4959 6069
rect 6501 6051 6639 6069
rect 13461 6051 13599 6069
rect 7461 5991 7539 6009
rect 10281 5991 10359 6009
rect 17121 5991 17319 6009
rect 1941 5931 2019 5949
rect 2661 5949 2700 5961
rect 2661 5919 2709 5949
rect 3141 5931 3219 5949
rect 5541 5931 5799 5949
rect 6861 5931 6999 5949
rect 7341 5931 7539 5949
rect 2691 5889 2709 5919
rect 12561 5931 12699 5949
rect 13761 5931 13869 5949
rect 5220 5889 5259 5901
rect 2691 5871 2769 5889
rect 2751 5781 2769 5871
rect 5211 5859 5259 5889
rect 6021 5889 6060 5901
rect 6021 5859 6069 5889
rect 8241 5889 8280 5901
rect 8340 5889 8379 5901
rect 8241 5859 8289 5889
rect 5211 5781 5229 5859
rect 6051 5781 6069 5859
rect 2721 5751 2769 5781
rect 2721 5739 2760 5751
rect 5181 5751 5229 5781
rect 5181 5739 5220 5751
rect 6021 5751 6069 5781
rect 6021 5739 6060 5751
rect 8271 5721 8289 5859
rect 8331 5859 8379 5889
rect 12981 5889 13020 5901
rect 12981 5859 13029 5889
rect 8331 5781 8349 5859
rect 8331 5751 8379 5781
rect 8340 5739 8379 5751
rect 13011 5778 13029 5859
rect 13851 5781 13869 5931
rect 15831 5931 15939 5949
rect 15831 5889 15849 5931
rect 16701 5931 16899 5949
rect 17121 5931 17259 5949
rect 13821 5751 13869 5781
rect 15771 5871 15849 5889
rect 13821 5739 13860 5751
rect 8271 5691 8319 5721
rect 8280 5679 8319 5691
rect 8931 5700 9099 5709
rect 8919 5691 9099 5700
rect 8919 5661 8961 5691
rect 13521 5691 13599 5709
rect 15771 5709 15789 5871
rect 16161 5889 16200 5901
rect 16800 5889 16839 5901
rect 16161 5859 16209 5889
rect 16191 5781 16209 5859
rect 16161 5751 16209 5781
rect 16791 5859 16839 5889
rect 17601 5871 17709 5889
rect 16791 5769 16809 5859
rect 17691 5781 17709 5871
rect 16791 5760 16869 5769
rect 16791 5751 16881 5760
rect 17691 5751 17739 5781
rect 16161 5739 16200 5751
rect 16839 5721 16881 5751
rect 17700 5739 17739 5751
rect 15771 5691 15939 5709
rect 17181 5691 17319 5709
rect 18429 5514 18609 7026
rect 18330 5466 18609 5514
rect 16101 5331 16179 5349
rect 561 5229 600 5241
rect 561 5199 609 5229
rect 1041 5211 1119 5229
rect 591 5121 609 5199
rect 4851 5121 4869 5319
rect 10761 5271 10959 5289
rect 5811 5211 5919 5229
rect 5271 5121 5289 5199
rect 591 5091 639 5121
rect 600 5079 639 5091
rect 4851 5091 4899 5121
rect 4860 5079 4899 5091
rect 5241 5091 5289 5121
rect 5811 5109 5829 5211
rect 6300 5229 6339 5241
rect 6291 5199 6339 5229
rect 6720 5229 6759 5241
rect 6711 5199 6759 5229
rect 10479 5229 10521 5259
rect 15741 5271 15819 5289
rect 11340 5229 11379 5241
rect 10431 5220 10521 5229
rect 10431 5211 10509 5220
rect 6291 5121 6309 5199
rect 5751 5091 5829 5109
rect 5241 5079 5280 5091
rect 5751 5049 5769 5091
rect 6261 5091 6309 5121
rect 6711 5121 6729 5199
rect 10431 5121 10449 5211
rect 11331 5199 11379 5229
rect 12420 5229 12459 5241
rect 12411 5199 12459 5229
rect 13641 5229 13680 5241
rect 13641 5199 13689 5229
rect 15681 5199 15729 5235
rect 11331 5121 11349 5199
rect 12411 5121 12429 5199
rect 6711 5091 6759 5121
rect 6261 5079 6300 5091
rect 6720 5079 6759 5091
rect 10431 5091 10479 5121
rect 10440 5079 10479 5091
rect 11331 5091 11379 5121
rect 11340 5079 11379 5091
rect 12411 5091 12459 5121
rect 12420 5079 12459 5091
rect 5661 5031 5769 5049
rect 6201 5031 6399 5049
rect 8241 5031 8319 5049
rect 13341 5031 13419 5049
rect 13671 5049 13689 5199
rect 15711 5121 15729 5199
rect 16371 5211 16479 5229
rect 16371 5121 16389 5211
rect 15711 5091 15759 5121
rect 15720 5079 15759 5091
rect 16341 5091 16389 5121
rect 16341 5079 16380 5091
rect 13671 5031 13779 5049
rect 5061 4971 5319 4989
rect -189 4686 90 4734
rect -189 3174 -9 4686
rect 10341 4611 10479 4629
rect 5661 4431 5919 4449
rect 3441 4371 3699 4389
rect 4881 4371 4959 4389
rect 5241 4371 5439 4389
rect 12801 4371 13119 4389
rect 14241 4371 14379 4389
rect 18141 4371 18219 4389
rect 5880 4329 5919 4341
rect 5871 4299 5919 4329
rect 6621 4329 6660 4341
rect 8700 4329 8739 4341
rect 6621 4299 6669 4329
rect 5871 4221 5889 4299
rect 6651 4221 6669 4299
rect 1761 4191 1839 4209
rect 5871 4191 5919 4221
rect 5880 4179 5919 4191
rect 6621 4191 6669 4221
rect 8691 4299 8739 4329
rect 9861 4329 9900 4341
rect 9861 4299 9909 4329
rect 10281 4329 10320 4341
rect 10281 4299 10329 4329
rect 8691 4221 8709 4299
rect 8691 4191 8739 4221
rect 6621 4179 6660 4191
rect 8700 4179 8739 4191
rect 9891 4209 9909 4299
rect 10311 4221 10329 4299
rect 13851 4311 13959 4329
rect 13851 4221 13869 4311
rect 15621 4311 15729 4329
rect 9831 4200 9909 4209
rect 9819 4191 9909 4200
rect 9819 4161 9861 4191
rect 10281 4191 10329 4221
rect 10281 4179 10320 4191
rect 13821 4191 13869 4221
rect 15711 4221 15729 4311
rect 15981 4329 16020 4341
rect 15981 4299 16029 4329
rect 16011 4221 16029 4299
rect 15711 4191 15759 4221
rect 13821 4179 13860 4191
rect 15720 4179 15759 4191
rect 16011 4191 16059 4221
rect 16020 4179 16059 4191
rect 18201 4191 18339 4209
rect 4461 4131 4599 4149
rect 10341 4131 10479 4149
rect 17841 4071 17979 4089
rect 18429 3954 18609 5466
rect 18330 3906 18609 3954
rect 13341 3711 13419 3729
rect 6861 3669 6900 3681
rect 9060 3669 9099 3681
rect 6861 3639 6909 3669
rect 141 3609 180 3621
rect 141 3579 189 3609
rect 171 3561 189 3579
rect 171 3531 219 3561
rect 180 3519 219 3531
rect 6891 3549 6909 3639
rect 9051 3639 9099 3669
rect 10881 3669 10920 3681
rect 10881 3639 10929 3669
rect 11181 3669 11220 3681
rect 11280 3669 11319 3681
rect 11181 3639 11229 3669
rect 9051 3561 9069 3639
rect 10911 3561 10929 3639
rect 6891 3531 7059 3549
rect 9051 3531 9099 3561
rect 9060 3519 9099 3531
rect 10911 3531 10959 3561
rect 10920 3519 10959 3531
rect 1761 3471 1839 3489
rect 3621 3471 3699 3489
rect 11211 3489 11229 3639
rect 11271 3639 11319 3669
rect 16539 3669 16581 3699
rect 16491 3660 16581 3669
rect 16491 3651 16569 3660
rect 11271 3561 11289 3639
rect 11271 3531 11319 3561
rect 11280 3519 11319 3531
rect 16491 3549 16509 3651
rect 16401 3531 16509 3549
rect 11211 3471 11379 3489
rect 11721 3471 11859 3489
rect 15681 3471 15879 3489
rect 18231 3441 18249 3579
rect -189 3126 90 3174
rect -189 1614 -9 3126
rect 9501 3051 9579 3069
rect 6519 2889 6561 2919
rect 6381 2880 6561 2889
rect 6381 2871 6549 2880
rect 15201 2871 15279 2889
rect 381 2811 759 2829
rect 3081 2811 3219 2829
rect 3621 2811 3939 2829
rect 4521 2811 4659 2829
rect 7641 2811 7899 2829
rect 12543 2811 12639 2829
rect 12921 2811 13179 2829
rect 17001 2811 17079 2829
rect 4761 2751 4839 2769
rect 5961 2751 6039 2769
rect 12141 2769 12180 2781
rect 15240 2769 15279 2781
rect 12141 2739 12189 2769
rect 12171 2649 12189 2739
rect 15231 2739 15279 2769
rect 15660 2769 15699 2781
rect 15651 2739 15699 2769
rect 16401 2769 16440 2781
rect 16401 2739 16449 2769
rect 15231 2661 15249 2739
rect 15651 2661 15669 2739
rect 16431 2661 16449 2739
rect 12171 2640 12249 2649
rect 12171 2631 12261 2640
rect 15231 2631 15279 2661
rect 12219 2601 12261 2631
rect 15240 2619 15279 2631
rect 15621 2631 15669 2661
rect 15621 2619 15660 2631
rect 16401 2631 16449 2661
rect 16401 2619 16440 2631
rect 9861 2571 9999 2589
rect 18429 2394 18609 3906
rect 18330 2346 18609 2394
rect 5601 2151 5679 2169
rect 8961 2151 9159 2169
rect 11781 2151 11919 2169
rect 12801 2151 12999 2169
rect 14700 2169 14739 2181
rect 14691 2139 14739 2169
rect 3861 2109 3900 2121
rect 3861 2079 3909 2109
rect 5181 2109 5220 2121
rect 5181 2079 5229 2109
rect 3891 2001 3909 2079
rect 3891 1971 3939 2001
rect 3900 1959 3939 1971
rect 5211 1989 5229 2079
rect 6111 2091 6219 2109
rect 6111 2001 6129 2091
rect 6660 2109 6699 2121
rect 6651 2079 6699 2109
rect 8901 2091 9039 2109
rect 14691 2109 14709 2139
rect 17460 2109 17499 2121
rect 14631 2091 14709 2109
rect 6651 2049 6669 2079
rect 6591 2031 6669 2049
rect 6591 2001 6609 2031
rect 9459 2001 9501 2019
rect 9531 2001 9549 2079
rect 5211 1980 5349 1989
rect 5211 1971 5361 1980
rect 5319 1941 5361 1971
rect 6081 1971 6129 2001
rect 6081 1959 6120 1971
rect 6561 1971 6609 2001
rect 6561 1959 6600 1971
rect 9441 1980 9501 2001
rect 9441 1971 9489 1980
rect 9441 1959 9480 1971
rect 11181 1971 11259 1989
rect 11331 1941 11349 2019
rect 14631 2001 14649 2091
rect 17451 2079 17499 2109
rect 17451 2001 17469 2079
rect 14601 1971 14649 2001
rect 14601 1959 14640 1971
rect 17421 1971 17469 2001
rect 17421 1959 17460 1971
rect 4641 1911 5019 1929
rect 11541 1911 11859 1929
rect -189 1566 90 1614
rect -189 54 -9 1566
rect 1401 1251 1479 1269
rect 6381 1251 6819 1269
rect 8181 1251 8379 1269
rect 8421 1251 8619 1269
rect 17601 1251 17739 1269
rect 4551 1191 4779 1209
rect 6600 1209 6639 1221
rect 6591 1179 6639 1209
rect 9681 1209 9720 1221
rect 9780 1209 9819 1221
rect 9681 1179 9729 1209
rect 6591 1089 6609 1179
rect 9711 1101 9729 1179
rect 6531 1080 6609 1089
rect 6519 1071 6609 1080
rect 6519 1041 6561 1071
rect 9681 1071 9729 1101
rect 9771 1179 9819 1209
rect 9681 1059 9720 1071
rect 9771 1041 9789 1179
rect 2661 1011 2799 1029
rect 5121 1011 5379 1029
rect 9720 1038 9789 1041
rect 9741 1011 9789 1038
rect 9741 999 9780 1011
rect 10881 1011 11019 1029
rect 6081 951 6159 969
rect 5061 891 5259 909
rect 18429 834 18609 2346
rect 18330 786 18609 834
rect 4881 711 5019 729
rect 8541 591 8739 609
rect 4461 531 4599 549
rect 7620 549 7659 561
rect 7611 519 7659 549
rect 8901 549 8940 561
rect 8901 519 8949 549
rect 12441 549 12480 561
rect 13320 549 13359 561
rect 12441 519 12489 549
rect 7611 441 7629 519
rect 6321 411 6399 429
rect 7581 411 7629 441
rect 8931 441 8949 519
rect 12000 489 12039 501
rect 11991 471 12039 489
rect 12000 459 12039 471
rect 8931 411 8979 441
rect 7581 399 7620 411
rect 8940 399 8979 411
rect 12471 429 12489 519
rect 13311 519 13359 549
rect 13311 441 13329 519
rect 11541 411 11709 429
rect 12471 411 12549 429
rect 1761 351 2019 369
rect 3021 351 3279 369
rect 3498 339 3501 360
rect 3561 351 3759 369
rect 6261 351 6579 369
rect 12531 369 12549 411
rect 13281 411 13329 441
rect 13281 399 13320 411
rect 12531 351 12639 369
rect 17961 351 18219 369
rect 3459 309 3501 339
rect 3459 300 3699 309
rect 3471 291 3699 300
rect 8421 111 8499 129
rect -189 6 90 54
rect 18429 6 18609 786
<< m2contact >>
rect 6819 18402 6861 18444
rect 6999 18399 7041 18441
rect 7599 18399 7641 18441
rect 7959 18399 8001 18441
rect 11739 18399 11781 18441
rect 16779 18399 16821 18441
rect 17079 18399 17121 18441
rect 12039 18339 12081 18381
rect 17739 18339 17781 18381
rect 13719 18279 13761 18321
rect 11739 18219 11781 18261
rect 12159 18219 12201 18261
rect 14199 18219 14241 18261
rect 17739 18219 17781 18261
rect 15519 18159 15561 18201
rect 15759 18159 15801 18201
rect 8541 17799 8583 17841
rect 8679 17799 8721 17841
rect 6399 17739 6441 17781
rect 6579 17739 6621 17781
rect 8379 17739 8421 17781
rect 8559 17739 8601 17781
rect 12819 17739 12861 17781
rect 13059 17739 13101 17781
rect 579 17679 621 17721
rect 11139 17679 11181 17721
rect 15879 17679 15921 17721
rect 579 17559 621 17601
rect 8919 17559 8961 17601
rect 9039 17559 9081 17601
rect 11019 17556 11061 17598
rect 15879 17559 15921 17601
rect 16899 17679 16941 17721
rect 16899 17559 16941 17601
rect 7719 17499 7761 17541
rect 7959 17499 8001 17541
rect 12519 17499 12561 17541
rect 12699 17499 12741 17541
rect 16299 17499 16341 17541
rect 16539 17499 16581 17541
rect 1119 16839 1161 16881
rect 1299 16839 1341 16881
rect 6639 16839 6681 16881
rect 6759 16839 6801 16881
rect 6879 16839 6921 16881
rect 8979 16839 9021 16881
rect 9159 16839 9201 16881
rect 14619 16839 14661 16881
rect 14739 16842 14781 16884
rect 1539 16779 1581 16821
rect 1539 16659 1581 16701
rect 1659 16659 1701 16701
rect 13119 16779 13161 16821
rect 14439 16779 14481 16821
rect 15939 16719 15981 16761
rect 16479 16719 16521 16761
rect 6819 16659 6861 16701
rect 13359 16659 13401 16701
rect 14679 16659 14721 16701
rect 1659 16596 1701 16638
rect 3279 16599 3321 16641
rect 3459 16599 3501 16641
rect 10341 16599 10383 16641
rect 10479 16599 10521 16641
rect 15399 16599 15441 16641
rect 15579 16599 15621 16641
rect 15699 16599 15741 16641
rect 4899 16539 4941 16581
rect 5139 16539 5181 16581
rect 5739 16479 5781 16521
rect 5919 16479 5961 16521
rect 3219 16179 3261 16221
rect 7839 16119 7881 16161
rect 8079 16119 8121 16161
rect 8499 16119 8541 16161
rect 3399 15999 3441 16041
rect 4659 15999 4701 16041
rect 7839 15999 7881 16041
rect 8079 15999 8121 16041
rect 8499 15999 8541 16041
rect 8919 16119 8961 16161
rect 9519 16119 9561 16161
rect 8919 15999 8961 16041
rect 9519 15999 9561 16041
rect 10179 16119 10221 16161
rect 10899 16119 10941 16161
rect 13059 16119 13101 16161
rect 16899 16119 16941 16161
rect 10179 15999 10221 16041
rect 10899 15999 10941 16041
rect 12699 15999 12741 16041
rect 12819 15999 12861 16041
rect 13059 15999 13101 16041
rect 16719 15999 16761 16041
rect 3339 15939 3381 15981
rect 3459 15939 3501 15981
rect 5919 15939 5961 15981
rect 6159 15939 6201 15981
rect 7119 15939 7161 15981
rect 7539 15939 7581 15981
rect 9579 15939 9621 15981
rect 9819 15939 9861 15981
rect 9939 15939 9981 15981
rect 10119 15936 10161 15978
rect 14079 15939 14121 15981
rect 14319 15939 14361 15981
rect 7659 15879 7701 15921
rect 7899 15879 7941 15921
rect 12459 15519 12501 15561
rect 12579 15519 12621 15561
rect 5079 15219 5121 15261
rect 7299 15219 7341 15261
rect 7779 15219 7821 15261
rect 9579 15219 9621 15261
rect 9699 15219 9741 15261
rect 10539 15219 10581 15261
rect 10659 15216 10701 15258
rect 10959 15219 11001 15261
rect 12159 15279 12201 15321
rect 3459 15099 3501 15141
rect 3579 15099 3621 15141
rect 5079 15099 5121 15141
rect 7419 15099 7461 15141
rect 7959 15099 8001 15141
rect 8199 15099 8241 15141
rect 8319 15099 8361 15141
rect 10959 15099 11001 15141
rect 11919 15099 11961 15141
rect 12579 15219 12621 15261
rect 13959 15219 14001 15261
rect 14259 15219 14301 15261
rect 15339 15279 15381 15321
rect 15579 15219 15621 15261
rect 12579 15099 12621 15141
rect 13959 15099 14001 15141
rect 14379 15099 14421 15141
rect 15099 15099 15141 15141
rect 4179 15039 4221 15081
rect 4659 15039 4701 15081
rect 9639 15039 9681 15081
rect 9759 15039 9801 15081
rect 16179 15219 16221 15261
rect 15999 15099 16041 15141
rect 15759 15039 15801 15081
rect 17139 14739 17181 14781
rect 17259 14739 17301 14781
rect 6279 14619 6321 14661
rect 6399 14619 6441 14661
rect 7839 14616 7881 14658
rect 8019 14619 8061 14661
rect 8199 14559 8241 14601
rect 7839 14439 7881 14481
rect 8199 14439 8241 14481
rect 8439 14559 8481 14601
rect 9159 14559 9201 14601
rect 2739 14379 2781 14421
rect 3039 14379 3081 14421
rect 6819 14379 6861 14421
rect 6999 14379 7041 14421
rect 10119 14559 10161 14601
rect 10779 14559 10821 14601
rect 8379 14376 8421 14418
rect 9399 14379 9441 14421
rect 9939 14379 9981 14421
rect 10779 14439 10821 14481
rect 12459 14619 12501 14661
rect 13899 14619 13941 14661
rect 14079 14619 14121 14661
rect 12999 14559 13041 14601
rect 13599 14559 13641 14601
rect 14019 14559 14061 14601
rect 14439 14559 14481 14601
rect 14739 14559 14781 14601
rect 12279 14439 12321 14481
rect 12999 14439 13041 14481
rect 13479 14439 13521 14481
rect 13899 14439 13941 14481
rect 14439 14439 14481 14481
rect 15459 14559 15501 14601
rect 15999 14619 16041 14661
rect 14919 14439 14961 14481
rect 15459 14439 15501 14481
rect 15759 14439 15801 14481
rect 16359 14559 16401 14601
rect 17559 14559 17601 14601
rect 18219 14499 18261 14541
rect 16359 14439 16401 14481
rect 17559 14439 17601 14481
rect 17679 14439 17721 14481
rect 15159 14379 15201 14421
rect 15339 14379 15381 14421
rect 17019 14379 17061 14421
rect 17259 14379 17301 14421
rect 13419 14259 13461 14301
rect 13539 14259 13581 14301
rect 17979 14139 18021 14181
rect 15519 13959 15561 14001
rect 15759 13959 15801 14001
rect 13959 13839 14001 13881
rect 14199 13839 14241 13881
rect 1179 13722 1221 13764
rect 1419 13719 1461 13761
rect 8739 13719 8781 13761
rect 15159 13719 15201 13761
rect 17979 13719 18021 13761
rect 3879 13659 3921 13701
rect 7299 13659 7341 13701
rect 1839 13599 1881 13641
rect 2979 13599 3021 13641
rect 8379 13659 8421 13701
rect 7839 13599 7881 13641
rect 1959 13539 2001 13581
rect 2439 13539 2481 13581
rect 3999 13539 4041 13581
rect 4239 13539 4281 13581
rect 4359 13539 4401 13581
rect 8259 13539 8301 13581
rect 10539 13659 10581 13701
rect 14019 13659 14061 13701
rect 9999 13599 10041 13641
rect 10479 13599 10521 13641
rect 8679 13539 8721 13581
rect 14199 13599 14241 13641
rect 14019 13539 14061 13581
rect 14739 13539 14781 13581
rect 15039 13539 15081 13581
rect 15219 13659 15261 13701
rect 16419 13659 16461 13701
rect 15219 13539 15261 13581
rect 16899 13659 16941 13701
rect 5079 13479 5121 13521
rect 5319 13479 5361 13521
rect 5979 13479 6021 13521
rect 6159 13479 6201 13521
rect 10479 13479 10521 13521
rect 17679 13539 17721 13581
rect 17919 13539 17961 13581
rect 16659 13479 16701 13521
rect 3699 13179 3741 13221
rect 3819 13179 3861 13221
rect 13779 13119 13821 13161
rect 1299 12999 1341 13041
rect 7359 12999 7401 13041
rect 8019 12999 8061 13041
rect 4719 12939 4761 12981
rect 2859 12879 2901 12921
rect 4299 12876 4341 12918
rect 7479 12939 7521 12981
rect 13299 12999 13341 13041
rect 13659 12996 13701 13038
rect 14019 13059 14061 13101
rect 14319 13059 14361 13101
rect 15639 13059 15681 13101
rect 15879 13059 15921 13101
rect 14139 12999 14181 13041
rect 15039 12999 15081 13041
rect 15339 12999 15381 13041
rect 1479 12819 1521 12861
rect 4059 12819 4101 12861
rect 14319 12879 14361 12921
rect 14859 12879 14901 12921
rect 16059 12999 16101 13041
rect 16539 12999 16581 13041
rect 16659 12999 16701 13041
rect 17139 12999 17181 13041
rect 17439 12999 17481 13041
rect 15519 12879 15561 12921
rect 16059 12879 16101 12921
rect 6039 12819 6081 12861
rect 6339 12819 6381 12861
rect 7539 12819 7581 12861
rect 13539 12819 13581 12861
rect 13779 12819 13821 12861
rect 13959 12819 14001 12861
rect 14259 12819 14301 12861
rect 17199 12819 17241 12861
rect 17379 12819 17421 12861
rect 7719 12579 7761 12621
rect 7959 12279 8001 12321
rect 8019 12279 8061 12321
rect 579 12159 621 12201
rect 819 12159 861 12201
rect 5319 12159 5361 12201
rect 5559 12159 5601 12201
rect 5859 12159 5901 12201
rect 6039 12159 6081 12201
rect 7059 12159 7101 12201
rect 7179 12159 7221 12201
rect 12219 12159 12261 12201
rect 12459 12159 12501 12201
rect 12939 12159 12981 12201
rect 13239 12156 13281 12198
rect 15579 12159 15621 12201
rect 15879 12159 15921 12201
rect 17079 12159 17121 12201
rect 17259 12156 17301 12198
rect 17739 12162 17781 12204
rect 17979 12159 18021 12201
rect 2679 12099 2721 12141
rect 4779 12099 4821 12141
rect 4959 12099 5001 12141
rect 3279 12039 3321 12081
rect 1359 11979 1401 12021
rect 1539 11979 1581 12021
rect 4779 11979 4821 12021
rect 5619 12099 5661 12141
rect 5979 12099 6021 12141
rect 5199 11979 5241 12021
rect 5499 11979 5541 12021
rect 6399 12099 6441 12141
rect 8319 12099 8361 12141
rect 6219 11979 6261 12021
rect 8319 11979 8361 12021
rect 8859 12099 8901 12141
rect 12699 12099 12741 12141
rect 13839 12099 13881 12141
rect 8859 11979 8901 12021
rect 5859 11919 5901 11961
rect 6999 11919 7041 11961
rect 7119 11919 7161 11961
rect 12759 11919 12801 11961
rect 13479 11919 13521 11961
rect 13659 11919 13701 11961
rect 15339 12099 15381 12141
rect 16179 12099 16221 12141
rect 18219 12162 18261 12204
rect 16659 12039 16701 12081
rect 14739 11979 14781 12021
rect 15339 11979 15381 12021
rect 15999 11979 16041 12021
rect 18039 11979 18081 12021
rect 13899 11856 13941 11898
rect 7839 11619 7881 11661
rect 7959 11616 8001 11658
rect 7899 11556 7941 11598
rect 8139 11559 8181 11601
rect 17019 11559 17061 11601
rect 17139 11559 17181 11601
rect 4479 11499 4521 11541
rect 2319 11439 2361 11481
rect 2559 11439 2601 11481
rect 2679 11439 2721 11481
rect 3699 11439 3741 11481
rect 4059 11439 4101 11481
rect 4839 11499 4881 11541
rect 5799 11499 5841 11541
rect 14859 11499 14901 11541
rect 14979 11499 15021 11541
rect 15099 11499 15141 11541
rect 17379 11499 17421 11541
rect 17619 11499 17661 11541
rect 2319 11319 2361 11361
rect 3699 11319 3741 11361
rect 4119 11319 4161 11361
rect 4659 11319 4701 11361
rect 4899 11319 4941 11361
rect 5679 11319 5721 11361
rect 5859 11439 5901 11481
rect 6399 11439 6441 11481
rect 8439 11439 8481 11481
rect 11919 11439 11961 11481
rect 17019 11439 17061 11481
rect 5859 11319 5901 11361
rect 6159 11319 6201 11361
rect 2739 11259 2781 11301
rect 2919 11259 2961 11301
rect 5139 11253 5181 11295
rect 5259 11259 5301 11301
rect 6219 11259 6261 11301
rect 6399 11259 6441 11301
rect 17439 11439 17481 11481
rect 17799 11439 17841 11481
rect 11979 11316 12021 11358
rect 17199 11319 17241 11361
rect 17559 11319 17601 11361
rect 17799 11319 17841 11361
rect 8379 11256 8421 11298
rect 9159 11259 9201 11301
rect 9399 11259 9441 11301
rect 16839 11259 16881 11301
rect 17259 11259 17301 11301
rect 17379 11253 17421 11295
rect 17619 11259 17661 11301
rect 8019 10839 8061 10881
rect 8139 10839 8181 10881
rect 5559 10719 5601 10761
rect 5799 10719 5841 10761
rect 4659 10659 4701 10701
rect 4959 10659 5001 10701
rect 159 10599 201 10641
rect 399 10599 441 10641
rect 1479 10599 1521 10641
rect 1779 10599 1821 10641
rect 4899 10539 4941 10581
rect 5859 10599 5901 10641
rect 8379 10599 8421 10641
rect 8559 10599 8601 10641
rect 16419 10599 16461 10641
rect 16599 10599 16641 10641
rect 5679 10476 5721 10518
rect 6159 10539 6201 10581
rect 11319 10539 11361 10581
rect 11439 10539 11481 10581
rect 13419 10539 13461 10581
rect 15999 10539 16041 10581
rect 4899 10419 4941 10461
rect 6159 10419 6201 10461
rect 13299 10419 13341 10461
rect 17139 10599 17181 10641
rect 18039 10539 18081 10581
rect 15999 10419 16041 10461
rect 16899 10419 16941 10461
rect 17859 10419 17901 10461
rect 6759 10359 6801 10401
rect 7059 10359 7101 10401
rect 7479 10059 7521 10101
rect 7659 10059 7701 10101
rect 9099 10059 9141 10101
rect 7119 9939 7161 9981
rect 9099 9939 9141 9981
rect 15459 9939 15501 9981
rect 1779 9879 1821 9921
rect 1779 9759 1821 9801
rect 1959 9879 2001 9921
rect 2259 9879 2301 9921
rect 2259 9759 2301 9801
rect 4659 9879 4701 9921
rect 4839 9879 4881 9921
rect 5799 9879 5841 9921
rect 4659 9759 4701 9801
rect 1359 9699 1401 9741
rect 1539 9699 1581 9741
rect 1899 9699 1941 9741
rect 3579 9699 3621 9741
rect 3819 9699 3861 9741
rect 5799 9759 5841 9801
rect 7179 9879 7221 9921
rect 7899 9879 7941 9921
rect 8619 9879 8661 9921
rect 10119 9879 10161 9921
rect 12159 9879 12201 9921
rect 7179 9759 7221 9801
rect 7899 9759 7941 9801
rect 14619 9879 14661 9921
rect 8799 9759 8841 9801
rect 10119 9759 10161 9801
rect 12159 9759 12201 9801
rect 13239 9759 13281 9801
rect 14439 9759 14481 9801
rect 15279 9759 15321 9801
rect 16599 9879 16641 9921
rect 17859 9876 17901 9918
rect 16599 9759 16641 9801
rect 5079 9699 5121 9741
rect 6999 9699 7041 9741
rect 7239 9699 7281 9741
rect 7479 9699 7521 9741
rect 7659 9693 7701 9735
rect 11619 9699 11661 9741
rect 11979 9699 12021 9741
rect 13239 9696 13281 9738
rect 13359 9699 13401 9741
rect 14799 9699 14841 9741
rect 15039 9699 15081 9741
rect 13179 9636 13221 9678
rect 18099 9636 18141 9678
rect 16899 9576 16941 9618
rect 17019 9579 17061 9621
rect 6279 9279 6321 9321
rect 6459 9279 6501 9321
rect 819 9039 861 9081
rect 1179 9039 1221 9081
rect 4959 9039 5001 9081
rect 5139 9039 5181 9081
rect 5799 9039 5841 9081
rect 6099 9039 6141 9081
rect 8139 9039 8181 9081
rect 8259 9039 8301 9081
rect 8439 9042 8481 9084
rect 8679 9036 8721 9078
rect 3219 8979 3261 9021
rect 4239 8979 4281 9021
rect 5439 8976 5481 9018
rect 5559 8979 5601 9021
rect 5859 8979 5901 9021
rect 2379 8859 2421 8901
rect 2559 8859 2601 8901
rect 3219 8859 3261 8901
rect 3999 8859 4041 8901
rect 6519 8979 6561 9021
rect 7719 8979 7761 9021
rect 9159 8979 9201 9021
rect 9519 8979 9561 9021
rect 9819 8979 9861 9021
rect 6519 8859 6561 8901
rect 5919 8799 5961 8841
rect 6699 8799 6741 8841
rect 6999 8799 7041 8841
rect 7779 8799 7821 8841
rect 9519 8859 9561 8901
rect 9819 8859 9861 8901
rect 12039 8979 12081 9021
rect 12279 8979 12321 9021
rect 12819 8979 12861 9021
rect 15999 8979 16041 9021
rect 16959 8979 17001 9021
rect 12039 8859 12081 8901
rect 12519 8859 12561 8901
rect 12939 8859 12981 8901
rect 14799 8859 14841 8901
rect 14919 8859 14961 8901
rect 15999 8859 16041 8901
rect 16779 8859 16821 8901
rect 9099 8796 9141 8838
rect 15459 8799 15501 8841
rect 15639 8799 15681 8841
rect 17439 8739 17481 8781
rect 17619 8739 17661 8781
rect 16599 8499 16641 8541
rect 17019 8499 17061 8541
rect 4899 8439 4941 8481
rect 5139 8439 5181 8481
rect 16659 8439 16701 8481
rect 16959 8439 17001 8481
rect 4419 8379 4461 8421
rect 4539 8379 4581 8421
rect 2919 8319 2961 8361
rect 2919 8199 2961 8241
rect 1239 8139 1281 8181
rect 1599 8139 1641 8181
rect 2619 8139 2661 8181
rect 2859 8139 2901 8181
rect 4779 8376 4821 8418
rect 5739 8379 5781 8421
rect 5979 8379 6021 8421
rect 7359 8379 7401 8421
rect 7599 8379 7641 8421
rect 16059 8379 16101 8421
rect 16299 8376 16341 8418
rect 16539 8379 16581 8421
rect 5139 8319 5181 8361
rect 6339 8319 6381 8361
rect 6759 8319 6801 8361
rect 6279 8256 6321 8298
rect 4899 8199 4941 8241
rect 7539 8319 7581 8361
rect 8379 8319 8421 8361
rect 9099 8319 9141 8361
rect 7779 8259 7821 8301
rect 9879 8319 9921 8361
rect 15339 8319 15381 8361
rect 15639 8319 15681 8361
rect 15999 8319 16041 8361
rect 9279 8259 9321 8301
rect 9759 8259 9801 8301
rect 6759 8199 6801 8241
rect 7359 8199 7401 8241
rect 7719 8199 7761 8241
rect 8259 8199 8301 8241
rect 9099 8199 9141 8241
rect 15219 8256 15261 8298
rect 16239 8319 16281 8361
rect 16119 8259 16161 8301
rect 17259 8379 17301 8421
rect 17439 8379 17481 8421
rect 17679 8382 17721 8424
rect 9879 8199 9921 8241
rect 15279 8199 15321 8241
rect 15759 8199 15801 8241
rect 15999 8199 16041 8241
rect 16599 8199 16641 8241
rect 17019 8319 17061 8361
rect 17379 8319 17421 8361
rect 17019 8199 17061 8241
rect 17379 8199 17421 8241
rect 17739 8199 17781 8241
rect 4599 8136 4641 8178
rect 6519 8139 6561 8181
rect 6639 8139 6681 8181
rect 7419 8139 7461 8181
rect 7599 8139 7641 8181
rect 7839 8139 7881 8181
rect 7959 8139 8001 8181
rect 15339 8139 15381 8181
rect 15939 8133 15981 8175
rect 16119 8139 16161 8181
rect 2799 8019 2841 8061
rect 2919 8019 2961 8061
rect 5859 7599 5901 7641
rect 6099 7599 6141 7641
rect 3279 7539 3321 7581
rect 3519 7539 3561 7581
rect 4059 7479 4101 7521
rect 4299 7479 4341 7521
rect 5901 7479 5943 7521
rect 6159 7479 6201 7521
rect 8079 7479 8121 7521
rect 8559 7479 8601 7521
rect 10959 7479 11001 7521
rect 11199 7482 11241 7524
rect 13119 7479 13161 7521
rect 459 7419 501 7461
rect 3099 7419 3141 7461
rect 3639 7419 3681 7461
rect 3759 7419 3801 7461
rect 7239 7419 7281 7461
rect 579 7299 621 7341
rect 2919 7239 2961 7281
rect 3699 7356 3741 7398
rect 8319 7419 8361 7461
rect 8739 7419 8781 7461
rect 9279 7419 9321 7461
rect 10059 7419 10101 7461
rect 3819 7299 3861 7341
rect 7419 7299 7461 7341
rect 8139 7299 8181 7341
rect 8739 7299 8781 7341
rect 14019 7419 14061 7461
rect 14439 7419 14481 7461
rect 15279 7419 15321 7461
rect 17019 7419 17061 7461
rect 9399 7299 9441 7341
rect 10179 7299 10221 7341
rect 13179 7299 13221 7341
rect 14199 7299 14241 7341
rect 14439 7299 14481 7341
rect 17619 7419 17661 7461
rect 18039 7479 18081 7521
rect 15399 7299 15441 7341
rect 17139 7299 17181 7341
rect 17439 7299 17481 7341
rect 17859 7299 17901 7341
rect 8139 7236 8181 7278
rect 8439 7239 8481 7281
rect 15219 6939 15261 6981
rect 15339 6939 15381 6981
rect 5019 6879 5061 6921
rect 5199 6879 5241 6921
rect 6519 6819 6561 6861
rect 7179 6819 7221 6861
rect 7359 6819 7401 6861
rect 219 6759 261 6801
rect 1479 6759 1521 6801
rect 639 6699 681 6741
rect 519 6639 561 6681
rect 3399 6759 3441 6801
rect 5079 6759 5121 6801
rect 5619 6759 5661 6801
rect 6159 6759 6201 6801
rect 1599 6639 1641 6681
rect 2499 6639 2541 6681
rect 2619 6639 2661 6681
rect 279 6573 321 6615
rect 3099 6579 3141 6621
rect 4659 6639 4701 6681
rect 4839 6639 4881 6681
rect 5199 6639 5241 6681
rect 7119 6759 7161 6801
rect 8079 6759 8121 6801
rect 9639 6759 9681 6801
rect 11619 6759 11661 6801
rect 12039 6759 12081 6801
rect 5439 6579 5481 6621
rect 6159 6639 6201 6681
rect 6579 6639 6621 6681
rect 7299 6636 7341 6678
rect 8139 6636 8181 6678
rect 9639 6639 9681 6681
rect 5679 6579 5721 6621
rect 12039 6639 12081 6681
rect 12219 6759 12261 6801
rect 14559 6759 14601 6801
rect 14679 6759 14721 6801
rect 15159 6759 15201 6801
rect 12219 6639 12261 6681
rect 15399 6639 15441 6681
rect 11799 6579 11841 6621
rect 15999 6519 16041 6561
rect 16239 6519 16281 6561
rect 5919 6459 5961 6501
rect 6219 6459 6261 6501
rect 4719 6039 4761 6081
rect 4959 6039 5001 6081
rect 6459 6039 6501 6081
rect 6639 6039 6681 6081
rect 13419 6039 13461 6081
rect 13599 6039 13641 6081
rect 7419 5979 7461 6021
rect 7539 5979 7581 6021
rect 10239 5979 10281 6021
rect 10359 5979 10401 6021
rect 17079 5979 17121 6021
rect 17319 5976 17361 6018
rect 1899 5919 1941 5961
rect 2019 5919 2061 5961
rect 2619 5919 2661 5961
rect 3099 5919 3141 5961
rect 3219 5919 3261 5961
rect 5499 5919 5541 5961
rect 5799 5919 5841 5961
rect 6819 5919 6861 5961
rect 6999 5919 7041 5961
rect 7299 5919 7341 5961
rect 7539 5916 7581 5958
rect 12519 5919 12561 5961
rect 12699 5919 12741 5961
rect 13719 5919 13761 5961
rect 5259 5859 5301 5901
rect 5979 5859 6021 5901
rect 8199 5859 8241 5901
rect 2679 5739 2721 5781
rect 5139 5739 5181 5781
rect 5979 5739 6021 5781
rect 8379 5859 8421 5901
rect 12939 5859 12981 5901
rect 8379 5739 8421 5781
rect 15939 5919 15981 5961
rect 16659 5919 16701 5961
rect 16899 5919 16941 5961
rect 17079 5916 17121 5958
rect 17259 5919 17301 5961
rect 12999 5736 13041 5778
rect 13779 5739 13821 5781
rect 8319 5679 8361 5721
rect 9099 5679 9141 5721
rect 13479 5679 13521 5721
rect 13599 5679 13641 5721
rect 16119 5859 16161 5901
rect 16119 5739 16161 5781
rect 16839 5859 16881 5901
rect 17559 5859 17601 5901
rect 17739 5739 17781 5781
rect 15939 5679 15981 5721
rect 16839 5679 16881 5721
rect 17139 5679 17181 5721
rect 17319 5679 17361 5721
rect 8919 5619 8961 5661
rect 4839 5319 4881 5361
rect 16059 5319 16101 5361
rect 16179 5319 16221 5361
rect 519 5199 561 5241
rect 999 5199 1041 5241
rect 1119 5199 1161 5241
rect 10479 5259 10521 5301
rect 10719 5259 10761 5301
rect 10959 5259 11001 5301
rect 5259 5199 5301 5241
rect 639 5079 681 5121
rect 4899 5079 4941 5121
rect 5199 5079 5241 5121
rect 5919 5199 5961 5241
rect 6339 5199 6381 5241
rect 6759 5199 6801 5241
rect 15699 5256 15741 5298
rect 15819 5259 15861 5301
rect 5619 5019 5661 5061
rect 6219 5079 6261 5121
rect 11379 5199 11421 5241
rect 12459 5199 12501 5241
rect 13599 5199 13641 5241
rect 15639 5199 15681 5241
rect 6759 5079 6801 5121
rect 10479 5079 10521 5121
rect 11379 5079 11421 5121
rect 12459 5079 12501 5121
rect 6159 5019 6201 5061
rect 6399 5019 6441 5061
rect 8199 5013 8241 5055
rect 8319 5019 8361 5061
rect 13299 5019 13341 5061
rect 13419 5019 13461 5061
rect 16479 5199 16521 5241
rect 15759 5079 15801 5121
rect 16299 5079 16341 5121
rect 13779 5013 13821 5055
rect 5019 4959 5061 5001
rect 5319 4959 5361 5001
rect 17013 4779 17055 4821
rect 10299 4599 10341 4641
rect 10479 4599 10521 4641
rect 17739 4551 17781 4593
rect 5619 4419 5661 4461
rect 5919 4419 5961 4461
rect 3399 4359 3441 4401
rect 3699 4359 3741 4401
rect 4839 4359 4881 4401
rect 4959 4359 5001 4401
rect 5199 4359 5241 4401
rect 5439 4359 5481 4401
rect 12759 4359 12801 4401
rect 13119 4359 13161 4401
rect 14199 4359 14241 4401
rect 14379 4359 14421 4401
rect 18099 4359 18141 4401
rect 18219 4359 18261 4401
rect 5919 4299 5961 4341
rect 6579 4299 6621 4341
rect 1719 4179 1761 4221
rect 1839 4179 1881 4221
rect 5919 4179 5961 4221
rect 6579 4179 6621 4221
rect 8739 4299 8781 4341
rect 9819 4299 9861 4341
rect 10239 4299 10281 4341
rect 8739 4179 8781 4221
rect 13959 4299 14001 4341
rect 15579 4299 15621 4341
rect 10239 4179 10281 4221
rect 13779 4179 13821 4221
rect 15939 4299 15981 4341
rect 15759 4179 15801 4221
rect 16059 4179 16101 4221
rect 18159 4179 18201 4221
rect 18339 4179 18381 4221
rect 4419 4119 4461 4161
rect 4599 4119 4641 4161
rect 9819 4119 9861 4161
rect 10299 4116 10341 4158
rect 10479 4119 10521 4161
rect 17799 4059 17841 4101
rect 17979 4059 18021 4101
rect 13299 3699 13341 3741
rect 13419 3699 13461 3741
rect 16539 3699 16581 3741
rect 6819 3639 6861 3681
rect 99 3579 141 3621
rect 219 3519 261 3561
rect 9099 3639 9141 3681
rect 10839 3639 10881 3681
rect 11139 3639 11181 3681
rect 7059 3519 7101 3561
rect 9099 3519 9141 3561
rect 10959 3519 11001 3561
rect 1719 3459 1761 3501
rect 1839 3453 1881 3495
rect 3579 3459 3621 3501
rect 3699 3459 3741 3501
rect 11319 3639 11361 3681
rect 11319 3519 11361 3561
rect 16359 3519 16401 3561
rect 18219 3579 18261 3621
rect 11379 3459 11421 3501
rect 11679 3459 11721 3501
rect 11859 3459 11901 3501
rect 15639 3459 15681 3501
rect 15879 3459 15921 3501
rect 18219 3399 18261 3441
rect 18027 3279 18069 3321
rect 9459 3036 9501 3078
rect 9579 3039 9621 3081
rect 6519 2919 6561 2961
rect 6339 2859 6381 2901
rect 15159 2859 15201 2901
rect 15279 2859 15321 2901
rect 339 2799 381 2841
rect 759 2799 801 2841
rect 3039 2799 3081 2841
rect 3219 2799 3261 2841
rect 3579 2799 3621 2841
rect 3939 2799 3981 2841
rect 4479 2799 4521 2841
rect 4659 2799 4701 2841
rect 7599 2799 7641 2841
rect 7899 2799 7941 2841
rect 12501 2799 12543 2841
rect 12639 2799 12681 2841
rect 12879 2802 12921 2844
rect 13179 2799 13221 2841
rect 16959 2799 17001 2841
rect 17079 2802 17121 2844
rect 4719 2736 4761 2778
rect 4839 2739 4881 2781
rect 5919 2739 5961 2781
rect 6039 2739 6081 2781
rect 12099 2739 12141 2781
rect 15279 2739 15321 2781
rect 15699 2739 15741 2781
rect 16359 2739 16401 2781
rect 15279 2619 15321 2661
rect 15579 2619 15621 2661
rect 16359 2619 16401 2661
rect 9819 2559 9861 2601
rect 9999 2559 10041 2601
rect 12219 2559 12261 2601
rect 5559 2139 5601 2181
rect 5679 2139 5721 2181
rect 8919 2139 8961 2181
rect 9159 2139 9201 2181
rect 11739 2139 11781 2181
rect 11919 2139 11961 2181
rect 12759 2139 12801 2181
rect 12999 2139 13041 2181
rect 14739 2139 14781 2181
rect 3819 2079 3861 2121
rect 5139 2079 5181 2121
rect 3939 1959 3981 2001
rect 6219 2079 6261 2121
rect 6699 2079 6741 2121
rect 8859 2079 8901 2121
rect 9039 2079 9081 2121
rect 9519 2079 9561 2121
rect 9459 2019 9501 2061
rect 11319 2019 11361 2061
rect 6039 1959 6081 2001
rect 6519 1959 6561 2001
rect 9399 1959 9441 2001
rect 9519 1959 9561 2001
rect 11139 1959 11181 2001
rect 11259 1959 11301 2001
rect 17499 2079 17541 2121
rect 14559 1959 14601 2001
rect 17379 1959 17421 2001
rect 4599 1899 4641 1941
rect 5019 1899 5061 1941
rect 5319 1899 5361 1941
rect 11319 1899 11361 1941
rect 11499 1899 11541 1941
rect 11859 1899 11901 1941
rect 1359 1239 1401 1281
rect 1479 1239 1521 1281
rect 6339 1239 6381 1281
rect 6819 1239 6861 1281
rect 8139 1239 8181 1281
rect 8379 1239 8421 1281
rect 8619 1239 8661 1281
rect 17559 1239 17601 1281
rect 17739 1239 17781 1281
rect 4779 1179 4821 1221
rect 6639 1179 6681 1221
rect 9639 1179 9681 1221
rect 9639 1059 9681 1101
rect 9819 1179 9861 1221
rect 2619 999 2661 1041
rect 2799 999 2841 1041
rect 5079 999 5121 1041
rect 5379 999 5421 1041
rect 6519 999 6561 1041
rect 9699 996 9741 1038
rect 10839 999 10881 1041
rect 11019 993 11061 1035
rect 6039 939 6081 981
rect 6159 939 6201 981
rect 5019 879 5061 921
rect 5259 879 5301 921
rect 4839 699 4881 741
rect 5019 699 5061 741
rect 8499 579 8541 621
rect 8739 579 8781 621
rect 4419 519 4461 561
rect 4599 519 4641 561
rect 7659 519 7701 561
rect 8859 519 8901 561
rect 12399 519 12441 561
rect 6279 399 6321 441
rect 6399 399 6441 441
rect 7539 399 7581 441
rect 12039 459 12081 501
rect 8979 399 9021 441
rect 11499 399 11541 441
rect 13359 519 13401 561
rect 1719 339 1761 381
rect 2019 339 2061 381
rect 2979 339 3021 381
rect 3279 339 3321 381
rect 3456 339 3498 381
rect 3519 339 3561 381
rect 3759 339 3801 381
rect 6219 339 6261 381
rect 6579 339 6621 381
rect 13239 399 13281 441
rect 12639 339 12681 381
rect 17919 339 17961 381
rect 18219 339 18261 381
rect 3699 276 3741 318
rect 8379 99 8421 141
rect 8499 99 8541 141
<< metal2 >>
rect 10008 18801 10032 18912
rect 14568 18801 14592 18912
rect 288 18348 312 18459
rect 768 18348 792 18459
rect 888 18381 912 18639
rect 528 18252 552 18342
rect 1188 18348 1212 18459
rect 1548 18384 1572 18519
rect 948 18261 972 18342
rect 1788 18261 1812 18399
rect 1968 18348 1992 18639
rect 2208 18372 2232 18519
rect 2268 18441 2292 18579
rect 2208 18348 2292 18372
rect 2379 18360 2421 18399
rect 2388 18348 2412 18360
rect 348 17781 372 18252
rect 528 18228 612 18252
rect 339 17700 381 17739
rect 348 17688 372 17700
rect 588 17721 612 18228
rect 828 17724 852 18216
rect 1128 17901 1152 18252
rect 1179 17724 1221 17742
rect 288 17481 312 17592
rect 288 16881 312 17439
rect 48 15741 72 16122
rect 108 15138 132 16539
rect 288 16461 312 16692
rect 408 16581 432 17592
rect 528 17361 552 17592
rect 588 17481 612 17559
rect 468 16452 492 17139
rect 648 17001 672 17679
rect 768 17361 792 17592
rect 888 17121 912 17556
rect 1008 17541 1032 17682
rect 1128 17481 1152 17592
rect 561 16812 600 16821
rect 561 16788 612 16812
rect 561 16779 600 16788
rect 441 16428 492 16452
rect 168 15264 192 16299
rect 408 16164 432 16419
rect 288 15861 312 16032
rect 468 16020 492 16032
rect 459 15981 501 16020
rect 588 15981 612 16359
rect 648 16038 672 16179
rect 768 16128 792 16299
rect 828 16221 852 16959
rect 1119 16800 1161 16839
rect 1188 16821 1212 17499
rect 1428 17481 1452 18216
rect 1608 18141 1632 18252
rect 2328 18141 2352 18216
rect 2568 18201 2592 18399
rect 2628 18321 2652 18459
rect 2748 18348 2772 18639
rect 10608 18621 10632 18699
rect 3288 18348 3312 18459
rect 1659 17700 1701 17739
rect 1668 17688 1692 17700
rect 1788 17688 1812 17979
rect 1908 17961 1932 18099
rect 2388 17961 2412 18039
rect 2568 18021 2592 18159
rect 2928 18081 2952 18252
rect 3048 17961 3072 18342
rect 1908 17928 1959 17961
rect 1920 17919 1959 17928
rect 1299 16824 1341 16839
rect 1128 16788 1152 16800
rect 888 16701 912 16782
rect 1428 16788 1452 17139
rect 1488 16872 1512 17679
rect 1848 17481 1872 17556
rect 1488 16860 1572 16872
rect 1488 16848 1581 16860
rect 1539 16821 1581 16848
rect 888 16401 912 16659
rect 1500 16692 1539 16701
rect 1188 16461 1212 16659
rect 1368 16461 1392 16692
rect 1488 16668 1539 16692
rect 1500 16659 1539 16668
rect 1608 16641 1632 16782
rect 1668 16701 1692 17439
rect 888 16128 912 16239
rect 948 15861 972 16032
rect 288 15228 312 15399
rect 348 15120 372 15132
rect 339 15081 381 15120
rect 588 14652 612 15639
rect 1008 15441 1032 15819
rect 1068 15681 1092 16419
rect 1248 16128 1272 16239
rect 1428 16032 1452 16599
rect 1668 16281 1692 16596
rect 1668 16128 1692 16239
rect 1728 16221 1752 16899
rect 1848 16872 1872 17139
rect 1908 16941 1932 17859
rect 3228 17841 3252 18252
rect 3588 17961 3612 18459
rect 4128 18348 4152 18459
rect 4308 18258 4332 18579
rect 4968 18348 4992 18459
rect 5088 18348 5199 18372
rect 5328 18348 5352 18459
rect 3768 18240 3792 18252
rect 3759 18201 3801 18240
rect 2148 17580 2172 17592
rect 2139 17541 2181 17580
rect 2328 17421 2352 17592
rect 1848 16848 1932 16872
rect 1908 16788 1932 16848
rect 2148 16701 2172 17379
rect 2448 17121 2472 17679
rect 2379 16872 2421 16899
rect 2328 16860 2421 16872
rect 2328 16848 2412 16860
rect 2328 16788 2352 16848
rect 2568 16761 2592 16959
rect 1968 16461 1992 16692
rect 2628 16581 2652 17592
rect 2748 17580 2772 17592
rect 2739 17541 2781 17580
rect 2808 16581 2832 16692
rect 2988 16341 3012 17799
rect 3468 17688 3612 17712
rect 3699 17700 3741 17739
rect 3708 17688 3732 17700
rect 3108 17580 3132 17592
rect 3099 17541 3141 17580
rect 3288 17061 3312 17592
rect 3108 16788 3132 16899
rect 3288 16788 3312 17019
rect 3408 16881 3432 17682
rect 3468 17061 3492 17688
rect 4008 17688 4032 18159
rect 4068 18021 4092 18252
rect 4188 18081 4212 18252
rect 4188 17841 4212 18039
rect 4068 17481 4092 17592
rect 3408 16701 3432 16839
rect 3468 16824 3492 17019
rect 3768 17001 3792 17439
rect 3699 16800 3741 16839
rect 3768 16821 3792 16959
rect 3708 16788 3732 16800
rect 1848 16038 1872 16179
rect 2019 16140 2061 16179
rect 2028 16128 2052 16140
rect 2268 16038 2292 16239
rect 2508 16128 2532 16239
rect 1188 15921 1212 16032
rect 828 14961 852 15132
rect 561 14628 612 14652
rect 288 14241 312 14472
rect 408 14460 432 14472
rect 399 14421 441 14460
rect 48 12972 72 13959
rect 228 13704 252 13779
rect 468 13704 492 14439
rect 528 14421 552 14619
rect 699 14580 741 14619
rect 708 14568 732 14580
rect 948 14478 972 14559
rect 528 13701 552 14379
rect 648 14241 672 14472
rect 768 14361 792 14472
rect 1008 14412 1032 15399
rect 1068 15081 1092 15279
rect 1248 15228 1272 15939
rect 1308 15801 1332 16032
rect 1428 16008 1512 16032
rect 1368 15228 1392 15399
rect 1188 14721 1212 15132
rect 1308 14961 1332 15132
rect 1488 15021 1512 16008
rect 1608 15861 1632 16032
rect 2088 15921 2112 16032
rect 1548 15264 1572 15579
rect 1668 15441 1692 15699
rect 2088 15621 2112 15879
rect 2328 15501 2352 16119
rect 2448 16020 2472 16032
rect 2439 15981 2481 16020
rect 2568 15921 2592 16032
rect 1668 15228 1692 15399
rect 2019 15240 2061 15279
rect 2028 15228 2052 15240
rect 1548 14901 1572 15222
rect 1728 14901 1752 15132
rect 1248 14568 1272 14859
rect 948 14388 1032 14412
rect 108 13032 132 13662
rect 288 13401 312 13572
rect 108 13008 159 13032
rect 468 13041 492 13662
rect 588 13668 612 14199
rect 708 13668 732 13779
rect 408 13008 459 13032
rect 48 12948 132 12972
rect 48 10881 72 11799
rect 48 8061 72 10839
rect 108 10341 132 12948
rect 168 12021 192 13002
rect 528 12921 552 13419
rect 708 13008 732 13119
rect 768 13101 792 13572
rect 888 13461 912 13659
rect 948 13581 972 14388
rect 1008 14181 1032 14319
rect 888 13101 912 13419
rect 1008 13041 1032 14139
rect 1188 13764 1212 14436
rect 1428 14061 1452 14562
rect 1488 13881 1512 14679
rect 1659 14580 1701 14619
rect 1668 14568 1692 14580
rect 1608 14241 1632 14472
rect 1248 13401 1272 13572
rect 348 12108 372 12219
rect 768 12201 792 12912
rect 948 12261 972 13002
rect 1128 13008 1152 13119
rect 1260 13032 1299 13041
rect 1248 13008 1299 13032
rect 1260 12999 1299 13008
rect 1188 12900 1212 12912
rect 1179 12861 1221 12900
rect 1308 12732 1332 12879
rect 1368 12801 1392 13059
rect 1428 13032 1452 13719
rect 1668 13704 1692 14379
rect 1728 14181 1752 14472
rect 1848 13641 1872 14019
rect 1608 13401 1632 13536
rect 1728 13401 1752 13572
rect 1908 13521 1932 14979
rect 1968 14481 1992 15132
rect 2088 15120 2112 15132
rect 2079 15081 2121 15120
rect 2268 14901 2292 15222
rect 2328 15081 2352 15459
rect 2748 15312 2772 16239
rect 3228 16221 3252 16656
rect 3468 16641 3492 16782
rect 2808 15741 2832 16122
rect 3108 15921 3132 16032
rect 3228 15921 3252 16116
rect 2928 15501 2952 15879
rect 3288 15621 3312 16599
rect 3348 15981 3372 16299
rect 3528 16128 3552 16239
rect 3828 16164 3852 17319
rect 4128 16812 4152 17499
rect 4068 16788 4152 16812
rect 4008 16581 4032 16692
rect 4188 16581 4212 17682
rect 4248 17601 4272 17919
rect 4488 17688 4512 18099
rect 4608 17361 4632 18252
rect 4728 18021 4752 18342
rect 4908 17841 4932 18252
rect 5148 17688 5172 18216
rect 5208 18081 5232 18342
rect 5508 18141 5532 18252
rect 5628 17901 5652 18459
rect 5988 18348 6012 18579
rect 5748 18258 5772 18342
rect 5928 18240 5952 18252
rect 4668 17481 4692 17682
rect 5208 17568 5292 17592
rect 4668 17172 4692 17439
rect 4608 17148 4692 17172
rect 4608 16701 4632 17148
rect 4839 16800 4881 16839
rect 4848 16788 4872 16800
rect 5208 16788 5232 17199
rect 5268 17181 5292 17568
rect 5328 17061 5352 17859
rect 5388 17241 5412 17559
rect 5628 17481 5652 17682
rect 5688 17172 5712 17799
rect 5748 17361 5772 18216
rect 5919 18201 5961 18240
rect 6108 18201 6132 18519
rect 6228 18348 6252 18579
rect 6708 18348 6732 18579
rect 6768 18441 6792 18519
rect 6768 18411 6819 18441
rect 6780 18402 6819 18411
rect 6780 18399 6840 18402
rect 6528 18261 6552 18342
rect 6999 18360 7041 18399
rect 7008 18348 7032 18360
rect 7128 18348 7152 18519
rect 5868 17688 5892 18039
rect 6168 17541 6192 17979
rect 6408 17901 6432 18252
rect 6339 17772 6381 17799
rect 6339 17760 6399 17772
rect 6348 17748 6399 17760
rect 6408 17688 6432 17739
rect 6579 17712 6621 17739
rect 6579 17700 6672 17712
rect 6588 17688 6672 17700
rect 7188 17712 7212 18252
rect 7188 17688 7272 17712
rect 6708 17241 6732 17592
rect 6828 17481 6852 17592
rect 7248 17181 7272 17688
rect 5688 17148 5739 17172
rect 4368 16521 4392 16692
rect 4488 16581 4512 16692
rect 4968 16698 4992 16779
rect 4899 16521 4941 16539
rect 4368 16401 4392 16479
rect 5088 16461 5112 16539
rect 5139 16521 5181 16539
rect 3468 16020 3492 16032
rect 3408 15741 3432 15999
rect 3459 15981 3501 16020
rect 3468 15861 3492 15939
rect 3768 15861 3792 16032
rect 3888 15921 3912 16032
rect 2748 15288 2832 15312
rect 2808 15228 2832 15288
rect 2928 15228 2952 15459
rect 3288 15264 3312 15459
rect 3048 15228 3192 15252
rect 2628 15081 2652 15219
rect 2079 14580 2121 14619
rect 2088 14568 2112 14580
rect 2148 14361 2172 14472
rect 2208 13761 2232 14199
rect 2268 14181 2292 14472
rect 2328 14001 2352 14079
rect 1428 13008 1512 13032
rect 1308 12708 1392 12732
rect 579 12144 621 12159
rect 819 12120 861 12159
rect 828 12108 852 12120
rect 408 12000 432 12012
rect 399 11961 441 12000
rect 168 11358 192 11499
rect 348 11448 372 11739
rect 468 11448 492 11679
rect 588 11481 612 12102
rect 1188 12108 1212 12219
rect 408 10641 432 11352
rect 528 11241 552 11352
rect 168 10455 192 10599
rect 588 10548 612 10779
rect 648 10572 672 11979
rect 768 11961 792 12012
rect 768 11541 792 11919
rect 828 11448 852 11679
rect 888 11481 912 12012
rect 1008 11781 1032 12099
rect 1368 12021 1392 12708
rect 1128 11661 1152 12012
rect 1248 11841 1272 12012
rect 1428 11901 1452 12879
rect 1488 12261 1512 12819
rect 1548 12801 1572 12912
rect 1668 12900 1692 12912
rect 1659 12861 1701 12900
rect 1788 12741 1812 13479
rect 1968 13221 1992 13539
rect 1848 12861 1872 13179
rect 2208 13101 2232 13572
rect 2328 13512 2352 13659
rect 2388 13581 2412 14859
rect 2448 14481 2472 14859
rect 2628 14652 2652 15039
rect 2748 14961 2772 15132
rect 2868 14901 2892 15132
rect 2628 14628 2712 14652
rect 2688 14568 2712 14628
rect 2988 14568 3012 15039
rect 3048 14841 3072 15228
rect 3468 15141 3492 15339
rect 3228 14961 3252 15132
rect 3048 14661 3072 14799
rect 3108 14568 3252 14592
rect 2448 13701 2472 14439
rect 2748 14460 2772 14472
rect 2739 14421 2781 14460
rect 3039 14421 3081 14436
rect 2628 13941 2652 14319
rect 2268 13488 2352 13512
rect 1968 12621 1992 12912
rect 2088 12441 2112 12879
rect 2148 12741 2172 12912
rect 2268 12741 2292 13488
rect 2448 13461 2472 13539
rect 2328 12861 2352 13359
rect 2568 13161 2592 13419
rect 2928 13281 2952 13839
rect 3108 13701 3132 13779
rect 3168 13752 3192 14139
rect 3228 13821 3252 14568
rect 3348 14601 3372 15132
rect 3528 14961 3552 15579
rect 3708 15228 3732 15699
rect 4068 15381 4092 16359
rect 4419 16332 4461 16359
rect 4368 16320 4461 16332
rect 4368 16308 4452 16320
rect 4368 16128 4392 16308
rect 4188 15561 4212 16119
rect 4668 16041 4692 16119
rect 5088 16032 5112 16419
rect 5268 16281 5292 16692
rect 5388 16281 5412 16839
rect 5748 16701 5772 17139
rect 5808 16824 5832 17079
rect 5808 16521 5832 16782
rect 5868 16641 5892 16839
rect 5988 16788 6012 17019
rect 7308 17001 7332 17859
rect 7368 17721 7392 18342
rect 7428 18252 7452 18519
rect 8001 18432 8040 18441
rect 8001 18399 8052 18432
rect 7599 18360 7641 18399
rect 7608 18348 7632 18360
rect 8028 18348 8052 18399
rect 8328 18384 8352 18459
rect 8568 18348 8592 18459
rect 7428 18228 7512 18252
rect 7488 17688 7512 18228
rect 7668 17841 7692 18252
rect 8328 18252 8352 18342
rect 9288 18348 9312 18519
rect 9588 18348 9612 18579
rect 9108 18258 9132 18339
rect 8328 18228 8412 18252
rect 8148 18141 8172 18216
rect 7908 17688 7932 17799
rect 7548 17481 7572 17592
rect 7728 17541 7752 17682
rect 8268 17688 8292 18099
rect 8388 17781 8412 18228
rect 8508 17841 8532 18252
rect 8379 17700 8421 17739
rect 8388 17688 8412 17700
rect 7959 17541 8001 17556
rect 6639 16824 6681 16839
rect 5721 16479 5739 16521
rect 5928 16401 5952 16479
rect 5388 16128 5412 16239
rect 5868 16128 5892 16359
rect 6048 16341 6072 16692
rect 4428 15801 4452 15972
rect 3621 15132 3660 15141
rect 3621 15108 3672 15132
rect 3768 15120 3792 15132
rect 3621 15099 3660 15108
rect 3759 15081 3801 15120
rect 3888 15081 3912 15279
rect 3999 15240 4041 15279
rect 4008 15228 4032 15240
rect 4128 15228 4152 15459
rect 4368 15264 4392 15459
rect 4188 15120 4212 15132
rect 3288 14301 3312 14562
rect 3588 14121 3612 14559
rect 3648 14001 3672 15039
rect 3828 14568 3852 14799
rect 3948 14601 3972 14739
rect 3768 14361 3792 14472
rect 3888 14121 3912 14472
rect 4008 14421 4032 15039
rect 4068 14604 4092 15096
rect 4179 15081 4221 15120
rect 4368 14841 4392 15222
rect 4428 15081 4452 15279
rect 4068 14241 4092 14562
rect 4188 14361 4212 14472
rect 4368 14421 4392 14472
rect 4188 14181 4212 14319
rect 3168 13728 3252 13752
rect 3228 13668 3252 13728
rect 2988 13221 3012 13599
rect 2619 13140 2661 13179
rect 2628 13128 2652 13140
rect 1488 11841 1512 12102
rect 1539 11961 1581 11979
rect 1239 11460 1281 11499
rect 1248 11448 1272 11460
rect 948 11241 972 11352
rect 648 10548 699 10572
rect 228 9924 252 10419
rect 468 10428 552 10452
rect 348 9888 372 10179
rect 468 9921 492 10359
rect 108 8898 132 9879
rect 288 8988 312 9756
rect 408 9681 432 9792
rect 528 9672 552 10428
rect 708 10401 732 10539
rect 588 9732 612 9939
rect 699 9900 741 9939
rect 828 9924 852 10719
rect 1008 10548 1032 10839
rect 1068 10761 1092 11439
rect 1548 11358 1572 11619
rect 1788 11541 1812 12012
rect 1128 10548 1152 11259
rect 1308 10881 1332 11352
rect 1788 11181 1812 11352
rect 1848 10641 1872 11319
rect 1479 10584 1521 10599
rect 1599 10560 1641 10599
rect 1779 10560 1821 10599
rect 1908 10584 1932 11499
rect 1968 11481 1992 12012
rect 2088 12000 2172 12012
rect 2088 11988 2181 12000
rect 2139 11961 2181 11988
rect 2181 11928 2232 11952
rect 2028 11781 2052 11859
rect 2088 11448 2112 11799
rect 2208 11481 2232 11928
rect 2268 11772 2292 12219
rect 2328 12108 2352 12579
rect 2388 12561 2412 13059
rect 2568 13008 2592 13119
rect 2868 12921 2892 13179
rect 2988 13008 3012 13179
rect 3108 13008 3132 13539
rect 3168 13461 3192 13572
rect 3408 13281 3432 13719
rect 3468 13401 3492 13899
rect 3639 13680 3681 13719
rect 3648 13668 3672 13680
rect 3888 13701 3912 13959
rect 4068 13668 4092 14136
rect 4188 13668 4212 13899
rect 3948 13581 3972 13662
rect 4368 13581 4392 14379
rect 4488 14061 4512 15699
rect 4608 15321 4632 15579
rect 4599 15240 4641 15279
rect 4608 15228 4632 15240
rect 4728 15228 4752 15759
rect 4848 15501 4872 16032
rect 4968 15741 4992 16032
rect 5028 16008 5112 16032
rect 4668 15081 4692 15132
rect 4668 14721 4692 15039
rect 4728 14652 4752 14979
rect 4788 14961 4812 15096
rect 4968 14781 4992 15222
rect 5028 15021 5052 16008
rect 5328 15801 5352 16032
rect 5268 15264 5292 15339
rect 5121 15252 5160 15261
rect 5121 15228 5172 15252
rect 5121 15219 5160 15228
rect 5088 14721 5112 15099
rect 4668 14628 4752 14652
rect 4668 14568 4692 14628
rect 4788 14301 4812 14559
rect 5148 14481 5172 14799
rect 4908 14361 4932 14472
rect 4668 13704 4692 14259
rect 5028 14061 5052 14472
rect 3528 13341 3552 13536
rect 3288 12918 3312 13059
rect 2688 12141 2712 12399
rect 2448 11841 2472 12012
rect 2268 11748 2352 11772
rect 2268 11358 2292 11679
rect 2328 11481 2352 11748
rect 2508 11661 2532 11892
rect 2439 11460 2481 11499
rect 2568 11481 2592 11739
rect 2448 11448 2472 11460
rect 2028 11181 2052 11316
rect 1608 10548 1632 10560
rect 1788 10548 1812 10560
rect 2028 10581 2052 10659
rect 1308 10461 1332 10542
rect 1428 10092 1452 10452
rect 1848 10392 1872 10452
rect 1968 10440 1992 10452
rect 1959 10401 2001 10440
rect 1848 10368 1932 10392
rect 1908 10332 1932 10368
rect 2028 10332 2052 10419
rect 1908 10308 2052 10332
rect 1368 10068 1452 10092
rect 1128 9924 1152 10059
rect 708 9888 732 9900
rect 1248 9888 1272 9999
rect 1368 9861 1392 10068
rect 588 9708 672 9732
rect 528 9648 579 9672
rect 528 9024 552 9339
rect 408 8328 432 8679
rect 528 8481 552 8982
rect 168 7821 192 8319
rect 348 8220 372 8232
rect 339 8181 381 8220
rect 588 8232 612 9639
rect 648 9024 672 9708
rect 768 9681 792 9792
rect 819 9024 861 9039
rect 948 8988 972 9459
rect 1188 9381 1212 9756
rect 1368 9741 1392 9819
rect 1428 9561 1452 9999
rect 1608 9888 1632 10059
rect 1788 9921 1812 10299
rect 2088 10281 2112 10959
rect 2268 10632 2292 10779
rect 2328 10701 2352 11319
rect 2508 11241 2532 11352
rect 2268 10608 2352 10632
rect 2328 10548 2352 10608
rect 2508 10461 2532 10542
rect 1548 9780 1572 9792
rect 1539 9741 1581 9780
rect 1848 9798 1872 9999
rect 1788 9681 1812 9759
rect 1908 9792 1932 10239
rect 2148 10041 2172 10239
rect 2268 10221 2292 10452
rect 2568 10401 2592 11319
rect 2628 11001 2652 11799
rect 2688 11481 2712 11559
rect 2748 11481 2772 12519
rect 2808 11532 2832 12819
rect 3228 12321 3252 12699
rect 3348 12561 3372 13239
rect 3708 13221 3732 13419
rect 3828 13221 3852 13572
rect 3948 13341 3972 13539
rect 4008 13341 4032 13539
rect 4239 13512 4281 13539
rect 4188 13500 4281 13512
rect 4188 13488 4272 13500
rect 3501 13068 3579 13092
rect 3408 12888 3492 12912
rect 3408 12681 3432 12888
rect 3408 12492 3432 12639
rect 3348 12468 3432 12492
rect 3288 12081 3312 12399
rect 2808 11508 2892 11532
rect 2868 11484 2892 11508
rect 2988 11448 3012 11799
rect 3348 11721 3372 12468
rect 3468 12108 3492 12759
rect 3588 12621 3612 12912
rect 3648 12441 3672 12879
rect 3708 12741 3732 13179
rect 3999 13020 4041 13059
rect 4008 13008 4032 13020
rect 4188 12981 4212 13488
rect 4428 13461 4452 13539
rect 4488 13392 4512 13572
rect 4401 13368 4512 13392
rect 4248 12981 4272 13299
rect 4728 12981 4752 13119
rect 3828 12612 3852 12939
rect 3948 12900 3972 12912
rect 4068 12900 4092 12912
rect 3939 12861 3981 12900
rect 4059 12861 4101 12900
rect 4668 12900 4692 12915
rect 3828 12588 3879 12612
rect 3528 11952 3552 12012
rect 3468 11928 3552 11952
rect 2688 11358 2712 11439
rect 2928 11340 2952 11352
rect 2919 11301 2961 11340
rect 2688 10932 2712 11139
rect 2628 10908 2712 10932
rect 2628 10341 2652 10908
rect 2748 10584 2772 11259
rect 3108 11181 3132 11679
rect 3468 11601 3492 11928
rect 3201 11352 3240 11361
rect 3201 11328 3252 11352
rect 3201 11319 3240 11328
rect 3348 11301 3372 11352
rect 3528 11301 3552 11679
rect 2868 10701 2892 10779
rect 2868 10548 2892 10659
rect 2988 10581 3012 11019
rect 2688 10281 2712 10419
rect 2928 10440 2952 10452
rect 2919 10401 2961 10440
rect 2268 10101 2292 10179
rect 2001 9912 2040 9921
rect 2001 9888 2052 9912
rect 2001 9879 2040 9888
rect 2268 9921 2292 10059
rect 2568 9888 2592 10179
rect 2688 9921 2712 10239
rect 1908 9768 1992 9792
rect 768 8601 792 8892
rect 648 8361 672 8559
rect 828 8412 852 8679
rect 768 8388 852 8412
rect 768 8328 792 8388
rect 528 8208 612 8232
rect 48 741 72 7719
rect 108 7161 132 7539
rect 468 7461 492 8019
rect 108 6321 132 6759
rect 108 3621 132 5559
rect 168 5421 192 7239
rect 288 7161 312 7332
rect 348 7041 372 7299
rect 528 7281 552 8208
rect 648 7581 672 7899
rect 828 7701 852 8232
rect 648 7428 672 7539
rect 768 7464 792 7599
rect 579 7281 621 7299
rect 228 6801 252 6999
rect 348 6768 372 6879
rect 228 6261 252 6579
rect 288 6081 312 6573
rect 408 6381 432 6672
rect 588 6672 612 6999
rect 708 6804 732 7332
rect 888 7161 912 8019
rect 768 6921 792 7119
rect 780 6852 819 6861
rect 768 6819 819 6852
rect 648 6780 699 6792
rect 639 6768 699 6780
rect 639 6741 681 6768
rect 768 6768 792 6819
rect 888 6768 912 6999
rect 948 6861 972 8139
rect 1008 8061 1032 8439
rect 1068 8181 1092 9039
rect 1179 9000 1221 9039
rect 1188 8988 1212 9000
rect 1308 8988 1332 9459
rect 1488 8901 1512 9159
rect 1779 9000 1821 9039
rect 1908 9021 1932 9699
rect 1788 8988 1812 9000
rect 1188 8328 1212 8619
rect 1548 8601 1572 8982
rect 1728 8721 1752 8856
rect 1848 8781 1872 8892
rect 1488 8238 1512 8439
rect 1668 8364 1692 8499
rect 1368 8208 1479 8232
rect 1608 8220 1632 8232
rect 1239 8181 1281 8196
rect 1599 8181 1641 8220
rect 1548 7821 1572 8079
rect 1908 7701 1932 8799
rect 1968 7881 1992 9768
rect 2220 9792 2259 9801
rect 2208 9768 2259 9792
rect 2220 9759 2259 9768
rect 2148 9561 2172 9699
rect 2328 9501 2352 9882
rect 2508 9780 2532 9792
rect 2499 9741 2541 9780
rect 2748 9621 2772 10299
rect 3048 10221 3072 10659
rect 3228 10548 3252 10779
rect 3348 10701 3372 11259
rect 3348 10548 3372 10659
rect 3108 10440 3192 10452
rect 3099 10428 3192 10440
rect 3099 10401 3141 10428
rect 3288 10341 3312 10452
rect 3468 10221 3492 11139
rect 2988 9888 3012 10059
rect 3108 9888 3132 10059
rect 3348 9981 3372 10059
rect 3468 9981 3492 10059
rect 3468 9888 3492 9939
rect 3528 9921 3552 10779
rect 3588 10701 3612 11799
rect 3648 11358 3672 12012
rect 3768 11901 3792 12279
rect 3708 11481 3732 11799
rect 3828 11721 3852 12102
rect 3888 12021 3912 12579
rect 4008 12201 4032 12519
rect 4308 12321 4332 12876
rect 4659 12861 4701 12900
rect 4008 12108 4032 12159
rect 4128 12108 4152 12279
rect 3828 11448 3852 11559
rect 4068 11481 4092 12012
rect 4188 11532 4212 11859
rect 4248 11841 4272 12099
rect 4308 11661 4332 12159
rect 4428 12144 4452 12699
rect 4788 12681 4812 13899
rect 4848 12681 4872 14019
rect 5208 14001 5232 14859
rect 5148 13704 5172 13839
rect 4968 13281 4992 13572
rect 5088 13560 5112 13572
rect 5079 13521 5121 13560
rect 5079 13461 5121 13479
rect 5028 13008 5052 13179
rect 4608 12108 4632 12459
rect 4188 11508 4272 11532
rect 4248 11448 4272 11508
rect 4368 11448 4392 11859
rect 4488 11541 4512 11976
rect 3708 10821 3732 11319
rect 3768 10941 3792 11316
rect 4008 10701 4032 11319
rect 4068 11241 4092 11376
rect 4128 10761 4152 11319
rect 4188 11241 4212 11352
rect 3768 10584 3792 10659
rect 3888 10548 3912 10659
rect 4488 10572 4512 11436
rect 4548 11358 4572 11559
rect 4608 11241 4632 11619
rect 4668 11481 4692 11979
rect 4728 11901 4752 12519
rect 4788 12141 4812 12576
rect 4908 12312 4932 12879
rect 4968 12381 4992 12912
rect 4908 12288 4992 12312
rect 4968 12141 4992 12288
rect 5028 12012 5052 12759
rect 5088 12741 5112 12912
rect 5148 12672 5172 12879
rect 5208 12801 5232 13479
rect 5268 13461 5292 14979
rect 5328 14961 5352 15099
rect 5388 15081 5412 15939
rect 5448 15921 5472 16032
rect 5628 15981 5652 16122
rect 5808 15921 5832 16032
rect 5928 16020 5952 16032
rect 5919 15981 5961 16020
rect 5448 15261 5472 15879
rect 5808 15741 5832 15879
rect 6048 15801 6072 16122
rect 6228 15981 6252 16032
rect 6201 15948 6252 15981
rect 6201 15939 6240 15948
rect 5748 15621 5772 15699
rect 5628 15228 5652 15579
rect 6048 15228 6072 15639
rect 5568 15120 5592 15132
rect 5559 15081 5601 15120
rect 5448 14604 5472 14679
rect 5388 14232 5412 14472
rect 5688 14352 5712 15099
rect 5748 15081 5772 15222
rect 6168 15141 6192 15759
rect 6228 15681 6252 15879
rect 6348 15801 6372 16599
rect 6408 15561 6432 16479
rect 6468 15921 6492 16539
rect 6588 16521 6612 16692
rect 6708 16581 6732 16839
rect 6768 16701 6792 16839
rect 6879 16800 6921 16839
rect 6888 16788 6912 16800
rect 6948 16680 6972 16692
rect 6828 16581 6852 16659
rect 6939 16641 6981 16680
rect 7068 16581 7092 16692
rect 7188 16641 7212 16839
rect 7479 16800 7521 16839
rect 7488 16788 7512 16800
rect 6648 16128 6672 16299
rect 6768 16128 6792 16479
rect 6948 16401 6972 16536
rect 6828 16161 6852 16239
rect 6948 16164 6972 16359
rect 7188 16332 7212 16479
rect 7308 16461 7332 16692
rect 7188 16308 7272 16332
rect 7068 16128 7092 16239
rect 7248 16041 7272 16308
rect 7428 16212 7452 16692
rect 7608 16221 7632 16782
rect 7428 16188 7512 16212
rect 7488 16164 7512 16188
rect 7668 16152 7692 16839
rect 7788 16788 7812 16899
rect 7848 16521 7872 16692
rect 7608 16128 7752 16152
rect 6588 15741 6612 16032
rect 6708 15801 6732 16032
rect 5868 14568 5892 15039
rect 5928 14961 5952 15132
rect 5808 14460 5832 14472
rect 5661 14328 5712 14352
rect 5388 14208 5472 14232
rect 5388 13668 5412 14139
rect 5448 14121 5472 14208
rect 5628 13701 5652 14319
rect 5748 13881 5772 14436
rect 5799 14421 5841 14460
rect 5961 14448 6012 14472
rect 5808 14061 5832 14379
rect 5988 14361 6012 14448
rect 5688 13581 5712 13839
rect 5988 13668 6012 14199
rect 5319 13521 5361 13539
rect 5568 13461 5592 13572
rect 5448 13008 5472 13119
rect 5568 13008 5592 13239
rect 5628 13041 5652 13179
rect 4788 11841 4812 11979
rect 4848 11952 4872 12012
rect 4968 11988 5052 12012
rect 5088 12648 5172 12672
rect 4848 11928 4932 11952
rect 4788 11448 4812 11679
rect 4848 11541 4872 11859
rect 4908 11721 4932 11928
rect 4908 11481 4932 11559
rect 4428 10548 4512 10572
rect 4608 10548 4632 11019
rect 4668 10821 4692 11319
rect 4848 11121 4872 11352
rect 4659 10701 4701 10716
rect 4728 10584 4752 10659
rect 3708 10152 3732 10452
rect 3828 10341 3852 10452
rect 4128 10272 4152 10452
rect 4248 10341 4272 10452
rect 4368 10341 4392 10419
rect 4128 10248 4212 10272
rect 3708 10128 3792 10152
rect 2139 9000 2181 9039
rect 2148 8988 2172 9000
rect 2268 8988 2292 9159
rect 2388 9021 2412 9219
rect 2028 8781 2052 8979
rect 2340 8892 2379 8901
rect 2208 8541 2232 8892
rect 2328 8868 2379 8892
rect 2340 8859 2379 8868
rect 2448 8841 2472 8982
rect 2319 8340 2361 8379
rect 2328 8328 2352 8340
rect 2028 8001 2052 8319
rect 2148 7761 2172 8232
rect 2448 7881 2472 8619
rect 2508 8361 2532 9579
rect 3048 9381 3072 9792
rect 3168 9681 3192 9792
rect 3588 9780 3612 9792
rect 3579 9741 3621 9780
rect 3708 9792 3732 10059
rect 3768 10041 3792 10128
rect 3708 9768 3852 9792
rect 3579 9681 3621 9699
rect 2748 8988 2772 9099
rect 2868 9021 2892 9339
rect 3048 8988 3072 9219
rect 3180 9012 3219 9021
rect 3168 8988 3219 9012
rect 3180 8979 3219 8988
rect 3288 8901 3312 9039
rect 3648 9012 3672 9759
rect 3861 9699 3879 9741
rect 3648 8988 3732 9012
rect 2559 8841 2601 8859
rect 2688 8661 2712 8892
rect 2928 8868 3012 8892
rect 2559 8340 2601 8379
rect 2568 8328 2592 8340
rect 2688 8328 2712 8619
rect 2928 8481 2952 8868
rect 3228 8781 3252 8859
rect 2928 8361 2952 8439
rect 2628 8220 2652 8232
rect 1188 7428 1212 7539
rect 1128 7272 1152 7332
rect 1248 7320 1272 7332
rect 1068 7248 1152 7272
rect 1239 7281 1281 7320
rect 1068 7041 1092 7248
rect 588 6648 672 6672
rect 528 5901 552 6639
rect 648 6441 672 6648
rect 708 6561 732 6636
rect 828 6381 852 6672
rect 468 5868 519 5892
rect 288 5601 312 5772
rect 348 5541 372 5679
rect 408 5601 432 5772
rect 528 5241 552 5739
rect 588 5721 612 6339
rect 888 6201 912 6579
rect 888 5904 912 6039
rect 108 3321 132 3516
rect 108 2181 132 3039
rect 168 3021 192 5199
rect 588 5118 612 5679
rect 648 5241 672 5739
rect 708 5421 732 5772
rect 828 5541 852 5772
rect 768 5208 792 5319
rect 948 5301 972 5739
rect 1008 5601 1032 6519
rect 1068 5901 1092 6819
rect 1128 6678 1152 6879
rect 1188 6801 1212 6999
rect 1368 6861 1392 7419
rect 1428 7332 1452 7659
rect 1428 7308 1512 7332
rect 1428 6768 1452 7119
rect 1488 6801 1512 7308
rect 1608 7161 1632 7332
rect 1728 7041 1752 7359
rect 1848 7161 1872 7332
rect 1968 7281 1992 7332
rect 1968 7248 2019 7281
rect 1980 7239 2019 7248
rect 1548 6678 1572 6819
rect 1728 6768 1752 6999
rect 1179 5880 1221 5919
rect 1308 5904 1332 6579
rect 1368 6501 1392 6672
rect 1608 6081 1632 6639
rect 1788 6561 1812 6672
rect 1788 6381 1812 6519
rect 1188 5868 1212 5880
rect 1479 5880 1521 5919
rect 1488 5868 1512 5880
rect 1788 5778 1812 6159
rect 1128 5760 1152 5772
rect 288 4761 312 5112
rect 681 5112 720 5121
rect 681 5088 732 5112
rect 681 5079 720 5088
rect 1008 4701 1032 5199
rect 348 4308 372 4539
rect 468 4308 492 4659
rect 648 4308 672 4539
rect 768 4308 792 4479
rect 288 3741 312 4212
rect 408 4101 432 4212
rect 348 3648 372 3939
rect 828 3801 852 4212
rect 948 4101 972 4479
rect 1008 4218 1032 4659
rect 588 3558 612 3759
rect 228 2841 252 3519
rect 948 3552 972 3996
rect 1068 3981 1092 5739
rect 1119 5721 1161 5760
rect 1668 5661 1692 5772
rect 1161 5232 1200 5241
rect 1161 5208 1212 5232
rect 1308 5208 1332 5499
rect 1668 5301 1692 5619
rect 1161 5199 1200 5208
rect 1488 5118 1512 5259
rect 1128 4941 1152 5079
rect 1188 4308 1212 4779
rect 1248 4761 1272 5076
rect 1308 4581 1332 5019
rect 1248 3684 1272 4212
rect 1428 4041 1452 4659
rect 1668 4401 1692 5112
rect 1788 4821 1812 5079
rect 1668 4308 1692 4359
rect 1848 4221 1872 6039
rect 1899 5901 1941 5919
rect 1968 5904 1992 6759
rect 2028 5961 2052 6819
rect 2088 6801 2112 7299
rect 2148 7281 2172 7656
rect 2148 6768 2172 7119
rect 2208 7101 2232 7839
rect 2508 7701 2532 8199
rect 2619 8181 2661 8220
rect 2748 8121 2772 8232
rect 2868 8181 2892 8319
rect 2919 8181 2961 8199
rect 2748 8061 2772 8079
rect 2748 8028 2799 8061
rect 2760 8019 2799 8028
rect 2961 8019 2979 8061
rect 2268 7221 2292 7539
rect 2448 7428 2472 7539
rect 2388 7101 2412 7332
rect 2508 6921 2532 7332
rect 2259 6780 2301 6819
rect 2268 6768 2292 6780
rect 2508 6681 2532 6816
rect 2088 6561 2112 6639
rect 2208 6561 2232 6672
rect 2328 6441 2352 6636
rect 2568 6561 2592 7179
rect 2628 6861 2652 7779
rect 2688 7221 2712 7599
rect 2808 7428 2832 7539
rect 2928 7428 2952 7659
rect 3108 7461 3132 7599
rect 3168 7464 3192 8499
rect 3228 8061 3252 8739
rect 3288 8361 3312 8796
rect 3468 8661 3492 8892
rect 3708 8712 3732 8988
rect 3648 8688 3732 8712
rect 3408 8328 3432 8619
rect 3519 8340 3561 8379
rect 3528 8328 3552 8340
rect 3348 7641 3372 8196
rect 3468 8061 3492 8232
rect 3519 7581 3561 7599
rect 2868 7041 2892 7332
rect 3048 7281 3072 7422
rect 3288 7428 3312 7539
rect 2748 6768 2772 6999
rect 2361 6072 2400 6081
rect 2361 6060 2412 6072
rect 2361 6039 2421 6060
rect 1938 5880 1941 5901
rect 2088 5868 2112 6039
rect 2379 6021 2421 6039
rect 2628 5961 2652 6639
rect 1908 5241 1932 5739
rect 2148 5541 2172 5772
rect 2148 5208 2172 5379
rect 2268 5244 2292 5859
rect 2328 5661 2352 5919
rect 2688 5901 2712 6099
rect 2748 5781 2772 5979
rect 2388 5301 2412 5739
rect 2508 5661 2532 5772
rect 2568 5481 2592 5679
rect 2628 5118 2652 5259
rect 2088 4941 2112 5112
rect 2388 5100 2412 5112
rect 2379 5061 2421 5100
rect 1908 4428 2139 4452
rect 1908 4344 1932 4428
rect 1959 4320 2001 4359
rect 2079 4320 2121 4359
rect 1968 4308 1992 4320
rect 2088 4308 2112 4320
rect 1488 3648 1512 3879
rect 1608 3861 1632 4212
rect 828 3528 972 3552
rect 288 3201 312 3516
rect 168 2808 219 2832
rect 168 2601 192 2808
rect 339 2760 381 2799
rect 348 2748 372 2760
rect 468 2748 492 2979
rect 588 2781 612 3516
rect 759 2841 801 2859
rect 639 2760 681 2799
rect 648 2748 672 2760
rect 768 2748 792 2799
rect 108 1881 132 2139
rect 168 1998 192 2259
rect 288 2181 312 2652
rect 408 2640 432 2652
rect 399 2601 441 2640
rect 948 2658 972 2979
rect 348 2088 372 2199
rect 528 2124 552 2619
rect 828 2361 852 2652
rect 468 2088 519 2112
rect 408 1881 432 1992
rect 348 1188 372 1419
rect 459 1200 501 1239
rect 588 1221 612 2199
rect 828 2172 852 2319
rect 828 2148 912 2172
rect 648 2088 792 2112
rect 888 2088 912 2148
rect 1008 2112 1032 3639
rect 1188 3441 1212 3552
rect 1308 3261 1332 3552
rect 1188 2841 1212 3159
rect 1248 2748 1272 3039
rect 1428 2658 1452 3519
rect 1548 2748 1572 3516
rect 1668 3441 1692 3699
rect 1728 3501 1752 4179
rect 2028 4152 2052 4212
rect 1968 4128 2052 4152
rect 1908 3648 1932 3759
rect 1968 3741 1992 4128
rect 2079 4101 2121 4119
rect 2148 4101 2172 4212
rect 2061 4080 2121 4101
rect 2061 4068 2112 4080
rect 2061 4059 2100 4068
rect 2028 3648 2052 3996
rect 2268 3861 2292 5019
rect 2508 4701 2532 5112
rect 2448 4308 2472 4419
rect 2628 4218 2652 4359
rect 2388 4101 2412 4212
rect 2688 4152 2712 5739
rect 2748 4461 2772 5379
rect 2808 5241 2832 6639
rect 2868 5904 2892 6936
rect 2928 6681 2952 7239
rect 3108 6981 3132 7299
rect 3168 6804 3192 7239
rect 3228 7101 3252 7332
rect 3408 7221 3432 7539
rect 3579 7440 3621 7479
rect 3648 7461 3672 8688
rect 3708 7461 3732 8619
rect 3768 8541 3792 9579
rect 4068 9501 4092 9879
rect 4128 9432 4152 10179
rect 4068 9408 4152 9432
rect 3888 8781 3912 8892
rect 4008 8661 4032 8859
rect 4068 8832 4092 9408
rect 4128 8901 4152 9159
rect 4068 8808 4152 8832
rect 4008 8328 4032 8439
rect 3828 7881 3852 8232
rect 3948 7821 3972 8232
rect 4128 7701 4152 8808
rect 4188 8781 4212 10248
rect 4428 10221 4452 10548
rect 4548 9921 4572 10452
rect 4848 10161 4872 10779
rect 4908 10581 4932 11319
rect 4968 11001 4992 11988
rect 5088 11721 5112 12648
rect 5028 11688 5079 11712
rect 5028 11481 5052 11688
rect 5088 11448 5112 11559
rect 5148 11541 5172 12279
rect 5208 12201 5232 12696
rect 5388 12261 5412 12912
rect 5688 12741 5712 13476
rect 5748 12204 5772 13419
rect 5928 13281 5952 13572
rect 5988 13101 6012 13479
rect 6108 13452 6132 14979
rect 6228 14721 6252 15519
rect 6348 15228 6372 15339
rect 6468 15264 6492 15579
rect 6408 14961 6432 15132
rect 6588 15021 6612 15519
rect 6828 15228 6852 15819
rect 6888 15741 6912 15999
rect 6768 14961 6792 15132
rect 6888 14901 6912 15099
rect 6279 14580 6321 14619
rect 6288 14568 6312 14580
rect 6348 14181 6372 14319
rect 6408 14301 6432 14619
rect 6288 13668 6312 14079
rect 6468 13761 6492 14679
rect 6948 14652 6972 15939
rect 7008 15921 7032 16032
rect 7128 16020 7152 16032
rect 7119 15981 7161 16020
rect 7008 15201 7032 15699
rect 7008 14661 7032 15159
rect 7068 15081 7092 15279
rect 7179 15240 7221 15279
rect 7308 15261 7332 15879
rect 7188 15228 7212 15240
rect 7368 15138 7392 15999
rect 7428 15861 7452 16032
rect 7548 15981 7572 16032
rect 7548 15501 7572 15939
rect 7728 15921 7752 16128
rect 7668 15801 7692 15879
rect 7728 15381 7752 15759
rect 7788 15561 7812 16239
rect 7839 16161 7881 16179
rect 7968 16128 7992 16359
rect 8028 16221 8052 16659
rect 8088 16161 8112 16959
rect 8148 16281 8172 17679
rect 8568 17421 8592 17739
rect 8688 17688 8712 17799
rect 8928 17781 8952 18252
rect 8928 17601 8952 17739
rect 8988 17661 9012 18099
rect 9348 17952 9372 18252
rect 9681 18228 9732 18252
rect 9288 17928 9372 17952
rect 8208 16821 8232 17379
rect 8268 16788 8292 16899
rect 8388 16128 8412 16599
rect 8508 16161 8532 17139
rect 8568 16401 8592 17079
rect 8628 16641 8652 17556
rect 8748 17481 8772 17592
rect 9048 17121 9072 17559
rect 9168 17301 9192 17592
rect 9288 17301 9312 17928
rect 9459 17700 9501 17739
rect 9468 17688 9492 17700
rect 8748 16788 8772 17079
rect 8979 16824 9021 16839
rect 8808 16521 8832 16692
rect 8568 16368 8619 16401
rect 8580 16359 8619 16368
rect 7848 15801 7872 15999
rect 7941 15879 7959 15921
rect 7761 15348 7812 15372
rect 7548 15228 7572 15339
rect 7788 15261 7812 15348
rect 7848 15321 7872 15579
rect 8028 15501 8052 15996
rect 8088 15381 8112 15999
rect 8148 15621 8172 16122
rect 8328 16020 8352 16032
rect 8319 15981 8361 16020
rect 8568 16038 8592 16299
rect 8868 16041 8892 16599
rect 8988 16572 9012 16782
rect 9048 16581 9072 17079
rect 9159 16800 9201 16839
rect 9168 16788 9192 16800
rect 9288 16788 9312 16899
rect 8928 16548 9012 16572
rect 8928 16161 8952 16548
rect 8988 16128 9012 16359
rect 9108 16161 9132 16359
rect 7248 15120 7272 15132
rect 7239 15081 7281 15120
rect 7248 14961 7272 15039
rect 6888 14628 6972 14652
rect 6828 14421 6852 14559
rect 6888 14478 6912 14628
rect 7068 14568 7092 14679
rect 7188 14568 7212 14739
rect 7008 14460 7032 14472
rect 7128 14460 7152 14472
rect 6168 13521 6192 13662
rect 6108 13428 6192 13452
rect 5979 13032 6021 13059
rect 5928 13020 6021 13032
rect 5928 13008 6012 13020
rect 5868 12201 5892 12912
rect 6048 12900 6072 12912
rect 6039 12861 6081 12900
rect 5928 12621 5952 12819
rect 5319 12120 5361 12159
rect 5328 12108 5352 12120
rect 5208 11712 5232 11979
rect 5268 11781 5292 12012
rect 5361 11952 5400 11958
rect 5361 11940 5412 11952
rect 5361 11919 5421 11940
rect 5379 11901 5421 11919
rect 5508 11901 5532 11979
rect 5208 11700 5292 11712
rect 5208 11688 5301 11700
rect 5259 11661 5301 11688
rect 5208 11448 5232 11559
rect 5328 11481 5352 11799
rect 5508 11532 5532 11859
rect 5568 11841 5592 12159
rect 5619 12141 5661 12159
rect 5868 12012 5892 12159
rect 5988 12141 6012 12639
rect 6168 12381 6192 13428
rect 6228 12861 6252 13419
rect 6468 13401 6492 13572
rect 6528 13461 6552 13539
rect 6588 13521 6612 14019
rect 6408 13008 6432 13179
rect 6348 12861 6372 12912
rect 6348 12732 6372 12819
rect 6348 12708 6432 12732
rect 5808 11988 5892 12012
rect 5448 11508 5532 11532
rect 5448 11448 5472 11508
rect 5568 11448 5592 11559
rect 5688 11481 5712 11619
rect 5268 11340 5292 11352
rect 5028 11241 5052 11316
rect 5259 11301 5301 11340
rect 5121 11259 5139 11295
rect 4968 10701 4992 10896
rect 5148 10641 5172 10959
rect 5208 10761 5232 10839
rect 5268 10821 5292 11196
rect 5328 11181 5352 11319
rect 5640 11352 5679 11361
rect 5628 11328 5679 11352
rect 5640 11319 5679 11328
rect 5508 11292 5532 11316
rect 5748 11301 5772 11559
rect 5808 11541 5832 11988
rect 5868 11481 5892 11919
rect 5928 11901 5952 12102
rect 6039 12120 6081 12159
rect 6048 12108 6072 12120
rect 6288 12021 6312 12699
rect 6408 12552 6432 12708
rect 6468 12612 6492 12912
rect 6588 12741 6612 13416
rect 6468 12588 6552 12612
rect 6408 12528 6492 12552
rect 6108 11841 6132 12012
rect 6048 11448 6072 11559
rect 5508 11268 5592 11292
rect 5388 11121 5412 11199
rect 5508 11121 5532 11199
rect 5568 11172 5592 11268
rect 5568 11148 5652 11172
rect 4248 9021 4272 9399
rect 4368 9381 4392 9792
rect 4488 9024 4512 9579
rect 4428 8781 4452 8892
rect 4461 8748 4512 8772
rect 4488 8421 4512 8748
rect 4548 8421 4572 8859
rect 4608 8412 4632 10119
rect 4668 9921 4692 9999
rect 4848 9921 4872 9999
rect 4800 9912 4839 9921
rect 4788 9888 4839 9912
rect 4800 9879 4839 9888
rect 4668 8841 4692 9759
rect 4908 9441 4932 10419
rect 4968 10341 4992 10416
rect 5148 10401 5172 10599
rect 5208 10521 5232 10719
rect 5448 10548 5472 11019
rect 5628 11001 5652 11148
rect 5559 10701 5601 10719
rect 5208 10341 5232 10479
rect 4968 9981 4992 10299
rect 5139 9900 5181 9939
rect 5148 9888 5172 9900
rect 5268 9888 5292 9999
rect 5328 9921 5352 10359
rect 5388 10341 5412 10452
rect 5508 10392 5532 10416
rect 5448 10368 5532 10392
rect 4968 9621 4992 9876
rect 5061 9768 5112 9792
rect 5028 9561 5052 9759
rect 5088 9441 5112 9699
rect 5148 9381 5172 9639
rect 5208 9621 5232 9792
rect 4848 9141 4872 9219
rect 5028 9201 5052 9279
rect 4848 8988 4872 9099
rect 4959 9000 5001 9039
rect 5088 9021 5112 9159
rect 4968 8988 4992 9000
rect 5139 9000 5181 9039
rect 5148 8988 5172 9000
rect 5268 8988 5292 9219
rect 5328 9201 5352 9759
rect 5388 9621 5412 9939
rect 5448 9081 5472 10368
rect 5628 10341 5652 10959
rect 5688 10581 5712 10779
rect 5808 10761 5832 11436
rect 5868 11121 5892 11319
rect 6108 11340 6132 11352
rect 6099 11301 6141 11340
rect 5748 10572 5772 10719
rect 5868 10641 5892 10839
rect 5748 10548 5832 10572
rect 5928 10548 5952 10899
rect 6168 10581 6192 11319
rect 6228 11301 6252 11979
rect 6288 11301 6312 11859
rect 6348 11181 6372 12339
rect 6399 12141 6441 12159
rect 6468 12144 6492 12528
rect 6528 12381 6552 12588
rect 6648 12201 6672 13719
rect 6768 13668 6792 14199
rect 6888 13881 6912 14436
rect 6999 14421 7041 14460
rect 7119 14421 7161 14460
rect 6888 13461 6912 13572
rect 6888 13008 6912 13239
rect 6768 12441 6792 12912
rect 6768 12108 6792 12336
rect 7008 12261 7032 13959
rect 7068 13704 7092 14079
rect 7188 14001 7212 14199
rect 7248 14121 7272 14439
rect 7308 14181 7332 14679
rect 7128 13668 7152 13779
rect 7308 13701 7332 13839
rect 7368 13641 7392 15096
rect 7428 14781 7452 15099
rect 7608 14781 7632 15132
rect 7548 14568 7572 14739
rect 7788 14661 7812 14739
rect 7848 14721 7872 15216
rect 7848 14481 7872 14616
rect 7839 14421 7881 14439
rect 7608 14301 7632 14412
rect 7608 13821 7632 14259
rect 7848 13641 7872 13779
rect 7248 13548 7332 13572
rect 7068 13041 7092 13479
rect 7308 13332 7332 13548
rect 7368 13401 7392 13599
rect 7308 13308 7419 13332
rect 7608 13281 7632 13452
rect 7248 13041 7272 13179
rect 7308 13101 7332 13239
rect 7368 13041 7392 13119
rect 7308 13008 7359 13032
rect 7068 12912 7092 12999
rect 7488 12981 7512 13239
rect 7908 13221 7932 15339
rect 8001 15132 8040 15141
rect 8001 15108 8052 15132
rect 8001 15099 8040 15108
rect 8061 14652 8100 14661
rect 8061 14619 8112 14652
rect 8088 14568 8112 14619
rect 8208 14601 8232 15099
rect 8268 14652 8292 15519
rect 8328 15141 8352 15639
rect 8508 15321 8532 15999
rect 8748 16020 8772 16032
rect 8619 15972 8661 15999
rect 8739 15981 8781 16020
rect 8619 15960 8712 15972
rect 8628 15948 8712 15960
rect 8628 15228 8652 15819
rect 8688 15801 8712 15948
rect 8748 15141 8772 15579
rect 8268 14628 8352 14652
rect 8268 14478 8292 14559
rect 7968 13341 7992 13779
rect 8088 13668 8112 13959
rect 8208 13941 8232 14439
rect 7068 12888 7152 12912
rect 7128 12681 7152 12888
rect 6888 12108 6912 12219
rect 7059 12132 7101 12159
rect 7041 12120 7101 12132
rect 7041 12108 7092 12120
rect 6528 11988 6612 12012
rect 6408 11481 6432 11859
rect 6528 11448 6552 11619
rect 6588 11481 6612 11988
rect 6648 11541 6672 12096
rect 6708 11481 6732 11739
rect 6828 11661 6852 12012
rect 6948 11952 6972 12012
rect 6948 11928 6999 11952
rect 6468 11340 6492 11352
rect 6459 11301 6501 11340
rect 6618 11316 6621 11340
rect 6579 11295 6621 11316
rect 6579 11280 6639 11295
rect 6588 11268 6639 11280
rect 6288 10548 6312 11139
rect 6408 11121 6432 11259
rect 6600 11253 6639 11268
rect 5508 9921 5532 10299
rect 5688 10161 5712 10476
rect 5628 9888 5652 10059
rect 5808 9921 5832 10239
rect 5988 10161 6012 10452
rect 6108 10281 6132 10539
rect 6159 10401 6201 10419
rect 6048 10101 6072 10179
rect 6048 9924 6072 9996
rect 6168 9981 6192 10359
rect 6228 10221 6252 10452
rect 6348 10440 6372 10452
rect 6339 10401 6381 10440
rect 6408 10341 6432 10419
rect 6468 9981 6492 10959
rect 6588 10548 6612 10719
rect 6768 10632 6792 11499
rect 6828 11361 6852 11619
rect 7008 11481 7032 11919
rect 7068 11484 7092 11979
rect 7128 11961 7152 12639
rect 7188 12201 7212 12912
rect 7248 12132 7272 12879
rect 7488 12801 7512 12939
rect 7968 12861 7992 13299
rect 8028 13041 8052 13179
rect 8088 13101 8112 13299
rect 8208 13281 8232 13572
rect 8148 13008 8172 13179
rect 8208 13161 8232 13239
rect 8268 13092 8292 13539
rect 8328 13221 8352 14628
rect 8388 14481 8412 14679
rect 8448 14601 8472 15039
rect 8508 14901 8532 15132
rect 8808 15132 8832 15759
rect 8928 15561 8952 15999
rect 9048 15741 9072 16032
rect 9108 15612 9132 15999
rect 9168 15681 9192 16539
rect 9228 16401 9252 16692
rect 9408 16461 9432 16899
rect 9528 16824 9552 17556
rect 9588 16788 9612 17439
rect 9708 17421 9732 18228
rect 9708 17061 9732 17259
rect 9708 16788 9732 17019
rect 9768 16941 9792 18579
rect 9888 18261 9912 18399
rect 9999 18360 10041 18399
rect 10008 18348 10032 18360
rect 10128 18348 10152 18519
rect 10608 18348 10632 18579
rect 10068 17841 10092 18252
rect 10188 18141 10212 18252
rect 10368 18141 10392 18342
rect 9828 17361 9852 17799
rect 10488 17688 10512 17919
rect 10548 17781 10572 18252
rect 10668 17601 10692 17979
rect 10728 17961 10752 18342
rect 10908 18141 10932 18252
rect 11148 18141 11172 18459
rect 11448 18348 11472 18459
rect 11268 17961 11292 18252
rect 10839 17700 10881 17739
rect 10848 17688 10872 17700
rect 11028 17661 11052 17739
rect 11181 17712 11220 17721
rect 11181 17688 11232 17712
rect 11328 17688 11352 18039
rect 11388 18021 11412 18252
rect 11181 17679 11220 17688
rect 10008 16824 10032 17199
rect 10068 17001 10092 17493
rect 10188 17481 10212 17592
rect 10128 16788 10152 17139
rect 9528 16221 9552 16479
rect 9399 16140 9441 16179
rect 9519 16161 9561 16179
rect 9408 16128 9432 16140
rect 9588 16041 9612 16239
rect 9288 15861 9312 16032
rect 9528 15741 9552 15999
rect 9579 15981 9621 15999
rect 9648 15861 9672 16299
rect 9108 15588 9192 15612
rect 8928 15264 8952 15456
rect 9048 15264 9072 15519
rect 8808 15108 8892 15132
rect 8508 14604 8532 14679
rect 8388 13701 8412 14376
rect 8688 14241 8712 14472
rect 8388 13161 8412 13299
rect 8268 13080 8412 13092
rect 8268 13068 8421 13080
rect 8379 13041 8421 13068
rect 8448 13032 8472 13479
rect 8628 13401 8652 13899
rect 8688 13701 8712 14199
rect 8748 13761 8772 14079
rect 8808 13941 8832 14919
rect 8868 14901 8892 15108
rect 9168 15132 9192 15588
rect 9348 15228 9372 15459
rect 9468 15228 9492 15459
rect 9168 15108 9252 15132
rect 9168 14901 9192 15039
rect 8988 14568 9012 14679
rect 9168 14601 9192 14679
rect 8928 14460 8952 14472
rect 8919 14421 8961 14460
rect 8841 13812 8880 13821
rect 8841 13800 8892 13812
rect 8841 13779 8901 13800
rect 8859 13761 8901 13779
rect 8781 13752 8820 13761
rect 8781 13719 8832 13752
rect 8808 13668 8832 13719
rect 8928 13668 8952 14379
rect 9048 14181 9072 14472
rect 9108 14121 9132 14379
rect 9048 13578 9072 13719
rect 8688 13092 8712 13539
rect 8748 13161 8772 13419
rect 9108 13341 9132 14079
rect 9228 14001 9252 15108
rect 9288 14472 9312 15096
rect 9408 14781 9432 15132
rect 9528 14841 9552 15096
rect 9588 14721 9612 15219
rect 9648 15081 9672 15699
rect 9708 15261 9732 16419
rect 9828 16341 9852 16779
rect 9879 16140 9921 16179
rect 10008 16161 10032 16539
rect 10068 16461 10092 16692
rect 9888 16128 9912 16140
rect 9828 16020 9852 16032
rect 9768 15672 9792 15999
rect 9819 15981 9861 16020
rect 9939 15981 9981 15996
rect 9768 15648 9852 15672
rect 9768 15228 9792 15579
rect 9828 15441 9852 15648
rect 10008 15228 10032 15699
rect 10068 15681 10092 16356
rect 10128 16041 10152 16179
rect 10188 16161 10212 16419
rect 10248 16221 10272 17379
rect 10428 17361 10452 17592
rect 11088 17598 11112 17679
rect 10308 16641 10332 16959
rect 10548 16788 10572 16959
rect 10668 16824 10692 17439
rect 10788 17361 10812 17592
rect 10908 17352 10932 17556
rect 10848 17328 10932 17352
rect 10488 16680 10512 16692
rect 10479 16641 10521 16680
rect 10308 16128 10332 16599
rect 10488 16521 10512 16599
rect 10428 16128 10452 16479
rect 10488 16221 10512 16416
rect 10608 16401 10632 16692
rect 10608 16161 10632 16239
rect 10668 16128 10692 16599
rect 10728 16461 10752 16659
rect 10788 16401 10812 17256
rect 10848 16272 10872 17328
rect 10968 16788 10992 17319
rect 11028 17001 11052 17556
rect 11268 17532 11292 17592
rect 11208 17508 11292 17532
rect 11088 16824 11112 17139
rect 10908 16572 10932 16659
rect 10908 16548 10959 16572
rect 10908 16341 10932 16476
rect 10848 16248 10932 16272
rect 10908 16161 10932 16248
rect 9948 15120 9972 15132
rect 9939 15081 9981 15120
rect 9288 14448 9372 14472
rect 9408 14460 9432 14472
rect 9528 14460 9552 14472
rect 9288 13701 9312 13779
rect 9348 13668 9372 14448
rect 9399 14421 9441 14460
rect 9519 14421 9561 14460
rect 9588 14352 9612 14436
rect 9648 14361 9672 14859
rect 9528 14328 9612 14352
rect 8688 13068 8772 13092
rect 8448 13008 8532 13032
rect 7188 12108 7272 12132
rect 7308 12108 7332 12399
rect 7428 12201 7452 12279
rect 7419 12120 7461 12159
rect 7428 12108 7452 12120
rect 6828 10761 6852 11319
rect 7008 11241 7032 11319
rect 6768 10608 6852 10632
rect 6828 10548 6852 10608
rect 6888 10581 6912 11199
rect 6648 10392 6672 10452
rect 6768 10440 6792 10452
rect 6759 10401 6801 10440
rect 6648 10368 6732 10392
rect 6708 10272 6732 10368
rect 6759 10341 6801 10359
rect 6708 10248 6819 10272
rect 6888 10272 6912 10419
rect 6861 10248 6912 10272
rect 4668 8481 4692 8619
rect 4608 8388 4692 8412
rect 4419 8340 4461 8379
rect 4428 8328 4452 8340
rect 4608 8241 4632 8319
rect 4248 8061 4272 8232
rect 4368 8121 4392 8232
rect 3759 7461 3801 7479
rect 3588 7428 3612 7440
rect 4059 7440 4101 7479
rect 4068 7428 4092 7440
rect 3288 7101 3312 7179
rect 3108 6660 3132 6672
rect 3099 6621 3141 6660
rect 3108 6201 3132 6579
rect 3228 6561 3252 6672
rect 3348 6501 3372 7119
rect 3468 6972 3492 7119
rect 3528 6981 3552 7332
rect 3708 7161 3732 7356
rect 3861 7332 3900 7341
rect 3861 7308 3912 7332
rect 3861 7299 3900 7308
rect 4128 7221 4152 7299
rect 3408 6948 3492 6972
rect 3408 6801 3432 6948
rect 3501 6888 3579 6912
rect 3828 6678 3852 6939
rect 4008 6804 4032 6999
rect 4128 6768 4152 7179
rect 4188 7041 4212 7719
rect 4248 6981 4272 7539
rect 4308 6861 4332 7479
rect 4479 7440 4521 7479
rect 4488 7428 4512 7440
rect 4608 7428 4632 8136
rect 4668 7761 4692 8388
rect 4728 8361 4752 8859
rect 4788 8481 4812 8892
rect 4908 8880 4932 8892
rect 4899 8841 4941 8880
rect 4848 8412 4872 8559
rect 4908 8481 4932 8619
rect 4821 8388 4872 8412
rect 4788 8328 4812 8376
rect 4719 8172 4761 8199
rect 4719 8160 4812 8172
rect 4728 8148 4812 8160
rect 4428 7101 4452 7332
rect 4548 7320 4572 7332
rect 4539 7281 4581 7320
rect 4368 6792 4392 6999
rect 4308 6768 4392 6792
rect 4479 6780 4521 6819
rect 4488 6768 4512 6780
rect 3468 6561 3492 6672
rect 3588 6501 3612 6672
rect 3828 6501 3852 6636
rect 3948 6561 3972 6636
rect 2988 5868 3012 5979
rect 3948 5961 3972 6339
rect 4068 6141 4092 6672
rect 3099 5904 3141 5919
rect 3048 5712 3072 5736
rect 2988 5688 3072 5712
rect 2868 5208 2892 5379
rect 2988 5244 3012 5688
rect 3228 5661 3252 5919
rect 3459 5880 3501 5919
rect 3468 5868 3492 5880
rect 3948 5868 3972 5919
rect 4068 5901 4092 6099
rect 3408 5712 3432 5772
rect 3408 5688 3492 5712
rect 3228 5208 3252 5439
rect 3048 5100 3072 5112
rect 3039 5061 3081 5100
rect 3408 5061 3432 5619
rect 3468 5412 3492 5688
rect 3708 5472 3732 5862
rect 3708 5448 3759 5472
rect 3468 5388 3552 5412
rect 2988 4701 3012 4779
rect 2859 4320 2901 4359
rect 2868 4308 2892 4320
rect 2988 4308 3012 4659
rect 2628 4128 2712 4152
rect 2148 3558 2172 3819
rect 2448 3648 2472 3759
rect 2568 3681 2592 3879
rect 1668 2748 1692 3399
rect 1068 2361 1092 2619
rect 1188 2301 1212 2652
rect 1308 2541 1332 2652
rect 1848 2541 1872 3453
rect 1548 2328 1692 2352
rect 1008 2088 1092 2112
rect 648 1281 672 2088
rect 1068 1998 1092 2088
rect 828 1761 852 1992
rect 1248 1980 1272 1992
rect 1068 1881 1092 1956
rect 1239 1941 1281 1980
rect 1368 1881 1392 1992
rect 468 1188 492 1200
rect 621 1188 672 1212
rect 768 1188 792 1419
rect 288 861 312 1092
rect 708 981 732 1092
rect 288 528 312 699
rect 408 528 432 819
rect 828 741 852 1092
rect 948 981 972 1239
rect 1248 1188 1272 1479
rect 1488 1341 1512 2079
rect 1479 1281 1521 1299
rect 1359 1200 1401 1239
rect 1548 1224 1572 2328
rect 1608 2121 1632 2259
rect 1668 2241 1692 2328
rect 1728 2088 1752 2319
rect 1848 2088 1872 2199
rect 1908 2121 1932 2799
rect 1788 1980 1812 1992
rect 1779 1941 1821 1980
rect 1788 1761 1812 1899
rect 1368 1188 1392 1200
rect 1668 1188 1692 1479
rect 1188 981 1212 1092
rect 768 528 792 639
rect 828 561 852 699
rect 1188 621 1212 939
rect 1608 921 1632 1092
rect 1248 564 1272 699
rect 1488 528 1512 819
rect 1608 528 1632 759
rect 948 201 972 519
rect 1428 420 1452 432
rect 1548 420 1572 432
rect 1419 381 1461 420
rect 1539 381 1581 420
rect 1728 381 1752 1056
rect 1848 921 1872 1299
rect 1908 1101 1932 1182
rect 1968 1041 1992 3399
rect 2208 2748 2232 3639
rect 2508 3261 2532 3516
rect 2628 3441 2652 4128
rect 2808 4101 2832 4212
rect 2868 3648 2892 4119
rect 2928 3801 2952 4212
rect 2808 3540 2832 3552
rect 2799 3501 2841 3540
rect 2568 3201 2592 3279
rect 2328 2661 2352 2859
rect 2559 2760 2601 2799
rect 2568 2748 2592 2760
rect 2148 2301 2172 2652
rect 2808 2658 2832 3459
rect 2928 3141 2952 3552
rect 2868 3108 2919 3132
rect 2628 2541 2652 2652
rect 2268 2088 2292 2199
rect 2388 2088 2412 2319
rect 2448 2121 2472 2499
rect 2808 2361 2832 2616
rect 2868 2601 2892 3108
rect 2988 3021 3012 3519
rect 3048 3501 3072 3999
rect 3108 3921 3132 4779
rect 3168 4161 3192 4419
rect 3228 3981 3252 4539
rect 3468 4461 3492 5319
rect 3528 4581 3552 5388
rect 3648 5208 3672 5319
rect 3768 5208 3792 5439
rect 3888 5241 3912 5772
rect 4128 5661 4152 6579
rect 4188 6501 4212 6672
rect 4308 6621 4332 6768
rect 4668 6681 4692 7059
rect 4188 5901 4212 6219
rect 4248 5868 4272 6159
rect 4368 5868 4392 6099
rect 4428 6021 4452 6636
rect 4608 6441 4632 6639
rect 4728 6201 4752 7659
rect 4788 7641 4812 8148
rect 4908 7941 4932 8199
rect 4968 8121 4992 8499
rect 5028 8181 5052 8679
rect 5088 8241 5112 8859
rect 5148 8481 5172 8799
rect 5208 8781 5232 8892
rect 5328 8421 5352 8892
rect 5448 8841 5472 8976
rect 5508 8721 5532 9759
rect 5568 9441 5592 9792
rect 5868 9792 5892 9882
rect 5868 9768 5952 9792
rect 5568 9021 5592 9279
rect 5688 8988 5712 9099
rect 5748 9081 5772 9279
rect 5808 9141 5832 9759
rect 5748 9045 5799 9081
rect 5760 9039 5799 9045
rect 5868 9021 5892 9339
rect 5628 8661 5652 8892
rect 5928 8892 5952 9768
rect 6168 9780 6192 9792
rect 6159 9741 6201 9780
rect 6219 9732 6261 9759
rect 6348 9741 6372 9792
rect 6219 9720 6312 9732
rect 6228 9708 6312 9720
rect 6348 9708 6399 9741
rect 6048 9501 6072 9699
rect 5868 8868 5952 8892
rect 5868 8841 5892 8868
rect 5328 8388 5379 8421
rect 5340 8382 5379 8388
rect 5181 8352 5220 8361
rect 5181 8328 5232 8352
rect 5181 8319 5220 8328
rect 5739 8340 5781 8379
rect 5748 8328 5772 8340
rect 4968 7428 4992 7719
rect 5088 7464 5112 7779
rect 4908 7320 4932 7332
rect 4899 7281 4941 7320
rect 5028 7161 5052 7332
rect 4788 6501 4812 7119
rect 5088 7041 5112 7299
rect 5148 7281 5172 7479
rect 5208 7221 5232 8139
rect 5508 8121 5532 8322
rect 5568 8001 5592 8259
rect 5481 7788 5559 7812
rect 5421 7728 5532 7752
rect 5268 7461 5292 7599
rect 5448 7581 5472 7659
rect 5508 7641 5532 7728
rect 5319 7440 5361 7479
rect 5328 7428 5352 7440
rect 5388 7320 5412 7332
rect 4968 6921 4992 6999
rect 4899 6780 4941 6819
rect 4908 6768 4932 6780
rect 5028 6768 5052 6879
rect 5088 6801 5112 6936
rect 5208 6921 5232 7116
rect 5268 6921 5292 7296
rect 5379 7281 5421 7320
rect 5628 7221 5652 8139
rect 5688 8121 5712 8232
rect 5688 7461 5712 7959
rect 5748 7464 5772 7779
rect 5868 7641 5892 8799
rect 5928 8361 5952 8799
rect 5988 8421 6012 9099
rect 6048 9021 6072 9459
rect 6099 9081 6141 9099
rect 6168 8988 6192 9579
rect 6228 9201 6252 9639
rect 6288 9321 6312 9708
rect 6360 9699 6399 9708
rect 6348 9021 6372 9579
rect 6468 9501 6492 9792
rect 6528 9561 6552 9759
rect 6588 9741 6612 9999
rect 6648 9381 6672 10179
rect 6768 10101 6792 10179
rect 6948 10161 6972 11139
rect 7008 10041 7032 11079
rect 7128 10941 7152 11259
rect 7188 11241 7212 12108
rect 7368 11481 7392 12012
rect 7548 11541 7572 12819
rect 8088 12681 8112 12879
rect 8208 12801 8232 12912
rect 7608 11721 7632 12519
rect 7728 12501 7752 12579
rect 7839 12120 7881 12159
rect 7908 12141 7932 12339
rect 7968 12321 7992 12639
rect 8061 12279 8079 12321
rect 7848 12108 7872 12120
rect 7968 11721 7992 12159
rect 7839 11661 7881 11679
rect 7860 11598 7920 11601
rect 7419 11460 7461 11499
rect 7428 11448 7452 11460
rect 7668 11448 7692 11559
rect 7881 11559 7899 11598
rect 7068 10581 7092 10899
rect 7128 10548 7152 10719
rect 7248 10581 7272 11019
rect 7308 11001 7332 11352
rect 6828 9888 6852 9999
rect 6708 9621 6732 9759
rect 6768 9501 6792 9792
rect 6948 9621 6972 9792
rect 6408 8952 6432 9279
rect 6348 8928 6432 8952
rect 6108 8880 6132 8892
rect 6099 8841 6141 8880
rect 6048 8328 6072 8619
rect 6288 8592 6312 8859
rect 6228 8568 6312 8592
rect 6168 8481 6192 8559
rect 6048 8061 6072 8139
rect 5859 7440 5901 7479
rect 5868 7428 5892 7440
rect 5340 6912 5379 6921
rect 5328 6879 5379 6912
rect 5328 6804 5352 6879
rect 5448 6768 5472 6939
rect 5568 6861 5592 7119
rect 5628 6801 5652 6999
rect 5688 6801 5712 7299
rect 5748 7041 5772 7239
rect 5808 7221 5832 7332
rect 4848 6441 4872 6639
rect 5148 6561 5172 6762
rect 5799 6780 5841 6819
rect 5868 6801 5892 7119
rect 5928 7101 5952 7299
rect 5988 6852 6012 7359
rect 6048 7341 6072 8019
rect 6108 7881 6132 8232
rect 6228 7821 6252 8568
rect 6288 8361 6312 8499
rect 6348 8361 6372 8928
rect 6408 8481 6432 8859
rect 6468 8661 6492 9279
rect 6528 9021 6552 9099
rect 6588 8988 6612 9219
rect 6828 9201 6852 9579
rect 6948 9321 6972 9516
rect 7008 9252 7032 9699
rect 7068 9561 7092 10359
rect 7308 10161 7332 10779
rect 7128 9981 7152 10119
rect 7188 9921 7212 10119
rect 7368 10101 7392 11259
rect 7428 10692 7452 10839
rect 7488 10821 7512 11319
rect 7608 11121 7632 11352
rect 7428 10668 7512 10692
rect 7488 10548 7512 10668
rect 7668 10581 7692 11259
rect 7728 11241 7752 11352
rect 7728 10641 7752 11199
rect 7908 10992 7932 11439
rect 7968 11301 7992 11616
rect 7908 10968 7992 10992
rect 7608 10548 7659 10572
rect 7908 10572 7932 10899
rect 7968 10821 7992 10968
rect 8028 10881 8052 12216
rect 8148 12108 8172 12459
rect 8328 12141 8352 12912
rect 8088 11601 8112 11976
rect 8319 11961 8361 11979
rect 8088 11481 8112 11559
rect 8139 11541 8181 11559
rect 8139 11460 8181 11499
rect 8148 11448 8172 11460
rect 8268 11448 8292 11619
rect 8388 11601 8412 12819
rect 8448 12201 8472 12879
rect 8499 12261 8541 12279
rect 8499 12240 8559 12261
rect 8508 12228 8559 12240
rect 8520 12219 8559 12228
rect 8628 12132 8652 12519
rect 8688 12501 8712 12999
rect 8628 12108 8712 12132
rect 8448 11988 8499 12012
rect 8388 11361 8412 11496
rect 8448 11481 8472 11988
rect 8628 11901 8652 11979
rect 8688 11541 8712 12108
rect 8748 12021 8772 13068
rect 8808 13041 8832 13299
rect 9168 13032 9192 13239
rect 9168 13008 9252 13032
rect 8880 12912 8919 12921
rect 8868 12888 8919 12912
rect 8880 12879 8919 12888
rect 9048 12801 9072 12912
rect 9408 12612 9432 13479
rect 9348 12588 9432 12612
rect 8868 12141 8892 12579
rect 9048 12108 9072 12459
rect 8808 11892 8832 12099
rect 8748 11868 8832 11892
rect 8748 11661 8772 11868
rect 8748 11472 8772 11619
rect 8688 11448 8772 11472
rect 7908 10548 8052 10572
rect 7548 10440 7572 10452
rect 7428 9921 7452 10419
rect 7539 10401 7581 10440
rect 7728 10341 7752 10479
rect 8028 10452 8052 10548
rect 7479 10041 7521 10059
rect 7128 9441 7152 9876
rect 7248 9780 7272 9792
rect 7188 9681 7212 9759
rect 7239 9741 7281 9780
rect 6948 9228 7032 9252
rect 6888 8988 6912 9099
rect 6948 9081 6972 9228
rect 6528 8781 6552 8859
rect 6528 8421 6552 8559
rect 6588 8472 6612 8799
rect 6648 8541 6672 8892
rect 6699 8781 6741 8799
rect 6588 8448 6672 8472
rect 6528 8328 6552 8379
rect 6048 6921 6072 7059
rect 5988 6828 6039 6852
rect 5808 6768 5832 6780
rect 5241 6672 5280 6681
rect 5241 6648 5292 6672
rect 5388 6660 5412 6672
rect 5241 6639 5280 6648
rect 5379 6621 5421 6660
rect 4608 5904 4632 6159
rect 4788 6141 4812 6219
rect 4848 6141 4872 6336
rect 4968 6201 4992 6519
rect 4968 6081 4992 6159
rect 4728 5868 4752 6039
rect 5028 6012 5052 6399
rect 5148 6021 5172 6279
rect 4968 5988 5052 6012
rect 4968 5868 4992 5988
rect 3288 4341 3312 4419
rect 3399 4320 3441 4359
rect 3588 4344 3612 5079
rect 3828 5001 3852 5112
rect 3948 4641 3972 5619
rect 4008 5181 4032 5259
rect 4188 5208 4212 5379
rect 4308 5301 4332 5772
rect 4488 5361 4512 5859
rect 4128 5001 4152 5112
rect 3699 4401 3741 4419
rect 3408 4308 3432 4320
rect 3528 4308 3579 4332
rect 3708 4308 3732 4359
rect 3168 3948 3219 3972
rect 3108 2841 3132 3639
rect 3168 3501 3192 3948
rect 3288 3861 3312 4179
rect 3348 4041 3372 4212
rect 3468 4200 3492 4212
rect 3768 4200 3792 4212
rect 3459 4161 3501 4200
rect 3759 4161 3801 4200
rect 3408 3648 3432 3819
rect 3039 2784 3081 2799
rect 3168 2748 3192 2979
rect 3228 2961 3252 3519
rect 3348 3261 3372 3552
rect 3468 3540 3492 3552
rect 3459 3501 3501 3540
rect 3588 3501 3612 3819
rect 3768 3648 3792 3939
rect 3888 3801 3912 4212
rect 4008 4161 4032 4419
rect 3708 3540 3732 3552
rect 3699 3501 3741 3540
rect 3828 3381 3852 3552
rect 3828 3261 3852 3339
rect 3228 2841 3252 2919
rect 3588 2841 3612 2979
rect 2028 1941 2052 2079
rect 2328 1881 2352 1992
rect 2508 1761 2532 2199
rect 2388 1101 2412 1419
rect 2568 1401 2592 2199
rect 2988 2124 3012 2652
rect 3108 2640 3132 2652
rect 3099 2601 3141 2640
rect 3288 2421 3312 2799
rect 3459 2760 3501 2799
rect 3579 2760 3621 2799
rect 3468 2748 3492 2760
rect 3588 2748 3612 2760
rect 3708 2658 3732 2919
rect 3888 2748 3912 2859
rect 3948 2841 3972 3519
rect 4008 3141 4032 3759
rect 4068 3501 4092 3879
rect 4128 3558 4152 4419
rect 4248 4308 4272 4779
rect 4308 4461 4332 5139
rect 4368 4461 4392 5319
rect 4608 5208 4632 5619
rect 4668 5481 4692 5772
rect 4728 5241 4752 5379
rect 4548 4941 4572 5112
rect 4788 4761 4812 5439
rect 4848 5361 4872 5862
rect 4848 5001 4872 5256
rect 4908 5241 4932 5739
rect 4968 5208 4992 5439
rect 5028 5421 5052 5772
rect 5208 5772 5232 6459
rect 5268 5901 5292 6579
rect 5448 5952 5472 6579
rect 5508 6321 5532 6672
rect 5388 5928 5472 5952
rect 5388 5868 5412 5928
rect 5499 5880 5541 5919
rect 5568 5901 5592 6639
rect 5508 5868 5532 5880
rect 5208 5748 5352 5772
rect 5088 5481 5112 5619
rect 5148 5601 5172 5739
rect 5328 5712 5352 5748
rect 5328 5688 5412 5712
rect 5079 5220 5121 5259
rect 5268 5241 5292 5679
rect 5388 5601 5412 5688
rect 5088 5208 5112 5220
rect 4368 4419 4419 4461
rect 4368 4308 4392 4419
rect 4488 4401 4512 4599
rect 4908 4581 4932 5079
rect 5148 5100 5172 5112
rect 5139 5061 5181 5100
rect 4548 4218 4572 4479
rect 4668 4308 4692 4539
rect 4788 4308 4812 4479
rect 4848 4401 4872 4539
rect 4728 4200 4752 4212
rect 4401 4119 4419 4161
rect 4548 3801 4572 4176
rect 4719 4161 4761 4200
rect 4641 4119 4659 4161
rect 4668 3648 4692 3879
rect 4848 3792 4872 4176
rect 4848 3768 4932 3792
rect 4848 3621 4872 3699
rect 4368 3540 4392 3552
rect 4248 3321 4272 3516
rect 4359 3501 4401 3540
rect 4428 3381 4452 3519
rect 4548 3321 4572 3552
rect 4008 2901 4032 3099
rect 4728 2961 4752 3552
rect 4161 2928 4212 2952
rect 4128 2784 4152 2919
rect 3288 2088 3312 2199
rect 2628 1641 2652 1959
rect 2988 1992 3012 2082
rect 2748 1821 2772 1956
rect 2868 1761 2892 1992
rect 2988 1968 3132 1992
rect 3228 1761 3252 1992
rect 2628 1272 2652 1599
rect 3408 1581 3432 2079
rect 3468 1881 3492 2379
rect 3528 2241 3552 2652
rect 3708 2124 3732 2199
rect 3819 2121 3861 2139
rect 3888 1998 3912 2199
rect 4068 2124 4092 2652
rect 4188 2541 4212 2928
rect 4701 2799 4719 2841
rect 4479 2760 4521 2799
rect 4488 2748 4512 2760
rect 4848 2781 4872 3219
rect 4908 3081 4932 3768
rect 4908 2784 4932 2859
rect 4968 2841 4992 4359
rect 5028 4221 5052 4959
rect 5208 4881 5232 5079
rect 5268 4941 5292 5136
rect 5328 5001 5352 5559
rect 5448 5481 5472 5772
rect 5499 5220 5541 5259
rect 5508 5208 5532 5220
rect 5628 5208 5652 6639
rect 5901 6672 5940 6681
rect 5901 6639 5952 6672
rect 5679 6561 5721 6579
rect 5928 6501 5952 6639
rect 5688 5841 5712 6339
rect 5928 6261 5952 6396
rect 5988 6321 6012 6639
rect 6048 6321 6072 6816
rect 6108 6501 6132 7599
rect 6288 7521 6312 8256
rect 6468 8220 6492 8232
rect 6348 7752 6372 8199
rect 6459 8181 6501 8220
rect 6648 8181 6672 8448
rect 6348 7728 6399 7752
rect 6408 7641 6432 7719
rect 6201 7512 6240 7521
rect 6201 7479 6252 7512
rect 6228 7428 6252 7479
rect 6399 7440 6441 7479
rect 6468 7461 6492 7959
rect 6408 7428 6432 7440
rect 6168 6801 6192 7179
rect 6288 7101 6312 7296
rect 6348 6981 6372 7059
rect 6528 6861 6552 8139
rect 6588 6921 6612 7479
rect 6648 7461 6672 7839
rect 6708 7752 6732 8619
rect 6768 8361 6792 8499
rect 6828 8421 6852 8859
rect 6948 8541 6972 8892
rect 7068 8880 7092 8892
rect 7059 8841 7101 8880
rect 7008 8601 7032 8799
rect 7128 8772 7152 8859
rect 7188 8841 7212 9159
rect 7068 8748 7152 8772
rect 6888 8328 6912 8439
rect 7068 8361 7092 8748
rect 7248 8721 7272 9279
rect 7308 8781 7332 9639
rect 7368 9441 7392 9792
rect 7428 9321 7452 9759
rect 7488 9741 7512 9999
rect 7548 9561 7572 10179
rect 7659 10101 7701 10119
rect 7428 8988 7452 9099
rect 7608 9012 7632 10059
rect 7788 10041 7812 10419
rect 7848 10392 7872 10452
rect 7968 10428 8052 10452
rect 7848 10368 7932 10392
rect 7908 10281 7932 10368
rect 7668 9921 7692 9996
rect 7908 9921 7932 10239
rect 7848 9780 7872 9792
rect 7839 9741 7881 9780
rect 7701 9699 7719 9735
rect 7728 9021 7752 9339
rect 7608 8988 7692 9012
rect 7188 8352 7212 8559
rect 7368 8421 7392 8799
rect 7188 8328 7239 8352
rect 6768 8121 6792 8199
rect 6828 7941 6852 8232
rect 6948 8172 6972 8232
rect 6888 8148 6972 8172
rect 6708 7728 6792 7752
rect 6708 7428 6732 7659
rect 6768 7461 6792 7728
rect 6888 7641 6912 8148
rect 6828 7308 6912 7332
rect 5799 5904 5841 5919
rect 5940 5892 5979 5901
rect 5928 5868 5979 5892
rect 5940 5859 5979 5868
rect 5808 5118 5832 5439
rect 5448 5100 5472 5112
rect 5439 5061 5481 5100
rect 5160 4392 5199 4401
rect 5148 4359 5199 4392
rect 5148 4344 5181 4359
rect 5328 3921 5352 4719
rect 5388 4581 5412 4719
rect 5568 4701 5592 5112
rect 5388 4341 5412 4539
rect 5568 4401 5592 4539
rect 5628 4461 5652 5019
rect 5688 4401 5712 5112
rect 5748 4641 5772 4899
rect 5868 4821 5892 5259
rect 5928 5241 5952 5619
rect 5988 5481 6012 5739
rect 6048 5304 6072 6279
rect 6108 6141 6132 6219
rect 6168 5952 6192 6639
rect 6348 6552 6372 6672
rect 6348 6528 6432 6552
rect 6228 6081 6252 6459
rect 6288 6141 6312 6219
rect 6348 5961 6372 6219
rect 6108 5928 6192 5952
rect 6108 5661 6132 5928
rect 6219 5892 6261 5919
rect 6408 5904 6432 6528
rect 6468 6261 6492 6759
rect 6648 6768 6672 7239
rect 6768 6861 6792 7299
rect 6888 6861 6912 7308
rect 6948 7161 6972 7779
rect 7008 7461 7032 8199
rect 7128 7941 7152 8232
rect 7248 7821 7272 8139
rect 7368 8112 7392 8199
rect 7428 8181 7452 8739
rect 7368 8088 7452 8112
rect 7059 7440 7101 7479
rect 7248 7461 7272 7716
rect 7308 7701 7332 8079
rect 7068 7428 7092 7440
rect 7308 7338 7332 7419
rect 7008 7221 7032 7299
rect 6768 6768 6912 6792
rect 7068 6768 7092 6999
rect 7119 6801 7161 6819
rect 6528 6552 6552 6756
rect 6579 6621 6621 6639
rect 6618 6600 6621 6621
rect 6528 6528 6612 6552
rect 6459 6081 6501 6099
rect 6168 5880 6261 5892
rect 6168 5868 6252 5880
rect 6168 5721 6192 5868
rect 6468 5868 6492 5976
rect 6288 5244 6312 5559
rect 6348 5541 6372 5772
rect 6588 5541 6612 6528
rect 6648 6381 6672 6579
rect 6708 6501 6732 6672
rect 6639 6081 6681 6099
rect 6708 6021 6732 6159
rect 6828 5961 6852 6519
rect 6888 6501 6912 6768
rect 7008 6621 7032 6672
rect 7008 6588 7059 6621
rect 7020 6579 7059 6588
rect 7101 6588 7152 6612
rect 7008 6081 7032 6519
rect 6888 5892 6912 5979
rect 6828 5868 6912 5892
rect 6348 5241 6372 5319
rect 6108 5061 6132 5112
rect 6219 5061 6261 5079
rect 6108 5028 6159 5061
rect 6120 5019 6159 5028
rect 6288 4821 6312 5202
rect 6528 5208 6552 5319
rect 6648 5241 6672 5559
rect 6348 4572 6372 5079
rect 6408 4812 6432 5019
rect 6468 4881 6492 5076
rect 6408 4788 6492 4812
rect 6468 4641 6492 4788
rect 6348 4548 6396 4572
rect 5481 4392 5520 4401
rect 5481 4359 5532 4392
rect 5508 4308 5532 4359
rect 5619 4320 5661 4356
rect 5628 4308 5652 4320
rect 5568 4200 5592 4212
rect 5559 4161 5601 4200
rect 5748 4161 5772 4302
rect 5808 4221 5832 4539
rect 5928 4341 5952 4419
rect 6168 4308 6192 4479
rect 6408 4308 6432 4539
rect 6468 4401 6492 4536
rect 6588 4341 6612 5076
rect 6708 4941 6732 5679
rect 6768 5241 6792 5772
rect 6948 5361 6972 5799
rect 7008 5601 7032 5919
rect 6768 4521 6792 5079
rect 6828 5001 6852 5112
rect 6888 4701 6912 4899
rect 6648 4221 6672 4479
rect 5448 3981 5472 4059
rect 5928 3981 5952 4179
rect 5988 4152 6012 4212
rect 5988 4128 6072 4152
rect 5079 3660 5121 3699
rect 5568 3684 5592 3759
rect 5928 3732 5952 3939
rect 5868 3708 5952 3732
rect 5088 3648 5112 3660
rect 5868 3648 5892 3708
rect 5988 3648 6012 4059
rect 6048 3681 6072 4128
rect 6159 3660 6201 3699
rect 6168 3648 6192 3660
rect 6288 3648 6312 4176
rect 6348 4101 6372 4212
rect 6468 4101 6492 4212
rect 6348 3981 6372 4059
rect 6348 3888 6459 3912
rect 6348 3741 6372 3888
rect 5388 3558 5412 3639
rect 4728 2658 4752 2736
rect 5088 2658 5112 3039
rect 5148 3021 5172 3552
rect 5148 2784 5172 2979
rect 5268 2901 5292 3552
rect 5388 2748 5412 3516
rect 5508 2658 5532 3516
rect 4428 2121 4452 2652
rect 4548 2088 4572 2379
rect 4968 2124 4992 2319
rect 5100 2112 5139 2121
rect 5088 2088 5139 2112
rect 5100 2079 5139 2088
rect 3648 1980 3672 1992
rect 3639 1941 3681 1980
rect 3981 1992 4020 2001
rect 3981 1968 4032 1992
rect 3981 1959 4020 1968
rect 2568 1248 2652 1272
rect 2568 1188 2592 1248
rect 2688 1188 2712 1359
rect 2148 1080 2172 1092
rect 2028 981 2052 1059
rect 2139 1041 2181 1080
rect 1788 438 1812 639
rect 1968 528 1992 819
rect 2208 612 2232 759
rect 2268 681 2292 1092
rect 2808 1092 2832 1359
rect 2868 1101 2892 1479
rect 2988 1188 3012 1539
rect 3108 1188 3132 1479
rect 2628 1080 2652 1092
rect 2619 1041 2661 1080
rect 2748 1068 2832 1092
rect 2448 621 2472 939
rect 2748 861 2772 1068
rect 2799 981 2841 999
rect 2208 588 2292 612
rect 2088 528 2232 552
rect 2028 420 2052 432
rect 2019 381 2061 420
rect 2208 261 2232 528
rect 2268 141 2292 588
rect 2508 528 2532 759
rect 2628 561 2652 639
rect 2688 321 2712 759
rect 2748 501 2772 819
rect 2808 441 2832 939
rect 3168 801 3192 1092
rect 2988 564 3012 759
rect 3288 741 3312 1539
rect 3528 1401 3552 1479
rect 3381 1212 3420 1221
rect 3381 1188 3432 1212
rect 3528 1188 3552 1359
rect 3648 1221 3672 1599
rect 3381 1179 3420 1188
rect 3828 1188 3852 1359
rect 3348 981 3372 1059
rect 3288 612 3312 699
rect 3228 588 3312 612
rect 3228 528 3252 588
rect 3288 420 3312 432
rect 2928 381 2961 396
rect 3279 381 3321 420
rect 3468 381 3492 519
rect 3528 381 3552 699
rect 3708 528 3732 819
rect 3828 528 3852 939
rect 3888 741 3912 1092
rect 4128 981 4152 1479
rect 4248 1401 4272 1959
rect 4428 1881 4452 2079
rect 5208 2001 5232 2439
rect 5328 2361 5352 2652
rect 5448 2241 5472 2319
rect 5568 2181 5592 3279
rect 5748 3261 5772 3639
rect 5748 3141 5772 3219
rect 5688 2748 5712 2919
rect 5799 2760 5841 2799
rect 5928 2781 5952 3552
rect 6468 3558 6492 3759
rect 6588 3732 6612 4179
rect 6648 3741 6672 4116
rect 6948 4101 6972 4779
rect 7068 4692 7092 6459
rect 7128 6321 7152 6588
rect 7188 6021 7212 6819
rect 7248 6501 7272 6879
rect 7308 6741 7332 6879
rect 7368 6861 7392 8019
rect 7428 7461 7452 8088
rect 7488 8061 7512 8679
rect 7548 8361 7572 8439
rect 7608 8421 7632 8619
rect 7668 8481 7692 8988
rect 7788 8988 7812 9459
rect 7908 9381 7932 9759
rect 7908 8988 7932 9159
rect 7968 9081 7992 10428
rect 8028 9912 8052 9999
rect 8088 9981 8112 11319
rect 8208 10941 8232 11352
rect 8808 11358 8832 11679
rect 8868 11481 8892 11979
rect 9108 11988 9192 12012
rect 9108 11601 9132 11988
rect 9348 11721 9372 12588
rect 9468 12132 9492 13659
rect 9528 13521 9552 14328
rect 9708 13701 9732 14559
rect 9768 13941 9792 15039
rect 9888 14841 9912 14919
rect 9948 14604 9972 14679
rect 9828 14001 9852 14079
rect 9768 13668 9792 13899
rect 9648 13281 9672 13572
rect 9888 13281 9912 14259
rect 9948 13701 9972 14379
rect 10068 14301 10092 15096
rect 10128 14601 10152 15936
rect 10188 15621 10212 15999
rect 10308 15501 10332 15939
rect 10368 15801 10392 16032
rect 10488 15741 10512 15996
rect 10848 15921 10872 15996
rect 10308 15228 10332 15459
rect 10548 15261 10572 15579
rect 10908 15561 10932 15999
rect 10188 14901 10212 15219
rect 10608 15141 10632 15519
rect 10668 15321 10692 15399
rect 10788 15264 10812 15399
rect 10908 15228 10932 15519
rect 10968 15261 10992 16539
rect 10368 14781 10392 15132
rect 10428 14841 10452 14919
rect 10188 14568 10212 14739
rect 10308 14568 10332 14679
rect 10488 14472 10512 14979
rect 10668 14961 10692 15216
rect 10788 14601 10812 14919
rect 10248 14361 10272 14472
rect 10368 14361 10392 14472
rect 10488 14448 10572 14472
rect 9948 13572 9972 13659
rect 10008 13641 10032 14139
rect 10488 13641 10512 13779
rect 10548 13701 10572 14448
rect 10728 14241 10752 14472
rect 10668 13941 10692 14019
rect 10728 13941 10752 14199
rect 10788 13668 10812 14439
rect 10848 14361 10872 14559
rect 10848 13701 10872 14079
rect 9948 13548 10032 13572
rect 9588 12741 9612 12912
rect 9768 12888 9852 12912
rect 9828 12801 9852 12888
rect 9768 12381 9792 12579
rect 9408 12108 9492 12132
rect 9408 11601 9432 12108
rect 9828 12072 9852 12759
rect 9888 12261 9912 13119
rect 9948 12321 9972 13419
rect 10008 13161 10032 13548
rect 10248 13221 10272 13452
rect 10008 12108 10032 12219
rect 10068 12201 10092 12912
rect 10188 12132 10212 12912
rect 10368 12741 10392 13119
rect 10488 13044 10512 13479
rect 10668 13461 10692 13572
rect 10608 13008 10632 13119
rect 10728 13041 10752 13299
rect 10548 12381 10572 12912
rect 10728 12621 10752 12819
rect 10788 12441 10812 13179
rect 10848 12801 10872 13419
rect 10908 13101 10932 15039
rect 10968 14961 10992 15099
rect 11028 15081 11052 16479
rect 11208 16401 11232 17508
rect 11388 17301 11412 17379
rect 11568 17361 11592 18699
rect 11328 16461 11352 16692
rect 11508 16161 11532 16779
rect 11568 16701 11592 17139
rect 11628 16821 11652 18759
rect 11688 18384 11712 18459
rect 11739 18384 11781 18399
rect 12048 18381 12072 18459
rect 11688 18261 11712 18342
rect 11739 18192 11781 18219
rect 11928 18240 11952 18252
rect 11919 18201 11961 18240
rect 11739 18180 11832 18192
rect 11748 18168 11832 18180
rect 11808 17688 11832 18168
rect 11928 17688 11952 17799
rect 11868 17541 11892 17592
rect 12048 17541 12072 18159
rect 12108 17841 12132 18342
rect 12201 18252 12240 18261
rect 12201 18228 12252 18252
rect 12201 18219 12240 18228
rect 12408 18201 12432 18339
rect 12468 18081 12492 18342
rect 12648 18141 12672 18252
rect 12888 18252 12912 18459
rect 13068 18384 13092 18639
rect 13128 18621 13152 18699
rect 13188 18348 13212 18459
rect 12828 18228 12912 18252
rect 12708 18021 12732 18159
rect 12768 18072 12792 18216
rect 12828 18141 12852 18228
rect 12768 18048 12852 18072
rect 12588 17901 12612 17979
rect 12408 17724 12432 17799
rect 12828 17781 12852 18048
rect 12888 17781 12912 18159
rect 13008 18081 13032 18252
rect 12759 17700 12801 17739
rect 12768 17688 12792 17700
rect 11688 16788 11712 17199
rect 11808 17061 11832 17259
rect 11868 17121 11892 17499
rect 12228 17481 12252 17556
rect 12348 17421 12372 17592
rect 12558 17559 12561 17580
rect 12519 17541 12561 17559
rect 12708 17580 12732 17592
rect 12699 17541 12741 17580
rect 13008 17598 13032 17976
rect 13068 17781 13092 17979
rect 13128 17781 13152 18252
rect 13188 17688 13212 18099
rect 13308 18021 13332 18699
rect 14388 18348 14412 18459
rect 13668 18258 13692 18339
rect 13368 17901 13392 18216
rect 13548 18141 13572 18216
rect 13299 17700 13341 17739
rect 13308 17688 13332 17700
rect 13428 17598 13452 17919
rect 13488 17841 13512 18099
rect 13608 17688 13632 17799
rect 13668 17772 13692 18216
rect 13728 18141 13752 18279
rect 13668 17748 13752 17772
rect 13728 17688 13752 17748
rect 13848 17721 13872 17799
rect 13908 17598 13932 17919
rect 12828 17421 12852 17559
rect 13248 17481 13272 17592
rect 13188 17448 13239 17472
rect 11568 16128 11592 16539
rect 11628 16521 11652 16659
rect 11748 16461 11772 16692
rect 11868 16512 11892 16659
rect 11988 16581 12012 17079
rect 12048 16821 12072 16959
rect 12108 16941 12132 17259
rect 12168 16788 12192 17319
rect 12708 16788 12732 17139
rect 13128 16941 13152 17379
rect 13128 16821 13152 16899
rect 11868 16488 11952 16512
rect 11688 16128 11712 16359
rect 11928 16341 11952 16488
rect 11808 16161 11832 16299
rect 12048 16212 12072 16659
rect 12108 16581 12132 16692
rect 12228 16581 12252 16692
rect 12408 16452 12432 16782
rect 12528 16680 12552 16692
rect 12519 16641 12561 16680
rect 12648 16461 12672 16692
rect 12408 16428 12459 16452
rect 12048 16188 12132 16212
rect 11841 16128 11892 16152
rect 12108 16128 12132 16188
rect 11208 15801 11232 16032
rect 11148 15501 11172 15699
rect 11328 15681 11352 16032
rect 11448 15921 11472 16119
rect 11628 15972 11652 16032
rect 11568 15948 11652 15972
rect 11481 15468 11532 15492
rect 11088 14661 11112 15339
rect 11328 15228 11352 15339
rect 11448 15228 11472 15459
rect 11508 15381 11532 15468
rect 11148 15021 11172 15099
rect 11268 15072 11292 15132
rect 11268 15048 11352 15072
rect 11268 14601 11292 14919
rect 11328 14841 11352 15048
rect 11388 15021 11412 15132
rect 11568 15081 11592 15948
rect 11748 15801 11772 15996
rect 11808 15741 11832 15996
rect 11628 15261 11652 15699
rect 11868 15612 11892 16128
rect 12228 15921 12252 16299
rect 11928 15741 11952 15819
rect 11808 15588 11892 15612
rect 11688 15228 11712 15399
rect 11808 15261 11832 15588
rect 11868 15381 11892 15519
rect 11928 15252 11952 15699
rect 11868 15228 11952 15252
rect 11748 15120 11772 15132
rect 11739 15081 11781 15120
rect 11448 14841 11472 14919
rect 11388 14568 11412 14739
rect 10968 14361 10992 14559
rect 11088 14121 11112 14472
rect 10968 13032 10992 14019
rect 11088 13668 11112 14016
rect 11328 13581 11352 14139
rect 11148 13341 11172 13572
rect 11148 13092 11172 13179
rect 11148 13068 11232 13092
rect 11208 13050 11232 13068
rect 10908 13008 10992 13032
rect 10908 12561 10932 13008
rect 10968 12621 10992 12879
rect 11028 12801 11052 12912
rect 10161 12108 10212 12132
rect 9828 12048 9879 12072
rect 8979 11460 9021 11499
rect 8988 11448 9012 11460
rect 8388 11121 8412 11256
rect 8148 10101 8172 10839
rect 8388 10641 8412 11079
rect 8568 10761 8592 11259
rect 8628 10881 8652 11352
rect 9168 11301 9192 11499
rect 8688 11061 8712 11259
rect 8259 10560 8301 10599
rect 8268 10548 8292 10560
rect 8388 10548 8412 10599
rect 8559 10581 8601 10599
rect 8619 10560 8661 10599
rect 8628 10548 8652 10560
rect 8748 10548 8772 10959
rect 8988 10584 9012 11079
rect 8328 10281 8352 10452
rect 8208 9921 8232 10119
rect 8028 9888 8112 9912
rect 8028 9381 8052 9759
rect 8148 9681 8172 9792
rect 8028 9012 8052 9339
rect 8088 9141 8112 9579
rect 8028 8988 8112 9012
rect 8088 8901 8112 8988
rect 7848 8880 7872 8892
rect 7839 8841 7881 8880
rect 7599 8340 7641 8379
rect 7608 8328 7632 8340
rect 7788 8301 7812 8799
rect 7968 8601 7992 8892
rect 8148 8781 8172 9039
rect 8208 9021 8232 9759
rect 8268 9321 8292 9939
rect 8328 9741 8352 10059
rect 8448 9981 8472 10299
rect 8508 10101 8532 10479
rect 8808 10221 8832 10452
rect 8619 9921 8661 9939
rect 8688 9741 8712 10119
rect 8928 10041 8952 10359
rect 8988 10341 9012 10542
rect 9048 10161 9072 10719
rect 9108 10101 9132 11019
rect 9168 10572 9192 10899
rect 9228 10701 9252 11559
rect 9468 11448 9492 11979
rect 9888 11901 9912 12039
rect 10488 12012 10512 12279
rect 10188 11781 10212 11979
rect 9588 11601 9612 11679
rect 9588 11448 9612 11559
rect 9648 11481 9672 11619
rect 9681 11472 9720 11481
rect 9681 11448 9732 11472
rect 9681 11439 9720 11448
rect 9288 11301 9312 11439
rect 9408 11340 9432 11352
rect 9399 11301 9441 11340
rect 9528 11241 9552 11316
rect 9528 10821 9552 10899
rect 9588 10821 9612 11079
rect 9648 10701 9672 11259
rect 9888 11232 9912 11739
rect 10248 11721 10272 11859
rect 10488 11841 10512 11970
rect 10548 11781 10572 12099
rect 10908 11901 10932 11979
rect 9948 11361 9972 11499
rect 10308 11481 10332 11739
rect 10368 11352 10392 11679
rect 9888 11208 9939 11232
rect 10128 11232 10152 11319
rect 10428 11301 10452 11619
rect 10521 11508 10692 11532
rect 10668 11448 10692 11508
rect 10068 11208 10152 11232
rect 9948 11001 9972 11199
rect 10068 11061 10092 11208
rect 9168 10548 9252 10572
rect 9468 10581 9492 10659
rect 9708 10548 9732 10779
rect 9768 10581 9792 10899
rect 8328 9501 8352 9699
rect 8268 9081 8292 9279
rect 8448 9084 8472 9459
rect 8508 9261 8532 9339
rect 8268 8832 8292 8892
rect 8268 8808 8352 8832
rect 8208 8421 8232 8499
rect 8199 8340 8241 8379
rect 8208 8328 8232 8340
rect 7548 7641 7572 8139
rect 7599 8121 7641 8139
rect 7668 8061 7692 8232
rect 7728 8001 7752 8199
rect 7848 8181 7872 8319
rect 7908 8112 7932 8259
rect 8328 8238 8352 8808
rect 8388 8781 8412 8892
rect 8388 8361 8412 8676
rect 8508 8364 8532 8859
rect 8568 8721 8592 9579
rect 8628 9381 8652 9639
rect 8688 9141 8712 9519
rect 8748 9201 8772 9999
rect 8808 9681 8832 9759
rect 8679 9000 8721 9036
rect 8688 8988 8712 9000
rect 8808 8988 8832 9459
rect 8988 9261 9012 9792
rect 8919 9000 8961 9039
rect 8988 9021 9012 9219
rect 8928 8988 8952 9000
rect 8628 8601 8652 8859
rect 8868 8661 8892 8892
rect 9048 8781 9072 9639
rect 9108 9621 9132 9939
rect 9228 9888 9252 9999
rect 9288 9981 9312 10452
rect 9408 10281 9432 10452
rect 9468 10341 9492 10419
rect 9348 9888 9372 10179
rect 9408 10041 9432 10239
rect 9288 9681 9312 9792
rect 9141 9408 9219 9432
rect 9108 8901 9132 9159
rect 9168 9021 9192 9339
rect 9408 9321 9432 9519
rect 9528 9321 9552 10419
rect 9588 10221 9612 10359
rect 9648 10341 9672 10452
rect 9768 10281 9792 10419
rect 9828 10401 9852 10959
rect 10488 10881 10512 11319
rect 10608 10881 10632 11352
rect 10728 11241 10752 11352
rect 10848 10881 10872 11679
rect 10968 11541 10992 12399
rect 11028 11721 11052 12339
rect 11088 12141 11112 12759
rect 11148 12501 11172 12879
rect 11148 12108 11172 12459
rect 11328 12432 11352 12579
rect 11388 12501 11412 14379
rect 11568 14361 11592 14472
rect 11448 13704 11472 13839
rect 11628 13821 11652 14439
rect 11688 13752 11712 15039
rect 11748 14061 11772 14679
rect 11808 14181 11832 14739
rect 11928 14661 11952 15099
rect 11988 14781 12012 15879
rect 12108 15561 12132 15639
rect 12048 15381 12072 15459
rect 12108 15228 12132 15519
rect 12198 15339 12201 15360
rect 12159 15321 12201 15339
rect 12228 15228 12252 15339
rect 12288 15321 12312 16239
rect 12468 16128 12492 16419
rect 12768 16041 12792 16599
rect 12828 16041 12852 16782
rect 13020 16152 13059 16161
rect 13008 16128 13059 16152
rect 13020 16119 13059 16128
rect 13128 16041 13152 16539
rect 13188 16341 13212 17448
rect 13668 17061 13692 17592
rect 13248 16281 13272 17019
rect 13548 16788 13572 16899
rect 13788 16788 13812 17079
rect 13968 16812 13992 18132
rect 14028 17721 14052 18099
rect 14208 17961 14232 18219
rect 14568 18021 14592 18252
rect 14688 18021 14712 18342
rect 14808 18141 14832 18639
rect 14868 18621 14892 18912
rect 15348 18741 15372 18912
rect 14928 18348 14952 18459
rect 15039 18360 15081 18399
rect 15048 18348 15072 18360
rect 14241 17928 14292 17952
rect 14148 17688 14172 17859
rect 14268 17721 14292 17928
rect 14328 17598 14352 17859
rect 14388 17721 14412 17979
rect 14988 17961 15012 18252
rect 14508 17688 14532 17799
rect 14448 17241 14472 17439
rect 13968 16788 14052 16812
rect 13308 16581 13332 16782
rect 13368 16521 13392 16659
rect 13608 16521 13632 16692
rect 13848 16680 13872 16692
rect 13839 16641 13881 16680
rect 13608 16341 13632 16479
rect 13788 16164 13812 16539
rect 13908 16461 13932 16539
rect 13968 16392 13992 16659
rect 14028 16461 14052 16788
rect 14088 16521 14112 16899
rect 14208 16788 14232 17139
rect 14448 16821 14472 17019
rect 13968 16368 14052 16392
rect 12348 15441 12372 15999
rect 12648 15921 12672 16032
rect 12861 16020 12912 16032
rect 12861 16008 12921 16020
rect 12648 15732 12672 15879
rect 12708 15801 12732 15999
rect 12879 15981 12921 16008
rect 13488 16038 13512 16119
rect 13068 15921 13092 15999
rect 12648 15708 12732 15732
rect 12468 15561 12492 15639
rect 12408 15321 12432 15459
rect 12048 14961 12072 15099
rect 12168 14781 12192 15132
rect 12099 14580 12141 14619
rect 12228 14604 12252 15039
rect 12288 14961 12312 15132
rect 12348 14781 12372 14979
rect 12408 14841 12432 15099
rect 12468 14661 12492 15399
rect 12528 14721 12552 15579
rect 12621 15552 12660 15561
rect 12621 15519 12672 15552
rect 12588 15261 12612 15456
rect 12648 15228 12672 15519
rect 12708 15321 12732 15708
rect 13008 15621 13032 15699
rect 12768 15228 12792 15519
rect 12888 15228 12912 15579
rect 13068 15252 13092 15879
rect 13248 15861 13272 16032
rect 13368 15921 13392 16032
rect 13008 15228 13092 15252
rect 13128 15228 13152 15639
rect 13248 15441 13272 15819
rect 13239 15240 13281 15279
rect 13248 15228 13272 15240
rect 12588 14901 12612 15099
rect 12588 14661 12612 14739
rect 12108 14568 12132 14580
rect 12540 14598 12600 14601
rect 12540 14589 12579 14598
rect 12528 14565 12579 14589
rect 12228 14481 12252 14562
rect 12540 14559 12579 14565
rect 12648 14541 12672 14979
rect 12828 14961 12852 15132
rect 12948 14901 12972 15099
rect 12348 14460 12372 14472
rect 11868 14112 11892 14259
rect 11808 14088 11892 14112
rect 11628 13728 11712 13752
rect 11628 13668 11652 13728
rect 11328 12408 11412 12432
rect 11268 12108 11292 12219
rect 11388 12012 11412 12408
rect 11448 12381 11472 13662
rect 11508 13041 11532 13539
rect 11568 13461 11592 13572
rect 11688 13461 11712 13572
rect 11808 13401 11832 14088
rect 11988 14001 12012 14079
rect 12048 13704 12072 14436
rect 11868 13548 11952 13572
rect 11868 13221 11892 13548
rect 11580 12912 11619 12921
rect 11568 12888 11619 12912
rect 11580 12879 11619 12888
rect 11508 12312 11532 12879
rect 11748 12801 11772 12912
rect 11328 11988 11412 12012
rect 11448 12288 11532 12312
rect 10968 11340 10992 11352
rect 10959 11301 11001 11340
rect 10008 10584 10032 10839
rect 10128 10584 10152 10839
rect 10968 10821 10992 11259
rect 11088 11121 11112 11352
rect 9948 10440 9972 10452
rect 9888 10161 9912 10419
rect 9939 10401 9981 10440
rect 9588 9141 9612 9939
rect 9648 9798 9672 9999
rect 9768 9888 9792 10119
rect 9708 9201 9732 9699
rect 9768 9381 9792 9519
rect 9528 9021 9552 9099
rect 9141 8868 9192 8892
rect 8688 8241 8712 8439
rect 8928 8328 8952 8439
rect 9108 8361 9132 8796
rect 7848 8088 7932 8112
rect 8259 8172 8301 8199
rect 7959 8112 8001 8139
rect 8208 8160 8301 8172
rect 8208 8148 8292 8160
rect 7959 8100 8052 8112
rect 7968 8088 8052 8100
rect 7548 7428 7572 7536
rect 7668 7428 7692 7839
rect 7428 6981 7452 7299
rect 7488 7161 7512 7332
rect 7788 7101 7812 7899
rect 7848 7464 7872 8088
rect 7908 7521 7932 8019
rect 8028 7932 8052 8088
rect 8208 8052 8232 8148
rect 8148 8028 8232 8052
rect 8148 8001 8172 8028
rect 8121 7968 8172 8001
rect 8121 7959 8160 7968
rect 8028 7908 8139 7932
rect 8088 7761 8112 7839
rect 8268 7812 8292 8079
rect 8208 7788 8292 7812
rect 8028 7521 8052 7659
rect 8028 7482 8079 7521
rect 7908 7428 7932 7479
rect 8148 7461 8172 7539
rect 8100 7332 8139 7341
rect 7968 7101 7992 7332
rect 8088 7299 8139 7332
rect 7488 6768 7512 7056
rect 7308 6441 7332 6636
rect 7428 6381 7452 6672
rect 7248 5868 7272 6339
rect 7548 6201 7572 6339
rect 7608 6261 7632 6672
rect 7668 6321 7692 6579
rect 7641 6228 7692 6252
rect 7359 6141 7401 6159
rect 7341 6120 7401 6141
rect 7341 6108 7392 6120
rect 7341 6099 7380 6108
rect 7299 5961 7341 5979
rect 7368 5868 7392 6039
rect 7581 5979 7599 6021
rect 7428 5901 7452 5979
rect 7668 5952 7692 6228
rect 7788 5961 7812 6939
rect 8028 6768 8052 6999
rect 8088 6801 8112 7299
rect 8139 7221 8181 7236
rect 8148 6741 8172 6879
rect 8148 6552 8172 6636
rect 8208 6621 8232 7788
rect 8268 7335 8292 7479
rect 8328 7461 8352 8196
rect 8448 8121 8472 8232
rect 8388 7761 8412 7959
rect 8568 7821 8592 8196
rect 8748 8172 8772 8319
rect 8688 8148 8772 8172
rect 8688 8001 8712 8148
rect 8868 8121 8892 8232
rect 8508 7428 8532 7539
rect 8568 7521 8592 7659
rect 8748 7461 8772 8079
rect 8868 8001 8892 8079
rect 8808 7401 8832 7719
rect 8928 7512 8952 8019
rect 9108 7521 9132 8199
rect 9168 7761 9192 8868
rect 9348 8781 9372 8892
rect 9468 8841 9492 8982
rect 9828 9021 9852 9579
rect 9888 8901 9912 9699
rect 9948 9501 9972 9792
rect 10068 9081 10092 10452
rect 10308 10452 10332 10542
rect 10728 10458 10752 10659
rect 11208 10641 11232 11499
rect 11328 11481 11352 11988
rect 11448 11481 11472 12288
rect 11748 12108 11772 12219
rect 11868 12141 11892 13059
rect 11928 12801 11952 13239
rect 11988 12918 12012 13479
rect 12048 13341 12072 13419
rect 12168 13281 12192 14139
rect 12228 13101 12252 14319
rect 12288 14001 12312 14439
rect 12339 14421 12381 14460
rect 12468 13668 12492 13839
rect 12528 13701 12552 14379
rect 12588 14181 12612 14439
rect 12648 14121 12672 14499
rect 12708 14241 12732 14859
rect 12888 14568 12912 14799
rect 13008 14601 13032 15228
rect 12828 14241 12852 14472
rect 13008 14361 13032 14439
rect 12588 13578 12612 13959
rect 12828 13881 12852 14199
rect 13068 14121 13092 15099
rect 13128 14301 13152 14919
rect 13188 14721 13212 15132
rect 13308 14604 13332 15039
rect 13368 14961 13392 15639
rect 13428 14661 13452 15759
rect 13488 15261 13512 15699
rect 13548 15264 13572 15579
rect 13668 15381 13692 15519
rect 13728 15501 13752 16032
rect 13488 14601 13512 15099
rect 13440 14472 13479 14481
rect 13428 14448 13479 14472
rect 13440 14439 13479 14448
rect 13368 14361 13392 14439
rect 13548 14301 13572 14619
rect 13608 14601 13632 15099
rect 13668 14901 13692 15132
rect 13668 14721 13692 14859
rect 13848 14841 13872 16239
rect 14028 16128 14052 16368
rect 14268 16332 14292 16692
rect 14388 16521 14412 16692
rect 14328 16401 14352 16479
rect 14448 16332 14472 16659
rect 14508 16581 14532 16899
rect 14568 16521 14592 17079
rect 14748 16884 14772 17799
rect 14808 17061 14832 17679
rect 14868 17592 14892 17739
rect 14868 17568 15012 17592
rect 14628 16401 14652 16839
rect 14868 16788 14892 17199
rect 14268 16308 14472 16332
rect 14148 16152 14172 16299
rect 14568 16281 14592 16359
rect 14148 16128 14232 16152
rect 14088 16020 14112 16032
rect 14079 15981 14121 16020
rect 13908 15081 13932 15459
rect 13968 15261 13992 15639
rect 14148 15312 14172 15939
rect 14208 15681 14232 16128
rect 14268 15981 14292 16239
rect 14508 16128 14532 16239
rect 14361 15939 14379 15981
rect 14148 15288 14232 15312
rect 14208 15261 14232 15288
rect 14208 15228 14259 15261
rect 14220 15219 14259 15228
rect 13968 14772 13992 15099
rect 14028 14961 14052 15132
rect 14328 15081 14352 15519
rect 14448 15321 14472 16032
rect 14628 15921 14652 16122
rect 14688 15801 14712 16659
rect 14748 15621 14772 16419
rect 14928 16392 14952 16692
rect 15048 16521 15072 17559
rect 15228 17061 15252 18699
rect 15288 17541 15312 18159
rect 15348 18141 15372 18216
rect 15468 18081 15492 18252
rect 15519 18201 15561 18219
rect 15588 18201 15612 18759
rect 15648 18261 15672 18399
rect 15828 18348 15852 18459
rect 15768 18240 15792 18252
rect 15759 18201 15801 18240
rect 15648 18021 15672 18099
rect 15348 17721 15372 17859
rect 15648 17721 15672 17979
rect 15768 17688 15792 17799
rect 15888 17721 15912 18219
rect 15528 17568 15612 17592
rect 15159 16800 15201 16839
rect 15168 16788 15192 16800
rect 15288 16788 15312 17259
rect 15348 16941 15372 17319
rect 15468 17241 15492 17319
rect 15408 16788 15432 17079
rect 15468 16821 15492 16959
rect 14928 16368 15012 16392
rect 14988 16161 15012 16368
rect 15039 16212 15081 16239
rect 15108 16212 15132 16539
rect 15039 16200 15132 16212
rect 15048 16188 15132 16200
rect 15048 16128 15072 16188
rect 14928 16020 14952 16032
rect 14919 15981 14961 16020
rect 15108 16008 15192 16032
rect 14928 15681 14952 15759
rect 14988 15501 15012 15999
rect 14508 15228 14532 15339
rect 14199 15012 14241 15039
rect 14148 15000 14241 15012
rect 14148 14988 14232 15000
rect 14148 14952 14172 14988
rect 14088 14928 14172 14952
rect 13968 14748 14052 14772
rect 13908 14661 13932 14739
rect 13608 14301 13632 14439
rect 13008 13941 13032 14019
rect 12948 13668 13092 13692
rect 12408 13560 12432 13572
rect 12399 13521 12441 13560
rect 12438 13500 12441 13521
rect 12468 13008 12492 13479
rect 12888 13461 12912 13662
rect 12948 13461 12972 13668
rect 12048 12261 12072 12459
rect 12228 12381 12252 12912
rect 11508 12021 11532 12102
rect 11508 11448 11532 11799
rect 11568 11481 11592 11919
rect 11688 11781 11712 12012
rect 11808 11781 11832 12012
rect 11268 11241 11292 11439
rect 11388 11292 11412 11316
rect 11328 11268 11412 11292
rect 11088 10458 11112 10599
rect 11328 10581 11352 11268
rect 11568 11172 11592 11319
rect 11508 11148 11592 11172
rect 10308 10428 10392 10452
rect 10128 9921 10152 10359
rect 10188 10041 10212 10419
rect 10308 9981 10332 10239
rect 10368 9888 10392 10428
rect 10428 9921 10452 10179
rect 10488 9798 10512 9939
rect 10128 9621 10152 9759
rect 10188 9501 10212 9792
rect 10548 9681 10572 10452
rect 10728 10341 10752 10416
rect 11208 10341 11232 10452
rect 10659 9900 10701 9939
rect 10668 9888 10692 9900
rect 10848 9801 10872 9939
rect 11079 9900 11121 9939
rect 11199 9900 11241 9939
rect 11088 9888 11112 9900
rect 11208 9888 11232 9900
rect 11328 9798 11352 10419
rect 11388 10041 11412 10539
rect 11448 9912 11472 10539
rect 11508 10281 11532 11148
rect 11628 10641 11652 11559
rect 11928 11481 11952 12219
rect 12048 12108 12072 12219
rect 12159 12120 12201 12159
rect 12219 12141 12261 12159
rect 12168 12108 12192 12120
rect 12288 11961 12312 12759
rect 12408 12621 12432 12879
rect 11988 11421 12012 11919
rect 12228 11448 12252 11559
rect 12348 11541 12372 12219
rect 12408 12141 12432 12579
rect 12528 12381 12552 12912
rect 12588 12561 12612 12879
rect 12648 12201 12672 13419
rect 13128 13341 13152 13536
rect 12708 12501 12732 13239
rect 12888 13008 12912 13119
rect 12768 12741 12792 12912
rect 12948 12381 12972 12852
rect 12459 12120 12501 12159
rect 12468 12108 12492 12120
rect 12708 12141 12732 12339
rect 12900 12192 12939 12201
rect 12888 12159 12939 12192
rect 12888 12108 12912 12159
rect 12408 11472 12432 11979
rect 12528 11721 12552 12012
rect 12768 12012 12792 12102
rect 13068 12018 13092 12279
rect 12708 11988 12792 12012
rect 12648 11781 12672 11976
rect 12348 11448 12432 11472
rect 11688 11061 11712 11319
rect 11748 10992 11772 11352
rect 12048 11352 12072 11448
rect 12648 11361 12672 11676
rect 12048 11328 12132 11352
rect 11868 11292 11892 11316
rect 11688 10968 11772 10992
rect 11808 11268 11892 11292
rect 11688 10941 11712 10968
rect 11688 10572 11712 10899
rect 11808 10581 11832 11268
rect 11988 11112 12012 11316
rect 11988 11088 12039 11112
rect 11628 10548 11712 10572
rect 12048 10521 12072 11079
rect 11748 10221 11772 10452
rect 12108 10401 12132 11328
rect 12168 11061 12192 11352
rect 12288 11181 12312 11352
rect 12219 10560 12261 10599
rect 12468 10572 12492 10959
rect 12228 10548 12252 10560
rect 12408 10548 12492 10572
rect 11388 9888 11472 9912
rect 9228 7581 9252 8739
rect 9528 8721 9552 8859
rect 9519 8460 9561 8499
rect 9528 8448 9552 8460
rect 9708 8277 9732 8799
rect 9288 8001 9312 8259
rect 9699 8238 9741 8259
rect 9768 8052 9792 8259
rect 9828 8061 9852 8859
rect 9888 8361 9912 8679
rect 9948 8421 9972 9039
rect 10068 8601 10092 8892
rect 10188 8601 10212 8892
rect 10188 8361 10212 8559
rect 9708 8028 9792 8052
rect 9261 7548 9312 7572
rect 8868 7488 8952 7512
rect 8439 7281 8481 7299
rect 8568 7161 8592 7332
rect 8739 7281 8781 7299
rect 8508 6981 8532 7059
rect 8448 6768 8472 6879
rect 8808 6804 8832 7359
rect 8301 6672 8340 6681
rect 8301 6648 8352 6672
rect 8301 6639 8340 6648
rect 8148 6528 8232 6552
rect 7539 5904 7581 5916
rect 7488 5868 7539 5892
rect 7488 5778 7512 5868
rect 7608 5928 7692 5952
rect 7608 5868 7632 5928
rect 7188 5760 7212 5772
rect 7179 5721 7221 5760
rect 7668 5601 7692 5772
rect 7128 5118 7152 5499
rect 7188 5301 7212 5439
rect 7248 5361 7272 5439
rect 7248 5208 7272 5319
rect 7368 5208 7392 5559
rect 7308 5052 7332 5112
rect 7308 5028 7392 5052
rect 7041 4668 7092 4692
rect 6528 3720 6612 3732
rect 6519 3708 6612 3720
rect 6519 3681 6561 3708
rect 6558 3660 6561 3681
rect 6699 3660 6741 3699
rect 6828 3681 6852 4059
rect 6948 3921 6972 4059
rect 7008 3792 7032 4659
rect 7248 4308 7272 4599
rect 7308 4461 7332 4539
rect 6948 3768 7032 3792
rect 6708 3648 6732 3660
rect 6888 3558 6912 3639
rect 6228 3540 6252 3552
rect 6108 3261 6132 3519
rect 6219 3501 6261 3540
rect 5808 2748 5832 2760
rect 5988 2658 6012 2859
rect 6108 2784 6132 3219
rect 6228 2748 6252 2979
rect 6288 2832 6312 3099
rect 6381 2859 6399 2901
rect 6288 2808 6372 2832
rect 6348 2748 6372 2808
rect 5868 2361 5892 2439
rect 5838 2319 5841 2340
rect 5799 2292 5841 2319
rect 5799 2280 5892 2292
rect 5808 2268 5892 2280
rect 5499 2100 5541 2139
rect 5508 2088 5532 2100
rect 4608 1980 4632 1992
rect 4599 1941 4641 1980
rect 4488 1821 4512 1899
rect 4908 1881 4932 1992
rect 5019 1941 5061 1956
rect 5268 1941 5292 2079
rect 5319 1941 5361 1959
rect 4188 1041 4212 1239
rect 4428 801 4452 972
rect 3768 420 3792 432
rect 3759 381 3801 420
rect 2928 348 2979 381
rect 2940 339 2979 348
rect 3720 318 3780 321
rect 3639 252 3681 279
rect 3741 279 3759 318
rect 3828 252 3852 339
rect 3639 240 3852 252
rect 3648 228 3852 240
rect 4008 141 4032 522
rect 4428 438 4452 519
rect 4128 420 4152 432
rect 4119 381 4161 420
rect 4488 261 4512 879
rect 4548 438 4572 699
rect 4608 561 4632 819
rect 4728 528 4752 1299
rect 4848 1221 4872 1659
rect 4968 1224 4992 1719
rect 5448 1641 5472 1992
rect 4821 1188 4872 1221
rect 4821 1179 4860 1188
rect 4848 561 4872 699
rect 4908 681 4932 1092
rect 5088 1041 5112 1479
rect 5568 1461 5592 1956
rect 5688 1761 5712 2139
rect 5748 2121 5772 2259
rect 5868 2088 5892 2268
rect 5988 2088 6012 2199
rect 6048 2112 6072 2739
rect 6468 2658 6492 2919
rect 6519 2901 6561 2919
rect 6168 2640 6192 2652
rect 6159 2601 6201 2640
rect 6228 2121 6252 2379
rect 6048 2088 6132 2112
rect 5928 1821 5952 1992
rect 6048 1641 6072 1959
rect 6108 1701 6132 2088
rect 6468 2088 6492 2379
rect 6588 2361 6612 2979
rect 6888 2781 6912 3516
rect 6948 3501 6972 3768
rect 7188 3741 7212 4212
rect 7008 3321 7032 3699
rect 7248 3648 7272 4119
rect 7368 3732 7392 5028
rect 7428 4401 7452 5079
rect 7488 5001 7512 5379
rect 7848 5118 7872 6459
rect 7908 5421 7932 6519
rect 8028 5904 8052 6279
rect 8148 5868 8172 6039
rect 8208 5901 8232 6528
rect 8268 5841 8292 6219
rect 8328 5772 8352 6579
rect 8868 6441 8892 7488
rect 9141 7488 9192 7512
rect 9168 7428 9192 7488
rect 9288 7461 9312 7548
rect 8928 7221 8952 7419
rect 9108 7320 9132 7332
rect 8928 6501 8952 7059
rect 8988 6981 9012 7299
rect 9099 7281 9141 7320
rect 9108 6768 9132 6939
rect 9228 6804 9252 7233
rect 9348 7101 9372 7779
rect 9441 7332 9480 7341
rect 9441 7308 9492 7332
rect 9441 7299 9480 7308
rect 9408 6768 9432 7119
rect 9648 6801 9672 7719
rect 8988 6681 9012 6762
rect 9600 6672 9639 6681
rect 9168 6660 9192 6672
rect 9468 6660 9492 6672
rect 9159 6621 9201 6660
rect 9459 6621 9501 6660
rect 9588 6648 9639 6672
rect 9600 6639 9639 6648
rect 8421 5892 8460 5901
rect 8421 5868 8472 5892
rect 8559 5880 8601 5919
rect 8568 5868 8592 5880
rect 8421 5859 8460 5868
rect 9348 5868 9492 5892
rect 7908 5121 7932 5259
rect 7968 5241 7992 5739
rect 8088 5421 8112 5772
rect 8268 5748 8352 5772
rect 8148 5361 8172 5499
rect 8268 5481 8292 5748
rect 7488 4401 7512 4959
rect 7728 4941 7752 5112
rect 7848 4941 7872 5076
rect 8328 5061 8352 5679
rect 8388 5421 8412 5739
rect 8508 5601 8532 5772
rect 8628 5760 8652 5772
rect 8619 5721 8661 5760
rect 8748 5721 8772 5862
rect 8958 5673 8961 5700
rect 8919 5661 8961 5673
rect 8568 5208 8592 5319
rect 7719 4320 7761 4359
rect 7899 4320 7941 4359
rect 8028 4344 8052 4959
rect 7728 4308 7752 4320
rect 7908 4308 7932 4320
rect 7428 3801 7452 4296
rect 7548 3741 7572 4059
rect 7368 3708 7452 3732
rect 6828 2748 6879 2772
rect 7008 2748 7032 3216
rect 7068 3141 7092 3519
rect 7428 3552 7452 3708
rect 7539 3660 7581 3699
rect 7548 3648 7572 3660
rect 7848 3552 7872 4059
rect 7968 3921 7992 4212
rect 8208 4101 8232 5013
rect 8448 4941 8472 5076
rect 8628 4641 8652 5112
rect 8499 4320 8541 4359
rect 8508 4308 8532 4320
rect 8268 4161 8292 4302
rect 8220 4032 8259 4041
rect 8208 3999 8259 4032
rect 8028 3648 8052 3939
rect 8139 3660 8181 3699
rect 8208 3681 8232 3999
rect 8388 3921 8412 4119
rect 8448 4041 8472 4212
rect 8568 4041 8592 4212
rect 8148 3648 8172 3660
rect 7368 3528 7452 3552
rect 7608 3540 7632 3552
rect 7728 3540 7752 3552
rect 7128 3201 7152 3279
rect 7368 3081 7392 3528
rect 7599 3501 7641 3540
rect 7719 3501 7761 3540
rect 7788 3528 7872 3552
rect 6768 2481 6792 2652
rect 6768 2241 6792 2439
rect 5028 741 5052 879
rect 5148 861 5172 1359
rect 5448 1188 5472 1359
rect 5928 1188 5952 1299
rect 5208 1041 5232 1182
rect 5388 1080 5412 1092
rect 5379 1041 5421 1080
rect 5988 981 6012 1092
rect 6108 1041 6132 1539
rect 6168 1224 6192 2079
rect 6288 1980 6312 1992
rect 6279 1941 6321 1980
rect 6408 1821 6432 1992
rect 6339 1200 6381 1239
rect 6528 1212 6552 1959
rect 6588 1941 6612 2199
rect 6648 1998 6672 2139
rect 6741 2112 6780 2121
rect 6741 2088 6792 2112
rect 6888 2088 6912 2199
rect 6741 2079 6780 2088
rect 6828 1281 6852 1659
rect 7068 1641 7092 2199
rect 7128 2121 7152 2259
rect 7188 2088 7212 2379
rect 7308 2352 7332 2739
rect 7368 2661 7392 2859
rect 7548 2748 7572 3159
rect 7599 2841 7641 2859
rect 7668 2784 7692 2919
rect 7248 2328 7332 2352
rect 7248 2181 7272 2328
rect 7308 2088 7332 2199
rect 7428 2121 7452 2439
rect 7248 1881 7272 1992
rect 7488 1881 7512 2652
rect 7788 2601 7812 3528
rect 7908 3201 7932 3639
rect 7899 2760 7941 2799
rect 7908 2748 7932 2760
rect 8028 2748 8052 3159
rect 8088 2961 8112 3552
rect 8268 3501 8292 3879
rect 8268 2658 8292 3459
rect 8328 2772 8352 3819
rect 8628 3792 8652 4179
rect 8688 4161 8712 5076
rect 8748 4821 8772 5499
rect 8988 5361 9012 5679
rect 9048 5541 9072 5862
rect 9468 5781 9492 5868
rect 9168 5721 9192 5772
rect 9141 5688 9192 5721
rect 9141 5679 9180 5688
rect 8988 5208 9012 5319
rect 8808 4941 8832 5199
rect 8928 4701 8952 5112
rect 8781 4332 8820 4341
rect 8781 4308 8832 4332
rect 8919 4320 8961 4359
rect 9108 4341 9132 5559
rect 9228 5208 9252 5379
rect 9288 5301 9312 5772
rect 9348 5361 9372 5619
rect 9348 5208 9372 5319
rect 9468 5001 9492 5619
rect 9228 4401 9252 4839
rect 8928 4308 8952 4320
rect 8781 4299 8820 4308
rect 9219 4320 9261 4359
rect 9228 4308 9252 4320
rect 9528 4341 9552 6519
rect 9648 6321 9672 6639
rect 9708 6561 9732 8028
rect 9828 7641 9852 8019
rect 9888 7821 9912 8199
rect 9948 8181 9972 8232
rect 9948 7941 9972 8139
rect 9948 7632 9972 7719
rect 10008 7701 10032 8199
rect 10128 7941 10152 8232
rect 9948 7608 10032 7632
rect 9879 7440 9921 7479
rect 10008 7464 10032 7608
rect 9888 7428 9912 7440
rect 10068 7461 10092 7599
rect 9948 7320 9972 7332
rect 9939 7281 9981 7320
rect 10128 6981 10152 7779
rect 10188 7464 10212 8199
rect 10248 7641 10272 8379
rect 10308 8361 10332 9579
rect 10368 8898 10392 9099
rect 10608 8988 10632 9159
rect 10788 8898 10812 9279
rect 10968 8988 10992 9699
rect 11148 9381 11172 9792
rect 11388 9321 11412 9888
rect 11628 9888 11652 9999
rect 11808 9798 11832 9939
rect 11988 9888 12012 10059
rect 12168 9921 12192 10239
rect 11928 9780 11952 9792
rect 11919 9741 11961 9780
rect 11619 9672 11661 9699
rect 11541 9660 11661 9672
rect 11979 9681 12021 9699
rect 11541 9648 11652 9660
rect 11508 9441 11532 9519
rect 11448 9024 11472 9219
rect 10368 8328 10392 8559
rect 10428 8220 10452 8232
rect 10419 8181 10461 8220
rect 10668 7521 10692 8892
rect 10728 7821 10752 8799
rect 11028 8601 11052 8892
rect 11208 8868 11259 8892
rect 11208 8721 11232 8868
rect 11448 8661 11472 8982
rect 11508 8892 11532 9399
rect 12168 9381 12192 9759
rect 12228 9561 12252 10359
rect 12528 9981 12552 10719
rect 12648 10161 12672 11256
rect 12708 11181 12732 11988
rect 12768 11481 12792 11919
rect 13008 11328 13092 11352
rect 12708 10581 12732 11139
rect 13068 11001 13092 11328
rect 12768 10548 12792 10839
rect 13008 10452 13032 10899
rect 13128 10761 13152 12219
rect 13188 12141 13212 13059
rect 13248 12261 13272 14259
rect 13428 13821 13452 14259
rect 13488 14001 13512 14139
rect 13368 13704 13392 13779
rect 13488 13668 13512 13959
rect 13548 13761 13572 14139
rect 13608 13881 13632 14259
rect 13428 13281 13452 13572
rect 13548 13548 13632 13572
rect 13368 13041 13392 13179
rect 13341 13008 13392 13041
rect 13488 13008 13512 13359
rect 13548 13161 13572 13299
rect 13608 13161 13632 13548
rect 13668 13101 13692 14379
rect 13728 14361 13752 14472
rect 13848 14061 13872 14472
rect 13908 14181 13932 14439
rect 13968 14301 13992 14679
rect 14028 14601 14052 14748
rect 14088 14661 14112 14928
rect 14148 14661 14172 14859
rect 14208 14841 14232 14919
rect 14328 14841 14352 15039
rect 14148 14622 14199 14661
rect 14388 14601 14412 15099
rect 14568 15021 14592 15132
rect 14388 14568 14439 14601
rect 14400 14559 14439 14568
rect 14028 14361 14052 14496
rect 14208 14412 14232 14472
rect 14148 14388 14232 14412
rect 13728 13701 13752 13779
rect 13848 13668 13872 13956
rect 13959 13881 14001 13899
rect 13908 13761 13932 13839
rect 13980 13692 14019 13701
rect 13968 13668 14019 13692
rect 13980 13659 14019 13668
rect 13761 13572 13800 13581
rect 13761 13548 13812 13572
rect 13761 13539 13800 13548
rect 13341 12999 13380 13008
rect 13668 12921 13692 12996
rect 13728 12921 13752 13419
rect 13788 13341 13812 13479
rect 13848 13281 13872 13419
rect 13908 13341 13932 13572
rect 14088 13578 14112 14139
rect 14148 14121 14172 14388
rect 14208 13881 14232 14079
rect 14448 14061 14472 14439
rect 14508 13872 14532 14919
rect 14559 14592 14601 14619
rect 14748 14601 14772 15279
rect 14808 14721 14832 15459
rect 14979 15312 15021 15339
rect 14928 15300 15021 15312
rect 14928 15288 15012 15300
rect 14928 15228 14952 15288
rect 15048 15228 15072 15939
rect 15108 15561 15132 15879
rect 15168 15801 15192 16008
rect 15228 15861 15252 16359
rect 15408 16161 15432 16599
rect 15468 16341 15492 16479
rect 15468 16128 15492 16299
rect 15528 16161 15552 17499
rect 15588 17481 15612 17568
rect 15888 17481 15912 17559
rect 15588 17301 15612 17439
rect 15588 16641 15612 17019
rect 15708 16881 15732 17139
rect 15768 16788 15792 17079
rect 15828 16821 15852 16959
rect 15888 16941 15912 17199
rect 15948 17121 15972 17682
rect 15948 16761 15972 17079
rect 15681 16668 15732 16692
rect 15588 16461 15612 16536
rect 14559 14580 14652 14592
rect 14568 14568 14652 14580
rect 14628 14061 14652 14319
rect 14688 14301 14712 14436
rect 14448 13860 14532 13872
rect 14439 13848 14532 13860
rect 14439 13821 14481 13848
rect 13779 13101 13821 13119
rect 13848 13032 13872 13239
rect 13908 13221 13932 13299
rect 13968 13281 13992 13479
rect 14028 13461 14052 13539
rect 14088 13101 14112 13536
rect 14019 13044 14061 13059
rect 13788 13008 13872 13032
rect 13428 12741 13452 12912
rect 13548 12900 13572 12912
rect 13539 12861 13581 12900
rect 13788 12861 13812 13008
rect 14148 13041 14172 13719
rect 14208 13641 14232 13776
rect 14208 13281 14232 13599
rect 14388 13428 14472 13452
rect 13968 12900 13992 12912
rect 13239 12120 13281 12156
rect 13248 12108 13272 12120
rect 13368 12108 13392 12339
rect 13548 12012 13572 12639
rect 13668 12108 13692 12339
rect 13848 12141 13872 12879
rect 13959 12861 14001 12900
rect 13908 12441 13932 12819
rect 13188 11301 13212 11979
rect 13248 11484 13272 11799
rect 13308 11721 13332 12012
rect 13428 12000 13512 12012
rect 13428 11988 13521 12000
rect 13548 11988 13632 12012
rect 13479 11961 13521 11988
rect 13248 11181 13272 11442
rect 13608 11352 13632 11988
rect 13701 11940 13812 11952
rect 13701 11928 13821 11940
rect 13779 11901 13821 11928
rect 13668 11481 13692 11856
rect 13848 11661 13872 11979
rect 13908 11961 13932 12336
rect 13968 12321 13992 12819
rect 14028 12381 14052 12819
rect 14208 12501 14232 13176
rect 14268 12861 14292 13359
rect 14328 13221 14352 13419
rect 14388 13152 14412 13428
rect 14448 13161 14472 13359
rect 14328 13140 14412 13152
rect 14319 13128 14412 13140
rect 14319 13101 14361 13128
rect 14688 13044 14712 13719
rect 14808 13668 14832 14559
rect 14868 13761 14892 14919
rect 14988 14604 15012 14799
rect 15108 14781 15132 15099
rect 15168 15081 15192 15639
rect 15228 14601 15252 15579
rect 15288 15261 15312 15999
rect 15348 15501 15372 16032
rect 15408 15312 15432 15699
rect 15588 15381 15612 16179
rect 15648 16161 15672 16656
rect 15741 16632 15780 16641
rect 15741 16599 15792 16632
rect 15708 16221 15732 16359
rect 15768 16281 15792 16599
rect 15699 16140 15741 16179
rect 15819 16140 15861 16179
rect 15708 16128 15732 16140
rect 15828 16128 15852 16140
rect 15561 15348 15612 15381
rect 15561 15339 15600 15348
rect 15381 15288 15432 15312
rect 15348 15228 15372 15279
rect 15459 15240 15501 15279
rect 15579 15261 15621 15279
rect 15468 15228 15492 15240
rect 14928 13821 14952 14439
rect 14988 13752 15012 14379
rect 15048 14181 15072 14472
rect 15168 14460 15192 14472
rect 15159 14421 15201 14460
rect 15228 13992 15252 14439
rect 15168 13968 15252 13992
rect 15168 13761 15192 13968
rect 14928 13728 15012 13752
rect 14928 13668 14952 13728
rect 15228 13701 15252 13899
rect 15288 13881 15312 15099
rect 15408 14901 15432 15132
rect 15348 14478 15372 14739
rect 15468 14601 15492 15039
rect 15528 14661 15552 15096
rect 15648 14961 15672 15819
rect 15948 15681 15972 16479
rect 16008 16401 16032 18579
rect 16779 18441 16821 18459
rect 16461 18408 16539 18432
rect 16299 18360 16341 18399
rect 16308 18348 16332 18360
rect 16659 18360 16701 18399
rect 16779 18381 16821 18399
rect 16668 18348 16692 18360
rect 16128 18021 16152 18219
rect 16248 18141 16272 18252
rect 16428 18081 16452 18219
rect 16248 17688 16272 17979
rect 16308 17580 16332 17592
rect 16299 17541 16341 17580
rect 16428 17481 16452 17682
rect 16368 17121 16392 17319
rect 16428 17181 16452 17439
rect 16488 16761 16512 17799
rect 16608 17724 16632 17859
rect 16548 17301 16572 17499
rect 16848 17112 16872 18519
rect 16908 17721 16932 18459
rect 16968 18141 16992 18699
rect 17448 18441 17472 18912
rect 17568 18801 17592 18912
rect 17747 18888 17772 18912
rect 17079 18360 17121 18399
rect 17088 18348 17112 18360
rect 17508 18348 17532 18519
rect 17268 18240 17292 18252
rect 17259 18201 17301 18240
rect 17208 17961 17232 18099
rect 17388 18021 17412 18279
rect 16968 17688 16992 17859
rect 17088 17688 17112 17799
rect 16908 17172 16932 17559
rect 17028 17421 17052 17556
rect 16908 17148 16992 17172
rect 16848 17088 16932 17112
rect 16248 16560 16272 16572
rect 16239 16521 16281 16560
rect 16008 16041 16032 16239
rect 16068 16161 16092 16239
rect 16179 16140 16221 16179
rect 16308 16164 16332 16539
rect 16488 16512 16512 16656
rect 16548 16641 16572 16779
rect 16488 16488 16572 16512
rect 16188 16128 16212 16140
rect 16488 16128 16512 16359
rect 16548 16212 16572 16488
rect 16608 16281 16632 17079
rect 16848 16821 16872 17019
rect 16548 16188 16632 16212
rect 16608 16128 16632 16188
rect 16728 16161 16752 16599
rect 16248 15861 16272 15996
rect 16248 15741 16272 15819
rect 15768 15264 15792 15579
rect 16128 15561 16152 15639
rect 16188 15261 16212 15519
rect 15828 15072 15852 15132
rect 15801 15048 15852 15072
rect 15699 14580 15741 14619
rect 15768 14601 15792 15039
rect 15948 15021 15972 15132
rect 16008 14961 16032 15099
rect 16068 14901 16092 15222
rect 16128 14961 16152 15222
rect 16368 15261 16392 15459
rect 15999 14661 16041 14679
rect 15708 14568 15732 14580
rect 15339 14421 15381 14436
rect 15408 14361 15432 14559
rect 15468 13941 15492 14439
rect 15648 14241 15672 14472
rect 15828 14478 15852 14619
rect 16008 14568 16032 14619
rect 16128 14568 16152 14799
rect 16248 14478 16272 14979
rect 15528 14001 15552 14199
rect 15648 13941 15672 14079
rect 14748 13341 14772 13539
rect 14988 13560 15012 13572
rect 14979 13521 15021 13560
rect 14748 13008 14772 13179
rect 14268 12018 14292 12099
rect 13968 11988 14052 12012
rect 13368 11340 13392 11352
rect 13359 11301 13401 11340
rect 13548 11328 13632 11352
rect 11628 8988 11652 9099
rect 11508 8868 11592 8892
rect 10221 7332 10260 7341
rect 10221 7308 10272 7332
rect 10221 7299 10260 7308
rect 9828 6621 9852 6759
rect 9648 5868 9672 6039
rect 9768 5904 9792 6459
rect 9948 6381 9972 6672
rect 10188 6201 10212 6762
rect 10248 6021 10272 6819
rect 10428 6801 10452 7299
rect 10488 6861 10512 7479
rect 10848 7428 10872 8019
rect 10908 7941 10932 8232
rect 10548 7281 10572 7359
rect 10668 7221 10692 7332
rect 10548 6792 10572 6939
rect 10488 6768 10572 6792
rect 10368 6261 10392 6672
rect 10368 6072 10392 6219
rect 10368 6048 10452 6072
rect 10068 5904 10092 5979
rect 10128 5868 10152 5979
rect 9588 4401 9612 5736
rect 9888 5721 9912 5862
rect 9888 5601 9912 5679
rect 10188 5481 10212 5772
rect 9768 5244 9792 5319
rect 10008 5121 10032 5379
rect 10368 5241 10392 5979
rect 9708 4881 9732 5112
rect 10428 5118 10452 6048
rect 10548 6021 10572 6639
rect 10608 6621 10632 6879
rect 10788 6861 10812 7332
rect 10968 7041 10992 7479
rect 11028 7341 11052 8232
rect 11088 7941 11112 8196
rect 11148 7452 11172 8319
rect 11208 7524 11232 8559
rect 11268 8061 11292 8439
rect 11328 8361 11352 8619
rect 11268 7641 11292 7779
rect 11088 7428 11172 7452
rect 11088 7032 11112 7428
rect 11328 7428 11352 7659
rect 11508 7461 11532 8196
rect 11568 8121 11592 8868
rect 11808 8328 11832 8439
rect 11928 8421 11952 8988
rect 11988 8901 12012 9159
rect 12048 9021 12072 9279
rect 12288 9021 12312 9939
rect 12888 9924 12912 10452
rect 13008 10428 13092 10452
rect 13068 9921 13092 10428
rect 13248 10440 13272 10452
rect 12348 9681 12372 9756
rect 11988 8352 12012 8679
rect 11928 8328 12012 8352
rect 11628 8241 11652 8322
rect 11508 7041 11532 7419
rect 11088 7008 11172 7032
rect 10668 6141 10692 6819
rect 10848 6804 10872 6999
rect 10728 6321 10752 6579
rect 10788 6561 10812 6672
rect 11148 6501 11172 7008
rect 10548 5868 10572 5979
rect 10659 5880 10701 5919
rect 10668 5868 10692 5880
rect 10788 5868 10812 6219
rect 10908 5778 10932 5919
rect 10608 5661 10632 5736
rect 10728 5601 10752 5772
rect 10761 5568 10812 5592
rect 10479 5244 10521 5259
rect 10719 5241 10761 5259
rect 9768 4521 9792 4779
rect 8601 3768 8652 3792
rect 8568 3648 8592 3759
rect 8748 3684 8772 4179
rect 9021 4188 9072 4212
rect 8868 3648 8892 3999
rect 8748 3558 8772 3642
rect 8508 3540 8532 3552
rect 8388 3081 8412 3519
rect 8499 3501 8541 3540
rect 9048 3501 9072 4188
rect 9288 4101 9312 4212
rect 9108 3681 9132 3759
rect 9288 3741 9312 3879
rect 9408 3672 9432 4059
rect 9468 4041 9492 4302
rect 9579 4320 9621 4359
rect 9588 4308 9612 4320
rect 9828 4341 9852 4539
rect 9888 4221 9912 4359
rect 10008 4341 10032 5016
rect 10248 4701 10272 5079
rect 10308 4932 10332 5112
rect 10788 5118 10812 5568
rect 10968 5421 10992 6099
rect 11208 5892 11232 6999
rect 11568 6801 11592 7959
rect 11808 7632 11832 8079
rect 11868 7701 11892 8232
rect 11988 8001 12012 8199
rect 12048 7641 12072 8859
rect 12288 8661 12312 8859
rect 12348 8721 12372 9459
rect 12408 9261 12432 9792
rect 12408 8961 12432 9099
rect 12468 8841 12492 9639
rect 12648 9321 12672 9519
rect 12528 9012 12552 9159
rect 12708 9141 12732 9879
rect 12768 9801 12792 9882
rect 13008 9780 13032 9792
rect 12948 9261 12972 9759
rect 12999 9741 13041 9780
rect 13068 9441 13092 9759
rect 13128 9681 13152 9939
rect 13188 9741 13212 10419
rect 13239 10401 13281 10440
rect 13248 10221 13272 10359
rect 13308 10341 13332 10419
rect 13248 9801 13272 9999
rect 13368 9981 13392 11139
rect 13488 10941 13512 11199
rect 13548 10821 13572 11328
rect 13908 11181 13932 11856
rect 13968 11841 13992 11988
rect 13968 11241 13992 11799
rect 13608 10701 13632 10899
rect 13428 10581 13452 10659
rect 13608 10548 13632 10659
rect 13668 10581 13692 11139
rect 13428 10041 13452 10419
rect 13548 10221 13572 10452
rect 13668 10428 13752 10452
rect 13368 9780 13392 9792
rect 13359 9741 13401 9780
rect 13221 9738 13260 9741
rect 13221 9699 13239 9738
rect 13188 9201 13212 9636
rect 12528 8988 12612 9012
rect 12828 9021 12852 9099
rect 12108 8121 12132 8499
rect 12288 8361 12312 8619
rect 12528 8601 12552 8859
rect 12768 8880 12792 8892
rect 12759 8841 12801 8880
rect 12828 8661 12852 8859
rect 12888 8781 12912 9159
rect 13248 9081 13272 9339
rect 13308 9021 13332 9699
rect 13488 9381 13512 9792
rect 12768 8481 12792 8559
rect 12339 8340 12381 8379
rect 12348 8328 12372 8340
rect 12828 8361 12852 8619
rect 12948 8532 12972 8859
rect 13008 8781 13032 8892
rect 13128 8781 13152 8892
rect 13239 8832 13281 8859
rect 13188 8820 13281 8832
rect 13308 8868 13359 8892
rect 13188 8808 13272 8820
rect 12888 8508 12972 8532
rect 11808 7608 11892 7632
rect 11748 7221 11772 7332
rect 11868 7161 11892 7608
rect 12048 7512 12072 7599
rect 11988 7488 12072 7512
rect 11988 7428 12012 7488
rect 12099 7440 12141 7479
rect 12228 7461 12252 7719
rect 12108 7428 12132 7440
rect 12168 7320 12192 7332
rect 12159 7281 12201 7320
rect 11628 6801 11652 6879
rect 11799 6780 11841 6819
rect 11808 6768 11832 6780
rect 12048 6801 12072 7119
rect 11328 6441 11352 6672
rect 11628 6501 11652 6696
rect 11688 6432 11712 6639
rect 11748 6561 11772 6672
rect 11808 6501 11832 6579
rect 12048 6561 12072 6639
rect 11601 6408 11712 6432
rect 11748 5961 11772 6339
rect 11208 5868 11292 5892
rect 11148 5541 11172 5736
rect 10308 4908 10392 4932
rect 10299 4581 10341 4599
rect 9408 3648 9492 3672
rect 9141 3552 9180 3561
rect 9141 3528 9192 3552
rect 9141 3519 9180 3528
rect 8328 2748 8412 2772
rect 8508 2748 8532 2919
rect 8688 2901 8712 3099
rect 9408 3021 9432 3519
rect 9468 3141 9492 3648
rect 7668 2088 7692 2259
rect 7728 1641 7752 1992
rect 7068 1461 7092 1599
rect 6639 1221 6681 1239
rect 6348 1188 6372 1200
rect 6468 1188 6612 1212
rect 6588 1098 6612 1188
rect 6819 1200 6861 1239
rect 6828 1188 6852 1200
rect 7128 1101 7152 1299
rect 7368 1188 7392 1299
rect 7848 1101 7872 1299
rect 6558 1056 6561 1080
rect 6519 1041 6561 1056
rect 5988 948 6039 981
rect 6000 939 6039 948
rect 6201 939 6219 981
rect 5301 879 5319 921
rect 4788 321 4812 432
rect 4968 321 4992 579
rect 5088 528 5112 639
rect 5208 564 5232 879
rect 5988 681 6012 819
rect 5268 420 5292 432
rect 5148 201 5172 396
rect 5259 381 5301 420
rect 5388 261 5412 639
rect 5808 321 5832 519
rect 5868 438 5892 579
rect 6048 528 6072 759
rect 6288 441 6312 639
rect 6348 438 6372 759
rect 7308 741 7332 1092
rect 6519 540 6561 579
rect 6528 528 6552 540
rect 6648 528 6672 639
rect 6768 438 6792 699
rect 7281 648 7359 672
rect 7299 540 7341 579
rect 7308 528 7332 540
rect 7668 561 7692 759
rect 6219 381 6261 396
rect 6408 141 6432 399
rect 6579 381 6621 396
rect 7068 321 7092 522
rect 7500 432 7539 441
rect 7248 201 7272 339
rect 7368 321 7392 432
rect 7488 408 7539 432
rect 7500 399 7539 408
rect 7608 381 7632 522
rect 7788 528 7812 819
rect 7908 621 7932 2559
rect 7968 1701 7992 2379
rect 8088 2301 8112 2652
rect 8079 2172 8121 2196
rect 8079 2160 8139 2172
rect 8088 2148 8139 2160
rect 8148 2088 8172 2139
rect 8268 2088 8412 2112
rect 8208 1761 8232 1992
rect 7968 1101 7992 1539
rect 8139 1200 8181 1239
rect 8268 1224 8292 1359
rect 8388 1281 8412 2088
rect 8448 2001 8472 2652
rect 8688 2088 8712 2859
rect 8988 2748 9012 2859
rect 9168 2658 9192 2919
rect 9348 2784 9372 2859
rect 8928 2481 8952 2652
rect 9408 2421 9432 2499
rect 8919 2121 8961 2139
rect 8568 1341 8592 1956
rect 8748 1881 8772 1992
rect 8868 1761 8892 2079
rect 8988 1998 9012 2139
rect 9048 2121 9072 2199
rect 9159 2100 9201 2139
rect 9168 2088 9192 2100
rect 9468 2061 9492 3036
rect 9528 2658 9552 4179
rect 9588 3681 9612 3999
rect 9648 3741 9672 4179
rect 9858 4176 9861 4200
rect 9819 4161 9861 4176
rect 9948 4101 9972 4302
rect 10239 4341 10281 4359
rect 10308 4221 10332 4539
rect 9708 3648 9732 3759
rect 9828 3648 9972 3672
rect 9588 3081 9612 3459
rect 9759 2760 9801 2799
rect 9948 2784 9972 3648
rect 10008 3621 10032 3819
rect 10248 3741 10272 4179
rect 10308 3648 10332 4116
rect 10368 3861 10392 4908
rect 10488 4641 10512 5079
rect 10668 4941 10692 5112
rect 10848 5112 10872 5319
rect 11001 5292 11040 5301
rect 11001 5259 11052 5292
rect 11028 5208 11052 5259
rect 10848 5088 10992 5112
rect 11148 5088 11232 5112
rect 10548 4308 10572 4479
rect 10428 4101 10452 4302
rect 10848 4221 10872 4659
rect 10908 4461 10932 5088
rect 10968 4308 10992 4779
rect 11208 4521 11232 5088
rect 10479 4161 10521 4179
rect 10428 3681 10452 4059
rect 10608 3921 10632 4212
rect 10728 4101 10752 4212
rect 11028 4101 11052 4212
rect 10068 2841 10092 3639
rect 10488 3558 10512 3699
rect 10599 3660 10641 3699
rect 10608 3648 10632 3660
rect 10728 3648 10752 3759
rect 10848 3681 10872 3879
rect 10908 3558 10932 4059
rect 11028 3648 11052 4059
rect 11148 3681 11172 4179
rect 10368 3441 10392 3552
rect 9768 2748 9792 2760
rect 9888 2748 9939 2772
rect 10068 2748 10092 2799
rect 10668 2748 10692 2979
rect 10788 2748 10812 3099
rect 10968 2841 10992 3519
rect 11088 3441 11112 3516
rect 11208 3501 11232 4479
rect 11268 3192 11292 5868
rect 11328 4344 11352 5619
rect 11448 5601 11472 5772
rect 11388 5241 11412 5379
rect 11568 5361 11592 5772
rect 11688 5661 11712 5862
rect 11748 5292 11772 5919
rect 11868 5904 11892 6519
rect 11988 5868 12012 6219
rect 12108 5781 12132 6762
rect 11928 5661 11952 5772
rect 12168 5601 12192 6999
rect 12228 6801 12252 7296
rect 12288 6861 12312 7599
rect 12468 7521 12492 8319
rect 12648 8121 12672 8232
rect 12768 8061 12792 8232
rect 12348 7341 12372 7479
rect 12528 7428 12552 7839
rect 12828 7464 12852 8199
rect 12468 7320 12492 7332
rect 12459 7281 12501 7320
rect 12588 7101 12612 7332
rect 12888 7041 12912 8508
rect 12948 7641 12972 8439
rect 13008 7761 13032 8619
rect 13188 8328 13212 8808
rect 13308 8661 13332 8868
rect 13548 8481 13572 9399
rect 13608 8721 13632 10359
rect 13668 9981 13692 10428
rect 13908 10401 13932 10779
rect 13968 10452 13992 11079
rect 14028 10581 14052 11919
rect 14328 10941 14352 12879
rect 14568 12801 14592 12912
rect 14868 12801 14892 12879
rect 14388 12561 14412 12639
rect 14388 11841 14412 12456
rect 14508 12144 14532 12639
rect 14628 12108 14652 12279
rect 14688 12141 14712 12759
rect 14808 12381 14832 12459
rect 14928 12261 14952 12999
rect 14988 12681 15012 13059
rect 15048 13041 15072 13539
rect 15108 13101 15132 13599
rect 15168 13521 15192 13656
rect 15168 13008 15192 13119
rect 15228 13101 15252 13539
rect 15288 13461 15312 13572
rect 15408 13341 15432 13572
rect 15288 13044 15312 13299
rect 15348 13041 15372 13119
rect 15048 12381 15072 12879
rect 15108 12741 15132 12912
rect 15168 12561 15192 12759
rect 15228 12441 15252 12912
rect 14508 11448 14532 11919
rect 14568 11901 14592 12012
rect 14388 11328 14472 11352
rect 14388 10821 14412 11328
rect 14088 10548 14112 10659
rect 13968 10428 14052 10452
rect 13728 9924 13752 10119
rect 13839 9900 13881 9939
rect 13848 9888 13872 9900
rect 13668 9681 13692 9759
rect 13908 9681 13932 9792
rect 14028 9621 14052 10428
rect 14388 10428 14472 10452
rect 14088 9681 14112 10359
rect 14388 10341 14412 10428
rect 14628 10212 14652 11799
rect 14748 11781 14772 11979
rect 14688 11472 14712 11619
rect 14988 11541 15012 11892
rect 15048 11601 15072 11739
rect 15228 11661 15252 12219
rect 15288 12018 15312 12819
rect 15408 12321 15432 13179
rect 15528 13032 15552 13539
rect 15588 13221 15612 13839
rect 15648 13341 15672 13899
rect 15501 13008 15552 13032
rect 15639 13044 15681 13059
rect 15708 13032 15732 14379
rect 15768 14241 15792 14439
rect 16068 14361 16092 14472
rect 15768 14001 15792 14079
rect 16068 13821 16092 13959
rect 15939 13680 15981 13719
rect 16128 13701 16152 14199
rect 16248 13821 16272 14436
rect 15948 13668 15972 13680
rect 16248 13668 16272 13779
rect 16308 13761 16332 14919
rect 16359 14601 16401 14619
rect 16428 14568 16452 15339
rect 16488 15261 16512 15879
rect 16548 15228 16572 15579
rect 16728 15312 16752 15999
rect 16788 15501 16812 16419
rect 16908 16332 16932 17088
rect 16968 16461 16992 17148
rect 17028 16821 17052 17379
rect 17148 17301 17172 17556
rect 17268 17121 17292 17979
rect 17388 17688 17412 17916
rect 17568 17901 17592 18252
rect 17448 17421 17472 17592
rect 17568 17481 17592 17592
rect 17148 16788 17172 17019
rect 17508 16824 17532 16899
rect 17568 16872 17592 17079
rect 17628 16941 17652 17559
rect 17688 17541 17712 18639
rect 17748 18381 17772 18888
rect 18008 18681 18032 18912
rect 17799 18360 17841 18399
rect 17808 18348 17832 18360
rect 17568 16848 17652 16872
rect 17628 16788 17652 16848
rect 17061 16692 17100 16701
rect 17061 16668 17112 16692
rect 17208 16680 17232 16692
rect 17061 16659 17100 16668
rect 17199 16641 17241 16680
rect 17421 16668 17472 16692
rect 16848 16308 16932 16332
rect 16848 15432 16872 16308
rect 17208 16281 17232 16599
rect 16908 16161 16932 16239
rect 17088 16128 17112 16239
rect 17388 16221 17412 16659
rect 17748 16692 17772 18219
rect 17808 17841 17832 17919
rect 17868 17724 17892 18159
rect 17928 18021 17952 18252
rect 17928 17772 17952 17979
rect 17928 17748 18012 17772
rect 17988 17688 18012 17748
rect 18108 17601 18132 17799
rect 17808 16701 17832 17019
rect 17688 16668 17772 16692
rect 17508 16452 17532 16539
rect 17508 16428 17592 16452
rect 17439 16332 17481 16359
rect 17439 16320 17532 16332
rect 17448 16308 17532 16320
rect 17028 15921 17052 16032
rect 17148 15861 17172 16032
rect 17208 15621 17232 15999
rect 17268 15801 17292 16179
rect 17379 16140 17421 16179
rect 17508 16161 17532 16308
rect 17388 16128 17412 16140
rect 17568 16041 17592 16428
rect 17028 15441 17052 15519
rect 16848 15408 16932 15432
rect 16668 15288 16752 15312
rect 16668 15228 16692 15288
rect 16848 15138 16872 15339
rect 16608 14952 16632 15096
rect 16608 14928 16692 14952
rect 16668 14601 16692 14928
rect 16368 13704 16392 14439
rect 16428 13701 16452 14079
rect 16608 13941 16632 14472
rect 16668 14121 16692 14439
rect 16728 13881 16752 14619
rect 16788 14601 16812 14799
rect 16848 14661 16872 15096
rect 16908 14721 16932 15408
rect 17028 15228 17052 15399
rect 17328 15132 17352 15699
rect 17208 15021 17232 15132
rect 17268 15108 17352 15132
rect 16848 14568 16872 14619
rect 16968 14568 16992 14919
rect 17088 14601 17112 14859
rect 17148 14781 17172 14919
rect 17268 14901 17292 15108
rect 17388 14841 17412 15819
rect 17448 14901 17472 15879
rect 17628 15741 17652 16539
rect 17688 15921 17712 16668
rect 17868 16581 17892 17499
rect 17988 16788 18012 16899
rect 18228 16701 18252 18759
rect 17868 16128 17892 16239
rect 17568 15264 17592 15399
rect 17988 15381 18012 16419
rect 18048 15861 18072 16659
rect 18108 16341 18132 16692
rect 18288 16461 18312 17559
rect 18288 16128 18312 16299
rect 18348 16161 18372 17859
rect 18168 15912 18192 16032
rect 18108 15888 18192 15912
rect 18108 15621 18132 15888
rect 18168 15681 18192 15819
rect 17961 15312 18000 15321
rect 17961 15279 18012 15312
rect 17679 15240 17721 15279
rect 17688 15228 17712 15240
rect 17988 15228 18012 15279
rect 17628 15021 17652 15132
rect 17748 15120 17832 15132
rect 17748 15108 17841 15120
rect 17799 15081 17841 15108
rect 16908 14361 16932 14436
rect 17028 14421 17052 14472
rect 16968 14388 17019 14412
rect 16968 14061 16992 14388
rect 17088 14352 17112 14439
rect 17028 14328 17112 14352
rect 15768 13461 15792 13539
rect 15708 13008 15792 13032
rect 15468 12741 15492 12999
rect 15528 12681 15552 12879
rect 15339 12141 15381 12159
rect 15459 12120 15501 12159
rect 15528 12132 15552 12279
rect 15588 12201 15612 12912
rect 15768 12861 15792 13008
rect 15828 12921 15852 13119
rect 15888 13101 15912 13572
rect 16008 13401 16032 13572
rect 16068 13041 16092 13539
rect 16188 13521 16212 13572
rect 16308 13512 16332 13572
rect 16248 13488 16332 13512
rect 15948 12741 15972 12876
rect 16068 12381 16092 12879
rect 16128 12621 16152 13419
rect 16188 13341 16212 13479
rect 16248 13044 16272 13488
rect 16428 13461 16452 13539
rect 16488 13041 16512 13659
rect 16548 13401 16572 13839
rect 16668 13668 16692 13779
rect 16908 13701 16932 13959
rect 16308 12441 16332 12912
rect 15468 12108 15492 12120
rect 15528 12108 15612 12132
rect 15348 11901 15372 11979
rect 15288 11721 15312 11799
rect 14688 11448 14772 11472
rect 14859 11460 14901 11499
rect 14868 11448 14892 11460
rect 14688 10821 14712 11316
rect 14568 10188 14652 10212
rect 14208 9888 14232 9999
rect 14328 9888 14352 10059
rect 14448 9921 14472 10179
rect 14400 9792 14439 9801
rect 14388 9768 14439 9792
rect 14400 9759 14439 9768
rect 14508 9732 14532 9939
rect 14448 9708 14532 9732
rect 13908 8988 13932 9099
rect 13968 9021 13992 9219
rect 14028 8868 14079 8892
rect 13668 8781 13692 8859
rect 13608 8541 13632 8679
rect 13668 8328 13692 8439
rect 13248 8172 13272 8232
rect 13188 8148 13272 8172
rect 13188 7761 13212 8148
rect 13080 7512 13119 7521
rect 13068 7479 13119 7512
rect 13068 7428 13092 7479
rect 13188 7461 13212 7656
rect 12861 7008 12912 7041
rect 12948 7308 12999 7332
rect 12861 6999 12900 7008
rect 12348 6768 12372 6939
rect 12468 6768 12492 6939
rect 12288 6660 12312 6672
rect 12228 6381 12252 6639
rect 12279 6621 12321 6660
rect 12288 5961 12312 6579
rect 12408 6012 12432 6636
rect 12348 5988 12432 6012
rect 12348 5868 12372 5988
rect 12468 5868 12492 6039
rect 12519 5961 12561 5979
rect 11748 5268 11832 5292
rect 11808 5244 11832 5268
rect 11928 5241 11952 5556
rect 11388 4581 11412 5079
rect 11448 4821 11472 5112
rect 11688 4992 11712 5202
rect 11628 4968 11712 4992
rect 11328 3681 11352 4119
rect 11388 4101 11412 4212
rect 11568 4101 11592 4779
rect 11628 4041 11652 4968
rect 11748 4881 11772 5079
rect 11868 4401 11892 5112
rect 11928 4344 11952 5079
rect 11988 4332 12012 5379
rect 12168 5301 12192 5496
rect 12408 5412 12432 5772
rect 12408 5388 12492 5412
rect 12228 5208 12252 5379
rect 12408 5118 12432 5319
rect 12468 5241 12492 5388
rect 12588 5301 12612 6939
rect 12648 6261 12672 6819
rect 12888 6768 12912 6939
rect 12948 6801 12972 7308
rect 13248 7338 13272 8079
rect 13308 7941 13332 8199
rect 13368 7881 13392 8319
rect 13488 7701 13512 8232
rect 13608 7761 13632 8196
rect 13728 8121 13752 8199
rect 13368 7464 13392 7599
rect 13488 7428 13512 7539
rect 13788 7524 13812 8559
rect 13968 8481 13992 8859
rect 14028 8652 14052 8868
rect 14028 8628 14112 8652
rect 14028 8328 14052 8559
rect 14088 8361 14112 8628
rect 14268 8601 14292 9579
rect 14328 8541 14352 9639
rect 14388 9021 14412 9339
rect 14448 8988 14472 9708
rect 14568 9321 14592 10188
rect 14688 10101 14712 10659
rect 14808 10548 14832 11253
rect 15048 11241 15072 11559
rect 15108 11061 15132 11499
rect 15588 11472 15612 12108
rect 15648 11781 15672 12339
rect 15879 12120 15921 12159
rect 15888 12108 15912 12120
rect 15960 12012 15999 12021
rect 15708 11601 15732 11979
rect 15828 11901 15852 12012
rect 15948 11988 15999 12012
rect 15960 11979 15999 11988
rect 15528 11448 15612 11472
rect 15048 10881 15072 10959
rect 15168 10872 15192 11319
rect 15228 11121 15252 11352
rect 15408 11328 15492 11352
rect 15108 10848 15192 10872
rect 15048 10692 15072 10839
rect 14988 10668 15072 10692
rect 14988 10590 15012 10668
rect 15108 10581 15132 10848
rect 15108 10428 15159 10452
rect 15048 10212 15072 10419
rect 14988 10188 15072 10212
rect 14619 9921 14661 9939
rect 14739 9900 14781 9939
rect 14748 9888 14772 9900
rect 14628 9768 14712 9792
rect 14628 9561 14652 9768
rect 14928 9792 14952 9879
rect 14799 9741 14841 9756
rect 14868 9768 14952 9792
rect 14868 9561 14892 9768
rect 14628 9030 14652 9099
rect 14688 9081 14712 9459
rect 14688 8721 14712 8856
rect 14088 7932 14112 8199
rect 14148 7941 14172 8439
rect 14028 7908 14112 7932
rect 13848 7641 13872 7779
rect 13908 7581 13932 7839
rect 13068 7161 13092 7239
rect 13008 6321 13032 7059
rect 13068 6801 13092 7119
rect 13188 6768 13212 7299
rect 13608 7041 13632 7359
rect 13428 6792 13452 6999
rect 13428 6768 13512 6792
rect 13128 6501 13152 6672
rect 13248 6261 13272 6672
rect 13368 6381 13392 6672
rect 13428 6081 13452 6639
rect 12648 5988 12759 6012
rect 12648 5901 12672 5988
rect 12699 5880 12741 5919
rect 12708 5868 12732 5880
rect 12948 5901 12972 5979
rect 13008 5841 13032 5919
rect 12888 5661 12912 5772
rect 12648 5232 12672 5619
rect 12588 5208 12672 5232
rect 12288 5100 12312 5112
rect 12279 5061 12321 5100
rect 11988 4308 12072 4332
rect 11748 3981 11772 4176
rect 11868 4101 11892 4212
rect 12048 3801 12072 4308
rect 12108 4218 12132 5019
rect 12468 5001 12492 5079
rect 12708 5100 12732 5112
rect 12699 5061 12741 5100
rect 12528 3861 12552 4539
rect 12828 4461 12852 5559
rect 12948 5481 12972 5739
rect 13128 5760 13152 5772
rect 12999 5721 13041 5736
rect 13068 5361 13092 5739
rect 13119 5721 13161 5760
rect 13248 5601 13272 5772
rect 12888 4701 12912 5259
rect 13248 5112 13272 5319
rect 13008 4881 13032 5112
rect 13068 4761 13092 4959
rect 13128 4821 13152 5112
rect 13188 5088 13272 5112
rect 12081 3768 12132 3792
rect 11361 3552 11400 3561
rect 11361 3528 11412 3552
rect 11508 3540 11532 3552
rect 11361 3519 11400 3528
rect 11499 3501 11541 3540
rect 11688 3501 11712 3759
rect 11868 3648 11892 3759
rect 12108 3558 12132 3768
rect 12348 3648 12372 3759
rect 11268 3168 11352 3192
rect 10908 2808 10959 2832
rect 10908 2721 10932 2808
rect 11028 2748 11052 2979
rect 11139 2760 11181 2799
rect 11268 2781 11292 3099
rect 11148 2748 11172 2760
rect 9708 2361 9732 2652
rect 9819 2601 9861 2616
rect 9999 2601 10041 2616
rect 9528 2121 9552 2319
rect 10248 2241 10272 2652
rect 9648 2088 9672 2199
rect 9768 2088 9792 2199
rect 10068 2088 10092 2199
rect 8148 1188 8172 1200
rect 8508 1188 8532 1299
rect 8619 1200 8661 1239
rect 8628 1188 8652 1200
rect 8928 1161 8952 1779
rect 9228 1341 9252 1992
rect 9348 1701 9372 1992
rect 9561 1998 9600 2001
rect 9561 1959 9579 1998
rect 9408 1821 9432 1959
rect 9828 1881 9852 1992
rect 10008 1881 10032 1992
rect 10128 1821 10152 1992
rect 10308 1941 10332 2079
rect 10368 1821 10392 2616
rect 10548 2088 10572 2499
rect 11208 2481 11232 2652
rect 10668 2241 10692 2439
rect 10668 2088 10692 2199
rect 10788 2001 10812 2439
rect 10848 2121 10872 2199
rect 10908 2088 10932 2319
rect 11019 2100 11061 2139
rect 11028 2088 11052 2100
rect 10488 1821 10512 1992
rect 11208 1998 11232 2139
rect 11268 2001 11292 2079
rect 11328 2061 11352 3168
rect 11388 2361 11412 3459
rect 11859 3441 11901 3459
rect 11508 2748 11532 2919
rect 11868 2661 11892 3219
rect 12108 2781 12132 2859
rect 12168 2784 12192 3639
rect 12288 3441 12312 3552
rect 12408 3540 12432 3552
rect 12399 3501 12441 3540
rect 12588 3441 12612 4419
rect 12759 4344 12801 4359
rect 12948 4332 12972 4479
rect 13188 4401 13212 5088
rect 13308 5061 13332 5679
rect 13428 5601 13452 5976
rect 13488 5721 13512 6339
rect 13668 6081 13692 7479
rect 13908 7428 13932 7539
rect 14028 7461 14052 7908
rect 14208 7872 14232 8499
rect 14448 8328 14472 8439
rect 14508 8361 14532 8559
rect 14748 8481 14772 9339
rect 14808 8901 14832 9459
rect 14928 9261 14952 9699
rect 14988 9681 15012 10188
rect 15108 10101 15132 10428
rect 15228 9888 15252 10179
rect 15039 9741 15081 9759
rect 14928 9141 14952 9219
rect 15048 9021 15072 9099
rect 14148 7848 14232 7872
rect 14088 7338 14112 7719
rect 13848 6852 13872 7332
rect 13968 7161 13992 7296
rect 14148 7281 14172 7848
rect 14268 7701 14292 8199
rect 14388 8121 14412 8232
rect 14568 8220 14592 8232
rect 14448 8061 14472 8139
rect 14448 7461 14472 8019
rect 14508 7521 14532 8199
rect 14559 8181 14601 8220
rect 14868 8181 14892 8979
rect 14928 8112 14952 8859
rect 15108 8841 15132 9639
rect 15168 9381 15192 9792
rect 15288 9501 15312 9759
rect 15348 9432 15372 10659
rect 15408 10221 15432 11199
rect 15468 11181 15492 11328
rect 15468 10581 15492 11019
rect 15528 10641 15552 11448
rect 15768 11361 15792 11739
rect 15828 11541 15852 11679
rect 15648 10881 15672 11352
rect 15828 11292 15852 11499
rect 15768 11268 15852 11292
rect 15768 11001 15792 11268
rect 15540 10572 15579 10581
rect 15528 10548 15579 10572
rect 15540 10539 15579 10548
rect 15768 10572 15792 10839
rect 15828 10821 15852 11199
rect 15708 10548 15792 10572
rect 15408 9621 15432 10059
rect 15468 9981 15492 10419
rect 15768 10221 15792 10419
rect 15828 10281 15852 10779
rect 15888 10701 15912 11619
rect 16128 11481 16152 12159
rect 16188 12141 16212 12399
rect 16428 12321 16452 12813
rect 16548 12561 16572 12999
rect 16608 12918 16632 13479
rect 16668 13041 16692 13479
rect 16728 13401 16752 13572
rect 16908 13281 16932 13539
rect 16788 13008 16812 13239
rect 16908 13008 16932 13119
rect 16968 13101 16992 13839
rect 17028 13041 17052 14328
rect 17148 13992 17172 14676
rect 17268 14661 17292 14739
rect 17508 14652 17532 14979
rect 17508 14640 17592 14652
rect 17508 14628 17601 14640
rect 17559 14601 17601 14628
rect 17259 14421 17301 14439
rect 17388 14361 17412 14472
rect 17088 13968 17172 13992
rect 16848 12900 16872 12912
rect 16839 12861 16881 12900
rect 16608 12201 16632 12399
rect 16668 12081 16692 12699
rect 15888 10458 15912 10596
rect 15648 9888 15672 9999
rect 15768 9888 15792 10116
rect 15948 10041 15972 11259
rect 16068 11241 16092 11352
rect 16188 10581 16212 12036
rect 16428 11601 16452 11892
rect 16248 11241 16272 11559
rect 16479 11460 16521 11499
rect 16488 11448 16512 11460
rect 16608 11481 16632 11559
rect 16581 11442 16632 11481
rect 16728 11472 16752 12519
rect 16788 12021 16812 12699
rect 16848 12141 16872 12219
rect 16908 12108 16932 12819
rect 16968 12681 16992 12912
rect 17028 12741 17052 12879
rect 17088 12201 17112 13968
rect 17508 13941 17532 14436
rect 17148 13761 17172 13899
rect 17148 13341 17172 13479
rect 17328 13221 17352 13452
rect 17148 13041 17172 13179
rect 17199 13020 17241 13059
rect 17208 13008 17232 13020
rect 17448 13041 17472 13299
rect 17508 12912 17532 13479
rect 17268 12900 17292 12912
rect 17388 12900 17412 12912
rect 17088 12132 17112 12159
rect 17028 12108 17112 12132
rect 16560 11439 16632 11442
rect 16428 11181 16452 11352
rect 16041 10572 16080 10581
rect 16041 10548 16092 10572
rect 16041 10539 16080 10548
rect 16299 10560 16341 10599
rect 16419 10560 16461 10599
rect 16308 10548 16332 10560
rect 16428 10548 16452 10560
rect 16008 10161 16032 10419
rect 15288 9408 15372 9432
rect 15168 8421 15192 9159
rect 15228 8781 15252 9279
rect 15141 8388 15192 8421
rect 15141 8379 15180 8388
rect 15108 8328 15219 8352
rect 14868 8100 14952 8112
rect 14859 8088 14952 8100
rect 14859 8061 14901 8088
rect 14619 7440 14661 7479
rect 14628 7428 14652 7440
rect 14748 7428 14772 8019
rect 14808 7452 14832 7779
rect 14868 7512 14892 7899
rect 14928 7728 15072 7752
rect 14928 7641 14952 7728
rect 14868 7488 14952 7512
rect 14808 7428 14892 7452
rect 14268 7320 14292 7332
rect 13848 6840 13932 6852
rect 13848 6828 13941 6840
rect 13899 6801 13941 6828
rect 13728 6672 13752 6762
rect 14148 6672 14172 6999
rect 13728 6648 13812 6672
rect 13788 6501 13812 6648
rect 14028 6648 14172 6672
rect 13848 6321 13872 6399
rect 13599 6012 13641 6039
rect 13599 6000 13692 6012
rect 13608 5988 13692 6000
rect 13668 5952 13692 5988
rect 13668 5928 13719 5952
rect 13599 5880 13641 5919
rect 13608 5868 13632 5880
rect 13728 5868 13752 5919
rect 13788 5901 13812 6219
rect 14148 6141 14172 6279
rect 13428 5208 13452 5439
rect 13548 5244 13572 5619
rect 13608 5241 13632 5679
rect 13488 5100 13512 5112
rect 13479 5061 13521 5100
rect 13248 4521 13272 5019
rect 13419 4992 13461 5019
rect 13419 4980 13539 4992
rect 13428 4968 13539 4980
rect 13668 4821 13692 5619
rect 13788 5301 13812 5739
rect 13848 5601 13872 6039
rect 14208 5961 14232 7299
rect 14259 7281 14301 7320
rect 14448 7041 14472 7299
rect 14448 6768 14472 6936
rect 14508 6804 14532 7359
rect 14388 6501 14412 6672
rect 14568 6561 14592 6759
rect 13908 5661 13932 5919
rect 13908 5208 13932 5439
rect 13968 5301 13992 5859
rect 12888 4308 12972 4332
rect 12708 3741 12732 4212
rect 12828 4101 12852 4212
rect 13008 3912 13032 4359
rect 13119 4320 13161 4359
rect 13128 4308 13152 4320
rect 13248 4308 13272 4479
rect 13719 4320 13761 4359
rect 13788 4341 13812 5013
rect 13728 4308 13752 4320
rect 13188 4101 13212 4212
rect 13461 4188 13572 4212
rect 13008 3888 13092 3912
rect 12648 2961 12672 3639
rect 12648 2841 12672 2919
rect 12768 2901 12792 3552
rect 12888 3261 12912 3552
rect 13008 3381 13032 3819
rect 13068 3261 13092 3888
rect 13260 3732 13299 3741
rect 13248 3699 13299 3732
rect 13248 3648 13272 3699
rect 12888 3081 12912 3219
rect 13008 2901 13032 3159
rect 12768 2808 12879 2832
rect 12459 2760 12501 2799
rect 12468 2748 12492 2760
rect 12168 2658 12192 2742
rect 12768 2748 12792 2808
rect 12588 2661 12612 2739
rect 13008 2661 13032 2859
rect 12228 2640 12279 2652
rect 12219 2628 12279 2640
rect 12219 2601 12261 2628
rect 11568 2088 11592 2199
rect 10128 1701 10152 1779
rect 9048 1188 9072 1299
rect 9159 1200 9201 1239
rect 9459 1200 9501 1239
rect 9168 1188 9192 1200
rect 9468 1188 9492 1200
rect 9588 1188 9612 1359
rect 9648 1221 9672 1299
rect 8388 1041 8412 1119
rect 9708 1101 9732 1182
rect 8028 438 8052 639
rect 8148 528 8172 879
rect 8268 528 8292 999
rect 7728 420 7752 432
rect 7719 381 7761 420
rect 8328 420 8352 432
rect 8319 381 8361 420
rect 8448 201 8472 819
rect 8508 621 8532 939
rect 8688 861 8712 1092
rect 9228 1080 9252 1092
rect 9408 1080 9432 1092
rect 9219 1041 9261 1080
rect 9399 1041 9441 1080
rect 9528 981 9552 1092
rect 9639 1041 9681 1059
rect 9699 981 9741 996
rect 9768 921 9792 1239
rect 9828 1221 9852 1359
rect 9879 1200 9921 1239
rect 9888 1188 9912 1200
rect 10128 1188 10152 1539
rect 11088 1461 11112 1539
rect 10428 1098 10452 1419
rect 10599 1200 10641 1239
rect 10608 1188 10632 1200
rect 10728 1188 10752 1359
rect 10908 1098 10932 1239
rect 11088 1188 11112 1419
rect 11148 1281 11172 1959
rect 11499 1941 11541 1956
rect 11328 1401 11352 1899
rect 11628 1881 11652 1992
rect 11748 1881 11772 2139
rect 11919 2100 11961 2139
rect 11928 2088 11952 2100
rect 12048 2088 12072 2259
rect 11868 1980 11892 1992
rect 11859 1941 11901 1980
rect 11448 1188 11472 1299
rect 11928 1188 11952 1299
rect 9948 981 9972 1092
rect 10308 981 10332 1092
rect 8781 579 8799 621
rect 8508 438 8532 579
rect 9108 564 9132 879
rect 9741 828 9819 852
rect 8820 552 8859 561
rect 8808 528 8859 552
rect 8820 519 8859 528
rect 9648 528 9672 759
rect 9768 528 9792 759
rect 10068 528 10092 939
rect 10128 561 10152 639
rect 10248 528 10272 699
rect 8928 438 8952 519
rect 9408 438 9432 519
rect 8988 321 9012 399
rect 9468 321 9492 459
rect 10548 441 10572 879
rect 10668 861 10692 1092
rect 10788 1041 10812 1092
rect 10788 1008 10839 1041
rect 10800 999 10839 1008
rect 11061 999 11079 1035
rect 11268 981 11292 1182
rect 9588 261 9612 396
rect 10188 141 10212 399
rect 10368 141 10392 432
rect 10608 381 10632 699
rect 10668 561 10692 639
rect 10728 528 10752 879
rect 10968 561 10992 939
rect 11388 801 11412 1092
rect 11508 1080 11532 1092
rect 11868 1080 11892 1092
rect 11499 1041 11541 1080
rect 11859 1041 11901 1080
rect 11808 648 11832 939
rect 12108 681 12132 1179
rect 12168 981 12192 2439
rect 12228 1998 12252 2199
rect 12288 1821 12312 2319
rect 12408 2241 12432 2652
rect 12708 2640 12732 2652
rect 12699 2601 12741 2640
rect 12768 2181 12792 2259
rect 12768 2088 12792 2139
rect 12348 1581 12372 2019
rect 12660 1992 12699 2001
rect 12468 1761 12492 1992
rect 12648 1968 12699 1992
rect 12660 1959 12699 1968
rect 12468 1341 12492 1719
rect 12888 1224 12912 2139
rect 12948 1998 12972 2319
rect 13068 2181 13092 3219
rect 13128 2781 13152 2919
rect 13221 2832 13260 2841
rect 13221 2799 13272 2832
rect 13248 2748 13272 2799
rect 13308 2772 13332 3399
rect 13428 3381 13452 3699
rect 13488 3681 13512 4119
rect 13539 3660 13581 3699
rect 13548 3648 13572 3660
rect 13368 3192 13392 3339
rect 13368 3168 13452 3192
rect 13308 2748 13392 2772
rect 13368 2421 13392 2748
rect 13428 2241 13452 3168
rect 13488 2781 13512 3039
rect 13608 2832 13632 3516
rect 13548 2808 13632 2832
rect 13548 2748 13572 2808
rect 13668 2748 13692 3159
rect 13788 3141 13812 4179
rect 13848 4101 13872 5079
rect 13968 5001 13992 5112
rect 13908 4218 13932 4419
rect 13968 4341 13992 4719
rect 14028 4392 14052 5079
rect 14088 4461 14112 5319
rect 14148 5301 14172 5772
rect 14208 5208 14232 5739
rect 14268 5301 14292 6159
rect 14508 5868 14532 6399
rect 14628 6081 14652 6819
rect 14688 6801 14712 7332
rect 14868 7221 14892 7428
rect 14748 6768 14772 7119
rect 14928 7101 14952 7488
rect 14988 7461 15012 7659
rect 15048 7512 15072 7728
rect 15168 7521 15192 8199
rect 15228 7821 15252 8256
rect 15288 8241 15312 9408
rect 15348 9081 15372 9279
rect 15468 9261 15492 9876
rect 15588 9561 15612 9792
rect 15708 9681 15732 9792
rect 15501 9228 15552 9252
rect 15441 8799 15459 8841
rect 15348 8361 15372 8739
rect 15408 8328 15432 8559
rect 15468 8421 15492 8679
rect 15528 8541 15552 9228
rect 15828 9081 15852 9639
rect 15588 8661 15612 9039
rect 15828 8988 15852 9039
rect 15948 9024 15972 9519
rect 16128 9492 16152 9639
rect 16188 9561 16212 10239
rect 16128 9468 16212 9492
rect 16008 9021 16032 9459
rect 16068 9072 16092 9399
rect 16188 9141 16212 9468
rect 16248 9261 16272 10299
rect 16368 10281 16392 10452
rect 16308 9921 16332 10179
rect 16368 9888 16392 10119
rect 16488 9984 16512 10359
rect 16548 10221 16572 11199
rect 16608 10641 16632 11439
rect 16668 11448 16752 11472
rect 16788 11448 16812 11559
rect 16908 11448 16932 11619
rect 16968 11541 16992 12012
rect 17028 11481 17052 11559
rect 16668 10821 16692 11448
rect 16728 10761 16752 11319
rect 17088 11352 17112 11979
rect 17148 11601 17172 12879
rect 17259 12861 17301 12900
rect 17379 12861 17421 12900
rect 17448 12888 17532 12912
rect 17208 12141 17232 12819
rect 17388 12381 17412 12819
rect 17448 12801 17472 12888
rect 17568 12852 17592 14439
rect 17628 13521 17652 14859
rect 17688 14481 17712 14799
rect 17688 13701 17712 13959
rect 17748 13881 17772 14979
rect 18048 14781 18072 15132
rect 18228 15021 18252 15222
rect 18288 15081 18312 15339
rect 18348 14592 18372 15999
rect 18408 15561 18432 17079
rect 18321 14568 18372 14592
rect 18228 14412 18252 14499
rect 18168 14388 18252 14412
rect 18168 14301 18192 14388
rect 17988 13761 18012 14139
rect 18288 14001 18312 14559
rect 18408 13761 18432 14679
rect 17988 13668 18132 13692
rect 17688 13461 17712 13539
rect 17748 13101 17772 13536
rect 17868 13281 17892 13572
rect 17808 13008 17832 13119
rect 17928 13041 17952 13539
rect 17988 13401 18012 13668
rect 18288 13461 18312 13572
rect 18048 13008 18072 13239
rect 17628 12861 17652 12999
rect 17748 12900 17772 12912
rect 17508 12828 17592 12852
rect 17268 12261 17292 12339
rect 17259 12120 17301 12156
rect 17388 12144 17412 12276
rect 17268 12108 17292 12120
rect 16839 11301 16881 11316
rect 16968 11241 16992 11352
rect 17028 11328 17112 11352
rect 16599 10581 16641 10599
rect 16659 10560 16701 10599
rect 16668 10548 16692 10560
rect 16788 10548 16812 10959
rect 16608 9921 16632 10419
rect 16068 9060 16152 9072
rect 16068 9048 16161 9060
rect 16119 9021 16161 9048
rect 15528 8328 15552 8436
rect 15648 8361 15672 8799
rect 15048 7488 15132 7512
rect 15108 7428 15132 7488
rect 15288 7461 15312 8136
rect 14988 7041 15012 7299
rect 14808 6321 14832 6672
rect 14328 5208 14352 5499
rect 14508 5241 14532 5679
rect 14628 5481 14652 6039
rect 14928 5961 14952 6819
rect 14988 6792 15012 6999
rect 15048 6861 15072 7332
rect 15168 6801 15192 6999
rect 15228 6981 15252 7179
rect 15288 6981 15312 7299
rect 15348 7161 15372 8139
rect 15588 8121 15612 8232
rect 15708 7881 15732 8619
rect 15948 8601 15972 8982
rect 16188 8988 16212 9099
rect 15768 8361 15792 8439
rect 16008 8361 16032 8859
rect 16248 8721 16272 8859
rect 16068 8421 16092 8619
rect 15408 7461 15432 7839
rect 15768 7812 15792 8199
rect 15828 8172 15852 8232
rect 15828 8148 15939 8172
rect 15708 7788 15792 7812
rect 15528 7428 15552 7539
rect 15339 6981 15381 6999
rect 14988 6768 15072 6792
rect 15228 6672 15252 6819
rect 15288 6741 15312 6939
rect 15408 6792 15432 7299
rect 15648 7152 15672 7659
rect 15588 7128 15672 7152
rect 15348 6768 15432 6792
rect 15468 6768 15492 6939
rect 15588 6768 15612 7128
rect 15708 7092 15732 7788
rect 16008 7701 16032 8199
rect 16068 8121 16092 8316
rect 16128 8181 16152 8259
rect 15768 7281 15792 7599
rect 16128 7461 16152 7659
rect 15948 7320 15972 7332
rect 15648 7068 15732 7092
rect 15648 6861 15672 7068
rect 15768 7041 15792 7119
rect 15708 7008 15759 7032
rect 15168 6648 15252 6672
rect 14688 5472 14712 5919
rect 14688 5448 14772 5472
rect 14559 5220 14601 5259
rect 14568 5208 14592 5220
rect 14268 4581 14292 5112
rect 14508 4701 14532 5079
rect 14028 4368 14112 4392
rect 14088 4308 14112 4368
rect 14199 4320 14241 4359
rect 14208 4308 14232 4320
rect 14028 4041 14052 4176
rect 14148 3921 14172 4212
rect 14328 3690 14352 4299
rect 14388 4221 14412 4359
rect 14688 4308 14712 4479
rect 14748 4401 14772 5448
rect 14808 5112 14832 5679
rect 14868 5241 14892 5739
rect 14928 5481 14952 5772
rect 15048 5481 15072 5919
rect 15108 5472 15132 6519
rect 15168 5721 15192 6648
rect 15348 6321 15372 6768
rect 15399 6621 15441 6639
rect 15228 5901 15252 6159
rect 15528 6021 15552 6672
rect 15279 5880 15321 5919
rect 15288 5868 15312 5880
rect 15528 5712 15552 5772
rect 15528 5688 15612 5712
rect 15108 5448 15192 5472
rect 14928 5361 14952 5439
rect 15168 5241 15192 5448
rect 14808 5088 14892 5112
rect 14808 4341 14832 5019
rect 14868 4581 14892 5088
rect 14928 4941 14952 5112
rect 15108 5100 15132 5112
rect 15099 5061 15141 5100
rect 14748 4101 14772 4212
rect 13908 3321 13932 3552
rect 14388 3441 14412 3999
rect 14448 3681 14472 3879
rect 14481 3552 14520 3561
rect 14808 3552 14832 4179
rect 14868 4161 14892 4476
rect 14481 3528 14532 3552
rect 14481 3519 14520 3528
rect 14721 3528 14832 3552
rect 13728 2361 13752 2616
rect 13848 2481 13872 2979
rect 14028 2901 14052 3339
rect 14088 3261 14112 3339
rect 14148 2748 14172 2859
rect 13908 2661 13932 2742
rect 14268 2661 14292 3219
rect 14328 2541 14352 2919
rect 14508 2748 14532 2979
rect 14448 2541 14472 2652
rect 12999 2112 13041 2139
rect 12999 2100 13092 2112
rect 13008 2088 13092 2100
rect 13128 1581 13152 1992
rect 13368 1881 13392 2079
rect 13548 1980 13572 1992
rect 13428 1761 13452 1959
rect 13539 1941 13581 1980
rect 13728 1641 13752 2199
rect 13908 2088 13932 2499
rect 13848 1881 13872 1992
rect 13968 1980 13992 1992
rect 13959 1941 14001 1980
rect 13788 1701 13812 1779
rect 12288 801 12312 1092
rect 11208 528 11232 639
rect 10788 420 10812 432
rect 10779 381 10821 420
rect 11088 321 11112 459
rect 11508 441 11532 639
rect 11268 141 11292 432
rect 12048 201 12072 459
rect 12108 438 12132 639
rect 12399 561 12441 579
rect 12228 261 12252 396
rect 12348 321 12372 432
rect 12468 321 12492 522
rect 12639 321 12681 339
rect 12888 201 12912 1182
rect 12948 1101 12972 1419
rect 13068 1188 13092 1359
rect 13179 1200 13221 1239
rect 13188 1188 13212 1200
rect 13488 1092 13512 1479
rect 14088 1212 14112 2139
rect 14208 1761 14232 2379
rect 14319 2100 14361 2139
rect 14328 2088 14352 2100
rect 14448 2088 14472 2319
rect 14568 2121 14592 2652
rect 14748 2181 14772 3528
rect 14868 3501 14892 3999
rect 14868 3201 14892 3459
rect 14859 2961 14901 2979
rect 14841 2940 14901 2961
rect 14841 2928 14892 2940
rect 14841 2919 14880 2928
rect 14868 2748 14892 2859
rect 14928 2841 14952 4359
rect 15108 4308 15132 4539
rect 15168 4401 15192 5079
rect 15228 4941 15252 5499
rect 15048 4200 15072 4212
rect 15039 4161 15081 4200
rect 15168 4101 15192 4212
rect 14988 2784 15012 3159
rect 15168 2901 15192 3639
rect 15228 2841 15252 4179
rect 15288 3021 15312 5679
rect 15348 4461 15372 5379
rect 15528 5208 15552 5559
rect 15588 5541 15612 5688
rect 15648 5241 15672 5739
rect 15708 5361 15732 7008
rect 15828 6981 15852 7299
rect 15939 7281 15981 7320
rect 16188 7332 16212 8559
rect 16248 8361 16272 8679
rect 16308 8481 16332 9519
rect 16368 8421 16392 9099
rect 16548 8988 16572 9159
rect 16608 9021 16632 9759
rect 16668 9561 16692 10179
rect 16728 9921 16752 10059
rect 16788 9972 16812 10359
rect 16848 10041 16872 10452
rect 16908 10101 16932 10419
rect 16788 9948 16872 9972
rect 16848 9888 16872 9948
rect 16968 9924 16992 10299
rect 16728 9441 16752 9759
rect 16788 9621 16812 9792
rect 16908 9681 16932 9792
rect 17028 9621 17052 11328
rect 17148 11292 17172 11496
rect 17208 11481 17232 11979
rect 17328 11901 17352 12012
rect 17328 11448 17352 11559
rect 17388 11541 17412 11619
rect 17448 11481 17472 11979
rect 17508 11841 17532 12828
rect 17268 11340 17292 11352
rect 17088 11268 17172 11292
rect 17088 10581 17112 11268
rect 17208 10881 17232 11319
rect 17259 11301 17301 11340
rect 17148 10641 17172 10779
rect 17328 10584 17352 11259
rect 17388 10761 17412 11253
rect 17088 9741 17112 10419
rect 17148 10281 17172 10452
rect 17148 10041 17172 10119
rect 17268 9981 17292 10119
rect 17328 9888 17352 10239
rect 17388 9921 17412 10416
rect 16668 9201 16692 9279
rect 16728 8988 16752 9219
rect 16428 8541 16452 8979
rect 16779 8841 16821 8859
rect 16848 8661 16872 8979
rect 16908 8901 16932 9576
rect 16968 9021 16992 9519
rect 17268 9501 17292 9792
rect 16608 8541 16632 8619
rect 16848 8541 16872 8619
rect 17028 8541 17052 8892
rect 17148 8832 17172 8856
rect 17088 8808 17172 8832
rect 16659 8481 16701 8499
rect 16299 8340 16341 8376
rect 16308 8328 16332 8340
rect 16539 8340 16581 8379
rect 16548 8328 16572 8340
rect 16248 7461 16272 8199
rect 16368 7941 16392 8232
rect 16668 8238 16692 8376
rect 16839 8340 16881 8379
rect 16848 8328 16872 8340
rect 16608 7872 16632 8199
rect 16788 8220 16812 8232
rect 16779 8181 16821 8220
rect 16548 7848 16632 7872
rect 16308 7428 16332 7599
rect 16479 7440 16521 7479
rect 16548 7461 16572 7848
rect 16488 7428 16512 7440
rect 16608 7341 16632 7659
rect 16128 7308 16212 7332
rect 15978 7260 15981 7281
rect 15888 6768 15912 7059
rect 16008 6801 16032 7239
rect 15828 6612 15852 6672
rect 15828 6588 15912 6612
rect 15468 5001 15492 5112
rect 15408 4308 15432 4539
rect 15528 4344 15552 4659
rect 15588 4641 15612 5112
rect 15588 4341 15612 4419
rect 15348 3261 15372 4179
rect 15468 3801 15492 4212
rect 15648 3732 15672 5079
rect 15708 4821 15732 5256
rect 15768 5241 15792 6219
rect 15828 5901 15852 6519
rect 15888 6201 15912 6588
rect 15948 5961 15972 6672
rect 16008 6561 16032 6639
rect 16068 6261 16092 6999
rect 16128 6561 16152 7308
rect 16428 7041 16452 7299
rect 16668 7281 16692 7479
rect 16788 7428 16812 7959
rect 16908 7521 16932 8199
rect 16968 8001 16992 8439
rect 17088 8412 17112 8808
rect 17268 8721 17292 9279
rect 17328 9021 17352 9699
rect 17388 9561 17412 9759
rect 17448 9741 17472 10539
rect 17508 10281 17532 11559
rect 17568 11541 17592 12759
rect 17688 12501 17712 12879
rect 17739 12861 17781 12900
rect 17748 12204 17772 12819
rect 17868 12741 17892 12912
rect 17868 12108 17892 12339
rect 17928 12141 17952 12879
rect 18108 12741 18132 12912
rect 18048 12708 18099 12732
rect 17628 11901 17652 11979
rect 17688 11601 17712 12012
rect 17808 11901 17832 12012
rect 17661 11532 17700 11541
rect 17661 11499 17712 11532
rect 17679 11484 17712 11499
rect 17808 11481 17832 11559
rect 17628 11340 17652 11352
rect 17568 11241 17592 11319
rect 17619 11301 17661 11340
rect 17748 11241 17772 11352
rect 17568 10161 17592 10839
rect 17628 10581 17652 10959
rect 17808 10821 17832 11319
rect 17688 10548 17712 10659
rect 17808 10548 17832 10779
rect 17868 10581 17892 11439
rect 17628 10041 17652 10419
rect 17748 10341 17772 10452
rect 17388 8988 17412 9159
rect 17508 9021 17532 9999
rect 17808 9981 17832 10359
rect 17868 9981 17892 10419
rect 17679 9900 17721 9939
rect 17820 9918 17880 9921
rect 17820 9909 17859 9918
rect 17688 9888 17712 9900
rect 17808 9885 17859 9909
rect 17820 9879 17859 9885
rect 17628 9780 17652 9792
rect 17619 9741 17661 9780
rect 17028 8400 17112 8412
rect 17019 8388 17112 8400
rect 17019 8361 17061 8388
rect 17148 8328 17172 8499
rect 17328 8421 17352 8859
rect 17448 8781 17472 8892
rect 17508 8481 17532 8859
rect 17568 8781 17592 9339
rect 17628 9141 17652 9519
rect 17688 9381 17712 9639
rect 17748 9621 17772 9792
rect 17688 8988 17712 9276
rect 17808 9252 17832 9699
rect 17748 9228 17832 9252
rect 17748 9081 17772 9228
rect 17808 8988 17832 9159
rect 17868 9021 17892 9759
rect 17628 8601 17652 8739
rect 17259 8340 17301 8379
rect 17388 8361 17412 8439
rect 17688 8424 17712 8799
rect 17748 8601 17772 8892
rect 17268 8328 17292 8340
rect 17448 8241 17472 8379
rect 17088 8220 17112 8232
rect 16899 7440 16941 7479
rect 17028 7461 17052 8199
rect 17079 8181 17121 8220
rect 17208 7572 17232 8232
rect 17148 7548 17232 7572
rect 16908 7428 16932 7440
rect 16488 6972 16512 7059
rect 16788 7041 16812 7239
rect 16968 7221 16992 7332
rect 16428 6948 16512 6972
rect 16428 6768 16452 6948
rect 16728 6861 16752 6939
rect 16248 6612 16272 6672
rect 16188 6588 16272 6612
rect 16128 5901 16152 6279
rect 16188 6201 16212 6588
rect 16548 6561 16572 6762
rect 16248 6381 16272 6519
rect 15948 5721 15972 5772
rect 15828 5301 15852 5679
rect 15948 5421 15972 5679
rect 16128 5541 16152 5739
rect 16188 5361 16212 5979
rect 16248 5781 16272 6339
rect 16308 5901 16332 6459
rect 16728 6201 16752 6279
rect 16368 5868 16392 6039
rect 16599 5880 16641 5919
rect 16659 5901 16701 5919
rect 16608 5868 16632 5880
rect 16728 5778 16752 6159
rect 16788 5961 16812 6579
rect 16848 5901 16872 6672
rect 16968 6501 16992 6999
rect 17028 6201 17052 7299
rect 17088 7281 17112 7479
rect 17148 7461 17172 7548
rect 17268 7512 17292 7719
rect 17328 7641 17352 8232
rect 17388 7521 17412 8199
rect 17448 7941 17472 8199
rect 17748 7881 17772 8199
rect 17268 7488 17352 7512
rect 17199 7440 17241 7479
rect 17208 7428 17232 7440
rect 17328 7428 17352 7488
rect 17148 7221 17172 7299
rect 17208 6852 17232 7239
rect 17268 6912 17292 7332
rect 17508 7338 17532 7659
rect 17268 6888 17352 6912
rect 17208 6828 17292 6852
rect 17268 6768 17292 6828
rect 17328 6801 17352 6888
rect 17448 6792 17472 7299
rect 17388 6768 17472 6792
rect 17508 6768 17532 7179
rect 17568 6981 17592 7479
rect 17628 7461 17652 7779
rect 17748 7428 17772 7719
rect 17808 7521 17832 8739
rect 17868 8601 17892 8859
rect 17928 8412 17952 11799
rect 17988 11481 18012 12159
rect 18048 12141 18072 12708
rect 18108 12108 18132 12339
rect 18228 12204 18252 13119
rect 18288 12261 18312 13356
rect 18348 13281 18372 13539
rect 18348 12132 18372 13239
rect 18408 12201 18432 13656
rect 18348 12108 18432 12132
rect 18048 11661 18072 11979
rect 18108 11541 18132 11919
rect 18288 11781 18312 12012
rect 18408 11901 18432 12108
rect 18348 11868 18399 11892
rect 18048 11508 18099 11532
rect 18048 11448 18072 11508
rect 18168 11481 18192 11739
rect 18048 10581 18072 11019
rect 18108 10941 18132 11352
rect 18168 10692 18192 11319
rect 18228 10701 18252 11619
rect 18288 11001 18312 11499
rect 18348 11061 18372 11868
rect 18108 10680 18192 10692
rect 18099 10668 18192 10680
rect 18099 10641 18141 10668
rect 18228 10632 18252 10659
rect 18168 10608 18252 10632
rect 18168 10548 18192 10608
rect 18288 10548 18312 10779
rect 18348 10581 18372 10899
rect 17988 9681 18012 10539
rect 18048 9921 18072 10119
rect 18108 9981 18132 10452
rect 18168 9888 18192 9999
rect 18108 9780 18132 9792
rect 17988 8841 18012 9459
rect 18048 9021 18072 9759
rect 18099 9741 18141 9780
rect 18108 9201 18132 9636
rect 18228 9501 18252 9792
rect 18168 8988 18192 9099
rect 18288 9081 18312 9699
rect 18348 9621 18372 9999
rect 18348 9012 18372 9459
rect 18408 9201 18432 11739
rect 18288 8988 18372 9012
rect 18408 8898 18432 9039
rect 18048 8481 18072 8859
rect 18108 8721 18132 8892
rect 17901 8388 17952 8412
rect 17868 8232 17892 8379
rect 17979 8340 18021 8379
rect 17988 8328 18012 8340
rect 17868 8208 17952 8232
rect 17928 7341 17952 8208
rect 18048 8001 18072 8196
rect 17988 7461 18012 7719
rect 18048 7521 18072 7839
rect 18168 7761 18192 8439
rect 18048 7428 18072 7479
rect 18168 7428 18192 7599
rect 18228 7461 18252 7959
rect 17628 6792 17652 7299
rect 17688 7221 17712 7332
rect 17868 6981 17892 7299
rect 17748 6801 17772 6939
rect 17628 6768 17712 6792
rect 17208 6561 17232 6672
rect 17328 6081 17352 6339
rect 17061 5979 17079 6021
rect 16899 5961 16941 5979
rect 17079 5880 17121 5916
rect 17088 5868 17112 5880
rect 15819 5220 15861 5259
rect 15939 5220 15981 5259
rect 15828 5208 15852 5220
rect 15948 5208 15972 5220
rect 16068 5112 16092 5319
rect 16179 5220 16221 5256
rect 16308 5241 16332 5736
rect 16368 5601 16392 5679
rect 16788 5661 16812 5799
rect 16839 5721 16881 5739
rect 16188 5208 16212 5220
rect 15768 4341 15792 5079
rect 15888 5001 15912 5112
rect 16008 5088 16092 5112
rect 15828 4641 15852 4839
rect 15828 4308 15852 4599
rect 15948 4341 15972 4599
rect 15588 3708 15672 3732
rect 15108 2658 15132 2739
rect 15108 2541 15132 2616
rect 14919 2100 14961 2139
rect 14928 2088 14952 2100
rect 14388 1872 14412 1992
rect 14439 1872 14481 1899
rect 14388 1860 14481 1872
rect 14388 1848 14472 1860
rect 14028 1188 14112 1212
rect 14139 1200 14181 1239
rect 14148 1188 14172 1200
rect 13128 981 13152 1092
rect 13248 1080 13272 1092
rect 13239 1041 13281 1080
rect 13488 1068 13572 1092
rect 13068 528 13092 759
rect 12948 381 12972 519
rect 13239 381 13281 399
rect 13308 321 13332 522
rect 13401 552 13440 561
rect 13401 528 13452 552
rect 13548 528 13572 1068
rect 13668 564 13692 1056
rect 14028 981 14052 1188
rect 14448 1041 14472 1848
rect 14568 1230 14592 1959
rect 14628 1941 14652 2082
rect 14688 1968 14772 1992
rect 14688 1188 14712 1968
rect 13401 519 13440 528
rect 14508 432 14532 639
rect 14568 432 14592 1188
rect 14748 801 14772 1092
rect 14868 681 14892 1992
rect 14928 1461 14952 1839
rect 14988 1761 15012 1992
rect 15048 1188 15072 1659
rect 15108 1281 15132 2079
rect 15168 1941 15192 2796
rect 15288 2781 15312 2859
rect 15408 2841 15432 3519
rect 15468 3261 15492 3552
rect 15378 2799 15381 2820
rect 15339 2760 15381 2799
rect 15348 2748 15372 2760
rect 15468 2748 15492 2919
rect 15588 2901 15612 3708
rect 15708 3672 15732 4299
rect 15768 3732 15792 4179
rect 15888 4101 15912 4212
rect 15768 3708 15852 3732
rect 15648 3648 15732 3672
rect 15828 3648 15852 3708
rect 15648 3501 15672 3648
rect 16008 3681 16032 5088
rect 16068 4341 16092 5019
rect 16128 4572 16152 5079
rect 16128 4548 16212 4572
rect 16128 4308 16152 4479
rect 16188 4401 16212 4548
rect 16248 4521 16272 5112
rect 16308 4641 16332 5079
rect 16368 4461 16392 5559
rect 16428 5112 16452 5619
rect 16848 5361 16872 5616
rect 16908 5541 16932 5772
rect 17139 5661 17181 5679
rect 17208 5601 17232 5862
rect 17268 5781 17292 5919
rect 17328 5892 17352 5976
rect 17388 5961 17412 6768
rect 17448 5952 17472 6639
rect 17568 6321 17592 6672
rect 17448 5928 17532 5952
rect 17328 5868 17412 5892
rect 17508 5868 17532 5928
rect 17559 5901 17601 5919
rect 17361 5679 17379 5721
rect 16908 5421 16932 5499
rect 16488 5241 16512 5319
rect 16779 5160 16821 5202
rect 16788 5148 16812 5160
rect 16428 5088 16512 5112
rect 16428 4881 16452 5019
rect 16488 4401 16512 5088
rect 16608 4941 16632 5112
rect 16728 4278 16752 5019
rect 17022 4821 17046 5019
rect 17088 4941 17112 5499
rect 17448 5481 17472 5772
rect 17628 5721 17652 5859
rect 17568 5481 17592 5619
rect 17688 5481 17712 6768
rect 17928 6768 17952 7059
rect 17988 6861 18012 7299
rect 18048 7092 18072 7179
rect 18108 7161 18132 7332
rect 18048 7068 18132 7092
rect 18048 6801 18072 6939
rect 17748 5901 17772 6639
rect 17808 6201 17832 6672
rect 17868 5868 17892 6039
rect 17988 5868 18012 6672
rect 18048 5892 18072 6639
rect 18108 6081 18132 7068
rect 18168 6981 18192 7179
rect 18048 5868 18132 5892
rect 17748 5541 17772 5739
rect 17928 5661 17952 5772
rect 17901 5508 18012 5532
rect 17148 5061 17172 5259
rect 17928 5241 17952 5439
rect 17988 5181 18012 5508
rect 17901 5172 17940 5181
rect 17901 5148 17952 5172
rect 17901 5139 17940 5148
rect 18108 5172 18132 5868
rect 18168 5232 18192 6819
rect 18228 5778 18252 7299
rect 18288 7221 18312 8799
rect 18168 5208 18252 5232
rect 18108 5148 18192 5172
rect 17148 4581 17172 4719
rect 17688 4551 17739 4572
rect 17688 4548 17772 4551
rect 17688 4368 17712 4548
rect 15768 3540 15792 3552
rect 15888 3540 15912 3552
rect 15759 3501 15801 3540
rect 15879 3501 15921 3540
rect 15228 2241 15252 2736
rect 15288 2421 15312 2619
rect 15408 2532 15432 2652
rect 15648 2658 15672 3099
rect 15828 2832 15852 3399
rect 16068 3381 16092 4179
rect 16308 3792 16332 4212
rect 16428 4101 16452 4236
rect 16308 3768 16392 3792
rect 16248 3648 16272 3759
rect 16368 3681 16392 3768
rect 16128 3561 16152 3639
rect 16428 3561 16452 3819
rect 15888 2901 15912 3339
rect 16308 3021 16332 3516
rect 16368 3141 16392 3519
rect 16488 3141 16512 4179
rect 16608 3921 16632 4119
rect 16668 3861 16692 4059
rect 16728 3981 16752 4236
rect 16788 4161 16812 4359
rect 16539 3684 16581 3699
rect 17028 3624 17052 3939
rect 17088 3681 17112 3879
rect 17148 3672 17172 3939
rect 17568 3921 17592 4236
rect 17808 4101 17832 4419
rect 17868 4041 17892 4539
rect 17928 3981 17952 4959
rect 18048 4344 18072 5052
rect 18108 4401 18132 5019
rect 18168 4461 18192 5148
rect 18228 4581 18252 5208
rect 17988 3681 18012 4059
rect 17148 3648 17232 3672
rect 16548 3540 16599 3552
rect 16539 3528 16599 3540
rect 16539 3501 16581 3528
rect 17148 3492 17172 3582
rect 17208 3501 17232 3648
rect 18048 3621 18072 3999
rect 18168 3681 18192 4179
rect 18228 3621 18252 4359
rect 18288 3912 18312 7059
rect 18348 7032 18372 8739
rect 18408 7821 18432 8559
rect 18408 7101 18432 7599
rect 18348 7008 18432 7032
rect 18348 4221 18372 6939
rect 18288 3888 18372 3912
rect 17961 3612 18000 3621
rect 17961 3588 18012 3612
rect 17961 3579 18000 3588
rect 18288 3552 18312 3819
rect 18228 3528 18312 3552
rect 17088 3468 17172 3492
rect 15828 2808 15912 2832
rect 15888 2784 15912 2808
rect 15741 2772 15780 2781
rect 15741 2748 15792 2772
rect 15741 2739 15780 2748
rect 16008 2781 16032 2859
rect 16068 2661 16092 2799
rect 16188 2748 16212 2979
rect 16320 2772 16359 2781
rect 16308 2748 16359 2772
rect 16320 2739 16359 2748
rect 15588 2532 15612 2619
rect 15408 2508 15612 2532
rect 15279 2100 15321 2139
rect 15288 2088 15312 2100
rect 15408 2088 15432 2199
rect 15708 2088 15732 2379
rect 15828 2361 15852 2616
rect 15828 2241 15852 2319
rect 15948 2124 15972 2652
rect 16359 2601 16401 2619
rect 16428 2124 16452 2679
rect 15168 1188 15192 1299
rect 15348 1212 15372 1956
rect 15468 1521 15492 1992
rect 15648 1881 15672 1992
rect 16128 1980 16152 1992
rect 15768 1821 15792 1956
rect 16119 1941 16161 1980
rect 16248 1521 16272 1992
rect 16368 1761 16392 1992
rect 16488 1701 16512 2979
rect 16548 2421 16572 3339
rect 16659 2760 16701 2799
rect 16668 2748 16692 2760
rect 16788 2748 16812 3279
rect 17088 2952 17112 3468
rect 18228 3492 18252 3528
rect 18108 3468 18252 3492
rect 17148 3021 17172 3399
rect 18036 3321 18060 3399
rect 17568 3021 17592 3219
rect 17088 2940 17172 2952
rect 17088 2928 17181 2940
rect 17088 2844 17112 2928
rect 17139 2901 17181 2928
rect 16728 2241 16752 2652
rect 16848 2640 16872 2652
rect 16839 2601 16881 2640
rect 16788 2268 16899 2292
rect 16668 2088 16692 2199
rect 16788 2088 16812 2268
rect 16968 2232 16992 2799
rect 17208 2640 17232 2652
rect 17199 2601 17241 2640
rect 16908 2208 16992 2232
rect 16848 2121 16872 2199
rect 16728 1821 16752 1992
rect 16908 1512 16932 2208
rect 16968 1821 16992 2139
rect 17148 2088 17172 2259
rect 17259 2100 17301 2139
rect 17268 2088 17292 2100
rect 16848 1488 16932 1512
rect 17028 1512 17052 1959
rect 17088 1641 17112 1992
rect 17028 1488 17112 1512
rect 15348 1188 15432 1212
rect 15228 1080 15252 1092
rect 15219 1041 15261 1080
rect 15408 1041 15432 1188
rect 15468 801 15492 1299
rect 16128 1188 16152 1479
rect 16299 1200 16341 1239
rect 16479 1200 16521 1239
rect 16308 1188 16332 1200
rect 16488 1188 16512 1200
rect 16668 1188 16692 1359
rect 16788 1161 16812 1419
rect 16848 1281 16872 1488
rect 17088 1221 17112 1488
rect 15048 564 15072 759
rect 15588 552 15612 759
rect 15648 681 15672 1092
rect 15588 528 15672 552
rect 16128 564 16152 639
rect 16788 564 16812 1119
rect 17061 1068 17112 1092
rect 15648 432 15672 528
rect 17088 552 17112 1068
rect 17148 921 17172 1659
rect 17208 1401 17232 1992
rect 17328 1980 17352 1992
rect 17319 1941 17361 1980
rect 17319 1572 17361 1599
rect 17268 1560 17361 1572
rect 17268 1548 17352 1560
rect 17268 1188 17292 1548
rect 17328 1272 17352 1479
rect 17388 1461 17412 1959
rect 17448 1281 17472 2979
rect 17568 2748 17592 2859
rect 17541 2112 17580 2121
rect 17541 2088 17592 2112
rect 17541 2079 17580 2088
rect 17628 1761 17652 1992
rect 17748 1281 17772 2379
rect 17808 1641 17832 3219
rect 17988 2784 18012 2979
rect 17988 1980 18012 1992
rect 17979 1941 18021 1980
rect 17328 1248 17412 1272
rect 17388 1188 17412 1248
rect 17448 921 17472 1092
rect 17088 528 17172 552
rect 17328 528 17352 879
rect 17568 438 17592 1239
rect 17628 1098 17652 1239
rect 17808 1188 17832 1299
rect 17868 1032 17892 1092
rect 17868 1008 17952 1032
rect 17868 528 17892 939
rect 17928 861 17952 1008
rect 18048 981 18072 1479
rect 18108 1098 18132 3099
rect 18168 861 18192 3339
rect 18228 1341 18252 3399
rect 13608 201 13632 432
rect 8361 99 8379 141
rect 8541 99 8559 141
rect 14028 -48 14052 432
rect 15168 -48 15192 432
rect 16248 -48 16272 432
rect 16668 -48 16692 432
rect 13968 -72 14052 -48
rect 15108 -72 15192 -48
rect 16188 -72 16272 -48
rect 16608 -72 16692 -48
rect 17028 -72 17052 432
rect 17448 -48 17472 432
rect 17928 420 17952 432
rect 17919 381 17961 420
rect 18228 381 18252 1299
rect 18288 1224 18312 3459
rect 18348 1521 18372 3888
rect 18408 3381 18432 7008
rect 18408 921 18432 3219
rect 17388 -72 17472 -48
<< m3contact >>
rect 9999 18759 10041 18801
rect 11619 18759 11661 18801
rect 14559 18759 14601 18801
rect 10599 18699 10641 18741
rect 11559 18699 11601 18741
rect 879 18639 921 18681
rect 1959 18639 2001 18681
rect 2739 18639 2781 18681
rect 279 18459 321 18501
rect 759 18459 801 18501
rect 519 18342 561 18384
rect 639 18342 681 18384
rect 1539 18519 1581 18561
rect 1179 18459 1221 18501
rect 876 18339 918 18381
rect 939 18342 981 18384
rect 1059 18342 1101 18384
rect 1779 18399 1821 18441
rect 1539 18342 1581 18384
rect 2259 18579 2301 18621
rect 2199 18519 2241 18561
rect 2079 18342 2121 18384
rect 2619 18459 2661 18501
rect 2259 18399 2301 18441
rect 2379 18399 2421 18441
rect 2559 18399 2601 18441
rect 339 17739 381 17781
rect 459 17682 501 17724
rect 699 18216 741 18258
rect 819 18216 861 18258
rect 939 18219 981 18261
rect 1239 18216 1281 18258
rect 1419 18216 1461 18258
rect 1119 17859 1161 17901
rect 1179 17742 1221 17784
rect 639 17679 681 17721
rect 819 17682 861 17724
rect 999 17682 1041 17724
rect 1179 17682 1221 17724
rect 1299 17682 1341 17724
rect 279 17439 321 17481
rect 279 16839 321 16881
rect 219 16782 261 16824
rect 99 16539 141 16581
rect 39 16122 81 16164
rect 39 15699 81 15741
rect 579 17439 621 17481
rect 519 17319 561 17361
rect 459 17139 501 17181
rect 399 16539 441 16581
rect 279 16419 321 16461
rect 399 16419 441 16461
rect 879 17556 921 17598
rect 759 17319 801 17361
rect 999 17499 1041 17541
rect 1239 17556 1281 17598
rect 1179 17499 1221 17541
rect 1119 17439 1161 17481
rect 879 17079 921 17121
rect 639 16959 681 17001
rect 819 16959 861 17001
rect 519 16779 561 16821
rect 699 16782 741 16824
rect 639 16656 681 16698
rect 159 16299 201 16341
rect 579 16359 621 16401
rect 399 16122 441 16164
rect 759 16299 801 16341
rect 639 16179 681 16221
rect 879 16782 921 16824
rect 999 16782 1041 16824
rect 1779 18219 1821 18261
rect 1899 18216 1941 18258
rect 2019 18216 2061 18258
rect 2319 18216 2361 18258
rect 2439 18216 2481 18258
rect 4299 18579 4341 18621
rect 5979 18579 6021 18621
rect 6219 18579 6261 18621
rect 6699 18579 6741 18621
rect 9579 18579 9621 18621
rect 9759 18579 9801 18621
rect 10599 18579 10641 18621
rect 3279 18459 3321 18501
rect 3579 18459 3621 18501
rect 4119 18459 4161 18501
rect 2859 18342 2901 18384
rect 3039 18342 3081 18384
rect 3399 18342 3441 18384
rect 2619 18279 2661 18321
rect 2799 18216 2841 18258
rect 2559 18159 2601 18201
rect 1599 18099 1641 18141
rect 1899 18099 1941 18141
rect 2319 18099 2361 18141
rect 1779 17979 1821 18021
rect 1659 17739 1701 17781
rect 1479 17679 1521 17721
rect 2379 18039 2421 18081
rect 2919 18039 2961 18081
rect 2559 17979 2601 18021
rect 1959 17919 2001 17961
rect 2379 17919 2421 17961
rect 3039 17919 3081 17961
rect 1899 17859 1941 17901
rect 1419 17439 1461 17481
rect 1419 17139 1461 17181
rect 1179 16779 1221 16821
rect 1299 16782 1341 16824
rect 1599 17556 1641 17598
rect 1719 17556 1761 17598
rect 1839 17556 1881 17598
rect 1659 17439 1701 17481
rect 1839 17439 1881 17481
rect 1599 16782 1641 16824
rect 879 16659 921 16701
rect 1059 16656 1101 16698
rect 1179 16659 1221 16701
rect 1839 17139 1881 17181
rect 1719 16899 1761 16941
rect 1419 16599 1461 16641
rect 1599 16599 1641 16641
rect 1059 16419 1101 16461
rect 1179 16419 1221 16461
rect 1359 16419 1401 16461
rect 879 16359 921 16401
rect 879 16239 921 16281
rect 819 16179 861 16221
rect 639 15996 681 16038
rect 819 15996 861 16038
rect 459 15939 501 15981
rect 579 15939 621 15981
rect 279 15819 321 15861
rect 936 15819 978 15861
rect 999 15819 1041 15861
rect 579 15639 621 15681
rect 279 15399 321 15441
rect 159 15222 201 15264
rect 399 15222 441 15264
rect 99 15096 141 15138
rect 459 15096 501 15138
rect 339 15039 381 15081
rect 519 14619 561 14661
rect 1239 16239 1281 16281
rect 1659 16239 1701 16281
rect 1539 16122 1581 16164
rect 3339 18216 3381 18258
rect 3699 18342 3741 18384
rect 3999 18342 4041 18384
rect 4959 18459 5001 18501
rect 5319 18459 5361 18501
rect 5619 18459 5661 18501
rect 4419 18342 4461 18384
rect 4539 18342 4581 18384
rect 4719 18342 4761 18384
rect 5199 18342 5241 18384
rect 5439 18342 5481 18384
rect 3759 18159 3801 18201
rect 3999 18159 4041 18201
rect 3579 17919 3621 17961
rect 2979 17799 3021 17841
rect 3219 17799 3261 17841
rect 2199 17682 2241 17724
rect 2439 17679 2481 17721
rect 2679 17682 2721 17724
rect 2799 17682 2841 17724
rect 2139 17499 2181 17541
rect 2139 17379 2181 17421
rect 2319 17379 2361 17421
rect 1899 16899 1941 16941
rect 2019 16782 2061 16824
rect 2439 17079 2481 17121
rect 2559 16959 2601 17001
rect 2379 16899 2421 16941
rect 2439 16782 2481 16824
rect 2559 16719 2601 16761
rect 1839 16656 1881 16698
rect 2139 16659 2181 16701
rect 2259 16656 2301 16698
rect 2379 16656 2421 16698
rect 2739 17499 2781 17541
rect 2739 16782 2781 16824
rect 2619 16539 2661 16581
rect 2799 16539 2841 16581
rect 1959 16419 2001 16461
rect 3699 17739 3741 17781
rect 3159 17682 3201 17724
rect 3399 17682 3441 17724
rect 3099 17499 3141 17541
rect 3279 17019 3321 17061
rect 3099 16899 3141 16941
rect 3879 17682 3921 17724
rect 4299 18216 4341 18258
rect 4479 18216 4521 18258
rect 4479 18099 4521 18141
rect 4179 18039 4221 18081
rect 4059 17979 4101 18021
rect 4239 17919 4281 17961
rect 4179 17799 4221 17841
rect 4179 17682 4221 17724
rect 3639 17556 3681 17598
rect 3939 17556 3981 17598
rect 4119 17499 4161 17541
rect 3759 17439 3801 17481
rect 4059 17439 4101 17481
rect 3459 17019 3501 17061
rect 3399 16839 3441 16881
rect 3819 17319 3861 17361
rect 3759 16959 3801 17001
rect 3699 16839 3741 16881
rect 3459 16782 3501 16824
rect 3579 16782 3621 16824
rect 3219 16656 3261 16698
rect 3399 16659 3441 16701
rect 2979 16299 3021 16341
rect 2259 16239 2301 16281
rect 2499 16239 2541 16281
rect 2739 16239 2781 16281
rect 1719 16179 1761 16221
rect 1839 16179 1881 16221
rect 2019 16179 2061 16221
rect 2139 16122 2181 16164
rect 2319 16119 2361 16161
rect 2619 16122 2661 16164
rect 1239 15939 1281 15981
rect 1179 15879 1221 15921
rect 1059 15639 1101 15681
rect 999 15399 1041 15441
rect 759 15222 801 15264
rect 879 15222 921 15264
rect 699 15096 741 15138
rect 819 14919 861 14961
rect 699 14619 741 14661
rect 339 14562 381 14604
rect 459 14439 501 14481
rect 399 14379 441 14421
rect 279 14199 321 14241
rect 39 13959 81 14001
rect 219 13779 261 13821
rect 819 14562 861 14604
rect 939 14559 981 14601
rect 519 14379 561 14421
rect 99 13662 141 13704
rect 219 13662 261 13704
rect 339 13662 381 13704
rect 456 13662 498 13704
rect 939 14436 981 14478
rect 1059 15279 1101 15321
rect 1299 15759 1341 15801
rect 1359 15399 1401 15441
rect 1059 15039 1101 15081
rect 1719 15996 1761 16038
rect 1839 15996 1881 16038
rect 1959 15996 2001 16038
rect 2259 15996 2301 16038
rect 2079 15879 2121 15921
rect 1599 15819 1641 15861
rect 1659 15699 1701 15741
rect 1539 15579 1581 15621
rect 2079 15579 2121 15621
rect 2439 15939 2481 15981
rect 2559 15879 2601 15921
rect 2319 15459 2361 15501
rect 1659 15399 1701 15441
rect 1539 15222 1581 15264
rect 2019 15279 2061 15321
rect 2139 15222 2181 15264
rect 2259 15222 2301 15264
rect 1479 14979 1521 15021
rect 1299 14919 1341 14961
rect 1899 14979 1941 15021
rect 1239 14859 1281 14901
rect 1539 14859 1581 14901
rect 1719 14859 1761 14901
rect 1179 14679 1221 14721
rect 1119 14562 1161 14604
rect 1479 14679 1521 14721
rect 1419 14562 1461 14604
rect 1179 14436 1221 14478
rect 1299 14436 1341 14478
rect 759 14319 801 14361
rect 579 14199 621 14241
rect 639 14199 681 14241
rect 279 13359 321 13401
rect 159 13002 201 13044
rect 279 13002 321 13044
rect 519 13659 561 13701
rect 699 13779 741 13821
rect 879 13659 921 13701
rect 639 13536 681 13578
rect 519 13419 561 13461
rect 39 11799 81 11841
rect 39 10839 81 10881
rect 459 12999 501 13041
rect 699 13119 741 13161
rect 999 14319 1041 14361
rect 999 14139 1041 14181
rect 939 13539 981 13581
rect 879 13419 921 13461
rect 759 13059 801 13101
rect 879 13059 921 13101
rect 819 13002 861 13044
rect 936 13002 978 13044
rect 1419 14019 1461 14061
rect 1659 14619 1701 14661
rect 1779 14562 1821 14604
rect 1659 14379 1701 14421
rect 1599 14199 1641 14241
rect 1479 13839 1521 13881
rect 1179 13659 1221 13701
rect 1299 13662 1341 13704
rect 1119 13536 1161 13578
rect 1239 13359 1281 13401
rect 1119 13119 1161 13161
rect 339 12876 381 12918
rect 519 12879 561 12921
rect 639 12876 681 12918
rect 339 12219 381 12261
rect 999 12999 1041 13041
rect 1359 13059 1401 13101
rect 1059 12876 1101 12918
rect 1299 12879 1341 12921
rect 1179 12819 1221 12861
rect 1719 14139 1761 14181
rect 1839 14019 1881 14061
rect 1539 13662 1581 13704
rect 1659 13662 1701 13704
rect 1599 13536 1641 13578
rect 2079 15039 2121 15081
rect 3759 16779 3801 16821
rect 3639 16656 3681 16698
rect 2799 16122 2841 16164
rect 2919 16122 2961 16164
rect 3039 16122 3081 16164
rect 3219 16116 3261 16158
rect 2979 15996 3021 16038
rect 2919 15879 2961 15921
rect 3099 15879 3141 15921
rect 3219 15879 3261 15921
rect 2799 15699 2841 15741
rect 3339 16299 3381 16341
rect 3519 16239 3561 16281
rect 3939 16782 3981 16824
rect 4239 17559 4281 17601
rect 4419 17556 4461 17598
rect 4719 17979 4761 18021
rect 5019 18216 5061 18258
rect 5139 18216 5181 18258
rect 4899 17799 4941 17841
rect 4659 17682 4701 17724
rect 4839 17682 4881 17724
rect 5019 17682 5061 17724
rect 5379 18216 5421 18258
rect 5499 18099 5541 18141
rect 5199 18039 5241 18081
rect 5739 18342 5781 18384
rect 5859 18342 5901 18384
rect 6099 18519 6141 18561
rect 5739 18216 5781 18258
rect 5319 17859 5361 17901
rect 5619 17859 5661 17901
rect 4779 17556 4821 17598
rect 5079 17556 5121 17598
rect 4659 17439 4701 17481
rect 4599 17319 4641 17361
rect 5199 17199 5241 17241
rect 4419 16782 4461 16824
rect 4839 16839 4881 16881
rect 4719 16782 4761 16824
rect 4959 16779 5001 16821
rect 5259 17139 5301 17181
rect 5679 17799 5721 17841
rect 5439 17682 5481 17724
rect 5619 17682 5661 17724
rect 5379 17559 5421 17601
rect 5499 17556 5541 17598
rect 5619 17439 5661 17481
rect 5379 17199 5421 17241
rect 6339 18342 6381 18384
rect 6519 18342 6561 18384
rect 6759 18519 6801 18561
rect 7119 18519 7161 18561
rect 7419 18519 7461 18561
rect 9279 18519 9321 18561
rect 6819 18339 6861 18381
rect 7359 18342 7401 18384
rect 6279 18216 6321 18258
rect 5919 18159 5961 18201
rect 6099 18159 6141 18201
rect 5859 18039 5901 18081
rect 6159 17979 6201 18021
rect 5979 17682 6021 17724
rect 5919 17556 5961 17598
rect 6039 17556 6081 17598
rect 6519 18219 6561 18261
rect 6759 18216 6801 18258
rect 7059 18216 7101 18258
rect 6399 17859 6441 17901
rect 6339 17799 6381 17841
rect 6759 17682 6801 17724
rect 7059 17682 7101 17724
rect 7299 17859 7341 17901
rect 6339 17556 6381 17598
rect 6159 17499 6201 17541
rect 5739 17319 5781 17361
rect 7119 17556 7161 17598
rect 6819 17439 6861 17481
rect 6699 17199 6741 17241
rect 5739 17139 5781 17181
rect 7239 17139 7281 17181
rect 5319 17019 5361 17061
rect 5379 16839 5421 16881
rect 3999 16539 4041 16581
rect 4179 16539 4221 16581
rect 4599 16659 4641 16701
rect 4779 16656 4821 16698
rect 4959 16656 5001 16698
rect 5139 16656 5181 16698
rect 4479 16539 4521 16581
rect 5079 16539 5121 16581
rect 4359 16479 4401 16521
rect 4899 16479 4941 16521
rect 5139 16479 5181 16521
rect 5079 16419 5121 16461
rect 4059 16359 4101 16401
rect 4356 16359 4398 16401
rect 4419 16359 4461 16401
rect 3819 16122 3861 16164
rect 3939 16122 3981 16164
rect 3579 15996 3621 16038
rect 3879 15879 3921 15921
rect 3459 15819 3501 15861
rect 3759 15819 3801 15861
rect 3399 15699 3441 15741
rect 3699 15699 3741 15741
rect 3279 15579 3321 15621
rect 3519 15579 3561 15621
rect 2919 15459 2961 15501
rect 3279 15459 3321 15501
rect 2439 15222 2481 15264
rect 2619 15219 2661 15261
rect 3459 15339 3501 15381
rect 2499 15096 2541 15138
rect 2319 15039 2361 15081
rect 2619 15039 2661 15081
rect 2259 14859 2301 14901
rect 2376 14859 2418 14901
rect 2439 14859 2481 14901
rect 2079 14619 2121 14661
rect 2199 14562 2241 14604
rect 1959 14439 2001 14481
rect 2139 14319 2181 14361
rect 2199 14199 2241 14241
rect 2259 14139 2301 14181
rect 2319 14079 2361 14121
rect 2319 13959 2361 14001
rect 2199 13719 2241 13761
rect 2019 13662 2061 13704
rect 2139 13662 2181 13704
rect 2319 13659 2361 13701
rect 1779 13479 1821 13521
rect 1899 13479 1941 13521
rect 1599 13359 1641 13401
rect 1719 13359 1761 13401
rect 1599 13002 1641 13044
rect 1419 12879 1461 12921
rect 1359 12759 1401 12801
rect 939 12219 981 12261
rect 1179 12219 1221 12261
rect 759 12159 801 12201
rect 459 12102 501 12144
rect 579 12102 621 12144
rect 699 12102 741 12144
rect 159 11979 201 12021
rect 279 11976 321 12018
rect 399 11919 441 11961
rect 339 11739 381 11781
rect 159 11499 201 11541
rect 459 11679 501 11721
rect 999 12099 1041 12141
rect 639 11979 681 12021
rect 579 11439 621 11481
rect 159 11316 201 11358
rect 279 11316 321 11358
rect 519 11199 561 11241
rect 579 10779 621 10821
rect 399 10536 441 10578
rect 759 11919 801 11961
rect 819 11679 861 11721
rect 759 11499 801 11541
rect 999 11739 1041 11781
rect 1659 12819 1701 12861
rect 1539 12759 1581 12801
rect 2079 13536 2121 13578
rect 1839 13179 1881 13221
rect 1959 13179 2001 13221
rect 2739 14919 2781 14961
rect 2979 15039 3021 15081
rect 2859 14859 2901 14901
rect 2559 14562 2601 14604
rect 3279 15222 3321 15264
rect 3219 14919 3261 14961
rect 3039 14799 3081 14841
rect 3039 14619 3081 14661
rect 2439 14439 2481 14481
rect 2619 14436 2661 14478
rect 2919 14436 2961 14478
rect 3039 14436 3081 14478
rect 2619 14319 2661 14361
rect 3159 14139 3201 14181
rect 2619 13899 2661 13941
rect 2919 13839 2961 13881
rect 2439 13659 2481 13701
rect 2379 13539 2421 13581
rect 2199 13059 2241 13101
rect 2019 13002 2061 13044
rect 1839 12819 1881 12861
rect 1779 12699 1821 12741
rect 2079 12879 2121 12921
rect 1959 12579 2001 12621
rect 2679 13479 2721 13521
rect 2439 13419 2481 13461
rect 2559 13419 2601 13461
rect 2319 13359 2361 13401
rect 3099 13779 3141 13821
rect 3279 14562 3321 14604
rect 4179 16119 4221 16161
rect 4659 16119 4701 16161
rect 4899 16122 4941 16164
rect 5499 16782 5541 16824
rect 5619 16782 5661 16824
rect 5799 17079 5841 17121
rect 5979 17019 6021 17061
rect 5859 16839 5901 16881
rect 5799 16782 5841 16824
rect 5559 16656 5601 16698
rect 5739 16659 5781 16701
rect 8319 18459 8361 18501
rect 8559 18459 8601 18501
rect 7719 18342 7761 18384
rect 8199 18342 8241 18384
rect 8319 18342 8361 18384
rect 8439 18342 8481 18384
rect 8859 18342 8901 18384
rect 7359 17679 7401 17721
rect 7539 18216 7581 18258
rect 8139 18216 8181 18258
rect 9099 18339 9141 18381
rect 8139 18099 8181 18141
rect 8259 18099 8301 18141
rect 7659 17799 7701 17841
rect 7899 17799 7941 17841
rect 7599 17682 7641 17724
rect 7719 17682 7761 17724
rect 8019 17682 8061 17724
rect 7419 17556 7461 17598
rect 8139 17679 8181 17721
rect 8499 17799 8541 17841
rect 7839 17556 7881 17598
rect 7959 17556 8001 17598
rect 7539 17439 7581 17481
rect 7299 16959 7341 17001
rect 8079 16959 8121 17001
rect 7779 16899 7821 16941
rect 6699 16839 6741 16881
rect 7179 16839 7221 16881
rect 7479 16839 7521 16881
rect 7659 16839 7701 16881
rect 6159 16782 6201 16824
rect 6399 16782 6441 16824
rect 6519 16782 6561 16824
rect 6639 16782 6681 16824
rect 5859 16599 5901 16641
rect 5679 16479 5721 16521
rect 5799 16479 5841 16521
rect 5856 16359 5898 16401
rect 5919 16359 5961 16401
rect 5259 16239 5301 16281
rect 5379 16239 5421 16281
rect 5259 16122 5301 16164
rect 5499 16122 5541 16164
rect 5619 16122 5661 16164
rect 5739 16122 5781 16164
rect 6459 16656 6501 16698
rect 6339 16599 6381 16641
rect 6039 16299 6081 16341
rect 6039 16122 6081 16164
rect 6159 16122 6201 16164
rect 4419 15759 4461 15801
rect 4719 15759 4761 15801
rect 4479 15699 4521 15741
rect 4179 15519 4221 15561
rect 4119 15459 4161 15501
rect 4359 15459 4401 15501
rect 4059 15339 4101 15381
rect 3879 15279 3921 15321
rect 3999 15279 4041 15321
rect 4419 15279 4461 15321
rect 4239 15222 4281 15264
rect 4359 15222 4401 15264
rect 4059 15096 4101 15138
rect 3639 15039 3681 15081
rect 3759 15039 3801 15081
rect 3879 15039 3921 15081
rect 3999 15039 4041 15081
rect 3519 14919 3561 14961
rect 3339 14559 3381 14601
rect 3399 14562 3441 14604
rect 3579 14559 3621 14601
rect 3459 14436 3501 14478
rect 3279 14259 3321 14301
rect 3579 14079 3621 14121
rect 3819 14799 3861 14841
rect 3939 14739 3981 14781
rect 3939 14559 3981 14601
rect 3759 14319 3801 14361
rect 4419 15039 4461 15081
rect 4359 14799 4401 14841
rect 4059 14562 4101 14604
rect 4239 14562 4281 14604
rect 3999 14379 4041 14421
rect 4359 14379 4401 14421
rect 4179 14319 4221 14361
rect 4059 14199 4101 14241
rect 4059 14136 4101 14178
rect 4179 14139 4221 14181
rect 3879 14079 3921 14121
rect 3639 13959 3681 14001
rect 3879 13959 3921 14001
rect 3459 13899 3501 13941
rect 3219 13779 3261 13821
rect 3099 13659 3141 13701
rect 3399 13719 3441 13761
rect 2919 13239 2961 13281
rect 3099 13539 3141 13581
rect 2619 13179 2661 13221
rect 2859 13179 2901 13221
rect 2979 13179 3021 13221
rect 2559 13119 2601 13161
rect 2379 13059 2421 13101
rect 2319 12819 2361 12861
rect 2139 12699 2181 12741
rect 2259 12699 2301 12741
rect 2319 12579 2361 12621
rect 2079 12399 2121 12441
rect 1479 12219 1521 12261
rect 2259 12219 2301 12261
rect 1479 12102 1521 12144
rect 1599 12102 1641 12144
rect 1719 12102 1761 12144
rect 2019 12102 2061 12144
rect 1419 11859 1461 11901
rect 1659 11976 1701 12018
rect 1539 11919 1581 11961
rect 1239 11799 1281 11841
rect 1479 11799 1521 11841
rect 1119 11619 1161 11661
rect 1539 11619 1581 11661
rect 1239 11499 1281 11541
rect 879 11439 921 11481
rect 1059 11439 1101 11481
rect 759 11316 801 11358
rect 939 11199 981 11241
rect 999 10839 1041 10881
rect 819 10719 861 10761
rect 699 10539 741 10581
rect 159 10413 201 10455
rect 219 10419 261 10461
rect 99 10299 141 10341
rect 279 10413 321 10455
rect 459 10359 501 10401
rect 339 10179 381 10221
rect 99 9879 141 9921
rect 219 9882 261 9924
rect 459 9879 501 9921
rect 279 9756 321 9798
rect 399 9639 441 9681
rect 699 10359 741 10401
rect 579 9939 621 9981
rect 699 9939 741 9981
rect 1779 11499 1821 11541
rect 1899 11499 1941 11541
rect 1719 11442 1761 11484
rect 1179 11316 1221 11358
rect 1119 11259 1161 11301
rect 1059 10719 1101 10761
rect 1539 11316 1581 11358
rect 1659 11316 1701 11358
rect 1839 11319 1881 11361
rect 1779 11139 1821 11181
rect 1299 10839 1341 10881
rect 1299 10542 1341 10584
rect 1479 10542 1521 10584
rect 1599 10599 1641 10641
rect 1839 10599 1881 10641
rect 2139 11919 2181 11961
rect 2019 11859 2061 11901
rect 2079 11799 2121 11841
rect 2019 11739 2061 11781
rect 1959 11439 2001 11481
rect 3279 13536 3321 13578
rect 3159 13419 3201 13461
rect 3639 13719 3681 13761
rect 3759 13662 3801 13704
rect 3939 13662 3981 13704
rect 4179 13899 4221 13941
rect 4599 15579 4641 15621
rect 4599 15279 4641 15321
rect 4959 15699 5001 15741
rect 4839 15459 4881 15501
rect 4839 15222 4881 15264
rect 4959 15222 5001 15264
rect 4779 15096 4821 15138
rect 4719 14979 4761 15021
rect 4659 14679 4701 14721
rect 4779 14919 4821 14961
rect 5379 15939 5421 15981
rect 5319 15759 5361 15801
rect 5259 15339 5301 15381
rect 5259 15222 5301 15264
rect 5019 14979 5061 15021
rect 4959 14739 5001 14781
rect 5199 15096 5241 15138
rect 5319 15099 5361 15141
rect 5259 14979 5301 15021
rect 5199 14859 5241 14901
rect 5139 14799 5181 14841
rect 5079 14679 5121 14721
rect 4779 14559 4821 14601
rect 4959 14562 5001 14604
rect 4599 14436 4641 14478
rect 4899 14319 4941 14361
rect 4659 14259 4701 14301
rect 4779 14259 4821 14301
rect 4479 14019 4521 14061
rect 5139 14439 5181 14481
rect 4839 14019 4881 14061
rect 5019 14019 5061 14061
rect 4779 13899 4821 13941
rect 4539 13662 4581 13704
rect 4659 13662 4701 13704
rect 3516 13536 3558 13578
rect 3579 13536 3621 13578
rect 3699 13536 3741 13578
rect 3459 13359 3501 13401
rect 3699 13419 3741 13461
rect 3519 13299 3561 13341
rect 3336 13239 3378 13281
rect 3399 13239 3441 13281
rect 3279 13059 3321 13101
rect 2439 12876 2481 12918
rect 3039 12876 3081 12918
rect 3159 12876 3201 12918
rect 3279 12876 3321 12918
rect 2799 12819 2841 12861
rect 2379 12519 2421 12561
rect 2739 12519 2781 12561
rect 2679 12399 2721 12441
rect 2319 12039 2361 12081
rect 2439 11799 2481 11841
rect 2259 11679 2301 11721
rect 2199 11439 2241 11481
rect 2619 11799 2661 11841
rect 2559 11739 2601 11781
rect 2499 11619 2541 11661
rect 2439 11499 2481 11541
rect 2019 11316 2061 11358
rect 2139 11316 2181 11358
rect 2259 11316 2301 11358
rect 2019 11139 2061 11181
rect 2079 10959 2121 11001
rect 2019 10659 2061 10701
rect 1899 10542 1941 10584
rect 2019 10539 2061 10581
rect 1059 10416 1101 10458
rect 1299 10419 1341 10461
rect 1119 10059 1161 10101
rect 1539 10416 1581 10458
rect 2019 10419 2061 10461
rect 1779 10299 1821 10341
rect 1959 10359 2001 10401
rect 1239 9999 1281 10041
rect 819 9882 861 9924
rect 1119 9882 1161 9924
rect 1599 10059 1641 10101
rect 1419 9999 1461 10041
rect 1359 9819 1401 9861
rect 579 9639 621 9681
rect 519 9339 561 9381
rect 399 8982 441 9024
rect 519 8982 561 9024
rect 99 8856 141 8898
rect 219 8856 261 8898
rect 339 8856 381 8898
rect 399 8679 441 8721
rect 159 8319 201 8361
rect 279 8322 321 8364
rect 519 8439 561 8481
rect 39 8019 81 8061
rect 459 8196 501 8238
rect 879 9756 921 9798
rect 1059 9756 1101 9798
rect 1179 9756 1221 9798
rect 759 9639 801 9681
rect 939 9459 981 9501
rect 639 8982 681 9024
rect 819 8982 861 9024
rect 1719 9882 1761 9924
rect 2259 10779 2301 10821
rect 2379 11316 2421 11358
rect 2559 11319 2601 11361
rect 2499 11199 2541 11241
rect 2319 10659 2361 10701
rect 2199 10542 2241 10584
rect 2499 10542 2541 10584
rect 1899 10239 1941 10281
rect 2076 10239 2118 10281
rect 2139 10239 2181 10281
rect 1839 9999 1881 10041
rect 1659 9756 1701 9798
rect 1839 9756 1881 9798
rect 2379 10416 2421 10458
rect 2499 10419 2541 10461
rect 2679 11559 2721 11601
rect 3219 12699 3261 12741
rect 3939 13539 3981 13581
rect 4119 13536 4161 13578
rect 4419 13539 4461 13581
rect 3936 13299 3978 13341
rect 3999 13299 4041 13341
rect 3459 13059 3501 13101
rect 3579 13059 3621 13101
rect 3519 13002 3561 13044
rect 3459 12759 3501 12801
rect 3399 12639 3441 12681
rect 3339 12519 3381 12561
rect 3279 12399 3321 12441
rect 3219 12279 3261 12321
rect 2859 12036 2901 12078
rect 3039 11919 3081 11961
rect 2979 11799 3021 11841
rect 2739 11439 2781 11481
rect 2859 11442 2901 11484
rect 3639 12879 3681 12921
rect 3579 12579 3621 12621
rect 3999 13059 4041 13101
rect 4419 13419 4461 13461
rect 4359 13359 4401 13401
rect 4599 13536 4641 13578
rect 4239 13299 4281 13341
rect 4479 13119 4521 13161
rect 4719 13119 4761 13161
rect 3819 12939 3861 12981
rect 4176 12939 4218 12981
rect 4239 12939 4281 12981
rect 3699 12699 3741 12741
rect 3939 12819 3981 12861
rect 3879 12579 3921 12621
rect 3639 12399 3681 12441
rect 3759 12279 3801 12321
rect 3579 12102 3621 12144
rect 3099 11679 3141 11721
rect 3339 11679 3381 11721
rect 2679 11316 2721 11358
rect 2799 11316 2841 11358
rect 2679 11139 2721 11181
rect 2619 10959 2661 11001
rect 2559 10359 2601 10401
rect 3579 11799 3621 11841
rect 3519 11679 3561 11721
rect 3459 11559 3501 11601
rect 3279 11442 3321 11484
rect 3399 11442 3441 11484
rect 3159 11319 3201 11361
rect 3339 11259 3381 11301
rect 3519 11259 3561 11301
rect 3099 11139 3141 11181
rect 2979 11019 3021 11061
rect 2859 10779 2901 10821
rect 2859 10659 2901 10701
rect 2739 10542 2781 10584
rect 3219 10779 3261 10821
rect 3039 10659 3081 10701
rect 2979 10539 3021 10581
rect 2679 10419 2721 10461
rect 2619 10299 2661 10341
rect 2799 10416 2841 10458
rect 2919 10359 2961 10401
rect 2739 10299 2781 10341
rect 2679 10239 2721 10281
rect 2259 10179 2301 10221
rect 2559 10179 2601 10221
rect 2259 10059 2301 10101
rect 2139 9999 2181 10041
rect 2139 9882 2181 9924
rect 2319 9882 2361 9924
rect 2439 9882 2481 9924
rect 1779 9639 1821 9681
rect 1419 9519 1461 9561
rect 1299 9459 1341 9501
rect 1179 9339 1221 9381
rect 1059 9039 1101 9081
rect 879 8856 921 8898
rect 819 8679 861 8721
rect 639 8559 681 8601
rect 759 8559 801 8601
rect 999 8439 1041 8481
rect 639 8319 681 8361
rect 879 8322 921 8364
rect 339 8139 381 8181
rect 459 8019 501 8061
rect 159 7779 201 7821
rect 39 7719 81 7761
rect 99 7539 141 7581
rect 219 7422 261 7464
rect 399 7422 441 7464
rect 159 7239 201 7281
rect 99 7119 141 7161
rect 99 6759 141 6801
rect 99 6279 141 6321
rect 99 5559 141 5601
rect 339 7299 381 7341
rect 279 7119 321 7161
rect 699 8196 741 8238
rect 639 7899 681 7941
rect 939 8139 981 8181
rect 879 8019 921 8061
rect 819 7659 861 7701
rect 759 7599 801 7641
rect 639 7539 681 7581
rect 759 7422 801 7464
rect 516 7239 558 7281
rect 579 7239 621 7281
rect 219 6999 261 7041
rect 339 6999 381 7041
rect 579 6999 621 7041
rect 339 6879 381 6921
rect 459 6762 501 6804
rect 279 6636 321 6678
rect 219 6579 261 6621
rect 219 6219 261 6261
rect 759 7119 801 7161
rect 879 7119 921 7161
rect 879 6999 921 7041
rect 759 6879 801 6921
rect 819 6819 861 6861
rect 699 6762 741 6804
rect 1479 9159 1521 9201
rect 1779 9039 1821 9081
rect 1539 8982 1581 9024
rect 1659 8982 1701 9024
rect 1239 8856 1281 8898
rect 1359 8856 1401 8898
rect 1479 8859 1521 8901
rect 1179 8619 1221 8661
rect 1899 8979 1941 9021
rect 1719 8856 1761 8898
rect 1899 8799 1941 8841
rect 1839 8739 1881 8781
rect 1719 8679 1761 8721
rect 1539 8559 1581 8601
rect 1659 8499 1701 8541
rect 1479 8439 1521 8481
rect 1299 8322 1341 8364
rect 1659 8322 1701 8364
rect 1779 8322 1821 8364
rect 1239 8196 1281 8238
rect 1479 8196 1521 8238
rect 1059 8139 1101 8181
rect 1719 8196 1761 8238
rect 1539 8079 1581 8121
rect 999 8019 1041 8061
rect 1539 7779 1581 7821
rect 2079 9756 2121 9798
rect 2139 9699 2181 9741
rect 2139 9519 2181 9561
rect 2679 9879 2721 9921
rect 2619 9756 2661 9798
rect 2499 9699 2541 9741
rect 3459 11139 3501 11181
rect 3339 10659 3381 10701
rect 3099 10359 3141 10401
rect 3279 10299 3321 10341
rect 3519 10779 3561 10821
rect 3039 10179 3081 10221
rect 3459 10179 3501 10221
rect 2979 10059 3021 10101
rect 3099 10059 3141 10101
rect 3339 10059 3381 10101
rect 3459 10059 3501 10101
rect 3339 9939 3381 9981
rect 3459 9939 3501 9981
rect 3819 12102 3861 12144
rect 3759 11859 3801 11901
rect 3699 11799 3741 11841
rect 3999 12519 4041 12561
rect 4659 12819 4701 12861
rect 4419 12699 4461 12741
rect 4119 12279 4161 12321
rect 4299 12279 4341 12321
rect 3999 12159 4041 12201
rect 4299 12159 4341 12201
rect 4239 12099 4281 12141
rect 3879 11979 3921 12021
rect 3819 11679 3861 11721
rect 3819 11559 3861 11601
rect 3939 11442 3981 11484
rect 4179 11859 4221 11901
rect 4239 11799 4281 11841
rect 5199 13959 5241 14001
rect 5139 13839 5181 13881
rect 5019 13662 5061 13704
rect 5139 13662 5181 13704
rect 5199 13479 5241 13521
rect 5079 13419 5121 13461
rect 4959 13239 5001 13281
rect 5019 13179 5061 13221
rect 4899 12879 4941 12921
rect 4776 12639 4818 12681
rect 4839 12639 4881 12681
rect 4779 12576 4821 12618
rect 4719 12519 4761 12561
rect 4599 12459 4641 12501
rect 4419 12102 4461 12144
rect 4479 11976 4521 12018
rect 4659 11979 4701 12021
rect 4359 11859 4401 11901
rect 4299 11619 4341 11661
rect 4599 11619 4641 11661
rect 4539 11559 4581 11601
rect 4479 11436 4521 11478
rect 4059 11376 4101 11418
rect 3639 11316 3681 11358
rect 3759 11316 3801 11358
rect 3879 11316 3921 11358
rect 3999 11319 4041 11361
rect 3759 10899 3801 10941
rect 3699 10779 3741 10821
rect 4059 11199 4101 11241
rect 4299 11316 4341 11358
rect 4179 11199 4221 11241
rect 4119 10719 4161 10761
rect 3579 10659 3621 10701
rect 3759 10659 3801 10701
rect 3879 10659 3921 10701
rect 3999 10659 4041 10701
rect 3759 10542 3801 10584
rect 4179 10542 4221 10584
rect 4299 10542 4341 10584
rect 4539 11316 4581 11358
rect 5019 12759 5061 12801
rect 4959 12339 5001 12381
rect 4899 12102 4941 12144
rect 5139 12879 5181 12921
rect 5079 12699 5121 12741
rect 5619 15939 5661 15981
rect 5439 15879 5481 15921
rect 5799 15879 5841 15921
rect 6219 15879 6261 15921
rect 6039 15759 6081 15801
rect 6159 15759 6201 15801
rect 5736 15699 5778 15741
rect 5799 15699 5841 15741
rect 6039 15639 6081 15681
rect 5619 15579 5661 15621
rect 5739 15579 5781 15621
rect 5436 15219 5478 15261
rect 5499 15222 5541 15264
rect 5739 15222 5781 15264
rect 5859 15222 5901 15264
rect 5679 15099 5721 15141
rect 5379 15039 5421 15081
rect 5559 15039 5601 15081
rect 5319 14919 5361 14961
rect 5439 14679 5481 14721
rect 5439 14562 5481 14604
rect 5559 14436 5601 14478
rect 5619 14319 5661 14361
rect 6459 16539 6501 16581
rect 6399 16479 6441 16521
rect 6339 15759 6381 15801
rect 6219 15639 6261 15681
rect 6999 16782 7041 16824
rect 6759 16659 6801 16701
rect 6939 16599 6981 16641
rect 7359 16782 7401 16824
rect 7599 16782 7641 16824
rect 7179 16599 7221 16641
rect 6699 16539 6741 16581
rect 6819 16539 6861 16581
rect 6939 16536 6981 16578
rect 7059 16539 7101 16581
rect 6579 16479 6621 16521
rect 6759 16479 6801 16521
rect 6639 16299 6681 16341
rect 7179 16479 7221 16521
rect 6939 16359 6981 16401
rect 6819 16239 6861 16281
rect 7299 16419 7341 16461
rect 7059 16239 7101 16281
rect 6819 16119 6861 16161
rect 6939 16122 6981 16164
rect 7599 16179 7641 16221
rect 7479 16122 7521 16164
rect 7959 16782 8001 16824
rect 8019 16659 8061 16701
rect 7839 16479 7881 16521
rect 7959 16359 8001 16401
rect 7779 16239 7821 16281
rect 6459 15879 6501 15921
rect 6879 15999 6921 16041
rect 6819 15819 6861 15861
rect 6699 15759 6741 15801
rect 6579 15699 6621 15741
rect 6459 15579 6501 15621
rect 6219 15519 6261 15561
rect 6399 15519 6441 15561
rect 5739 15039 5781 15081
rect 5859 15039 5901 15081
rect 6159 15099 6201 15141
rect 6099 14979 6141 15021
rect 5919 14919 5961 14961
rect 5739 14436 5781 14478
rect 5379 14139 5421 14181
rect 5439 14079 5481 14121
rect 5499 13662 5541 13704
rect 5919 14436 5961 14478
rect 5799 14379 5841 14421
rect 5979 14319 6021 14361
rect 5979 14199 6021 14241
rect 5799 14019 5841 14061
rect 5676 13839 5718 13881
rect 5739 13839 5781 13881
rect 5619 13659 5661 13701
rect 5859 13662 5901 13704
rect 5319 13539 5361 13581
rect 5439 13536 5481 13578
rect 5679 13539 5721 13581
rect 5679 13476 5721 13518
rect 5259 13419 5301 13461
rect 5559 13419 5601 13461
rect 5559 13239 5601 13281
rect 5439 13119 5481 13161
rect 5319 13002 5361 13044
rect 5619 13179 5661 13221
rect 5619 12999 5661 13041
rect 5199 12759 5241 12801
rect 5199 12696 5241 12738
rect 4719 11859 4761 11901
rect 4839 11859 4881 11901
rect 4779 11799 4821 11841
rect 4779 11679 4821 11721
rect 4659 11439 4701 11481
rect 4899 11679 4941 11721
rect 4899 11559 4941 11601
rect 4899 11439 4941 11481
rect 4599 11199 4641 11241
rect 4599 11019 4641 11061
rect 4719 11316 4761 11358
rect 4839 11079 4881 11121
rect 4659 10779 4701 10821
rect 4839 10779 4881 10821
rect 4659 10716 4701 10758
rect 4719 10659 4761 10701
rect 3819 10299 3861 10341
rect 4359 10419 4401 10461
rect 4239 10299 4281 10341
rect 4359 10299 4401 10341
rect 4119 10179 4161 10221
rect 3699 10059 3741 10101
rect 3519 9879 3561 9921
rect 2919 9756 2961 9798
rect 2499 9579 2541 9621
rect 2739 9579 2781 9621
rect 2319 9459 2361 9501
rect 2379 9219 2421 9261
rect 2259 9159 2301 9201
rect 2139 9039 2181 9081
rect 2019 8979 2061 9021
rect 2376 8979 2418 9021
rect 2439 8982 2481 9024
rect 2019 8739 2061 8781
rect 2439 8799 2481 8841
rect 2439 8619 2481 8661
rect 2199 8499 2241 8541
rect 2319 8379 2361 8421
rect 2019 8319 2061 8361
rect 2199 8322 2241 8364
rect 2019 7959 2061 8001
rect 1959 7839 2001 7881
rect 2259 8196 2301 8238
rect 3399 9756 3441 9798
rect 3639 9759 3681 9801
rect 3759 9999 3801 10041
rect 3879 9882 3921 9924
rect 4059 9879 4101 9921
rect 3159 9639 3201 9681
rect 3579 9639 3621 9681
rect 2859 9339 2901 9381
rect 3039 9339 3081 9381
rect 2739 9099 2781 9141
rect 2619 8982 2661 9024
rect 3039 9219 3081 9261
rect 2859 8979 2901 9021
rect 3279 9039 3321 9081
rect 3399 8982 3441 9024
rect 3519 8982 3561 9024
rect 3939 9756 3981 9798
rect 3879 9699 3921 9741
rect 3759 9579 3801 9621
rect 2559 8799 2601 8841
rect 2799 8856 2841 8898
rect 2679 8619 2721 8661
rect 2559 8379 2601 8421
rect 2499 8319 2541 8361
rect 3099 8856 3141 8898
rect 3279 8859 3321 8901
rect 3279 8796 3321 8838
rect 3219 8739 3261 8781
rect 3159 8499 3201 8541
rect 2919 8439 2961 8481
rect 2859 8319 2901 8361
rect 2979 8322 3021 8364
rect 2499 8199 2541 8241
rect 2199 7839 2241 7881
rect 2439 7839 2481 7881
rect 2139 7719 2181 7761
rect 1419 7659 1461 7701
rect 1899 7659 1941 7701
rect 1179 7539 1221 7581
rect 1059 7422 1101 7464
rect 1359 7419 1401 7461
rect 1239 7239 1281 7281
rect 1059 6999 1101 7041
rect 1179 6999 1221 7041
rect 1119 6879 1161 6921
rect 939 6819 981 6861
rect 1059 6819 1101 6861
rect 399 6339 441 6381
rect 279 6039 321 6081
rect 339 5862 381 5904
rect 699 6636 741 6678
rect 699 6519 741 6561
rect 639 6399 681 6441
rect 939 6636 981 6678
rect 879 6579 921 6621
rect 579 6339 621 6381
rect 819 6339 861 6381
rect 519 5859 561 5901
rect 339 5679 381 5721
rect 279 5559 321 5601
rect 519 5739 561 5781
rect 399 5559 441 5601
rect 339 5499 381 5541
rect 159 5379 201 5421
rect 159 5199 201 5241
rect 339 5202 381 5244
rect 459 5202 501 5244
rect 999 6519 1041 6561
rect 879 6159 921 6201
rect 879 6039 921 6081
rect 759 5862 801 5904
rect 879 5862 921 5904
rect 639 5739 681 5781
rect 579 5679 621 5721
rect 99 3516 141 3558
rect 99 3279 141 3321
rect 99 3039 141 3081
rect 939 5739 981 5781
rect 819 5499 861 5541
rect 699 5379 741 5421
rect 759 5319 801 5361
rect 639 5199 681 5241
rect 2139 7656 2181 7698
rect 1539 7422 1581 7464
rect 1899 7422 1941 7464
rect 2019 7422 2061 7464
rect 1719 7359 1761 7401
rect 1419 7119 1461 7161
rect 1359 6819 1401 6861
rect 1179 6759 1221 6801
rect 1299 6762 1341 6804
rect 1599 7119 1641 7161
rect 2079 7299 2121 7341
rect 2019 7239 2061 7281
rect 1839 7119 1881 7161
rect 1719 6999 1761 7041
rect 1539 6819 1581 6861
rect 2019 6819 2061 6861
rect 1839 6762 1881 6804
rect 1959 6759 2001 6801
rect 1119 6636 1161 6678
rect 1239 6636 1281 6678
rect 1299 6579 1341 6621
rect 1179 5919 1221 5961
rect 1059 5859 1101 5901
rect 1539 6636 1581 6678
rect 1359 6459 1401 6501
rect 1659 6636 1701 6678
rect 1779 6519 1821 6561
rect 1779 6339 1821 6381
rect 1779 6159 1821 6201
rect 1599 6039 1641 6081
rect 1479 5919 1521 5961
rect 1299 5862 1341 5904
rect 1599 5862 1641 5904
rect 1059 5739 1101 5781
rect 1839 6039 1881 6081
rect 999 5559 1041 5601
rect 939 5259 981 5301
rect 879 5202 921 5244
rect 399 5076 441 5118
rect 579 5076 621 5118
rect 819 5076 861 5118
rect 279 4719 321 4761
rect 459 4659 501 4701
rect 999 4659 1041 4701
rect 339 4539 381 4581
rect 639 4539 681 4581
rect 759 4479 801 4521
rect 939 4479 981 4521
rect 699 4176 741 4218
rect 399 4059 441 4101
rect 339 3939 381 3981
rect 279 3699 321 3741
rect 999 4176 1041 4218
rect 939 4059 981 4101
rect 939 3996 981 4038
rect 579 3759 621 3801
rect 819 3759 861 3801
rect 459 3642 501 3684
rect 759 3642 801 3684
rect 159 2979 201 3021
rect 279 3516 321 3558
rect 399 3516 441 3558
rect 579 3516 621 3558
rect 699 3516 741 3558
rect 1239 5736 1281 5778
rect 1539 5736 1581 5778
rect 1119 5679 1161 5721
rect 1779 5736 1821 5778
rect 1659 5619 1701 5661
rect 1299 5499 1341 5541
rect 1479 5259 1521 5301
rect 1659 5259 1701 5301
rect 1119 5079 1161 5121
rect 1719 5202 1761 5244
rect 1239 5076 1281 5118
rect 1359 5076 1401 5118
rect 1479 5076 1521 5118
rect 1119 4899 1161 4941
rect 1179 4779 1221 4821
rect 1299 5019 1341 5061
rect 1239 4719 1281 4761
rect 1419 4659 1461 4701
rect 1299 4539 1341 4581
rect 1299 4302 1341 4344
rect 1059 3939 1101 3981
rect 1779 5079 1821 5121
rect 1779 4779 1821 4821
rect 1659 4359 1701 4401
rect 1539 4302 1581 4344
rect 2139 7239 2181 7281
rect 2139 7119 2181 7161
rect 2079 6759 2121 6801
rect 3039 8196 3081 8238
rect 2919 8139 2961 8181
rect 2739 8079 2781 8121
rect 2979 8019 3021 8061
rect 2619 7779 2661 7821
rect 2499 7659 2541 7701
rect 2259 7539 2301 7581
rect 2439 7539 2481 7581
rect 2259 7179 2301 7221
rect 2199 7059 2241 7101
rect 2379 7059 2421 7101
rect 2559 7179 2601 7221
rect 2499 6879 2541 6921
rect 2259 6819 2301 6861
rect 2499 6816 2541 6858
rect 2079 6639 2121 6681
rect 2319 6636 2361 6678
rect 2079 6519 2121 6561
rect 2199 6519 2241 6561
rect 2919 7659 2961 7701
rect 2679 7599 2721 7641
rect 2799 7539 2841 7581
rect 3099 7599 3141 7641
rect 3039 7422 3081 7464
rect 3579 8856 3621 8898
rect 3399 8619 3441 8661
rect 3459 8619 3501 8661
rect 3279 8319 3321 8361
rect 3519 8379 3561 8421
rect 3339 8196 3381 8238
rect 3219 8019 3261 8061
rect 3459 8019 3501 8061
rect 3339 7599 3381 7641
rect 3519 7599 3561 7641
rect 3399 7539 3441 7581
rect 2679 7179 2721 7221
rect 3159 7422 3201 7464
rect 3099 7299 3141 7341
rect 3039 7239 3081 7281
rect 2739 6999 2781 7041
rect 2859 6999 2901 7041
rect 2619 6819 2661 6861
rect 2859 6936 2901 6978
rect 2559 6519 2601 6561
rect 2319 6399 2361 6441
rect 2079 6039 2121 6081
rect 2319 6039 2361 6081
rect 1896 5859 1938 5901
rect 1959 5862 2001 5904
rect 2379 5979 2421 6021
rect 2679 6636 2721 6678
rect 2799 6639 2841 6681
rect 2679 6099 2721 6141
rect 2319 5919 2361 5961
rect 2259 5859 2301 5901
rect 1899 5739 1941 5781
rect 2019 5736 2061 5778
rect 2139 5499 2181 5541
rect 2139 5379 2181 5421
rect 1899 5199 1941 5241
rect 2019 5202 2061 5244
rect 2439 5862 2481 5904
rect 2559 5862 2601 5904
rect 2739 5979 2781 6021
rect 2679 5859 2721 5901
rect 2379 5739 2421 5781
rect 2319 5619 2361 5661
rect 2619 5736 2661 5778
rect 2739 5739 2781 5781
rect 2559 5679 2601 5721
rect 2499 5619 2541 5661
rect 2559 5439 2601 5481
rect 2379 5259 2421 5301
rect 2619 5259 2661 5301
rect 2259 5202 2301 5244
rect 2439 5202 2481 5244
rect 1959 5076 2001 5118
rect 2199 5076 2241 5118
rect 2259 5019 2301 5061
rect 2379 5019 2421 5061
rect 2079 4899 2121 4941
rect 2139 4419 2181 4461
rect 1959 4359 2001 4401
rect 1899 4302 1941 4344
rect 2079 4359 2121 4401
rect 1419 3999 1461 4041
rect 1479 3879 1521 3921
rect 999 3639 1041 3681
rect 1119 3642 1161 3684
rect 1239 3642 1281 3684
rect 1599 3819 1641 3861
rect 1659 3699 1701 3741
rect 279 3159 321 3201
rect 459 2979 501 3021
rect 219 2799 261 2841
rect 939 2979 981 3021
rect 759 2859 801 2901
rect 639 2799 681 2841
rect 579 2739 621 2781
rect 159 2559 201 2601
rect 159 2259 201 2301
rect 99 2139 141 2181
rect 519 2619 561 2661
rect 399 2559 441 2601
rect 339 2199 381 2241
rect 279 2139 321 2181
rect 699 2616 741 2658
rect 939 2616 981 2658
rect 819 2319 861 2361
rect 579 2199 621 2241
rect 519 2082 561 2124
rect 159 1956 201 1998
rect 279 1956 321 1998
rect 99 1839 141 1881
rect 399 1839 441 1881
rect 339 1419 381 1461
rect 459 1239 501 1281
rect 1179 3399 1221 3441
rect 1419 3519 1461 3561
rect 1299 3219 1341 3261
rect 1179 3159 1221 3201
rect 1239 3039 1281 3081
rect 1179 2799 1221 2841
rect 1119 2742 1161 2784
rect 1059 2619 1101 2661
rect 1539 3516 1581 3558
rect 1899 3759 1941 3801
rect 2079 4119 2121 4161
rect 2019 4059 2061 4101
rect 2139 4059 2181 4101
rect 2019 3996 2061 4038
rect 1959 3699 2001 3741
rect 2619 5076 2661 5118
rect 2499 4659 2541 4701
rect 2439 4419 2481 4461
rect 2619 4359 2661 4401
rect 2499 4176 2541 4218
rect 2619 4176 2661 4218
rect 2739 5379 2781 5421
rect 3159 7239 3201 7281
rect 3099 6939 3141 6981
rect 3579 7479 3621 7521
rect 3699 8619 3741 8661
rect 4059 9459 4101 9501
rect 3939 8982 3981 9024
rect 3879 8739 3921 8781
rect 4119 9159 4161 9201
rect 4119 8859 4161 8901
rect 3999 8619 4041 8661
rect 3759 8499 3801 8541
rect 3999 8439 4041 8481
rect 3879 8322 3921 8364
rect 3819 7839 3861 7881
rect 3939 7779 3981 7821
rect 4719 10542 4761 10584
rect 4419 10179 4461 10221
rect 4299 9882 4341 9924
rect 4419 9882 4461 9924
rect 4659 10416 4701 10458
rect 5139 12279 5181 12321
rect 5079 11679 5121 11721
rect 5079 11559 5121 11601
rect 5019 11439 5061 11481
rect 5499 12876 5541 12918
rect 5739 13419 5781 13461
rect 5679 12699 5721 12741
rect 5379 12219 5421 12261
rect 5919 13239 5961 13281
rect 6339 15339 6381 15381
rect 6579 15519 6621 15561
rect 6459 15222 6501 15264
rect 6939 15939 6981 15981
rect 6879 15699 6921 15741
rect 6579 14979 6621 15021
rect 6879 15099 6921 15141
rect 6399 14919 6441 14961
rect 6759 14919 6801 14961
rect 6879 14859 6921 14901
rect 6219 14679 6261 14721
rect 6459 14679 6501 14721
rect 6219 14436 6261 14478
rect 6339 14319 6381 14361
rect 6399 14259 6441 14301
rect 6339 14139 6381 14181
rect 6279 14079 6321 14121
rect 6159 13662 6201 13704
rect 7239 15999 7281 16041
rect 7359 15999 7401 16041
rect 6999 15879 7041 15921
rect 7299 15879 7341 15921
rect 6999 15699 7041 15741
rect 7059 15279 7101 15321
rect 7179 15279 7221 15321
rect 6999 15159 7041 15201
rect 7419 15819 7461 15861
rect 7719 15879 7761 15921
rect 7656 15759 7698 15801
rect 7719 15759 7761 15801
rect 7539 15459 7581 15501
rect 7839 16179 7881 16221
rect 8019 16179 8061 16221
rect 8319 17556 8361 17598
rect 9099 18216 9141 18258
rect 9219 18216 9261 18258
rect 8979 18099 9021 18141
rect 8919 17739 8961 17781
rect 9639 18216 9681 18258
rect 9099 17682 9141 17724
rect 8979 17619 9021 17661
rect 8619 17556 8661 17598
rect 8199 17379 8241 17421
rect 8559 17379 8601 17421
rect 8499 17139 8541 17181
rect 8259 16899 8301 16941
rect 8199 16779 8241 16821
rect 8379 16782 8421 16824
rect 8319 16656 8361 16698
rect 8379 16599 8421 16641
rect 8139 16239 8181 16281
rect 8139 16122 8181 16164
rect 8259 16122 8301 16164
rect 8559 17079 8601 17121
rect 8739 17439 8781 17481
rect 9459 17739 9501 17781
rect 9579 17682 9621 17724
rect 9399 17556 9441 17598
rect 9519 17556 9561 17598
rect 9159 17259 9201 17301
rect 9279 17259 9321 17301
rect 8739 17079 8781 17121
rect 9039 17079 9081 17121
rect 8859 16782 8901 16824
rect 8979 16782 9021 16824
rect 8619 16599 8661 16641
rect 8859 16599 8901 16641
rect 8799 16479 8841 16521
rect 8619 16359 8661 16401
rect 8559 16299 8601 16341
rect 7899 15996 7941 16038
rect 8019 15996 8061 16038
rect 7959 15879 8001 15921
rect 7839 15759 7881 15801
rect 7839 15579 7881 15621
rect 7779 15519 7821 15561
rect 7539 15339 7581 15381
rect 7719 15339 7761 15381
rect 7659 15222 7701 15264
rect 8019 15459 8061 15501
rect 8439 15996 8481 16038
rect 8679 16122 8721 16164
rect 9279 16899 9321 16941
rect 9399 16899 9441 16941
rect 9039 16539 9081 16581
rect 9159 16539 9201 16581
rect 8979 16359 9021 16401
rect 9099 16359 9141 16401
rect 9099 16119 9141 16161
rect 8319 15939 8361 15981
rect 8319 15639 8361 15681
rect 8139 15579 8181 15621
rect 8259 15519 8301 15561
rect 7899 15339 7941 15381
rect 8079 15339 8121 15381
rect 7839 15279 7881 15321
rect 7839 15216 7881 15258
rect 7359 15096 7401 15138
rect 7059 15039 7101 15081
rect 7239 15039 7281 15081
rect 7239 14919 7281 14961
rect 7179 14739 7221 14781
rect 7059 14679 7101 14721
rect 6639 14562 6681 14604
rect 6819 14559 6861 14601
rect 6579 14436 6621 14478
rect 6699 14436 6741 14478
rect 6999 14619 7041 14661
rect 7299 14679 7341 14721
rect 6879 14436 6921 14478
rect 6759 14199 6801 14241
rect 6579 14019 6621 14061
rect 6459 13719 6501 13761
rect 6399 13662 6441 13704
rect 6339 13536 6381 13578
rect 5979 13059 6021 13101
rect 5199 12159 5241 12201
rect 5619 12159 5661 12201
rect 5739 12162 5781 12204
rect 5919 12819 5961 12861
rect 5979 12639 6021 12681
rect 5919 12579 5961 12621
rect 5439 12102 5481 12144
rect 5379 11976 5421 12018
rect 5319 11919 5361 11961
rect 5379 11859 5421 11901
rect 5499 11859 5541 11901
rect 5319 11799 5361 11841
rect 5259 11739 5301 11781
rect 5259 11619 5301 11661
rect 5199 11559 5241 11601
rect 5139 11499 5181 11541
rect 5739 12099 5781 12141
rect 5679 11976 5721 12018
rect 5919 12102 5961 12144
rect 6219 13419 6261 13461
rect 6519 13539 6561 13581
rect 6639 13719 6681 13761
rect 6579 13479 6621 13521
rect 6516 13419 6558 13461
rect 6579 13416 6621 13458
rect 6459 13359 6501 13401
rect 6399 13179 6441 13221
rect 6219 12819 6261 12861
rect 6279 12699 6321 12741
rect 6159 12339 6201 12381
rect 5559 11799 5601 11841
rect 5679 11619 5721 11661
rect 5559 11559 5601 11601
rect 5319 11439 5361 11481
rect 5739 11559 5781 11601
rect 5679 11439 5721 11481
rect 5019 11316 5061 11358
rect 5139 11316 5181 11358
rect 5319 11319 5361 11361
rect 5079 11253 5121 11295
rect 5019 11199 5061 11241
rect 5259 11196 5301 11238
rect 4959 10959 5001 11001
rect 5139 10959 5181 11001
rect 4959 10896 5001 10938
rect 5199 10839 5241 10881
rect 5499 11316 5541 11358
rect 6159 12102 6201 12144
rect 6579 12699 6621 12741
rect 6339 12339 6381 12381
rect 5919 11859 5961 11901
rect 6279 11979 6321 12021
rect 6099 11799 6141 11841
rect 6039 11559 6081 11601
rect 5799 11436 5841 11478
rect 5919 11442 5961 11484
rect 5379 11199 5421 11241
rect 5499 11199 5541 11241
rect 5319 11139 5361 11181
rect 5739 11259 5781 11301
rect 5379 11079 5421 11121
rect 5499 11079 5541 11121
rect 5439 11019 5481 11061
rect 5259 10779 5301 10821
rect 5199 10719 5241 10761
rect 5139 10599 5181 10641
rect 5019 10542 5061 10584
rect 4599 10119 4641 10161
rect 4839 10119 4881 10161
rect 4539 9879 4581 9921
rect 4239 9399 4281 9441
rect 4479 9756 4521 9798
rect 4479 9579 4521 9621
rect 4359 9339 4401 9381
rect 4359 8982 4401 9024
rect 4479 8982 4521 9024
rect 4299 8856 4341 8898
rect 4539 8859 4581 8901
rect 4179 8739 4221 8781
rect 4419 8739 4461 8781
rect 4479 8379 4521 8421
rect 4659 9999 4701 10041
rect 4839 9999 4881 10041
rect 4719 9756 4761 9798
rect 4959 10416 5001 10458
rect 5319 10542 5361 10584
rect 5619 10959 5661 11001
rect 5559 10659 5601 10701
rect 5199 10479 5241 10521
rect 5139 10359 5181 10401
rect 5319 10359 5361 10401
rect 4959 10299 5001 10341
rect 5199 10299 5241 10341
rect 5259 9999 5301 10041
rect 4959 9939 5001 9981
rect 5139 9939 5181 9981
rect 4959 9876 5001 9918
rect 5499 10416 5541 10458
rect 5379 10299 5421 10341
rect 5379 9939 5421 9981
rect 5319 9879 5361 9921
rect 5019 9759 5061 9801
rect 4959 9579 5001 9621
rect 5019 9519 5061 9561
rect 5139 9639 5181 9681
rect 4899 9399 4941 9441
rect 5079 9399 5121 9441
rect 5319 9759 5361 9801
rect 5199 9579 5241 9621
rect 5139 9339 5181 9381
rect 5019 9279 5061 9321
rect 4839 9219 4881 9261
rect 5259 9219 5301 9261
rect 5016 9159 5058 9201
rect 5079 9159 5121 9201
rect 4839 9099 4881 9141
rect 5181 9039 5223 9081
rect 5079 8979 5121 9021
rect 5379 9579 5421 9621
rect 5319 9159 5361 9201
rect 5679 10779 5721 10821
rect 5979 11316 6021 11358
rect 6099 11259 6141 11301
rect 5859 11079 5901 11121
rect 5919 10899 5961 10941
rect 5859 10839 5901 10881
rect 5739 10719 5781 10761
rect 5679 10539 5721 10581
rect 6279 11859 6321 11901
rect 6279 11259 6321 11301
rect 6399 12159 6441 12201
rect 6519 12339 6561 12381
rect 7239 14439 7281 14481
rect 7119 14379 7161 14421
rect 7179 14199 7221 14241
rect 7059 14079 7101 14121
rect 6999 13959 7041 14001
rect 6879 13839 6921 13881
rect 6879 13419 6921 13461
rect 6879 13239 6921 13281
rect 6759 12399 6801 12441
rect 6759 12336 6801 12378
rect 6639 12159 6681 12201
rect 6459 12102 6501 12144
rect 6639 12096 6681 12138
rect 7299 14139 7341 14181
rect 7239 14079 7281 14121
rect 7179 13959 7221 14001
rect 7299 13839 7341 13881
rect 7119 13779 7161 13821
rect 7059 13662 7101 13704
rect 7479 15096 7521 15138
rect 7719 15096 7761 15138
rect 7419 14739 7461 14781
rect 7536 14739 7578 14781
rect 7599 14739 7641 14781
rect 7779 14739 7821 14781
rect 7839 14679 7881 14721
rect 7779 14619 7821 14661
rect 7839 14379 7881 14421
rect 7599 14259 7641 14301
rect 7599 13779 7641 13821
rect 7839 13779 7881 13821
rect 7359 13599 7401 13641
rect 7059 13479 7101 13521
rect 7359 13359 7401 13401
rect 7419 13299 7461 13341
rect 7299 13239 7341 13281
rect 7479 13239 7521 13281
rect 7599 13239 7641 13281
rect 7239 13179 7281 13221
rect 7359 13119 7401 13161
rect 7299 13059 7341 13101
rect 7059 12999 7101 13041
rect 7239 12999 7281 13041
rect 8079 15222 8121 15264
rect 8139 15096 8181 15138
rect 8559 15996 8601 16038
rect 8619 15999 8661 16041
rect 8859 15999 8901 16041
rect 8619 15819 8661 15861
rect 8499 15279 8541 15321
rect 8439 15222 8481 15264
rect 8739 15939 8781 15981
rect 8679 15759 8721 15801
rect 8799 15759 8841 15801
rect 8739 15579 8781 15621
rect 8439 15039 8481 15081
rect 8379 14679 8421 14721
rect 8259 14559 8301 14601
rect 8019 14436 8061 14478
rect 8139 14436 8181 14478
rect 8079 13959 8121 14001
rect 7959 13779 8001 13821
rect 8259 14436 8301 14478
rect 8199 13899 8241 13941
rect 7959 13299 8001 13341
rect 8079 13299 8121 13341
rect 7899 13179 7941 13221
rect 7119 12639 7161 12681
rect 6879 12219 6921 12261
rect 6999 12219 7041 12261
rect 6999 12102 7041 12144
rect 6399 11859 6441 11901
rect 6519 11619 6561 11661
rect 6699 11739 6741 11781
rect 6639 11499 6681 11541
rect 7059 11979 7101 12021
rect 6819 11619 6861 11661
rect 6759 11499 6801 11541
rect 6579 11439 6621 11481
rect 6699 11439 6741 11481
rect 6576 11316 6618 11358
rect 6639 11316 6681 11358
rect 6459 11259 6501 11301
rect 6276 11139 6318 11181
rect 6339 11139 6381 11181
rect 6099 10539 6141 10581
rect 6639 11253 6681 11295
rect 6399 11079 6441 11121
rect 6459 10959 6501 11001
rect 5499 10299 5541 10341
rect 5619 10299 5661 10341
rect 5859 10416 5901 10458
rect 5799 10239 5841 10281
rect 5679 10119 5721 10161
rect 5619 10059 5661 10101
rect 5499 9879 5541 9921
rect 5739 9882 5781 9924
rect 6159 10359 6201 10401
rect 6099 10239 6141 10281
rect 6039 10179 6081 10221
rect 5979 10119 6021 10161
rect 6039 10059 6081 10101
rect 6039 9996 6081 10038
rect 6399 10419 6441 10461
rect 6339 10359 6381 10401
rect 6399 10299 6441 10341
rect 6219 10179 6261 10221
rect 6579 10719 6621 10761
rect 7239 12879 7281 12921
rect 8019 13179 8061 13221
rect 8199 13239 8241 13281
rect 8139 13179 8181 13221
rect 8079 13059 8121 13101
rect 8199 13119 8241 13161
rect 8739 15099 8781 15141
rect 9099 15999 9141 16041
rect 9039 15699 9081 15741
rect 9579 17439 9621 17481
rect 9519 16782 9561 16824
rect 9699 17379 9741 17421
rect 9699 17259 9741 17301
rect 9699 17019 9741 17061
rect 10119 18519 10161 18561
rect 9879 18399 9921 18441
rect 9999 18399 10041 18441
rect 10359 18342 10401 18384
rect 10479 18342 10521 18384
rect 11139 18459 11181 18501
rect 11439 18459 11481 18501
rect 10719 18342 10761 18384
rect 10839 18342 10881 18384
rect 10959 18342 11001 18384
rect 9879 18219 9921 18261
rect 10179 18099 10221 18141
rect 10359 18099 10401 18141
rect 10479 17919 10521 17961
rect 9819 17799 9861 17841
rect 10059 17799 10101 17841
rect 9999 17682 10041 17724
rect 10119 17682 10161 17724
rect 10359 17682 10401 17724
rect 10659 17979 10701 18021
rect 10539 17739 10581 17781
rect 11019 18216 11061 18258
rect 11319 18342 11361 18384
rect 10899 18099 10941 18141
rect 11139 18099 11181 18141
rect 11319 18039 11361 18081
rect 10719 17919 10761 17961
rect 11259 17919 11301 17961
rect 10839 17739 10881 17781
rect 11019 17739 11061 17781
rect 11079 17679 11121 17721
rect 11379 17979 11421 18021
rect 11019 17619 11061 17661
rect 9939 17556 9981 17598
rect 10059 17556 10101 17598
rect 10059 17493 10101 17535
rect 9819 17319 9861 17361
rect 9999 17199 10041 17241
rect 9759 16899 9801 16941
rect 10179 17439 10221 17481
rect 10239 17379 10281 17421
rect 10119 17139 10161 17181
rect 10059 16959 10101 17001
rect 9819 16779 9861 16821
rect 9999 16782 10041 16824
rect 9639 16656 9681 16698
rect 9519 16479 9561 16521
rect 9399 16419 9441 16461
rect 9219 16359 9261 16401
rect 9699 16419 9741 16461
rect 9639 16299 9681 16341
rect 9579 16239 9621 16281
rect 9399 16179 9441 16221
rect 9519 16179 9561 16221
rect 9459 15996 9501 16038
rect 9579 15999 9621 16041
rect 9279 15819 9321 15861
rect 9639 15819 9681 15861
rect 9519 15699 9561 15741
rect 9639 15699 9681 15741
rect 9159 15639 9201 15681
rect 8919 15519 8961 15561
rect 9039 15519 9081 15561
rect 8919 15456 8961 15498
rect 8919 15222 8961 15264
rect 9039 15222 9081 15264
rect 8799 14919 8841 14961
rect 8499 14859 8541 14901
rect 8499 14679 8541 14721
rect 8499 14562 8541 14604
rect 8619 14562 8661 14604
rect 8379 14439 8421 14481
rect 8559 14436 8601 14478
rect 8679 14199 8721 14241
rect 8619 13899 8661 13941
rect 8439 13662 8481 13704
rect 8499 13536 8541 13578
rect 8439 13479 8481 13521
rect 8379 13299 8421 13341
rect 8319 13179 8361 13221
rect 8379 13119 8421 13161
rect 8259 13002 8301 13044
rect 8379 12999 8421 13041
rect 8739 14079 8781 14121
rect 8979 15096 9021 15138
rect 9339 15459 9381 15501
rect 9459 15459 9501 15501
rect 9159 15039 9201 15081
rect 8859 14859 8901 14901
rect 9159 14859 9201 14901
rect 8979 14679 9021 14721
rect 9159 14679 9201 14721
rect 9099 14562 9141 14604
rect 8919 14379 8961 14421
rect 8799 13899 8841 13941
rect 8799 13779 8841 13821
rect 8859 13719 8901 13761
rect 8679 13659 8721 13701
rect 9099 14379 9141 14421
rect 9039 14139 9081 14181
rect 9099 14079 9141 14121
rect 9039 13719 9081 13761
rect 8619 13359 8661 13401
rect 8739 13536 8781 13578
rect 8859 13536 8901 13578
rect 9039 13536 9081 13578
rect 8739 13419 8781 13461
rect 9279 15096 9321 15138
rect 9519 15096 9561 15138
rect 9519 14799 9561 14841
rect 9399 14739 9441 14781
rect 9939 16656 9981 16698
rect 9999 16539 10041 16581
rect 9819 16299 9861 16341
rect 9879 16179 9921 16221
rect 10059 16419 10101 16461
rect 10179 16419 10221 16461
rect 10059 16356 10101 16398
rect 9999 16119 10041 16161
rect 9759 15999 9801 16041
rect 9939 15996 9981 16038
rect 9999 15699 10041 15741
rect 9759 15579 9801 15621
rect 9819 15399 9861 15441
rect 9879 15222 9921 15264
rect 10119 16179 10161 16221
rect 10539 17556 10581 17598
rect 10659 17559 10701 17601
rect 10659 17439 10701 17481
rect 10419 17319 10461 17361
rect 10299 16959 10341 17001
rect 10539 16959 10581 17001
rect 10419 16782 10461 16824
rect 10899 17556 10941 17598
rect 11079 17556 11121 17598
rect 10779 17319 10821 17361
rect 10779 17256 10821 17298
rect 10659 16782 10701 16824
rect 10299 16599 10341 16641
rect 10239 16179 10281 16221
rect 10416 16479 10458 16521
rect 10479 16479 10521 16521
rect 10479 16416 10521 16458
rect 10719 16659 10761 16701
rect 10659 16599 10701 16641
rect 10599 16359 10641 16401
rect 10599 16239 10641 16281
rect 10479 16179 10521 16221
rect 10599 16119 10641 16161
rect 10719 16419 10761 16461
rect 10779 16359 10821 16401
rect 10959 17319 11001 17361
rect 11379 17556 11421 17598
rect 11079 17139 11121 17181
rect 11019 16959 11061 17001
rect 11079 16782 11121 16824
rect 10899 16659 10941 16701
rect 11019 16656 11061 16698
rect 10959 16539 11001 16581
rect 10899 16476 10941 16518
rect 10899 16299 10941 16341
rect 10779 16122 10821 16164
rect 10119 15999 10161 16041
rect 10059 15639 10101 15681
rect 9819 15096 9861 15138
rect 10059 15096 10101 15138
rect 9939 15039 9981 15081
rect 9639 14859 9681 14901
rect 9579 14679 9621 14721
rect 9459 14562 9501 14604
rect 9219 13959 9261 14001
rect 9279 13779 9321 13821
rect 9279 13659 9321 13701
rect 9579 14436 9621 14478
rect 9519 14379 9561 14421
rect 9699 14559 9741 14601
rect 9459 13659 9501 13701
rect 9219 13536 9261 13578
rect 9399 13479 9441 13521
rect 8799 13299 8841 13341
rect 9099 13299 9141 13341
rect 8739 13119 8781 13161
rect 8679 12999 8721 13041
rect 8079 12879 8121 12921
rect 7959 12819 8001 12861
rect 7479 12759 7521 12801
rect 7299 12399 7341 12441
rect 7419 12279 7461 12321
rect 7419 12159 7461 12201
rect 6996 11439 7038 11481
rect 7059 11442 7101 11484
rect 6819 11319 6861 11361
rect 6936 11316 6978 11358
rect 6999 11319 7041 11361
rect 7119 11259 7161 11301
rect 6879 11199 6921 11241
rect 6999 11199 7041 11241
rect 6819 10719 6861 10761
rect 6699 10542 6741 10584
rect 6939 11139 6981 11181
rect 6879 10539 6921 10581
rect 6879 10419 6921 10461
rect 6759 10299 6801 10341
rect 6819 10239 6861 10281
rect 6639 10179 6681 10221
rect 6759 10179 6801 10221
rect 6579 9999 6621 10041
rect 6159 9939 6201 9981
rect 6459 9939 6501 9981
rect 5859 9882 5901 9924
rect 6039 9882 6081 9924
rect 6399 9882 6441 9924
rect 5499 9759 5541 9801
rect 5439 9039 5481 9081
rect 4719 8859 4761 8901
rect 4659 8799 4701 8841
rect 4659 8619 4701 8661
rect 4659 8439 4701 8481
rect 4299 8322 4341 8364
rect 4599 8319 4641 8361
rect 4479 8196 4521 8238
rect 4599 8199 4641 8241
rect 4359 8079 4401 8121
rect 4239 8019 4281 8061
rect 4179 7719 4221 7761
rect 4119 7659 4161 7701
rect 3759 7479 3801 7521
rect 3699 7419 3741 7461
rect 3939 7422 3981 7464
rect 3279 7179 3321 7221
rect 3399 7179 3441 7221
rect 3339 7119 3381 7161
rect 3459 7119 3501 7161
rect 3216 7059 3258 7101
rect 3279 7059 3321 7101
rect 3039 6762 3081 6804
rect 3159 6762 3201 6804
rect 2919 6639 2961 6681
rect 3219 6519 3261 6561
rect 3999 7296 4041 7338
rect 4119 7299 4161 7341
rect 4119 7179 4161 7221
rect 3699 7119 3741 7161
rect 3999 6999 4041 7041
rect 3519 6939 3561 6981
rect 3819 6939 3861 6981
rect 3459 6879 3501 6921
rect 3579 6879 3621 6921
rect 3519 6762 3561 6804
rect 3639 6762 3681 6804
rect 3999 6762 4041 6804
rect 4239 7539 4281 7581
rect 4179 6999 4221 7041
rect 4479 7479 4521 7521
rect 4239 6939 4281 6981
rect 5079 8859 5121 8901
rect 4899 8799 4941 8841
rect 5019 8679 5061 8721
rect 4899 8619 4941 8661
rect 4839 8559 4881 8601
rect 4779 8439 4821 8481
rect 4959 8499 5001 8541
rect 4719 8319 4761 8361
rect 4719 8199 4761 8241
rect 4839 8196 4881 8238
rect 4659 7719 4701 7761
rect 4719 7659 4761 7701
rect 4539 7239 4581 7281
rect 4419 7059 4461 7101
rect 4659 7059 4701 7101
rect 4359 6999 4401 7041
rect 4299 6819 4341 6861
rect 4479 6819 4521 6861
rect 3459 6519 3501 6561
rect 3699 6636 3741 6678
rect 3819 6636 3861 6678
rect 3939 6636 3981 6678
rect 3939 6519 3981 6561
rect 3339 6459 3381 6501
rect 3579 6459 3621 6501
rect 3819 6459 3861 6501
rect 3939 6339 3981 6381
rect 3099 6159 3141 6201
rect 2979 5979 3021 6021
rect 2859 5862 2901 5904
rect 4119 6579 4161 6621
rect 4059 6099 4101 6141
rect 3459 5919 3501 5961
rect 3939 5919 3981 5961
rect 3099 5862 3141 5904
rect 2919 5736 2961 5778
rect 3039 5736 3081 5778
rect 2859 5379 2901 5421
rect 2799 5199 2841 5241
rect 3339 5862 3381 5904
rect 3699 5862 3741 5904
rect 3819 5862 3861 5904
rect 3519 5736 3561 5778
rect 3219 5619 3261 5661
rect 3399 5619 3441 5661
rect 3219 5439 3261 5481
rect 2979 5202 3021 5244
rect 2919 5076 2961 5118
rect 3279 5076 3321 5118
rect 4059 5859 4101 5901
rect 3759 5439 3801 5481
rect 3459 5319 3501 5361
rect 3039 5019 3081 5061
rect 3399 5019 3441 5061
rect 2979 4779 3021 4821
rect 3099 4779 3141 4821
rect 2979 4659 3021 4701
rect 2739 4419 2781 4461
rect 2859 4359 2901 4401
rect 2379 4059 2421 4101
rect 2559 3879 2601 3921
rect 2139 3819 2181 3861
rect 2259 3819 2301 3861
rect 2439 3759 2481 3801
rect 2199 3639 2241 3681
rect 2319 3642 2361 3684
rect 2559 3639 2601 3681
rect 1839 3516 1881 3558
rect 1959 3516 2001 3558
rect 2139 3516 2181 3558
rect 1659 3399 1701 3441
rect 1059 2319 1101 2361
rect 1419 2616 1461 2658
rect 1599 2616 1641 2658
rect 1719 2616 1761 2658
rect 1959 3399 2001 3441
rect 1899 2799 1941 2841
rect 1299 2499 1341 2541
rect 1839 2499 1881 2541
rect 1179 2259 1221 2301
rect 1179 2082 1221 2124
rect 1299 2082 1341 2124
rect 1479 2079 1521 2121
rect 939 1956 981 1998
rect 1059 1956 1101 1998
rect 1239 1899 1281 1941
rect 1059 1839 1101 1881
rect 1359 1839 1401 1881
rect 819 1719 861 1761
rect 1239 1479 1281 1521
rect 759 1419 801 1461
rect 639 1239 681 1281
rect 579 1179 621 1221
rect 939 1239 981 1281
rect 399 1056 441 1098
rect 699 939 741 981
rect 279 819 321 861
rect 399 819 441 861
rect 39 699 81 741
rect 279 699 321 741
rect 1479 1299 1521 1341
rect 1599 2259 1641 2301
rect 1719 2319 1761 2361
rect 1659 2199 1701 2241
rect 1599 2079 1641 2121
rect 1839 2199 1881 2241
rect 1899 2079 1941 2121
rect 1659 1956 1701 1998
rect 1779 1899 1821 1941
rect 1779 1719 1821 1761
rect 1659 1479 1701 1521
rect 1539 1182 1581 1224
rect 1839 1299 1881 1341
rect 1299 1056 1341 1098
rect 939 939 981 981
rect 1179 939 1221 981
rect 819 699 861 741
rect 759 639 801 681
rect 1719 1056 1761 1098
rect 1599 879 1641 921
rect 1479 819 1521 861
rect 1239 699 1281 741
rect 1179 579 1221 621
rect 819 519 861 561
rect 939 519 981 561
rect 1119 522 1161 564
rect 1239 522 1281 564
rect 1599 759 1641 801
rect 339 396 381 438
rect 459 396 501 438
rect 699 396 741 438
rect 1059 396 1101 438
rect 1179 396 1221 438
rect 1419 339 1461 381
rect 1899 1182 1941 1224
rect 1899 1059 1941 1101
rect 2079 2742 2121 2784
rect 2379 3516 2421 3558
rect 2499 3516 2541 3558
rect 2859 4119 2901 4161
rect 2799 4059 2841 4101
rect 2739 3642 2781 3684
rect 3039 3999 3081 4041
rect 2919 3759 2961 3801
rect 2799 3459 2841 3501
rect 2619 3399 2661 3441
rect 2559 3279 2601 3321
rect 2499 3219 2541 3261
rect 2559 3159 2601 3201
rect 2319 2859 2361 2901
rect 2559 2799 2601 2841
rect 2679 2742 2721 2784
rect 2319 2619 2361 2661
rect 2979 3519 3021 3561
rect 2499 2616 2541 2658
rect 2799 2616 2841 2658
rect 2439 2499 2481 2541
rect 2619 2499 2661 2541
rect 2379 2319 2421 2361
rect 2139 2259 2181 2301
rect 2259 2199 2301 2241
rect 2019 2079 2061 2121
rect 2919 3099 2961 3141
rect 3219 4539 3261 4581
rect 3159 4419 3201 4461
rect 3159 4119 3201 4161
rect 3639 5319 3681 5361
rect 3999 5736 4041 5778
rect 4419 6636 4461 6678
rect 4536 6636 4578 6678
rect 4599 6639 4641 6681
rect 4299 6579 4341 6621
rect 4179 6459 4221 6501
rect 4179 6219 4221 6261
rect 4239 6159 4281 6201
rect 4179 5859 4221 5901
rect 4359 6099 4401 6141
rect 4599 6399 4641 6441
rect 5139 8799 5181 8841
rect 5199 8739 5241 8781
rect 5439 8799 5481 8841
rect 5679 9756 5721 9798
rect 5559 9399 5601 9441
rect 5559 9279 5601 9321
rect 5739 9279 5781 9321
rect 5679 9099 5721 9141
rect 5859 9339 5901 9381
rect 5799 9099 5841 9141
rect 5799 8979 5841 9021
rect 5499 8679 5541 8721
rect 5739 8856 5781 8898
rect 5979 9756 6021 9798
rect 6039 9699 6081 9741
rect 6159 9699 6201 9741
rect 6219 9759 6261 9801
rect 6219 9639 6261 9681
rect 6159 9579 6201 9621
rect 6039 9459 6081 9501
rect 5979 9099 6021 9141
rect 5859 8799 5901 8841
rect 5619 8619 5661 8661
rect 5379 8379 5421 8421
rect 5319 8322 5361 8364
rect 5499 8322 5541 8364
rect 5079 8199 5121 8241
rect 5259 8196 5301 8238
rect 5379 8196 5421 8238
rect 5019 8139 5061 8181
rect 5196 8139 5238 8181
rect 4959 8079 5001 8121
rect 4899 7899 4941 7941
rect 5079 7779 5121 7821
rect 4959 7719 5001 7761
rect 4779 7599 4821 7641
rect 4839 7422 4881 7464
rect 5139 7479 5181 7521
rect 5079 7422 5121 7464
rect 4899 7239 4941 7281
rect 5079 7299 5121 7341
rect 4779 7119 4821 7161
rect 5019 7119 5061 7161
rect 5139 7239 5181 7281
rect 5559 8259 5601 8301
rect 5499 8079 5541 8121
rect 5619 8139 5661 8181
rect 5559 7959 5601 8001
rect 5439 7779 5481 7821
rect 5559 7779 5601 7821
rect 5379 7719 5421 7761
rect 5439 7659 5481 7701
rect 5259 7599 5301 7641
rect 5499 7599 5541 7641
rect 5439 7539 5481 7581
rect 5319 7479 5361 7521
rect 5259 7419 5301 7461
rect 5439 7422 5481 7464
rect 5259 7296 5301 7338
rect 5199 7179 5241 7221
rect 5199 7116 5241 7158
rect 4959 6999 5001 7041
rect 5079 6999 5121 7041
rect 5079 6936 5121 6978
rect 4959 6879 5001 6921
rect 4899 6819 4941 6861
rect 5499 7296 5541 7338
rect 5379 7239 5421 7281
rect 5679 8079 5721 8121
rect 5679 7959 5721 8001
rect 5739 7779 5781 7821
rect 6099 9099 6141 9141
rect 6039 8979 6081 9021
rect 6399 9699 6441 9741
rect 6339 9579 6381 9621
rect 6219 9159 6261 9201
rect 6519 9759 6561 9801
rect 6579 9699 6621 9741
rect 6519 9519 6561 9561
rect 6459 9459 6501 9501
rect 6999 11079 7041 11121
rect 6939 10119 6981 10161
rect 6759 10059 6801 10101
rect 8199 12759 8241 12801
rect 7959 12639 8001 12681
rect 8079 12639 8121 12681
rect 7599 12519 7641 12561
rect 7719 12459 7761 12501
rect 7899 12339 7941 12381
rect 7839 12159 7881 12201
rect 8139 12459 8181 12501
rect 8079 12279 8121 12321
rect 8019 12216 8061 12258
rect 7959 12159 8001 12201
rect 7899 12099 7941 12141
rect 7719 11976 7761 12018
rect 7599 11679 7641 11721
rect 7839 11679 7881 11721
rect 7959 11679 8001 11721
rect 7659 11559 7701 11601
rect 7419 11499 7461 11541
rect 7539 11499 7581 11541
rect 7359 11439 7401 11481
rect 7839 11556 7881 11598
rect 7779 11442 7821 11484
rect 7899 11439 7941 11481
rect 7179 11199 7221 11241
rect 7239 11019 7281 11061
rect 7056 10899 7098 10941
rect 7119 10899 7161 10941
rect 7119 10719 7161 10761
rect 7059 10539 7101 10581
rect 7479 11319 7521 11361
rect 7359 11259 7401 11301
rect 7299 10959 7341 11001
rect 7299 10779 7341 10821
rect 7239 10539 7281 10581
rect 7179 10416 7221 10458
rect 6819 9999 6861 10041
rect 6999 9999 7041 10041
rect 6699 9759 6741 9801
rect 6699 9579 6741 9621
rect 6819 9579 6861 9621
rect 6939 9579 6981 9621
rect 6759 9459 6801 9501
rect 6639 9339 6681 9381
rect 6399 9279 6441 9321
rect 6339 8979 6381 9021
rect 6216 8856 6258 8898
rect 6279 8859 6321 8901
rect 6099 8799 6141 8841
rect 6039 8619 6081 8661
rect 5919 8319 5961 8361
rect 6159 8559 6201 8601
rect 6159 8439 6201 8481
rect 5979 8196 6021 8238
rect 6039 8139 6081 8181
rect 6039 8019 6081 8061
rect 5859 7479 5901 7521
rect 5676 7419 5718 7461
rect 5739 7422 5781 7464
rect 5979 7359 6021 7401
rect 5679 7299 5721 7341
rect 5619 7179 5661 7221
rect 5559 7119 5601 7161
rect 5439 6939 5481 6981
rect 5259 6879 5301 6921
rect 5379 6879 5421 6921
rect 5139 6762 5181 6804
rect 5319 6762 5361 6804
rect 5619 6999 5661 7041
rect 5556 6819 5598 6861
rect 5739 7239 5781 7281
rect 5919 7299 5961 7341
rect 5799 7179 5841 7221
rect 5859 7119 5901 7161
rect 5739 6999 5781 7041
rect 5799 6819 5841 6861
rect 4779 6459 4821 6501
rect 4959 6636 5001 6678
rect 5679 6759 5721 6801
rect 5919 7059 5961 7101
rect 6099 7839 6141 7881
rect 6279 8499 6321 8541
rect 6399 8859 6441 8901
rect 6579 9219 6621 9261
rect 6519 9099 6561 9141
rect 6939 9516 6981 9558
rect 6939 9279 6981 9321
rect 7116 10119 7158 10161
rect 7179 10119 7221 10161
rect 7299 10119 7341 10161
rect 7419 10839 7461 10881
rect 7659 11259 7701 11301
rect 7599 11079 7641 11121
rect 7479 10779 7521 10821
rect 7719 11199 7761 11241
rect 7959 11259 8001 11301
rect 7899 10899 7941 10941
rect 7719 10599 7761 10641
rect 7659 10539 7701 10581
rect 8259 12102 8301 12144
rect 8439 12879 8481 12921
rect 8379 12819 8421 12861
rect 8079 11976 8121 12018
rect 8199 11976 8241 12018
rect 8319 11919 8361 11961
rect 8259 11619 8301 11661
rect 8079 11559 8121 11601
rect 8139 11499 8181 11541
rect 8079 11439 8121 11481
rect 8619 12519 8661 12561
rect 8499 12279 8541 12321
rect 8559 12219 8601 12261
rect 8439 12159 8481 12201
rect 8559 12102 8601 12144
rect 8679 12459 8721 12501
rect 8379 11559 8421 11601
rect 8379 11496 8421 11538
rect 8499 11976 8541 12018
rect 8619 11979 8661 12021
rect 8619 11859 8661 11901
rect 9159 13239 9201 13281
rect 8799 12999 8841 13041
rect 8919 12879 8961 12921
rect 9039 12759 9081 12801
rect 8859 12579 8901 12621
rect 9039 12459 9081 12501
rect 8799 12099 8841 12141
rect 8739 11979 8781 12021
rect 8799 11679 8841 11721
rect 8739 11619 8781 11661
rect 8679 11499 8721 11541
rect 8559 11442 8601 11484
rect 8079 11319 8121 11361
rect 7959 10779 8001 10821
rect 7719 10479 7761 10521
rect 7419 10419 7461 10461
rect 7359 10059 7401 10101
rect 7119 9876 7161 9918
rect 7299 9882 7341 9924
rect 7539 10359 7581 10401
rect 7779 10419 7821 10461
rect 7719 10299 7761 10341
rect 7539 10179 7581 10221
rect 7479 9999 7521 10041
rect 7419 9879 7461 9921
rect 7059 9519 7101 9561
rect 7179 9639 7221 9681
rect 7299 9639 7341 9681
rect 7119 9399 7161 9441
rect 7239 9279 7281 9321
rect 6819 9159 6861 9201
rect 6879 9099 6921 9141
rect 6699 8982 6741 9024
rect 7179 9159 7221 9201
rect 6939 9039 6981 9081
rect 6999 8982 7041 9024
rect 6579 8799 6621 8841
rect 6519 8739 6561 8781
rect 6459 8619 6501 8661
rect 6519 8559 6561 8601
rect 6399 8439 6441 8481
rect 6819 8859 6861 8901
rect 6699 8739 6741 8781
rect 6699 8619 6741 8661
rect 6639 8499 6681 8541
rect 6519 8379 6561 8421
rect 6279 8319 6321 8361
rect 6399 8322 6441 8364
rect 6219 7779 6261 7821
rect 6039 7299 6081 7341
rect 6039 7059 6081 7101
rect 6039 6879 6081 6921
rect 6039 6816 6081 6858
rect 5859 6759 5901 6801
rect 5259 6579 5301 6621
rect 5379 6579 5421 6621
rect 4959 6519 5001 6561
rect 5139 6519 5181 6561
rect 4839 6399 4881 6441
rect 4839 6336 4881 6378
rect 4779 6219 4821 6261
rect 4599 6159 4641 6201
rect 4719 6159 4761 6201
rect 4419 5979 4461 6021
rect 5199 6459 5241 6501
rect 5019 6399 5061 6441
rect 4959 6159 5001 6201
rect 4776 6099 4818 6141
rect 4839 6099 4881 6141
rect 4479 5859 4521 5901
rect 4599 5862 4641 5904
rect 5139 6279 5181 6321
rect 4839 5862 4881 5904
rect 5139 5979 5181 6021
rect 5079 5862 5121 5904
rect 3939 5619 3981 5661
rect 4119 5619 4161 5661
rect 3879 5199 3921 5241
rect 3579 5079 3621 5121
rect 3519 4539 3561 4581
rect 3279 4419 3321 4461
rect 3459 4419 3501 4461
rect 3279 4299 3321 4341
rect 3699 5076 3741 5118
rect 3819 4959 3861 5001
rect 4179 5379 4221 5421
rect 3999 5259 4041 5301
rect 4599 5619 4641 5661
rect 4359 5319 4401 5361
rect 4479 5319 4521 5361
rect 4299 5259 4341 5301
rect 3999 5139 4041 5181
rect 4299 5139 4341 5181
rect 4119 4959 4161 5001
rect 4239 4779 4281 4821
rect 3939 4599 3981 4641
rect 3699 4419 3741 4461
rect 3999 4419 4041 4461
rect 4119 4419 4161 4461
rect 3579 4302 3621 4344
rect 3819 4302 3861 4344
rect 3279 4179 3321 4221
rect 3099 3879 3141 3921
rect 3099 3639 3141 3681
rect 3039 3459 3081 3501
rect 2979 2979 3021 3021
rect 3219 3939 3261 3981
rect 3459 4119 3501 4161
rect 3759 4119 3801 4161
rect 3339 3999 3381 4041
rect 3759 3939 3801 3981
rect 3279 3819 3321 3861
rect 3399 3819 3441 3861
rect 3579 3819 3621 3861
rect 3279 3642 3321 3684
rect 3219 3519 3261 3561
rect 3159 3459 3201 3501
rect 3159 2979 3201 3021
rect 3099 2799 3141 2841
rect 3039 2742 3081 2784
rect 3999 4119 4041 4161
rect 4059 3879 4101 3921
rect 3879 3759 3921 3801
rect 3999 3759 4041 3801
rect 3879 3642 3921 3684
rect 3459 3459 3501 3501
rect 3939 3519 3981 3561
rect 3819 3339 3861 3381
rect 3339 3219 3381 3261
rect 3819 3219 3861 3261
rect 3579 2979 3621 3021
rect 3219 2919 3261 2961
rect 3699 2919 3741 2961
rect 3279 2799 3321 2841
rect 3459 2799 3501 2841
rect 2859 2559 2901 2601
rect 2799 2319 2841 2361
rect 2496 2199 2538 2241
rect 2559 2199 2601 2241
rect 2439 2079 2481 2121
rect 2199 1956 2241 1998
rect 2019 1899 2061 1941
rect 2319 1839 2361 1881
rect 2499 1719 2541 1761
rect 2379 1419 2421 1461
rect 2079 1182 2121 1224
rect 2199 1182 2241 1224
rect 3099 2559 3141 2601
rect 3879 2859 3921 2901
rect 4479 5202 4521 5244
rect 4659 5439 4701 5481
rect 4779 5439 4821 5481
rect 4719 5379 4761 5421
rect 4719 5199 4761 5241
rect 4659 5076 4701 5118
rect 4539 4899 4581 4941
rect 4899 5739 4941 5781
rect 4839 5256 4881 5298
rect 4959 5439 5001 5481
rect 4899 5199 4941 5241
rect 5556 6639 5598 6681
rect 5619 6639 5661 6681
rect 5499 6279 5541 6321
rect 5559 5859 5601 5901
rect 5079 5619 5121 5661
rect 5259 5679 5301 5721
rect 5139 5559 5181 5601
rect 5079 5439 5121 5481
rect 5019 5379 5061 5421
rect 5079 5259 5121 5301
rect 5316 5559 5358 5601
rect 5379 5559 5421 5601
rect 5259 5136 5301 5178
rect 4839 4959 4881 5001
rect 4779 4719 4821 4761
rect 4479 4599 4521 4641
rect 4299 4419 4341 4461
rect 4419 4419 4461 4461
rect 5019 5076 5061 5118
rect 5139 5019 5181 5061
rect 4659 4539 4701 4581
rect 4836 4539 4878 4581
rect 4899 4539 4941 4581
rect 4539 4479 4581 4521
rect 4479 4359 4521 4401
rect 4779 4479 4821 4521
rect 4299 4176 4341 4218
rect 4539 4176 4581 4218
rect 4359 4119 4401 4161
rect 4839 4176 4881 4218
rect 4659 4119 4701 4161
rect 4719 4119 4761 4161
rect 4659 3879 4701 3921
rect 4539 3759 4581 3801
rect 4299 3642 4341 3684
rect 4839 3699 4881 3741
rect 4839 3579 4881 3621
rect 4119 3516 4161 3558
rect 4239 3516 4281 3558
rect 4059 3459 4101 3501
rect 4419 3519 4461 3561
rect 4359 3459 4401 3501
rect 4419 3339 4461 3381
rect 4239 3279 4281 3321
rect 4539 3279 4581 3321
rect 3999 3099 4041 3141
rect 4839 3219 4881 3261
rect 4119 2919 4161 2961
rect 3999 2859 4041 2901
rect 3999 2742 4041 2784
rect 4119 2742 4161 2784
rect 3399 2616 3441 2658
rect 3279 2379 3321 2421
rect 3459 2379 3501 2421
rect 3279 2199 3321 2241
rect 2679 2082 2721 2124
rect 2799 2082 2841 2124
rect 2979 2082 3021 2124
rect 3159 2082 3201 2124
rect 2619 1959 2661 2001
rect 2739 1956 2781 1998
rect 3399 2079 3441 2121
rect 2739 1779 2781 1821
rect 2859 1719 2901 1761
rect 3219 1719 3261 1761
rect 2619 1599 2661 1641
rect 2559 1359 2601 1401
rect 3699 2616 3741 2658
rect 3939 2616 3981 2658
rect 3519 2199 3561 2241
rect 3699 2199 3741 2241
rect 3879 2199 3921 2241
rect 3819 2139 3861 2181
rect 3579 2082 3621 2124
rect 3699 2082 3741 2124
rect 4719 2919 4761 2961
rect 4719 2799 4761 2841
rect 4599 2742 4641 2784
rect 4899 3039 4941 3081
rect 4899 2859 4941 2901
rect 5439 5439 5481 5481
rect 5499 5259 5541 5301
rect 5739 6636 5781 6678
rect 5859 6639 5901 6681
rect 5979 6639 6021 6681
rect 5679 6519 5721 6561
rect 5919 6396 5961 6438
rect 5679 6339 5721 6381
rect 6339 8199 6381 8241
rect 6459 8139 6501 8181
rect 6459 7959 6501 8001
rect 6399 7719 6441 7761
rect 6399 7599 6441 7641
rect 6279 7479 6321 7521
rect 6399 7479 6441 7521
rect 6459 7419 6501 7461
rect 6279 7296 6321 7338
rect 6159 7179 6201 7221
rect 6276 7059 6318 7101
rect 6339 7059 6381 7101
rect 6339 6939 6381 6981
rect 6639 7839 6681 7881
rect 6579 7479 6621 7521
rect 6759 8499 6801 8541
rect 7119 8859 7161 8901
rect 7059 8799 7101 8841
rect 7179 8799 7221 8841
rect 6999 8559 7041 8601
rect 6939 8499 6981 8541
rect 6879 8439 6921 8481
rect 6819 8379 6861 8421
rect 7419 9759 7461 9801
rect 7359 9399 7401 9441
rect 7659 10119 7701 10161
rect 7599 10059 7641 10101
rect 7539 9519 7581 9561
rect 7419 9279 7461 9321
rect 7419 9099 7461 9141
rect 7899 10239 7941 10281
rect 7659 9996 7701 10038
rect 7779 9999 7821 10041
rect 7659 9879 7701 9921
rect 7779 9882 7821 9924
rect 7719 9756 7761 9798
rect 7719 9693 7761 9735
rect 7839 9699 7881 9741
rect 7779 9459 7821 9501
rect 7719 9339 7761 9381
rect 7539 8856 7581 8898
rect 7359 8799 7401 8841
rect 7299 8739 7341 8781
rect 7239 8679 7281 8721
rect 7179 8559 7221 8601
rect 7059 8319 7101 8361
rect 7419 8739 7461 8781
rect 7239 8322 7281 8364
rect 6759 8079 6801 8121
rect 6999 8199 7041 8241
rect 6819 7899 6861 7941
rect 6699 7659 6741 7701
rect 6639 7419 6681 7461
rect 6939 7779 6981 7821
rect 6879 7599 6921 7641
rect 6759 7419 6801 7461
rect 6759 7299 6801 7341
rect 6639 7239 6681 7281
rect 6579 6879 6621 6921
rect 6279 6762 6321 6804
rect 6456 6759 6498 6801
rect 6099 6459 6141 6501
rect 5976 6279 6018 6321
rect 6039 6279 6081 6321
rect 5919 6219 5961 6261
rect 5799 5862 5841 5904
rect 5679 5799 5721 5841
rect 5859 5736 5901 5778
rect 5919 5619 5961 5661
rect 5799 5439 5841 5481
rect 5859 5259 5901 5301
rect 5439 5019 5481 5061
rect 5259 4899 5301 4941
rect 5199 4839 5241 4881
rect 5316 4719 5358 4761
rect 5379 4719 5421 4761
rect 5139 4302 5181 4344
rect 5019 4179 5061 4221
rect 5199 4176 5241 4218
rect 5559 4659 5601 4701
rect 5379 4539 5421 4581
rect 5559 4539 5601 4581
rect 5799 5076 5841 5118
rect 5739 4899 5781 4941
rect 5979 5439 6021 5481
rect 6099 6219 6141 6261
rect 6099 6099 6141 6141
rect 6219 6636 6261 6678
rect 6276 6219 6318 6261
rect 6339 6219 6381 6261
rect 6279 6099 6321 6141
rect 6219 6039 6261 6081
rect 6219 5919 6261 5961
rect 6339 5919 6381 5961
rect 6519 6756 6561 6798
rect 7299 8196 7341 8238
rect 7239 8139 7281 8181
rect 7119 7899 7161 7941
rect 7299 8079 7341 8121
rect 7479 8679 7521 8721
rect 7239 7779 7281 7821
rect 7239 7716 7281 7758
rect 7059 7479 7101 7521
rect 6999 7419 7041 7461
rect 7359 8019 7401 8061
rect 7299 7659 7341 7701
rect 7299 7419 7341 7461
rect 6999 7299 7041 7341
rect 7179 7296 7221 7338
rect 7299 7296 7341 7338
rect 6999 7179 7041 7221
rect 6939 7119 6981 7161
rect 7059 6999 7101 7041
rect 6759 6819 6801 6861
rect 6879 6819 6921 6861
rect 7236 6879 7278 6921
rect 7299 6879 7341 6921
rect 7119 6819 7161 6861
rect 6576 6579 6618 6621
rect 6639 6579 6681 6621
rect 6459 6219 6501 6261
rect 6459 6099 6501 6141
rect 6459 5976 6501 6018
rect 6279 5862 6321 5904
rect 6399 5862 6441 5904
rect 6159 5679 6201 5721
rect 6099 5619 6141 5661
rect 6279 5559 6321 5601
rect 6039 5262 6081 5304
rect 6819 6519 6861 6561
rect 6699 6459 6741 6501
rect 6639 6339 6681 6381
rect 6699 6159 6741 6201
rect 6639 6099 6681 6141
rect 6699 5979 6741 6021
rect 7059 6579 7101 6621
rect 6999 6519 7041 6561
rect 6879 6459 6921 6501
rect 7059 6459 7101 6501
rect 6999 6039 7041 6081
rect 6879 5979 6921 6021
rect 6699 5862 6741 5904
rect 6939 5799 6981 5841
rect 6699 5679 6741 5721
rect 6639 5559 6681 5601
rect 6339 5499 6381 5541
rect 6579 5499 6621 5541
rect 6339 5319 6381 5361
rect 6519 5319 6561 5361
rect 6039 5199 6081 5241
rect 6159 5202 6201 5244
rect 6279 5202 6321 5244
rect 5979 5076 6021 5118
rect 6219 5019 6261 5061
rect 6399 5202 6441 5244
rect 6639 5199 6681 5241
rect 6339 5079 6381 5121
rect 5859 4779 5901 4821
rect 6279 4779 6321 4821
rect 5739 4599 5781 4641
rect 5799 4539 5841 4581
rect 6459 5076 6501 5118
rect 6579 5076 6621 5118
rect 6459 4839 6501 4881
rect 6459 4599 6501 4641
rect 6396 4539 6438 4581
rect 5556 4359 5598 4401
rect 5379 4299 5421 4341
rect 5619 4356 5661 4398
rect 5679 4359 5721 4401
rect 5739 4302 5781 4344
rect 5439 4176 5481 4218
rect 6159 4479 6201 4521
rect 6039 4302 6081 4344
rect 6459 4536 6501 4578
rect 6459 4359 6501 4401
rect 6519 4302 6561 4344
rect 6999 5559 7041 5601
rect 6939 5319 6981 5361
rect 6879 5202 6921 5244
rect 6699 4899 6741 4941
rect 6939 5076 6981 5118
rect 6819 4959 6861 5001
rect 6879 4899 6921 4941
rect 6939 4779 6981 4821
rect 6879 4659 6921 4701
rect 6639 4479 6681 4521
rect 6759 4479 6801 4521
rect 6819 4302 6861 4344
rect 5799 4179 5841 4221
rect 5559 4119 5601 4161
rect 5739 4119 5781 4161
rect 5439 4059 5481 4101
rect 6099 4176 6141 4218
rect 6279 4176 6321 4218
rect 5979 4059 6021 4101
rect 5439 3939 5481 3981
rect 5919 3939 5961 3981
rect 5319 3879 5361 3921
rect 5559 3759 5601 3801
rect 5079 3699 5121 3741
rect 5199 3642 5241 3684
rect 5379 3639 5421 3681
rect 5559 3642 5601 3684
rect 5739 3639 5781 3681
rect 6159 3699 6201 3741
rect 6039 3639 6081 3681
rect 6639 4179 6681 4221
rect 6339 4059 6381 4101
rect 6459 4059 6501 4101
rect 6339 3939 6381 3981
rect 6459 3879 6501 3921
rect 6459 3759 6501 3801
rect 6339 3699 6381 3741
rect 5079 3039 5121 3081
rect 4959 2799 5001 2841
rect 4899 2742 4941 2784
rect 5139 2979 5181 3021
rect 5379 3516 5421 3558
rect 5499 3516 5541 3558
rect 5259 2859 5301 2901
rect 5139 2742 5181 2784
rect 5259 2742 5301 2784
rect 5559 3279 5601 3321
rect 4179 2499 4221 2541
rect 4059 2082 4101 2124
rect 4179 2082 4221 2124
rect 4539 2616 4581 2658
rect 4719 2616 4761 2658
rect 4959 2616 5001 2658
rect 5079 2616 5121 2658
rect 5199 2616 5241 2658
rect 5199 2439 5241 2481
rect 4539 2379 4581 2421
rect 4419 2079 4461 2121
rect 4959 2319 5001 2361
rect 4659 2082 4701 2124
rect 4959 2082 5001 2124
rect 3759 1956 3801 1998
rect 3879 1956 3921 1998
rect 4119 1956 4161 1998
rect 4239 1959 4281 2001
rect 3639 1899 3681 1941
rect 3459 1839 3501 1881
rect 3639 1599 3681 1641
rect 2979 1539 3021 1581
rect 3279 1539 3321 1581
rect 3399 1539 3441 1581
rect 2859 1479 2901 1521
rect 2679 1359 2721 1401
rect 2799 1359 2841 1401
rect 2019 1059 2061 1101
rect 1959 999 2001 1041
rect 2139 999 2181 1041
rect 2019 939 2061 981
rect 1839 879 1881 921
rect 1959 819 2001 861
rect 1779 639 1821 681
rect 2199 759 2241 801
rect 2379 1059 2421 1101
rect 2499 1056 2541 1098
rect 3099 1479 3141 1521
rect 2439 939 2481 981
rect 2259 639 2301 681
rect 2859 1059 2901 1101
rect 3039 1056 3081 1098
rect 2799 939 2841 981
rect 2739 819 2781 861
rect 2499 759 2541 801
rect 2679 759 2721 801
rect 1779 396 1821 438
rect 1899 396 1941 438
rect 1539 339 1581 381
rect 1677 339 1719 381
rect 2199 219 2241 261
rect 939 159 981 201
rect 2439 579 2481 621
rect 2379 522 2421 564
rect 2619 639 2661 681
rect 2619 519 2661 561
rect 2439 396 2481 438
rect 2559 396 2601 438
rect 2739 459 2781 501
rect 2979 759 3021 801
rect 3159 759 3201 801
rect 3519 1479 3561 1521
rect 3519 1359 3561 1401
rect 3339 1179 3381 1221
rect 4119 1479 4161 1521
rect 3819 1359 3861 1401
rect 3639 1179 3681 1221
rect 3939 1182 3981 1224
rect 3339 1059 3381 1101
rect 3459 1056 3501 1098
rect 3579 1056 3621 1098
rect 3759 1056 3801 1098
rect 3339 939 3381 981
rect 3819 939 3861 981
rect 3699 819 3741 861
rect 3279 699 3321 741
rect 3519 699 3561 741
rect 2979 522 3021 564
rect 3339 522 3381 564
rect 3459 519 3501 561
rect 2799 399 2841 441
rect 2919 396 2961 438
rect 3159 396 3201 438
rect 5499 2616 5541 2658
rect 5319 2319 5361 2361
rect 5439 2319 5481 2361
rect 5439 2199 5481 2241
rect 5739 3219 5781 3261
rect 5739 3099 5781 3141
rect 5679 2919 5721 2961
rect 5799 2799 5841 2841
rect 6099 3519 6141 3561
rect 6759 4176 6801 4218
rect 6639 4116 6681 4158
rect 6999 4659 7041 4701
rect 7119 6279 7161 6321
rect 7599 8619 7641 8661
rect 7539 8439 7581 8481
rect 7899 9339 7941 9381
rect 7899 9159 7941 9201
rect 8019 9999 8061 10041
rect 8379 11319 8421 11361
rect 8919 11976 8961 12018
rect 9639 14319 9681 14361
rect 9879 14919 9921 14961
rect 9879 14799 9921 14841
rect 9939 14679 9981 14721
rect 9939 14562 9981 14604
rect 9879 14436 9921 14478
rect 9879 14259 9921 14301
rect 9819 14079 9861 14121
rect 9819 13959 9861 14001
rect 9759 13899 9801 13941
rect 9699 13659 9741 13701
rect 9519 13479 9561 13521
rect 10239 15996 10281 16038
rect 10299 15939 10341 15981
rect 10179 15579 10221 15621
rect 10479 15996 10521 16038
rect 10719 15996 10761 16038
rect 10839 15996 10881 16038
rect 10359 15759 10401 15801
rect 10839 15879 10881 15921
rect 10479 15699 10521 15741
rect 10539 15579 10581 15621
rect 10299 15459 10341 15501
rect 10179 15219 10221 15261
rect 10419 15222 10461 15264
rect 10599 15519 10641 15561
rect 10899 15519 10941 15561
rect 10659 15399 10701 15441
rect 10779 15399 10821 15441
rect 10659 15279 10701 15321
rect 10779 15222 10821 15264
rect 11019 16479 11061 16521
rect 10179 14859 10221 14901
rect 10479 15096 10521 15138
rect 10599 15099 10641 15141
rect 10479 14979 10521 15021
rect 10419 14919 10461 14961
rect 10419 14799 10461 14841
rect 10179 14739 10221 14781
rect 10359 14739 10401 14781
rect 10299 14679 10341 14721
rect 10839 15096 10881 15138
rect 10899 15039 10941 15081
rect 10659 14919 10701 14961
rect 10779 14919 10821 14961
rect 10659 14562 10701 14604
rect 10839 14559 10881 14601
rect 10239 14319 10281 14361
rect 10359 14319 10401 14361
rect 10059 14259 10101 14301
rect 9999 14139 10041 14181
rect 9939 13659 9981 13701
rect 10479 13779 10521 13821
rect 10599 14436 10641 14478
rect 10719 14199 10761 14241
rect 10659 14019 10701 14061
rect 10656 13899 10698 13941
rect 10719 13899 10761 13941
rect 10839 14319 10881 14361
rect 10839 14079 10881 14121
rect 10839 13659 10881 13701
rect 9939 13419 9981 13461
rect 9639 13239 9681 13281
rect 9879 13239 9921 13281
rect 9879 13119 9921 13161
rect 9819 12759 9861 12801
rect 9579 12699 9621 12741
rect 9759 12579 9801 12621
rect 9759 12339 9801 12381
rect 9519 12108 9561 12150
rect 9699 12108 9741 12150
rect 9339 11679 9381 11721
rect 10239 13179 10281 13221
rect 9999 13119 10041 13161
rect 10359 13119 10401 13161
rect 10119 13002 10161 13044
rect 10239 13002 10281 13044
rect 9939 12279 9981 12321
rect 9879 12219 9921 12261
rect 9999 12219 10041 12261
rect 10059 12159 10101 12201
rect 10119 12102 10161 12144
rect 10659 13419 10701 13461
rect 10839 13419 10881 13461
rect 10719 13299 10761 13341
rect 10599 13119 10641 13161
rect 10479 13002 10521 13044
rect 10779 13179 10821 13221
rect 10719 12999 10761 13041
rect 10359 12699 10401 12741
rect 10659 12876 10701 12918
rect 10719 12819 10761 12861
rect 10719 12579 10761 12621
rect 11379 17379 11421 17421
rect 11559 17319 11601 17361
rect 11379 17259 11421 17301
rect 11559 17139 11601 17181
rect 11379 16782 11421 16824
rect 11499 16779 11541 16821
rect 11319 16419 11361 16461
rect 11199 16359 11241 16401
rect 11139 16122 11181 16164
rect 11259 16122 11301 16164
rect 13119 18699 13161 18741
rect 13299 18699 13341 18741
rect 13059 18639 13101 18681
rect 11679 18459 11721 18501
rect 12039 18459 12081 18501
rect 12879 18459 12921 18501
rect 11676 18342 11718 18384
rect 11739 18342 11781 18384
rect 11859 18342 11901 18384
rect 11979 18342 12021 18384
rect 12099 18342 12141 18384
rect 12279 18342 12321 18384
rect 11679 18219 11721 18261
rect 11799 18216 11841 18258
rect 11919 18159 11961 18201
rect 12039 18159 12081 18201
rect 11919 17799 11961 17841
rect 11739 17556 11781 17598
rect 12396 18339 12438 18381
rect 12459 18342 12501 18384
rect 12579 18342 12621 18384
rect 12699 18342 12741 18384
rect 12399 18159 12441 18201
rect 12759 18216 12801 18258
rect 13119 18579 13161 18621
rect 13179 18459 13221 18501
rect 13059 18342 13101 18384
rect 12699 18159 12741 18201
rect 12639 18099 12681 18141
rect 12459 18039 12501 18081
rect 12879 18159 12921 18201
rect 12819 18099 12861 18141
rect 12579 17979 12621 18021
rect 12699 17979 12741 18021
rect 12579 17859 12621 17901
rect 12099 17799 12141 17841
rect 12399 17799 12441 17841
rect 12999 18039 13041 18081
rect 12996 17976 13038 18018
rect 13059 17979 13101 18021
rect 12759 17739 12801 17781
rect 12879 17739 12921 17781
rect 12279 17682 12321 17724
rect 12399 17682 12441 17724
rect 12639 17682 12681 17724
rect 12219 17556 12261 17598
rect 11859 17499 11901 17541
rect 12039 17499 12081 17541
rect 11799 17259 11841 17301
rect 11679 17199 11721 17241
rect 11619 16779 11661 16821
rect 12219 17439 12261 17481
rect 12516 17559 12558 17601
rect 12579 17556 12621 17598
rect 12819 17559 12861 17601
rect 13179 18099 13221 18141
rect 13119 17739 13161 17781
rect 14799 18639 14841 18681
rect 14379 18459 14421 18501
rect 13479 18342 13521 18384
rect 13659 18339 13701 18381
rect 14499 18342 14541 18384
rect 14679 18342 14721 18384
rect 13359 18216 13401 18258
rect 13539 18216 13581 18258
rect 13659 18216 13701 18258
rect 13299 17979 13341 18021
rect 13476 18099 13518 18141
rect 13539 18099 13581 18141
rect 13419 17919 13461 17961
rect 13359 17859 13401 17901
rect 13299 17739 13341 17781
rect 13479 17799 13521 17841
rect 13599 17799 13641 17841
rect 13719 18099 13761 18141
rect 13899 17919 13941 17961
rect 13839 17799 13881 17841
rect 13839 17679 13881 17721
rect 12999 17556 13041 17598
rect 13119 17556 13161 17598
rect 13419 17556 13461 17598
rect 13539 17556 13581 17598
rect 12339 17379 12381 17421
rect 12819 17379 12861 17421
rect 13119 17379 13161 17421
rect 12159 17319 12201 17361
rect 12099 17259 12141 17301
rect 11859 17079 11901 17121
rect 11979 17079 12021 17121
rect 11799 17019 11841 17061
rect 11799 16782 11841 16824
rect 11556 16659 11598 16701
rect 11619 16659 11661 16701
rect 11559 16539 11601 16581
rect 11436 16119 11478 16161
rect 11499 16119 11541 16161
rect 11619 16479 11661 16521
rect 11859 16659 11901 16701
rect 12039 16959 12081 17001
rect 12099 16899 12141 16941
rect 12039 16779 12081 16821
rect 12699 17139 12741 17181
rect 12279 16782 12321 16824
rect 12399 16782 12441 16824
rect 12579 16782 12621 16824
rect 13119 16899 13161 16941
rect 12819 16782 12861 16824
rect 12939 16782 12981 16824
rect 13059 16782 13101 16824
rect 12039 16659 12081 16701
rect 11979 16539 12021 16581
rect 11739 16419 11781 16461
rect 11679 16359 11721 16401
rect 11799 16299 11841 16341
rect 11919 16299 11961 16341
rect 12099 16539 12141 16581
rect 12219 16539 12261 16581
rect 12519 16599 12561 16641
rect 12759 16599 12801 16641
rect 12459 16419 12501 16461
rect 12639 16419 12681 16461
rect 12219 16299 12261 16341
rect 11799 16119 11841 16161
rect 11199 15759 11241 15801
rect 11139 15699 11181 15741
rect 11736 15996 11778 16038
rect 11799 15996 11841 16038
rect 11439 15879 11481 15921
rect 11319 15639 11361 15681
rect 11139 15459 11181 15501
rect 11439 15459 11481 15501
rect 11079 15339 11121 15381
rect 11319 15339 11361 15381
rect 11019 15039 11061 15081
rect 10959 14919 11001 14961
rect 11199 15222 11241 15264
rect 11499 15339 11541 15381
rect 11139 15099 11181 15141
rect 11139 14979 11181 15021
rect 11259 14919 11301 14961
rect 11079 14619 11121 14661
rect 10959 14559 11001 14601
rect 11139 14562 11181 14604
rect 11739 15759 11781 15801
rect 11619 15699 11661 15741
rect 11799 15699 11841 15741
rect 12039 15996 12081 16038
rect 12279 16239 12321 16281
rect 11979 15879 12021 15921
rect 12219 15879 12261 15921
rect 11919 15819 11961 15861
rect 11919 15699 11961 15741
rect 11679 15399 11721 15441
rect 11619 15219 11661 15261
rect 11859 15519 11901 15561
rect 11859 15339 11901 15381
rect 11799 15219 11841 15261
rect 11559 15039 11601 15081
rect 11676 15039 11718 15081
rect 11739 15039 11781 15081
rect 11379 14979 11421 15021
rect 11439 14919 11481 14961
rect 11319 14799 11361 14841
rect 11439 14799 11481 14841
rect 11379 14739 11421 14781
rect 11259 14559 11301 14601
rect 11499 14562 11541 14604
rect 10959 14319 11001 14361
rect 11199 14436 11241 14478
rect 11439 14436 11481 14478
rect 11379 14379 11421 14421
rect 11319 14139 11361 14181
rect 11079 14079 11121 14121
rect 10959 14019 11001 14061
rect 10899 13059 10941 13101
rect 11079 14016 11121 14058
rect 11199 13662 11241 13704
rect 11319 13539 11361 13581
rect 11139 13299 11181 13341
rect 11139 13179 11181 13221
rect 10839 12759 10881 12801
rect 11079 13002 11121 13044
rect 11199 13008 11241 13050
rect 10959 12879 11001 12921
rect 11139 12879 11181 12921
rect 11016 12759 11058 12801
rect 11079 12759 11121 12801
rect 10959 12579 11001 12621
rect 10899 12519 10941 12561
rect 10779 12399 10821 12441
rect 10959 12399 11001 12441
rect 10539 12339 10581 12381
rect 10479 12279 10521 12321
rect 9879 12039 9921 12081
rect 9459 11979 9501 12021
rect 9099 11559 9141 11601
rect 9219 11559 9261 11601
rect 9399 11559 9441 11601
rect 8979 11499 9021 11541
rect 9159 11499 9201 11541
rect 8859 11439 8901 11481
rect 8499 11316 8541 11358
rect 8559 11259 8601 11301
rect 8379 11079 8421 11121
rect 8199 10899 8241 10941
rect 8799 11316 8841 11358
rect 8919 11316 8961 11358
rect 9039 11316 9081 11358
rect 8679 11259 8721 11301
rect 8979 11079 9021 11121
rect 8679 11019 8721 11061
rect 8739 10959 8781 11001
rect 8619 10839 8661 10881
rect 8559 10719 8601 10761
rect 8259 10599 8301 10641
rect 8559 10539 8601 10581
rect 8619 10599 8661 10641
rect 9099 11019 9141 11061
rect 9039 10719 9081 10761
rect 8859 10542 8901 10584
rect 8979 10542 9021 10584
rect 8499 10479 8541 10521
rect 8439 10299 8481 10341
rect 8319 10239 8361 10281
rect 8199 10119 8241 10161
rect 8139 10059 8181 10101
rect 8079 9939 8121 9981
rect 8319 10059 8361 10101
rect 8259 9939 8301 9981
rect 8199 9879 8241 9921
rect 8019 9759 8061 9801
rect 8199 9759 8241 9801
rect 8139 9639 8181 9681
rect 8079 9579 8121 9621
rect 8019 9339 8061 9381
rect 7959 9039 8001 9081
rect 8079 9099 8121 9141
rect 7839 8799 7881 8841
rect 7659 8439 7701 8481
rect 8079 8859 8121 8901
rect 8679 10416 8721 10458
rect 8919 10359 8961 10401
rect 8799 10179 8841 10221
rect 8679 10119 8721 10161
rect 8499 10059 8541 10101
rect 8439 9939 8481 9981
rect 8619 9939 8661 9981
rect 8499 9882 8541 9924
rect 8439 9756 8481 9798
rect 8559 9756 8601 9798
rect 8979 10299 9021 10341
rect 9039 10119 9081 10161
rect 9159 10899 9201 10941
rect 9279 11439 9321 11481
rect 10059 11976 10101 12018
rect 10179 11979 10221 12021
rect 10539 12099 10581 12141
rect 10659 12108 10701 12150
rect 10839 12108 10881 12150
rect 9879 11859 9921 11901
rect 10299 11970 10341 12012
rect 10479 11970 10521 12012
rect 10239 11859 10281 11901
rect 9879 11739 9921 11781
rect 10179 11739 10221 11781
rect 9579 11679 9621 11721
rect 9639 11619 9681 11661
rect 9579 11559 9621 11601
rect 9639 11439 9681 11481
rect 9519 11316 9561 11358
rect 9279 11259 9321 11301
rect 9639 11259 9681 11301
rect 9519 11199 9561 11241
rect 9579 11079 9621 11121
rect 9519 10899 9561 10941
rect 9516 10779 9558 10821
rect 9579 10779 9621 10821
rect 10479 11799 10521 11841
rect 10899 11979 10941 12021
rect 10899 11859 10941 11901
rect 10299 11739 10341 11781
rect 10539 11739 10581 11781
rect 10239 11679 10281 11721
rect 9939 11499 9981 11541
rect 10359 11679 10401 11721
rect 10839 11679 10881 11721
rect 10299 11439 10341 11481
rect 9939 11319 9981 11361
rect 10056 11310 10098 11352
rect 10119 11319 10161 11361
rect 10419 11619 10461 11661
rect 9939 11199 9981 11241
rect 10239 11310 10281 11352
rect 10359 11310 10401 11352
rect 10479 11499 10521 11541
rect 10539 11442 10581 11484
rect 10479 11319 10521 11361
rect 10419 11259 10461 11301
rect 10059 11019 10101 11061
rect 9819 10959 9861 11001
rect 9939 10959 9981 11001
rect 9759 10899 9801 10941
rect 9699 10779 9741 10821
rect 9219 10659 9261 10701
rect 9459 10659 9501 10701
rect 9639 10659 9681 10701
rect 9339 10542 9381 10584
rect 9459 10539 9501 10581
rect 9579 10542 9621 10584
rect 9759 10539 9801 10581
rect 8739 9999 8781 10041
rect 8919 9999 8961 10041
rect 9219 9999 9261 10041
rect 8319 9699 8361 9741
rect 8679 9699 8721 9741
rect 8619 9639 8661 9681
rect 8559 9579 8601 9621
rect 8319 9459 8361 9501
rect 8439 9459 8481 9501
rect 8259 9279 8301 9321
rect 8499 9339 8541 9381
rect 8499 9219 8541 9261
rect 8199 8979 8241 9021
rect 8319 8982 8361 9024
rect 8439 8979 8481 9021
rect 8139 8739 8181 8781
rect 7959 8559 8001 8601
rect 8199 8499 8241 8541
rect 8199 8379 8241 8421
rect 7839 8319 7881 8361
rect 8079 8322 8121 8364
rect 7539 8139 7581 8181
rect 7479 8019 7521 8061
rect 7599 8079 7641 8121
rect 7659 8019 7701 8061
rect 7899 8259 7941 8301
rect 8019 8196 8061 8238
rect 8139 8196 8181 8238
rect 8499 8859 8541 8901
rect 8379 8739 8421 8781
rect 8379 8676 8421 8718
rect 8679 9519 8721 9561
rect 8619 9339 8661 9381
rect 8919 9882 8961 9924
rect 8859 9756 8901 9798
rect 8799 9639 8841 9681
rect 8799 9459 8841 9501
rect 8739 9159 8781 9201
rect 8679 9099 8721 9141
rect 9039 9639 9081 9681
rect 8979 9219 9021 9261
rect 8919 9039 8961 9081
rect 8979 8979 9021 9021
rect 8619 8859 8661 8901
rect 8559 8679 8601 8721
rect 8739 8856 8781 8898
rect 9456 10419 9498 10461
rect 9519 10419 9561 10461
rect 9459 10299 9501 10341
rect 9399 10239 9441 10281
rect 9339 10179 9381 10221
rect 9279 9939 9321 9981
rect 9399 9999 9441 10041
rect 9399 9756 9441 9798
rect 9279 9639 9321 9681
rect 9099 9579 9141 9621
rect 9399 9519 9441 9561
rect 9099 9399 9141 9441
rect 9219 9399 9261 9441
rect 9159 9339 9201 9381
rect 9099 9159 9141 9201
rect 9579 10359 9621 10401
rect 9759 10419 9801 10461
rect 9639 10299 9681 10341
rect 10719 11199 10761 11241
rect 11019 12339 11061 12381
rect 11319 12579 11361 12621
rect 11139 12459 11181 12501
rect 11079 12099 11121 12141
rect 11619 14439 11661 14481
rect 11559 14319 11601 14361
rect 11439 13839 11481 13881
rect 11619 13779 11661 13821
rect 11799 14739 11841 14781
rect 11739 14679 11781 14721
rect 12099 15639 12141 15681
rect 12099 15519 12141 15561
rect 12039 15459 12081 15501
rect 12039 15339 12081 15381
rect 12156 15339 12198 15381
rect 12219 15339 12261 15381
rect 12579 16122 12621 16164
rect 12999 16656 13041 16698
rect 13119 16539 13161 16581
rect 13239 17439 13281 17481
rect 13779 17556 13821 17598
rect 13899 17556 13941 17598
rect 13779 17079 13821 17121
rect 13239 17019 13281 17061
rect 13659 17019 13701 17061
rect 13179 16299 13221 16341
rect 13539 16899 13581 16941
rect 13299 16782 13341 16824
rect 13419 16782 13461 16824
rect 13899 16782 13941 16824
rect 14019 18099 14061 18141
rect 14439 18216 14481 18258
rect 15579 18759 15621 18801
rect 15219 18699 15261 18741
rect 15339 18699 15381 18741
rect 14859 18579 14901 18621
rect 14919 18459 14961 18501
rect 15039 18399 15081 18441
rect 14799 18099 14841 18141
rect 14379 17979 14421 18021
rect 14559 17979 14601 18021
rect 14679 17979 14721 18021
rect 14199 17919 14241 17961
rect 14139 17859 14181 17901
rect 14019 17679 14061 17721
rect 14319 17859 14361 17901
rect 14259 17679 14301 17721
rect 15099 18216 15141 18258
rect 14979 17919 15021 17961
rect 14499 17799 14541 17841
rect 14739 17799 14781 17841
rect 14379 17679 14421 17721
rect 14619 17682 14661 17724
rect 14079 17556 14121 17598
rect 14199 17556 14241 17598
rect 14319 17556 14361 17598
rect 14439 17556 14481 17598
rect 14559 17556 14601 17598
rect 14439 17439 14481 17481
rect 14439 17199 14481 17241
rect 14199 17139 14241 17181
rect 14079 16899 14121 16941
rect 13299 16539 13341 16581
rect 13479 16656 13521 16698
rect 13959 16659 14001 16701
rect 13839 16599 13881 16641
rect 13779 16539 13821 16581
rect 13899 16539 13941 16581
rect 13359 16479 13401 16521
rect 13599 16479 13641 16521
rect 13599 16299 13641 16341
rect 13239 16239 13281 16281
rect 13899 16419 13941 16461
rect 14559 17079 14601 17121
rect 14439 17019 14481 17061
rect 14319 16782 14361 16824
rect 14499 16899 14541 16941
rect 14079 16479 14121 16521
rect 14019 16419 14061 16461
rect 13839 16239 13881 16281
rect 13299 16122 13341 16164
rect 13479 16119 13521 16161
rect 13659 16122 13701 16164
rect 13779 16122 13821 16164
rect 12336 15999 12378 16041
rect 12399 15996 12441 16038
rect 12519 15996 12561 16038
rect 12759 15999 12801 16041
rect 12639 15879 12681 15921
rect 12939 15996 12981 16038
rect 13119 15999 13161 16041
rect 12879 15939 12921 15981
rect 13059 15879 13101 15921
rect 12699 15759 12741 15801
rect 12459 15639 12501 15681
rect 12519 15579 12561 15621
rect 12399 15459 12441 15501
rect 12339 15399 12381 15441
rect 12459 15399 12501 15441
rect 12279 15279 12321 15321
rect 12399 15279 12441 15321
rect 12339 15222 12381 15264
rect 12039 15099 12081 15141
rect 12039 14919 12081 14961
rect 12219 15039 12261 15081
rect 11979 14739 12021 14781
rect 12159 14739 12201 14781
rect 11919 14619 11961 14661
rect 12099 14619 12141 14661
rect 11979 14562 12021 14604
rect 12399 15099 12441 15141
rect 12339 14979 12381 15021
rect 12279 14919 12321 14961
rect 12399 14799 12441 14841
rect 12339 14739 12381 14781
rect 12579 15456 12621 15498
rect 12999 15699 13041 15741
rect 12879 15579 12921 15621
rect 12999 15579 13041 15621
rect 12759 15519 12801 15561
rect 12699 15279 12741 15321
rect 13479 15996 13521 16038
rect 13599 15996 13641 16038
rect 13359 15879 13401 15921
rect 13239 15819 13281 15861
rect 13119 15639 13161 15681
rect 13419 15759 13461 15801
rect 13359 15639 13401 15681
rect 13239 15399 13281 15441
rect 13239 15279 13281 15321
rect 12699 15096 12741 15138
rect 12639 14979 12681 15021
rect 12579 14859 12621 14901
rect 12579 14739 12621 14781
rect 12519 14679 12561 14721
rect 12579 14619 12621 14661
rect 12219 14562 12261 14604
rect 12399 14562 12441 14604
rect 12579 14556 12621 14598
rect 12939 15099 12981 15141
rect 12819 14919 12861 14961
rect 12699 14859 12741 14901
rect 12939 14859 12981 14901
rect 12639 14499 12681 14541
rect 11919 14436 11961 14478
rect 12039 14436 12081 14478
rect 12219 14439 12261 14481
rect 11859 14259 11901 14301
rect 11799 14139 11841 14181
rect 11739 14019 11781 14061
rect 11439 13662 11481 13704
rect 11379 12459 11421 12501
rect 11259 12219 11301 12261
rect 11199 11976 11241 12018
rect 11499 13539 11541 13581
rect 11559 13419 11601 13461
rect 11679 13419 11721 13461
rect 11979 14079 12021 14121
rect 11979 13959 12021 14001
rect 12219 14319 12261 14361
rect 12159 14139 12201 14181
rect 12039 13662 12081 13704
rect 11799 13359 11841 13401
rect 11979 13479 12021 13521
rect 11919 13239 11961 13281
rect 11859 13179 11901 13221
rect 11859 13059 11901 13101
rect 11499 12999 11541 13041
rect 11499 12879 11541 12921
rect 11619 12879 11661 12921
rect 11439 12339 11481 12381
rect 11739 12759 11781 12801
rect 11019 11679 11061 11721
rect 10959 11499 11001 11541
rect 11199 11499 11241 11541
rect 11019 11442 11061 11484
rect 10959 11259 11001 11301
rect 9999 10839 10041 10881
rect 10119 10839 10161 10881
rect 10479 10839 10521 10881
rect 10599 10839 10641 10881
rect 10839 10839 10881 10881
rect 11079 11079 11121 11121
rect 10959 10779 11001 10821
rect 10719 10659 10761 10701
rect 9999 10542 10041 10584
rect 10119 10542 10161 10584
rect 10299 10542 10341 10584
rect 10479 10542 10521 10584
rect 10599 10542 10641 10584
rect 9879 10419 9921 10461
rect 9819 10359 9861 10401
rect 9759 10239 9801 10281
rect 9579 10179 9621 10221
rect 9939 10359 9981 10401
rect 9759 10119 9801 10161
rect 9879 10119 9921 10161
rect 9639 9999 9681 10041
rect 9579 9939 9621 9981
rect 9399 9279 9441 9321
rect 9519 9279 9561 9321
rect 9879 9882 9921 9924
rect 9639 9756 9681 9798
rect 9819 9756 9861 9798
rect 9699 9699 9741 9741
rect 9879 9699 9921 9741
rect 9819 9579 9861 9621
rect 9759 9519 9801 9561
rect 9759 9339 9801 9381
rect 9699 9159 9741 9201
rect 9516 9099 9558 9141
rect 9579 9099 9621 9141
rect 9279 8982 9321 9024
rect 9459 8982 9501 9024
rect 9099 8859 9141 8901
rect 9039 8739 9081 8781
rect 8859 8619 8901 8661
rect 8619 8559 8661 8601
rect 8679 8439 8721 8481
rect 8919 8439 8961 8481
rect 8499 8322 8541 8364
rect 8739 8319 8781 8361
rect 9039 8322 9081 8364
rect 8319 8196 8361 8238
rect 7719 7959 7761 8001
rect 7779 7899 7821 7941
rect 7659 7839 7701 7881
rect 7539 7599 7581 7641
rect 7539 7536 7581 7578
rect 7419 7419 7461 7461
rect 7599 7296 7641 7338
rect 7479 7119 7521 7161
rect 7899 8019 7941 8061
rect 8259 8079 8301 8121
rect 8079 7959 8121 8001
rect 8139 7899 8181 7941
rect 8079 7839 8121 7881
rect 8079 7719 8121 7761
rect 8019 7659 8061 7701
rect 8139 7539 8181 7581
rect 7899 7479 7941 7521
rect 7839 7422 7881 7464
rect 8019 7422 8061 7464
rect 8139 7419 8181 7461
rect 7479 7056 7521 7098
rect 7779 7059 7821 7101
rect 7959 7059 8001 7101
rect 7419 6939 7461 6981
rect 8019 6999 8061 7041
rect 7779 6939 7821 6981
rect 7299 6699 7341 6741
rect 7239 6459 7281 6501
rect 7299 6399 7341 6441
rect 7239 6339 7281 6381
rect 7419 6339 7461 6381
rect 7539 6339 7581 6381
rect 7179 5979 7221 6021
rect 7659 6579 7701 6621
rect 7659 6279 7701 6321
rect 7599 6219 7641 6261
rect 7359 6159 7401 6201
rect 7539 6159 7581 6201
rect 7299 6099 7341 6141
rect 7359 6039 7401 6081
rect 7299 5979 7341 6021
rect 7599 5979 7641 6021
rect 8139 7179 8181 7221
rect 8139 6879 8181 6921
rect 8139 6699 8181 6741
rect 7899 6636 7941 6678
rect 7899 6519 7941 6561
rect 8259 7479 8301 7521
rect 8559 8196 8601 8238
rect 8679 8199 8721 8241
rect 8439 8079 8481 8121
rect 8379 7959 8421 8001
rect 8979 8196 9021 8238
rect 8739 8079 8781 8121
rect 8859 8079 8901 8121
rect 8679 7959 8721 8001
rect 8559 7779 8601 7821
rect 8379 7719 8421 7761
rect 8559 7659 8601 7701
rect 8499 7539 8541 7581
rect 8919 8019 8961 8061
rect 8859 7959 8901 8001
rect 8799 7719 8841 7761
rect 8679 7419 8721 7461
rect 9219 8856 9261 8898
rect 9579 8982 9621 9024
rect 9699 8982 9741 9024
rect 9939 9459 9981 9501
rect 10179 10419 10221 10461
rect 11739 12219 11781 12261
rect 11499 12102 11541 12144
rect 11619 12102 11661 12144
rect 12039 13419 12081 13461
rect 12039 13299 12081 13341
rect 12159 13239 12201 13281
rect 12459 14436 12501 14478
rect 12579 14439 12621 14481
rect 12339 14379 12381 14421
rect 12519 14379 12561 14421
rect 12279 13959 12321 14001
rect 12459 13839 12501 13881
rect 12339 13662 12381 13704
rect 12579 14139 12621 14181
rect 12879 14799 12921 14841
rect 13059 15099 13101 15141
rect 12939 14436 12981 14478
rect 12999 14319 13041 14361
rect 12699 14199 12741 14241
rect 12819 14199 12861 14241
rect 12639 14079 12681 14121
rect 12579 13959 12621 14001
rect 12519 13659 12561 13701
rect 13119 14919 13161 14961
rect 13299 15039 13341 15081
rect 13179 14679 13221 14721
rect 13359 14919 13401 14961
rect 13479 15699 13521 15741
rect 13539 15579 13581 15621
rect 13659 15519 13701 15561
rect 13719 15459 13761 15501
rect 13659 15339 13701 15381
rect 13476 15219 13518 15261
rect 13539 15222 13581 15264
rect 13719 15222 13761 15264
rect 13479 15099 13521 15141
rect 13599 15099 13641 15141
rect 13419 14619 13461 14661
rect 13299 14562 13341 14604
rect 13539 14619 13581 14661
rect 13479 14559 13521 14601
rect 13239 14436 13281 14478
rect 13359 14439 13401 14481
rect 13359 14319 13401 14361
rect 13659 14859 13701 14901
rect 14139 16299 14181 16341
rect 14439 16659 14481 16701
rect 14316 16479 14358 16521
rect 14379 16479 14421 16521
rect 14319 16359 14361 16401
rect 14499 16539 14541 16581
rect 14859 17739 14901 17781
rect 14799 17679 14841 17721
rect 15099 17682 15141 17724
rect 15039 17559 15081 17601
rect 14859 17199 14901 17241
rect 14799 17019 14841 17061
rect 14559 16479 14601 16521
rect 14739 16779 14781 16821
rect 14556 16359 14598 16401
rect 14619 16359 14661 16401
rect 14259 16239 14301 16281
rect 14496 16239 14538 16281
rect 14559 16239 14601 16281
rect 13959 15996 14001 16038
rect 14139 15939 14181 15981
rect 13959 15639 14001 15681
rect 13899 15459 13941 15501
rect 14379 16122 14421 16164
rect 14619 16122 14661 16164
rect 14259 15939 14301 15981
rect 14379 15939 14421 15981
rect 14199 15639 14241 15681
rect 14319 15519 14361 15561
rect 14079 15222 14121 15264
rect 13899 15039 13941 15081
rect 13839 14799 13881 14841
rect 13899 14739 13941 14781
rect 14139 15096 14181 15138
rect 14619 15879 14661 15921
rect 14799 16656 14841 16698
rect 14739 16419 14781 16461
rect 14679 15759 14721 15801
rect 15399 18342 15441 18384
rect 15339 18216 15381 18258
rect 15279 18159 15321 18201
rect 15339 18099 15381 18141
rect 15519 18219 15561 18261
rect 16959 18699 17001 18741
rect 15999 18579 16041 18621
rect 15819 18459 15861 18501
rect 15639 18399 15681 18441
rect 15639 18219 15681 18261
rect 15879 18219 15921 18261
rect 15579 18159 15621 18201
rect 15639 18099 15681 18141
rect 15459 18039 15501 18081
rect 15639 17979 15681 18021
rect 15339 17859 15381 17901
rect 15339 17679 15381 17721
rect 15459 17682 15501 17724
rect 15759 17799 15801 17841
rect 15639 17679 15681 17721
rect 15939 17682 15981 17724
rect 15399 17556 15441 17598
rect 15279 17499 15321 17541
rect 15519 17499 15561 17541
rect 15339 17319 15381 17361
rect 15459 17319 15501 17361
rect 15279 17259 15321 17301
rect 15219 17019 15261 17061
rect 15159 16839 15201 16881
rect 15459 17199 15501 17241
rect 15399 17079 15441 17121
rect 15339 16899 15381 16941
rect 15459 16959 15501 17001
rect 15459 16779 15501 16821
rect 15219 16656 15261 16698
rect 15339 16656 15381 16698
rect 15099 16539 15141 16581
rect 15039 16479 15081 16521
rect 14859 16122 14901 16164
rect 15039 16239 15081 16281
rect 15219 16359 15261 16401
rect 14979 16119 15021 16161
rect 14979 15999 15021 16041
rect 14919 15939 14961 15981
rect 14919 15759 14961 15801
rect 14919 15639 14961 15681
rect 14739 15579 14781 15621
rect 15039 15939 15081 15981
rect 14799 15459 14841 15501
rect 14979 15459 15021 15501
rect 14499 15339 14541 15381
rect 14439 15279 14481 15321
rect 14739 15279 14781 15321
rect 14619 15222 14661 15264
rect 14199 15039 14241 15081
rect 14319 15039 14361 15081
rect 14019 14919 14061 14961
rect 13659 14679 13701 14721
rect 13959 14679 14001 14721
rect 13659 14562 13701 14604
rect 13779 14562 13821 14604
rect 13599 14439 13641 14481
rect 13659 14379 13701 14421
rect 13119 14259 13161 14301
rect 13239 14259 13281 14301
rect 13599 14259 13641 14301
rect 13059 14079 13101 14121
rect 12999 14019 13041 14061
rect 12999 13899 13041 13941
rect 12819 13839 12861 13881
rect 12759 13662 12801 13704
rect 12879 13662 12921 13704
rect 12579 13536 12621 13578
rect 12699 13536 12741 13578
rect 12396 13479 12438 13521
rect 12459 13479 12501 13521
rect 12219 13059 12261 13101
rect 12159 13002 12201 13044
rect 12279 13002 12321 13044
rect 13119 13536 13161 13578
rect 12639 13419 12681 13461
rect 12876 13419 12918 13461
rect 12939 13419 12981 13461
rect 11979 12876 12021 12918
rect 12099 12876 12141 12918
rect 11919 12759 11961 12801
rect 12039 12459 12081 12501
rect 12399 12879 12441 12921
rect 12279 12759 12321 12801
rect 12219 12339 12261 12381
rect 11919 12219 11961 12261
rect 12039 12219 12081 12261
rect 11859 12099 11901 12141
rect 11499 11979 11541 12021
rect 11559 11919 11601 11961
rect 11499 11799 11541 11841
rect 11256 11439 11298 11481
rect 11319 11439 11361 11481
rect 11439 11439 11481 11481
rect 11679 11739 11721 11781
rect 11799 11739 11841 11781
rect 11619 11559 11661 11601
rect 11559 11439 11601 11481
rect 11379 11316 11421 11358
rect 11559 11319 11601 11361
rect 11259 11199 11301 11241
rect 11079 10599 11121 10641
rect 11199 10599 11241 10641
rect 10899 10542 10941 10584
rect 11259 10542 11301 10584
rect 11379 10539 11421 10581
rect 10119 10359 10161 10401
rect 10299 10239 10341 10281
rect 10179 9999 10221 10041
rect 10299 9939 10341 9981
rect 10239 9882 10281 9924
rect 10419 10416 10461 10458
rect 10419 10179 10461 10221
rect 10479 9939 10521 9981
rect 10419 9879 10461 9921
rect 10119 9579 10161 9621
rect 10299 9756 10341 9798
rect 10479 9756 10521 9798
rect 10719 10416 10761 10458
rect 10959 10416 11001 10458
rect 11079 10416 11121 10458
rect 11319 10419 11361 10461
rect 10719 10299 10761 10341
rect 11199 10299 11241 10341
rect 10659 9939 10701 9981
rect 10839 9939 10881 9981
rect 11079 9939 11121 9981
rect 11199 9939 11241 9981
rect 10719 9756 10761 9798
rect 10839 9759 10881 9801
rect 11379 9999 11421 10041
rect 11799 11442 11841 11484
rect 12159 12159 12201 12201
rect 12219 12099 12261 12141
rect 12099 11976 12141 12018
rect 12399 12579 12441 12621
rect 12339 12219 12381 12261
rect 11979 11919 12021 11961
rect 12279 11919 12321 11961
rect 12219 11559 12261 11601
rect 12039 11448 12081 11490
rect 12579 12879 12621 12921
rect 12579 12519 12621 12561
rect 12519 12339 12561 12381
rect 13119 13299 13161 13341
rect 12699 13239 12741 13281
rect 12879 13119 12921 13161
rect 13179 13059 13221 13101
rect 12759 12699 12801 12741
rect 12699 12459 12741 12501
rect 12699 12339 12741 12381
rect 12939 12339 12981 12381
rect 12639 12159 12681 12201
rect 12399 12099 12441 12141
rect 12579 12102 12621 12144
rect 13059 12279 13101 12321
rect 12759 12102 12801 12144
rect 12399 11979 12441 12021
rect 12339 11499 12381 11541
rect 12639 11976 12681 12018
rect 13119 12219 13161 12261
rect 12639 11739 12681 11781
rect 12519 11679 12561 11721
rect 12639 11676 12681 11718
rect 12459 11448 12501 11490
rect 11979 11379 12021 11421
rect 11679 11319 11721 11361
rect 11679 11019 11721 11061
rect 11859 11316 11901 11358
rect 11679 10899 11721 10941
rect 11619 10599 11661 10641
rect 12039 11079 12081 11121
rect 11799 10539 11841 10581
rect 12039 10479 12081 10521
rect 11499 10239 11541 10281
rect 11859 10410 11901 10452
rect 12639 11319 12681 11361
rect 12639 11256 12681 11298
rect 12279 11139 12321 11181
rect 12159 11019 12201 11061
rect 12459 10959 12501 11001
rect 12219 10599 12261 10641
rect 12519 10719 12561 10761
rect 12099 10359 12141 10401
rect 12219 10359 12261 10401
rect 12159 10239 12201 10281
rect 11739 10179 11781 10221
rect 11979 10059 12021 10101
rect 11619 9999 11661 10041
rect 11019 9756 11061 9798
rect 10959 9699 11001 9741
rect 10539 9639 10581 9681
rect 10299 9579 10341 9621
rect 10179 9459 10221 9501
rect 9939 9039 9981 9081
rect 10059 9039 10101 9081
rect 9459 8799 9501 8841
rect 9219 8739 9261 8781
rect 9339 8739 9381 8781
rect 9159 7719 9201 7761
rect 9639 8856 9681 8898
rect 9759 8856 9801 8898
rect 9879 8859 9921 8901
rect 9699 8799 9741 8841
rect 9519 8679 9561 8721
rect 9519 8499 9561 8541
rect 9699 8196 9741 8238
rect 9879 8679 9921 8721
rect 10119 8982 10161 9024
rect 10059 8559 10101 8601
rect 10179 8559 10221 8601
rect 9939 8379 9981 8421
rect 10059 8322 10101 8364
rect 10239 8379 10281 8421
rect 10179 8319 10221 8361
rect 9279 7959 9321 8001
rect 9339 7779 9381 7821
rect 9219 7539 9261 7581
rect 8799 7359 8841 7401
rect 8259 7293 8301 7335
rect 8376 7293 8418 7335
rect 8439 7299 8481 7341
rect 8739 7239 8781 7281
rect 8559 7119 8601 7161
rect 8499 7059 8541 7101
rect 8499 6939 8541 6981
rect 8439 6879 8481 6921
rect 8679 6762 8721 6804
rect 8799 6762 8841 6804
rect 8259 6639 8301 6681
rect 8739 6636 8781 6678
rect 8199 6579 8241 6621
rect 8319 6579 8361 6621
rect 7839 6459 7881 6501
rect 7416 5859 7458 5901
rect 7539 5862 7581 5904
rect 7779 5919 7821 5961
rect 7719 5862 7761 5904
rect 7299 5736 7341 5778
rect 7479 5736 7521 5778
rect 7179 5679 7221 5721
rect 7359 5559 7401 5601
rect 7659 5559 7701 5601
rect 7119 5499 7161 5541
rect 7176 5439 7218 5481
rect 7239 5439 7281 5481
rect 7239 5319 7281 5361
rect 7179 5259 7221 5301
rect 7479 5379 7521 5421
rect 7119 5076 7161 5118
rect 7419 5079 7461 5121
rect 6819 4059 6861 4101
rect 6939 4059 6981 4101
rect 6636 3699 6678 3741
rect 6699 3699 6741 3741
rect 6516 3639 6558 3681
rect 6579 3642 6621 3684
rect 6939 3879 6981 3921
rect 7239 4599 7281 4641
rect 7119 4302 7161 4344
rect 7299 4539 7341 4581
rect 7299 4419 7341 4461
rect 6879 3639 6921 3681
rect 6339 3516 6381 3558
rect 6459 3516 6501 3558
rect 6639 3516 6681 3558
rect 6759 3516 6801 3558
rect 6879 3516 6921 3558
rect 6219 3459 6261 3501
rect 6099 3219 6141 3261
rect 5979 2859 6021 2901
rect 6279 3099 6321 3141
rect 6219 2979 6261 3021
rect 6099 2742 6141 2784
rect 6579 2979 6621 3021
rect 6459 2919 6501 2961
rect 6399 2859 6441 2901
rect 5739 2616 5781 2658
rect 5859 2616 5901 2658
rect 5979 2616 6021 2658
rect 5859 2439 5901 2481
rect 5796 2319 5838 2361
rect 5859 2319 5901 2361
rect 5739 2259 5781 2301
rect 5499 2139 5541 2181
rect 5259 2079 5301 2121
rect 5379 2082 5421 2124
rect 4719 1956 4761 1998
rect 4479 1899 4521 1941
rect 4419 1839 4461 1881
rect 5019 1956 5061 1998
rect 5199 1959 5241 2001
rect 5319 1959 5361 2001
rect 5259 1899 5301 1941
rect 4899 1839 4941 1881
rect 4479 1779 4521 1821
rect 4959 1719 5001 1761
rect 4839 1659 4881 1701
rect 4239 1359 4281 1401
rect 4719 1299 4761 1341
rect 4179 1239 4221 1281
rect 4419 1182 4461 1224
rect 4239 1119 4281 1161
rect 4179 999 4221 1041
rect 4119 939 4161 981
rect 4479 879 4521 921
rect 4419 759 4461 801
rect 3879 699 3921 741
rect 3999 522 4041 564
rect 4179 522 4221 564
rect 4299 522 4341 564
rect 3639 396 3681 438
rect 3819 339 3861 381
rect 2679 279 2721 321
rect 3639 279 3681 321
rect 3759 276 3801 318
rect 4239 396 4281 438
rect 4419 396 4461 438
rect 4119 339 4161 381
rect 4599 819 4641 861
rect 4539 699 4581 741
rect 5559 1956 5601 1998
rect 5439 1599 5481 1641
rect 5079 1479 5121 1521
rect 4959 1182 5001 1224
rect 5739 2079 5781 2121
rect 5979 2199 6021 2241
rect 6519 2859 6561 2901
rect 6279 2616 6321 2658
rect 6459 2616 6501 2658
rect 6159 2559 6201 2601
rect 6219 2379 6261 2421
rect 6459 2379 6501 2421
rect 5799 1956 5841 1998
rect 5919 1779 5961 1821
rect 5679 1719 5721 1761
rect 6159 2079 6201 2121
rect 6339 2082 6381 2124
rect 6699 2742 6741 2784
rect 7239 4119 7281 4161
rect 6999 3699 7041 3741
rect 7179 3699 7221 3741
rect 6939 3459 6981 3501
rect 7119 3642 7161 3684
rect 7659 5202 7701 5244
rect 8019 6279 8061 6321
rect 8139 6039 8181 6081
rect 8019 5862 8061 5904
rect 8259 6219 8301 6261
rect 8259 5799 8301 5841
rect 7959 5739 8001 5781
rect 9099 7479 9141 7521
rect 8919 7419 8961 7461
rect 9039 7422 9081 7464
rect 8979 7299 9021 7341
rect 8919 7179 8961 7221
rect 8919 7059 8961 7101
rect 9219 7296 9261 7338
rect 9099 7239 9141 7281
rect 9219 7233 9261 7275
rect 8979 6939 9021 6981
rect 9099 6939 9141 6981
rect 8979 6762 9021 6804
rect 9639 7719 9681 7761
rect 9519 7422 9561 7464
rect 9399 7119 9441 7161
rect 9339 7059 9381 7101
rect 9219 6762 9261 6804
rect 9519 6762 9561 6804
rect 8979 6639 9021 6681
rect 9159 6579 9201 6621
rect 9459 6579 9501 6621
rect 9519 6519 9561 6561
rect 8919 6459 8961 6501
rect 8859 6399 8901 6441
rect 8559 5919 8601 5961
rect 8739 5862 8781 5904
rect 8859 5862 8901 5904
rect 9039 5862 9081 5904
rect 9219 5862 9261 5904
rect 7899 5379 7941 5421
rect 7899 5259 7941 5301
rect 8139 5499 8181 5541
rect 8079 5379 8121 5421
rect 8259 5439 8301 5481
rect 8139 5319 8181 5361
rect 7959 5199 8001 5241
rect 8079 5202 8121 5244
rect 7599 5076 7641 5118
rect 7479 4959 7521 5001
rect 7836 5076 7878 5118
rect 7899 5079 7941 5121
rect 8019 5076 8061 5118
rect 8199 5076 8241 5118
rect 8919 5736 8961 5778
rect 8619 5679 8661 5721
rect 8739 5679 8781 5721
rect 8916 5673 8958 5715
rect 8979 5679 9021 5721
rect 8499 5559 8541 5601
rect 8739 5499 8781 5541
rect 8379 5379 8421 5421
rect 8559 5319 8601 5361
rect 8439 5076 8481 5118
rect 8019 4959 8061 5001
rect 7719 4899 7761 4941
rect 7839 4899 7881 4941
rect 7416 4359 7458 4401
rect 7479 4359 7521 4401
rect 7719 4359 7761 4401
rect 7419 4296 7461 4338
rect 7539 4302 7581 4344
rect 7899 4359 7941 4401
rect 8019 4302 8061 4344
rect 7599 4176 7641 4218
rect 7539 4059 7581 4101
rect 7839 4059 7881 4101
rect 7419 3759 7461 3801
rect 6999 3279 7041 3321
rect 6999 3216 7041 3258
rect 6879 2739 6921 2781
rect 7179 3516 7221 3558
rect 7299 3516 7341 3558
rect 7539 3699 7581 3741
rect 7659 3642 7701 3684
rect 8439 4899 8481 4941
rect 8679 5076 8721 5118
rect 8619 4599 8661 4641
rect 8499 4359 8541 4401
rect 8259 4302 8301 4344
rect 8379 4302 8421 4344
rect 8259 4119 8301 4161
rect 8379 4119 8421 4161
rect 8199 4059 8241 4101
rect 8259 3999 8301 4041
rect 8019 3939 8061 3981
rect 7959 3879 8001 3921
rect 7899 3639 7941 3681
rect 8139 3699 8181 3741
rect 8619 4179 8661 4221
rect 8439 3999 8481 4041
rect 8559 3999 8601 4041
rect 8259 3879 8301 3921
rect 8379 3879 8421 3921
rect 8199 3639 8241 3681
rect 7119 3279 7161 3321
rect 7119 3159 7161 3201
rect 7059 3099 7101 3141
rect 7599 3459 7641 3501
rect 7719 3459 7761 3501
rect 7539 3159 7581 3201
rect 7359 3039 7401 3081
rect 7359 2859 7401 2901
rect 7179 2742 7221 2784
rect 7299 2739 7341 2781
rect 7119 2616 7161 2658
rect 6759 2439 6801 2481
rect 6579 2319 6621 2361
rect 7179 2379 7221 2421
rect 7119 2259 7161 2301
rect 6579 2199 6621 2241
rect 6759 2199 6801 2241
rect 6879 2199 6921 2241
rect 7059 2199 7101 2241
rect 6099 1659 6141 1701
rect 6039 1599 6081 1641
rect 6099 1539 6141 1581
rect 5559 1419 5601 1461
rect 5139 1359 5181 1401
rect 5439 1359 5481 1401
rect 5199 1182 5241 1224
rect 5319 1182 5361 1224
rect 5919 1299 5961 1341
rect 5559 1182 5601 1224
rect 5799 1182 5841 1224
rect 5499 1056 5541 1098
rect 5859 1056 5901 1098
rect 5199 999 5241 1041
rect 6279 1899 6321 1941
rect 6399 1779 6441 1821
rect 6159 1182 6201 1224
rect 6639 2139 6681 2181
rect 6639 1956 6681 1998
rect 6819 1956 6861 1998
rect 6939 1956 6981 1998
rect 6579 1899 6621 1941
rect 6819 1659 6861 1701
rect 7119 2079 7161 2121
rect 7659 2919 7701 2961
rect 7599 2859 7641 2901
rect 7659 2742 7701 2784
rect 7359 2619 7401 2661
rect 7419 2439 7461 2481
rect 7299 2199 7341 2241
rect 7239 2139 7281 2181
rect 7419 2079 7461 2121
rect 7359 1956 7401 1998
rect 7599 2616 7641 2658
rect 7899 3159 7941 3201
rect 8019 3159 8061 3201
rect 8319 3819 8361 3861
rect 8259 3459 8301 3501
rect 8079 2919 8121 2961
rect 8559 3759 8601 3801
rect 9099 5559 9141 5601
rect 9039 5499 9081 5541
rect 8979 5319 9021 5361
rect 8799 5199 8841 5241
rect 8799 4899 8841 4941
rect 8739 4779 8781 4821
rect 8919 4659 8961 4701
rect 8919 4359 8961 4401
rect 9219 5379 9261 5421
rect 9459 5739 9501 5781
rect 9339 5619 9381 5661
rect 9459 5619 9501 5661
rect 9339 5319 9381 5361
rect 9279 5259 9321 5301
rect 9279 5076 9321 5118
rect 9459 4959 9501 5001
rect 9219 4839 9261 4881
rect 9219 4359 9261 4401
rect 9099 4299 9141 4341
rect 9339 4302 9381 4344
rect 9456 4302 9498 4344
rect 9819 8019 9861 8061
rect 9999 8199 10041 8241
rect 9939 8139 9981 8181
rect 9939 7899 9981 7941
rect 9879 7779 9921 7821
rect 9939 7719 9981 7761
rect 9819 7599 9861 7641
rect 10179 8199 10221 8241
rect 10119 7899 10161 7941
rect 10119 7779 10161 7821
rect 9999 7659 10041 7701
rect 9879 7479 9921 7521
rect 10059 7599 10101 7641
rect 9999 7422 10041 7464
rect 9819 7296 9861 7338
rect 9939 7239 9981 7281
rect 10779 9279 10821 9321
rect 10599 9159 10641 9201
rect 10359 9099 10401 9141
rect 10479 8982 10521 9024
rect 11319 9756 11361 9798
rect 11139 9339 11181 9381
rect 11499 9882 11541 9924
rect 11799 9939 11841 9981
rect 12099 9882 12141 9924
rect 11559 9756 11601 9798
rect 11679 9756 11721 9798
rect 11799 9756 11841 9798
rect 12039 9756 12081 9798
rect 11919 9699 11961 9741
rect 11499 9639 11541 9681
rect 11979 9639 12021 9681
rect 11499 9519 11541 9561
rect 11499 9399 11541 9441
rect 11379 9279 11421 9321
rect 11439 9219 11481 9261
rect 11079 8982 11121 9024
rect 11439 8982 11481 9024
rect 10359 8856 10401 8898
rect 10539 8856 10581 8898
rect 10359 8559 10401 8601
rect 10299 8319 10341 8361
rect 10479 8322 10521 8364
rect 10539 8196 10581 8238
rect 10419 8139 10461 8181
rect 10239 7599 10281 7641
rect 10779 8856 10821 8898
rect 10899 8856 10941 8898
rect 10719 8799 10761 8841
rect 11259 8850 11301 8892
rect 11199 8679 11241 8721
rect 12939 11976 12981 12018
rect 13059 11976 13101 12018
rect 12759 11439 12801 11481
rect 12819 11310 12861 11352
rect 12699 11139 12741 11181
rect 13059 10959 13101 11001
rect 12999 10899 13041 10941
rect 12759 10839 12801 10881
rect 12699 10539 12741 10581
rect 13476 14139 13518 14181
rect 13539 14139 13581 14181
rect 13479 13959 13521 14001
rect 13356 13779 13398 13821
rect 13419 13779 13461 13821
rect 13359 13662 13401 13704
rect 13599 13839 13641 13881
rect 13539 13719 13581 13761
rect 13479 13359 13521 13401
rect 13419 13239 13461 13281
rect 13359 13179 13401 13221
rect 13539 13299 13581 13341
rect 13536 13119 13578 13161
rect 13599 13119 13641 13161
rect 13719 14319 13761 14361
rect 14199 14919 14241 14961
rect 14139 14859 14181 14901
rect 14199 14799 14241 14841
rect 14319 14799 14361 14841
rect 14199 14619 14241 14661
rect 14139 14562 14181 14604
rect 14259 14562 14301 14604
rect 14439 15096 14481 15138
rect 14559 14979 14601 15021
rect 14499 14919 14541 14961
rect 14019 14496 14061 14538
rect 14319 14436 14361 14478
rect 14019 14319 14061 14361
rect 13959 14259 14001 14301
rect 13899 14139 13941 14181
rect 14079 14139 14121 14181
rect 13839 14019 13881 14061
rect 13839 13956 13881 13998
rect 13719 13779 13761 13821
rect 13719 13659 13761 13701
rect 13959 13899 14001 13941
rect 13899 13839 13941 13881
rect 13899 13719 13941 13761
rect 13719 13539 13761 13581
rect 13779 13479 13821 13521
rect 13719 13419 13761 13461
rect 13659 13059 13701 13101
rect 13839 13419 13881 13461
rect 13779 13299 13821 13341
rect 14136 14079 14178 14121
rect 14199 14079 14241 14121
rect 14439 14019 14481 14061
rect 14559 14619 14601 14661
rect 14979 15339 15021 15381
rect 15099 15879 15141 15921
rect 15459 16479 15501 16521
rect 15459 16299 15501 16341
rect 15399 16119 15441 16161
rect 15699 17556 15741 17598
rect 15819 17556 15861 17598
rect 15579 17439 15621 17481
rect 15879 17439 15921 17481
rect 15579 17259 15621 17301
rect 15879 17199 15921 17241
rect 15699 17139 15741 17181
rect 15579 17019 15621 17061
rect 15759 17079 15801 17121
rect 15699 16839 15741 16881
rect 15819 16959 15861 17001
rect 15939 17079 15981 17121
rect 15879 16899 15921 16941
rect 15819 16779 15861 16821
rect 15639 16656 15681 16698
rect 15579 16536 15621 16578
rect 15579 16419 15621 16461
rect 15579 16179 15621 16221
rect 15519 16119 15561 16161
rect 15279 15999 15321 16041
rect 15219 15819 15261 15861
rect 15159 15759 15201 15801
rect 15159 15639 15201 15681
rect 15099 15519 15141 15561
rect 14979 15096 15021 15138
rect 14859 14919 14901 14961
rect 14799 14679 14841 14721
rect 14799 14559 14841 14601
rect 14679 14436 14721 14478
rect 14619 14319 14661 14361
rect 14679 14259 14721 14301
rect 14619 14019 14661 14061
rect 14199 13776 14241 13818
rect 14439 13779 14481 13821
rect 14139 13719 14181 13761
rect 13959 13479 14001 13521
rect 13899 13299 13941 13341
rect 13839 13239 13881 13281
rect 13779 13059 13821 13101
rect 14079 13536 14121 13578
rect 14019 13419 14061 13461
rect 13959 13239 14001 13281
rect 13899 13179 13941 13221
rect 14079 13059 14121 13101
rect 13656 12879 13698 12921
rect 13719 12879 13761 12921
rect 13899 13002 13941 13044
rect 14019 13002 14061 13044
rect 14679 13719 14721 13761
rect 14319 13419 14361 13461
rect 14259 13359 14301 13401
rect 14199 13239 14241 13281
rect 14199 13176 14241 13218
rect 13839 12879 13881 12921
rect 13419 12699 13461 12741
rect 13539 12639 13581 12681
rect 13359 12339 13401 12381
rect 13239 12219 13281 12261
rect 13179 12099 13221 12141
rect 13179 11979 13221 12021
rect 13659 12339 13701 12381
rect 13779 12102 13821 12144
rect 14079 12876 14121 12918
rect 13899 12819 13941 12861
rect 14019 12819 14061 12861
rect 13899 12399 13941 12441
rect 13899 12336 13941 12378
rect 13239 11799 13281 11841
rect 13299 11679 13341 11721
rect 13239 11442 13281 11484
rect 13479 11442 13521 11484
rect 13179 11259 13221 11301
rect 13719 11976 13761 12018
rect 13839 11979 13881 12021
rect 13659 11856 13701 11898
rect 13779 11859 13821 11901
rect 14319 13179 14361 13221
rect 14439 13359 14481 13401
rect 14439 13119 14481 13161
rect 14979 14799 15021 14841
rect 15219 15579 15261 15621
rect 15159 15039 15201 15081
rect 15099 14739 15141 14781
rect 14979 14562 15021 14604
rect 15099 14562 15141 14604
rect 15399 15699 15441 15741
rect 15339 15459 15381 15501
rect 15699 16359 15741 16401
rect 15939 16479 15981 16521
rect 15759 16239 15801 16281
rect 15699 16179 15741 16221
rect 15639 16119 15681 16161
rect 15819 16179 15861 16221
rect 15759 15996 15801 16038
rect 15639 15819 15681 15861
rect 15519 15339 15561 15381
rect 15459 15279 15501 15321
rect 15279 15219 15321 15261
rect 15579 15279 15621 15321
rect 15279 15099 15321 15141
rect 15219 14559 15261 14601
rect 14979 14379 15021 14421
rect 14919 13779 14961 13821
rect 14859 13719 14901 13761
rect 15219 14439 15261 14481
rect 15039 14139 15081 14181
rect 15219 13899 15261 13941
rect 15519 15096 15561 15138
rect 15459 15039 15501 15081
rect 15399 14859 15441 14901
rect 15339 14739 15381 14781
rect 16839 18519 16881 18561
rect 16779 18459 16821 18501
rect 16299 18399 16341 18441
rect 16419 18399 16461 18441
rect 16539 18399 16581 18441
rect 16659 18399 16701 18441
rect 16179 18342 16221 18384
rect 16479 18342 16521 18384
rect 16779 18339 16821 18381
rect 16119 18219 16161 18261
rect 16419 18219 16461 18261
rect 16239 18099 16281 18141
rect 16539 18216 16581 18258
rect 16719 18216 16761 18258
rect 16419 18039 16461 18081
rect 16119 17979 16161 18021
rect 16239 17979 16281 18021
rect 16119 17682 16161 17724
rect 16599 17859 16641 17901
rect 16479 17799 16521 17841
rect 16419 17682 16461 17724
rect 16179 17556 16221 17598
rect 16419 17439 16461 17481
rect 16359 17319 16401 17361
rect 16419 17139 16461 17181
rect 16359 17079 16401 17121
rect 16599 17682 16641 17724
rect 16719 17682 16761 17724
rect 16659 17556 16701 17598
rect 16539 17259 16581 17301
rect 16599 17079 16641 17121
rect 16899 18459 16941 18501
rect 17559 18759 17601 18801
rect 17679 18639 17721 18681
rect 17499 18519 17541 18561
rect 17439 18399 17481 18441
rect 17199 18342 17241 18384
rect 17379 18279 17421 18321
rect 17139 18216 17181 18258
rect 17259 18159 17301 18201
rect 16959 18099 17001 18141
rect 17199 18099 17241 18141
rect 17259 17979 17301 18021
rect 17379 17979 17421 18021
rect 17199 17919 17241 17961
rect 16959 17859 17001 17901
rect 17079 17799 17121 17841
rect 17019 17556 17061 17598
rect 17139 17556 17181 17598
rect 17019 17379 17061 17421
rect 16539 16779 16581 16821
rect 16479 16656 16521 16698
rect 16299 16539 16341 16581
rect 16239 16479 16281 16521
rect 15999 16359 16041 16401
rect 15996 16239 16038 16281
rect 16059 16239 16101 16281
rect 16179 16179 16221 16221
rect 16059 16119 16101 16161
rect 16539 16599 16581 16641
rect 16479 16359 16521 16401
rect 16299 16122 16341 16164
rect 16839 17019 16881 17061
rect 16719 16782 16761 16824
rect 16839 16779 16881 16821
rect 16779 16656 16821 16698
rect 16719 16599 16761 16641
rect 16599 16239 16641 16281
rect 16779 16419 16821 16461
rect 16719 16119 16761 16161
rect 15999 15999 16041 16041
rect 16119 15996 16161 16038
rect 16239 15996 16281 16038
rect 16539 15996 16581 16038
rect 16659 15996 16701 16038
rect 16479 15879 16521 15921
rect 16239 15819 16281 15861
rect 16239 15699 16281 15741
rect 15939 15639 15981 15681
rect 16119 15639 16161 15681
rect 15759 15579 15801 15621
rect 16116 15519 16158 15561
rect 16179 15519 16221 15561
rect 15759 15222 15801 15264
rect 15879 15222 15921 15264
rect 16056 15222 16098 15264
rect 16119 15222 16161 15264
rect 16359 15459 16401 15501
rect 15639 14919 15681 14961
rect 15519 14619 15561 14661
rect 15699 14619 15741 14661
rect 15399 14559 15441 14601
rect 15579 14562 15621 14604
rect 15939 14979 15981 15021
rect 15999 14919 16041 14961
rect 16239 15222 16281 15264
rect 16419 15339 16461 15381
rect 16359 15219 16401 15261
rect 16299 15096 16341 15138
rect 16239 14979 16281 15021
rect 16119 14919 16161 14961
rect 16059 14859 16101 14901
rect 16119 14799 16161 14841
rect 15999 14679 16041 14721
rect 15819 14619 15861 14661
rect 15759 14559 15801 14601
rect 15339 14436 15381 14478
rect 15399 14319 15441 14361
rect 15519 14436 15561 14478
rect 16299 14919 16341 14961
rect 15699 14379 15741 14421
rect 15519 14199 15561 14241
rect 15639 14199 15681 14241
rect 15639 14079 15681 14121
rect 15459 13899 15501 13941
rect 15639 13899 15681 13941
rect 15279 13839 15321 13881
rect 15579 13839 15621 13881
rect 15159 13656 15201 13698
rect 15339 13662 15381 13704
rect 15459 13662 15501 13704
rect 15099 13599 15141 13641
rect 14859 13536 14901 13578
rect 14979 13479 15021 13521
rect 14739 13299 14781 13341
rect 14739 13179 14781 13221
rect 14379 13002 14421 13044
rect 14499 13002 14541 13044
rect 14679 13002 14721 13044
rect 14979 13059 15021 13101
rect 14919 12999 14961 13041
rect 14199 12459 14241 12501
rect 14019 12339 14061 12381
rect 13959 12279 14001 12321
rect 14079 12102 14121 12144
rect 14259 12099 14301 12141
rect 13899 11919 13941 11961
rect 13839 11619 13881 11661
rect 13659 11439 13701 11481
rect 13359 11259 13401 11301
rect 13479 11199 13521 11241
rect 13239 11139 13281 11181
rect 13359 11139 13401 11181
rect 13119 10719 13161 10761
rect 13119 10542 13161 10584
rect 12639 10119 12681 10161
rect 12279 9939 12321 9981
rect 12519 9939 12561 9981
rect 12219 9519 12261 9561
rect 12159 9339 12201 9381
rect 12039 9279 12081 9321
rect 11979 9159 12021 9201
rect 11619 9099 11661 9141
rect 11799 8988 11841 9030
rect 11919 8988 11961 9030
rect 11319 8619 11361 8661
rect 11439 8619 11481 8661
rect 11019 8559 11061 8601
rect 11199 8559 11241 8601
rect 10839 8322 10881 8364
rect 10959 8322 11001 8364
rect 11139 8319 11181 8361
rect 10839 8019 10881 8061
rect 10719 7779 10761 7821
rect 10479 7479 10521 7521
rect 10659 7479 10701 7521
rect 10179 7422 10221 7464
rect 10359 7422 10401 7464
rect 10419 7299 10461 7341
rect 10119 6939 10161 6981
rect 10239 6819 10281 6861
rect 9819 6759 9861 6801
rect 10059 6762 10101 6804
rect 10179 6762 10221 6804
rect 9819 6579 9861 6621
rect 9699 6519 9741 6561
rect 9759 6459 9801 6501
rect 9639 6279 9681 6321
rect 9639 6039 9681 6081
rect 9939 6339 9981 6381
rect 10179 6159 10221 6201
rect 10719 7422 10761 7464
rect 10899 7899 10941 7941
rect 10539 7359 10581 7401
rect 10539 7239 10581 7281
rect 10659 7179 10701 7221
rect 10539 6939 10581 6981
rect 10479 6819 10521 6861
rect 10419 6759 10461 6801
rect 10599 6879 10641 6921
rect 10539 6639 10581 6681
rect 10359 6219 10401 6261
rect 10056 5979 10098 6021
rect 10119 5979 10161 6021
rect 9759 5862 9801 5904
rect 9879 5862 9921 5904
rect 10059 5862 10101 5904
rect 10239 5862 10281 5904
rect 9579 5736 9621 5778
rect 9699 5736 9741 5778
rect 9879 5679 9921 5721
rect 9879 5559 9921 5601
rect 10179 5439 10221 5481
rect 9999 5379 10041 5421
rect 9759 5319 9801 5361
rect 9759 5202 9801 5244
rect 10179 5202 10221 5244
rect 10359 5199 10401 5241
rect 9879 5076 9921 5118
rect 9999 5079 10041 5121
rect 10119 5076 10161 5118
rect 10239 5079 10281 5121
rect 11079 8196 11121 8238
rect 11079 7899 11121 7941
rect 11259 8439 11301 8481
rect 11319 8319 11361 8361
rect 11439 8322 11481 8364
rect 11379 8196 11421 8238
rect 11499 8196 11541 8238
rect 11259 8019 11301 8061
rect 11259 7779 11301 7821
rect 11319 7659 11361 7701
rect 11259 7599 11301 7641
rect 11019 7299 11061 7341
rect 10839 6999 10881 7041
rect 10959 6999 11001 7041
rect 11199 7419 11241 7461
rect 11799 8439 11841 8481
rect 11619 8322 11661 8364
rect 12099 8982 12141 9024
rect 12219 8982 12261 9024
rect 12459 9882 12501 9924
rect 12579 9882 12621 9924
rect 12696 9879 12738 9921
rect 12759 9882 12801 9924
rect 12879 9882 12921 9924
rect 13179 10419 13221 10461
rect 13119 9939 13161 9981
rect 12339 9756 12381 9798
rect 12339 9639 12381 9681
rect 12339 9459 12381 9501
rect 11979 8859 12021 8901
rect 11979 8679 12021 8721
rect 11919 8379 11961 8421
rect 11619 8199 11661 8241
rect 11739 8196 11781 8238
rect 11559 8079 11601 8121
rect 11799 8079 11841 8121
rect 11559 7959 11601 8001
rect 11499 7419 11541 7461
rect 11259 7296 11301 7338
rect 11379 7296 11421 7338
rect 10659 6819 10701 6861
rect 10779 6819 10821 6861
rect 10599 6579 10641 6621
rect 10839 6762 10881 6804
rect 10959 6768 11001 6810
rect 10719 6579 10761 6621
rect 10779 6519 10821 6561
rect 11199 6999 11241 7041
rect 11499 6999 11541 7041
rect 11139 6459 11181 6501
rect 10719 6279 10761 6321
rect 10779 6219 10821 6261
rect 10659 6099 10701 6141
rect 10539 5979 10581 6021
rect 10659 5919 10701 5961
rect 10959 6099 11001 6141
rect 10899 5919 10941 5961
rect 10599 5736 10641 5778
rect 10599 5619 10641 5661
rect 10899 5736 10941 5778
rect 10719 5559 10761 5601
rect 10479 5202 10521 5244
rect 10599 5202 10641 5244
rect 10719 5199 10761 5241
rect 9999 5016 10041 5058
rect 9699 4839 9741 4881
rect 9759 4779 9801 4821
rect 9819 4539 9861 4581
rect 9759 4479 9801 4521
rect 9579 4359 9621 4401
rect 8679 4119 8721 4161
rect 8439 3642 8481 3684
rect 8859 4176 8901 4218
rect 8979 4176 9021 4218
rect 8859 3999 8901 4041
rect 8739 3642 8781 3684
rect 8379 3519 8421 3561
rect 8619 3516 8661 3558
rect 8739 3516 8781 3558
rect 8919 3516 8961 3558
rect 9159 4176 9201 4218
rect 9279 4059 9321 4101
rect 9399 4059 9441 4101
rect 9279 3879 9321 3921
rect 9099 3759 9141 3801
rect 9279 3699 9321 3741
rect 9219 3642 9261 3684
rect 9339 3642 9381 3684
rect 9519 4299 9561 4341
rect 9759 4302 9801 4344
rect 9879 4359 9921 4401
rect 9936 4302 9978 4344
rect 10419 5076 10461 5118
rect 11079 5862 11121 5904
rect 11979 8199 12021 8241
rect 11979 7959 12021 8001
rect 11859 7659 11901 7701
rect 12159 8856 12201 8898
rect 12279 8859 12321 8901
rect 12519 9756 12561 9798
rect 12459 9639 12501 9681
rect 12399 9219 12441 9261
rect 12399 9099 12441 9141
rect 12399 8919 12441 8961
rect 12639 9519 12681 9561
rect 12639 9279 12681 9321
rect 12519 9159 12561 9201
rect 13059 9879 13101 9921
rect 12759 9759 12801 9801
rect 12939 9759 12981 9801
rect 13059 9759 13101 9801
rect 12999 9699 13041 9741
rect 13239 10359 13281 10401
rect 13299 10299 13341 10341
rect 13239 10179 13281 10221
rect 13239 9999 13281 10041
rect 13479 10899 13521 10941
rect 13719 11316 13761 11358
rect 14139 11976 14181 12018
rect 14259 11976 14301 12018
rect 14019 11919 14061 11961
rect 13959 11799 14001 11841
rect 13959 11199 14001 11241
rect 13659 11139 13701 11181
rect 13899 11139 13941 11181
rect 13599 10899 13641 10941
rect 13539 10779 13581 10821
rect 13419 10659 13461 10701
rect 13599 10659 13641 10701
rect 13479 10542 13521 10584
rect 13959 11079 14001 11121
rect 13899 10779 13941 10821
rect 13659 10539 13701 10581
rect 13419 10419 13461 10461
rect 13599 10359 13641 10401
rect 13539 10179 13581 10221
rect 13419 9999 13461 10041
rect 13359 9939 13401 9981
rect 13419 9882 13461 9924
rect 13179 9699 13221 9741
rect 13299 9699 13341 9741
rect 13119 9639 13161 9681
rect 13059 9399 13101 9441
rect 12939 9219 12981 9261
rect 13239 9339 13281 9381
rect 12879 9159 12921 9201
rect 13179 9159 13221 9201
rect 12699 9099 12741 9141
rect 12819 9099 12861 9141
rect 12699 8982 12741 9024
rect 12459 8799 12501 8841
rect 12339 8679 12381 8721
rect 12279 8619 12321 8661
rect 12099 8499 12141 8541
rect 12639 8856 12681 8898
rect 12819 8859 12861 8901
rect 12759 8799 12801 8841
rect 13239 9039 13281 9081
rect 13059 8982 13101 9024
rect 13179 8982 13221 9024
rect 13539 9399 13581 9441
rect 13479 9339 13521 9381
rect 13299 8979 13341 9021
rect 12879 8739 12921 8781
rect 12819 8619 12861 8661
rect 12519 8559 12561 8601
rect 12759 8559 12801 8601
rect 12759 8439 12801 8481
rect 12339 8379 12381 8421
rect 12279 8319 12321 8361
rect 12459 8319 12501 8361
rect 12579 8322 12621 8364
rect 12699 8322 12741 8364
rect 13239 8859 13281 8901
rect 12999 8739 13041 8781
rect 13119 8739 13161 8781
rect 12999 8619 13041 8661
rect 12819 8319 12861 8361
rect 12219 8196 12261 8238
rect 12099 8079 12141 8121
rect 12219 7719 12261 7761
rect 11679 7422 11721 7464
rect 11739 7179 11781 7221
rect 12039 7599 12081 7641
rect 12099 7479 12141 7521
rect 12279 7599 12321 7641
rect 12219 7419 12261 7461
rect 12039 7296 12081 7338
rect 12219 7296 12261 7338
rect 12159 7239 12201 7281
rect 11859 7119 11901 7161
rect 12039 7119 12081 7161
rect 11619 6879 11661 6921
rect 11799 6819 11841 6861
rect 11559 6759 11601 6801
rect 11919 6762 11961 6804
rect 12159 6999 12201 7041
rect 12099 6762 12141 6804
rect 11619 6696 11661 6738
rect 11499 6630 11541 6672
rect 11679 6639 11721 6681
rect 11619 6459 11661 6501
rect 11319 6399 11361 6441
rect 11559 6399 11601 6441
rect 11859 6636 11901 6678
rect 11979 6636 12021 6678
rect 11739 6519 11781 6561
rect 11859 6519 11901 6561
rect 12039 6519 12081 6561
rect 11799 6459 11841 6501
rect 11739 6339 11781 6381
rect 11739 5919 11781 5961
rect 11139 5736 11181 5778
rect 11139 5499 11181 5541
rect 10959 5379 11001 5421
rect 10839 5319 10881 5361
rect 10239 4659 10281 4701
rect 10299 4539 10341 4581
rect 10239 4359 10281 4401
rect 9519 4179 9561 4221
rect 9636 4179 9678 4221
rect 9459 3999 9501 4041
rect 9279 3516 9321 3558
rect 9399 3519 9441 3561
rect 8499 3459 8541 3501
rect 9039 3459 9081 3501
rect 8679 3099 8721 3141
rect 8379 3039 8421 3081
rect 8499 2919 8541 2961
rect 9459 3099 9501 3141
rect 9399 2979 9441 3021
rect 9159 2919 9201 2961
rect 8679 2859 8721 2901
rect 8979 2859 9021 2901
rect 7959 2616 8001 2658
rect 7779 2559 7821 2601
rect 7899 2559 7941 2601
rect 7659 2259 7701 2301
rect 7779 2082 7821 2124
rect 7599 1956 7641 1998
rect 7239 1839 7281 1881
rect 7479 1839 7521 1881
rect 7059 1599 7101 1641
rect 7719 1599 7761 1641
rect 7059 1419 7101 1461
rect 7119 1299 7161 1341
rect 7359 1299 7401 1341
rect 7839 1299 7881 1341
rect 6639 1239 6681 1281
rect 6699 1182 6741 1224
rect 7239 1182 7281 1224
rect 7719 1182 7761 1224
rect 6279 1056 6321 1098
rect 6399 1056 6441 1098
rect 6516 1056 6558 1098
rect 6579 1056 6621 1098
rect 6759 1056 6801 1098
rect 6879 1056 6921 1098
rect 7119 1059 7161 1101
rect 6099 999 6141 1041
rect 6219 939 6261 981
rect 5199 879 5241 921
rect 5319 879 5361 921
rect 5139 819 5181 861
rect 4899 639 4941 681
rect 5079 639 5121 681
rect 4959 579 5001 621
rect 4839 519 4881 561
rect 4539 396 4581 438
rect 4659 396 4701 438
rect 5979 819 6021 861
rect 6039 759 6081 801
rect 6339 759 6381 801
rect 5379 639 5421 681
rect 5979 639 6021 681
rect 5199 522 5241 564
rect 5139 396 5181 438
rect 4779 279 4821 321
rect 4959 279 5001 321
rect 4479 219 4521 261
rect 5259 339 5301 381
rect 5859 579 5901 621
rect 5559 522 5601 564
rect 5679 522 5721 564
rect 5799 519 5841 561
rect 5499 396 5541 438
rect 5619 396 5661 438
rect 6279 639 6321 681
rect 6159 522 6201 564
rect 5859 396 5901 438
rect 5979 396 6021 438
rect 6099 396 6141 438
rect 6219 396 6261 438
rect 7419 1056 7461 1098
rect 7659 1056 7701 1098
rect 7839 1059 7881 1101
rect 7779 819 7821 861
rect 7659 759 7701 801
rect 6759 699 6801 741
rect 7299 699 7341 741
rect 6639 639 6681 681
rect 6519 579 6561 621
rect 6339 396 6381 438
rect 7239 639 7281 681
rect 7359 639 7401 681
rect 7299 579 7341 621
rect 6879 522 6921 564
rect 7059 522 7101 564
rect 7419 522 7461 564
rect 7599 522 7641 564
rect 5799 279 5841 321
rect 5379 219 5421 261
rect 5139 159 5181 201
rect 6459 396 6501 438
rect 6579 396 6621 438
rect 6759 396 6801 438
rect 6939 396 6981 438
rect 7239 339 7281 381
rect 7059 279 7101 321
rect 7959 2379 8001 2421
rect 8259 2616 8301 2658
rect 8079 2259 8121 2301
rect 8079 2196 8121 2238
rect 8139 2139 8181 2181
rect 8079 1956 8121 1998
rect 8199 1719 8241 1761
rect 7959 1659 8001 1701
rect 7959 1539 8001 1581
rect 8259 1359 8301 1401
rect 8859 2742 8901 2784
rect 9339 2859 9381 2901
rect 9339 2742 9381 2784
rect 8799 2616 8841 2658
rect 9159 2616 9201 2658
rect 9279 2616 9321 2658
rect 9399 2499 9441 2541
rect 8919 2439 8961 2481
rect 9399 2379 9441 2421
rect 9039 2199 9081 2241
rect 8979 2139 9021 2181
rect 8919 2079 8961 2121
rect 8439 1959 8481 2001
rect 8559 1956 8601 1998
rect 8739 1839 8781 1881
rect 9279 2082 9321 2124
rect 9579 3999 9621 4041
rect 9699 4176 9741 4218
rect 9816 4176 9858 4218
rect 9879 4179 9921 4221
rect 9999 4299 10041 4341
rect 10119 4302 10161 4344
rect 10059 4176 10101 4218
rect 10179 4176 10221 4218
rect 10299 4179 10341 4221
rect 9939 4059 9981 4101
rect 9999 3819 10041 3861
rect 9699 3759 9741 3801
rect 9639 3699 9681 3741
rect 9579 3639 9621 3681
rect 9639 3516 9681 3558
rect 9759 3516 9801 3558
rect 9579 3459 9621 3501
rect 9759 2799 9801 2841
rect 10239 3699 10281 3741
rect 10059 3639 10101 3681
rect 10179 3642 10221 3684
rect 10539 5076 10581 5118
rect 10779 5076 10821 5118
rect 10659 4899 10701 4941
rect 10839 4659 10881 4701
rect 10539 4479 10581 4521
rect 10419 4302 10461 4344
rect 10659 4302 10701 4344
rect 10959 4779 11001 4821
rect 10899 4419 10941 4461
rect 11199 4479 11241 4521
rect 11079 4302 11121 4344
rect 10479 4179 10521 4221
rect 10419 4059 10461 4101
rect 10359 3819 10401 3861
rect 10839 4179 10881 4221
rect 11139 4179 11181 4221
rect 10719 4059 10761 4101
rect 10899 4059 10941 4101
rect 11019 4059 11061 4101
rect 10599 3879 10641 3921
rect 10839 3879 10881 3921
rect 10719 3759 10761 3801
rect 10479 3699 10521 3741
rect 10599 3699 10641 3741
rect 10419 3639 10461 3681
rect 9999 3579 10041 3621
rect 10239 3516 10281 3558
rect 10479 3516 10521 3558
rect 10659 3516 10701 3558
rect 10779 3516 10821 3558
rect 10899 3516 10941 3558
rect 10359 3399 10401 3441
rect 10779 3099 10821 3141
rect 10659 2979 10701 3021
rect 10059 2799 10101 2841
rect 9939 2742 9981 2784
rect 10179 2742 10221 2784
rect 11079 3516 11121 3558
rect 11199 3459 11241 3501
rect 11079 3399 11121 3441
rect 11379 5862 11421 5904
rect 11499 5862 11541 5904
rect 11679 5862 11721 5904
rect 11319 5619 11361 5661
rect 11439 5559 11481 5601
rect 11379 5379 11421 5421
rect 11679 5619 11721 5661
rect 11559 5319 11601 5361
rect 11979 6219 12021 6261
rect 11859 5862 11901 5904
rect 12099 5739 12141 5781
rect 11919 5619 11961 5661
rect 12639 8079 12681 8121
rect 12819 8199 12861 8241
rect 12759 8019 12801 8061
rect 12519 7839 12561 7881
rect 12339 7479 12381 7521
rect 12459 7479 12501 7521
rect 12639 7422 12681 7464
rect 12819 7422 12861 7464
rect 12339 7299 12381 7341
rect 12459 7239 12501 7281
rect 12579 7059 12621 7101
rect 12939 8439 12981 8481
rect 13359 8850 13401 8892
rect 13299 8619 13341 8661
rect 14139 11316 14181 11358
rect 14439 12876 14481 12918
rect 14799 12876 14841 12918
rect 14559 12759 14601 12801
rect 14679 12759 14721 12801
rect 14859 12759 14901 12801
rect 14379 12639 14421 12681
rect 14499 12639 14541 12681
rect 14379 12519 14421 12561
rect 14379 12456 14421 12498
rect 14619 12279 14661 12321
rect 14499 12102 14541 12144
rect 14799 12459 14841 12501
rect 14799 12339 14841 12381
rect 15159 13479 15201 13521
rect 15159 13119 15201 13161
rect 15099 13059 15141 13101
rect 15279 13419 15321 13461
rect 15519 13539 15561 13581
rect 15279 13299 15321 13341
rect 15399 13299 15441 13341
rect 15219 13059 15261 13101
rect 15399 13179 15441 13221
rect 15339 13119 15381 13161
rect 15279 13002 15321 13044
rect 15039 12879 15081 12921
rect 14979 12639 15021 12681
rect 15159 12759 15201 12801
rect 15099 12699 15141 12741
rect 15159 12519 15201 12561
rect 15279 12819 15321 12861
rect 15219 12399 15261 12441
rect 15039 12339 15081 12381
rect 14919 12219 14961 12261
rect 15219 12219 15261 12261
rect 14679 12099 14721 12141
rect 14499 11919 14541 11961
rect 14379 11799 14421 11841
rect 14559 11859 14601 11901
rect 14619 11799 14661 11841
rect 14319 10899 14361 10941
rect 14379 10779 14421 10821
rect 14079 10659 14121 10701
rect 14019 10539 14061 10581
rect 14259 10548 14301 10590
rect 13899 10359 13941 10401
rect 13719 10119 13761 10161
rect 13659 9939 13701 9981
rect 13839 9939 13881 9981
rect 13719 9882 13761 9924
rect 13659 9759 13701 9801
rect 13779 9756 13821 9798
rect 13659 9639 13701 9681
rect 13899 9639 13941 9681
rect 14079 10359 14121 10401
rect 14379 10299 14421 10341
rect 14439 10179 14481 10221
rect 14739 11739 14781 11781
rect 14679 11619 14721 11661
rect 15039 11739 15081 11781
rect 15459 12999 15501 13041
rect 15639 13299 15681 13341
rect 15579 13179 15621 13221
rect 15639 13002 15681 13044
rect 15819 14436 15861 14478
rect 15939 14436 15981 14478
rect 16239 14436 16281 14478
rect 16059 14319 16101 14361
rect 15759 14199 15801 14241
rect 16119 14199 16161 14241
rect 15759 14079 15801 14121
rect 16059 13959 16101 14001
rect 16059 13779 16101 13821
rect 15939 13719 15981 13761
rect 15819 13662 15861 13704
rect 16239 13779 16281 13821
rect 16119 13659 16161 13701
rect 16359 14619 16401 14661
rect 16539 15579 16581 15621
rect 16479 15219 16521 15261
rect 17139 17259 17181 17301
rect 17379 17916 17421 17958
rect 17559 17859 17601 17901
rect 17499 17682 17541 17724
rect 17619 17559 17661 17601
rect 17559 17439 17601 17481
rect 17439 17379 17481 17421
rect 17259 17079 17301 17121
rect 17559 17079 17601 17121
rect 17139 17019 17181 17061
rect 17019 16779 17061 16821
rect 17499 16899 17541 16941
rect 18219 18759 18261 18801
rect 17999 18639 18041 18681
rect 17799 18399 17841 18441
rect 17679 17499 17721 17541
rect 17619 16899 17661 16941
rect 17259 16782 17301 16824
rect 17499 16782 17541 16824
rect 17019 16659 17061 16701
rect 17379 16659 17421 16701
rect 17199 16599 17241 16641
rect 16959 16419 17001 16461
rect 16779 15459 16821 15501
rect 16899 16239 16941 16281
rect 17079 16239 17121 16281
rect 17199 16239 17241 16281
rect 16959 16122 17001 16164
rect 17559 16656 17601 16698
rect 17859 18159 17901 18201
rect 17799 17919 17841 17961
rect 17799 17799 17841 17841
rect 17919 17979 17961 18021
rect 18099 17799 18141 17841
rect 17859 17682 17901 17724
rect 17919 17556 17961 17598
rect 18099 17559 18141 17601
rect 17859 17499 17901 17541
rect 17799 17019 17841 17061
rect 17499 16539 17541 16581
rect 17619 16539 17661 16581
rect 17439 16359 17481 16401
rect 17259 16179 17301 16221
rect 17379 16179 17421 16221
rect 17019 15879 17061 15921
rect 17199 15999 17241 16041
rect 17139 15819 17181 15861
rect 17499 16119 17541 16161
rect 17439 15996 17481 16038
rect 17559 15999 17601 16041
rect 17439 15879 17481 15921
rect 17379 15819 17421 15861
rect 17259 15759 17301 15801
rect 17319 15699 17361 15741
rect 17199 15579 17241 15621
rect 17019 15519 17061 15561
rect 16839 15339 16881 15381
rect 16599 15096 16641 15138
rect 16719 15096 16761 15138
rect 16839 15096 16881 15138
rect 16539 14562 16581 14604
rect 16779 14799 16821 14841
rect 16719 14619 16761 14661
rect 16659 14559 16701 14601
rect 16299 13719 16341 13761
rect 16479 14436 16521 14478
rect 16419 14079 16461 14121
rect 16359 13662 16401 13704
rect 16659 14439 16701 14481
rect 16659 14079 16701 14121
rect 16599 13899 16641 13941
rect 17019 15399 17061 15441
rect 17139 15222 17181 15264
rect 17079 15096 17121 15138
rect 17199 14979 17241 15021
rect 16959 14919 17001 14961
rect 17139 14919 17181 14961
rect 16899 14679 16941 14721
rect 16839 14619 16881 14661
rect 16779 14559 16821 14601
rect 17079 14859 17121 14901
rect 17259 14859 17301 14901
rect 17799 16659 17841 16701
rect 17979 16899 18021 16941
rect 18339 17859 18381 17901
rect 18279 17559 18321 17601
rect 18039 16659 18081 16701
rect 17859 16539 17901 16581
rect 17979 16419 18021 16461
rect 17859 16239 17901 16281
rect 17799 15996 17841 16038
rect 17679 15879 17721 15921
rect 17619 15699 17661 15741
rect 17559 15399 17601 15441
rect 18219 16659 18261 16701
rect 18279 16419 18321 16461
rect 18099 16299 18141 16341
rect 18279 16299 18321 16341
rect 18399 17079 18441 17121
rect 18339 16119 18381 16161
rect 18339 15999 18381 16041
rect 18039 15819 18081 15861
rect 18159 15819 18201 15861
rect 18159 15639 18201 15681
rect 18099 15579 18141 15621
rect 17979 15339 18021 15381
rect 18279 15339 18321 15381
rect 17679 15279 17721 15321
rect 17919 15279 17961 15321
rect 17559 15222 17601 15264
rect 18099 15222 18141 15264
rect 18219 15222 18261 15264
rect 17919 15096 17961 15138
rect 17799 15039 17841 15081
rect 17499 14979 17541 15021
rect 17619 14979 17661 15021
rect 17739 14979 17781 15021
rect 17439 14859 17481 14901
rect 17379 14799 17421 14841
rect 17139 14676 17181 14718
rect 17079 14559 17121 14601
rect 16899 14436 16941 14478
rect 17079 14439 17121 14481
rect 16899 14319 16941 14361
rect 16959 14019 17001 14061
rect 16899 13959 16941 14001
rect 16539 13839 16581 13881
rect 16719 13839 16761 13881
rect 16479 13659 16521 13701
rect 15759 13539 15801 13581
rect 15759 13419 15801 13461
rect 15819 13119 15861 13161
rect 15459 12699 15501 12741
rect 15519 12639 15561 12681
rect 15399 12279 15441 12321
rect 15519 12279 15561 12321
rect 15339 12159 15381 12201
rect 15459 12159 15501 12201
rect 16059 13539 16101 13581
rect 15999 13359 16041 13401
rect 15999 13002 16041 13044
rect 16179 13479 16221 13521
rect 16419 13539 16461 13581
rect 16119 13419 16161 13461
rect 15819 12879 15861 12921
rect 15939 12876 15981 12918
rect 15759 12819 15801 12861
rect 15939 12699 15981 12741
rect 16179 13299 16221 13341
rect 16419 13419 16461 13461
rect 16239 13002 16281 13044
rect 16359 13002 16401 13044
rect 16659 13779 16701 13821
rect 16839 13662 16881 13704
rect 16959 13839 17001 13881
rect 16599 13479 16641 13521
rect 16539 13359 16581 13401
rect 16479 12999 16521 13041
rect 16119 12579 16161 12621
rect 16419 12876 16461 12918
rect 16419 12813 16461 12855
rect 16179 12399 16221 12441
rect 16299 12399 16341 12441
rect 15639 12339 15681 12381
rect 16059 12339 16101 12381
rect 15279 11976 15321 12018
rect 15399 11976 15441 12018
rect 15339 11859 15381 11901
rect 15279 11799 15321 11841
rect 15279 11679 15321 11721
rect 15219 11619 15261 11661
rect 15039 11559 15081 11601
rect 14679 11316 14721 11358
rect 14799 11316 14841 11358
rect 14799 11253 14841 11295
rect 14679 10779 14721 10821
rect 14679 10659 14721 10701
rect 14319 10059 14361 10101
rect 14199 9999 14241 10041
rect 14499 9939 14541 9981
rect 14439 9879 14481 9921
rect 14259 9756 14301 9798
rect 14079 9639 14121 9681
rect 14319 9639 14361 9681
rect 14019 9579 14061 9621
rect 14259 9579 14301 9621
rect 13959 9219 14001 9261
rect 13899 9099 13941 9141
rect 13719 8988 13761 9030
rect 13959 8979 14001 9021
rect 13659 8859 13701 8901
rect 13959 8859 14001 8901
rect 13659 8739 13701 8781
rect 13599 8679 13641 8721
rect 13779 8559 13821 8601
rect 13599 8499 13641 8541
rect 13539 8439 13581 8481
rect 13659 8439 13701 8481
rect 13359 8319 13401 8361
rect 13539 8322 13581 8364
rect 13119 8196 13161 8238
rect 13299 8199 13341 8241
rect 13239 8079 13281 8121
rect 12999 7719 13041 7761
rect 13179 7719 13221 7761
rect 13179 7656 13221 7698
rect 12939 7599 12981 7641
rect 13179 7419 13221 7461
rect 12819 6999 12861 7041
rect 12339 6939 12381 6981
rect 12459 6939 12501 6981
rect 12579 6939 12621 6981
rect 12879 6939 12921 6981
rect 12279 6819 12321 6861
rect 12399 6636 12441 6678
rect 12279 6579 12321 6621
rect 12219 6339 12261 6381
rect 12459 6039 12501 6081
rect 12279 5919 12321 5961
rect 12519 5979 12561 6021
rect 12279 5736 12321 5778
rect 11919 5556 11961 5598
rect 12159 5559 12201 5601
rect 11499 5202 11541 5244
rect 11679 5202 11721 5244
rect 11799 5202 11841 5244
rect 12159 5496 12201 5538
rect 11979 5379 12021 5421
rect 11559 5076 11601 5118
rect 11919 5199 11961 5241
rect 11739 5079 11781 5121
rect 11439 4779 11481 4821
rect 11559 4779 11601 4821
rect 11379 4539 11421 4581
rect 11319 4302 11361 4344
rect 11439 4302 11481 4344
rect 11319 4119 11361 4161
rect 11379 4059 11421 4101
rect 11559 4059 11601 4101
rect 11739 4839 11781 4881
rect 11919 5079 11961 5121
rect 11859 4359 11901 4401
rect 11799 4302 11841 4344
rect 11919 4302 11961 4344
rect 12219 5379 12261 5421
rect 12159 5259 12201 5301
rect 12099 5202 12141 5244
rect 12399 5319 12441 5361
rect 12639 6819 12681 6861
rect 12759 6762 12801 6804
rect 12999 7296 13041 7338
rect 13119 7296 13161 7338
rect 13299 7899 13341 7941
rect 13359 7839 13401 7881
rect 13599 8196 13641 8238
rect 13719 8199 13761 8241
rect 13719 8079 13761 8121
rect 13599 7719 13641 7761
rect 13479 7659 13521 7701
rect 13359 7599 13401 7641
rect 13479 7539 13521 7581
rect 13359 7422 13401 7464
rect 14079 8850 14121 8892
rect 14019 8559 14061 8601
rect 13959 8439 14001 8481
rect 13899 8322 13941 8364
rect 14259 8559 14301 8601
rect 14379 9339 14421 9381
rect 14379 8979 14421 9021
rect 15039 11199 15081 11241
rect 15279 11442 15321 11484
rect 16119 12159 16161 12201
rect 15759 12102 15801 12144
rect 15699 11979 15741 12021
rect 15639 11739 15681 11781
rect 15819 11859 15861 11901
rect 15759 11739 15801 11781
rect 15699 11559 15741 11601
rect 15159 11319 15201 11361
rect 15099 11019 15141 11061
rect 15039 10959 15081 11001
rect 15039 10839 15081 10881
rect 15399 11199 15441 11241
rect 15219 11079 15261 11121
rect 14979 10548 15021 10590
rect 15339 10659 15381 10701
rect 15099 10539 15141 10581
rect 15036 10419 15078 10461
rect 14679 10059 14721 10101
rect 14619 9939 14661 9981
rect 14739 9939 14781 9981
rect 14919 9879 14961 9921
rect 14799 9756 14841 9798
rect 14919 9699 14961 9741
rect 14619 9519 14661 9561
rect 14859 9519 14901 9561
rect 14679 9459 14721 9501
rect 14799 9459 14841 9501
rect 14559 9279 14601 9321
rect 14619 9099 14661 9141
rect 14739 9339 14781 9381
rect 14679 9039 14721 9081
rect 14619 8988 14661 9030
rect 14679 8856 14721 8898
rect 14679 8679 14721 8721
rect 14499 8559 14541 8601
rect 14199 8499 14241 8541
rect 14319 8499 14361 8541
rect 14139 8439 14181 8481
rect 14079 8319 14121 8361
rect 13959 8196 14001 8238
rect 14079 8199 14121 8241
rect 13899 7839 13941 7881
rect 13839 7779 13881 7821
rect 13839 7599 13881 7641
rect 13899 7539 13941 7581
rect 13659 7479 13701 7521
rect 13779 7482 13821 7524
rect 13599 7359 13641 7401
rect 13059 7239 13101 7281
rect 13059 7119 13101 7161
rect 12999 7059 13041 7101
rect 12939 6759 12981 6801
rect 12819 6636 12861 6678
rect 13059 6759 13101 6801
rect 13239 7296 13281 7338
rect 13419 7296 13461 7338
rect 13419 6999 13461 7041
rect 13599 6999 13641 7041
rect 13299 6762 13341 6804
rect 13119 6459 13161 6501
rect 12999 6279 13041 6321
rect 13419 6639 13461 6681
rect 13359 6339 13401 6381
rect 12639 6219 12681 6261
rect 13239 6219 13281 6261
rect 13479 6339 13521 6381
rect 12759 5979 12801 6021
rect 12939 5979 12981 6021
rect 12741 5919 12783 5961
rect 12639 5859 12681 5901
rect 12819 5862 12861 5904
rect 13419 5976 13461 6018
rect 12999 5919 13041 5961
rect 13179 5862 13221 5904
rect 13299 5862 13341 5904
rect 12999 5799 13041 5841
rect 12759 5736 12801 5778
rect 12939 5739 12981 5781
rect 12639 5619 12681 5661
rect 12879 5619 12921 5661
rect 12579 5259 12621 5301
rect 12819 5559 12861 5601
rect 12159 5076 12201 5118
rect 12399 5076 12441 5118
rect 12099 5019 12141 5061
rect 12279 5019 12321 5061
rect 11739 4176 11781 4218
rect 11619 3999 11661 4041
rect 11859 4059 11901 4101
rect 11739 3939 11781 3981
rect 12519 5076 12561 5118
rect 12699 5019 12741 5061
rect 12459 4959 12501 5001
rect 12519 4539 12561 4581
rect 12219 4302 12261 4344
rect 12399 4302 12441 4344
rect 12099 4176 12141 4218
rect 12279 4176 12321 4218
rect 13059 5739 13101 5781
rect 12999 5679 13041 5721
rect 12939 5439 12981 5481
rect 13119 5679 13161 5721
rect 13299 5679 13341 5721
rect 13239 5559 13281 5601
rect 13059 5319 13101 5361
rect 13239 5319 13281 5361
rect 12879 5259 12921 5301
rect 13059 5202 13101 5244
rect 13059 4959 13101 5001
rect 12999 4839 13041 4881
rect 13119 4779 13161 4821
rect 13059 4719 13101 4761
rect 12879 4659 12921 4701
rect 12939 4479 12981 4521
rect 12579 4419 12621 4461
rect 12819 4419 12861 4461
rect 12519 3819 12561 3861
rect 11679 3759 11721 3801
rect 11859 3759 11901 3801
rect 12039 3759 12081 3801
rect 11439 3642 11481 3684
rect 11559 3642 11601 3684
rect 11979 3642 12021 3684
rect 12339 3759 12381 3801
rect 12159 3639 12201 3681
rect 12459 3642 12501 3684
rect 11799 3516 11841 3558
rect 11919 3516 11961 3558
rect 12099 3516 12141 3558
rect 11499 3459 11541 3501
rect 11259 3099 11301 3141
rect 11019 2979 11061 3021
rect 10959 2799 11001 2841
rect 11139 2799 11181 2841
rect 11259 2739 11301 2781
rect 10899 2679 10941 2721
rect 9519 2616 9561 2658
rect 9819 2616 9861 2658
rect 9999 2616 10041 2658
rect 10119 2616 10161 2658
rect 9519 2319 9561 2361
rect 9699 2319 9741 2361
rect 10359 2616 10401 2658
rect 10599 2616 10641 2658
rect 10719 2616 10761 2658
rect 11079 2616 11121 2658
rect 9639 2199 9681 2241
rect 9759 2199 9801 2241
rect 10059 2199 10101 2241
rect 10239 2199 10281 2241
rect 10179 2082 10221 2124
rect 10299 2079 10341 2121
rect 8979 1956 9021 1998
rect 9099 1956 9141 1998
rect 8919 1779 8961 1821
rect 8859 1719 8901 1761
rect 8499 1299 8541 1341
rect 8559 1299 8601 1341
rect 8259 1182 8301 1224
rect 9579 1956 9621 1998
rect 9699 1956 9741 1998
rect 9819 1839 9861 1881
rect 9999 1839 10041 1881
rect 10299 1899 10341 1941
rect 10539 2499 10581 2541
rect 10659 2439 10701 2481
rect 10779 2439 10821 2481
rect 11199 2439 11241 2481
rect 10659 2199 10701 2241
rect 10899 2319 10941 2361
rect 10839 2199 10881 2241
rect 10839 2079 10881 2121
rect 11019 2139 11061 2181
rect 11199 2139 11241 2181
rect 10599 1956 10641 1998
rect 10779 1959 10821 2001
rect 10959 1956 11001 1998
rect 11079 1956 11121 1998
rect 11259 2079 11301 2121
rect 11859 3399 11901 3441
rect 11859 3219 11901 3261
rect 11499 2919 11541 2961
rect 11619 2742 11661 2784
rect 12099 2859 12141 2901
rect 11979 2742 12021 2784
rect 12399 3459 12441 3501
rect 12759 4302 12801 4344
rect 13779 7419 13821 7461
rect 14139 7899 14181 7941
rect 14439 8439 14481 8481
rect 14319 8322 14361 8364
rect 15159 10410 15201 10452
rect 15219 10179 15261 10221
rect 15099 10059 15141 10101
rect 15099 9882 15141 9924
rect 15039 9759 15081 9801
rect 14979 9639 15021 9681
rect 15099 9639 15141 9681
rect 14919 9219 14961 9261
rect 14919 9099 14961 9141
rect 15039 9099 15081 9141
rect 14859 8979 14901 9021
rect 14976 8982 15018 9024
rect 15039 8979 15081 9021
rect 14739 8439 14781 8481
rect 14499 8319 14541 8361
rect 14259 8199 14301 8241
rect 14079 7719 14121 7761
rect 13959 7296 14001 7338
rect 14079 7296 14121 7338
rect 14499 8199 14541 8241
rect 14439 8139 14481 8181
rect 14379 8079 14421 8121
rect 14439 8019 14481 8061
rect 14259 7659 14301 7701
rect 14319 7422 14361 7464
rect 14739 8190 14781 8232
rect 14559 8139 14601 8181
rect 14859 8139 14901 8181
rect 15279 9459 15321 9501
rect 15459 11139 15501 11181
rect 15459 11019 15501 11061
rect 15819 11679 15861 11721
rect 15879 11619 15921 11661
rect 15819 11499 15861 11541
rect 15759 11319 15801 11361
rect 15819 11199 15861 11241
rect 15759 10959 15801 11001
rect 15639 10839 15681 10881
rect 15759 10839 15801 10881
rect 15519 10599 15561 10641
rect 15459 10539 15501 10581
rect 15579 10539 15621 10581
rect 15819 10779 15861 10821
rect 15459 10419 15501 10461
rect 15759 10419 15801 10461
rect 15399 10179 15441 10221
rect 15399 10059 15441 10101
rect 16899 13539 16941 13581
rect 16719 13359 16761 13401
rect 16779 13239 16821 13281
rect 16899 13239 16941 13281
rect 16899 13119 16941 13161
rect 16959 13059 17001 13101
rect 17259 14619 17301 14661
rect 17619 14859 17661 14901
rect 17319 14562 17361 14604
rect 17439 14562 17481 14604
rect 17259 14439 17301 14481
rect 17499 14436 17541 14478
rect 17379 14319 17421 14361
rect 17019 12999 17061 13041
rect 16599 12876 16641 12918
rect 16719 12876 16761 12918
rect 16839 12819 16881 12861
rect 16899 12819 16941 12861
rect 16659 12699 16701 12741
rect 16779 12699 16821 12741
rect 16539 12519 16581 12561
rect 16599 12399 16641 12441
rect 16419 12279 16461 12321
rect 16599 12159 16641 12201
rect 16719 12519 16761 12561
rect 16179 12036 16221 12078
rect 16119 11439 16161 11481
rect 15939 11259 15981 11301
rect 15879 10659 15921 10701
rect 15879 10596 15921 10638
rect 15879 10416 15921 10458
rect 15819 10239 15861 10281
rect 15759 10179 15801 10221
rect 15759 10116 15801 10158
rect 15639 9999 15681 10041
rect 15459 9876 15501 9918
rect 16059 11199 16101 11241
rect 16239 11559 16281 11601
rect 16419 11559 16461 11601
rect 16599 11559 16641 11601
rect 16479 11499 16521 11541
rect 16359 11442 16401 11484
rect 16539 11442 16581 11484
rect 16839 12219 16881 12261
rect 16839 12099 16881 12141
rect 17019 12879 17061 12921
rect 17019 12699 17061 12741
rect 16959 12639 17001 12681
rect 17139 13899 17181 13941
rect 17499 13899 17541 13941
rect 17139 13719 17181 13761
rect 17139 13479 17181 13521
rect 17499 13479 17541 13521
rect 17139 13299 17181 13341
rect 17439 13299 17481 13341
rect 17139 13179 17181 13221
rect 17319 13179 17361 13221
rect 17199 13059 17241 13101
rect 17319 13002 17361 13044
rect 17139 12879 17181 12921
rect 16779 11979 16821 12021
rect 16899 11619 16941 11661
rect 16779 11559 16821 11601
rect 16239 11199 16281 11241
rect 16539 11199 16581 11241
rect 16419 11139 16461 11181
rect 16299 10599 16341 10641
rect 16179 10539 16221 10581
rect 16119 10416 16161 10458
rect 16239 10299 16281 10341
rect 16179 10239 16221 10281
rect 15999 10119 16041 10161
rect 15939 9999 15981 10041
rect 15939 9882 15981 9924
rect 15399 9579 15441 9621
rect 15159 9339 15201 9381
rect 15219 9279 15261 9321
rect 15159 9159 15201 9201
rect 15099 8799 15141 8841
rect 15219 8739 15261 8781
rect 15099 8379 15141 8421
rect 15219 8319 15261 8361
rect 15159 8199 15201 8241
rect 14739 8019 14781 8061
rect 14859 8019 14901 8061
rect 14499 7479 14541 7521
rect 14619 7479 14661 7521
rect 14859 7899 14901 7941
rect 14799 7779 14841 7821
rect 14979 7659 15021 7701
rect 14919 7599 14961 7641
rect 14499 7359 14541 7401
rect 14139 7239 14181 7281
rect 13959 7119 14001 7161
rect 14139 6999 14181 7041
rect 13719 6762 13761 6804
rect 13899 6759 13941 6801
rect 13839 6630 13881 6672
rect 13779 6459 13821 6501
rect 13839 6399 13881 6441
rect 13839 6279 13881 6321
rect 14139 6279 14181 6321
rect 13779 6219 13821 6261
rect 13659 6039 13701 6081
rect 13599 5919 13641 5961
rect 14139 6099 14181 6141
rect 13839 6039 13881 6081
rect 13779 5859 13821 5901
rect 13659 5736 13701 5778
rect 13539 5619 13581 5661
rect 13419 5559 13461 5601
rect 13419 5439 13461 5481
rect 13539 5202 13581 5244
rect 13659 5619 13701 5661
rect 13239 5019 13281 5061
rect 13479 5019 13521 5061
rect 13539 4959 13581 5001
rect 14379 7296 14421 7338
rect 14259 7239 14301 7281
rect 14439 6999 14481 7041
rect 14439 6936 14481 6978
rect 14319 6762 14361 6804
rect 14619 6819 14661 6861
rect 14499 6762 14541 6804
rect 14559 6519 14601 6561
rect 14379 6459 14421 6501
rect 14499 6399 14541 6441
rect 14259 6159 14301 6201
rect 13899 5919 13941 5961
rect 14199 5919 14241 5961
rect 13959 5859 14001 5901
rect 14079 5862 14121 5904
rect 13899 5619 13941 5661
rect 13839 5559 13881 5601
rect 13899 5439 13941 5481
rect 13779 5259 13821 5301
rect 14079 5319 14121 5361
rect 13959 5259 14001 5301
rect 13776 5076 13818 5118
rect 13839 5079 13881 5121
rect 13659 4779 13701 4821
rect 13239 4479 13281 4521
rect 12999 4359 13041 4401
rect 13179 4359 13221 4401
rect 12819 4059 12861 4101
rect 13719 4359 13761 4401
rect 13599 4302 13641 4344
rect 13779 4299 13821 4341
rect 13299 4176 13341 4218
rect 13419 4179 13461 4221
rect 13659 4176 13701 4218
rect 13479 4119 13521 4161
rect 13179 4059 13221 4101
rect 12999 3819 13041 3861
rect 12699 3699 12741 3741
rect 12639 3639 12681 3681
rect 12819 3642 12861 3684
rect 12279 3399 12321 3441
rect 12579 3399 12621 3441
rect 12639 2919 12681 2961
rect 12999 3339 13041 3381
rect 13179 3516 13221 3558
rect 13299 3516 13341 3558
rect 13299 3399 13341 3441
rect 12879 3219 12921 3261
rect 13059 3219 13101 3261
rect 12999 3159 13041 3201
rect 12879 3039 12921 3081
rect 12759 2859 12801 2901
rect 12999 2859 13041 2901
rect 12459 2799 12501 2841
rect 12159 2742 12201 2784
rect 12339 2742 12381 2784
rect 11559 2616 11601 2658
rect 11679 2616 11721 2658
rect 11859 2619 11901 2661
rect 12579 2739 12621 2781
rect 12879 2739 12921 2781
rect 12039 2616 12081 2658
rect 12156 2616 12198 2658
rect 12279 2616 12321 2658
rect 12159 2439 12201 2481
rect 11379 2319 11421 2361
rect 12039 2259 12081 2301
rect 11559 2199 11601 2241
rect 11439 2082 11481 2124
rect 9399 1779 9441 1821
rect 10119 1779 10161 1821
rect 10359 1779 10401 1821
rect 10479 1779 10521 1821
rect 9339 1659 9381 1701
rect 10119 1659 10161 1701
rect 10119 1539 10161 1581
rect 11079 1539 11121 1581
rect 9579 1359 9621 1401
rect 9819 1359 9861 1401
rect 9039 1299 9081 1341
rect 9219 1299 9261 1341
rect 9159 1239 9201 1281
rect 9459 1239 9501 1281
rect 9639 1299 9681 1341
rect 9759 1239 9801 1281
rect 9699 1182 9741 1224
rect 8379 1119 8421 1161
rect 8919 1119 8961 1161
rect 7959 1059 8001 1101
rect 8079 1056 8121 1098
rect 8199 1056 8241 1098
rect 8559 1056 8601 1098
rect 8259 999 8301 1041
rect 8379 999 8421 1041
rect 8139 879 8181 921
rect 8019 639 8061 681
rect 7899 579 7941 621
rect 8499 939 8541 981
rect 8439 819 8481 861
rect 7839 396 7881 438
rect 8019 396 8061 438
rect 8199 396 8241 438
rect 7599 339 7641 381
rect 7719 339 7761 381
rect 8319 339 8361 381
rect 7359 279 7401 321
rect 9099 1056 9141 1098
rect 9219 999 9261 1041
rect 9399 999 9441 1041
rect 9699 1059 9741 1101
rect 9639 999 9681 1041
rect 9519 939 9561 981
rect 9699 939 9741 981
rect 9879 1239 9921 1281
rect 10419 1419 10461 1461
rect 11079 1419 11121 1461
rect 10239 1182 10281 1224
rect 10719 1359 10761 1401
rect 10599 1239 10641 1281
rect 10899 1239 10941 1281
rect 11199 1956 11241 1998
rect 11499 1956 11541 1998
rect 11979 1956 12021 1998
rect 11619 1839 11661 1881
rect 11739 1839 11781 1881
rect 11319 1359 11361 1401
rect 11439 1299 11481 1341
rect 11919 1299 11961 1341
rect 11139 1239 11181 1281
rect 11259 1182 11301 1224
rect 11559 1182 11601 1224
rect 11799 1182 11841 1224
rect 10179 1056 10221 1098
rect 10419 1056 10461 1098
rect 9939 939 9981 981
rect 10059 939 10101 981
rect 10299 939 10341 981
rect 9099 879 9141 921
rect 9759 879 9801 921
rect 8679 819 8721 861
rect 8799 579 8841 621
rect 9699 819 9741 861
rect 9819 819 9861 861
rect 9639 759 9681 801
rect 9759 759 9801 801
rect 8679 522 8721 564
rect 8919 519 8961 561
rect 9099 522 9141 564
rect 9219 522 9261 564
rect 9399 519 9441 561
rect 10539 879 10581 921
rect 10239 699 10281 741
rect 10119 639 10161 681
rect 10119 519 10161 561
rect 8499 396 8541 438
rect 8619 396 8661 438
rect 8739 396 8781 438
rect 8919 396 8961 438
rect 9459 459 9501 501
rect 9039 396 9081 438
rect 9159 396 9201 438
rect 9399 396 9441 438
rect 10899 1056 10941 1098
rect 11019 1056 11061 1098
rect 11079 999 11121 1041
rect 12099 1179 12141 1221
rect 10959 939 11001 981
rect 11259 939 11301 981
rect 10719 879 10761 921
rect 10659 819 10701 861
rect 10599 699 10641 741
rect 9579 396 9621 438
rect 9699 396 9741 438
rect 10179 399 10221 441
rect 8979 279 9021 321
rect 9459 279 9501 321
rect 9579 219 9621 261
rect 7239 159 7281 201
rect 8439 159 8481 201
rect 10539 399 10581 441
rect 10659 639 10701 681
rect 10659 519 10701 561
rect 10839 522 10881 564
rect 11499 999 11541 1041
rect 11979 1056 12021 1098
rect 11859 999 11901 1041
rect 11799 939 11841 981
rect 11379 759 11421 801
rect 11199 639 11241 681
rect 11499 639 11541 681
rect 12279 2319 12321 2361
rect 12219 2199 12261 2241
rect 12219 1956 12261 1998
rect 12579 2619 12621 2661
rect 12819 2616 12861 2658
rect 12999 2619 13041 2661
rect 12699 2559 12741 2601
rect 12939 2319 12981 2361
rect 12759 2259 12801 2301
rect 12399 2199 12441 2241
rect 12879 2139 12921 2181
rect 12579 2085 12621 2127
rect 12339 2019 12381 2061
rect 12279 1779 12321 1821
rect 12699 1959 12741 2001
rect 12459 1719 12501 1761
rect 12339 1539 12381 1581
rect 12459 1299 12501 1341
rect 13119 2919 13161 2961
rect 13119 2739 13161 2781
rect 13539 3699 13581 3741
rect 13479 3639 13521 3681
rect 13599 3516 13641 3558
rect 13356 3339 13398 3381
rect 13419 3339 13461 3381
rect 13179 2616 13221 2658
rect 13359 2379 13401 2421
rect 13479 3039 13521 3081
rect 13659 3159 13701 3201
rect 13479 2739 13521 2781
rect 14019 5079 14061 5121
rect 13959 4959 14001 5001
rect 13959 4719 14001 4761
rect 13899 4419 13941 4461
rect 14199 5739 14241 5781
rect 14139 5259 14181 5301
rect 14379 5862 14421 5904
rect 14859 7179 14901 7221
rect 14739 7119 14781 7161
rect 15339 9279 15381 9321
rect 16059 9756 16101 9798
rect 15699 9639 15741 9681
rect 15819 9639 15861 9681
rect 16119 9639 16161 9681
rect 15579 9519 15621 9561
rect 15459 9219 15501 9261
rect 15339 9039 15381 9081
rect 15399 8982 15441 9024
rect 15399 8799 15441 8841
rect 15339 8739 15381 8781
rect 15459 8679 15501 8721
rect 15399 8559 15441 8601
rect 15939 9519 15981 9561
rect 15579 9039 15621 9081
rect 15819 9039 15861 9081
rect 15999 9459 16041 9501
rect 16179 9519 16221 9561
rect 15939 8982 15981 9024
rect 16059 9399 16101 9441
rect 16479 10359 16521 10401
rect 16359 10239 16401 10281
rect 16299 10179 16341 10221
rect 16359 10119 16401 10161
rect 16299 9879 16341 9921
rect 17079 11979 17121 12021
rect 16959 11499 17001 11541
rect 16719 11319 16761 11361
rect 16659 10779 16701 10821
rect 16839 11316 16881 11358
rect 17259 12819 17301 12861
rect 17679 14799 17721 14841
rect 17679 13959 17721 14001
rect 18279 15039 18321 15081
rect 18219 14979 18261 15021
rect 18039 14739 18081 14781
rect 18279 14559 18321 14601
rect 18408 15519 18450 15561
rect 18399 14679 18441 14721
rect 18159 14259 18201 14301
rect 17739 13839 17781 13881
rect 18279 13959 18321 14001
rect 18399 13719 18441 13761
rect 17679 13659 17721 13701
rect 17799 13662 17841 13704
rect 17619 13479 17661 13521
rect 17739 13536 17781 13578
rect 17679 13419 17721 13461
rect 17859 13239 17901 13281
rect 17799 13119 17841 13161
rect 17739 13059 17781 13101
rect 17619 12999 17661 13041
rect 18219 13662 18261 13704
rect 18399 13656 18441 13698
rect 18159 13536 18201 13578
rect 18339 13539 18381 13581
rect 18279 13419 18321 13461
rect 17979 13359 18021 13401
rect 18279 13356 18321 13398
rect 18039 13239 18081 13281
rect 17919 12999 17961 13041
rect 18219 13119 18261 13161
rect 17679 12879 17721 12921
rect 17439 12759 17481 12801
rect 17259 12339 17301 12381
rect 17379 12339 17421 12381
rect 17379 12276 17421 12318
rect 17259 12219 17301 12261
rect 17199 12099 17241 12141
rect 17379 12102 17421 12144
rect 17199 11979 17241 12021
rect 17139 11496 17181 11538
rect 16959 11199 17001 11241
rect 16779 10959 16821 11001
rect 16719 10719 16761 10761
rect 16599 10539 16641 10581
rect 16659 10599 16701 10641
rect 16599 10419 16641 10461
rect 16539 10179 16581 10221
rect 16479 9942 16521 9984
rect 16719 10416 16761 10458
rect 16779 10359 16821 10401
rect 16659 10179 16701 10221
rect 16479 9879 16521 9921
rect 16419 9756 16461 9798
rect 16539 9756 16581 9798
rect 16299 9519 16341 9561
rect 16239 9219 16281 9261
rect 16179 9099 16221 9141
rect 15699 8856 15741 8898
rect 15579 8619 15621 8661
rect 15519 8499 15561 8541
rect 15519 8436 15561 8478
rect 15459 8379 15501 8421
rect 15699 8619 15741 8661
rect 15459 8196 15501 8238
rect 15279 8136 15321 8178
rect 15219 7779 15261 7821
rect 14979 7419 15021 7461
rect 15159 7479 15201 7521
rect 15219 7422 15261 7464
rect 14979 7299 15021 7341
rect 14919 7059 14961 7101
rect 14979 6999 15021 7041
rect 14919 6819 14961 6861
rect 14799 6279 14841 6321
rect 14619 6039 14661 6081
rect 14439 5736 14481 5778
rect 14499 5679 14541 5721
rect 14319 5499 14361 5541
rect 14259 5259 14301 5301
rect 15159 7296 15201 7338
rect 15279 7299 15321 7341
rect 15219 7179 15261 7221
rect 15159 6999 15201 7041
rect 15039 6819 15081 6861
rect 15579 8079 15621 8121
rect 16119 8979 16161 9021
rect 15939 8559 15981 8601
rect 15759 8439 15801 8481
rect 15759 8319 15801 8361
rect 15879 8322 15921 8364
rect 16059 8856 16101 8898
rect 16239 8859 16281 8901
rect 16239 8679 16281 8721
rect 16059 8619 16101 8661
rect 16179 8559 16221 8601
rect 16059 8316 16101 8358
rect 15399 7839 15441 7881
rect 15699 7839 15741 7881
rect 15939 8196 15981 8238
rect 15639 7659 15681 7701
rect 15519 7539 15561 7581
rect 15399 7419 15441 7461
rect 15339 7119 15381 7161
rect 15339 6999 15381 7041
rect 15279 6939 15321 6981
rect 15219 6819 15261 6861
rect 15099 6636 15141 6678
rect 15459 7296 15501 7338
rect 15459 6939 15501 6981
rect 16059 8079 16101 8121
rect 15999 7659 16041 7701
rect 16119 7659 16161 7701
rect 15759 7599 15801 7641
rect 15879 7422 15921 7464
rect 15999 7422 16041 7464
rect 16119 7419 16161 7461
rect 15819 7299 15861 7341
rect 15759 7239 15801 7281
rect 15759 7119 15801 7161
rect 15639 6819 15681 6861
rect 15279 6699 15321 6741
rect 15099 6519 15141 6561
rect 14679 5919 14721 5961
rect 14919 5919 14961 5961
rect 15039 5919 15081 5961
rect 14619 5439 14661 5481
rect 14799 5862 14841 5904
rect 14859 5739 14901 5781
rect 14799 5679 14841 5721
rect 14559 5259 14601 5301
rect 14499 5199 14541 5241
rect 14379 5076 14421 5118
rect 14499 5079 14541 5121
rect 14499 4659 14541 4701
rect 14259 4539 14301 4581
rect 14679 4479 14721 4521
rect 14079 4419 14121 4461
rect 14319 4299 14361 4341
rect 13899 4176 13941 4218
rect 14019 4176 14061 4218
rect 13839 4059 13881 4101
rect 14019 3999 14061 4041
rect 14139 3879 14181 3921
rect 14559 4302 14601 4344
rect 14919 5439 14961 5481
rect 15039 5439 15081 5481
rect 15399 6579 15441 6621
rect 15339 6279 15381 6321
rect 15219 6159 15261 6201
rect 15519 5979 15561 6021
rect 15279 5919 15321 5961
rect 15219 5859 15261 5901
rect 15579 5862 15621 5904
rect 15339 5736 15381 5778
rect 15159 5679 15201 5721
rect 15279 5679 15321 5721
rect 15639 5739 15681 5781
rect 15219 5499 15261 5541
rect 14919 5319 14961 5361
rect 14859 5199 14901 5241
rect 15159 5199 15201 5241
rect 14799 5019 14841 5061
rect 14739 4359 14781 4401
rect 15159 5079 15201 5121
rect 15099 5019 15141 5061
rect 14919 4899 14961 4941
rect 14859 4539 14901 4581
rect 15099 4539 15141 4581
rect 14859 4476 14901 4518
rect 14799 4299 14841 4341
rect 14379 4179 14421 4221
rect 14619 4176 14661 4218
rect 14799 4179 14841 4221
rect 14739 4059 14781 4101
rect 14379 3999 14421 4041
rect 14019 3642 14061 3684
rect 14139 3648 14181 3690
rect 14319 3648 14361 3690
rect 14439 3879 14481 3921
rect 14439 3639 14481 3681
rect 14439 3519 14481 3561
rect 14919 4359 14961 4401
rect 14859 4119 14901 4161
rect 14859 3999 14901 4041
rect 14679 3510 14721 3552
rect 14379 3399 14421 3441
rect 14016 3339 14058 3381
rect 14079 3339 14121 3381
rect 13899 3279 13941 3321
rect 13779 3099 13821 3141
rect 13839 2979 13881 3021
rect 13599 2616 13641 2658
rect 13719 2616 13761 2658
rect 14079 3219 14121 3261
rect 14259 3219 14301 3261
rect 14019 2859 14061 2901
rect 14139 2859 14181 2901
rect 13899 2742 13941 2784
rect 14019 2742 14061 2784
rect 14499 2979 14541 3021
rect 14319 2919 14361 2961
rect 13899 2619 13941 2661
rect 14079 2616 14121 2658
rect 14259 2619 14301 2661
rect 14619 2742 14661 2784
rect 13899 2499 13941 2541
rect 14319 2499 14361 2541
rect 14439 2499 14481 2541
rect 13839 2439 13881 2481
rect 13719 2319 13761 2361
rect 13419 2199 13461 2241
rect 13719 2199 13761 2241
rect 13059 2139 13101 2181
rect 13179 2082 13221 2124
rect 13359 2079 13401 2121
rect 13479 2082 13521 2124
rect 12939 1956 12981 1998
rect 13239 1956 13281 1998
rect 13419 1959 13461 2001
rect 13359 1839 13401 1881
rect 13539 1899 13581 1941
rect 13419 1719 13461 1761
rect 14199 2379 14241 2421
rect 14079 2139 14121 2181
rect 13959 1899 14001 1941
rect 13839 1839 13881 1881
rect 13779 1779 13821 1821
rect 13779 1659 13821 1701
rect 13719 1599 13761 1641
rect 13119 1539 13161 1581
rect 13479 1479 13521 1521
rect 12939 1419 12981 1461
rect 12339 1182 12381 1224
rect 12639 1182 12681 1224
rect 12759 1182 12801 1224
rect 12879 1182 12921 1224
rect 12159 939 12201 981
rect 12579 1056 12621 1098
rect 12699 1056 12741 1098
rect 12279 759 12321 801
rect 12099 639 12141 681
rect 10959 519 11001 561
rect 11319 522 11361 564
rect 11079 459 11121 501
rect 10899 396 10941 438
rect 10599 339 10641 381
rect 10779 339 10821 381
rect 11079 279 11121 321
rect 11379 396 11421 438
rect 12399 579 12441 621
rect 12279 522 12321 564
rect 12459 522 12501 564
rect 12639 522 12681 564
rect 12759 522 12801 564
rect 12099 396 12141 438
rect 12219 396 12261 438
rect 12579 396 12621 438
rect 12699 396 12741 438
rect 12339 279 12381 321
rect 12459 279 12501 321
rect 12639 279 12681 321
rect 12219 219 12261 261
rect 13059 1359 13101 1401
rect 13179 1239 13221 1281
rect 13299 1182 13341 1224
rect 12939 1059 12981 1101
rect 13599 1182 13641 1224
rect 14439 2319 14481 2361
rect 14319 2139 14361 2181
rect 14859 3459 14901 3501
rect 14859 3159 14901 3201
rect 14859 2979 14901 3021
rect 14799 2919 14841 2961
rect 14859 2859 14901 2901
rect 15219 4899 15261 4941
rect 15159 4359 15201 4401
rect 15039 4119 15081 4161
rect 15219 4179 15261 4221
rect 15159 4059 15201 4101
rect 15159 3639 15201 3681
rect 15039 3516 15081 3558
rect 14979 3159 15021 3201
rect 14919 2799 14961 2841
rect 15519 5559 15561 5601
rect 15339 5379 15381 5421
rect 15579 5499 15621 5541
rect 15759 6999 15801 7041
rect 16059 7296 16101 7338
rect 16539 9159 16581 9201
rect 16359 9099 16401 9141
rect 16299 8439 16341 8481
rect 16419 8979 16461 9021
rect 16719 10059 16761 10101
rect 16959 10299 17001 10341
rect 16899 10059 16941 10101
rect 16839 9999 16881 10041
rect 16719 9879 16761 9921
rect 16959 9882 17001 9924
rect 16719 9759 16761 9801
rect 16659 9519 16701 9561
rect 16899 9639 16941 9681
rect 17439 11979 17481 12021
rect 17319 11859 17361 11901
rect 17379 11619 17421 11661
rect 17319 11559 17361 11601
rect 17199 11439 17241 11481
rect 17619 12819 17661 12861
rect 17559 12759 17601 12801
rect 17499 11799 17541 11841
rect 17499 11559 17541 11601
rect 17379 11316 17421 11358
rect 17319 11259 17361 11301
rect 17199 10839 17241 10881
rect 17139 10779 17181 10821
rect 17379 10719 17421 10761
rect 17079 10539 17121 10581
rect 17199 10542 17241 10584
rect 17319 10542 17361 10584
rect 17439 10539 17481 10581
rect 17079 10419 17121 10461
rect 17259 10416 17301 10458
rect 17379 10416 17421 10458
rect 17139 10239 17181 10281
rect 17319 10239 17361 10281
rect 17139 10119 17181 10161
rect 17259 10119 17301 10161
rect 17139 9999 17181 10041
rect 17259 9939 17301 9981
rect 17199 9882 17241 9924
rect 17379 9879 17421 9921
rect 17079 9699 17121 9741
rect 16779 9579 16821 9621
rect 16719 9399 16761 9441
rect 16659 9279 16701 9321
rect 16719 9219 16761 9261
rect 16659 9159 16701 9201
rect 16599 8979 16641 9021
rect 16839 8979 16881 9021
rect 16659 8856 16701 8898
rect 16779 8799 16821 8841
rect 16959 9519 17001 9561
rect 17379 9759 17421 9801
rect 17319 9699 17361 9741
rect 17259 9459 17301 9501
rect 17259 9279 17301 9321
rect 17079 8982 17121 9024
rect 16899 8859 16941 8901
rect 16599 8619 16641 8661
rect 16839 8619 16881 8661
rect 17139 8856 17181 8898
rect 16419 8499 16461 8541
rect 16659 8499 16701 8541
rect 16839 8499 16881 8541
rect 16359 8379 16401 8421
rect 16419 8322 16461 8364
rect 16659 8376 16701 8418
rect 16839 8379 16881 8421
rect 16239 8199 16281 8241
rect 16479 8196 16521 8238
rect 16359 7899 16401 7941
rect 16659 8196 16701 8238
rect 16899 8199 16941 8241
rect 16779 8139 16821 8181
rect 16779 7959 16821 8001
rect 16299 7599 16341 7641
rect 16239 7419 16281 7461
rect 16479 7479 16521 7521
rect 16599 7659 16641 7701
rect 16539 7419 16581 7461
rect 16659 7479 16701 7521
rect 15936 7239 15978 7281
rect 15999 7239 16041 7281
rect 15879 7059 15921 7101
rect 15819 6939 15861 6981
rect 16059 6999 16101 7041
rect 15999 6759 16041 6801
rect 15819 6519 15861 6561
rect 15759 6219 15801 6261
rect 15699 5319 15741 5361
rect 15459 4959 15501 5001
rect 15519 4659 15561 4701
rect 15399 4539 15441 4581
rect 15339 4419 15381 4461
rect 15639 5079 15681 5121
rect 15579 4599 15621 4641
rect 15579 4419 15621 4461
rect 15519 4302 15561 4344
rect 15339 4179 15381 4221
rect 15459 3759 15501 3801
rect 15879 6159 15921 6201
rect 15999 6639 16041 6681
rect 16356 7296 16398 7338
rect 16419 7299 16461 7341
rect 16599 7299 16641 7341
rect 17739 12819 17781 12861
rect 17679 12459 17721 12501
rect 17919 12879 17961 12921
rect 17859 12699 17901 12741
rect 17859 12339 17901 12381
rect 17739 12099 17781 12141
rect 17919 12099 17961 12141
rect 17619 11979 17661 12021
rect 17619 11859 17661 11901
rect 17799 11859 17841 11901
rect 17919 11799 17961 11841
rect 17679 11559 17721 11601
rect 17799 11559 17841 11601
rect 17559 11499 17601 11541
rect 17679 11442 17721 11484
rect 17859 11439 17901 11481
rect 17559 11199 17601 11241
rect 17739 11199 17781 11241
rect 17619 10959 17661 11001
rect 17559 10839 17601 10881
rect 17499 10239 17541 10281
rect 17799 10779 17841 10821
rect 17679 10659 17721 10701
rect 17619 10539 17661 10581
rect 17859 10539 17901 10581
rect 17619 10419 17661 10461
rect 17559 10119 17601 10161
rect 17799 10359 17841 10401
rect 17739 10299 17781 10341
rect 17499 9999 17541 10041
rect 17619 9999 17661 10041
rect 17439 9699 17481 9741
rect 17379 9519 17421 9561
rect 17379 9159 17421 9201
rect 17319 8979 17361 9021
rect 17679 9939 17721 9981
rect 17796 9939 17838 9981
rect 17859 9939 17901 9981
rect 17619 9699 17661 9741
rect 17679 9639 17721 9681
rect 17619 9519 17661 9561
rect 17559 9339 17601 9381
rect 17499 8979 17541 9021
rect 17319 8859 17361 8901
rect 17259 8679 17301 8721
rect 17139 8499 17181 8541
rect 17499 8859 17541 8901
rect 17859 9759 17901 9801
rect 17799 9699 17841 9741
rect 17739 9579 17781 9621
rect 17679 9339 17721 9381
rect 17679 9276 17721 9318
rect 17619 9099 17661 9141
rect 17799 9159 17841 9201
rect 17739 9039 17781 9081
rect 17859 8979 17901 9021
rect 17679 8799 17721 8841
rect 17559 8739 17601 8781
rect 17619 8559 17661 8601
rect 17379 8439 17421 8481
rect 17499 8439 17541 8481
rect 17319 8379 17361 8421
rect 17859 8859 17901 8901
rect 17799 8739 17841 8781
rect 17739 8559 17781 8601
rect 17559 8322 17601 8364
rect 17679 8319 17721 8361
rect 16959 7959 17001 8001
rect 16899 7479 16941 7521
rect 17079 8139 17121 8181
rect 17259 7719 17301 7761
rect 17079 7479 17121 7521
rect 16839 7296 16881 7338
rect 16659 7239 16701 7281
rect 16779 7239 16821 7281
rect 16479 7059 16521 7101
rect 16419 6999 16461 7041
rect 17019 7299 17061 7341
rect 16959 7179 17001 7221
rect 16779 6999 16821 7041
rect 16959 6999 17001 7041
rect 16299 6762 16341 6804
rect 16719 6939 16761 6981
rect 16719 6819 16761 6861
rect 16539 6762 16581 6804
rect 16659 6762 16701 6804
rect 16779 6762 16821 6804
rect 16359 6636 16401 6678
rect 16119 6519 16161 6561
rect 16119 6279 16161 6321
rect 16059 6219 16101 6261
rect 15816 5859 15858 5901
rect 15879 5862 15921 5904
rect 15999 5862 16041 5904
rect 16719 6636 16761 6678
rect 16779 6579 16821 6621
rect 16539 6519 16581 6561
rect 16299 6459 16341 6501
rect 16239 6339 16281 6381
rect 16179 6159 16221 6201
rect 16179 5979 16221 6021
rect 16059 5736 16101 5778
rect 15819 5679 15861 5721
rect 16119 5499 16161 5541
rect 15939 5379 15981 5421
rect 16719 6279 16761 6321
rect 16719 6159 16761 6201
rect 16359 6039 16401 6081
rect 16299 5859 16341 5901
rect 16599 5919 16641 5961
rect 16479 5862 16521 5904
rect 16659 5859 16701 5901
rect 16236 5739 16278 5781
rect 16779 5919 16821 5961
rect 16959 6459 17001 6501
rect 17199 7479 17241 7521
rect 17439 8199 17481 8241
rect 17319 7599 17361 7641
rect 17619 8196 17661 8238
rect 17439 7899 17481 7941
rect 17739 7839 17781 7881
rect 17619 7779 17661 7821
rect 17499 7659 17541 7701
rect 17139 7419 17181 7461
rect 17379 7479 17421 7521
rect 17079 7239 17121 7281
rect 17199 7239 17241 7281
rect 17139 7179 17181 7221
rect 17379 7296 17421 7338
rect 17559 7479 17601 7521
rect 17319 6759 17361 6801
rect 17499 7296 17541 7338
rect 17499 7179 17541 7221
rect 17739 7719 17781 7761
rect 17859 8559 17901 8601
rect 17859 8379 17901 8421
rect 18099 12699 18141 12741
rect 18099 12339 18141 12381
rect 18039 12099 18081 12141
rect 18339 13239 18381 13281
rect 18279 12219 18321 12261
rect 18219 12099 18261 12141
rect 18399 12159 18441 12201
rect 18159 11976 18201 12018
rect 18099 11919 18141 11961
rect 18039 11619 18081 11661
rect 18159 11739 18201 11781
rect 18279 11739 18321 11781
rect 17979 11439 18021 11481
rect 18099 11499 18141 11541
rect 18219 11619 18261 11661
rect 18159 11439 18201 11481
rect 18039 11019 18081 11061
rect 18159 11319 18201 11361
rect 18099 10899 18141 10941
rect 18279 11499 18321 11541
rect 18399 11859 18441 11901
rect 18399 11739 18441 11781
rect 18339 11019 18381 11061
rect 18279 10959 18321 11001
rect 18339 10899 18381 10941
rect 18279 10779 18321 10821
rect 18219 10659 18261 10701
rect 18099 10599 18141 10641
rect 17979 10539 18021 10581
rect 18339 10539 18381 10581
rect 18039 10119 18081 10161
rect 18219 10416 18261 10458
rect 18159 9999 18201 10041
rect 18339 9999 18381 10041
rect 18099 9939 18141 9981
rect 18039 9879 18081 9921
rect 18039 9759 18081 9801
rect 17979 9639 18021 9681
rect 17979 9459 18021 9501
rect 18099 9699 18141 9741
rect 18279 9699 18321 9741
rect 18219 9459 18261 9501
rect 18099 9159 18141 9201
rect 18159 9099 18201 9141
rect 18039 8979 18081 9021
rect 18339 9579 18381 9621
rect 18339 9459 18381 9501
rect 18279 9039 18321 9081
rect 18399 9159 18441 9201
rect 18399 9039 18441 9081
rect 18039 8859 18081 8901
rect 17979 8799 18021 8841
rect 18219 8856 18261 8898
rect 18399 8856 18441 8898
rect 18279 8799 18321 8841
rect 18099 8679 18141 8721
rect 18039 8439 18081 8481
rect 18159 8439 18201 8481
rect 17979 8379 18021 8421
rect 17799 7479 17841 7521
rect 18039 8196 18081 8238
rect 18039 7959 18081 8001
rect 18039 7839 18081 7881
rect 17979 7719 18021 7761
rect 18219 7959 18261 8001
rect 18159 7719 18201 7761
rect 18159 7599 18201 7641
rect 17979 7419 18021 7461
rect 18219 7419 18261 7461
rect 17619 7299 17661 7341
rect 17559 6939 17601 6981
rect 17799 7296 17841 7338
rect 17919 7299 17961 7341
rect 17979 7299 18021 7341
rect 17679 7179 17721 7221
rect 17919 7059 17961 7101
rect 17739 6939 17781 6981
rect 17859 6939 17901 6981
rect 17199 6519 17241 6561
rect 17319 6339 17361 6381
rect 17019 6159 17061 6201
rect 17319 6039 17361 6081
rect 16899 5979 16941 6021
rect 17019 5979 17061 6021
rect 16959 5862 17001 5904
rect 17199 5862 17241 5904
rect 16779 5799 16821 5841
rect 16299 5736 16341 5778
rect 16419 5736 16461 5778
rect 16539 5736 16581 5778
rect 16719 5736 16761 5778
rect 15759 5199 15801 5241
rect 15939 5259 15981 5301
rect 16179 5256 16221 5298
rect 16359 5679 16401 5721
rect 16839 5739 16881 5781
rect 16419 5619 16461 5661
rect 16776 5619 16818 5661
rect 16359 5559 16401 5601
rect 16299 5199 16341 5241
rect 15699 4779 15741 4821
rect 15879 4959 15921 5001
rect 15819 4839 15861 4881
rect 15819 4599 15861 4641
rect 15939 4599 15981 4641
rect 15696 4299 15738 4341
rect 15759 4299 15801 4341
rect 15399 3519 15441 3561
rect 15339 3219 15381 3261
rect 15279 2979 15321 3021
rect 15156 2796 15198 2838
rect 15219 2799 15261 2841
rect 14979 2742 15021 2784
rect 15099 2739 15141 2781
rect 14919 2616 14961 2658
rect 15099 2616 15141 2658
rect 15099 2499 15141 2541
rect 14919 2139 14961 2181
rect 14556 2079 14598 2121
rect 14619 2082 14661 2124
rect 14799 2082 14841 2124
rect 14499 1956 14541 1998
rect 14439 1899 14481 1941
rect 14199 1719 14241 1761
rect 14139 1239 14181 1281
rect 14319 1188 14361 1230
rect 13239 999 13281 1041
rect 13119 939 13161 981
rect 13059 759 13101 801
rect 12939 519 12981 561
rect 13179 522 13221 564
rect 13299 522 13341 564
rect 13119 396 13161 438
rect 12939 339 12981 381
rect 13239 339 13281 381
rect 13659 1056 13701 1098
rect 13779 1050 13821 1092
rect 15099 2079 15141 2121
rect 14619 1899 14661 1941
rect 14559 1188 14601 1230
rect 14439 999 14481 1041
rect 14019 939 14061 981
rect 14499 639 14541 681
rect 13659 522 13701 564
rect 13899 522 13941 564
rect 13479 396 13521 438
rect 14739 759 14781 801
rect 14919 1839 14961 1881
rect 14979 1719 15021 1761
rect 15039 1659 15081 1701
rect 14919 1419 14961 1461
rect 15459 3219 15501 3261
rect 15459 2919 15501 2961
rect 15336 2799 15378 2841
rect 15399 2799 15441 2841
rect 15219 2736 15261 2778
rect 15879 4059 15921 4101
rect 15936 3642 15978 3684
rect 16119 5079 16161 5121
rect 16059 5019 16101 5061
rect 16119 4479 16161 4521
rect 16059 4299 16101 4341
rect 16299 4599 16341 4641
rect 16239 4479 16281 4521
rect 16839 5616 16881 5658
rect 17019 5736 17061 5778
rect 17139 5619 17181 5661
rect 17439 6639 17481 6681
rect 17379 5919 17421 5961
rect 17559 6279 17601 6321
rect 17559 5919 17601 5961
rect 17619 5859 17661 5901
rect 17259 5739 17301 5781
rect 17379 5679 17421 5721
rect 17199 5559 17241 5601
rect 16899 5499 16941 5541
rect 17079 5499 17121 5541
rect 16899 5379 16941 5421
rect 16479 5319 16521 5361
rect 16839 5319 16881 5361
rect 16539 5202 16581 5244
rect 16659 5202 16701 5244
rect 16779 5202 16821 5244
rect 16959 5142 17001 5184
rect 16419 5019 16461 5061
rect 16419 4839 16461 4881
rect 16359 4419 16401 4461
rect 16719 5019 16761 5061
rect 17013 5019 17055 5061
rect 16599 4899 16641 4941
rect 16179 4359 16221 4401
rect 16479 4359 16521 4401
rect 16239 4302 16281 4344
rect 17619 5679 17661 5721
rect 17559 5619 17601 5661
rect 17739 6759 17781 6801
rect 18039 7179 18081 7221
rect 18219 7299 18261 7341
rect 18159 7179 18201 7221
rect 18099 7119 18141 7161
rect 18039 6939 18081 6981
rect 17979 6819 18021 6861
rect 18039 6759 18081 6801
rect 17739 6639 17781 6681
rect 17799 6159 17841 6201
rect 17859 6039 17901 6081
rect 17739 5859 17781 5901
rect 18039 6639 18081 6681
rect 18159 6939 18201 6981
rect 18159 6819 18201 6861
rect 18099 6039 18141 6081
rect 17799 5736 17841 5778
rect 17919 5619 17961 5661
rect 17739 5499 17781 5541
rect 17859 5499 17901 5541
rect 17439 5439 17481 5481
rect 17559 5439 17601 5481
rect 17679 5439 17721 5481
rect 17919 5439 17961 5481
rect 17139 5259 17181 5301
rect 17919 5199 17961 5241
rect 17559 5136 17601 5178
rect 17859 5139 17901 5181
rect 17979 5139 18021 5181
rect 18339 8739 18381 8781
rect 18279 7179 18321 7221
rect 18279 7059 18321 7101
rect 18219 5736 18261 5778
rect 17139 5019 17181 5061
rect 17919 4959 17961 5001
rect 17079 4899 17121 4941
rect 17139 4719 17181 4761
rect 17139 4539 17181 4581
rect 16779 4359 16821 4401
rect 17859 4539 17901 4581
rect 17799 4419 17841 4461
rect 16419 4236 16461 4278
rect 16599 4236 16641 4278
rect 16719 4236 16761 4278
rect 15999 3639 16041 3681
rect 15759 3459 15801 3501
rect 15921 3459 15963 3501
rect 15819 3399 15861 3441
rect 15639 3099 15681 3141
rect 15579 2859 15621 2901
rect 15519 2616 15561 2658
rect 16179 4176 16221 4218
rect 16239 3759 16281 3801
rect 16479 4179 16521 4221
rect 16419 4059 16461 4101
rect 16419 3819 16461 3861
rect 16119 3639 16161 3681
rect 16359 3639 16401 3681
rect 16119 3519 16161 3561
rect 16299 3516 16341 3558
rect 16419 3519 16461 3561
rect 15879 3339 15921 3381
rect 16059 3339 16101 3381
rect 16599 4119 16641 4161
rect 16659 4059 16701 4101
rect 16599 3879 16641 3921
rect 17199 4242 17241 4284
rect 17559 4236 17601 4278
rect 16779 4119 16821 4161
rect 16719 3939 16761 3981
rect 17019 3939 17061 3981
rect 17139 3939 17181 3981
rect 16659 3819 16701 3861
rect 16539 3642 16581 3684
rect 16659 3642 16701 3684
rect 17079 3879 17121 3921
rect 17079 3639 17121 3681
rect 17859 3999 17901 4041
rect 18099 5019 18141 5061
rect 18219 4539 18261 4581
rect 18159 4419 18201 4461
rect 18039 4302 18081 4344
rect 18099 4176 18141 4218
rect 17919 3939 17961 3981
rect 17559 3879 17601 3921
rect 18039 3999 18081 4041
rect 16839 3582 16881 3624
rect 17019 3582 17061 3624
rect 17139 3582 17181 3624
rect 16599 3516 16641 3558
rect 16539 3459 16581 3501
rect 17979 3639 18021 3681
rect 18159 3639 18201 3681
rect 18399 8559 18441 8601
rect 18399 7779 18441 7821
rect 18399 7599 18441 7641
rect 18399 7059 18441 7101
rect 18339 6939 18381 6981
rect 18279 3819 18321 3861
rect 17619 3576 17661 3618
rect 17919 3579 17961 3621
rect 18039 3579 18081 3621
rect 16539 3339 16581 3381
rect 16359 3099 16401 3141
rect 16479 3099 16521 3141
rect 16179 2979 16221 3021
rect 16299 2979 16341 3021
rect 16479 2979 16521 3021
rect 15879 2859 15921 2901
rect 15999 2859 16041 2901
rect 15879 2742 15921 2784
rect 16059 2799 16101 2841
rect 15999 2739 16041 2781
rect 16419 2679 16461 2721
rect 15639 2616 15681 2658
rect 15819 2616 15861 2658
rect 15279 2379 15321 2421
rect 15699 2379 15741 2421
rect 15219 2199 15261 2241
rect 15399 2199 15441 2241
rect 15279 2139 15321 2181
rect 15819 2319 15861 2361
rect 15819 2199 15861 2241
rect 16059 2619 16101 2661
rect 16239 2616 16281 2658
rect 16359 2559 16401 2601
rect 15819 2082 15861 2124
rect 15939 2082 15981 2124
rect 16179 2082 16221 2124
rect 16299 2082 16341 2124
rect 16419 2082 16461 2124
rect 15339 1956 15381 1998
rect 15159 1899 15201 1941
rect 15159 1299 15201 1341
rect 15099 1239 15141 1281
rect 15279 1182 15321 1224
rect 15759 1956 15801 1998
rect 15639 1839 15681 1881
rect 16119 1899 16161 1941
rect 15759 1779 15801 1821
rect 16359 1719 16401 1761
rect 16779 3279 16821 3321
rect 16659 2799 16701 2841
rect 17199 3459 17241 3501
rect 18279 3459 18321 3501
rect 17139 3399 17181 3441
rect 18027 3399 18069 3441
rect 18159 3339 18201 3381
rect 17559 3219 17601 3261
rect 17799 3219 17841 3261
rect 17139 2979 17181 3021
rect 17439 2979 17481 3021
rect 17559 2979 17601 3021
rect 17139 2859 17181 2901
rect 16539 2379 16581 2421
rect 16839 2559 16881 2601
rect 16656 2199 16698 2241
rect 16719 2199 16761 2241
rect 16899 2259 16941 2301
rect 16839 2199 16881 2241
rect 17079 2739 17121 2781
rect 17199 2559 17241 2601
rect 17139 2259 17181 2301
rect 16839 2079 16881 2121
rect 16599 1956 16641 1998
rect 16719 1779 16761 1821
rect 16479 1659 16521 1701
rect 15459 1479 15501 1521
rect 16119 1479 16161 1521
rect 16239 1479 16281 1521
rect 16959 2139 17001 2181
rect 17259 2139 17301 2181
rect 17019 1959 17061 2001
rect 16959 1779 17001 1821
rect 17139 1659 17181 1701
rect 17079 1599 17121 1641
rect 15459 1299 15501 1341
rect 15099 1056 15141 1098
rect 15219 999 15261 1041
rect 15399 999 15441 1041
rect 15579 1182 15621 1224
rect 16779 1419 16821 1461
rect 16659 1359 16701 1401
rect 16299 1239 16341 1281
rect 16479 1239 16521 1281
rect 16839 1239 16881 1281
rect 17079 1179 17121 1221
rect 16779 1119 16821 1161
rect 15039 759 15081 801
rect 15459 759 15501 801
rect 15579 759 15621 801
rect 14859 639 14901 681
rect 14739 528 14781 570
rect 15039 522 15081 564
rect 15759 1050 15801 1092
rect 15639 639 15681 681
rect 16119 639 16161 681
rect 15879 528 15921 570
rect 17019 1050 17061 1092
rect 16119 522 16161 564
rect 16539 522 16581 564
rect 16779 522 16821 564
rect 17319 1899 17361 1941
rect 17319 1599 17361 1641
rect 17199 1359 17241 1401
rect 17319 1479 17361 1521
rect 17379 1419 17421 1461
rect 17559 2859 17601 2901
rect 17739 2379 17781 2421
rect 17619 1719 17661 1761
rect 18099 3099 18141 3141
rect 17979 2979 18021 3021
rect 17979 2742 18021 2784
rect 17919 2082 17961 2124
rect 17979 1899 18021 1941
rect 17799 1599 17841 1641
rect 18039 1479 18081 1521
rect 17799 1299 17841 1341
rect 17439 1239 17481 1281
rect 17619 1239 17661 1281
rect 17319 1056 17361 1098
rect 17139 879 17181 921
rect 17319 879 17361 921
rect 17439 879 17481 921
rect 17919 1182 17961 1224
rect 17619 1056 17661 1098
rect 17739 1056 17781 1098
rect 17859 939 17901 981
rect 18099 1056 18141 1098
rect 18039 939 18081 981
rect 18219 1299 18261 1341
rect 17919 819 17961 861
rect 18159 819 18201 861
rect 13299 279 13341 321
rect 12039 159 12081 201
rect 12879 159 12921 201
rect 13599 159 13641 201
rect 2259 99 2301 141
rect 3999 99 4041 141
rect 6399 99 6441 141
rect 8319 99 8361 141
rect 8559 99 8601 141
rect 10179 99 10221 141
rect 10359 99 10401 141
rect 11259 99 11301 141
rect 14199 390 14241 432
rect 14379 390 14421 432
rect 14496 390 14538 432
rect 14559 390 14601 432
rect 15339 390 15381 432
rect 15519 390 15561 432
rect 15639 390 15681 432
rect 17559 396 17601 438
rect 17799 396 17841 438
rect 18399 3339 18441 3381
rect 18399 3219 18441 3261
rect 18339 1479 18381 1521
rect 18279 1182 18321 1224
rect 18399 879 18441 921
<< metal3 >>
rect 10041 18768 11619 18792
rect 14601 18768 15579 18792
rect 17601 18768 18219 18792
rect 10641 18708 11559 18732
rect 11601 18708 13119 18732
rect 13341 18708 14892 18732
rect 921 18648 1959 18672
rect 2001 18648 2739 18672
rect 13101 18648 14799 18672
rect 14868 18672 14892 18708
rect 15261 18708 15339 18732
rect 15408 18708 16959 18732
rect 15408 18672 15432 18708
rect 14868 18648 15432 18672
rect 17721 18648 17999 18672
rect 2301 18588 4299 18612
rect 4341 18588 5979 18612
rect 6021 18588 6219 18612
rect 6741 18588 7152 18612
rect 7128 18561 7152 18588
rect 9621 18588 9759 18612
rect 9801 18588 10599 18612
rect 13161 18588 14859 18612
rect 14901 18588 15999 18612
rect 1581 18528 2199 18552
rect 6141 18528 6759 18552
rect 7161 18528 7419 18552
rect 9321 18528 10119 18552
rect 16881 18528 17499 18552
rect 321 18468 759 18492
rect 801 18468 1179 18492
rect 2661 18468 3279 18492
rect 3621 18468 4119 18492
rect 5001 18468 5319 18492
rect 5361 18468 5619 18492
rect 8361 18468 8559 18492
rect 11181 18468 11439 18492
rect 11721 18468 12039 18492
rect 12921 18468 13179 18492
rect 13221 18468 14379 18492
rect 14421 18468 14919 18492
rect 15861 18468 16779 18492
rect 16941 18468 17472 18492
rect 17448 18441 17472 18468
rect 1821 18408 2259 18432
rect 2421 18408 2559 18432
rect 9921 18408 9999 18432
rect 15081 18408 15639 18432
rect 16341 18408 16419 18432
rect 16581 18408 16659 18432
rect 17481 18408 17799 18432
rect 561 18351 639 18375
rect 768 18348 876 18372
rect 768 18312 792 18348
rect 981 18351 1059 18375
rect 1581 18348 1932 18372
rect 708 18288 792 18312
rect 1908 18312 1932 18348
rect 2901 18351 3039 18375
rect 3441 18348 3699 18372
rect 4248 18348 4419 18372
rect 1908 18288 2052 18312
rect 708 18258 732 18288
rect 861 18228 939 18252
rect 1281 18225 1419 18249
rect 2028 18258 2052 18288
rect 1821 18228 1899 18252
rect 2088 18252 2112 18342
rect 2508 18288 2619 18312
rect 2088 18228 2319 18252
rect 2508 18252 2532 18288
rect 2481 18228 2532 18252
rect 2841 18228 3339 18252
rect 4008 18252 4032 18342
rect 3708 18228 4032 18252
rect 3708 18192 3732 18228
rect 2601 18168 3732 18192
rect 3801 18168 3999 18192
rect 4248 18192 4272 18348
rect 4581 18351 4719 18375
rect 5241 18351 5439 18375
rect 5781 18351 5859 18375
rect 6381 18351 6519 18375
rect 7401 18351 7719 18375
rect 8241 18351 8319 18375
rect 8901 18348 9099 18372
rect 4341 18225 4479 18249
rect 5061 18225 5139 18249
rect 5181 18228 5379 18252
rect 5781 18225 6279 18249
rect 6561 18228 6759 18252
rect 6828 18252 6852 18339
rect 6828 18228 7059 18252
rect 7101 18228 7539 18252
rect 8448 18252 8472 18342
rect 10401 18351 10479 18375
rect 10761 18351 10839 18375
rect 11001 18348 11319 18372
rect 11361 18351 11676 18375
rect 11781 18351 11859 18375
rect 12021 18351 12099 18375
rect 12321 18348 12396 18372
rect 12501 18351 12579 18375
rect 12741 18348 13059 18372
rect 11028 18288 11892 18312
rect 8181 18228 8472 18252
rect 9141 18225 9219 18249
rect 9681 18228 9879 18252
rect 11028 18258 11052 18288
rect 11721 18228 11799 18252
rect 11868 18252 11892 18288
rect 11868 18228 12759 18252
rect 4041 18168 4272 18192
rect 5961 18168 6099 18192
rect 11961 18168 12039 18192
rect 12441 18168 12699 18192
rect 13008 18192 13032 18348
rect 13521 18348 13659 18372
rect 14541 18351 14679 18375
rect 15108 18348 15399 18372
rect 15108 18258 15132 18348
rect 16608 18348 16779 18372
rect 16188 18261 16212 18342
rect 16488 18261 16512 18342
rect 16608 18312 16632 18348
rect 13401 18225 13539 18249
rect 13701 18225 14439 18249
rect 15381 18228 15519 18252
rect 15681 18228 15879 18252
rect 16161 18228 16212 18261
rect 16161 18219 16200 18228
rect 16461 18228 16512 18261
rect 16548 18288 16632 18312
rect 17208 18312 17232 18342
rect 17208 18288 17379 18312
rect 16548 18258 16572 18288
rect 16461 18219 16500 18228
rect 16761 18228 17139 18252
rect 12921 18168 13032 18192
rect 15321 18168 15579 18192
rect 17301 18168 17859 18192
rect 1641 18108 1899 18132
rect 2361 18108 4479 18132
rect 4521 18108 5499 18132
rect 5541 18108 8139 18132
rect 8181 18108 8259 18132
rect 9021 18108 10179 18132
rect 10221 18108 10359 18132
rect 10941 18108 11139 18132
rect 12681 18108 12819 18132
rect 13221 18108 13476 18132
rect 13581 18108 13719 18132
rect 13761 18108 14019 18132
rect 14841 18108 15339 18132
rect 15681 18108 16239 18132
rect 17001 18108 17199 18132
rect 2421 18048 2919 18072
rect 2961 18048 4179 18072
rect 5241 18048 5859 18072
rect 11361 18048 12459 18072
rect 12501 18048 12999 18072
rect 13041 18048 15459 18072
rect 15501 18048 16419 18072
rect 1821 17988 2559 18012
rect 4101 17988 4719 18012
rect 6201 17988 10659 18012
rect 11421 17988 12579 18012
rect 12741 17988 12996 18012
rect 13101 17988 13299 18012
rect 14421 17988 14559 18012
rect 14721 17988 15639 18012
rect 16161 17988 16239 18012
rect 17301 17988 17379 18012
rect 17421 17988 17919 18012
rect 2001 17928 2379 17952
rect 3081 17928 3579 17952
rect 3621 17928 4239 17952
rect 10521 17928 10719 17952
rect 10761 17928 11259 17952
rect 11301 17928 13419 17952
rect 13941 17928 14199 17952
rect 14241 17928 14979 17952
rect 17241 17928 17379 17952
rect 17421 17928 17799 17952
rect 1161 17868 1899 17892
rect 5361 17868 5619 17892
rect 6441 17868 7299 17892
rect 12621 17868 13359 17892
rect 14181 17868 14319 17892
rect 14448 17868 15339 17892
rect 3021 17808 3219 17832
rect 4221 17808 4899 17832
rect 5721 17808 6339 17832
rect 7701 17808 7899 17832
rect 7941 17808 8499 17832
rect 9861 17808 10059 17832
rect 11961 17808 12099 17832
rect 12141 17808 12399 17832
rect 12441 17808 13332 17832
rect 381 17748 1179 17772
rect 13308 17781 13332 17808
rect 13521 17808 13599 17832
rect 14448 17832 14472 17868
rect 16641 17868 16959 17892
rect 17601 17868 18339 17892
rect 13881 17808 14472 17832
rect 14541 17808 14739 17832
rect 14781 17808 15759 17832
rect 16521 17808 17079 17832
rect 17841 17808 18099 17832
rect 1221 17748 1659 17772
rect 3408 17748 3699 17772
rect 3408 17724 3432 17748
rect 8961 17748 9459 17772
rect 9501 17748 10092 17772
rect 468 17592 492 17682
rect 681 17688 819 17712
rect 1041 17691 1179 17715
rect 1341 17688 1479 17712
rect 2241 17688 2439 17712
rect 2481 17688 2679 17712
rect 3201 17691 3399 17715
rect 3921 17691 4179 17715
rect 4701 17691 4839 17715
rect 5661 17691 5979 17715
rect 6801 17688 7059 17712
rect 7101 17688 7359 17712
rect 2808 17652 2832 17682
rect 5028 17652 5052 17682
rect 5448 17652 5472 17682
rect 7401 17688 7572 17712
rect 2808 17628 3012 17652
rect 5028 17628 5472 17652
rect 468 17568 879 17592
rect 1281 17568 1599 17592
rect 1641 17568 1692 17592
rect 1041 17508 1179 17532
rect 1668 17532 1692 17568
rect 1761 17565 1839 17589
rect 2988 17592 3012 17628
rect 5448 17601 5472 17628
rect 2988 17568 3639 17592
rect 3681 17568 3939 17592
rect 4281 17568 4419 17592
rect 4821 17568 5079 17592
rect 5421 17568 5472 17601
rect 5421 17559 5460 17568
rect 5541 17568 5919 17592
rect 6081 17568 6339 17592
rect 7161 17568 7419 17592
rect 7548 17592 7572 17688
rect 7641 17691 7719 17715
rect 8061 17688 8139 17712
rect 9141 17688 9492 17712
rect 7548 17568 7839 17592
rect 8001 17568 8319 17592
rect 8979 17589 9021 17619
rect 8661 17565 9399 17589
rect 9468 17592 9492 17688
rect 9621 17688 9972 17712
rect 9948 17598 9972 17688
rect 10068 17712 10092 17748
rect 10581 17748 10692 17772
rect 10068 17688 10119 17712
rect 10668 17712 10692 17748
rect 10881 17748 11019 17772
rect 12801 17748 12879 17772
rect 13161 17748 13272 17772
rect 10668 17688 11079 17712
rect 9468 17568 9519 17592
rect 1668 17508 2139 17532
rect 2781 17508 3099 17532
rect 4161 17508 6159 17532
rect 10008 17535 10032 17682
rect 10368 17592 10392 17682
rect 12441 17688 12612 17712
rect 10548 17628 11019 17652
rect 10548 17598 10572 17628
rect 12288 17652 12312 17682
rect 12288 17640 12549 17652
rect 12288 17628 12561 17640
rect 12519 17601 12561 17628
rect 10101 17568 10392 17592
rect 10701 17568 10899 17592
rect 11121 17565 11379 17589
rect 11781 17568 12219 17592
rect 12558 17580 12561 17601
rect 12588 17598 12612 17688
rect 13248 17712 13272 17748
rect 13341 17748 14859 17772
rect 13248 17688 13839 17712
rect 12648 17592 12672 17682
rect 14061 17712 14100 17721
rect 14220 17712 14259 17721
rect 14061 17679 14112 17712
rect 12648 17568 12819 17592
rect 14088 17598 14112 17679
rect 14208 17679 14259 17712
rect 14421 17688 14592 17712
rect 14208 17598 14232 17679
rect 14568 17598 14592 17688
rect 14661 17688 14799 17712
rect 15108 17601 15132 17682
rect 15381 17712 15420 17721
rect 15381 17679 15432 17712
rect 15501 17688 15612 17712
rect 13041 17565 13119 17589
rect 13461 17565 13539 17589
rect 13821 17565 13899 17589
rect 14361 17565 14439 17589
rect 15081 17568 15132 17601
rect 15408 17598 15432 17679
rect 15081 17559 15120 17568
rect 15588 17592 15612 17688
rect 15681 17688 15852 17712
rect 15828 17598 15852 17688
rect 15981 17691 16119 17715
rect 16461 17691 16599 17715
rect 17148 17688 17499 17712
rect 15588 17568 15699 17592
rect 16221 17568 16659 17592
rect 16728 17592 16752 17682
rect 17148 17598 17172 17688
rect 17868 17652 17892 17682
rect 17628 17640 17892 17652
rect 17619 17628 17892 17640
rect 17619 17601 17661 17628
rect 16728 17568 17019 17592
rect 17961 17568 18099 17592
rect 18141 17568 18279 17592
rect 10008 17499 10059 17535
rect 11901 17508 12039 17532
rect 15321 17508 15519 17532
rect 17721 17508 17859 17532
rect 321 17448 579 17472
rect 621 17448 1119 17472
rect 1461 17448 1659 17472
rect 1701 17448 1839 17472
rect 3801 17448 4059 17472
rect 4701 17448 5619 17472
rect 5661 17448 6819 17472
rect 7581 17448 8739 17472
rect 9621 17448 10179 17472
rect 10221 17448 10659 17472
rect 12261 17448 13239 17472
rect 13281 17448 14439 17472
rect 15621 17448 15879 17472
rect 16461 17448 17559 17472
rect 2181 17388 2319 17412
rect 8241 17388 8559 17412
rect 9741 17388 10239 17412
rect 11421 17388 12339 17412
rect 12381 17388 12819 17412
rect 13161 17388 14772 17412
rect 561 17328 759 17352
rect 2148 17352 2172 17379
rect 801 17328 2172 17352
rect 3861 17328 4599 17352
rect 4641 17328 5739 17352
rect 9861 17328 10419 17352
rect 10821 17328 10959 17352
rect 11001 17328 11559 17352
rect 11601 17328 12159 17352
rect 14748 17352 14772 17388
rect 17061 17388 17439 17412
rect 14748 17328 15339 17352
rect 15501 17328 16359 17352
rect 9201 17268 9279 17292
rect 9321 17268 9699 17292
rect 10821 17268 11379 17292
rect 11841 17268 12099 17292
rect 15321 17268 15579 17292
rect 16581 17268 17139 17292
rect 5241 17208 5379 17232
rect 5421 17208 6699 17232
rect 10041 17208 11679 17232
rect 14481 17208 14859 17232
rect 14901 17208 15459 17232
rect 15921 17208 16692 17232
rect 501 17148 1419 17172
rect 1461 17148 1839 17172
rect 5301 17148 5739 17172
rect 7281 17148 8499 17172
rect 10161 17148 11079 17172
rect 11601 17148 12699 17172
rect 12741 17148 14199 17172
rect 15741 17148 16419 17172
rect 16668 17172 16692 17208
rect 16668 17148 18372 17172
rect 18348 17121 18372 17148
rect 921 17088 2439 17112
rect 5841 17088 8559 17112
rect 8601 17088 8739 17112
rect 9081 17088 11859 17112
rect 12021 17088 13779 17112
rect 14601 17088 15399 17112
rect 15801 17088 15939 17112
rect 16401 17088 16599 17112
rect 16641 17088 17259 17112
rect 17301 17088 17559 17112
rect 18348 17088 18399 17121
rect 18360 17079 18399 17088
rect 3321 17028 3459 17052
rect 5361 17028 5979 17052
rect 9741 17028 11799 17052
rect 13281 17028 13659 17052
rect 14481 17028 14799 17052
rect 15261 17028 15579 17052
rect 16881 17028 17139 17052
rect 17181 17028 17799 17052
rect 681 16968 819 16992
rect 2601 16968 3759 16992
rect 7341 16968 8079 16992
rect 10101 16968 10299 16992
rect 10581 16968 11019 16992
rect 15228 16992 15252 17019
rect 12081 16968 15252 16992
rect 15501 16968 15819 16992
rect 1761 16908 1899 16932
rect 2421 16908 3099 16932
rect 7488 16908 7779 16932
rect 7488 16881 7512 16908
rect 7908 16908 8259 16932
rect 321 16848 612 16872
rect 261 16788 519 16812
rect 588 16692 612 16848
rect 3441 16848 3699 16872
rect 4881 16848 5379 16872
rect 5568 16848 5859 16872
rect 741 16791 879 16815
rect 1008 16752 1032 16782
rect 1221 16812 1260 16821
rect 1221 16779 1272 16812
rect 1341 16791 1599 16815
rect 1641 16788 2019 16812
rect 2481 16788 2739 16812
rect 3501 16791 3579 16815
rect 4461 16788 4719 16812
rect 4761 16788 4959 16812
rect 1008 16728 1152 16752
rect 1128 16701 1152 16728
rect 588 16668 639 16692
rect 921 16668 1059 16692
rect 1128 16668 1179 16701
rect 1140 16659 1179 16668
rect 1248 16692 1272 16779
rect 2388 16728 2559 16752
rect 1248 16668 1839 16692
rect 2388 16698 2412 16728
rect 2181 16668 2259 16692
rect 3261 16668 3399 16692
rect 3768 16692 3792 16779
rect 3681 16668 3792 16692
rect 3948 16692 3972 16782
rect 5568 16812 5592 16848
rect 6399 16848 6699 16872
rect 6399 16824 6441 16848
rect 6741 16848 6852 16872
rect 5541 16788 5592 16812
rect 5661 16791 5799 16815
rect 6201 16788 6399 16812
rect 6561 16791 6639 16815
rect 6828 16812 6852 16848
rect 7221 16848 7479 16872
rect 7908 16872 7932 16908
rect 9321 16908 9399 16932
rect 9441 16908 9759 16932
rect 12141 16908 13119 16932
rect 13581 16908 14079 16932
rect 14541 16908 15072 16932
rect 7701 16848 7932 16872
rect 15048 16872 15072 16908
rect 15381 16908 15879 16932
rect 17541 16908 17619 16932
rect 17661 16908 17979 16932
rect 15048 16848 15159 16872
rect 15201 16848 15699 16872
rect 6828 16788 6999 16812
rect 7401 16791 7599 16815
rect 8001 16788 8052 16812
rect 5808 16752 5832 16782
rect 4188 16728 5832 16752
rect 4188 16692 4212 16728
rect 8028 16701 8052 16788
rect 8901 16791 8979 16815
rect 9561 16791 9819 16815
rect 8199 16752 8241 16779
rect 8199 16740 8352 16752
rect 8208 16728 8352 16740
rect 3948 16668 4212 16692
rect 4641 16668 4779 16692
rect 5001 16665 5139 16689
rect 5601 16668 5739 16692
rect 6501 16668 6759 16692
rect 8328 16698 8352 16728
rect 8388 16641 8412 16782
rect 9861 16791 9999 16815
rect 11421 16788 11499 16812
rect 9681 16668 9912 16692
rect 1461 16608 1599 16632
rect 5901 16608 6339 16632
rect 6981 16608 7179 16632
rect 8661 16608 8859 16632
rect 9888 16632 9912 16668
rect 10428 16692 10452 16782
rect 10668 16752 10692 16782
rect 11088 16752 11112 16782
rect 10668 16740 10752 16752
rect 10908 16740 11112 16752
rect 10668 16728 10761 16740
rect 9981 16668 10452 16692
rect 10719 16701 10761 16728
rect 10899 16728 11112 16740
rect 10899 16701 10941 16728
rect 11628 16701 11652 16779
rect 11808 16701 11832 16782
rect 12321 16791 12399 16815
rect 12861 16791 12939 16815
rect 13341 16791 13419 16815
rect 14268 16788 14319 16812
rect 12048 16701 12072 16779
rect 11061 16668 11556 16692
rect 11808 16668 11859 16701
rect 11820 16659 11859 16668
rect 12588 16692 12612 16782
rect 12588 16668 12999 16692
rect 13068 16692 13092 16782
rect 13908 16701 13932 16782
rect 13068 16668 13479 16692
rect 13908 16668 13959 16701
rect 13920 16659 13959 16668
rect 9888 16608 10299 16632
rect 10428 16608 10659 16632
rect 141 16548 399 16572
rect 2661 16548 2799 16572
rect 2841 16548 3999 16572
rect 4041 16548 4179 16572
rect 4521 16548 5079 16572
rect 6501 16548 6699 16572
rect 6861 16548 6939 16572
rect 6981 16548 7059 16572
rect 9081 16548 9159 16572
rect 10428 16572 10452 16608
rect 12561 16608 12759 16632
rect 14268 16632 14292 16788
rect 15108 16788 15459 16812
rect 14748 16752 14772 16779
rect 15108 16752 15132 16788
rect 15861 16788 16212 16812
rect 14448 16740 15132 16752
rect 14439 16728 15132 16740
rect 16188 16752 16212 16788
rect 16581 16788 16719 16812
rect 16800 16812 16839 16821
rect 16788 16779 16839 16812
rect 17448 16788 17499 16812
rect 16188 16728 16272 16752
rect 14439 16701 14481 16728
rect 14841 16668 15219 16692
rect 15381 16665 15639 16689
rect 16248 16692 16272 16728
rect 16788 16698 16812 16779
rect 17028 16701 17052 16779
rect 16248 16668 16479 16692
rect 17268 16692 17292 16782
rect 17268 16668 17379 16692
rect 13881 16608 14292 16632
rect 16581 16608 16719 16632
rect 17448 16632 17472 16788
rect 17601 16668 17799 16692
rect 18081 16668 18219 16692
rect 17241 16608 17472 16632
rect 10041 16548 10452 16572
rect 11001 16548 11559 16572
rect 12021 16548 12099 16572
rect 12261 16548 13119 16572
rect 13161 16548 13299 16572
rect 13341 16548 13779 16572
rect 13941 16548 14499 16572
rect 15141 16548 15579 16572
rect 16341 16548 17499 16572
rect 17661 16548 17859 16572
rect 4401 16488 4899 16512
rect 5181 16488 5679 16512
rect 5841 16488 6399 16512
rect 6621 16488 6759 16512
rect 6801 16488 7179 16512
rect 7881 16488 8799 16512
rect 9561 16488 10416 16512
rect 10521 16488 10899 16512
rect 11061 16488 11619 16512
rect 13401 16488 13599 16512
rect 14121 16488 14316 16512
rect 14421 16488 14559 16512
rect 15081 16488 15459 16512
rect 15981 16488 16239 16512
rect 321 16428 399 16452
rect 1101 16428 1179 16452
rect 1221 16428 1359 16452
rect 1401 16428 1959 16452
rect 5121 16428 7299 16452
rect 9441 16428 9699 16452
rect 10101 16428 10179 16452
rect 621 16368 879 16392
rect 4101 16368 4356 16392
rect 4461 16368 5856 16392
rect 5961 16368 6939 16392
rect 8001 16368 8412 16392
rect 201 16308 759 16332
rect 3021 16308 3339 16332
rect 6081 16308 6639 16332
rect 8388 16332 8412 16368
rect 8661 16368 8979 16392
rect 9021 16368 9099 16392
rect 9261 16368 10059 16392
rect 10188 16392 10212 16419
rect 10521 16428 10719 16452
rect 10761 16428 11319 16452
rect 11781 16428 12459 16452
rect 12681 16428 13899 16452
rect 14061 16428 14739 16452
rect 15621 16428 16512 16452
rect 16488 16401 16512 16428
rect 16821 16428 16959 16452
rect 18021 16428 18279 16452
rect 10188 16368 10599 16392
rect 10641 16368 10779 16392
rect 11241 16368 11679 16392
rect 14361 16368 14556 16392
rect 14661 16368 15219 16392
rect 15741 16368 15999 16392
rect 16521 16368 17439 16392
rect 8388 16308 8559 16332
rect 9681 16308 9819 16332
rect 10941 16308 11799 16332
rect 11961 16308 12219 16332
rect 12648 16308 13179 16332
rect 921 16248 1239 16272
rect 1701 16248 2259 16272
rect 2301 16248 2499 16272
rect 2781 16248 3519 16272
rect 5301 16248 5379 16272
rect 6861 16248 7059 16272
rect 7821 16248 8139 16272
rect 9621 16248 10599 16272
rect 12648 16272 12672 16308
rect 13641 16308 14139 16332
rect 15501 16308 18099 16332
rect 18141 16308 18279 16332
rect 18321 16308 18552 16332
rect 12321 16248 12672 16272
rect 13281 16248 13839 16272
rect 14301 16248 14496 16272
rect 14601 16248 15039 16272
rect 15801 16248 15996 16272
rect 16101 16248 16599 16272
rect 16941 16248 17079 16272
rect 17241 16248 17859 16272
rect 681 16188 819 16212
rect 1761 16188 1839 16212
rect 1881 16188 2019 16212
rect 7641 16188 7839 16212
rect 9441 16188 9519 16212
rect 9921 16188 10119 16212
rect 10281 16212 10320 16221
rect 10281 16179 10332 16212
rect 15621 16188 15699 16212
rect 15861 16188 16179 16212
rect 17301 16188 17379 16212
rect 81 16131 399 16155
rect 1248 16128 1539 16152
rect 681 16005 819 16029
rect 1248 15981 1272 16128
rect 2181 16128 2319 16152
rect 2661 16128 2772 16152
rect 2748 16092 2772 16128
rect 2841 16131 2919 16155
rect 3081 16128 3219 16152
rect 3588 16128 3819 16152
rect 2748 16068 2892 16092
rect 1761 16005 1839 16029
rect 2001 16005 2259 16029
rect 2868 16032 2892 16068
rect 3588 16038 3612 16128
rect 3981 16128 4179 16152
rect 4701 16128 4899 16152
rect 4941 16128 5259 16152
rect 5541 16128 5619 16152
rect 5661 16131 5739 16155
rect 6081 16131 6159 16155
rect 7521 16128 7632 16152
rect 2868 16008 2979 16032
rect 501 15948 579 15972
rect 1848 15972 1872 15996
rect 1848 15948 2439 15972
rect 5421 15948 5619 15972
rect 6828 15972 6852 16119
rect 6948 16092 6972 16122
rect 6888 16080 6972 16092
rect 6879 16068 6972 16080
rect 6879 16041 6921 16068
rect 7281 16008 7359 16032
rect 7608 16032 7632 16128
rect 8028 16038 8052 16179
rect 8181 16131 8259 16155
rect 8688 16041 8712 16122
rect 9141 16128 9552 16152
rect 9528 16092 9552 16128
rect 10308 16152 10332 16179
rect 10308 16128 10392 16152
rect 9528 16080 9792 16092
rect 9528 16068 9801 16080
rect 9759 16041 9801 16068
rect 7608 16008 7899 16032
rect 8481 16005 8559 16029
rect 8661 16008 8712 16041
rect 8661 15999 8700 16008
rect 8901 16008 9099 16032
rect 9501 16008 9579 16032
rect 10008 16032 10032 16119
rect 9981 16008 10032 16032
rect 10161 16005 10239 16029
rect 10368 15981 10392 16128
rect 10488 16038 10512 16179
rect 10641 16128 10752 16152
rect 10728 16038 10752 16128
rect 10821 16128 11139 16152
rect 11301 16128 11436 16152
rect 11541 16128 11772 16152
rect 11748 16092 11772 16128
rect 11841 16128 12432 16152
rect 11748 16080 12369 16092
rect 11748 16068 12381 16080
rect 12339 16041 12381 16068
rect 10881 16008 11736 16032
rect 11841 16005 12039 16029
rect 12378 16020 12381 16041
rect 12408 16038 12432 16128
rect 12621 16128 13299 16152
rect 13341 16128 13479 16152
rect 13701 16128 13752 16152
rect 13728 16092 13752 16128
rect 13821 16131 14379 16155
rect 14661 16131 14859 16155
rect 15108 16128 15399 16152
rect 13728 16068 13992 16092
rect 12561 16008 12759 16032
rect 12981 16008 13119 16032
rect 13968 16038 13992 16068
rect 14988 16041 15012 16119
rect 13521 16005 13599 16029
rect 15108 15981 15132 16128
rect 16101 16128 16212 16152
rect 15528 16032 15552 16119
rect 15321 16008 15552 16032
rect 15648 16032 15672 16119
rect 16188 16092 16212 16128
rect 16680 16152 16719 16161
rect 16341 16128 16572 16152
rect 16188 16068 16272 16092
rect 15648 16008 15759 16032
rect 16248 16038 16272 16068
rect 16548 16038 16572 16128
rect 16668 16119 16719 16152
rect 16668 16038 16692 16119
rect 16041 16008 16119 16032
rect 16968 16032 16992 16122
rect 18300 16152 18339 16161
rect 18288 16119 18339 16152
rect 16968 16008 17199 16032
rect 17508 16032 17532 16119
rect 18288 16041 18312 16119
rect 17481 16008 17532 16032
rect 17601 16008 17799 16032
rect 18288 16008 18339 16041
rect 18300 15999 18339 16008
rect 6828 15948 6939 15972
rect 8361 15948 8739 15972
rect 10341 15948 10392 15981
rect 10341 15939 10380 15948
rect 12921 15948 14139 15972
rect 14181 15948 14259 15972
rect 14421 15948 14919 15972
rect 15081 15948 15132 15981
rect 15081 15939 15120 15948
rect 588 15912 612 15939
rect 588 15888 1179 15912
rect 2121 15888 2559 15912
rect 2961 15888 3099 15912
rect 3261 15888 3879 15912
rect 5481 15888 5799 15912
rect 6261 15888 6459 15912
rect 6501 15888 6999 15912
rect 7341 15888 7719 15912
rect 8328 15912 8352 15939
rect 8001 15888 8352 15912
rect 10308 15912 10332 15939
rect 10308 15888 10839 15912
rect 11481 15888 11979 15912
rect 12261 15888 12639 15912
rect 13101 15888 13359 15912
rect 14268 15888 14619 15912
rect 321 15828 936 15852
rect 1041 15828 1599 15852
rect 3501 15828 3759 15852
rect 6861 15828 7419 15852
rect 8661 15828 9279 15852
rect 9321 15828 9639 15852
rect 9681 15828 11919 15852
rect 14268 15852 14292 15888
rect 14661 15888 15099 15912
rect 16521 15888 17019 15912
rect 17481 15888 17679 15912
rect 13281 15828 14292 15852
rect 15261 15828 15639 15852
rect 16281 15828 17139 15852
rect 17421 15828 18039 15852
rect 18201 15828 18633 15852
rect 1341 15768 4419 15792
rect 4761 15768 5319 15792
rect 5361 15768 6039 15792
rect 6201 15768 6339 15792
rect 6741 15768 7656 15792
rect 7761 15768 7839 15792
rect 7881 15768 8412 15792
rect 1308 15732 1332 15759
rect 81 15708 1332 15732
rect 1701 15708 2799 15732
rect 3441 15708 3699 15732
rect 4521 15708 4959 15732
rect 5001 15708 5736 15732
rect 5841 15708 6579 15732
rect 6921 15708 6999 15732
rect 8388 15732 8412 15768
rect 8721 15768 8799 15792
rect 10401 15768 11199 15792
rect 11781 15768 12699 15792
rect 13461 15768 14679 15792
rect 14961 15768 15159 15792
rect 15348 15768 17259 15792
rect 8388 15708 9039 15732
rect 9561 15708 9639 15732
rect 10041 15708 10479 15732
rect 10521 15708 11139 15732
rect 11661 15708 11799 15732
rect 11961 15708 12999 15732
rect 15348 15732 15372 15768
rect 13521 15708 15372 15732
rect 15441 15708 16239 15732
rect 17361 15708 17619 15732
rect 621 15648 1059 15672
rect 6081 15648 6219 15672
rect 8361 15648 9159 15672
rect 10101 15648 11319 15672
rect 12141 15648 12459 15672
rect 13161 15648 13359 15672
rect 14001 15648 14199 15672
rect 14241 15648 14919 15672
rect 15201 15648 15939 15672
rect 16161 15648 18159 15672
rect 1581 15588 2079 15612
rect 3321 15588 3519 15612
rect 4641 15588 5619 15612
rect 5781 15588 6459 15612
rect 7881 15588 8139 15612
rect 8781 15588 9759 15612
rect 10221 15588 10539 15612
rect 12561 15588 12879 15612
rect 13041 15588 13539 15612
rect 14781 15588 15219 15612
rect 15801 15588 16539 15612
rect 16581 15588 17199 15612
rect 17241 15588 18099 15612
rect 4221 15528 6219 15552
rect 6441 15528 6579 15552
rect 7821 15528 8259 15552
rect 8961 15528 9039 15552
rect 10641 15528 10899 15552
rect 11901 15528 12099 15552
rect 12801 15528 13659 15552
rect 14361 15528 15012 15552
rect 14988 15501 15012 15528
rect 15141 15528 16116 15552
rect 16221 15528 17019 15552
rect 18450 15528 18633 15552
rect 2361 15468 2919 15492
rect 3321 15468 4119 15492
rect 4401 15468 4839 15492
rect 7581 15468 8019 15492
rect 8961 15468 9339 15492
rect 9501 15468 10299 15492
rect 11181 15468 11439 15492
rect 12081 15468 12399 15492
rect 12621 15468 13719 15492
rect 13941 15468 14799 15492
rect 15021 15468 15339 15492
rect 16401 15468 16779 15492
rect 321 15408 999 15432
rect 1401 15408 1659 15432
rect 9861 15408 10659 15432
rect 10821 15408 11679 15432
rect 12381 15408 12459 15432
rect 12501 15408 13239 15432
rect 17061 15408 17559 15432
rect 3501 15348 4059 15372
rect 5301 15348 6339 15372
rect 6381 15348 6612 15372
rect 1101 15288 2019 15312
rect 3921 15288 3999 15312
rect 4461 15288 4599 15312
rect 6588 15312 6612 15348
rect 7581 15348 7719 15372
rect 7941 15348 8079 15372
rect 11121 15348 11319 15372
rect 11541 15348 11859 15372
rect 12000 15372 12039 15381
rect 11988 15339 12039 15372
rect 12198 15339 12201 15360
rect 12261 15348 12672 15372
rect 6588 15288 7059 15312
rect 7221 15288 7839 15312
rect 201 15231 399 15255
rect 441 15228 759 15252
rect 921 15231 1539 15255
rect 2181 15231 2259 15255
rect 2481 15228 2619 15252
rect 2688 15228 3279 15252
rect 2688 15192 2712 15228
rect 4281 15231 4359 15255
rect 4881 15231 4959 15255
rect 5001 15228 5259 15252
rect 5478 15219 5481 15240
rect 5781 15231 5859 15255
rect 6501 15228 6912 15252
rect 5439 15192 5481 15219
rect 2508 15168 2712 15192
rect 5268 15180 5481 15192
rect 5268 15168 5469 15180
rect 2508 15138 2532 15168
rect 141 15105 459 15129
rect 501 15108 699 15132
rect 4101 15108 4779 15132
rect 5268 15132 5292 15168
rect 5241 15108 5292 15132
rect 5508 15132 5532 15222
rect 6888 15141 6912 15228
rect 7668 15192 7692 15222
rect 7041 15168 7692 15192
rect 5361 15108 5532 15132
rect 5721 15108 6159 15132
rect 7728 15138 7752 15288
rect 8388 15288 8499 15312
rect 7881 15228 8079 15252
rect 8388 15192 8412 15288
rect 11988 15312 12012 15339
rect 10701 15288 12012 15312
rect 12159 15312 12201 15339
rect 12159 15300 12279 15312
rect 12165 15288 12279 15300
rect 12441 15288 12612 15312
rect 8481 15228 8919 15252
rect 9921 15228 10179 15252
rect 9048 15192 9072 15222
rect 10461 15228 10779 15252
rect 11388 15228 11619 15252
rect 11208 15192 11232 15222
rect 8388 15168 8472 15192
rect 9048 15168 9252 15192
rect 7401 15105 7479 15129
rect 7761 15108 8139 15132
rect 8448 15081 8472 15168
rect 8781 15108 8979 15132
rect 9228 15132 9252 15168
rect 11088 15168 11232 15192
rect 9228 15108 9279 15132
rect 9561 15105 9819 15129
rect 10101 15105 10479 15129
rect 10521 15108 10599 15132
rect 11088 15132 11112 15168
rect 10881 15108 11112 15132
rect 11388 15132 11412 15228
rect 11841 15252 11880 15261
rect 11841 15219 11892 15252
rect 11181 15108 11412 15132
rect 11868 15132 11892 15219
rect 12348 15141 12372 15222
rect 11868 15108 12039 15132
rect 12348 15108 12399 15141
rect 12360 15099 12399 15108
rect 12588 15132 12612 15288
rect 12648 15252 12672 15348
rect 13701 15348 14499 15372
rect 15021 15348 15519 15372
rect 16461 15348 16839 15372
rect 16881 15348 17979 15372
rect 18021 15348 18279 15372
rect 12741 15288 13032 15312
rect 13008 15252 13032 15288
rect 13281 15288 13761 15312
rect 13719 15264 13761 15288
rect 14481 15288 14739 15312
rect 15501 15288 15579 15312
rect 17508 15288 17679 15312
rect 12648 15228 12732 15252
rect 13008 15228 13476 15252
rect 12708 15192 12732 15228
rect 13068 15192 13092 15228
rect 13581 15228 13632 15252
rect 12708 15168 13032 15192
rect 13068 15168 13152 15192
rect 13008 15141 13032 15168
rect 12588 15108 12699 15132
rect 12741 15108 12939 15132
rect 13008 15108 13059 15141
rect 13020 15099 13059 15108
rect 13128 15132 13152 15168
rect 13608 15141 13632 15228
rect 13761 15228 14079 15252
rect 13128 15108 13479 15132
rect 14181 15108 14439 15132
rect 14628 15132 14652 15222
rect 15528 15228 15759 15252
rect 15288 15141 15312 15219
rect 14628 15108 14979 15132
rect 15528 15138 15552 15228
rect 15921 15231 16056 15255
rect 16161 15231 16239 15255
rect 16320 15252 16359 15261
rect 16308 15219 16359 15252
rect 16788 15228 17139 15252
rect 16308 15138 16332 15219
rect 16488 15132 16512 15219
rect 16788 15192 16812 15228
rect 17508 15252 17532 15288
rect 17721 15288 17919 15312
rect 17181 15228 17532 15252
rect 17601 15228 17952 15252
rect 16728 15168 16812 15192
rect 16728 15138 16752 15168
rect 17928 15138 17952 15228
rect 18141 15231 18219 15255
rect 16488 15108 16599 15132
rect 16881 15105 17079 15129
rect 381 15048 1059 15072
rect 2121 15048 2319 15072
rect 2661 15048 2979 15072
rect 3681 15048 3759 15072
rect 3921 15048 3999 15072
rect 4041 15048 4419 15072
rect 5421 15048 5559 15072
rect 5781 15048 5859 15072
rect 7101 15048 7239 15072
rect 9201 15048 9939 15072
rect 10941 15048 11019 15072
rect 11601 15048 11676 15072
rect 11781 15048 12219 15072
rect 13341 15048 13899 15072
rect 14241 15048 14319 15072
rect 15201 15048 15459 15072
rect 17841 15048 18279 15072
rect 1521 14988 1899 15012
rect 4761 14988 5019 15012
rect 5061 14988 5259 15012
rect 6141 14988 6579 15012
rect 10521 14988 11139 15012
rect 11748 15012 11772 15039
rect 11421 14988 11772 15012
rect 12381 14988 12639 15012
rect 14601 14988 15912 15012
rect 861 14928 1299 14952
rect 2781 14928 3192 14952
rect 1281 14868 1539 14892
rect 1761 14868 2259 14892
rect 2301 14868 2376 14892
rect 2481 14868 2859 14892
rect 3168 14892 3192 14928
rect 3261 14928 3519 14952
rect 4821 14928 5319 14952
rect 5961 14928 6399 14952
rect 6441 14928 6759 14952
rect 7281 14928 8799 14952
rect 9921 14928 10419 14952
rect 10701 14928 10779 14952
rect 11001 14928 11259 14952
rect 11481 14928 12039 14952
rect 12081 14928 12279 14952
rect 12321 14928 12819 14952
rect 13161 14928 13359 14952
rect 13401 14928 14019 14952
rect 14241 14928 14499 14952
rect 14901 14928 15639 14952
rect 15888 14952 15912 14988
rect 15981 14988 16239 15012
rect 17241 14988 17499 15012
rect 17661 14988 17739 15012
rect 17781 14988 18219 15012
rect 15888 14928 15999 14952
rect 16161 14928 16299 14952
rect 17001 14928 17139 14952
rect 3168 14868 5199 14892
rect 6921 14868 8499 14892
rect 8541 14868 8859 14892
rect 8901 14868 9159 14892
rect 9681 14868 10179 14892
rect 12621 14868 12699 14892
rect 12981 14868 13659 14892
rect 14028 14892 14052 14919
rect 14028 14868 14139 14892
rect 15441 14868 16059 14892
rect 17121 14868 17259 14892
rect 17481 14868 17619 14892
rect 3081 14808 3819 14832
rect 4401 14808 5139 14832
rect 9561 14808 9879 14832
rect 10461 14808 11319 14832
rect 11361 14808 11439 14832
rect 12441 14808 12879 14832
rect 13881 14808 14199 14832
rect 14361 14808 14979 14832
rect 16161 14808 16779 14832
rect 17421 14808 17679 14832
rect 3981 14748 4959 14772
rect 7221 14748 7419 14772
rect 7461 14748 7536 14772
rect 7641 14748 7779 14772
rect 9441 14748 10179 14772
rect 10401 14748 11379 14772
rect 11841 14748 11979 14772
rect 12201 14748 12339 14772
rect 12621 14748 13899 14772
rect 15141 14748 15339 14772
rect 18081 14748 18372 14772
rect 18348 14721 18372 14748
rect 1221 14688 1479 14712
rect 4701 14688 5079 14712
rect 5121 14688 5439 14712
rect 6261 14688 6459 14712
rect 7101 14688 7299 14712
rect 7881 14688 8379 14712
rect 8541 14688 8979 14712
rect 9021 14688 9159 14712
rect 9621 14688 9939 14712
rect 10341 14688 11739 14712
rect 12561 14688 13179 14712
rect 13701 14688 13959 14712
rect 14841 14688 15999 14712
rect 16941 14688 17139 14712
rect 18348 14688 18399 14721
rect 18360 14679 18399 14688
rect 561 14628 699 14652
rect 741 14628 1659 14652
rect 1701 14628 2079 14652
rect 2928 14628 3039 14652
rect 381 14568 492 14592
rect 468 14481 492 14568
rect 861 14568 939 14592
rect 1161 14571 1419 14595
rect 1728 14568 1779 14592
rect 1728 14532 1752 14568
rect 2241 14568 2559 14592
rect 2928 14532 2952 14628
rect 7821 14628 8052 14652
rect 3321 14571 3339 14595
rect 3381 14571 3399 14595
rect 3621 14568 3939 14592
rect 4101 14571 4239 14595
rect 4821 14568 4959 14592
rect 6681 14568 6819 14592
rect 1548 14508 1752 14532
rect 2628 14508 2952 14532
rect 5448 14532 5472 14562
rect 5448 14508 5892 14532
rect 981 14445 1179 14469
rect 1548 14472 1572 14508
rect 1341 14460 1692 14472
rect 1341 14448 1701 14460
rect 1659 14421 1701 14448
rect 2001 14448 2439 14472
rect 2628 14478 2652 14508
rect 2928 14478 2952 14508
rect 3081 14448 3459 14472
rect 4641 14448 5139 14472
rect 5181 14448 5559 14472
rect 5601 14445 5739 14469
rect 5868 14472 5892 14508
rect 5868 14448 5919 14472
rect 6261 14448 6579 14472
rect 6741 14445 6879 14469
rect 7008 14472 7032 14619
rect 7008 14448 7239 14472
rect 8028 14478 8052 14628
rect 11121 14628 11472 14652
rect 8301 14568 8499 14592
rect 9141 14568 9372 14592
rect 8628 14532 8652 14562
rect 8628 14508 9012 14532
rect 8181 14445 8259 14469
rect 8421 14445 8559 14469
rect 8988 14472 9012 14508
rect 8988 14448 9072 14472
rect 441 14388 519 14412
rect 4041 14388 4359 14412
rect 4401 14388 5799 14412
rect 7161 14388 7839 14412
rect 8559 14412 8601 14436
rect 9048 14421 9072 14448
rect 8559 14388 8919 14412
rect 9048 14388 9099 14421
rect 9060 14379 9099 14388
rect 9348 14412 9372 14568
rect 9501 14568 9699 14592
rect 9981 14568 10572 14592
rect 10548 14532 10572 14568
rect 10701 14568 10839 14592
rect 11001 14568 11139 14592
rect 10548 14508 10632 14532
rect 10608 14478 10632 14508
rect 9621 14445 9879 14469
rect 10641 14448 11199 14472
rect 9348 14388 9519 14412
rect 11268 14412 11292 14559
rect 11448 14478 11472 14628
rect 12141 14628 12579 14652
rect 11541 14568 11652 14592
rect 11628 14481 11652 14568
rect 11928 14478 11952 14619
rect 12021 14568 12192 14592
rect 12168 14532 12192 14568
rect 12261 14571 12399 14595
rect 12168 14508 12492 14532
rect 12081 14448 12219 14472
rect 12468 14478 12492 14508
rect 12528 14421 12552 14628
rect 13461 14628 13539 14652
rect 14241 14628 14559 14652
rect 15561 14628 15699 14652
rect 15741 14628 15819 14652
rect 16761 14628 16839 14652
rect 17301 14628 17412 14652
rect 12588 14481 12612 14556
rect 13308 14532 13332 14562
rect 13821 14568 14139 14592
rect 14208 14568 14259 14592
rect 12681 14508 13332 14532
rect 12981 14448 13239 14472
rect 13281 14448 13359 14472
rect 11268 14388 11379 14412
rect 12381 14388 12519 14412
rect 13488 14412 13512 14559
rect 13668 14532 13692 14562
rect 13608 14520 13692 14532
rect 13599 14508 13692 14520
rect 13599 14481 13641 14508
rect 14208 14532 14232 14568
rect 14841 14568 14979 14592
rect 15048 14568 15099 14592
rect 15048 14532 15072 14568
rect 15441 14568 15579 14592
rect 16359 14592 16401 14619
rect 16359 14580 16539 14592
rect 16368 14568 16539 14580
rect 14061 14508 14232 14532
rect 14988 14508 15072 14532
rect 14361 14448 14679 14472
rect 14988 14421 15012 14508
rect 15228 14481 15252 14559
rect 15381 14445 15519 14469
rect 15768 14472 15792 14559
rect 16668 14481 16692 14559
rect 16779 14532 16821 14559
rect 16779 14520 16932 14532
rect 16788 14508 16932 14520
rect 15708 14460 15792 14472
rect 15699 14448 15792 14460
rect 15699 14421 15741 14448
rect 15861 14445 15939 14469
rect 16281 14445 16479 14469
rect 16908 14478 16932 14508
rect 17088 14481 17112 14559
rect 17328 14532 17352 14562
rect 17268 14520 17352 14532
rect 17259 14508 17352 14520
rect 17388 14532 17412 14628
rect 17481 14568 18279 14592
rect 17388 14508 17532 14532
rect 17259 14481 17301 14508
rect 17508 14478 17532 14508
rect 13488 14388 13659 14412
rect 801 14328 999 14352
rect 2181 14328 2619 14352
rect 3801 14328 4179 14352
rect 4941 14328 5619 14352
rect 6021 14328 6339 14352
rect 9681 14328 10239 14352
rect 10401 14328 10839 14352
rect 11001 14328 11559 14352
rect 12261 14328 12999 14352
rect 13401 14328 13719 14352
rect 14061 14328 14619 14352
rect 15441 14328 16059 14352
rect 16941 14328 17379 14352
rect 3321 14268 4659 14292
rect 4701 14268 4779 14292
rect 6441 14268 7599 14292
rect 9921 14268 10059 14292
rect 11901 14268 13119 14292
rect 13161 14268 13239 14292
rect 13560 14292 13599 14301
rect 13548 14259 13599 14292
rect 14001 14268 14532 14292
rect 321 14208 579 14232
rect 621 14208 639 14232
rect 681 14208 1599 14232
rect 1641 14208 2199 14232
rect 4101 14208 5979 14232
rect 6021 14208 6759 14232
rect 6828 14208 7179 14232
rect 1041 14148 1719 14172
rect 2301 14148 3159 14172
rect 3768 14148 4059 14172
rect 2361 14088 3579 14112
rect 3768 14112 3792 14148
rect 4221 14148 5379 14172
rect 6828 14172 6852 14208
rect 8721 14208 10719 14232
rect 11748 14208 12699 14232
rect 6381 14148 6852 14172
rect 7341 14148 9039 14172
rect 9081 14148 9999 14172
rect 11748 14172 11772 14208
rect 13548 14232 13572 14259
rect 12861 14208 13572 14232
rect 14508 14232 14532 14268
rect 14721 14268 18159 14292
rect 14508 14208 15519 14232
rect 15681 14208 15759 14232
rect 15801 14208 16119 14232
rect 11361 14148 11772 14172
rect 11841 14148 12159 14172
rect 12621 14148 13476 14172
rect 13581 14148 13899 14172
rect 14121 14148 15039 14172
rect 3621 14088 3792 14112
rect 3921 14088 5439 14112
rect 5481 14088 6279 14112
rect 6528 14088 7059 14112
rect 1461 14028 1839 14052
rect 4521 14028 4839 14052
rect 4881 14028 5019 14052
rect 6528 14052 6552 14088
rect 7281 14088 8739 14112
rect 9141 14088 9819 14112
rect 10881 14088 11079 14112
rect 12021 14088 12639 14112
rect 13101 14088 14136 14112
rect 14241 14088 15639 14112
rect 15801 14088 16419 14112
rect 16461 14088 16659 14112
rect 5841 14028 6552 14052
rect 6621 14028 8832 14052
rect 81 13968 2319 13992
rect 3681 13968 3879 13992
rect 5241 13968 6999 13992
rect 7221 13968 8079 13992
rect 8808 13992 8832 14028
rect 10701 14028 10959 14052
rect 11001 14028 11079 14052
rect 11781 14028 12999 14052
rect 13881 14028 14439 14052
rect 14661 14028 16959 14052
rect 8808 13968 9219 13992
rect 9861 13968 11979 13992
rect 12321 13968 12579 13992
rect 13521 13968 13839 13992
rect 16101 13968 16899 13992
rect 17721 13968 18279 13992
rect 2661 13908 3459 13932
rect 4221 13908 4779 13932
rect 4821 13908 8199 13932
rect 8661 13908 8799 13932
rect 9801 13908 10656 13932
rect 10761 13908 12552 13932
rect 1521 13848 2919 13872
rect 5181 13848 5676 13872
rect 5781 13848 6552 13872
rect 261 13788 699 13812
rect 3141 13788 3219 13812
rect 6528 13812 6552 13848
rect 6921 13848 7299 13872
rect 11481 13848 12459 13872
rect 12528 13872 12552 13908
rect 13041 13908 13959 13932
rect 15261 13908 15459 13932
rect 15681 13908 16599 13932
rect 17181 13908 17499 13932
rect 12528 13848 12819 13872
rect 13641 13848 13899 13872
rect 15321 13848 15579 13872
rect 16581 13848 16719 13872
rect 17001 13848 17739 13872
rect 6528 13788 7119 13812
rect 7641 13788 7839 13812
rect 8001 13788 8799 13812
rect 9321 13788 10479 13812
rect 11661 13788 13356 13812
rect 13461 13788 13719 13812
rect 14241 13788 14439 13812
rect 14961 13788 16059 13812
rect 16281 13788 16659 13812
rect 2241 13728 3252 13752
rect 141 13671 219 13695
rect 381 13671 456 13695
rect 921 13668 1179 13692
rect 1341 13668 1539 13692
rect 1701 13668 2019 13692
rect 528 13572 552 13659
rect 1548 13632 1572 13662
rect 2148 13632 2172 13662
rect 2361 13668 2439 13692
rect 3141 13692 3180 13701
rect 3228 13692 3252 13728
rect 3441 13728 3639 13752
rect 6501 13728 6639 13752
rect 8901 13728 9039 13752
rect 13188 13728 13539 13752
rect 3141 13659 3192 13692
rect 3228 13668 3672 13692
rect 1548 13608 2172 13632
rect 3168 13632 3192 13659
rect 3168 13608 3612 13632
rect 528 13548 639 13572
rect 981 13548 1119 13572
rect 1641 13548 2079 13572
rect 1821 13488 1899 13512
rect 2148 13512 2172 13608
rect 2421 13548 3099 13572
rect 3588 13578 3612 13608
rect 3321 13545 3516 13569
rect 3648 13572 3672 13668
rect 3801 13671 3939 13695
rect 4701 13668 5019 13692
rect 5088 13668 5139 13692
rect 4548 13632 4572 13662
rect 5088 13632 5112 13668
rect 4428 13620 4572 13632
rect 4419 13608 4572 13620
rect 4608 13608 5112 13632
rect 4419 13581 4461 13608
rect 3648 13548 3699 13572
rect 3981 13548 4119 13572
rect 4608 13578 4632 13608
rect 5361 13548 5439 13572
rect 2148 13488 2679 13512
rect 5508 13512 5532 13662
rect 5661 13668 5859 13692
rect 5901 13671 6159 13695
rect 7101 13671 8439 13695
rect 8481 13668 8679 13692
rect 5721 13548 6339 13572
rect 6408 13572 6432 13662
rect 9168 13668 9279 13692
rect 9168 13632 9192 13668
rect 9501 13668 9699 13692
rect 9981 13668 10839 13692
rect 11241 13671 11439 13695
rect 12081 13668 12339 13692
rect 12480 13692 12519 13701
rect 12468 13659 12519 13692
rect 12801 13671 12879 13695
rect 7401 13608 8112 13632
rect 6408 13548 6519 13572
rect 8088 13572 8112 13608
rect 8988 13608 9192 13632
rect 8088 13548 8499 13572
rect 8541 13548 8739 13572
rect 8988 13572 9012 13608
rect 8901 13548 9012 13572
rect 9081 13545 9219 13569
rect 11361 13548 11499 13572
rect 12468 13521 12492 13659
rect 13188 13632 13212 13728
rect 13941 13728 14139 13752
rect 14721 13728 14859 13752
rect 15339 13728 15939 13752
rect 15339 13704 15381 13728
rect 18441 13752 18480 13761
rect 18441 13719 18492 13752
rect 13401 13668 13692 13692
rect 13128 13608 13212 13632
rect 13668 13632 13692 13668
rect 13761 13668 15072 13692
rect 15048 13641 15072 13668
rect 15201 13671 15339 13695
rect 16080 13692 16119 13701
rect 13668 13620 13752 13632
rect 13668 13608 13761 13620
rect 15048 13608 15099 13641
rect 13128 13578 13152 13608
rect 13719 13581 13761 13608
rect 15060 13599 15099 13608
rect 12621 13545 12699 13569
rect 15468 13581 15492 13662
rect 15828 13581 15852 13662
rect 16068 13659 16119 13692
rect 16068 13581 16092 13659
rect 14121 13545 14859 13569
rect 15468 13548 15519 13581
rect 15480 13539 15519 13548
rect 15801 13548 15852 13581
rect 15801 13539 15840 13548
rect 16308 13572 16332 13719
rect 16401 13668 16479 13692
rect 16881 13668 16932 13692
rect 16908 13581 16932 13668
rect 16308 13548 16419 13572
rect 17148 13521 17172 13719
rect 17841 13668 18192 13692
rect 17679 13632 17721 13659
rect 17679 13620 17772 13632
rect 17688 13608 17772 13620
rect 17748 13578 17772 13608
rect 18168 13578 18192 13668
rect 18261 13671 18399 13695
rect 18468 13632 18492 13719
rect 18348 13620 18492 13632
rect 18339 13608 18492 13620
rect 18339 13581 18381 13608
rect 5241 13488 5532 13512
rect 5721 13488 6579 13512
rect 7101 13488 8439 13512
rect 9441 13488 9519 13512
rect 12021 13488 12396 13512
rect 13821 13488 13959 13512
rect 15021 13488 15159 13512
rect 16221 13488 16599 13512
rect 17541 13488 17619 13512
rect 561 13428 879 13452
rect 2481 13428 2559 13452
rect 3201 13428 3699 13452
rect 4461 13428 5079 13452
rect 5301 13428 5559 13452
rect 5601 13428 5739 13452
rect 6261 13428 6516 13452
rect 6621 13428 6879 13452
rect 8781 13428 9939 13452
rect 9981 13428 10659 13452
rect 10881 13428 11559 13452
rect 11721 13428 12039 13452
rect 12681 13428 12876 13452
rect 12981 13428 13719 13452
rect 13881 13428 14019 13452
rect 14361 13428 15279 13452
rect 15321 13428 15759 13452
rect 16161 13428 16419 13452
rect 17721 13428 18279 13452
rect 321 13368 1239 13392
rect 1281 13368 1599 13392
rect 1761 13368 2319 13392
rect 3501 13368 4359 13392
rect 6501 13368 7359 13392
rect 8661 13368 11799 13392
rect 13521 13368 14259 13392
rect 14481 13368 15999 13392
rect 16041 13368 16539 13392
rect 16581 13368 16719 13392
rect 18021 13368 18279 13392
rect 3561 13308 3936 13332
rect 4041 13308 4239 13332
rect 7461 13308 7959 13332
rect 8121 13308 8379 13332
rect 8841 13308 9099 13332
rect 10761 13308 11139 13332
rect 12081 13308 13119 13332
rect 13581 13308 13779 13332
rect 13941 13308 14739 13332
rect 15321 13308 15399 13332
rect 15681 13308 16179 13332
rect 17181 13308 17439 13332
rect 2961 13248 3336 13272
rect 3441 13248 4959 13272
rect 5601 13248 5919 13272
rect 6921 13248 7299 13272
rect 7521 13248 7599 13272
rect 8241 13248 9159 13272
rect 9201 13248 9639 13272
rect 9921 13248 11919 13272
rect 12201 13248 12699 13272
rect 13461 13248 13839 13272
rect 14001 13248 14199 13272
rect 16821 13248 16899 13272
rect 17901 13248 18039 13272
rect 18081 13248 18339 13272
rect 1881 13188 1959 13212
rect 2001 13188 2619 13212
rect 2901 13188 2979 13212
rect 3021 13188 5019 13212
rect 5661 13188 6399 13212
rect 7281 13188 7899 13212
rect 8061 13188 8139 13212
rect 8181 13188 8319 13212
rect 10281 13188 10779 13212
rect 11181 13188 11859 13212
rect 13401 13188 13899 13212
rect 14241 13188 14319 13212
rect 14781 13188 15399 13212
rect 15441 13188 15579 13212
rect 17181 13188 17319 13212
rect 741 13128 1119 13152
rect 2601 13128 4479 13152
rect 4761 13128 5439 13152
rect 7401 13128 8199 13152
rect 8421 13128 8739 13152
rect 9921 13128 9999 13152
rect 10401 13128 10599 13152
rect 12921 13128 13536 13152
rect 13641 13128 14439 13152
rect 15201 13128 15339 13152
rect 15861 13128 16899 13152
rect 17841 13128 18219 13152
rect 921 13068 1359 13092
rect 2241 13068 2379 13092
rect 3321 13068 3459 13092
rect 3621 13068 3999 13092
rect 6021 13092 6060 13101
rect 6021 13059 6072 13092
rect 7341 13068 8079 13092
rect 11901 13068 12219 13092
rect 13221 13068 13659 13092
rect 13821 13068 14079 13092
rect 15021 13068 15099 13092
rect 17001 13068 17172 13092
rect 201 13011 279 13035
rect 501 13008 672 13032
rect 381 12888 519 12912
rect 648 12918 672 13008
rect 768 12972 792 13059
rect 861 13011 936 13035
rect 999 12972 1041 12999
rect 1428 13008 1599 13032
rect 768 12948 972 12972
rect 999 12960 1152 12972
rect 1008 12948 1152 12960
rect 948 12912 972 12948
rect 948 12888 1059 12912
rect 1128 12912 1152 12948
rect 1428 12921 1452 13008
rect 3561 13008 3612 13032
rect 2028 12921 2052 13002
rect 3588 12921 3612 13008
rect 5508 13008 5619 13032
rect 3861 12948 4176 12972
rect 1128 12888 1299 12912
rect 2028 12888 2079 12921
rect 2040 12879 2079 12888
rect 2481 12885 3039 12909
rect 3201 12885 3279 12909
rect 3588 12888 3639 12921
rect 3600 12879 3639 12888
rect 4239 12912 4281 12939
rect 4239 12900 4899 12912
rect 4248 12888 4899 12900
rect 5328 12912 5352 13002
rect 5508 12918 5532 13008
rect 6048 13032 6072 13059
rect 6048 13008 7059 13032
rect 8088 13008 8259 13032
rect 7248 12921 7272 12999
rect 8088 12921 8112 13008
rect 8421 13032 8460 13041
rect 8421 12999 8472 13032
rect 8721 13008 8799 13032
rect 8928 13008 10119 13032
rect 8448 12921 8472 12999
rect 8928 12921 8952 13008
rect 10281 13008 10479 13032
rect 10680 13032 10719 13041
rect 10668 12999 10719 13032
rect 5181 12888 5352 12912
rect 10668 12918 10692 12999
rect 10908 12921 10932 13059
rect 11088 12921 11112 13002
rect 10908 12888 10959 12921
rect 10920 12879 10959 12888
rect 11088 12888 11139 12921
rect 11100 12879 11139 12888
rect 1221 12828 1659 12852
rect 1701 12828 1839 12852
rect 2361 12828 2799 12852
rect 2841 12828 3012 12852
rect 1401 12768 1539 12792
rect 2988 12792 3012 12828
rect 3981 12828 4659 12852
rect 5961 12828 6219 12852
rect 8001 12828 8379 12852
rect 11208 12852 11232 13008
rect 14088 13008 14379 13032
rect 11508 12921 11532 12999
rect 12168 12972 12192 13002
rect 11928 12948 12192 12972
rect 11928 12912 11952 12948
rect 11661 12888 11952 12912
rect 12021 12885 12099 12909
rect 12288 12912 12312 13002
rect 12288 12888 12399 12912
rect 12621 12888 13656 12912
rect 13761 12888 13839 12912
rect 13908 12861 13932 13002
rect 14028 12861 14052 13002
rect 14088 12918 14112 13008
rect 14541 13011 14679 13035
rect 14721 13008 14919 13032
rect 15228 12972 15252 13059
rect 15048 12960 15252 12972
rect 15039 12948 15252 12960
rect 15039 12921 15081 12948
rect 14481 12888 14799 12912
rect 15288 12861 15312 13002
rect 15501 13008 15639 13032
rect 16041 13008 16239 13032
rect 15861 12888 15939 12912
rect 10761 12828 11232 12852
rect 15408 12828 15759 12852
rect 2988 12768 3459 12792
rect 5061 12768 5199 12792
rect 7521 12768 8199 12792
rect 9081 12768 9819 12792
rect 10881 12768 11016 12792
rect 11121 12768 11739 12792
rect 11961 12768 12279 12792
rect 14601 12768 14679 12792
rect 14721 12768 14859 12792
rect 15408 12792 15432 12828
rect 16368 12855 16392 13002
rect 16488 12912 16512 12999
rect 17028 12921 17052 12999
rect 17148 12921 17172 13068
rect 17241 13068 17739 13092
rect 17361 13008 17619 13032
rect 17688 12921 17712 13068
rect 17928 12921 17952 12999
rect 16461 12888 16512 12912
rect 16641 12885 16719 12909
rect 16368 12828 16419 12855
rect 16380 12819 16419 12828
rect 16881 12828 16899 12852
rect 16941 12828 17259 12852
rect 17661 12828 17739 12852
rect 15201 12768 15432 12792
rect 17481 12768 17559 12792
rect 1821 12708 2139 12732
rect 2301 12708 3219 12732
rect 3741 12708 4419 12732
rect 5121 12708 5199 12732
rect 5241 12708 5679 12732
rect 6321 12708 6579 12732
rect 9621 12708 10359 12732
rect 12801 12708 13419 12732
rect 15141 12708 15459 12732
rect 15981 12708 16659 12732
rect 16821 12708 17019 12732
rect 17901 12708 18099 12732
rect 3441 12648 4776 12672
rect 4881 12648 5979 12672
rect 7161 12648 7959 12672
rect 8121 12648 8352 12672
rect 2001 12588 2319 12612
rect 3621 12588 3879 12612
rect 4821 12588 5919 12612
rect 8328 12612 8352 12648
rect 13581 12648 14379 12672
rect 14541 12648 14979 12672
rect 15561 12648 16959 12672
rect 8328 12588 8859 12612
rect 9801 12588 10719 12612
rect 11001 12588 11319 12612
rect 12441 12588 16119 12612
rect 2421 12528 2739 12552
rect 3381 12528 3999 12552
rect 4761 12528 7599 12552
rect 8148 12528 8619 12552
rect 8148 12501 8172 12528
rect 10941 12528 12579 12552
rect 14421 12528 15159 12552
rect 16581 12528 16719 12552
rect 4641 12468 6792 12492
rect 6768 12441 6792 12468
rect 7761 12468 8139 12492
rect 8721 12468 9039 12492
rect 9348 12468 11139 12492
rect 2121 12408 2679 12432
rect 2721 12408 3279 12432
rect 3321 12408 3639 12432
rect 6801 12408 7299 12432
rect 9348 12432 9372 12468
rect 11421 12468 12039 12492
rect 12741 12468 14199 12492
rect 14421 12468 14799 12492
rect 17088 12468 17679 12492
rect 7341 12408 9372 12432
rect 10821 12408 10959 12432
rect 13941 12408 15219 12432
rect 16221 12408 16299 12432
rect 17088 12432 17112 12468
rect 16641 12408 17112 12432
rect 5001 12348 6159 12372
rect 6201 12348 6339 12372
rect 6561 12348 6759 12372
rect 6801 12348 7092 12372
rect 3261 12288 3759 12312
rect 3801 12288 4119 12312
rect 4341 12288 5139 12312
rect 7068 12312 7092 12348
rect 7941 12348 9759 12372
rect 10581 12348 11019 12372
rect 11061 12348 11439 12372
rect 11481 12348 12219 12372
rect 12561 12348 12699 12372
rect 12981 12348 13359 12372
rect 13401 12348 13659 12372
rect 13941 12348 14019 12372
rect 14841 12348 15039 12372
rect 15681 12348 16059 12372
rect 17301 12348 17379 12372
rect 17421 12348 17859 12372
rect 17901 12348 18099 12372
rect 7068 12288 7419 12312
rect 8121 12288 8499 12312
rect 9981 12288 10479 12312
rect 13101 12288 13959 12312
rect 14661 12288 15399 12312
rect 15441 12288 15519 12312
rect 16461 12288 17379 12312
rect 381 12228 939 12252
rect 981 12228 1179 12252
rect 1521 12228 2259 12252
rect 5421 12228 6879 12252
rect 648 12168 759 12192
rect 501 12111 579 12135
rect 648 12021 672 12168
rect 4041 12168 4299 12192
rect 4848 12168 5199 12192
rect 741 12108 999 12132
rect 1041 12108 1479 12132
rect 1521 12111 1599 12135
rect 1761 12108 2019 12132
rect 3621 12111 3819 12135
rect 4281 12108 4419 12132
rect 2361 12048 2859 12072
rect 201 11988 279 12012
rect 1548 12000 1659 12012
rect 1539 11988 1659 12000
rect 1539 11961 1581 11988
rect 3921 11988 4479 12012
rect 4848 12012 4872 12168
rect 5661 12168 5739 12192
rect 4941 12108 5439 12132
rect 5508 12108 5739 12132
rect 5508 12072 5532 12108
rect 5808 12072 5832 12228
rect 7041 12228 8019 12252
rect 8601 12228 9879 12252
rect 9921 12228 9999 12252
rect 11301 12228 11739 12252
rect 11781 12228 11919 12252
rect 12081 12228 12339 12252
rect 13161 12228 13239 12252
rect 14961 12228 15219 12252
rect 16881 12228 17259 12252
rect 17388 12252 17412 12276
rect 17388 12228 18279 12252
rect 6441 12168 6639 12192
rect 7461 12168 7839 12192
rect 7881 12168 7959 12192
rect 8208 12168 8439 12192
rect 5961 12111 6159 12135
rect 6501 12108 6639 12132
rect 6681 12108 6999 12132
rect 7899 12072 7941 12099
rect 5388 12048 5532 12072
rect 5688 12048 5832 12072
rect 7608 12060 7941 12072
rect 8208 12072 8232 12168
rect 12201 12168 12621 12192
rect 8301 12108 8559 12132
rect 8601 12108 8799 12132
rect 7608 12048 7932 12060
rect 8208 12048 8532 12072
rect 5388 12018 5412 12048
rect 5688 12018 5712 12048
rect 4701 11988 4872 12012
rect 6321 11988 7059 12012
rect 7608 12012 7632 12048
rect 8508 12018 8532 12048
rect 9528 12021 9552 12108
rect 9708 12072 9732 12108
rect 9708 12048 9879 12072
rect 7101 11988 7632 12012
rect 7761 11985 8079 12009
rect 8241 12000 8352 12012
rect 8241 11988 8361 12000
rect 8319 11961 8361 11988
rect 8661 11988 8739 12012
rect 8781 11988 8919 12012
rect 9501 11988 9552 12021
rect 10068 12018 10092 12159
rect 10128 12021 10152 12102
rect 10581 12108 10659 12132
rect 12579 12144 12621 12168
rect 12681 12168 12852 12192
rect 10881 12108 11079 12132
rect 10848 12021 10872 12108
rect 11541 12111 11619 12135
rect 12621 12111 12759 12135
rect 9501 11979 9540 11988
rect 10128 11988 10179 12021
rect 10140 11979 10179 11988
rect 10341 11979 10479 12003
rect 10848 11988 10899 12021
rect 10860 11979 10899 11988
rect 11241 11988 11499 12012
rect 441 11928 759 11952
rect 2181 11928 3039 11952
rect 5148 11928 5319 11952
rect 1461 11868 2019 11892
rect 3801 11868 4179 11892
rect 4401 11868 4719 11892
rect 5148 11892 5172 11928
rect 11868 11952 11892 12099
rect 12228 12012 12252 12099
rect 12408 12021 12432 12099
rect 12141 11988 12252 12012
rect 12828 12012 12852 12168
rect 15381 12168 15459 12192
rect 16161 12168 16599 12192
rect 17868 12168 18252 12192
rect 13821 12108 14079 12132
rect 14301 12108 14499 12132
rect 14568 12108 14679 12132
rect 13188 12021 13212 12099
rect 14568 12072 14592 12108
rect 15708 12108 15759 12132
rect 14508 12048 14592 12072
rect 12681 11988 12852 12012
rect 12981 11985 13059 12009
rect 13761 11988 13839 12012
rect 14181 11985 14259 12009
rect 14508 11961 14532 12048
rect 15708 12021 15732 12108
rect 16188 12120 16839 12132
rect 16179 12108 16839 12120
rect 16179 12078 16221 12108
rect 17421 12108 17472 12132
rect 17208 12021 17232 12099
rect 17448 12021 17472 12108
rect 17868 12132 17892 12168
rect 18228 12141 18252 12168
rect 17781 12108 17892 12132
rect 17961 12132 18000 12141
rect 17961 12099 18012 12132
rect 15321 11985 15399 12009
rect 16821 11988 17079 12012
rect 17748 12012 17772 12099
rect 17661 11988 17772 12012
rect 17988 12012 18012 12099
rect 18039 12072 18081 12099
rect 18039 12060 18192 12072
rect 18048 12048 18192 12060
rect 18168 12018 18192 12048
rect 17988 12000 18132 12012
rect 17988 11988 18141 12000
rect 18099 11961 18141 11988
rect 18408 12012 18432 12159
rect 18408 11988 18492 12012
rect 11601 11928 11892 11952
rect 12021 11928 12279 11952
rect 13941 11928 14019 11952
rect 4881 11868 5172 11892
rect 5421 11868 5499 11892
rect 5961 11868 6279 11892
rect 6441 11868 8619 11892
rect 9921 11868 10239 11892
rect 10281 11868 10899 11892
rect 10941 11868 13659 11892
rect 13821 11868 14559 11892
rect 15381 11868 15819 11892
rect 17361 11868 17619 11892
rect 17841 11868 18399 11892
rect 81 11808 1239 11832
rect 1521 11808 2079 11832
rect 2481 11808 2619 11832
rect 3021 11808 3579 11832
rect 3741 11808 4239 11832
rect 4821 11808 5319 11832
rect 5601 11808 6099 11832
rect 10308 11820 10479 11832
rect 10299 11808 10479 11820
rect 10299 11781 10341 11808
rect 11541 11808 13239 11832
rect 14001 11808 14379 11832
rect 14661 11808 15279 11832
rect 17541 11808 17919 11832
rect 18468 11781 18492 11988
rect 381 11748 999 11772
rect 2061 11748 2559 11772
rect 2688 11748 5259 11772
rect 501 11688 819 11712
rect 861 11688 2259 11712
rect 2688 11712 2712 11748
rect 6741 11748 7992 11772
rect 7968 11721 7992 11748
rect 9921 11748 10179 11772
rect 10581 11748 11679 11772
rect 11841 11748 12639 11772
rect 14781 11748 15039 11772
rect 15681 11748 15759 11772
rect 18201 11748 18279 11772
rect 18441 11748 18492 11781
rect 18441 11739 18480 11748
rect 2301 11688 2712 11712
rect 3141 11688 3339 11712
rect 3561 11688 3819 11712
rect 4821 11688 4899 11712
rect 4941 11688 5079 11712
rect 7641 11688 7839 11712
rect 8001 11688 8799 11712
rect 9381 11688 9579 11712
rect 10281 11688 10359 11712
rect 10881 11688 11019 11712
rect 12561 11688 12639 11712
rect 14748 11712 14772 11739
rect 13341 11688 14772 11712
rect 15321 11688 15819 11712
rect 1161 11628 1539 11652
rect 1581 11628 2499 11652
rect 4341 11628 4599 11652
rect 5301 11628 5679 11652
rect 6561 11628 6819 11652
rect 8301 11628 8739 11652
rect 9681 11628 10419 11652
rect 13881 11628 14679 11652
rect 15261 11628 15879 11652
rect 16941 11628 17379 11652
rect 18081 11628 18219 11652
rect 2721 11568 3459 11592
rect 3861 11568 4539 11592
rect 4941 11568 5079 11592
rect 5241 11568 5559 11592
rect 5781 11568 6039 11592
rect 7701 11568 7839 11592
rect 8121 11568 8379 11592
rect 8421 11568 9099 11592
rect 9261 11568 9399 11592
rect 9621 11568 10632 11592
rect 201 11508 759 11532
rect 801 11508 1239 11532
rect 1821 11508 1899 11532
rect 1941 11508 2439 11532
rect 6681 11508 6759 11532
rect 7461 11508 7539 11532
rect 8181 11508 8379 11532
rect 921 11448 1059 11472
rect 1761 11448 1812 11472
rect 201 11325 279 11349
rect 588 11352 612 11439
rect 1788 11361 1812 11448
rect 2160 11472 2199 11481
rect 2148 11439 2199 11472
rect 2568 11448 2739 11472
rect 588 11328 759 11352
rect 1221 11328 1539 11352
rect 1581 11325 1659 11349
rect 1788 11328 1839 11361
rect 1800 11319 1839 11328
rect 1968 11352 1992 11439
rect 2148 11358 2172 11439
rect 2568 11361 2592 11448
rect 2901 11448 3279 11472
rect 3441 11448 3912 11472
rect 1968 11328 2019 11352
rect 2301 11325 2379 11349
rect 2721 11325 2799 11349
rect 2841 11328 3159 11352
rect 3888 11358 3912 11448
rect 3948 11361 3972 11442
rect 4521 11448 4659 11472
rect 4728 11448 4899 11472
rect 4728 11412 4752 11448
rect 5061 11472 5100 11481
rect 5061 11439 5112 11472
rect 4101 11388 4752 11412
rect 3681 11325 3759 11349
rect 3948 11328 3999 11361
rect 3960 11319 3999 11328
rect 4341 11325 4539 11349
rect 4761 11325 5019 11349
rect 2139 11292 2181 11316
rect 1161 11268 2181 11292
rect 3381 11268 3519 11292
rect 5088 11295 5112 11439
rect 5148 11412 5172 11499
rect 8421 11508 8679 11532
rect 9021 11508 9159 11532
rect 9981 11508 10479 11532
rect 5319 11412 5361 11439
rect 5148 11388 5232 11412
rect 5319 11400 5412 11412
rect 5328 11388 5412 11400
rect 5208 11352 5232 11388
rect 5208 11328 5319 11352
rect 5388 11352 5412 11388
rect 5388 11328 5499 11352
rect 5688 11352 5712 11439
rect 5841 11451 5919 11475
rect 5961 11448 6579 11472
rect 7101 11448 7332 11472
rect 6699 11412 6741 11439
rect 6648 11400 6741 11412
rect 6648 11388 6732 11400
rect 6648 11358 6672 11388
rect 7005 11361 7029 11439
rect 5688 11328 5979 11352
rect 6021 11325 6576 11349
rect 6861 11328 6936 11352
rect 5148 11292 5172 11316
rect 7308 11301 7332 11448
rect 7821 11448 7899 11472
rect 7368 11352 7392 11439
rect 8088 11361 8112 11439
rect 7368 11328 7479 11352
rect 8421 11325 8499 11349
rect 8568 11301 8592 11442
rect 8901 11448 9279 11472
rect 9639 11412 9681 11439
rect 8748 11400 9681 11412
rect 10128 11448 10299 11472
rect 8748 11388 9672 11400
rect 8748 11301 8772 11388
rect 10128 11361 10152 11448
rect 10608 11472 10632 11568
rect 11661 11568 12219 11592
rect 15081 11568 15699 11592
rect 16281 11568 16419 11592
rect 16641 11568 16779 11592
rect 17361 11568 17499 11592
rect 17721 11568 17799 11592
rect 11001 11508 11199 11532
rect 15861 11508 16479 11532
rect 16848 11508 16959 11532
rect 10581 11448 10632 11472
rect 11061 11448 11256 11472
rect 11688 11448 11799 11472
rect 8841 11325 8919 11349
rect 9081 11328 9519 11352
rect 9981 11328 10056 11352
rect 10281 11319 10359 11343
rect 11328 11352 11352 11439
rect 10521 11328 11352 11352
rect 11448 11352 11472 11439
rect 11568 11361 11592 11439
rect 11688 11361 11712 11448
rect 12339 11481 12381 11499
rect 12081 11457 12459 11481
rect 12348 11448 12372 11457
rect 13281 11451 13479 11475
rect 12759 11412 12801 11439
rect 11421 11328 11472 11352
rect 11979 11352 12021 11379
rect 11901 11340 12021 11352
rect 12588 11400 12801 11412
rect 12588 11388 12792 11400
rect 11901 11328 12012 11340
rect 12588 11301 12612 11388
rect 13668 11352 13692 11439
rect 15288 11412 15312 11442
rect 16161 11448 16332 11472
rect 15108 11388 15312 11412
rect 16308 11412 16332 11448
rect 16401 11451 16539 11475
rect 16308 11400 16752 11412
rect 16308 11388 16761 11400
rect 12681 11319 12819 11343
rect 13668 11328 13719 11352
rect 14181 11325 14679 11349
rect 15108 11352 15132 11388
rect 16719 11361 16761 11388
rect 14841 11328 15132 11352
rect 15201 11328 15759 11352
rect 16848 11358 16872 11508
rect 17181 11508 17559 11532
rect 18141 11508 18279 11532
rect 17241 11448 17352 11472
rect 17328 11301 17352 11448
rect 17388 11448 17679 11472
rect 17388 11358 17412 11448
rect 17901 11448 17979 11472
rect 18168 11361 18192 11439
rect 5148 11268 5739 11292
rect 6141 11268 6279 11292
rect 6321 11268 6459 11292
rect 6681 11268 7119 11292
rect 7308 11268 7359 11301
rect 7320 11259 7359 11268
rect 7701 11268 7959 11292
rect 8721 11268 8772 11301
rect 8721 11259 8760 11268
rect 9321 11268 9639 11292
rect 10461 11268 10959 11292
rect 12588 11298 12660 11301
rect 12588 11268 12639 11298
rect 12600 11259 12639 11268
rect 13221 11268 13359 11292
rect 14841 11268 15939 11292
rect 561 11208 939 11232
rect 981 11208 2499 11232
rect 2541 11208 4059 11232
rect 4221 11208 4599 11232
rect 5061 11208 5259 11232
rect 5421 11208 5499 11232
rect 6921 11208 6999 11232
rect 7221 11208 7719 11232
rect 9561 11208 9939 11232
rect 10761 11208 11259 11232
rect 13521 11208 13959 11232
rect 15081 11208 15399 11232
rect 15861 11208 16059 11232
rect 16281 11208 16539 11232
rect 16581 11208 16959 11232
rect 17601 11208 17739 11232
rect 1821 11148 2019 11172
rect 2061 11148 2679 11172
rect 3141 11148 3459 11172
rect 5361 11148 6276 11172
rect 6381 11148 6939 11172
rect 12321 11148 12699 11172
rect 13281 11148 13359 11172
rect 13701 11148 13899 11172
rect 15501 11148 16419 11172
rect 4881 11088 5379 11112
rect 5541 11088 5859 11112
rect 5901 11088 6072 11112
rect 3021 11028 4599 11052
rect 4641 11028 5439 11052
rect 6048 11052 6072 11088
rect 6441 11088 6999 11112
rect 7641 11088 8379 11112
rect 9021 11088 9579 11112
rect 11121 11088 12039 11112
rect 14001 11088 15219 11112
rect 6048 11028 7239 11052
rect 7281 11028 8679 11052
rect 9141 11028 10059 11052
rect 11721 11028 12159 11052
rect 15141 11028 15459 11052
rect 18081 11028 18339 11052
rect 2121 10968 2619 10992
rect 5001 10968 5139 10992
rect 5661 10968 6432 10992
rect 3801 10908 4932 10932
rect 81 10848 999 10872
rect 1041 10848 1299 10872
rect 4908 10872 4932 10908
rect 5001 10908 5919 10932
rect 6408 10932 6432 10968
rect 6501 10968 7299 10992
rect 8781 10968 9819 10992
rect 9981 10968 10692 10992
rect 6408 10908 7056 10932
rect 7161 10908 7899 10932
rect 8241 10908 9159 10932
rect 9561 10908 9759 10932
rect 10668 10932 10692 10968
rect 12501 10968 13059 10992
rect 13101 10968 15039 10992
rect 15801 10968 16779 10992
rect 17661 10968 18279 10992
rect 10668 10908 11679 10932
rect 13041 10908 13479 10932
rect 13641 10908 14319 10932
rect 18141 10908 18339 10932
rect 4908 10848 5199 10872
rect 5901 10848 7419 10872
rect 8661 10848 9999 10872
rect 10161 10848 10479 10872
rect 10641 10848 10839 10872
rect 10881 10848 12759 10872
rect 15081 10848 15639 10872
rect 15681 10848 15759 10872
rect 17241 10848 17559 10872
rect 621 10788 2259 10812
rect 2901 10788 3219 10812
rect 3561 10788 3699 10812
rect 4701 10788 4839 10812
rect 5301 10788 5679 10812
rect 7341 10788 7479 10812
rect 8001 10788 9516 10812
rect 9621 10788 9699 10812
rect 11001 10788 13539 10812
rect 13941 10788 14379 10812
rect 14721 10788 15819 10812
rect 16701 10788 17139 10812
rect 17841 10788 18279 10812
rect 861 10728 1059 10752
rect 4161 10728 4659 10752
rect 5241 10728 5739 10752
rect 6621 10728 6819 10752
rect 6861 10728 7119 10752
rect 8601 10728 9039 10752
rect 12561 10728 13119 10752
rect 16761 10728 17379 10752
rect 1848 10668 2019 10692
rect 1848 10641 1872 10668
rect 2361 10668 2859 10692
rect 3081 10668 3339 10692
rect 3621 10668 3759 10692
rect 3921 10668 3999 10692
rect 4041 10668 4719 10692
rect 5268 10668 5559 10692
rect 1641 10608 1839 10632
rect 5268 10632 5292 10668
rect 9261 10668 9459 10692
rect 9681 10668 10719 10692
rect 13461 10668 13599 10692
rect 14121 10668 14679 10692
rect 15381 10668 15879 10692
rect 17721 10668 18219 10692
rect 5181 10608 5292 10632
rect 7761 10608 8259 10632
rect 8301 10608 8619 10632
rect 11121 10608 11199 10632
rect 11661 10608 12219 10632
rect 15561 10608 15879 10632
rect 15921 10608 16299 10632
rect 16341 10608 16659 10632
rect 18060 10632 18099 10641
rect 18048 10599 18099 10632
rect 441 10548 699 10572
rect 1341 10551 1479 10575
rect 1608 10548 1899 10572
rect 1608 10512 1632 10548
rect 2541 10551 2739 10575
rect 1548 10488 1632 10512
rect 201 10422 219 10446
rect 261 10422 279 10446
rect 1101 10428 1299 10452
rect 1548 10458 1572 10488
rect 2028 10461 2052 10539
rect 2208 10512 2232 10542
rect 3801 10548 4179 10572
rect 4761 10548 5019 10572
rect 2208 10488 2652 10512
rect 2628 10461 2652 10488
rect 2421 10428 2499 10452
rect 2628 10428 2679 10461
rect 2640 10419 2679 10428
rect 2988 10452 3012 10539
rect 2841 10428 3012 10452
rect 4308 10461 4332 10542
rect 4668 10488 5199 10512
rect 4308 10428 4359 10461
rect 4320 10419 4359 10428
rect 4668 10458 4692 10488
rect 5328 10452 5352 10542
rect 6141 10548 6699 10572
rect 7101 10548 7212 10572
rect 5679 10512 5721 10539
rect 5679 10500 5952 10512
rect 5688 10488 5952 10500
rect 5001 10428 5352 10452
rect 5541 10428 5859 10452
rect 5928 10452 5952 10488
rect 6888 10461 6912 10539
rect 5928 10428 6399 10452
rect 7188 10458 7212 10548
rect 8901 10551 8979 10575
rect 7239 10512 7281 10539
rect 7239 10500 7452 10512
rect 7248 10488 7461 10500
rect 7419 10461 7461 10488
rect 7668 10452 7692 10539
rect 7761 10488 8499 10512
rect 8559 10512 8601 10539
rect 8559 10500 8712 10512
rect 8568 10488 8712 10500
rect 7668 10428 7779 10452
rect 8688 10458 8712 10488
rect 9348 10452 9372 10542
rect 9459 10512 9501 10539
rect 9459 10500 9552 10512
rect 9468 10488 9561 10500
rect 9519 10461 9561 10488
rect 9348 10428 9456 10452
rect 9588 10401 9612 10542
rect 10341 10551 10479 10575
rect 10641 10548 10899 10572
rect 11301 10548 11379 10572
rect 9768 10461 9792 10539
rect 10008 10512 10032 10542
rect 9888 10500 10032 10512
rect 9879 10488 10032 10500
rect 9879 10461 9921 10488
rect 10128 10401 10152 10542
rect 12741 10548 13119 10572
rect 13161 10548 13479 10572
rect 14301 10548 14979 10572
rect 15621 10548 15792 10572
rect 11799 10512 11841 10539
rect 10368 10488 11892 10512
rect 10368 10452 10392 10488
rect 10221 10428 10392 10452
rect 10461 10425 10719 10449
rect 11001 10425 11079 10449
rect 11121 10428 11319 10452
rect 11868 10452 11892 10488
rect 12081 10488 13092 10512
rect 13068 10452 13092 10488
rect 13068 10428 13179 10452
rect 13668 10452 13692 10539
rect 13461 10428 13692 10452
rect 14028 10452 14052 10539
rect 15099 10512 15141 10539
rect 15099 10500 15192 10512
rect 15108 10488 15192 10500
rect 14028 10428 15036 10452
rect 15168 10452 15192 10488
rect 15468 10461 15492 10539
rect 15768 10461 15792 10548
rect 16641 10548 16752 10572
rect 16179 10512 16221 10539
rect 16179 10500 16632 10512
rect 16188 10488 16641 10500
rect 16599 10461 16641 10488
rect 15921 10425 16119 10449
rect 16728 10458 16752 10548
rect 17361 10548 17439 10572
rect 17088 10461 17112 10539
rect 501 10368 699 10392
rect 741 10368 1959 10392
rect 2601 10368 2919 10392
rect 2961 10368 3099 10392
rect 5181 10368 5319 10392
rect 6201 10368 6339 10392
rect 7581 10368 8919 10392
rect 9861 10368 9939 10392
rect 12141 10368 12219 10392
rect 13281 10368 13599 10392
rect 13941 10368 14079 10392
rect 16521 10368 16779 10392
rect 141 10308 1779 10332
rect 2661 10308 2739 10332
rect 3321 10308 3819 10332
rect 3861 10308 4239 10332
rect 4401 10308 4959 10332
rect 5241 10308 5379 10332
rect 5541 10308 5619 10332
rect 6441 10308 6759 10332
rect 6801 10308 7719 10332
rect 8481 10308 8979 10332
rect 9501 10308 9639 10332
rect 10761 10308 11199 10332
rect 13341 10308 14379 10332
rect 16281 10308 16959 10332
rect 17208 10332 17232 10542
rect 17901 10548 17979 10572
rect 17628 10461 17652 10539
rect 18048 10512 18072 10599
rect 17928 10488 18072 10512
rect 18228 10548 18339 10572
rect 17301 10425 17379 10449
rect 17928 10452 17952 10488
rect 18228 10458 18252 10548
rect 17808 10440 17952 10452
rect 17799 10428 17952 10440
rect 17799 10401 17841 10428
rect 17208 10308 17739 10332
rect 1941 10248 2076 10272
rect 2181 10248 2679 10272
rect 5841 10248 6099 10272
rect 6861 10248 7899 10272
rect 8361 10248 9399 10272
rect 9801 10248 10299 10272
rect 11541 10248 12159 10272
rect 15861 10248 16179 10272
rect 16401 10248 17139 10272
rect 17361 10248 17499 10272
rect 381 10188 2259 10212
rect 2601 10188 3039 10212
rect 3501 10188 4119 10212
rect 4461 10188 6039 10212
rect 6261 10188 6639 10212
rect 6801 10188 7539 10212
rect 8841 10188 9339 10212
rect 9381 10188 9579 10212
rect 9621 10188 10419 10212
rect 11781 10188 13239 10212
rect 13581 10188 14439 10212
rect 15261 10188 15399 10212
rect 15801 10188 16299 10212
rect 16581 10188 16659 10212
rect 4641 10128 4839 10152
rect 5721 10128 5979 10152
rect 6981 10128 7116 10152
rect 7221 10128 7299 10152
rect 7701 10128 8199 10152
rect 8721 10128 9039 10152
rect 9801 10128 9879 10152
rect 12681 10128 13719 10152
rect 15801 10128 15999 10152
rect 16041 10128 16359 10152
rect 17181 10128 17259 10152
rect 17601 10128 18039 10152
rect 1161 10068 1599 10092
rect 2301 10068 2979 10092
rect 3141 10068 3339 10092
rect 3501 10068 3699 10092
rect 3741 10068 5619 10092
rect 6081 10068 6759 10092
rect 7401 10068 7599 10092
rect 8181 10068 8319 10092
rect 8541 10068 9852 10092
rect 1281 10008 1419 10032
rect 1881 10008 2139 10032
rect 3801 10008 4659 10032
rect 4881 10008 5259 10032
rect 6081 10008 6579 10032
rect 6621 10008 6819 10032
rect 7041 10008 7479 10032
rect 7701 10008 7779 10032
rect 7821 10008 8019 10032
rect 8781 10008 8919 10032
rect 8961 10008 9219 10032
rect 9441 10008 9639 10032
rect 9828 10032 9852 10068
rect 11628 10068 11979 10092
rect 11628 10041 11652 10068
rect 14361 10068 14679 10092
rect 15141 10068 15399 10092
rect 16761 10068 16899 10092
rect 9828 10008 10179 10032
rect 11421 10008 11619 10032
rect 13281 10008 13419 10032
rect 13461 10008 14199 10032
rect 15681 10008 15939 10032
rect 16881 10008 17139 10032
rect 17541 10008 17619 10032
rect 18201 10008 18339 10032
rect 621 9948 699 9972
rect 3381 9948 3459 9972
rect 5001 9948 5139 9972
rect 5421 9948 5712 9972
rect 141 9888 219 9912
rect 288 9888 459 9912
rect 288 9798 312 9888
rect 861 9888 1119 9912
rect 1761 9888 2139 9912
rect 2181 9888 2292 9912
rect 1068 9828 1359 9852
rect 1068 9798 1092 9828
rect 2268 9852 2292 9888
rect 2361 9891 2439 9915
rect 2721 9888 3072 9912
rect 2268 9828 2352 9852
rect 921 9768 1059 9792
rect 1221 9768 1659 9792
rect 1881 9765 2079 9789
rect 2328 9792 2352 9828
rect 2328 9768 2619 9792
rect 2661 9768 2919 9792
rect 3048 9792 3072 9888
rect 3921 9888 4059 9912
rect 4128 9888 4299 9912
rect 3519 9852 3561 9879
rect 4128 9852 4152 9888
rect 3519 9840 3672 9852
rect 3528 9828 3681 9840
rect 3639 9801 3681 9828
rect 3048 9768 3399 9792
rect 3948 9828 4152 9852
rect 4428 9852 4452 9882
rect 4581 9888 4959 9912
rect 5688 9912 5712 9948
rect 6201 9972 6240 9981
rect 6201 9939 6252 9972
rect 6501 9948 6732 9972
rect 5688 9888 5739 9912
rect 5901 9891 6039 9915
rect 4428 9828 4812 9852
rect 3948 9798 3972 9828
rect 4521 9768 4719 9792
rect 4788 9792 4812 9828
rect 5328 9801 5352 9879
rect 5508 9801 5532 9879
rect 6228 9801 6252 9939
rect 6441 9888 6552 9912
rect 6528 9801 6552 9888
rect 6708 9801 6732 9948
rect 8301 9948 8439 9972
rect 9321 9948 9579 9972
rect 10341 9948 10479 9972
rect 10521 9948 10659 9972
rect 10881 9948 11079 9972
rect 11241 9948 11799 9972
rect 12321 9948 12519 9972
rect 13161 9948 13359 9972
rect 13401 9948 13659 9972
rect 13881 9948 14499 9972
rect 14661 9948 14739 9972
rect 16521 9972 16560 9981
rect 16521 9942 16572 9972
rect 16500 9939 16572 9942
rect 17301 9948 17679 9972
rect 18141 9972 18180 9981
rect 18141 9939 18192 9972
rect 7161 9888 7299 9912
rect 7821 9888 8052 9912
rect 7428 9801 7452 9879
rect 7659 9852 7701 9879
rect 7659 9840 7752 9852
rect 7668 9828 7752 9840
rect 4788 9768 5019 9792
rect 5721 9768 5979 9792
rect 7728 9798 7752 9828
rect 8028 9801 8052 9888
rect 8088 9792 8112 9939
rect 8241 9888 8412 9912
rect 8388 9852 8412 9888
rect 8619 9912 8661 9939
rect 8541 9900 8661 9912
rect 8541 9888 8652 9900
rect 8961 9888 9432 9912
rect 8388 9828 8472 9852
rect 8088 9768 8199 9792
rect 8448 9798 8472 9828
rect 9408 9798 9432 9888
rect 9921 9888 10239 9912
rect 8601 9768 8859 9792
rect 9681 9765 9819 9789
rect 3939 9741 3981 9756
rect 2181 9708 2499 9732
rect 3921 9699 3981 9741
rect 6081 9708 6159 9732
rect 6441 9708 6579 9732
rect 7761 9708 7839 9732
rect 8559 9732 8601 9756
rect 9888 9741 9912 9882
rect 10461 9888 11052 9912
rect 10341 9765 10479 9789
rect 10761 9768 10839 9792
rect 11028 9798 11052 9888
rect 11208 9888 11499 9912
rect 8361 9708 8601 9732
rect 8721 9708 9699 9732
rect 11208 9732 11232 9888
rect 12141 9888 12459 9912
rect 12621 9888 12696 9912
rect 12801 9891 12879 9915
rect 13461 9888 13512 9912
rect 13068 9801 13092 9879
rect 11361 9765 11559 9789
rect 11721 9765 11799 9789
rect 11841 9768 12039 9792
rect 12381 9765 12519 9789
rect 12801 9768 12939 9792
rect 13488 9792 13512 9888
rect 13488 9768 13659 9792
rect 11001 9708 11232 9732
rect 11559 9732 11601 9756
rect 11559 9708 11919 9732
rect 13041 9708 13179 9732
rect 13728 9732 13752 9882
rect 14481 9888 14919 9912
rect 15141 9888 15459 9912
rect 15528 9888 15939 9912
rect 15528 9852 15552 9888
rect 16341 9888 16479 9912
rect 14928 9828 15552 9852
rect 13821 9768 14259 9792
rect 14301 9768 14799 9792
rect 14928 9741 14952 9828
rect 16548 9798 16572 9939
rect 17001 9891 17199 9915
rect 16728 9801 16752 9879
rect 17388 9801 17412 9879
rect 15081 9768 16059 9792
rect 16101 9768 16419 9792
rect 17808 9741 17832 9939
rect 17868 9801 17892 9939
rect 18048 9801 18072 9879
rect 18168 9741 18192 9939
rect 13341 9708 13752 9732
rect 17121 9708 17319 9732
rect 17481 9708 17619 9732
rect 18141 9732 18192 9741
rect 18141 9708 18279 9732
rect 18141 9699 18180 9708
rect 441 9648 579 9672
rect 621 9648 759 9672
rect 1821 9648 2832 9672
rect 2541 9588 2739 9612
rect 2808 9612 2832 9648
rect 3201 9648 3579 9672
rect 5181 9648 6219 9672
rect 7221 9648 7299 9672
rect 8181 9648 8619 9672
rect 8841 9648 9039 9672
rect 9081 9648 9279 9672
rect 10581 9648 11499 9672
rect 12021 9648 12339 9672
rect 12501 9648 13119 9672
rect 13701 9648 13899 9672
rect 14121 9648 14319 9672
rect 15021 9648 15099 9672
rect 15741 9648 15819 9672
rect 16161 9648 16899 9672
rect 17721 9648 17979 9672
rect 2808 9588 3759 9612
rect 4521 9588 4959 9612
rect 5241 9588 5379 9612
rect 5421 9588 6159 9612
rect 6381 9588 6699 9612
rect 6861 9588 6939 9612
rect 8121 9588 8559 9612
rect 9141 9588 9819 9612
rect 10161 9588 10299 9612
rect 14061 9588 14259 9612
rect 15441 9588 16779 9612
rect 17781 9588 18339 9612
rect 1461 9528 2139 9552
rect 5061 9528 6519 9552
rect 6981 9528 7059 9552
rect 7581 9528 8679 9552
rect 9441 9528 9759 9552
rect 11541 9528 12219 9552
rect 12681 9528 14619 9552
rect 14901 9528 15579 9552
rect 15981 9528 16179 9552
rect 16341 9528 16659 9552
rect 17001 9528 17379 9552
rect 17421 9528 17619 9552
rect 981 9468 1299 9492
rect 1341 9468 2319 9492
rect 2361 9468 4059 9492
rect 6081 9468 6459 9492
rect 6501 9468 6759 9492
rect 7821 9468 8319 9492
rect 8361 9468 8439 9492
rect 8841 9468 9939 9492
rect 9981 9468 10179 9492
rect 12381 9468 14679 9492
rect 14841 9468 15279 9492
rect 16041 9468 17259 9492
rect 18021 9468 18219 9492
rect 18261 9468 18339 9492
rect 4281 9408 4899 9432
rect 5121 9408 5559 9432
rect 5601 9408 7119 9432
rect 7401 9408 9099 9432
rect 9261 9408 11499 9432
rect 13101 9408 13539 9432
rect 16101 9408 16719 9432
rect 561 9348 1179 9372
rect 2901 9348 3039 9372
rect 4401 9348 5139 9372
rect 5901 9348 6639 9372
rect 7761 9348 7899 9372
rect 8061 9348 8499 9372
rect 8661 9348 9159 9372
rect 9801 9348 11139 9372
rect 12201 9348 13239 9372
rect 13521 9348 14379 9372
rect 14781 9348 15159 9372
rect 17601 9348 17679 9372
rect 5061 9288 5532 9312
rect 2421 9228 3039 9252
rect 4881 9228 5259 9252
rect 5508 9252 5532 9288
rect 5601 9288 5739 9312
rect 6441 9288 6939 9312
rect 7281 9288 7419 9312
rect 8301 9288 9399 9312
rect 9561 9288 10779 9312
rect 11421 9288 12039 9312
rect 12081 9288 12639 9312
rect 14601 9288 15219 9312
rect 15381 9288 16659 9312
rect 17301 9288 17679 9312
rect 5508 9228 6579 9252
rect 8541 9228 8979 9252
rect 11481 9228 12399 9252
rect 12981 9228 13959 9252
rect 14001 9228 14919 9252
rect 15501 9228 16239 9252
rect 16281 9228 16719 9252
rect 1521 9168 2259 9192
rect 4161 9168 5016 9192
rect 5121 9168 5319 9192
rect 6261 9168 6819 9192
rect 7221 9168 7899 9192
rect 8781 9168 9099 9192
rect 9741 9168 10599 9192
rect 12021 9168 12519 9192
rect 12921 9168 13179 9192
rect 15201 9168 16539 9192
rect 16701 9168 17379 9192
rect 17841 9168 18099 9192
rect 18441 9192 18480 9201
rect 18441 9159 18492 9192
rect 2268 9132 2292 9159
rect 2268 9108 2739 9132
rect 4008 9108 4839 9132
rect 1101 9048 1779 9072
rect 1821 9048 2139 9072
rect 4008 9072 4032 9108
rect 5721 9108 5799 9132
rect 5841 9108 5979 9132
rect 6141 9108 6519 9132
rect 6561 9108 6879 9132
rect 7461 9108 8079 9132
rect 8721 9108 9516 9132
rect 9621 9108 10359 9132
rect 11661 9108 12399 9132
rect 12741 9108 12819 9132
rect 13941 9108 14619 9132
rect 14961 9108 15039 9132
rect 16221 9108 16359 9132
rect 17661 9108 18159 9132
rect 3321 9048 4032 9072
rect 5223 9048 5439 9072
rect 6900 9072 6939 9081
rect 6888 9039 6939 9072
rect 8961 9048 9321 9072
rect 441 8991 519 9015
rect 681 8991 819 9015
rect 1581 8991 1659 9015
rect 1860 9012 1899 9021
rect 1848 8979 1899 9012
rect 2061 8988 2376 9012
rect 2481 8991 2619 9015
rect 2820 9012 2859 9021
rect 2808 8979 2859 9012
rect 3561 8988 3939 9012
rect 4248 8988 4359 9012
rect 1848 8952 1872 8979
rect 1728 8928 1872 8952
rect 141 8865 219 8889
rect 381 8868 879 8892
rect 921 8868 1239 8892
rect 1401 8868 1479 8892
rect 1728 8898 1752 8928
rect 2808 8898 2832 8979
rect 3141 8868 3279 8892
rect 1941 8808 2439 8832
rect 2799 8832 2841 8856
rect 2601 8808 2841 8832
rect 3408 8832 3432 8982
rect 4248 8952 4272 8988
rect 4521 8988 4572 9012
rect 4068 8928 4272 8952
rect 4068 8892 4092 8928
rect 4548 8901 4572 8988
rect 5079 8952 5121 8979
rect 5028 8940 5121 8952
rect 5688 8988 5799 9012
rect 5028 8928 5112 8940
rect 3621 8868 4092 8892
rect 4161 8868 4299 8892
rect 5028 8892 5052 8928
rect 4761 8868 5052 8892
rect 5688 8892 5712 8988
rect 6300 9012 6339 9021
rect 6288 8979 6339 9012
rect 6888 9012 6912 9039
rect 6768 8988 6912 9012
rect 5121 8868 5712 8892
rect 6048 8892 6072 8979
rect 6288 8901 6312 8979
rect 6708 8952 6732 8982
rect 6408 8940 6732 8952
rect 6399 8928 6732 8940
rect 6399 8901 6441 8928
rect 5781 8868 6216 8892
rect 6768 8892 6792 8988
rect 7959 9012 8001 9039
rect 9279 9024 9321 9048
rect 9981 9048 10059 9072
rect 13281 9048 13392 9072
rect 7728 9000 8001 9012
rect 7728 8988 7992 9000
rect 7008 8952 7032 8982
rect 7728 8952 7752 8988
rect 8199 8952 8241 8979
rect 6948 8928 7032 8952
rect 7128 8940 7752 8952
rect 7119 8928 7752 8940
rect 7848 8940 8241 8952
rect 7848 8928 8232 8940
rect 6648 8868 6792 8892
rect 6648 8841 6672 8868
rect 6948 8892 6972 8928
rect 6861 8868 6972 8892
rect 7119 8901 7161 8928
rect 7848 8892 7872 8928
rect 7581 8868 7872 8892
rect 7908 8868 8079 8892
rect 7908 8841 7932 8868
rect 8328 8892 8352 8982
rect 8481 8988 8592 9012
rect 8568 8952 8592 8988
rect 8748 8988 8979 9012
rect 8568 8940 8652 8952
rect 8568 8928 8661 8940
rect 8619 8901 8661 8928
rect 8328 8868 8499 8892
rect 8748 8898 8772 8988
rect 9321 8988 9432 9012
rect 9408 8952 9432 8988
rect 9501 8991 9579 9015
rect 9741 8988 10119 9012
rect 10521 8988 11079 9012
rect 11121 8991 11439 9015
rect 11841 8997 11919 9021
rect 12741 8988 13059 9012
rect 12108 8952 12132 8982
rect 9408 8928 9672 8952
rect 9648 8898 9672 8928
rect 11928 8928 12132 8952
rect 9141 8865 9219 8889
rect 9801 8868 9879 8892
rect 10401 8865 10539 8889
rect 10821 8865 10899 8889
rect 11928 8892 11952 8928
rect 12228 8901 12252 8982
rect 12441 8928 12552 8952
rect 11301 8868 11952 8892
rect 12021 8868 12159 8892
rect 12228 8868 12279 8901
rect 12240 8859 12279 8868
rect 12528 8892 12552 8928
rect 12528 8868 12639 8892
rect 12708 8892 12732 8982
rect 13188 8901 13212 8982
rect 12708 8868 12819 8892
rect 13188 8868 13239 8901
rect 13200 8859 13239 8868
rect 3321 8808 3432 8832
rect 4701 8808 4899 8832
rect 5181 8808 5439 8832
rect 5901 8808 6099 8832
rect 6621 8808 6672 8841
rect 6621 8799 6660 8808
rect 7101 8808 7179 8832
rect 7221 8808 7359 8832
rect 7881 8808 7932 8841
rect 7881 8799 7920 8808
rect 9501 8808 9699 8832
rect 10761 8808 12459 8832
rect 13308 8832 13332 8979
rect 13368 8892 13392 9048
rect 14721 9048 15339 9072
rect 15621 9048 15819 9072
rect 17700 9072 17739 9081
rect 17688 9039 17739 9072
rect 18321 9048 18399 9072
rect 13728 8901 13752 8988
rect 14661 8988 14859 9012
rect 14901 8988 14976 9012
rect 15081 8988 15372 9012
rect 13968 8901 13992 8979
rect 13701 8868 13752 8901
rect 13701 8859 13740 8868
rect 14388 8892 14412 8979
rect 15348 8952 15372 8988
rect 15441 8991 15939 9015
rect 16461 8988 16599 9012
rect 16881 8988 17079 9012
rect 16119 8952 16161 8979
rect 15348 8928 16092 8952
rect 16119 8940 16272 8952
rect 16128 8928 16281 8940
rect 16068 8898 16092 8928
rect 16239 8901 16281 8928
rect 17328 8901 17352 8979
rect 17508 8901 17532 8979
rect 14121 8868 14412 8892
rect 14721 8865 15699 8889
rect 16701 8880 16812 8892
rect 16701 8868 16821 8880
rect 16779 8841 16821 8868
rect 16941 8868 17139 8892
rect 17688 8841 17712 9039
rect 17868 8901 17892 8979
rect 18048 8901 18072 8979
rect 18261 8865 18399 8889
rect 12801 8808 13332 8832
rect 15141 8808 15399 8832
rect 18021 8808 18279 8832
rect 1881 8748 2019 8772
rect 3261 8748 3879 8772
rect 4221 8748 4419 8772
rect 4908 8772 4932 8799
rect 4908 8748 5199 8772
rect 6561 8748 6699 8772
rect 7341 8748 7419 8772
rect 8181 8748 8379 8772
rect 9081 8748 9219 8772
rect 9261 8748 9339 8772
rect 12921 8748 12999 8772
rect 13161 8748 13659 8772
rect 15261 8748 15339 8772
rect 17601 8748 17799 8772
rect 18468 8772 18492 9159
rect 18381 8748 18492 8772
rect 441 8688 819 8712
rect 861 8688 1719 8712
rect 5061 8688 5499 8712
rect 7281 8688 7479 8712
rect 8421 8688 8559 8712
rect 9561 8688 9879 8712
rect 9921 8688 11199 8712
rect 12021 8688 12339 8712
rect 13641 8688 14679 8712
rect 15501 8688 16239 8712
rect 17301 8688 18099 8712
rect 1221 8628 2439 8652
rect 2721 8628 3399 8652
rect 3441 8628 3459 8652
rect 3741 8628 3999 8652
rect 4701 8628 4899 8652
rect 5661 8628 6039 8652
rect 6501 8628 6699 8652
rect 7641 8628 8859 8652
rect 11361 8628 11439 8652
rect 12321 8628 12819 8652
rect 13041 8628 13299 8652
rect 15621 8628 15699 8652
rect 15741 8628 16059 8652
rect 16641 8628 16839 8652
rect 681 8568 759 8592
rect 801 8568 1539 8592
rect 5628 8592 5652 8619
rect 4881 8568 5652 8592
rect 6201 8568 6519 8592
rect 7041 8568 7179 8592
rect 8001 8568 8619 8592
rect 9108 8568 10059 8592
rect 1701 8508 2199 8532
rect 3201 8508 3759 8532
rect 5001 8508 6279 8532
rect 6681 8508 6759 8532
rect 6828 8508 6939 8532
rect 561 8448 999 8472
rect 1521 8448 2919 8472
rect 4041 8448 4659 8472
rect 4821 8448 6159 8472
rect 6348 8448 6399 8472
rect 2361 8388 2559 8412
rect 3561 8388 3921 8412
rect 3879 8364 3921 8388
rect 4521 8400 4632 8412
rect 4521 8388 4641 8400
rect 201 8328 279 8352
rect 681 8352 720 8361
rect 681 8319 732 8352
rect 921 8328 1272 8352
rect 708 8238 732 8319
rect 1248 8238 1272 8328
rect 1341 8328 1659 8352
rect 1821 8328 1872 8352
rect 501 8208 699 8232
rect 1521 8205 1719 8229
rect 1848 8232 1872 8328
rect 2061 8328 2199 8352
rect 2901 8328 2979 8352
rect 3021 8328 3279 8352
rect 2508 8241 2532 8319
rect 3108 8292 3132 8328
rect 3921 8328 4299 8352
rect 4599 8361 4641 8388
rect 6348 8412 6372 8448
rect 6828 8472 6852 8508
rect 9108 8532 9132 8568
rect 10221 8568 10359 8592
rect 11061 8568 11199 8592
rect 12561 8568 12759 8592
rect 13608 8568 13779 8592
rect 13608 8541 13632 8568
rect 14061 8568 14259 8592
rect 14541 8568 15399 8592
rect 15981 8568 16179 8592
rect 17661 8568 17739 8592
rect 17901 8568 18399 8592
rect 8241 8508 9132 8532
rect 9561 8508 12099 8532
rect 12708 8508 13599 8532
rect 6441 8448 6852 8472
rect 6921 8448 7512 8472
rect 5421 8388 6372 8412
rect 6561 8388 6819 8412
rect 7488 8412 7512 8448
rect 7581 8448 7659 8472
rect 8721 8448 8919 8472
rect 11301 8448 11799 8472
rect 12708 8472 12732 8508
rect 14241 8508 14319 8532
rect 14388 8508 15519 8532
rect 12528 8448 12732 8472
rect 7488 8388 8199 8412
rect 9981 8388 10239 8412
rect 12528 8412 12552 8448
rect 12801 8448 12939 8472
rect 13581 8448 13659 8472
rect 14001 8448 14139 8472
rect 14388 8472 14412 8508
rect 16461 8508 16659 8532
rect 16881 8508 17139 8532
rect 14208 8448 14412 8472
rect 14208 8412 14232 8448
rect 14481 8448 14739 8472
rect 15048 8448 15519 8472
rect 15048 8412 15072 8448
rect 15801 8448 16299 8472
rect 17421 8448 17499 8472
rect 18081 8448 18159 8472
rect 12381 8388 12552 8412
rect 13968 8388 14232 8412
rect 14808 8388 15072 8412
rect 5361 8331 5499 8355
rect 6321 8331 6399 8355
rect 7281 8328 7812 8352
rect 3108 8268 3192 8292
rect 1848 8208 2259 8232
rect 2928 8220 3039 8232
rect 2919 8208 3039 8220
rect 2919 8181 2961 8208
rect 3168 8232 3192 8268
rect 4728 8241 4752 8319
rect 4968 8268 5412 8292
rect 3168 8208 3339 8232
rect 4521 8205 4599 8229
rect 4968 8232 4992 8268
rect 4881 8208 4992 8232
rect 5388 8238 5412 8268
rect 5919 8292 5961 8319
rect 7059 8292 7101 8319
rect 5601 8280 5961 8292
rect 6948 8280 7101 8292
rect 7788 8292 7812 8328
rect 7881 8328 8079 8352
rect 8148 8328 8499 8352
rect 5601 8268 5952 8280
rect 6948 8268 7092 8280
rect 7788 8268 7872 8292
rect 5121 8208 5259 8232
rect 6021 8220 6072 8232
rect 6021 8208 6081 8220
rect 381 8148 939 8172
rect 981 8148 1059 8172
rect 5061 8148 5196 8172
rect 5259 8172 5301 8196
rect 6039 8181 6081 8208
rect 6948 8232 6972 8268
rect 6381 8208 6972 8232
rect 7041 8208 7299 8232
rect 7848 8232 7872 8268
rect 8148 8292 8172 8328
rect 8781 8328 9039 8352
rect 10101 8328 10179 8352
rect 7941 8268 8172 8292
rect 10068 8241 10092 8322
rect 10521 8328 10839 8352
rect 11001 8328 11139 8352
rect 11481 8331 11619 8355
rect 7848 8208 8019 8232
rect 5259 8148 5619 8172
rect 6501 8148 7239 8172
rect 7848 8172 7872 8208
rect 8181 8205 8319 8229
rect 8601 8208 8679 8232
rect 9021 8205 9699 8229
rect 10041 8208 10092 8241
rect 10041 8199 10080 8208
rect 10308 8232 10332 8319
rect 10221 8208 10539 8232
rect 10581 8205 11079 8229
rect 11328 8232 11352 8319
rect 11928 8241 11952 8379
rect 12501 8328 12579 8352
rect 12741 8328 12792 8352
rect 11328 8208 11379 8232
rect 11541 8205 11619 8229
rect 11661 8205 11739 8229
rect 11928 8208 11979 8241
rect 11940 8199 11979 8208
rect 12288 8232 12312 8319
rect 12261 8208 12312 8232
rect 12768 8241 12792 8328
rect 12861 8328 13152 8352
rect 12768 8208 12819 8241
rect 12780 8199 12819 8208
rect 13128 8238 13152 8328
rect 13401 8328 13539 8352
rect 13608 8328 13899 8352
rect 13608 8238 13632 8328
rect 13968 8352 13992 8388
rect 13941 8328 13992 8352
rect 14268 8328 14319 8352
rect 14088 8241 14112 8319
rect 14268 8241 14292 8328
rect 14508 8241 14532 8319
rect 13341 8208 13599 8232
rect 13761 8208 13959 8232
rect 14808 8232 14832 8388
rect 15228 8400 15459 8412
rect 15099 8352 15141 8379
rect 15219 8388 15459 8400
rect 15219 8361 15261 8388
rect 16401 8388 16659 8412
rect 16701 8388 16839 8412
rect 17901 8388 17979 8412
rect 15099 8340 15192 8352
rect 15108 8328 15192 8340
rect 15168 8241 15192 8328
rect 15288 8328 15759 8352
rect 14781 8208 14832 8232
rect 7581 8148 7872 8172
rect 9981 8148 10419 8172
rect 14481 8148 14559 8172
rect 14601 8148 14859 8172
rect 15288 8178 15312 8328
rect 15921 8328 16059 8352
rect 16248 8328 16419 8352
rect 16248 8241 16272 8328
rect 17319 8352 17361 8379
rect 17319 8340 17559 8352
rect 17328 8328 17559 8340
rect 17328 8292 17352 8328
rect 16908 8280 17352 8292
rect 16899 8268 17352 8280
rect 16899 8241 16941 8268
rect 15501 8208 15939 8232
rect 16521 8205 16659 8229
rect 17481 8208 17619 8232
rect 17688 8232 17712 8319
rect 17688 8208 18039 8232
rect 15948 8172 15972 8196
rect 16479 8172 16521 8196
rect 15948 8148 16521 8172
rect 16821 8148 17079 8172
rect 1581 8088 2739 8112
rect 4401 8088 4959 8112
rect 5541 8088 5679 8112
rect 6801 8088 7299 8112
rect 7641 8088 8259 8112
rect 8481 8088 8739 8112
rect 8781 8088 8859 8112
rect 11601 8088 11799 8112
rect 12141 8088 12639 8112
rect 13281 8088 13719 8112
rect 13788 8088 14379 8112
rect 81 8028 459 8052
rect 921 8028 999 8052
rect 3021 8028 3219 8052
rect 3261 8028 3459 8052
rect 3501 8028 4239 8052
rect 6081 8028 7359 8052
rect 7401 8028 7479 8052
rect 7701 8028 7899 8052
rect 8961 8028 9819 8052
rect 10881 8028 11259 8052
rect 13788 8052 13812 8088
rect 15621 8088 16059 8112
rect 12801 8028 13812 8052
rect 14088 8028 14439 8052
rect 2061 7968 5352 7992
rect 681 7908 4899 7932
rect 5328 7932 5352 7968
rect 5601 7968 5679 7992
rect 6501 7968 7719 7992
rect 7788 7980 8079 7992
rect 7779 7968 8079 7980
rect 7779 7941 7821 7968
rect 8421 7968 8679 7992
rect 8901 7968 9279 7992
rect 11601 7968 11979 7992
rect 14088 7992 14112 8028
rect 14781 8028 14859 8052
rect 12021 7968 14112 7992
rect 16821 7968 16959 7992
rect 17001 7968 18039 7992
rect 18081 7968 18219 7992
rect 5328 7908 6819 7932
rect 6861 7908 7119 7932
rect 8181 7908 9939 7932
rect 10161 7908 10899 7932
rect 11121 7908 13299 7932
rect 14181 7908 14859 7932
rect 16401 7908 17439 7932
rect 2001 7848 2199 7872
rect 2481 7848 3819 7872
rect 6141 7848 6639 7872
rect 7701 7848 8079 7872
rect 12561 7848 13359 7872
rect 13941 7848 15399 7872
rect 15441 7848 15699 7872
rect 17781 7848 18039 7872
rect 201 7788 1539 7812
rect 2661 7788 3939 7812
rect 5121 7788 5439 7812
rect 5601 7788 5739 7812
rect 6261 7788 6939 7812
rect 7281 7788 8559 7812
rect 9381 7788 9879 7812
rect 10161 7788 10719 7812
rect 11301 7788 13839 7812
rect 14841 7788 15219 7812
rect 17661 7788 18399 7812
rect 81 7728 2139 7752
rect 4221 7728 4659 7752
rect 5001 7728 5379 7752
rect 6441 7728 7239 7752
rect 8121 7728 8379 7752
rect 8841 7728 9159 7752
rect 9681 7728 9939 7752
rect 12261 7728 12999 7752
rect 13041 7728 13179 7752
rect 13641 7728 14079 7752
rect 17301 7728 17739 7752
rect 18021 7728 18159 7752
rect 861 7668 1419 7692
rect 1461 7668 1899 7692
rect 2181 7668 2499 7692
rect 2961 7668 4119 7692
rect 4161 7668 4719 7692
rect 5481 7668 6699 7692
rect 7341 7668 8019 7692
rect 8601 7668 9999 7692
rect 11361 7668 11859 7692
rect 11901 7668 13179 7692
rect 13221 7668 13479 7692
rect 13521 7668 14259 7692
rect 14301 7668 14979 7692
rect 15681 7668 15999 7692
rect 16161 7668 16599 7692
rect 17328 7668 17499 7692
rect 17328 7641 17352 7668
rect 801 7608 2679 7632
rect 3141 7608 3339 7632
rect 3561 7608 4272 7632
rect 4248 7581 4272 7608
rect 4821 7608 5259 7632
rect 5541 7608 6399 7632
rect 6921 7608 7539 7632
rect 9861 7608 10059 7632
rect 10281 7608 11259 7632
rect 12081 7608 12279 7632
rect 12981 7608 13359 7632
rect 13881 7608 14919 7632
rect 15801 7608 16299 7632
rect 16908 7608 17319 7632
rect 141 7548 639 7572
rect 1221 7548 2259 7572
rect 2301 7548 2439 7572
rect 2841 7548 3399 7572
rect 4281 7548 5439 7572
rect 7581 7548 8139 7572
rect 8541 7548 9219 7572
rect 13521 7548 13899 7572
rect 16908 7572 16932 7608
rect 18201 7608 18399 7632
rect 15561 7548 16932 7572
rect 3621 7488 3759 7512
rect 4521 7488 5139 7512
rect 5361 7488 5859 7512
rect 6108 7488 6279 7512
rect 261 7428 372 7452
rect 348 7341 372 7428
rect 441 7428 759 7452
rect 1101 7428 1359 7452
rect 1401 7428 1539 7452
rect 3081 7431 3159 7455
rect 1908 7392 1932 7422
rect 1761 7368 1932 7392
rect 2028 7341 2052 7422
rect 3741 7431 3939 7455
rect 4881 7431 5079 7455
rect 5481 7428 5676 7452
rect 2028 7308 2079 7341
rect 2040 7299 2079 7308
rect 3141 7308 3999 7332
rect 4161 7308 5079 7332
rect 5268 7338 5292 7419
rect 5448 7392 5472 7422
rect 5448 7368 5652 7392
rect 5301 7305 5499 7329
rect 201 7248 516 7272
rect 621 7248 1239 7272
rect 2061 7248 2139 7272
rect 3081 7248 3159 7272
rect 4581 7248 4899 7272
rect 5181 7248 5379 7272
rect 5628 7272 5652 7368
rect 5748 7341 5772 7422
rect 6108 7392 6132 7488
rect 6441 7488 6579 7512
rect 6621 7488 7059 7512
rect 7608 7488 7899 7512
rect 6801 7452 6840 7461
rect 6801 7419 6852 7452
rect 7341 7428 7419 7452
rect 6459 7392 6501 7419
rect 6021 7368 6132 7392
rect 6288 7380 6501 7392
rect 6288 7368 6492 7380
rect 5721 7308 5772 7341
rect 5721 7299 5760 7308
rect 5961 7308 6039 7332
rect 6288 7338 6312 7368
rect 6648 7332 6672 7419
rect 6648 7308 6759 7332
rect 5628 7248 5739 7272
rect 6828 7272 6852 7419
rect 7008 7341 7032 7419
rect 7608 7338 7632 7488
rect 8301 7488 9099 7512
rect 9468 7488 9879 7512
rect 7881 7431 8019 7455
rect 8721 7428 8919 7452
rect 8139 7392 8181 7419
rect 8139 7380 8799 7392
rect 8148 7368 8799 7380
rect 9048 7341 9072 7422
rect 7221 7305 7299 7329
rect 8301 7302 8376 7326
rect 8481 7320 8772 7332
rect 8481 7308 8781 7320
rect 6681 7248 6852 7272
rect 8739 7281 8781 7308
rect 9021 7308 9072 7341
rect 9021 7299 9060 7308
rect 9468 7332 9492 7488
rect 10521 7488 10659 7512
rect 12141 7488 12339 7512
rect 12381 7488 12459 7512
rect 13701 7488 13779 7512
rect 14268 7488 14499 7512
rect 9561 7428 9852 7452
rect 9828 7338 9852 7428
rect 10041 7431 10179 7455
rect 10401 7428 10452 7452
rect 10428 7341 10452 7428
rect 10728 7392 10752 7422
rect 11241 7428 11499 7452
rect 11568 7428 11679 7452
rect 11568 7392 11592 7428
rect 12681 7431 12819 7455
rect 13008 7428 13179 7452
rect 10581 7368 10752 7392
rect 11388 7368 11592 7392
rect 9261 7308 9492 7332
rect 11388 7338 11412 7368
rect 12228 7338 12252 7419
rect 11061 7308 11259 7332
rect 12081 7305 12219 7329
rect 13008 7338 13032 7428
rect 13401 7428 13572 7452
rect 13548 7401 13572 7428
rect 14268 7452 14292 7488
rect 14541 7488 14619 7512
rect 16521 7488 16659 7512
rect 16941 7488 17079 7512
rect 17121 7488 17199 7512
rect 17421 7512 17460 7521
rect 17421 7479 17472 7512
rect 17601 7488 17799 7512
rect 14028 7428 14292 7452
rect 13548 7368 13599 7401
rect 13560 7359 13599 7368
rect 12381 7308 12852 7332
rect 9141 7248 9219 7272
rect 2301 7188 2559 7212
rect 2721 7188 3279 7212
rect 3441 7188 4119 7212
rect 5028 7188 5199 7212
rect 5028 7161 5052 7188
rect 5661 7188 5799 7212
rect 6648 7212 6672 7239
rect 9981 7248 10539 7272
rect 12201 7248 12459 7272
rect 12828 7272 12852 7308
rect 13161 7305 13239 7329
rect 13788 7332 13812 7419
rect 13461 7308 13812 7332
rect 14028 7332 14052 7428
rect 14361 7428 14472 7452
rect 14448 7401 14472 7428
rect 14448 7368 14499 7401
rect 14460 7359 14499 7368
rect 14988 7341 15012 7419
rect 14001 7308 14052 7332
rect 14121 7305 14379 7329
rect 15168 7338 15192 7479
rect 15228 7341 15252 7422
rect 15441 7452 15480 7461
rect 15441 7419 15492 7452
rect 15228 7308 15279 7341
rect 15240 7299 15279 7308
rect 15468 7338 15492 7419
rect 15828 7428 15879 7452
rect 15828 7341 15852 7428
rect 16008 7281 16032 7422
rect 16281 7428 16392 7452
rect 16119 7392 16161 7419
rect 16068 7380 16161 7392
rect 16068 7368 16152 7380
rect 16068 7338 16092 7368
rect 16368 7338 16392 7428
rect 16539 7392 16581 7419
rect 16428 7380 16581 7392
rect 16419 7368 16572 7380
rect 16419 7341 16461 7368
rect 16641 7308 16839 7332
rect 17148 7332 17172 7419
rect 17448 7392 17472 7479
rect 17448 7380 17652 7392
rect 17448 7368 17661 7380
rect 17619 7341 17661 7368
rect 17988 7341 18012 7419
rect 18228 7341 18252 7419
rect 17061 7308 17172 7332
rect 17421 7305 17499 7329
rect 17841 7308 17919 7332
rect 12828 7248 13059 7272
rect 14181 7248 14259 7272
rect 15801 7248 15936 7272
rect 16701 7248 16779 7272
rect 17121 7248 17199 7272
rect 6201 7188 6672 7212
rect 7041 7188 8139 7212
rect 8961 7188 10659 7212
rect 11781 7188 14859 7212
rect 14901 7188 15219 7212
rect 17001 7188 17139 7212
rect 17181 7188 17499 7212
rect 17721 7188 18039 7212
rect 18201 7188 18279 7212
rect 141 7128 279 7152
rect 801 7128 879 7152
rect 1461 7128 1599 7152
rect 1641 7128 1839 7152
rect 1881 7128 2139 7152
rect 2181 7128 3339 7152
rect 3501 7128 3699 7152
rect 4821 7128 5019 7152
rect 5241 7128 5559 7152
rect 5901 7128 6939 7152
rect 7521 7128 8559 7152
rect 8601 7128 9399 7152
rect 11901 7128 12039 7152
rect 13101 7128 13959 7152
rect 14781 7128 15339 7152
rect 15801 7128 18099 7152
rect 2241 7068 2379 7092
rect 2421 7068 3216 7092
rect 3321 7068 4419 7092
rect 4701 7068 5919 7092
rect 6081 7068 6276 7092
rect 6381 7068 7479 7092
rect 7521 7068 7779 7092
rect 8001 7068 8499 7092
rect 8961 7068 9339 7092
rect 12621 7068 12999 7092
rect 14961 7068 15879 7092
rect 16521 7068 17919 7092
rect 18321 7068 18399 7092
rect 261 7008 339 7032
rect 621 7008 879 7032
rect 921 7008 1059 7032
rect 1221 7008 1719 7032
rect 1761 7008 2739 7032
rect 2781 7008 2859 7032
rect 4041 7008 4179 7032
rect 4401 7008 4959 7032
rect 5121 7008 5472 7032
rect 5448 6981 5472 7008
rect 5661 7008 5739 7032
rect 5781 7008 7059 7032
rect 8061 7008 10839 7032
rect 11001 7008 11199 7032
rect 12201 7008 12819 7032
rect 13461 7008 13599 7032
rect 14181 7008 14439 7032
rect 15021 7008 15159 7032
rect 15381 7008 15759 7032
rect 16101 7008 16419 7032
rect 16821 7008 16959 7032
rect 2901 6948 3099 6972
rect 3561 6948 3819 6972
rect 3861 6948 4239 6972
rect 4281 6948 5079 6972
rect 5481 6948 6339 6972
rect 7461 6948 7779 6972
rect 8541 6948 8979 6972
rect 9021 6948 9099 6972
rect 9168 6948 10119 6972
rect 381 6888 759 6912
rect 1161 6888 1392 6912
rect 1368 6861 1392 6888
rect 2541 6888 3459 6912
rect 3621 6888 4332 6912
rect 4308 6861 4332 6888
rect 5001 6888 5259 6912
rect 5421 6888 6039 6912
rect 6621 6888 7236 6912
rect 7341 6888 8139 6912
rect 9168 6912 9192 6948
rect 10161 6948 10539 6972
rect 11499 6972 11541 6999
rect 11499 6960 12339 6972
rect 11508 6948 12339 6960
rect 12501 6948 12579 6972
rect 12621 6948 12879 6972
rect 14481 6948 15279 6972
rect 15321 6948 15459 6972
rect 15501 6948 15819 6972
rect 15861 6948 16719 6972
rect 17601 6948 17739 6972
rect 17901 6948 18039 6972
rect 18201 6948 18339 6972
rect 8481 6888 9192 6912
rect 10641 6888 11619 6912
rect 981 6828 1059 6852
rect 1401 6828 1539 6852
rect 2061 6828 2259 6852
rect -72 6768 99 6792
rect 501 6771 699 6795
rect 321 6645 699 6669
rect 828 6621 852 6819
rect 2541 6828 2619 6852
rect 4341 6828 4479 6852
rect 4521 6828 4899 6852
rect 5841 6828 6039 6852
rect 1221 6792 1260 6801
rect 1221 6759 1272 6792
rect 1341 6768 1392 6792
rect 1248 6678 1272 6759
rect 981 6645 1119 6669
rect 1368 6621 1392 6768
rect 1881 6768 1959 6792
rect 2121 6768 3039 6792
rect 3201 6768 3519 6792
rect 3681 6768 3999 6792
rect 4041 6768 4512 6792
rect 2088 6681 2112 6759
rect 1581 6645 1659 6669
rect 2361 6648 2679 6672
rect 2841 6648 2919 6672
rect 3741 6645 3819 6669
rect 3981 6648 4419 6672
rect 4488 6672 4512 6768
rect 5181 6771 5319 6795
rect 5565 6681 5589 6819
rect 6921 6828 7119 6852
rect 10281 6828 10479 6852
rect 10701 6828 10779 6852
rect 11841 6828 12192 6852
rect 6321 6768 6456 6792
rect 5679 6732 5721 6759
rect 5628 6720 5721 6732
rect 5628 6708 5712 6720
rect 5628 6681 5652 6708
rect 5868 6681 5892 6759
rect 6759 6792 6801 6819
rect 6561 6780 6801 6792
rect 6561 6768 6792 6780
rect 8721 6771 8799 6795
rect 9021 6771 9219 6795
rect 9561 6768 9819 6792
rect 10101 6771 10179 6795
rect 10881 6768 10959 6792
rect 11520 6792 11559 6801
rect 5988 6720 7299 6732
rect 5979 6708 7299 6720
rect 5979 6681 6021 6708
rect 10419 6732 10461 6759
rect 11508 6759 11559 6792
rect 11961 6771 12099 6795
rect 10419 6720 10572 6732
rect 10428 6708 10581 6720
rect 4488 6648 4536 6672
rect 4641 6648 4959 6672
rect 5661 6648 5739 6672
rect 6261 6660 6609 6672
rect 6648 6660 7899 6672
rect 6261 6648 6621 6660
rect 6579 6621 6621 6648
rect -72 6588 219 6612
rect 828 6588 879 6621
rect 840 6579 879 6588
rect 1341 6588 1392 6621
rect 1341 6579 1380 6588
rect 4161 6588 4299 6612
rect 5301 6588 5379 6612
rect 6618 6600 6621 6621
rect 6639 6648 7899 6660
rect 6639 6621 6681 6648
rect 8139 6672 8181 6699
rect 10539 6681 10581 6708
rect 8139 6660 8259 6672
rect 8148 6648 8259 6660
rect 8781 6648 8979 6672
rect 11508 6672 11532 6759
rect 12168 6732 12192 6828
rect 12321 6828 12639 6852
rect 12759 6828 14619 6852
rect 12759 6804 12801 6828
rect 14961 6828 15039 6852
rect 15261 6828 15639 6852
rect 18021 6828 18159 6852
rect 12768 6732 12792 6762
rect 13101 6768 13272 6792
rect 12939 6732 12981 6759
rect 11661 6708 12012 6732
rect 12168 6708 12792 6732
rect 12828 6720 12981 6732
rect 13248 6732 13272 6768
rect 13341 6771 13719 6795
rect 13860 6792 13899 6801
rect 13848 6759 13899 6792
rect 14361 6771 14499 6795
rect 16341 6768 16539 6792
rect 16581 6771 16659 6795
rect 13248 6720 13452 6732
rect 12828 6708 12972 6720
rect 13248 6708 13461 6720
rect 11988 6678 12012 6708
rect 11721 6648 11859 6672
rect 12708 6672 12732 6708
rect 12828 6678 12852 6708
rect 13419 6681 13461 6708
rect 12441 6648 12732 6672
rect 13848 6672 13872 6759
rect 15108 6708 15279 6732
rect 15108 6678 15132 6708
rect 16008 6681 16032 6759
rect 15648 6648 15912 6672
rect 7101 6588 7659 6612
rect 8241 6588 8319 6612
rect 9201 6588 9459 6612
rect 9861 6588 10599 6612
rect 10761 6588 12279 6612
rect 15648 6612 15672 6648
rect 15441 6588 15672 6612
rect 15888 6612 15912 6648
rect 16728 6678 16752 6819
rect 16821 6768 16872 6792
rect 16068 6648 16359 6672
rect 16068 6612 16092 6648
rect 16848 6621 16872 6768
rect 17361 6768 17472 6792
rect 17448 6681 17472 6768
rect 17748 6681 17772 6759
rect 18048 6681 18072 6759
rect 15888 6588 16092 6612
rect 16821 6588 16872 6621
rect 16821 6579 16860 6588
rect 741 6528 999 6552
rect 1821 6528 2079 6552
rect 2241 6528 2559 6552
rect 3261 6528 3459 6552
rect 3501 6528 3939 6552
rect 5001 6528 5139 6552
rect 5721 6528 6819 6552
rect 7041 6528 7899 6552
rect 9561 6528 9699 6552
rect 10821 6528 11739 6552
rect 11901 6528 12039 6552
rect 14601 6528 15099 6552
rect 15861 6528 16119 6552
rect 16581 6528 17199 6552
rect 2208 6492 2232 6519
rect 1401 6468 2232 6492
rect 3381 6468 3579 6492
rect 3861 6468 4179 6492
rect 4821 6468 5199 6492
rect 6141 6468 6699 6492
rect 6921 6468 7059 6492
rect 7281 6468 7839 6492
rect 8961 6468 9759 6492
rect 11181 6468 11619 6492
rect 11841 6468 13119 6492
rect 13821 6468 14379 6492
rect 16341 6468 16959 6492
rect 681 6408 2319 6432
rect 4248 6408 4599 6432
rect 441 6348 579 6372
rect 861 6348 1779 6372
rect 4248 6372 4272 6408
rect 4881 6408 5019 6432
rect 5961 6408 6972 6432
rect 3981 6348 4272 6372
rect 4308 6348 4839 6372
rect 4308 6312 4332 6348
rect 5721 6348 6639 6372
rect 6948 6372 6972 6408
rect 7341 6408 8859 6432
rect 11361 6408 11559 6432
rect 13881 6408 14499 6432
rect 6948 6348 7239 6372
rect 7281 6348 7419 6372
rect 7581 6348 9939 6372
rect 11781 6348 12219 6372
rect 13401 6348 13479 6372
rect 16281 6348 17319 6372
rect 141 6288 4332 6312
rect 4908 6288 5112 6312
rect 261 6228 4179 6252
rect 4908 6252 4932 6288
rect 4821 6228 4932 6252
rect 5088 6252 5112 6288
rect 5181 6288 5499 6312
rect 5541 6288 5976 6312
rect 6081 6288 7119 6312
rect 7701 6288 8019 6312
rect 9681 6288 10719 6312
rect 13041 6288 13839 6312
rect 14181 6288 14799 6312
rect 15381 6288 16119 6312
rect 16761 6288 17559 6312
rect 5088 6228 5919 6252
rect 6141 6228 6276 6252
rect 6381 6228 6459 6252
rect 7641 6228 8259 6252
rect 8301 6228 10359 6252
rect 10821 6228 11979 6252
rect 12021 6228 12639 6252
rect 13281 6228 13779 6252
rect 15801 6228 16059 6252
rect 921 6168 1779 6192
rect 3141 6168 4239 6192
rect 4641 6168 4719 6192
rect 5001 6168 6699 6192
rect 7401 6168 7539 6192
rect 10221 6168 14259 6192
rect 15261 6168 15879 6192
rect 16221 6168 16719 6192
rect 17061 6168 17799 6192
rect 2721 6108 4059 6132
rect 4401 6108 4776 6132
rect 4881 6108 6099 6132
rect 6321 6108 6459 6132
rect 6681 6108 7299 6132
rect 10701 6108 10959 6132
rect 13608 6108 14139 6132
rect 321 6048 879 6072
rect 1641 6048 1839 6072
rect 2121 6048 2319 6072
rect 6261 6048 6999 6072
rect 2421 5988 2739 6012
rect 3021 5988 3492 6012
rect 3468 5961 3492 5988
rect 4461 5988 5139 6012
rect 6459 6018 6501 6048
rect 7401 6048 8139 6072
rect 8181 6048 9639 6072
rect 9681 6048 10152 6072
rect 10128 6021 10152 6048
rect 13608 6072 13632 6108
rect 12501 6048 13152 6072
rect 6741 5988 6852 6012
rect 1221 5928 1479 5952
rect 1521 5928 2319 5952
rect 3501 5928 3939 5952
rect 6261 5928 6339 5952
rect 6828 5952 6852 5988
rect 6921 5988 7179 6012
rect 7641 5988 10056 6012
rect 10161 5988 10539 6012
rect 12801 5988 12939 6012
rect 13128 6012 13152 6048
rect 13548 6048 13632 6072
rect 13128 5988 13419 6012
rect 7299 5952 7341 5979
rect 6828 5940 7341 5952
rect 6828 5928 7332 5940
rect 7821 5928 8559 5952
rect 10701 5928 10899 5952
rect 11028 5928 11739 5952
rect 348 5721 372 5862
rect 921 5868 972 5892
rect 528 5781 552 5859
rect 768 5772 792 5862
rect 948 5781 972 5868
rect 1341 5868 1599 5892
rect 1938 5859 1941 5880
rect 2001 5868 2259 5892
rect 1068 5781 1092 5859
rect 1899 5832 1941 5859
rect 2448 5832 2472 5862
rect 1899 5820 1992 5832
rect 2388 5820 2472 5832
rect 1908 5808 1992 5820
rect 1968 5781 1992 5808
rect 681 5748 792 5772
rect 1281 5748 1539 5772
rect 1581 5745 1779 5769
rect 1941 5772 1992 5781
rect 2379 5808 2472 5820
rect 2379 5781 2421 5808
rect 1941 5748 2019 5772
rect 1941 5739 1980 5748
rect 2568 5721 2592 5862
rect 2901 5871 3099 5895
rect 3741 5871 3819 5895
rect 4020 5892 4059 5901
rect 2679 5832 2721 5859
rect 2628 5820 2721 5832
rect 2628 5808 2712 5820
rect 2628 5778 2652 5808
rect 2781 5748 2919 5772
rect 3348 5772 3372 5862
rect 4008 5859 4059 5892
rect 4521 5868 4599 5892
rect 4881 5871 5079 5895
rect 5601 5868 5772 5892
rect 4008 5778 4032 5859
rect 4179 5832 4221 5859
rect 4179 5820 5679 5832
rect 4188 5808 5679 5820
rect 5748 5832 5772 5868
rect 5841 5868 6279 5892
rect 6441 5871 6699 5895
rect 6741 5868 7416 5892
rect 7581 5871 7719 5895
rect 8781 5871 8859 5895
rect 9081 5871 9219 5895
rect 9801 5871 9879 5895
rect 10101 5871 10239 5895
rect 11028 5892 11052 5928
rect 12519 5952 12561 5979
rect 13548 5961 13572 6048
rect 13701 6048 13839 6072
rect 14661 6048 16359 6072
rect 17361 6048 17859 6072
rect 17901 6048 18099 6072
rect 15561 5988 16179 6012
rect 16941 5988 17019 6012
rect 12321 5940 12561 5952
rect 12321 5928 12552 5940
rect 12783 5928 12999 5952
rect 13548 5928 13599 5961
rect 13560 5919 13599 5928
rect 13941 5928 14199 5952
rect 14721 5928 14919 5952
rect 15081 5928 15279 5952
rect 16641 5928 16779 5952
rect 17421 5928 17559 5952
rect 10281 5868 11052 5892
rect 11121 5868 11379 5892
rect 11541 5871 11679 5895
rect 5748 5808 6939 5832
rect 8028 5781 8052 5862
rect 11868 5832 11892 5862
rect 8301 5808 8952 5832
rect 3081 5748 3372 5772
rect 3561 5748 3999 5772
rect 4941 5748 5859 5772
rect 7341 5745 7479 5769
rect 8001 5748 8052 5781
rect 8928 5778 8952 5808
rect 10848 5808 11892 5832
rect 8001 5739 8040 5748
rect 9501 5748 9579 5772
rect 9621 5745 9699 5769
rect 10848 5772 10872 5808
rect 10641 5748 10872 5772
rect 10941 5745 11139 5769
rect 12141 5748 12279 5772
rect 12648 5772 12672 5859
rect 12828 5832 12852 5862
rect 12828 5808 12912 5832
rect 12888 5781 12912 5808
rect 13041 5832 13080 5841
rect 13041 5820 13092 5832
rect 13041 5799 13101 5820
rect 13059 5781 13101 5799
rect 12648 5748 12759 5772
rect 12888 5748 12939 5781
rect 12900 5739 12939 5748
rect 621 5688 1119 5712
rect 5301 5688 6159 5712
rect 6741 5688 7179 5712
rect 8661 5688 8739 5712
rect 8781 5688 8916 5712
rect 9021 5688 9879 5712
rect 13041 5688 13119 5712
rect 13188 5712 13212 5862
rect 13308 5772 13332 5862
rect 13821 5868 13959 5892
rect 14421 5868 14652 5892
rect 13308 5748 13659 5772
rect 14088 5772 14112 5862
rect 14628 5832 14652 5868
rect 14808 5832 14832 5862
rect 15219 5832 15261 5859
rect 14628 5808 14832 5832
rect 14088 5748 14199 5772
rect 14481 5760 14532 5772
rect 14481 5748 14541 5760
rect 14499 5721 14541 5748
rect 14808 5721 14832 5808
rect 15108 5820 15261 5832
rect 15468 5868 15579 5892
rect 15108 5808 15252 5820
rect 15108 5772 15132 5808
rect 14901 5748 15132 5772
rect 15468 5772 15492 5868
rect 15381 5748 15492 5772
rect 15825 5772 15849 5859
rect 15681 5748 15849 5772
rect 15888 5721 15912 5862
rect 13188 5688 13299 5712
rect 15201 5688 15279 5712
rect 15861 5688 15912 5721
rect 16008 5712 16032 5862
rect 16521 5868 16659 5892
rect 17001 5871 17199 5895
rect 17661 5868 17739 5892
rect 16299 5832 16341 5859
rect 16299 5820 16779 5832
rect 16308 5808 16779 5820
rect 16101 5748 16236 5772
rect 16341 5745 16419 5769
rect 16581 5745 16719 5769
rect 16881 5748 17019 5772
rect 17301 5748 17799 5772
rect 17841 5745 18219 5769
rect 16008 5688 16359 5712
rect 15861 5679 15900 5688
rect 17421 5688 17619 5712
rect 1188 5628 1659 5652
rect 141 5568 279 5592
rect 441 5568 999 5592
rect 1188 5592 1212 5628
rect 2361 5628 2499 5652
rect 3261 5628 3399 5652
rect 3981 5628 4119 5652
rect 4641 5628 5079 5652
rect 5961 5628 6099 5652
rect 7668 5628 9339 5652
rect 7668 5601 7692 5628
rect 9501 5628 10599 5652
rect 10641 5628 11319 5652
rect 11721 5628 11919 5652
rect 11961 5628 12639 5652
rect 12681 5628 12879 5652
rect 12921 5628 13539 5652
rect 13701 5628 13899 5652
rect 16461 5628 16776 5652
rect 16881 5628 17139 5652
rect 17601 5628 17919 5652
rect 1041 5568 1212 5592
rect 5181 5568 5316 5592
rect 5421 5568 6279 5592
rect 6681 5568 6999 5592
rect 7401 5568 7659 5592
rect 8541 5568 9099 5592
rect 9921 5568 10719 5592
rect 11481 5568 11919 5592
rect 12201 5568 12819 5592
rect 13281 5568 13419 5592
rect 13881 5568 15519 5592
rect 16401 5568 17199 5592
rect 381 5508 819 5532
rect 861 5508 1299 5532
rect 1341 5508 2139 5532
rect 6381 5508 6579 5532
rect 6621 5508 7119 5532
rect 7161 5508 8139 5532
rect 8781 5508 9039 5532
rect 11181 5508 12159 5532
rect 14361 5508 15219 5532
rect 15621 5508 16119 5532
rect 16941 5508 17079 5532
rect 17781 5508 17859 5532
rect 2601 5448 3219 5472
rect 3261 5448 3759 5472
rect 3801 5448 4659 5472
rect 4821 5448 4959 5472
rect 5121 5448 5439 5472
rect 5841 5448 5979 5472
rect 6021 5448 7176 5472
rect 7281 5448 8259 5472
rect 10221 5448 12939 5472
rect 12981 5448 13419 5472
rect 13461 5448 13899 5472
rect 14661 5448 14919 5472
rect 15081 5448 15312 5472
rect 15288 5421 15312 5448
rect 17721 5448 17919 5472
rect 201 5388 699 5412
rect 2181 5388 2739 5412
rect 2781 5388 2859 5412
rect 4221 5388 4719 5412
rect 4761 5388 5019 5412
rect 7521 5388 7899 5412
rect 8121 5388 8379 5412
rect 8421 5388 9219 5412
rect 9261 5388 9999 5412
rect 11001 5388 11379 5412
rect 12021 5388 12219 5412
rect 15288 5388 15339 5421
rect 15300 5379 15339 5388
rect 15981 5388 16899 5412
rect 801 5328 1212 5352
rect 1188 5292 1212 5328
rect 3501 5328 3639 5352
rect 4401 5328 4479 5352
rect 6381 5328 6519 5352
rect 6981 5328 7239 5352
rect 8181 5328 8559 5352
rect 8601 5328 8979 5352
rect 9381 5328 9759 5352
rect 10881 5328 11559 5352
rect 11601 5328 12399 5352
rect 13101 5328 13239 5352
rect 14121 5328 14919 5352
rect 15660 5352 15699 5361
rect 15648 5319 15699 5352
rect 16521 5328 16839 5352
rect 981 5268 1152 5292
rect 1188 5268 1332 5292
rect 201 5208 339 5232
rect 501 5208 639 5232
rect 681 5208 879 5232
rect 1128 5232 1152 5268
rect 1128 5208 1272 5232
rect 441 5085 579 5109
rect 621 5088 819 5112
rect 888 5112 912 5202
rect 888 5088 1119 5112
rect 1248 5118 1272 5208
rect 1308 5061 1332 5268
rect 1521 5268 1659 5292
rect 2421 5268 2619 5292
rect 2661 5268 3999 5292
rect 4041 5268 4299 5292
rect 4881 5268 5079 5292
rect 5121 5268 5499 5292
rect 5901 5268 6039 5292
rect 7221 5268 7899 5292
rect 9321 5268 9492 5292
rect 1728 5121 1752 5202
rect 1941 5232 1980 5241
rect 1941 5199 1992 5232
rect 2061 5211 2259 5235
rect 2481 5208 2799 5232
rect 3588 5208 3879 5232
rect 1401 5085 1479 5109
rect 1728 5088 1779 5121
rect 1740 5079 1779 5088
rect 1968 5118 1992 5199
rect 2241 5088 2619 5112
rect 2661 5085 2919 5109
rect 2988 5112 3012 5202
rect 3588 5121 3612 5208
rect 4368 5208 4479 5232
rect 4368 5181 4392 5208
rect 4680 5232 4719 5241
rect 3708 5148 3999 5172
rect 2988 5088 3279 5112
rect 3708 5118 3732 5148
rect 4341 5148 4392 5181
rect 4668 5199 4719 5232
rect 4941 5208 5052 5232
rect 5268 5220 6039 5232
rect 4341 5139 4380 5148
rect 4668 5118 4692 5199
rect 5028 5118 5052 5208
rect 5259 5208 6039 5220
rect 5259 5178 5301 5208
rect 6321 5211 6399 5235
rect 6528 5208 6639 5232
rect 5841 5085 5979 5109
rect 6168 5112 6192 5202
rect 6528 5172 6552 5208
rect 6708 5208 6879 5232
rect 6708 5172 6732 5208
rect 7668 5172 7692 5202
rect 8001 5208 8079 5232
rect 8121 5208 8799 5232
rect 6468 5148 6552 5172
rect 6588 5148 6732 5172
rect 7488 5148 7692 5172
rect 6168 5088 6339 5112
rect 6468 5118 6492 5148
rect 6588 5118 6612 5148
rect 7488 5121 7512 5148
rect 6981 5085 7119 5109
rect 7461 5088 7512 5121
rect 7461 5079 7500 5088
rect 7641 5085 7836 5109
rect 7941 5088 8019 5112
rect 8241 5088 8439 5112
rect 8721 5085 9279 5109
rect 9468 5112 9492 5268
rect 12621 5268 12879 5292
rect 13821 5292 13860 5301
rect 13821 5259 13872 5292
rect 14001 5292 14040 5301
rect 14001 5259 14052 5292
rect 14181 5268 14259 5292
rect 14301 5268 14559 5292
rect 9801 5208 10179 5232
rect 10320 5232 10359 5241
rect 10308 5199 10359 5232
rect 10521 5211 10599 5235
rect 10641 5208 10719 5232
rect 11541 5211 11679 5235
rect 10308 5172 10332 5199
rect 11808 5172 11832 5202
rect 10248 5160 10332 5172
rect 11748 5160 11832 5172
rect 10239 5148 10332 5160
rect 11739 5148 11832 5160
rect 10239 5121 10281 5148
rect 9468 5088 9852 5112
rect 2301 5028 2379 5052
rect 3081 5028 3399 5052
rect 5181 5028 5439 5052
rect 5481 5028 6219 5052
rect 9828 5052 9852 5088
rect 9921 5088 9999 5112
rect 10041 5085 10119 5109
rect 11739 5121 11781 5148
rect 11928 5121 11952 5199
rect 10461 5085 10539 5109
rect 10821 5085 11559 5109
rect 12108 5061 12132 5202
rect 12168 5118 12192 5259
rect 12228 5208 13059 5232
rect 9828 5028 9999 5052
rect 3408 4992 3432 5019
rect 12228 5052 12252 5208
rect 12441 5085 12519 5109
rect 13548 5112 13572 5202
rect 13848 5121 13872 5259
rect 14028 5121 14052 5259
rect 14388 5208 14499 5232
rect 13548 5088 13776 5112
rect 14388 5118 14412 5208
rect 14859 5172 14901 5199
rect 14748 5160 14901 5172
rect 14748 5148 14892 5160
rect 14748 5112 14772 5148
rect 15168 5121 15192 5199
rect 15648 5121 15672 5319
rect 15981 5268 16179 5292
rect 16221 5268 16701 5292
rect 16659 5244 16701 5268
rect 17448 5292 17472 5439
rect 17181 5268 17472 5292
rect 16488 5208 16539 5232
rect 15759 5172 15801 5199
rect 15759 5160 16152 5172
rect 15768 5148 16161 5160
rect 16119 5121 16161 5148
rect 14541 5088 14772 5112
rect 12141 5028 12252 5052
rect 12321 5028 12699 5052
rect 13281 5028 13479 5052
rect 14841 5028 15099 5052
rect 16308 5052 16332 5199
rect 16488 5061 16512 5208
rect 16701 5211 16779 5235
rect 17568 5178 17592 5439
rect 16968 5112 16992 5142
rect 17628 5148 17859 5172
rect 17628 5112 17652 5148
rect 16848 5088 16992 5112
rect 17028 5100 17652 5112
rect 17019 5088 17652 5100
rect 16101 5028 16332 5052
rect 16461 5028 16512 5061
rect 16461 5019 16500 5028
rect 16848 5052 16872 5088
rect 17019 5061 17061 5088
rect 16761 5028 16872 5052
rect 17055 5040 17061 5061
rect 3408 4968 3819 4992
rect 4161 4968 4839 4992
rect 6861 4968 7479 4992
rect 7728 4968 8019 4992
rect 7728 4941 7752 4968
rect 8061 4968 9459 4992
rect 12501 4968 13059 4992
rect 13581 4968 13959 4992
rect 15501 4968 15879 4992
rect 1161 4908 2079 4932
rect 4581 4908 5259 4932
rect 5781 4908 6699 4932
rect 6921 4908 7719 4932
rect 7881 4908 8439 4932
rect 8841 4908 10659 4932
rect 14961 4908 15219 4932
rect 16641 4908 17079 4932
rect 3228 4848 5199 4872
rect 1221 4788 1779 4812
rect 1821 4788 2979 4812
rect 3228 4812 3252 4848
rect 6501 4848 7572 4872
rect 3141 4788 3252 4812
rect 4281 4788 5859 4812
rect 6321 4788 6939 4812
rect 7548 4812 7572 4848
rect 9261 4848 9699 4872
rect 11781 4848 12999 4872
rect 15861 4848 16419 4872
rect 7548 4788 8739 4812
rect 9801 4788 10959 4812
rect 11001 4788 11439 4812
rect 11481 4788 11559 4812
rect 11601 4788 13119 4812
rect 13161 4788 13659 4812
rect 15468 4788 15699 4812
rect 321 4728 1239 4752
rect 4821 4728 5316 4752
rect 5421 4728 6252 4752
rect 501 4668 999 4692
rect 1461 4668 2499 4692
rect 3021 4668 5559 4692
rect 6228 4692 6252 4728
rect 13101 4728 13959 4752
rect 15468 4752 15492 4788
rect 17148 4761 17172 5019
rect 17928 5001 17952 5199
rect 18021 5148 18132 5172
rect 18108 5061 18132 5148
rect 14001 4728 15492 4752
rect 6228 4668 6879 4692
rect 7041 4668 8919 4692
rect 10281 4668 10839 4692
rect 12921 4668 14499 4692
rect 14541 4668 15519 4692
rect 3981 4608 4479 4632
rect 4848 4608 5739 4632
rect 4848 4581 4872 4608
rect 7008 4632 7032 4659
rect 6501 4608 7032 4632
rect 7281 4608 8619 4632
rect 15621 4608 15819 4632
rect 15981 4608 16299 4632
rect 381 4548 639 4572
rect 681 4548 1299 4572
rect 3261 4548 3519 4572
rect 4701 4548 4836 4572
rect 4941 4548 5379 4572
rect 5601 4548 5799 4572
rect 5841 4548 6396 4572
rect 7248 4572 7272 4599
rect 6501 4548 7272 4572
rect 7341 4548 8592 4572
rect 801 4488 939 4512
rect 4581 4488 4779 4512
rect 6201 4488 6639 4512
rect 6681 4488 6759 4512
rect 8568 4512 8592 4548
rect 9861 4548 10299 4572
rect 11421 4548 12519 4572
rect 14301 4548 14859 4572
rect 14901 4548 15099 4572
rect 15141 4548 15399 4572
rect 17901 4548 18219 4572
rect 8568 4488 9759 4512
rect 10581 4488 11199 4512
rect 12981 4488 13239 4512
rect 14721 4488 14859 4512
rect 14901 4488 16119 4512
rect 16161 4488 16239 4512
rect 2181 4428 2439 4452
rect 2781 4428 3159 4452
rect 3321 4428 3459 4452
rect 3741 4428 3999 4452
rect 4161 4428 4299 4452
rect 4461 4428 7299 4452
rect 9888 4428 10899 4452
rect 9888 4401 9912 4428
rect 12621 4428 12819 4452
rect 13941 4428 14079 4452
rect 15381 4428 15579 4452
rect 16401 4428 16872 4452
rect 1701 4368 1959 4392
rect 2121 4368 2619 4392
rect 2661 4368 2859 4392
rect 2901 4368 4092 4392
rect 1341 4308 1539 4332
rect 1581 4311 1899 4335
rect 3621 4311 3819 4335
rect 4068 4332 4092 4368
rect 4521 4368 5556 4392
rect 5661 4368 5679 4392
rect 5721 4368 6459 4392
rect 6768 4368 7416 4392
rect 4068 4308 5139 4332
rect 5781 4311 6039 4335
rect 6768 4332 6792 4368
rect 7521 4368 7719 4392
rect 7761 4368 7899 4392
rect 8541 4368 8919 4392
rect 8961 4368 9219 4392
rect 9621 4368 9879 4392
rect 13041 4368 13179 4392
rect 13221 4368 13719 4392
rect 14781 4368 14919 4392
rect 15201 4392 15240 4401
rect 15201 4359 15252 4392
rect 16521 4368 16779 4392
rect 6561 4308 6792 4332
rect 6861 4308 7092 4332
rect 3288 4221 3312 4299
rect 5379 4272 5421 4299
rect 5328 4260 5421 4272
rect 5328 4248 5412 4260
rect 741 4185 999 4209
rect 2541 4185 2619 4209
rect 4341 4185 4539 4209
rect 4881 4188 5019 4212
rect 5328 4212 5352 4248
rect 5241 4188 5352 4212
rect 5481 4188 5799 4212
rect 6141 4185 6279 4209
rect 2121 4128 2859 4152
rect 3201 4128 3459 4152
rect 3501 4128 3759 4152
rect 4041 4128 4359 4152
rect 4701 4119 4719 4161
rect 5601 4128 5739 4152
rect 6528 4152 6552 4302
rect 7068 4272 7092 4308
rect 7161 4308 7419 4332
rect 7461 4308 7539 4332
rect 7668 4308 8019 4332
rect 7068 4248 7272 4272
rect 6681 4188 6759 4212
rect 7248 4161 7272 4248
rect 7668 4212 7692 4308
rect 8301 4311 8379 4335
rect 8868 4308 9099 4332
rect 8868 4272 8892 4308
rect 9381 4311 9456 4335
rect 9801 4311 9936 4335
rect 10041 4332 10080 4341
rect 10041 4299 10092 4332
rect 10239 4332 10281 4359
rect 10161 4320 10281 4332
rect 10161 4308 10272 4320
rect 10461 4311 10659 4335
rect 11121 4311 11319 4335
rect 11481 4308 11799 4332
rect 9519 4272 9561 4299
rect 10068 4272 10092 4299
rect 8808 4248 8892 4272
rect 8928 4248 9492 4272
rect 9519 4260 9612 4272
rect 9528 4248 9612 4260
rect 10068 4260 10512 4272
rect 10068 4248 10521 4260
rect 7641 4188 7692 4212
rect 8808 4212 8832 4248
rect 8661 4188 8832 4212
rect 8928 4212 8952 4248
rect 9468 4221 9492 4248
rect 9588 4221 9612 4248
rect 10479 4221 10521 4248
rect 8901 4188 8952 4212
rect 9021 4188 9159 4212
rect 9468 4188 9519 4221
rect 9480 4179 9519 4188
rect 9588 4188 9636 4221
rect 9600 4179 9636 4188
rect 9741 4185 9816 4209
rect 9921 4188 10059 4212
rect 10221 4188 10299 4212
rect 10881 4188 11139 4212
rect 6528 4128 6639 4152
rect 8301 4128 8379 4152
rect 8979 4152 9021 4176
rect 8721 4128 9021 4152
rect 10488 4152 10512 4179
rect 11868 4212 11892 4359
rect 11961 4308 12219 4332
rect 12441 4308 12759 4332
rect 11781 4188 11892 4212
rect 12141 4185 12279 4209
rect 13341 4188 13419 4212
rect 10488 4128 11319 4152
rect 13608 4152 13632 4302
rect 14361 4308 14559 4332
rect 13788 4212 13812 4299
rect 14808 4221 14832 4299
rect 15228 4221 15252 4359
rect 15561 4308 15696 4332
rect 13701 4188 13812 4212
rect 13941 4185 14019 4209
rect 14421 4188 14619 4212
rect 15768 4212 15792 4299
rect 15381 4188 15792 4212
rect 16068 4212 16092 4299
rect 16188 4272 16212 4359
rect 16281 4308 16392 4332
rect 16368 4272 16392 4308
rect 16188 4248 16332 4272
rect 16368 4248 16419 4272
rect 16068 4188 16179 4212
rect 16308 4212 16332 4248
rect 16641 4245 16719 4269
rect 16308 4188 16479 4212
rect 13521 4128 13632 4152
rect 14901 4128 15039 4152
rect 16641 4128 16779 4152
rect 441 4068 939 4092
rect 981 4068 2019 4092
rect 2181 4068 2379 4092
rect 2421 4068 2799 4092
rect 2841 4068 5439 4092
rect 6021 4068 6339 4092
rect 6501 4068 6819 4092
rect 6981 4068 7539 4092
rect 7881 4068 8199 4092
rect 9321 4068 9399 4092
rect 9981 4068 10419 4092
rect 10761 4068 10899 4092
rect 10941 4068 11019 4092
rect 11421 4068 11559 4092
rect 11901 4068 12819 4092
rect 12861 4068 13179 4092
rect 13881 4068 14712 4092
rect 981 4008 1419 4032
rect 1461 4008 2019 4032
rect 3081 4008 3339 4032
rect 8301 4008 8439 4032
rect 8601 4008 8859 4032
rect 8901 4008 9459 4032
rect 9501 4008 9579 4032
rect 9621 4008 11619 4032
rect 14061 4008 14379 4032
rect 14688 4032 14712 4068
rect 14781 4068 15159 4092
rect 15201 4068 15879 4092
rect 15921 4068 16419 4092
rect 16848 4092 16872 4428
rect 17148 4272 17172 4539
rect 17841 4428 18159 4452
rect 17748 4308 18039 4332
rect 17148 4248 17199 4272
rect 17748 4272 17772 4308
rect 17601 4248 17772 4272
rect 18141 4188 18633 4212
rect 16701 4068 16872 4092
rect 14688 4008 14859 4032
rect 17901 4008 18039 4032
rect 381 3948 1059 3972
rect 3261 3948 3759 3972
rect 5481 3948 5919 3972
rect 6381 3948 8019 3972
rect 8061 3948 11739 3972
rect 16761 3948 17019 3972
rect 17181 3948 17919 3972
rect 1521 3888 2559 3912
rect 2601 3888 3099 3912
rect 4101 3888 4659 3912
rect 4701 3888 5319 3912
rect 6501 3888 6939 3912
rect 8001 3888 8259 3912
rect 8421 3888 9279 3912
rect 9321 3888 10032 3912
rect 10008 3861 10032 3888
rect 10641 3888 10839 3912
rect 14181 3888 14439 3912
rect 16641 3888 17079 3912
rect 17601 3888 17892 3912
rect 1641 3828 2139 3852
rect 2181 3828 2259 3852
rect 3321 3828 3399 3852
rect 3441 3828 3579 3852
rect 7428 3828 8319 3852
rect 7428 3801 7452 3828
rect 10041 3828 10359 3852
rect 12561 3828 12999 3852
rect 16461 3828 16659 3852
rect 17868 3852 17892 3888
rect 17868 3828 18279 3852
rect 621 3768 819 3792
rect 1941 3768 2439 3792
rect 2481 3768 2919 3792
rect 3921 3768 3999 3792
rect 4581 3768 5559 3792
rect 6501 3768 7419 3792
rect 8601 3768 9099 3792
rect 9141 3768 9699 3792
rect 10761 3768 11679 3792
rect 11721 3768 11859 3792
rect 12081 3768 12339 3792
rect 15501 3768 16239 3792
rect 1701 3708 1959 3732
rect 4881 3708 5079 3732
rect 6201 3708 6339 3732
rect 6678 3699 6681 3720
rect 6741 3708 6999 3732
rect 7581 3708 8139 3732
rect 9468 3708 9639 3732
rect 288 3558 312 3699
rect 501 3648 759 3672
rect 801 3648 999 3672
rect 1068 3648 1119 3672
rect 1068 3612 1092 3648
rect 708 3588 1092 3612
rect 708 3558 732 3588
rect -72 3528 99 3552
rect 441 3525 579 3549
rect 1248 3552 1272 3642
rect 2241 3648 2319 3672
rect 2520 3672 2559 3681
rect 2508 3639 2559 3672
rect 1248 3528 1419 3552
rect 2508 3558 2532 3639
rect 2748 3612 2772 3642
rect 3141 3648 3279 3672
rect 3408 3648 3879 3672
rect 3408 3612 3432 3648
rect 3948 3648 4299 3672
rect 2748 3588 2892 3612
rect 3228 3600 3432 3612
rect 1581 3528 1839 3552
rect 2001 3525 2139 3549
rect 2181 3528 2379 3552
rect 2868 3552 2892 3588
rect 3219 3588 3432 3600
rect 3219 3561 3261 3588
rect 3948 3561 3972 3648
rect 5241 3648 5379 3672
rect 5601 3648 5739 3672
rect 6081 3672 6120 3681
rect 6081 3639 6132 3672
rect 6558 3639 6561 3660
rect 6639 3672 6681 3699
rect 6621 3660 6681 3672
rect 6621 3648 6669 3660
rect 6921 3648 7119 3672
rect 4428 3600 4839 3612
rect 4419 3588 4839 3600
rect 4419 3561 4461 3588
rect 6108 3561 6132 3639
rect 6519 3612 6561 3639
rect 6519 3600 6672 3612
rect 6528 3588 6672 3600
rect 2868 3528 2979 3552
rect 4161 3525 4239 3549
rect 5421 3525 5499 3549
rect 6648 3558 6672 3588
rect 7188 3558 7212 3699
rect 7308 3648 7659 3672
rect 7308 3558 7332 3648
rect 7941 3648 8199 3672
rect 8781 3651 9219 3675
rect 8448 3561 8472 3642
rect 6381 3525 6459 3549
rect 6801 3525 6879 3549
rect 8421 3528 8472 3561
rect 9288 3558 9312 3699
rect 9381 3648 9432 3672
rect 9408 3561 9432 3648
rect 9468 3612 9492 3708
rect 10281 3708 10479 3732
rect 10521 3708 10599 3732
rect 12741 3708 13539 3732
rect 10101 3648 10179 3672
rect 9468 3588 9552 3612
rect 8421 3519 8460 3528
rect 8661 3525 8739 3549
rect 8781 3528 8919 3552
rect 9528 3501 9552 3588
rect 9588 3552 9612 3639
rect 9768 3588 9999 3612
rect 9768 3558 9792 3588
rect 10419 3612 10461 3639
rect 11208 3648 11439 3672
rect 10419 3600 10572 3612
rect 10428 3588 10572 3600
rect 9588 3528 9639 3552
rect 10281 3525 10479 3549
rect 10548 3552 10572 3588
rect 10548 3528 10659 3552
rect 10821 3525 10899 3549
rect 11208 3552 11232 3648
rect 11601 3648 11832 3672
rect 11808 3558 11832 3648
rect 12021 3648 12159 3672
rect 12501 3648 12639 3672
rect 12861 3648 13212 3672
rect 13188 3558 13212 3648
rect 13308 3558 13332 3708
rect 14061 3648 14139 3672
rect 14181 3657 14319 3681
rect 15201 3648 15936 3672
rect 16041 3648 16119 3672
rect 16581 3651 16659 3675
rect 17121 3648 17232 3672
rect 11121 3528 11232 3552
rect 11961 3525 12099 3549
rect 13488 3552 13512 3639
rect 14448 3561 14472 3639
rect 16359 3612 16401 3639
rect 16359 3600 16839 3612
rect 16368 3588 16839 3600
rect 17061 3591 17139 3615
rect 17208 3612 17232 3648
rect 17808 3648 17979 3672
rect 17208 3588 17619 3612
rect 13488 3528 13599 3552
rect 2841 3468 3039 3492
rect 3201 3468 3459 3492
rect 4101 3468 4359 3492
rect 6261 3468 6939 3492
rect 6981 3468 7599 3492
rect 7761 3468 8259 3492
rect 8541 3468 9039 3492
rect 9528 3468 9579 3501
rect 9540 3459 9579 3468
rect 11241 3468 11499 3492
rect 11799 3492 11841 3516
rect 14721 3528 15039 3552
rect 15441 3528 16119 3552
rect 16341 3528 16419 3552
rect 16848 3552 16872 3582
rect 16641 3528 16872 3552
rect 11799 3468 12399 3492
rect 14901 3468 15759 3492
rect 15963 3468 16539 3492
rect 17160 3492 17199 3501
rect 17148 3480 17199 3492
rect 17139 3459 17199 3480
rect 17139 3441 17181 3459
rect 1221 3408 1659 3432
rect 2001 3408 2619 3432
rect 10401 3408 11079 3432
rect 11901 3408 12279 3432
rect 12621 3408 13299 3432
rect 14421 3408 15819 3432
rect 3861 3348 4419 3372
rect 13041 3348 13356 3372
rect 13461 3348 14016 3372
rect 14121 3348 15879 3372
rect 16101 3348 16539 3372
rect 141 3288 2559 3312
rect 4281 3288 4539 3312
rect 5601 3288 6999 3312
rect 7161 3288 13899 3312
rect 15288 3288 16779 3312
rect 1341 3228 2499 3252
rect 3381 3228 3819 3252
rect 4881 3228 5739 3252
rect 6141 3228 6999 3252
rect 11901 3228 12879 3252
rect 13101 3228 14079 3252
rect 15288 3252 15312 3288
rect 17808 3261 17832 3648
rect 18201 3648 18372 3672
rect 18081 3588 18312 3612
rect 17928 3432 17952 3579
rect 18288 3501 18312 3588
rect 17928 3408 18027 3432
rect 18348 3432 18372 3648
rect 18069 3408 18072 3432
rect 18348 3408 18492 3432
rect 18201 3348 18399 3372
rect 18468 3261 18492 3408
rect 14301 3228 15312 3252
rect 15381 3228 15459 3252
rect 15501 3228 17559 3252
rect 18441 3228 18492 3261
rect 18441 3219 18480 3228
rect 321 3168 1179 3192
rect 2601 3168 7119 3192
rect 7581 3168 7899 3192
rect 7941 3168 8019 3192
rect 13041 3168 13659 3192
rect 14901 3168 14979 3192
rect 2961 3108 3999 3132
rect 5781 3108 6279 3132
rect 7101 3108 8679 3132
rect 9501 3108 10779 3132
rect 10821 3108 11259 3132
rect 13821 3108 15639 3132
rect 15681 3108 16359 3132
rect 16521 3108 18099 3132
rect 141 3048 1239 3072
rect 4941 3048 5079 3072
rect 6528 3048 7359 3072
rect 201 2988 459 3012
rect 501 2988 939 3012
rect 3021 2988 3159 3012
rect 3201 2988 3579 3012
rect 5181 2988 6219 3012
rect 6528 3012 6552 3048
rect 7608 3048 8379 3072
rect 6261 2988 6552 3012
rect 7608 3012 7632 3048
rect 12921 3048 13479 3072
rect 6621 2988 7632 3012
rect 9441 2988 10659 3012
rect 10701 2988 11019 3012
rect 13881 2988 14499 3012
rect 14901 2988 15252 3012
rect 3261 2928 3699 2952
rect 4161 2928 4719 2952
rect 5268 2928 5679 2952
rect 5268 2901 5292 2928
rect 6501 2928 7659 2952
rect 8121 2928 8499 2952
rect 8541 2928 9159 2952
rect 9201 2928 11499 2952
rect 12681 2928 13119 2952
rect 14361 2928 14799 2952
rect 15228 2952 15252 2988
rect 15321 2988 16179 3012
rect 16341 2988 16479 3012
rect 17181 2988 17439 3012
rect 17601 2988 17979 3012
rect 15228 2928 15459 2952
rect 801 2868 2319 2892
rect 3921 2868 3999 2892
rect 4941 2868 5259 2892
rect 6021 2868 6399 2892
rect 6561 2868 7359 2892
rect 7401 2868 7599 2892
rect 8721 2868 8979 2892
rect 9381 2868 12099 2892
rect 12801 2868 12999 2892
rect 14061 2868 14139 2892
rect 14901 2868 15579 2892
rect 15921 2868 15999 2892
rect 17181 2868 17559 2892
rect 261 2808 639 2832
rect 1221 2808 1899 2832
rect 2601 2808 3099 2832
rect 3141 2808 3279 2832
rect 3321 2808 3459 2832
rect 4761 2808 4959 2832
rect 5001 2808 5799 2832
rect 9801 2808 10059 2832
rect 11001 2808 11139 2832
rect 11568 2808 12459 2832
rect 540 2772 579 2781
rect 528 2739 579 2772
rect 2721 2748 3039 2772
rect 4041 2751 4119 2775
rect 4641 2748 4899 2772
rect 5181 2751 5259 2775
rect 6141 2751 6699 2775
rect 528 2661 552 2739
rect 1128 2661 1152 2742
rect 741 2625 939 2649
rect 1101 2628 1152 2661
rect 1101 2619 1140 2628
rect 1461 2625 1599 2649
rect 2088 2652 2112 2742
rect 7221 2748 7299 2772
rect 7701 2748 7992 2772
rect 1761 2628 2112 2652
rect 2361 2628 2499 2652
rect 2841 2625 3399 2649
rect 3741 2625 3939 2649
rect 4581 2625 4719 2649
rect 5001 2628 5079 2652
rect 5121 2625 5199 2649
rect 5541 2625 5739 2649
rect 5901 2625 5979 2649
rect 6321 2625 6459 2649
rect 6888 2652 6912 2739
rect 6888 2628 7119 2652
rect 7968 2658 7992 2748
rect 8901 2748 9339 2772
rect 9981 2751 10179 2775
rect 11088 2748 11259 2772
rect 10728 2688 10899 2712
rect 10728 2658 10752 2688
rect 11088 2658 11112 2748
rect 11568 2658 11592 2808
rect 14961 2808 15156 2832
rect 15261 2808 15336 2832
rect 16101 2808 16659 2832
rect 11661 2748 11979 2772
rect 12201 2751 12339 2775
rect 12621 2748 12879 2772
rect 13161 2772 13200 2781
rect 13161 2739 13212 2772
rect 13521 2748 13632 2772
rect 7401 2628 7599 2652
rect 8301 2625 8799 2649
rect 9201 2625 9279 2649
rect 9561 2625 9819 2649
rect 10041 2625 10119 2649
rect 10401 2625 10599 2649
rect 11721 2628 11859 2652
rect 12081 2625 12156 2649
rect 12321 2628 12579 2652
rect 12861 2628 12999 2652
rect 13188 2658 13212 2739
rect 13608 2658 13632 2748
rect 13941 2751 14019 2775
rect 15021 2748 15099 2772
rect 13761 2628 13899 2652
rect 14121 2628 14259 2652
rect 14628 2652 14652 2742
rect 15399 2772 15441 2799
rect 15261 2760 15441 2772
rect 15261 2748 15432 2760
rect 15888 2712 15912 2742
rect 16041 2748 17079 2772
rect 18021 2748 18552 2772
rect 15888 2688 16419 2712
rect 14628 2628 14919 2652
rect 15141 2625 15519 2649
rect 15681 2625 15819 2649
rect 16101 2628 16239 2652
rect 201 2568 399 2592
rect 2901 2568 3099 2592
rect 5199 2592 5241 2616
rect 5199 2568 6159 2592
rect 7821 2568 7899 2592
rect 12168 2592 12192 2616
rect 12168 2568 12699 2592
rect 15519 2592 15561 2616
rect 15519 2568 16359 2592
rect 16401 2568 16839 2592
rect 16881 2568 17199 2592
rect 1341 2508 1839 2532
rect 2481 2508 2619 2532
rect 2661 2508 4179 2532
rect 9441 2508 10539 2532
rect 13941 2508 14319 2532
rect 14481 2508 15099 2532
rect 5241 2448 5859 2472
rect 6801 2448 7419 2472
rect 8961 2448 10659 2472
rect 10821 2448 11199 2472
rect 12201 2448 13839 2472
rect 3321 2388 3459 2412
rect 4581 2388 6219 2412
rect 6261 2388 6459 2412
rect 6501 2388 7179 2412
rect 8001 2388 9399 2412
rect 13401 2388 14199 2412
rect 15321 2388 15699 2412
rect 16581 2388 17739 2412
rect 861 2328 1059 2352
rect 1101 2328 1719 2352
rect 2421 2328 2799 2352
rect 5001 2328 5319 2352
rect 5481 2328 5796 2352
rect 5901 2328 6579 2352
rect 9561 2328 9699 2352
rect 9741 2328 10899 2352
rect 11421 2328 12279 2352
rect 12981 2328 13719 2352
rect 14481 2328 15819 2352
rect 201 2268 1179 2292
rect 1221 2268 1599 2292
rect 1641 2268 2139 2292
rect 5781 2268 7119 2292
rect 7161 2268 7659 2292
rect 7701 2268 8079 2292
rect 12081 2268 12759 2292
rect 16941 2268 17139 2292
rect 381 2208 579 2232
rect 1701 2208 1839 2232
rect 2301 2208 2496 2232
rect 2601 2208 3279 2232
rect 3561 2208 3699 2232
rect 3921 2208 5439 2232
rect 6021 2208 6579 2232
rect 6621 2208 6759 2232
rect 6921 2208 7059 2232
rect 7341 2208 8079 2232
rect 9081 2208 9639 2232
rect 9801 2208 10059 2232
rect 10101 2208 10239 2232
rect 10701 2208 10839 2232
rect 11601 2208 12219 2232
rect 12261 2208 12399 2232
rect 13461 2208 13719 2232
rect 15261 2208 15399 2232
rect 15861 2208 16656 2232
rect 16761 2208 16839 2232
rect 141 2148 279 2172
rect 5541 2148 6639 2172
rect 6681 2148 7239 2172
rect 7281 2148 7392 2172
rect 561 2091 1179 2115
rect 1341 2088 1479 2112
rect 1641 2112 1680 2121
rect 1641 2079 1692 2112
rect 1941 2088 2019 2112
rect 2208 2088 2439 2112
rect 1668 1998 1692 2079
rect 2208 1998 2232 2088
rect 2628 2088 2679 2112
rect 2628 2001 2652 2088
rect 2841 2091 2979 2115
rect 201 1965 279 1989
rect 981 1965 1059 1989
rect 3168 1992 3192 2082
rect 3441 2088 3579 2112
rect 3819 2112 3861 2139
rect 3741 2100 3861 2112
rect 3741 2088 3852 2100
rect 3888 2088 4059 2112
rect 3888 2052 3912 2088
rect 4221 2088 4272 2112
rect 3768 2028 3912 2052
rect 3768 1998 3792 2028
rect 4248 2001 4272 2088
rect 4461 2088 4659 2112
rect 2781 1968 3192 1992
rect 3921 1965 4119 1989
rect 4968 1992 4992 2082
rect 5301 2088 5379 2112
rect 5781 2112 5820 2121
rect 5781 2079 5832 2112
rect 6201 2088 6339 2112
rect 4761 1968 4992 1992
rect 5061 1968 5199 1992
rect 5808 1998 5832 2079
rect 5361 1968 5559 1992
rect 6681 1965 6819 1989
rect 7128 1992 7152 2079
rect 7368 1998 7392 2148
rect 8181 2148 8979 2172
rect 11061 2148 11199 2172
rect 12921 2148 13059 2172
rect 14121 2148 14319 2172
rect 14961 2148 15279 2172
rect 16428 2148 16959 2172
rect 7821 2088 8919 2112
rect 7419 2052 7461 2079
rect 7419 2040 7632 2052
rect 7428 2028 7632 2040
rect 7608 1998 7632 2028
rect 8088 1998 8112 2088
rect 10221 2088 10299 2112
rect 9288 2052 9312 2082
rect 10188 2052 10212 2082
rect 10881 2088 11052 2112
rect 9288 2028 9792 2052
rect 6981 1968 7152 1992
rect 8481 1968 8559 1992
rect 9021 1965 9099 1989
rect 9621 1965 9699 1989
rect 9768 1992 9792 2028
rect 10128 2028 10212 2052
rect 11028 2052 11052 2088
rect 11301 2088 11439 2112
rect 16428 2124 16452 2148
rect 17001 2148 17259 2172
rect 11028 2028 11112 2052
rect 10128 1992 10152 2028
rect 9768 1968 10152 1992
rect 10641 1968 10779 1992
rect 11088 1998 11112 2028
rect 12588 2052 12612 2085
rect 13221 2088 13359 2112
rect 14520 2112 14556 2121
rect 12381 2028 12612 2052
rect 12708 2040 12972 2052
rect 12699 2028 12972 2040
rect 12699 2001 12741 2028
rect 10821 1968 10959 1992
rect 11241 1965 11499 1989
rect 12021 1965 12219 1989
rect 12948 1998 12972 2028
rect 13488 2001 13512 2082
rect 12981 1965 13239 1989
rect 13461 1968 13512 2001
rect 14508 2079 14556 2112
rect 14661 2091 14799 2115
rect 15141 2088 15819 2112
rect 15981 2091 16179 2115
rect 16341 2091 16419 2115
rect 16608 2088 16839 2112
rect 14508 1998 14532 2079
rect 16608 1998 16632 2088
rect 17028 2088 17919 2112
rect 17028 2001 17052 2088
rect 13461 1959 13500 1968
rect 15381 1968 15759 1992
rect 1008 1908 1239 1932
rect 141 1848 399 1872
rect 1008 1872 1032 1908
rect 1821 1908 2019 1932
rect 3888 1932 3912 1956
rect 3681 1908 3912 1932
rect 4521 1908 5259 1932
rect 6321 1908 6579 1932
rect 10341 1908 10452 1932
rect 441 1848 1032 1872
rect 1101 1848 1359 1872
rect 2361 1848 3459 1872
rect 4461 1848 4899 1872
rect 7281 1848 7479 1872
rect 8781 1848 9819 1872
rect 9861 1848 9999 1872
rect 10428 1872 10452 1908
rect 13581 1908 13959 1932
rect 14481 1908 14619 1932
rect 15201 1908 16119 1932
rect 17361 1908 17979 1932
rect 10428 1848 11619 1872
rect 11661 1848 11739 1872
rect 13401 1848 13839 1872
rect 14961 1848 15639 1872
rect 2781 1788 4479 1812
rect 5961 1788 6399 1812
rect 7248 1812 7272 1839
rect 6441 1788 7272 1812
rect 8961 1788 9399 1812
rect 10161 1788 10359 1812
rect 10401 1788 10479 1812
rect 12321 1788 13779 1812
rect 15801 1788 16719 1812
rect 16761 1788 16959 1812
rect 861 1728 1779 1752
rect 2541 1728 2859 1752
rect 2901 1728 3219 1752
rect 5001 1728 5679 1752
rect 8241 1728 8859 1752
rect 12501 1728 13419 1752
rect 14241 1728 14979 1752
rect 16401 1728 17619 1752
rect 4881 1668 6099 1692
rect 6861 1668 7959 1692
rect 9381 1668 10119 1692
rect 13821 1668 15039 1692
rect 16521 1668 17139 1692
rect 2661 1608 3639 1632
rect 5481 1608 6039 1632
rect 7101 1608 7719 1632
rect 13761 1608 17079 1632
rect 17361 1608 17799 1632
rect 3021 1548 3279 1572
rect 3321 1548 3399 1572
rect 6141 1548 7959 1572
rect 8001 1548 10119 1572
rect 11121 1548 12339 1572
rect 12381 1548 13119 1572
rect 1281 1488 1659 1512
rect 1701 1488 2859 1512
rect 3141 1488 3519 1512
rect 4161 1488 5079 1512
rect 13521 1488 15459 1512
rect 16161 1488 16239 1512
rect 17361 1488 18039 1512
rect 18081 1488 18339 1512
rect 381 1428 759 1452
rect 801 1428 2379 1452
rect 5601 1428 7059 1452
rect 10461 1428 11079 1452
rect 12981 1428 14919 1452
rect 16821 1428 17379 1452
rect 2601 1368 2679 1392
rect 2721 1368 2799 1392
rect 3561 1368 3819 1392
rect 3861 1368 4239 1392
rect 5181 1368 5439 1392
rect 8301 1368 9579 1392
rect 9861 1368 10719 1392
rect 11361 1368 13059 1392
rect 16701 1368 17199 1392
rect 1521 1308 1839 1332
rect 4761 1308 5919 1332
rect 7161 1308 7359 1332
rect 7881 1308 8499 1332
rect 8541 1308 8559 1332
rect 8601 1308 9039 1332
rect 9261 1308 9639 1332
rect 11481 1308 11919 1332
rect 11961 1308 12459 1332
rect 15201 1308 15459 1332
rect 17841 1308 18219 1332
rect 501 1248 639 1272
rect 681 1248 939 1272
rect 3528 1248 4179 1272
rect 468 1188 579 1212
rect 468 1092 492 1188
rect 1308 1188 1539 1212
rect 1308 1098 1332 1188
rect 1941 1191 2079 1215
rect 441 1068 492 1092
rect 1761 1068 1899 1092
rect 2208 1092 2232 1182
rect 3348 1101 3372 1179
rect 3528 1152 3552 1248
rect 7368 1272 7392 1299
rect 7368 1248 9159 1272
rect 9201 1248 9459 1272
rect 9801 1248 9879 1272
rect 10641 1248 10899 1272
rect 10941 1248 11139 1272
rect 13221 1248 14139 1272
rect 16341 1248 16479 1272
rect 16521 1248 16839 1272
rect 17481 1248 17619 1272
rect 3600 1212 3639 1221
rect 3468 1128 3552 1152
rect 3588 1179 3639 1212
rect 3981 1191 4419 1215
rect 4668 1188 4959 1212
rect 2061 1068 2232 1092
rect 2421 1068 2499 1092
rect 2901 1068 3039 1092
rect 3468 1098 3492 1128
rect 3588 1098 3612 1179
rect 4668 1152 4692 1188
rect 5241 1191 5319 1215
rect 5601 1188 5799 1212
rect 6639 1215 6681 1239
rect 6201 1191 6699 1215
rect 6648 1188 6672 1191
rect 7761 1188 8259 1212
rect 9741 1191 10239 1215
rect 11301 1191 11559 1215
rect 11601 1188 11799 1212
rect 4281 1128 4692 1152
rect 5808 1152 5832 1182
rect 7248 1152 7272 1182
rect 12141 1188 12339 1212
rect 12381 1188 12639 1212
rect 12801 1191 12879 1215
rect 13341 1188 13599 1212
rect 14361 1197 14559 1221
rect 5808 1128 8232 1152
rect 3621 1068 3759 1092
rect 5541 1068 5859 1092
rect 5928 1092 5952 1128
rect 5928 1068 6279 1092
rect 6441 1065 6516 1089
rect 6621 1065 6759 1089
rect 6921 1068 7119 1092
rect 7461 1068 7659 1092
rect 7701 1068 7839 1092
rect 8208 1098 8232 1128
rect 8421 1128 8919 1152
rect 8001 1068 8079 1092
rect 8241 1068 8559 1092
rect 9141 1068 9699 1092
rect 10221 1065 10419 1089
rect 10941 1065 11019 1089
rect 12021 1068 12579 1092
rect 12741 1068 12939 1092
rect 15108 1098 15132 1239
rect 15321 1188 15579 1212
rect 17040 1212 17079 1221
rect 17028 1179 17079 1212
rect 17961 1191 18279 1215
rect 15768 1128 16779 1152
rect 13701 1068 13779 1092
rect 2001 1008 2139 1032
rect 4221 1008 5199 1032
rect 5859 1032 5901 1056
rect 15768 1092 15792 1128
rect 17028 1092 17052 1179
rect 17361 1065 17619 1089
rect 17781 1065 18099 1089
rect 5859 1008 6099 1032
rect 8301 1008 8379 1032
rect 9261 1008 9399 1032
rect 9441 1008 9639 1032
rect 11121 1008 11499 1032
rect 11541 1008 11859 1032
rect 13281 1008 14439 1032
rect 14481 1008 15219 1032
rect 15261 1008 15399 1032
rect 741 948 939 972
rect 1221 948 2019 972
rect 2061 948 2439 972
rect 2841 948 3339 972
rect 3861 948 4119 972
rect 6261 948 8499 972
rect 9561 948 9699 972
rect 9981 948 10059 972
rect 10101 948 10299 972
rect 10341 948 10959 972
rect 11001 948 11259 972
rect 11841 948 12159 972
rect 13161 948 14019 972
rect 17901 948 18039 972
rect 1641 888 1839 912
rect 4521 888 5199 912
rect 5361 888 8139 912
rect 9141 888 9759 912
rect 10581 888 10719 912
rect 17181 888 17319 912
rect 17481 888 18399 912
rect 321 828 399 852
rect 441 828 1479 852
rect 1521 828 1959 852
rect 2781 828 3699 852
rect 4641 828 5139 852
rect 5181 828 5979 852
rect 7821 828 8439 852
rect 8721 828 9699 852
rect 9861 828 10659 852
rect 17961 828 18159 852
rect 1641 768 2199 792
rect 2541 768 2679 792
rect 3021 768 3159 792
rect 3201 768 4419 792
rect 4548 768 6039 792
rect 4548 741 4572 768
rect 6081 768 6339 792
rect 7701 768 9639 792
rect 9801 768 11379 792
rect 11421 768 12279 792
rect 12321 768 13059 792
rect 14781 768 15039 792
rect 15501 768 15579 792
rect 81 708 279 732
rect 861 708 1239 732
rect 3321 708 3519 732
rect 3921 708 4539 732
rect 6801 708 7299 732
rect 7848 708 10239 732
rect 801 648 1779 672
rect 1821 648 2259 672
rect 2301 648 2619 672
rect 2661 648 4899 672
rect 5121 648 5379 672
rect 6021 648 6279 672
rect 6681 648 7239 672
rect 7848 672 7872 708
rect 10281 708 10599 732
rect 7401 648 7872 672
rect 8061 648 10119 672
rect 10701 648 11199 672
rect 11241 648 11499 672
rect 12141 648 12732 672
rect 5001 588 5859 612
rect 5901 588 6519 612
rect 7341 588 7899 612
rect 8760 612 8799 621
rect 8748 588 8799 612
rect 8760 579 8799 588
rect 8841 588 9192 612
rect 348 528 819 552
rect 348 438 372 528
rect 981 528 1119 552
rect 1188 438 1212 579
rect 1281 528 2379 552
rect 2448 438 2472 579
rect 2580 552 2619 561
rect 2568 519 2619 552
rect 3021 528 3252 552
rect 2568 438 2592 519
rect 3228 492 3252 528
rect 3381 528 3459 552
rect 4041 531 4179 555
rect 4341 528 4839 552
rect 5241 528 5559 552
rect 5721 528 5799 552
rect 5868 528 6159 552
rect 5868 492 5892 528
rect 6921 531 7059 555
rect 7461 531 7599 555
rect 8268 528 8679 552
rect 8268 492 8292 528
rect 8961 528 9099 552
rect 2781 468 3192 492
rect 3228 468 3312 492
rect 501 408 699 432
rect 741 408 1059 432
rect 1821 405 1899 429
rect 3168 438 3192 468
rect 2841 408 2919 432
rect 3288 432 3312 468
rect 5628 468 9072 492
rect 5628 438 5652 468
rect 9048 438 9072 468
rect 9168 438 9192 588
rect 9261 528 9399 552
rect 10161 528 10659 552
rect 10920 552 10959 561
rect 9501 468 9732 492
rect 9708 438 9732 468
rect 3288 408 3639 432
rect 4281 405 4419 429
rect 4581 405 4659 429
rect 5181 408 5499 432
rect 5901 405 5979 429
rect 6141 405 6219 429
rect 6381 405 6459 429
rect 6621 405 6759 429
rect 6981 408 7839 432
rect 8061 405 8199 429
rect 8541 405 8619 429
rect 8781 405 8919 429
rect 9441 405 9579 429
rect 10221 408 10539 432
rect 1059 372 1101 396
rect 1059 348 1419 372
rect 1581 348 1677 372
rect 3861 348 4119 372
rect 5619 372 5661 396
rect 5301 348 5661 372
rect 7281 348 7599 372
rect 7641 348 7719 372
rect 7839 372 7881 396
rect 7839 348 8319 372
rect 10641 348 10779 372
rect 10848 372 10872 522
rect 10908 519 10959 552
rect 12399 552 12441 579
rect 12321 540 12441 552
rect 12321 528 12432 540
rect 12501 531 12639 555
rect 10908 438 10932 519
rect 11328 492 11352 522
rect 11121 468 11352 492
rect 12708 438 12732 648
rect 14541 648 14859 672
rect 15681 648 16119 672
rect 12801 528 12939 552
rect 13221 531 13299 555
rect 13701 531 13899 555
rect 14781 528 15039 552
rect 15921 528 16119 552
rect 16581 531 16779 555
rect 14208 468 14592 492
rect 11421 405 12099 429
rect 12261 408 12579 432
rect 13161 408 13479 432
rect 14208 432 14232 468
rect 14568 432 14592 468
rect 14421 399 14496 423
rect 14601 399 15339 423
rect 15561 399 15639 423
rect 17601 405 17799 429
rect 10848 348 11052 372
rect 2721 288 3639 312
rect 3801 288 4779 312
rect 4821 288 4959 312
rect 5841 288 7059 312
rect 7101 288 7359 312
rect 9021 288 9459 312
rect 11028 312 11052 348
rect 12981 348 13239 372
rect 11028 288 11079 312
rect 11121 288 12339 312
rect 12381 288 12459 312
rect 12681 288 13299 312
rect 2241 228 4479 252
rect 5421 228 7032 252
rect 981 168 5139 192
rect 7008 192 7032 228
rect 9621 228 12219 252
rect 7008 168 7239 192
rect 8481 168 12039 192
rect 12921 168 13599 192
rect 2301 108 3999 132
rect 6441 108 8319 132
rect 8601 108 10179 132
rect 10401 108 11259 132
use INVX1  _889_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 16170 0 -1 5490
box -36 -24 216 816
use NOR2X1  _890_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 15210 0 1 3930
box -36 -24 276 816
use NAND2X1  _891_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 15570 0 1 3930
box -36 -24 276 816
use INVX1  _892_
timestamp 1727136778
transform 1 0 16230 0 -1 3930
box -36 -24 216 816
use INVX1  _893_
timestamp 1727136778
transform -1 0 15930 0 1 3930
box -36 -24 216 816
use INVX2  _894_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 16590 0 -1 3930
box -36 -24 216 816
use NOR2X1  _895_
timestamp 1727136778
transform -1 0 15990 0 -1 5490
box -36 -24 276 816
use NAND2X1  _896_
timestamp 1727136778
transform -1 0 15630 0 -1 5490
box -36 -24 276 816
use INVX1  _897_
timestamp 1727136778
transform 1 0 15450 0 1 7050
box -36 -24 216 816
use NOR2X1  _898_
timestamp 1727136778
transform -1 0 16710 0 -1 5490
box -36 -24 276 816
use AOI21X1  _899_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 15870 0 1 5490
box -36 -24 336 816
use NOR2X1  _900_
timestamp 1727136778
transform -1 0 17850 0 1 7050
box -36 -24 276 816
use OAI21X1  _901_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 17430 0 1 7050
box -36 -24 336 816
use INVX1  _902_
timestamp 1727136778
transform 1 0 17490 0 -1 7050
box -36 -24 216 816
use INVX4  _903_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 14790 0 1 5490
box -36 -24 276 816
use OAI21X1  _904_
timestamp 1727136778
transform -1 0 16350 0 1 3930
box -36 -24 336 816
use INVX1  _905_
timestamp 1727136778
transform -1 0 17310 0 -1 7050
box -36 -24 216 816
use NOR2X1  _906_
timestamp 1727136778
transform -1 0 12930 0 -1 7050
box -36 -24 276 816
use INVX1  _907_
timestamp 1727136778
transform 1 0 15030 0 -1 7050
box -36 -24 216 816
use INVX1  _908_
timestamp 1727136778
transform 1 0 17970 0 -1 8610
box -36 -24 216 816
use OAI21X1  _909_
timestamp 1727136778
transform 1 0 16890 0 1 5490
box -36 -24 336 816
use OAI21X1  _910_
timestamp 1727136778
transform 1 0 16650 0 -1 7050
box -36 -24 336 816
use AOI22X1  _911_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 16350 0 1 5490
box -42 -24 396 816
use NAND2X1  _912_
timestamp 1727136778
transform 1 0 17370 0 1 5490
box -36 -24 276 816
use OAI21X1  _913_
timestamp 1727136778
transform -1 0 17010 0 1 7050
box -36 -24 336 816
use OAI21X1  _914_
timestamp 1727136778
transform -1 0 16110 0 1 7050
box -36 -24 336 816
use NAND2X1  _915_
timestamp 1727136778
transform 1 0 15810 0 -1 7050
box -36 -24 276 816
use NOR2X1  _916_
timestamp 1727136778
transform -1 0 17190 0 1 8610
box -36 -24 276 816
use NOR2X1  _917_
timestamp 1727136778
transform 1 0 17550 0 -1 8610
box -36 -24 276 816
use OAI22X1  _918_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 16590 0 -1 8610
box -36 -24 396 816
use OR2X2  _919_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 16290 0 1 7050
box -36 -24 336 816
use INVX1  _920_
timestamp 1727136778
transform -1 0 16890 0 -1 8610
box -36 -24 216 816
use AOI22X1  _921_
timestamp 1727136778
transform 1 0 17070 0 -1 8610
box -42 -24 396 816
use NAND3X1  _922_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 16230 0 -1 7050
box -36 -24 336 816
use AND2X2  _923_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 17790 0 -1 7050
box -36 -24 336 819
use OAI21X1  _924_
timestamp 1727136778
transform 1 0 17790 0 1 5490
box -36 -24 336 816
use INVX1  _925_
timestamp 1727136778
transform -1 0 18150 0 1 3930
box -36 -24 216 816
use INVX1  _926_
timestamp 1727136778
transform -1 0 13170 0 1 13290
box -36 -24 216 816
use NAND2X1  _927_
timestamp 1727136778
transform 1 0 14670 0 -1 10170
box -36 -24 276 816
use OAI21X1  _928_
timestamp 1727136778
transform 1 0 14190 0 -1 10170
box -36 -24 336 816
use INVX1  _929_
timestamp 1727136778
transform 1 0 12690 0 1 13290
box -36 -24 216 816
use NAND2X1  _930_
timestamp 1727136778
transform 1 0 11130 0 1 11730
box -36 -24 276 816
use OAI21X1  _931_
timestamp 1727136778
transform -1 0 11850 0 1 11730
box -36 -24 336 816
use INVX1  _932_
timestamp 1727136778
transform 1 0 12450 0 -1 13290
box -36 -24 216 816
use NAND2X1  _933_
timestamp 1727136778
transform -1 0 13530 0 -1 10170
box -36 -24 276 816
use OAI21X1  _934_
timestamp 1727136778
transform 1 0 13710 0 -1 10170
box -36 -24 336 816
use INVX1  _935_
timestamp 1727136778
transform -1 0 16350 0 1 14850
box -36 -24 216 816
use NAND2X1  _936_
timestamp 1727136778
transform 1 0 12330 0 1 13290
box -36 -24 276 816
use OAI21X1  _937_
timestamp 1727136778
transform -1 0 12330 0 -1 13290
box -36 -24 336 816
use INVX1  _938_
timestamp 1727136778
transform -1 0 12150 0 -1 16410
box -36 -24 216 816
use NAND2X1  _939_
timestamp 1727136778
transform 1 0 11070 0 1 13290
box -36 -24 276 816
use OAI21X1  _940_
timestamp 1727136778
transform 1 0 10470 0 -1 13290
box -36 -24 336 816
use INVX1  _941_
timestamp 1727136778
transform -1 0 9990 0 -1 14850
box -36 -24 216 816
use NAND2X1  _942_
timestamp 1727136778
transform 1 0 10950 0 -1 11730
box -36 -24 276 816
use OAI21X1  _943_
timestamp 1727136778
transform 1 0 10530 0 -1 11730
box -36 -24 336 816
use INVX1  _944_
timestamp 1727136778
transform -1 0 16170 0 1 10170
box -36 -24 216 816
use NAND2X1  _945_
timestamp 1727136778
transform 1 0 16770 0 -1 10170
box -36 -24 276 816
use OAI21X1  _946_
timestamp 1727136778
transform 1 0 16350 0 -1 10170
box -36 -24 336 816
use INVX4  _947_
timestamp 1727136778
transform 1 0 17070 0 1 2370
box -36 -24 276 816
use NAND2X1  _948_
timestamp 1727136778
transform 1 0 15810 0 -1 8610
box -36 -24 276 816
use OAI21X1  _949_
timestamp 1727136778
transform 1 0 15390 0 -1 8610
box -36 -24 336 816
use INVX1  _950_
timestamp 1727136778
transform -1 0 14190 0 1 5490
box -36 -24 216 816
use INVX1  _951_
timestamp 1727136778
transform 1 0 11790 0 -1 5490
box -36 -24 216 816
use INVX2  _952_
timestamp 1727136778
transform 1 0 7110 0 1 10170
box -36 -24 216 816
use NOR2X1  _953_
timestamp 1727136778
transform 1 0 8010 0 -1 3930
box -36 -24 276 816
use AND2X2  _954_
timestamp 1727136778
transform -1 0 7770 0 1 3930
box -36 -24 336 819
use NAND2X1  _955_
timestamp 1727136778
transform 1 0 8370 0 1 2370
box -36 -24 276 816
use NAND2X1  _956_
timestamp 1727136778
transform 1 0 9630 0 1 5490
box -36 -24 276 816
use NAND2X1  _957_
timestamp 1727136778
transform 1 0 10530 0 -1 5490
box -36 -24 276 816
use OR2X2  _958_
timestamp 1727136778
transform 1 0 10950 0 -1 5490
box -36 -24 336 816
use NAND2X1  _959_
timestamp 1727136778
transform 1 0 10950 0 1 3930
box -36 -24 276 816
use AND2X2  _960_
timestamp 1727136778
transform 1 0 9570 0 1 3930
box -36 -24 336 819
use OAI21X1  _961_
timestamp 1727136778
transform -1 0 10770 0 1 3930
box -36 -24 336 816
use NAND2X1  _962_
timestamp 1727136778
transform 1 0 11430 0 -1 5490
box -36 -24 276 816
use INVX1  _963_
timestamp 1727136778
transform 1 0 8850 0 -1 3930
box -36 -24 216 816
use NAND2X1  _964_
timestamp 1727136778
transform -1 0 8190 0 1 5490
box -36 -24 276 816
use NAND2X1  _965_
timestamp 1727136778
transform 1 0 7590 0 1 5490
box -36 -24 276 816
use OR2X2  _966_
timestamp 1727136778
transform 1 0 10110 0 -1 5490
box -36 -24 336 816
use INVX1  _967_
timestamp 1727136778
transform -1 0 8970 0 1 5490
box -36 -24 216 816
use INVX1  _968_
timestamp 1727136778
transform 1 0 7830 0 1 10170
box -36 -24 216 816
use OAI21X1  _969_
timestamp 1727136778
transform -1 0 8670 0 1 5490
box -36 -24 336 816
use NAND3X1  _970_
timestamp 1727136778
transform 1 0 9150 0 -1 3930
box -36 -24 336 816
use NOR2X1  _971_
timestamp 1727136778
transform 1 0 9210 0 -1 5490
box -36 -24 276 816
use AND2X2  _972_
timestamp 1727136778
transform -1 0 9930 0 -1 5490
box -36 -24 336 819
use OAI21X1  _973_
timestamp 1727136778
transform 1 0 9150 0 1 3930
box -36 -24 336 816
use NAND3X1  _974_
timestamp 1727136778
transform -1 0 10830 0 1 2370
box -36 -24 336 816
use INVX1  _975_
timestamp 1727136778
transform 1 0 9270 0 1 2370
box -36 -24 216 816
use NAND2X1  _976_
timestamp 1727136778
transform 1 0 7890 0 1 3930
box -36 -24 276 816
use INVX2  _977_
timestamp 1727136778
transform 1 0 6450 0 1 11730
box -36 -24 216 816
use NAND2X1  _978_
timestamp 1727136778
transform 1 0 7590 0 -1 5490
box -36 -24 276 816
use OAI21X1  _979_
timestamp 1727136778
transform 1 0 6330 0 1 3930
box -36 -24 336 816
use OAI21X1  _980_
timestamp 1727136778
transform 1 0 8790 0 1 2370
box -36 -24 336 816
use AOI21X1  _981_
timestamp 1727136778
transform 1 0 11010 0 1 2370
box -36 -24 336 816
use OAI21X1  _982_
timestamp 1727136778
transform -1 0 10710 0 -1 2370
box -36 -24 336 816
use OAI21X1  _983_
timestamp 1727136778
transform -1 0 8610 0 1 3930
box -36 -24 336 816
use AND2X2  _984_
timestamp 1727136778
transform -1 0 7650 0 -1 7050
box -36 -24 336 819
use NAND3X1  _985_
timestamp 1727136778
transform -1 0 7410 0 1 5490
box -36 -24 336 816
use AOI22X1  _986_
timestamp 1727136778
transform -1 0 5550 0 -1 7050
box -42 -24 396 816
use INVX1  _987_
timestamp 1727136778
transform -1 0 5010 0 1 2370
box -36 -24 216 816
use NAND2X1  _988_
timestamp 1727136778
transform -1 0 4410 0 1 3930
box -36 -24 276 816
use INVX1  _989_
timestamp 1727136778
transform -1 0 5610 0 -1 3930
box -36 -24 216 816
use NAND3X1  _990_
timestamp 1727136778
transform 1 0 5670 0 1 2370
box -36 -24 336 816
use NAND2X1  _991_
timestamp 1727136778
transform 1 0 7290 0 1 11730
box -36 -24 276 816
use NOR2X1  _992_
timestamp 1727136778
transform -1 0 7410 0 -1 5490
box -36 -24 276 816
use OAI21X1  _993_
timestamp 1727136778
transform 1 0 6150 0 1 2370
box -36 -24 336 816
use NAND3X1  _994_
timestamp 1727136778
transform 1 0 7890 0 1 2370
box -36 -24 336 816
use AOI21X1  _995_
timestamp 1727136778
transform -1 0 8670 0 -1 3930
box -36 -24 336 816
use OAI21X1  _996_
timestamp 1727136778
transform 1 0 5190 0 1 2370
box -36 -24 336 816
use NAND3X1  _997_
timestamp 1727136778
transform -1 0 4650 0 1 2370
box -36 -24 336 816
use NAND3X1  _998_
timestamp 1727136778
transform 1 0 4890 0 -1 2370
box -36 -24 336 816
use NAND2X1  _999_
timestamp 1727136778
transform 1 0 6690 0 1 5490
box -36 -24 276 816
use INVX1  _1000_
timestamp 1727136778
transform 1 0 6750 0 1 3930
box -36 -24 216 816
use AND2X2  _1001_
timestamp 1727136778
transform 1 0 8430 0 -1 5490
box -36 -24 336 819
use NAND2X1  _1002_
timestamp 1727136778
transform 1 0 7110 0 1 3930
box -36 -24 276 816
use INVX1  _1003_
timestamp 1727136778
transform -1 0 9030 0 -1 5490
box -36 -24 216 816
use OAI21X1  _1004_
timestamp 1727136778
transform 1 0 7530 0 -1 3930
box -36 -24 336 816
use NAND3X1  _1005_
timestamp 1727136778
transform -1 0 7350 0 -1 3930
box -36 -24 336 816
use OAI21X1  _1006_
timestamp 1727136778
transform 1 0 6150 0 -1 3930
box -36 -24 336 816
use INVX1  _1007_
timestamp 1727136778
transform -1 0 5250 0 1 3930
box -36 -24 216 816
use OAI21X1  _1008_
timestamp 1727136778
transform 1 0 5430 0 1 3930
box -36 -24 336 816
use NAND3X1  _1009_
timestamp 1727136778
transform -1 0 6210 0 1 3930
box -36 -24 336 816
use AND2X2  _1010_
timestamp 1727136778
transform 1 0 6990 0 1 2370
box -36 -24 336 819
use NAND3X1  _1011_
timestamp 1727136778
transform -1 0 6990 0 -1 2370
box -36 -24 336 816
use AOI21X1  _1012_
timestamp 1727136778
transform -1 0 4770 0 -1 2370
box -36 -24 336 816
use AOI21X1  _1013_
timestamp 1727136778
transform -1 0 7710 0 1 2370
box -36 -24 336 816
use NAND2X1  _1014_
timestamp 1727136778
transform -1 0 6870 0 1 2370
box -36 -24 276 816
use OAI21X1  _1015_
timestamp 1727136778
transform -1 0 6510 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1016_
timestamp 1727136778
transform -1 0 6510 0 1 810
box -36 -24 336 816
use AOI21X1  _1017_
timestamp 1727136778
transform 1 0 6690 0 1 810
box -36 -24 336 816
use OAI21X1  _1018_
timestamp 1727136778
transform -1 0 7470 0 1 810
box -36 -24 336 816
use AOI21X1  _1019_
timestamp 1727136778
transform -1 0 5610 0 -1 2370
box -36 -24 336 816
use OAI21X1  _1020_
timestamp 1727136778
transform -1 0 4890 0 1 3930
box -36 -24 336 816
use AND2X2  _1021_
timestamp 1727136778
transform -1 0 4650 0 1 11730
box -36 -24 336 819
use NAND2X1  _1022_
timestamp 1727136778
transform -1 0 4410 0 1 5490
box -36 -24 276 816
use INVX1  _1023_
timestamp 1727136778
transform 1 0 3510 0 1 7050
box -36 -24 216 816
use INVX2  _1024_
timestamp 1727136778
transform 1 0 4590 0 -1 14850
box -36 -24 216 816
use NAND2X1  _1025_
timestamp 1727136778
transform 1 0 4410 0 -1 7050
box -36 -24 276 816
use OAI21X1  _1026_
timestamp 1727136778
transform 1 0 3870 0 1 7050
box -36 -24 336 816
use NAND2X1  _1027_
timestamp 1727136778
transform 1 0 4590 0 1 5490
box -36 -24 276 816
use INVX1  _1028_
timestamp 1727136778
transform 1 0 3210 0 -1 5490
box -36 -24 216 816
use NAND3X1  _1029_
timestamp 1727136778
transform -1 0 3090 0 -1 5490
box -36 -24 336 816
use NOR2X1  _1030_
timestamp 1727136778
transform -1 0 5070 0 -1 7050
box -36 -24 276 816
use AOI22X1  _1031_
timestamp 1727136778
transform 1 0 3930 0 -1 7050
box -42 -24 396 816
use OAI21X1  _1032_
timestamp 1727136778
transform -1 0 4050 0 1 5490
box -36 -24 336 816
use AOI21X1  _1033_
timestamp 1727136778
transform -1 0 3570 0 1 3930
box -36 -24 336 816
use AOI21X1  _1034_
timestamp 1727136778
transform -1 0 5310 0 -1 3930
box -36 -24 336 816
use OAI21X1  _1035_
timestamp 1727136778
transform -1 0 3570 0 1 5490
box -36 -24 336 816
use NAND3X1  _1036_
timestamp 1727136778
transform -1 0 3870 0 -1 5490
box -36 -24 336 816
use AOI21X1  _1037_
timestamp 1727136778
transform -1 0 3510 0 -1 3930
box -36 -24 336 816
use NAND2X1  _1038_
timestamp 1727136778
transform 1 0 4950 0 1 5490
box -36 -24 276 816
use INVX1  _1039_
timestamp 1727136778
transform -1 0 4230 0 -1 5490
box -36 -24 216 816
use AND2X2  _1040_
timestamp 1727136778
transform -1 0 6510 0 1 5490
box -36 -24 336 819
use AND2X2  _1041_
timestamp 1727136778
transform -1 0 8250 0 -1 5490
box -36 -24 336 819
use NAND2X1  _1042_
timestamp 1727136778
transform 1 0 5790 0 1 5490
box -36 -24 276 816
use INVX2  _1043_
timestamp 1727136778
transform 1 0 6990 0 -1 7050
box -36 -24 216 816
use NAND2X1  _1044_
timestamp 1727136778
transform 1 0 6810 0 -1 5490
box -36 -24 276 816
use OAI21X1  _1045_
timestamp 1727136778
transform 1 0 6390 0 -1 5490
box -36 -24 336 816
use NAND3X1  _1046_
timestamp 1727136778
transform -1 0 5190 0 -1 5490
box -36 -24 336 816
use OAI21X1  _1047_
timestamp 1727136778
transform 1 0 5310 0 1 5490
box -36 -24 336 816
use OAI21X1  _1048_
timestamp 1727136778
transform -1 0 6210 0 -1 5490
box -36 -24 336 816
use NAND3X1  _1049_
timestamp 1727136778
transform -1 0 4710 0 -1 5490
box -36 -24 336 816
use AND2X2  _1050_
timestamp 1727136778
transform 1 0 4530 0 -1 3930
box -36 -24 336 819
use OAI21X1  _1051_
timestamp 1727136778
transform -1 0 2430 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1052_
timestamp 1727136778
transform 1 0 3690 0 -1 3930
box -36 -24 336 816
use NAND3X1  _1053_
timestamp 1727136778
transform 1 0 3690 0 1 3930
box -36 -24 336 816
use NAND2X1  _1054_
timestamp 1727136778
transform -1 0 4410 0 -1 3930
box -36 -24 276 816
use NAND3X1  _1055_
timestamp 1727136778
transform -1 0 3210 0 1 2370
box -36 -24 336 816
use NAND3X1  _1056_
timestamp 1727136778
transform 1 0 3090 0 -1 2370
box -36 -24 336 816
use OAI21X1  _1057_
timestamp 1727136778
transform -1 0 6030 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1058_
timestamp 1727136778
transform 1 0 3870 0 1 2370
box -36 -24 336 816
use OAI21X1  _1059_
timestamp 1727136778
transform 1 0 3390 0 1 2370
box -36 -24 336 816
use NAND3X1  _1060_
timestamp 1727136778
transform -1 0 3810 0 -1 2370
box -36 -24 336 816
use INVX4  _1061_
timestamp 1727136778
transform -1 0 9090 0 1 11730
box -36 -24 276 816
use NOR2X1  _1062_
timestamp 1727136778
transform -1 0 6030 0 -1 3930
box -36 -24 276 816
use OAI21X1  _1063_
timestamp 1727136778
transform 1 0 6570 0 -1 3930
box -36 -24 336 816
use XNOR2X1  _1064_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727153789
transform 1 0 4230 0 1 810
box -36 -24 456 816
use INVX1  _1065_
timestamp 1727136778
transform -1 0 3030 0 -1 810
box -36 -24 216 816
use NAND3X1  _1066_
timestamp 1727136778
transform 1 0 3150 0 -1 810
box -36 -24 336 816
use AOI21X1  _1067_
timestamp 1727136778
transform 1 0 3990 0 -1 2370
box -36 -24 336 816
use AOI21X1  _1068_
timestamp 1727136778
transform -1 0 2910 0 -1 2370
box -36 -24 336 816
use OAI21X1  _1069_
timestamp 1727136778
transform 1 0 3750 0 1 810
box -36 -24 336 816
use NAND3X1  _1070_
timestamp 1727136778
transform 1 0 5970 0 -1 810
box -36 -24 336 816
use NAND2X1  _1071_
timestamp 1727136778
transform 1 0 4830 0 1 810
box -36 -24 276 816
use INVX1  _1072_
timestamp 1727136778
transform -1 0 810 0 -1 810
box -36 -24 216 816
use OAI21X1  _1073_
timestamp 1727136778
transform -1 0 3210 0 1 810
box -36 -24 336 816
use AOI21X1  _1074_
timestamp 1727136778
transform -1 0 2730 0 1 2370
box -36 -24 336 816
use OAI21X1  _1075_
timestamp 1727136778
transform -1 0 2670 0 1 5490
box -36 -24 336 816
use NAND3X1  _1076_
timestamp 1727136778
transform -1 0 3270 0 -1 7050
box -36 -24 336 816
use AOI22X1  _1077_
timestamp 1727136778
transform 1 0 3450 0 -1 7050
box -42 -24 396 816
use INVX1  _1078_
timestamp 1727136778
transform -1 0 1650 0 1 7050
box -36 -24 216 816
use NAND2X1  _1079_
timestamp 1727136778
transform -1 0 2970 0 1 7050
box -36 -24 276 816
use INVX1  _1080_
timestamp 1727136778
transform -1 0 2790 0 -1 7050
box -36 -24 216 816
use NAND3X1  _1081_
timestamp 1727136778
transform -1 0 990 0 -1 7050
box -36 -24 336 816
use NAND2X1  _1082_
timestamp 1727136778
transform -1 0 3330 0 1 7050
box -36 -24 276 816
use NOR2X1  _1083_
timestamp 1727136778
transform -1 0 2550 0 1 7050
box -36 -24 276 816
use OAI21X1  _1084_
timestamp 1727136778
transform -1 0 1470 0 -1 7050
box -36 -24 336 816
use AOI21X1  _1085_
timestamp 1727136778
transform -1 0 1350 0 1 5490
box -36 -24 336 816
use OAI21X1  _1086_
timestamp 1727136778
transform 1 0 2130 0 -1 7050
box -36 -24 336 816
use NAND3X1  _1087_
timestamp 1727136778
transform 1 0 1650 0 -1 7050
box -36 -24 336 816
use AOI22X1  _1088_
timestamp 1727136778
transform -1 0 2250 0 -1 5490
box -42 -24 396 816
use NAND2X1  _1089_
timestamp 1727136778
transform 1 0 5970 0 -1 8610
box -36 -24 276 816
use INVX1  _1090_
timestamp 1727136778
transform 1 0 4770 0 -1 8610
box -36 -24 216 816
use AND2X2  _1091_
timestamp 1727136778
transform -1 0 5970 0 -1 7050
box -36 -24 336 819
use AND2X2  _1092_
timestamp 1727136778
transform -1 0 6450 0 1 7050
box -36 -24 336 819
use NAND2X1  _1093_
timestamp 1727136778
transform 1 0 5730 0 1 7050
box -36 -24 276 816
use AOI22X1  _1094_
timestamp 1727136778
transform 1 0 6570 0 1 10170
box -42 -24 396 816
use INVX1  _1095_
timestamp 1727136778
transform -1 0 5790 0 -1 8610
box -36 -24 216 816
use NAND3X1  _1096_
timestamp 1727136778
transform -1 0 5430 0 -1 8610
box -36 -24 336 816
use OAI21X1  _1097_
timestamp 1727136778
transform -1 0 5070 0 1 7050
box -36 -24 336 816
use OAI21X1  _1098_
timestamp 1727136778
transform -1 0 5550 0 1 7050
box -36 -24 336 816
use NAND3X1  _1099_
timestamp 1727136778
transform -1 0 4650 0 1 7050
box -36 -24 336 816
use AND2X2  _1100_
timestamp 1727136778
transform -1 0 450 0 1 7050
box -36 -24 336 819
use OAI21X1  _1101_
timestamp 1727136778
transform -1 0 510 0 -1 5490
box -36 -24 336 816
use AOI21X1  _1102_
timestamp 1727136778
transform -1 0 3150 0 1 5490
box -36 -24 336 816
use NAND3X1  _1103_
timestamp 1727136778
transform 1 0 1950 0 1 5490
box -36 -24 336 816
use NAND3X1  _1104_
timestamp 1727136778
transform 1 0 1470 0 1 5490
box -36 -24 336 816
use NAND2X1  _1105_
timestamp 1727136778
transform 1 0 630 0 1 7050
box -36 -24 276 816
use NAND3X1  _1106_
timestamp 1727136778
transform -1 0 510 0 1 5490
box -36 -24 336 816
use NAND3X1  _1107_
timestamp 1727136778
transform 1 0 630 0 1 2370
box -36 -24 336 816
use OAI21X1  _1108_
timestamp 1727136778
transform 1 0 2730 0 -1 3930
box -36 -24 336 816
use NAND3X1  _1109_
timestamp 1727136778
transform -1 0 1410 0 -1 5490
box -36 -24 336 816
use OAI21X1  _1110_
timestamp 1727136778
transform -1 0 930 0 -1 5490
box -36 -24 336 816
use NAND3X1  _1111_
timestamp 1727136778
transform -1 0 510 0 1 3930
box -36 -24 336 816
use NAND2X1  _1112_
timestamp 1727136778
transform -1 0 6390 0 -1 7050
box -36 -24 276 816
use INVX1  _1113_
timestamp 1727136778
transform 1 0 1470 0 -1 3930
box -36 -24 216 816
use AOI22X1  _1114_
timestamp 1727136778
transform -1 0 5730 0 -1 5490
box -42 -24 396 816
use INVX1  _1115_
timestamp 1727136778
transform -1 0 1770 0 -1 5490
box -36 -24 216 816
use OAI21X1  _1116_
timestamp 1727136778
transform -1 0 2190 0 1 3930
box -36 -24 336 816
use NOR2X1  _1117_
timestamp 1727136778
transform 1 0 2370 0 1 3930
box -36 -24 276 816
use NAND2X1  _1118_
timestamp 1727136778
transform -1 0 1350 0 1 3930
box -36 -24 276 816
use NAND3X1  _1119_
timestamp 1727136778
transform 1 0 1530 0 1 2370
box -36 -24 336 816
use NAND2X1  _1120_
timestamp 1727136778
transform 1 0 1530 0 1 3930
box -36 -24 276 816
use OAI21X1  _1121_
timestamp 1727136778
transform 1 0 2790 0 1 3930
box -36 -24 336 816
use NAND3X1  _1122_
timestamp 1727136778
transform -1 0 2550 0 -1 3930
box -36 -24 336 816
use NAND2X1  _1123_
timestamp 1727136778
transform -1 0 2250 0 1 2370
box -36 -24 276 816
use NAND3X1  _1124_
timestamp 1727136778
transform 1 0 1650 0 -1 2370
box -36 -24 336 816
use AOI21X1  _1125_
timestamp 1727136778
transform 1 0 630 0 1 3930
box -36 -24 336 816
use AOI21X1  _1126_
timestamp 1727136778
transform -1 0 510 0 1 2370
box -36 -24 336 816
use NAND3X1  _1127_
timestamp 1727136778
transform 1 0 1830 0 -1 3930
box -36 -24 336 816
use NAND3X1  _1128_
timestamp 1727136778
transform -1 0 1350 0 -1 3930
box -36 -24 336 816
use NAND2X1  _1129_
timestamp 1727136778
transform -1 0 870 0 -1 3930
box -36 -24 276 816
use OAI21X1  _1130_
timestamp 1727136778
transform 1 0 1170 0 -1 2370
box -36 -24 336 816
use AOI21X1  _1131_
timestamp 1727136778
transform -1 0 1410 0 1 810
box -36 -24 336 816
use AOI21X1  _1132_
timestamp 1727136778
transform -1 0 2730 0 1 810
box -36 -24 336 816
use OAI21X1  _1133_
timestamp 1727136778
transform -1 0 510 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1134_
timestamp 1727136778
transform -1 0 990 0 -1 2370
box -36 -24 336 816
use AOI21X1  _1135_
timestamp 1727136778
transform 1 0 630 0 1 810
box -36 -24 336 816
use OAI21X1  _1136_
timestamp 1727136778
transform -1 0 1290 0 -1 810
box -36 -24 336 816
use NAND3X1  _1137_
timestamp 1727136778
transform -1 0 510 0 1 810
box -36 -24 336 816
use NAND3X1  _1138_
timestamp 1727136778
transform 1 0 1530 0 1 810
box -36 -24 336 816
use NAND3X1  _1139_
timestamp 1727136778
transform 1 0 1890 0 -1 810
box -36 -24 336 816
use AOI21X1  _1140_
timestamp 1727136778
transform 1 0 5490 0 -1 810
box -36 -24 336 816
use INVX1  _1141_
timestamp 1727136778
transform 1 0 6870 0 -1 810
box -36 -24 216 816
use INVX1  _1142_
timestamp 1727136778
transform 1 0 7650 0 1 810
box -36 -24 216 816
use NOR2X1  _1143_
timestamp 1727136778
transform 1 0 10050 0 1 3930
box -36 -24 276 816
use INVX1  _1144_
timestamp 1727136778
transform 1 0 11010 0 -1 3930
box -36 -24 216 816
use OAI21X1  _1145_
timestamp 1727136778
transform 1 0 9150 0 1 5490
box -36 -24 336 816
use AOI21X1  _1146_
timestamp 1727136778
transform -1 0 10410 0 -1 3930
box -36 -24 336 816
use OAI21X1  _1147_
timestamp 1727136778
transform -1 0 9030 0 1 3930
box -36 -24 336 816
use NAND3X1  _1148_
timestamp 1727136778
transform 1 0 9630 0 -1 3930
box -36 -24 336 816
use AOI21X1  _1149_
timestamp 1727136778
transform -1 0 9930 0 1 2370
box -36 -24 336 816
use AND2X2  _1150_
timestamp 1727136778
transform 1 0 8550 0 -1 2370
box -36 -24 336 819
use NAND3X1  _1151_
timestamp 1727136778
transform 1 0 10050 0 1 2370
box -36 -24 336 816
use AOI21X1  _1152_
timestamp 1727136778
transform -1 0 9870 0 -1 2370
box -36 -24 336 816
use OAI21X1  _1153_
timestamp 1727136778
transform 1 0 7170 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1154_
timestamp 1727136778
transform 1 0 7590 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1155_
timestamp 1727136778
transform 1 0 8070 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1156_
timestamp 1727136778
transform -1 0 8310 0 1 810
box -36 -24 336 816
use OAI21X1  _1157_
timestamp 1727136778
transform -1 0 3630 0 1 810
box -36 -24 336 816
use NAND3X1  _1158_
timestamp 1727136778
transform 1 0 3630 0 -1 810
box -36 -24 336 816
use AOI22X1  _1159_
timestamp 1727136778
transform -1 0 5610 0 1 810
box -42 -24 396 816
use NAND3X1  _1160_
timestamp 1727136778
transform 1 0 1410 0 -1 810
box -36 -24 336 816
use OAI21X1  _1161_
timestamp 1727136778
transform 1 0 2370 0 -1 810
box -36 -24 336 816
use AOI21X1  _1162_
timestamp 1727136778
transform 1 0 4110 0 -1 810
box -36 -24 336 816
use NAND3X1  _1163_
timestamp 1727136778
transform 1 0 9990 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1164_
timestamp 1727136778
transform 1 0 11370 0 -1 3930
box -36 -24 336 816
use NAND2X1  _1165_
timestamp 1727136778
transform -1 0 12030 0 1 5490
box -36 -24 276 816
use OR2X2  _1166_
timestamp 1727136778
transform 1 0 12510 0 -1 5490
box -36 -24 336 816
use NAND2X1  _1167_
timestamp 1727136778
transform 1 0 12990 0 -1 5490
box -36 -24 276 816
use AOI22X1  _1168_
timestamp 1727136778
transform -1 0 10830 0 1 5490
box -42 -24 396 816
use OAI21X1  _1169_
timestamp 1727136778
transform 1 0 12090 0 -1 5490
box -36 -24 336 816
use OAI21X1  _1170_
timestamp 1727136778
transform 1 0 10590 0 -1 3930
box -36 -24 336 816
use NAND3X1  _1171_
timestamp 1727136778
transform 1 0 12270 0 -1 3930
box -36 -24 336 816
use AOI21X1  _1172_
timestamp 1727136778
transform 1 0 11790 0 -1 3930
box -36 -24 336 816
use OAI21X1  _1173_
timestamp 1727136778
transform 1 0 12270 0 1 2370
box -36 -24 336 816
use OAI21X1  _1174_
timestamp 1727136778
transform 1 0 10890 0 -1 2370
box -36 -24 336 816
use NAND3X1  _1175_
timestamp 1727136778
transform -1 0 11670 0 -1 2370
box -36 -24 336 816
use INVX1  _1176_
timestamp 1727136778
transform 1 0 11010 0 1 810
box -36 -24 216 816
use AOI22X1  _1177_
timestamp 1727136778
transform -1 0 9390 0 -1 2370
box -42 -24 396 816
use OAI21X1  _1178_
timestamp 1727136778
transform -1 0 9270 0 1 810
box -36 -24 336 816
use NAND3X1  _1179_
timestamp 1727136778
transform 1 0 10110 0 1 810
box -36 -24 336 816
use AOI21X1  _1180_
timestamp 1727136778
transform 1 0 6450 0 -1 810
box -36 -24 336 816
use NOR3X1  _1181_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 9990 0 -1 810
box -36 -24 576 819
use INVX1  _1182_
timestamp 1727136778
transform -1 0 12090 0 1 2370
box -36 -24 216 816
use NAND3X1  _1183_
timestamp 1727136778
transform 1 0 11490 0 1 2370
box -36 -24 336 816
use INVX1  _1184_
timestamp 1727136778
transform -1 0 11190 0 1 5490
box -36 -24 216 816
use OAI21X1  _1185_
timestamp 1727136778
transform -1 0 11610 0 1 5490
box -36 -24 336 816
use OR2X2  _1186_
timestamp 1727136778
transform 1 0 12210 0 1 3930
box -36 -24 336 816
use NAND2X1  _1187_
timestamp 1727136778
transform -1 0 10290 0 1 5490
box -36 -24 276 816
use NOR2X1  _1188_
timestamp 1727136778
transform -1 0 13590 0 -1 5490
box -36 -24 276 816
use INVX1  _1189_
timestamp 1727136778
transform 1 0 11370 0 1 3930
box -36 -24 216 816
use OAI21X1  _1190_
timestamp 1727136778
transform 1 0 11730 0 1 3930
box -36 -24 336 816
use NAND3X1  _1191_
timestamp 1727136778
transform -1 0 12930 0 1 3930
box -36 -24 336 816
use INVX1  _1192_
timestamp 1727136778
transform 1 0 13530 0 -1 3930
box -36 -24 216 816
use INVX1  _1193_
timestamp 1727136778
transform 1 0 13170 0 1 2370
box -36 -24 216 816
use OAI21X1  _1194_
timestamp 1727136778
transform 1 0 12690 0 1 2370
box -36 -24 336 816
use NAND3X1  _1195_
timestamp 1727136778
transform 1 0 13530 0 1 2370
box -36 -24 336 816
use AOI21X1  _1196_
timestamp 1727136778
transform 1 0 11850 0 -1 2370
box -36 -24 336 816
use NOR3X1  _1197_
timestamp 1727136778
transform -1 0 12870 0 -1 2370
box -36 -24 576 819
use OAI21X1  _1198_
timestamp 1727136778
transform 1 0 9390 0 1 810
box -36 -24 336 816
use NAND3X1  _1199_
timestamp 1727136778
transform 1 0 8490 0 1 810
box -36 -24 336 816
use NAND3X1  _1200_
timestamp 1727136778
transform 1 0 10590 0 1 810
box -36 -24 336 816
use NAND3X1  _1201_
timestamp 1727136778
transform -1 0 11610 0 1 810
box -36 -24 336 816
use INVX1  _1202_
timestamp 1727136778
transform 1 0 12270 0 1 810
box -36 -24 216 816
use OAI21X1  _1203_
timestamp 1727136778
transform 1 0 10710 0 -1 810
box -36 -24 336 816
use AOI21X1  _1204_
timestamp 1727136778
transform -1 0 11430 0 -1 810
box -36 -24 336 816
use OAI21X1  _1205_
timestamp 1727136778
transform 1 0 8130 0 -1 810
box -36 -24 336 816
use AOI21X1  _1206_
timestamp 1727136778
transform -1 0 510 0 -1 810
box -36 -24 336 816
use NAND2X1  _1207_
timestamp 1727136778
transform 1 0 2370 0 -1 5490
box -36 -24 276 816
use OAI21X1  _1208_
timestamp 1727136778
transform -1 0 510 0 -1 3930
box -36 -24 336 816
use NAND2X1  _1209_
timestamp 1727136778
transform 1 0 7230 0 -1 10170
box -36 -24 276 816
use INVX1  _1210_
timestamp 1727136778
transform -1 0 4830 0 -1 10170
box -36 -24 216 816
use NOR2X1  _1211_
timestamp 1727136778
transform -1 0 6810 0 -1 7050
box -36 -24 276 816
use OAI21X1  _1212_
timestamp 1727136778
transform 1 0 5610 0 1 8610
box -36 -24 336 816
use NAND2X1  _1213_
timestamp 1727136778
transform 1 0 6330 0 -1 10170
box -36 -24 276 816
use OR2X2  _1214_
timestamp 1727136778
transform 1 0 6750 0 -1 10170
box -36 -24 336 816
use NAND3X1  _1215_
timestamp 1727136778
transform -1 0 4530 0 -1 10170
box -36 -24 336 816
use AND2X2  _1216_
timestamp 1727136778
transform -1 0 6210 0 -1 10170
box -36 -24 336 819
use NOR2X1  _1217_
timestamp 1727136778
transform 1 0 6090 0 1 8610
box -36 -24 276 816
use OAI21X1  _1218_
timestamp 1727136778
transform -1 0 5790 0 -1 10170
box -36 -24 336 816
use NAND2X1  _1219_
timestamp 1727136778
transform 1 0 3810 0 -1 10170
box -36 -24 276 816
use AOI21X1  _1220_
timestamp 1727136778
transform -1 0 930 0 1 5490
box -36 -24 336 816
use NAND2X1  _1221_
timestamp 1727136778
transform -1 0 4890 0 -1 11730
box -36 -24 276 816
use AND2X2  _1222_
timestamp 1727136778
transform -1 0 6090 0 -1 13290
box -36 -24 336 819
use OAI21X1  _1223_
timestamp 1727136778
transform 1 0 5430 0 -1 11730
box -36 -24 336 816
use AND2X2  _1224_
timestamp 1727136778
transform -1 0 6690 0 -1 11730
box -36 -24 336 819
use OAI21X1  _1225_
timestamp 1727136778
transform 1 0 5910 0 -1 11730
box -36 -24 336 816
use NAND3X1  _1226_
timestamp 1727136778
transform -1 0 5310 0 -1 11730
box -36 -24 336 816
use INVX1  _1227_
timestamp 1727136778
transform 1 0 4830 0 1 11730
box -36 -24 216 816
use NAND2X1  _1228_
timestamp 1727136778
transform 1 0 6030 0 1 11730
box -36 -24 276 816
use AOI22X1  _1229_
timestamp 1727136778
transform 1 0 6750 0 1 11730
box -42 -24 396 816
use INVX1  _1230_
timestamp 1727136778
transform 1 0 5670 0 1 11730
box -36 -24 216 816
use NAND3X1  _1231_
timestamp 1727136778
transform -1 0 5490 0 1 11730
box -36 -24 336 816
use NAND2X1  _1232_
timestamp 1727136778
transform 1 0 2370 0 -1 11730
box -36 -24 276 816
use AOI21X1  _1233_
timestamp 1727136778
transform 1 0 1050 0 1 7050
box -36 -24 336 816
use NAND2X1  _1234_
timestamp 1727136778
transform 1 0 3450 0 -1 13290
box -36 -24 276 816
use XOR2X1  _1235_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727152697
transform 1 0 2850 0 1 11730
box -36 -24 453 816
use NAND2X1  _1236_
timestamp 1727136778
transform -1 0 1170 0 1 10170
box -36 -24 276 816
use OAI21X1  _1237_
timestamp 1727136778
transform 1 0 1830 0 1 7050
box -36 -24 336 816
use XNOR2X1  _1238_
timestamp 1727153789
transform 1 0 2310 0 1 11730
box -36 -24 456 816
use NAND2X1  _1239_
timestamp 1727136778
transform -1 0 1830 0 -1 11730
box -36 -24 276 816
use NAND3X1  _1240_
timestamp 1727136778
transform -1 0 1650 0 1 10170
box -36 -24 336 816
use AND2X2  _1241_
timestamp 1727136778
transform -1 0 990 0 -1 11730
box -36 -24 336 819
use NAND2X1  _1242_
timestamp 1727136778
transform 1 0 2010 0 -1 11730
box -36 -24 276 816
use NAND2X1  _1243_
timestamp 1727136778
transform 1 0 1170 0 -1 11730
box -36 -24 276 816
use NAND3X1  _1244_
timestamp 1727136778
transform 1 0 690 0 1 11730
box -36 -24 336 816
use NAND3X1  _1245_
timestamp 1727136778
transform -1 0 930 0 -1 10170
box -36 -24 336 816
use OAI21X1  _1246_
timestamp 1727136778
transform -1 0 510 0 -1 7050
box -36 -24 336 816
use AOI22X1  _1247_
timestamp 1727136778
transform -1 0 570 0 -1 11730
box -42 -24 396 816
use AOI21X1  _1248_
timestamp 1727136778
transform 1 0 1770 0 1 10170
box -36 -24 336 816
use OAI21X1  _1249_
timestamp 1727136778
transform 1 0 210 0 1 8610
box -36 -24 336 816
use NAND3X1  _1250_
timestamp 1727136778
transform -1 0 990 0 1 8610
box -36 -24 336 816
use AND2X2  _1251_
timestamp 1727136778
transform -1 0 3630 0 -1 10170
box -36 -24 336 819
use NAND3X1  _1252_
timestamp 1727136778
transform 1 0 1530 0 -1 10170
box -36 -24 336 816
use OAI21X1  _1253_
timestamp 1727136778
transform 1 0 210 0 -1 10170
box -36 -24 336 816
use NAND3X1  _1254_
timestamp 1727136778
transform -1 0 2250 0 -1 10170
box -36 -24 336 816
use NAND3X1  _1255_
timestamp 1727136778
transform -1 0 510 0 -1 8610
box -36 -24 336 816
use AOI21X1  _1256_
timestamp 1727136778
transform 1 0 1110 0 1 2370
box -36 -24 336 816
use AOI22X1  _1257_
timestamp 1727136778
transform -1 0 3210 0 -1 10170
box -42 -24 396 816
use AOI21X1  _1258_
timestamp 1727136778
transform 1 0 1170 0 1 8610
box -36 -24 336 816
use OAI21X1  _1259_
timestamp 1727136778
transform -1 0 2850 0 1 8610
box -36 -24 336 816
use AOI21X1  _1260_
timestamp 1727136778
transform -1 0 2790 0 -1 8610
box -36 -24 336 816
use INVX1  _1261_
timestamp 1727136778
transform 1 0 2970 0 -1 8610
box -36 -24 216 816
use NAND3X1  _1262_
timestamp 1727136778
transform 1 0 690 0 -1 8610
box -36 -24 336 816
use OAI21X1  _1263_
timestamp 1727136778
transform -1 0 2370 0 1 8610
box -36 -24 336 816
use AOI21X1  _1264_
timestamp 1727136778
transform 1 0 1590 0 -1 8610
box -36 -24 336 816
use OAI21X1  _1265_
timestamp 1727136778
transform -1 0 2370 0 -1 8610
box -36 -24 336 816
use OAI21X1  _1266_
timestamp 1727136778
transform -1 0 2310 0 1 810
box -36 -24 336 816
use NAND3X1  _1267_
timestamp 1727136778
transform -1 0 1410 0 -1 8610
box -36 -24 336 816
use NAND3X1  _1268_
timestamp 1727136778
transform 1 0 3330 0 -1 8610
box -36 -24 336 816
use NAND3X1  _1269_
timestamp 1727136778
transform 1 0 3810 0 -1 8610
box -36 -24 336 816
use AND2X2  _1270_
timestamp 1727136778
transform 1 0 7110 0 -1 8610
box -36 -24 336 819
use XOR2X1  _1271_
timestamp 1727152697
transform -1 0 9750 0 -1 8610
box -36 -24 453 816
use NOR2X1  _1272_
timestamp 1727136778
transform 1 0 15090 0 -1 10170
box -36 -24 276 816
use NOR2X1  _1273_
timestamp 1727136778
transform -1 0 14490 0 -1 8610
box -36 -24 276 816
use OAI21X1  _1274_
timestamp 1727136778
transform 1 0 12570 0 -1 8610
box -36 -24 336 816
use AOI21X1  _1275_
timestamp 1727136778
transform 1 0 11970 0 1 7050
box -36 -24 336 816
use OAI21X1  _1276_
timestamp 1727136778
transform -1 0 13710 0 -1 8610
box -36 -24 336 816
use OAI21X1  _1277_
timestamp 1727136778
transform 1 0 12450 0 1 7050
box -36 -24 336 816
use NAND2X1  _1278_
timestamp 1727136778
transform 1 0 14370 0 1 5490
box -36 -24 276 816
use OAI21X1  _1279_
timestamp 1727136778
transform 1 0 14190 0 -1 5490
box -36 -24 336 816
use INVX1  _1280_
timestamp 1727136778
transform -1 0 10890 0 -1 7050
box -36 -24 216 816
use INVX1  _1281_
timestamp 1727136778
transform -1 0 11790 0 1 7050
box -36 -24 216 816
use OAI21X1  _1282_
timestamp 1727136778
transform -1 0 12510 0 -1 7050
box -36 -24 336 816
use OAI21X1  _1283_
timestamp 1727136778
transform -1 0 11430 0 1 7050
box -36 -24 336 816
use NAND3X1  _1284_
timestamp 1727136778
transform -1 0 5310 0 -1 810
box -36 -24 336 816
use INVX1  _1285_
timestamp 1727136778
transform -1 0 9990 0 1 810
box -36 -24 216 816
use NAND2X1  _1286_
timestamp 1727136778
transform -1 0 4830 0 -1 810
box -36 -24 276 816
use NAND3X1  _1287_
timestamp 1727136778
transform 1 0 5790 0 1 810
box -36 -24 336 816
use NAND3X1  _1288_
timestamp 1727136778
transform 1 0 9030 0 -1 810
box -36 -24 336 816
use AOI21X1  _1289_
timestamp 1727136778
transform 1 0 8610 0 -1 810
box -36 -24 336 816
use OAI21X1  _1290_
timestamp 1727136778
transform -1 0 9810 0 -1 810
box -36 -24 336 816
use AOI21X1  _1291_
timestamp 1727136778
transform -1 0 7530 0 -1 810
box -36 -24 336 816
use NAND2X1  _1292_
timestamp 1727136778
transform -1 0 6990 0 -1 8610
box -36 -24 276 816
use OAI21X1  _1293_
timestamp 1727136778
transform -1 0 8250 0 -1 8610
box -36 -24 336 816
use INVX1  _1294_
timestamp 1727136778
transform 1 0 3870 0 1 8610
box -36 -24 216 816
use AOI21X1  _1295_
timestamp 1727136778
transform 1 0 3390 0 1 8610
box -36 -24 336 816
use OAI21X1  _1296_
timestamp 1727136778
transform -1 0 5310 0 -1 10170
box -36 -24 336 816
use INVX1  _1297_
timestamp 1727136778
transform 1 0 4950 0 1 10170
box -36 -24 216 816
use AOI21X1  _1298_
timestamp 1727136778
transform 1 0 1050 0 -1 10170
box -36 -24 336 816
use OAI21X1  _1299_
timestamp 1727136778
transform 1 0 2430 0 -1 10170
box -36 -24 336 816
use NAND2X1  _1300_
timestamp 1727136778
transform -1 0 5130 0 -1 13290
box -36 -24 276 816
use NOR2X1  _1301_
timestamp 1727136778
transform 1 0 6210 0 1 10170
box -36 -24 276 816
use NAND2X1  _1302_
timestamp 1727136778
transform -1 0 6030 0 1 13290
box -36 -24 276 816
use NAND2X1  _1303_
timestamp 1727136778
transform -1 0 6510 0 -1 13290
box -36 -24 276 816
use OAI22X1  _1304_
timestamp 1727136778
transform -1 0 5610 0 -1 13290
box -36 -24 396 816
use XNOR2X1  _1305_
timestamp 1727153789
transform -1 0 4710 0 -1 13290
box -36 -24 456 816
use XNOR2X1  _1306_
timestamp 1727153789
transform 1 0 2430 0 -1 13290
box -36 -24 456 816
use NOR2X1  _1307_
timestamp 1727136778
transform 1 0 1110 0 1 11730
box -36 -24 276 816
use AOI21X1  _1308_
timestamp 1727136778
transform -1 0 510 0 1 11730
box -36 -24 336 816
use NAND2X1  _1309_
timestamp 1727136778
transform 1 0 4050 0 1 13290
box -36 -24 276 816
use NAND2X1  _1310_
timestamp 1727136778
transform 1 0 4890 0 -1 14850
box -36 -24 276 816
use INVX1  _1311_
timestamp 1727136778
transform 1 0 3390 0 -1 14850
box -36 -24 216 816
use AND2X2  _1312_
timestamp 1727136778
transform -1 0 5610 0 -1 14850
box -36 -24 336 819
use AND2X2  _1313_
timestamp 1727136778
transform -1 0 4410 0 -1 14850
box -36 -24 336 819
use NAND2X1  _1314_
timestamp 1727136778
transform -1 0 3930 0 -1 14850
box -36 -24 276 816
use AOI22X1  _1315_
timestamp 1727136778
transform 1 0 3990 0 1 14850
box -42 -24 396 816
use INVX1  _1316_
timestamp 1727136778
transform -1 0 2550 0 1 14850
box -36 -24 216 816
use AOI21X1  _1317_
timestamp 1727136778
transform 1 0 2910 0 -1 14850
box -36 -24 336 816
use INVX2  _1318_
timestamp 1727136778
transform 1 0 8430 0 1 13290
box -36 -24 216 816
use OAI21X1  _1319_
timestamp 1727136778
transform -1 0 6510 0 1 13290
box -36 -24 336 816
use OAI21X1  _1320_
timestamp 1727136778
transform -1 0 5610 0 1 13290
box -36 -24 336 816
use AOI21X1  _1321_
timestamp 1727136778
transform -1 0 5190 0 1 13290
box -36 -24 336 816
use OAI22X1  _1322_
timestamp 1727136778
transform -1 0 3870 0 1 13290
box -36 -24 396 816
use NAND3X1  _1323_
timestamp 1727136778
transform -1 0 4710 0 1 13290
box -36 -24 336 816
use NAND3X1  _1324_
timestamp 1727136778
transform -1 0 2790 0 -1 14850
box -36 -24 336 816
use NOR2X1  _1325_
timestamp 1727136778
transform -1 0 3330 0 1 13290
box -36 -24 276 816
use NAND3X1  _1326_
timestamp 1727136778
transform -1 0 2310 0 -1 14850
box -36 -24 336 816
use NAND2X1  _1327_
timestamp 1727136778
transform -1 0 450 0 -1 14850
box -36 -24 276 816
use NOR2X1  _1328_
timestamp 1727136778
transform -1 0 450 0 -1 13290
box -36 -24 276 816
use NOR2X1  _1329_
timestamp 1727136778
transform 1 0 1950 0 1 11730
box -36 -24 276 816
use OAI21X1  _1330_
timestamp 1727136778
transform -1 0 1830 0 1 11730
box -36 -24 336 816
use AOI21X1  _1331_
timestamp 1727136778
transform 1 0 630 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1332_
timestamp 1727136778
transform 1 0 1470 0 -1 13290
box -36 -24 336 816
use XOR2X1  _1333_
timestamp 1727152697
transform 1 0 2490 0 1 13290
box -36 -24 453 816
use NAND3X1  _1334_
timestamp 1727136778
transform 1 0 1590 0 -1 14850
box -36 -24 336 816
use NAND2X1  _1335_
timestamp 1727136778
transform -1 0 390 0 1 13290
box -36 -24 276 816
use NAND3X1  _1336_
timestamp 1727136778
transform 1 0 1530 0 1 13290
box -36 -24 336 816
use NAND3X1  _1337_
timestamp 1727136778
transform 1 0 3450 0 1 11730
box -36 -24 336 816
use NOR3X1  _1338_
timestamp 1727136778
transform 1 0 210 0 1 10170
box -36 -24 576 819
use AOI21X1  _1339_
timestamp 1727136778
transform 1 0 2190 0 1 10170
box -36 -24 336 816
use AOI21X1  _1340_
timestamp 1727136778
transform 1 0 2010 0 1 13290
box -36 -24 336 816
use NAND3X1  _1341_
timestamp 1727136778
transform 1 0 570 0 1 13290
box -36 -24 336 816
use OAI21X1  _1342_
timestamp 1727136778
transform -1 0 870 0 -1 13290
box -36 -24 336 816
use AOI21X1  _1343_
timestamp 1727136778
transform 1 0 1050 0 -1 13290
box -36 -24 336 816
use OAI21X1  _1344_
timestamp 1727136778
transform -1 0 2970 0 1 10170
box -36 -24 336 816
use NAND3X1  _1345_
timestamp 1727136778
transform -1 0 4770 0 1 10170
box -36 -24 336 816
use NAND3X1  _1346_
timestamp 1727136778
transform 1 0 2790 0 -1 11730
box -36 -24 336 816
use OAI21X1  _1347_
timestamp 1727136778
transform 1 0 3150 0 1 10170
box -36 -24 336 816
use NAND3X1  _1348_
timestamp 1727136778
transform -1 0 4350 0 1 10170
box -36 -24 336 816
use NAND3X1  _1349_
timestamp 1727136778
transform -1 0 4530 0 1 8610
box -36 -24 336 816
use AOI21X1  _1350_
timestamp 1727136778
transform 1 0 1650 0 1 8610
box -36 -24 336 816
use OAI21X1  _1351_
timestamp 1727136778
transform 1 0 2970 0 1 8610
box -36 -24 336 816
use NAND3X1  _1352_
timestamp 1727136778
transform 1 0 5310 0 1 10170
box -36 -24 336 816
use NAND3X1  _1353_
timestamp 1727136778
transform -1 0 3930 0 1 10170
box -36 -24 336 816
use NAND3X1  _1354_
timestamp 1727136778
transform 1 0 5130 0 1 8610
box -36 -24 336 816
use NAND2X1  _1355_
timestamp 1727136778
transform -1 0 6750 0 1 8610
box -36 -24 276 816
use AND2X2  _1356_
timestamp 1727136778
transform 1 0 9930 0 -1 8610
box -36 -24 336 819
use OAI21X1  _1357_
timestamp 1727136778
transform 1 0 10350 0 -1 8610
box -36 -24 336 816
use OAI21X1  _1358_
timestamp 1727136778
transform 1 0 10830 0 -1 8610
box -36 -24 336 816
use AND2X2  _1359_
timestamp 1727136778
transform 1 0 13770 0 -1 5490
box -36 -24 336 819
use NAND2X1  _1360_
timestamp 1727136778
transform 1 0 13590 0 1 5490
box -36 -24 276 816
use OAI21X1  _1361_
timestamp 1727136778
transform -1 0 12930 0 1 5490
box -36 -24 336 816
use OAI21X1  _1362_
timestamp 1727136778
transform 1 0 13110 0 1 5490
box -36 -24 336 816
use AOI21X1  _1363_
timestamp 1727136778
transform -1 0 12510 0 1 5490
box -36 -24 336 816
use AOI22X1  _1364_
timestamp 1727136778
transform 1 0 11730 0 -1 7050
box -42 -24 396 816
use OAI21X1  _1365_
timestamp 1727136778
transform -1 0 14790 0 1 3930
box -36 -24 336 816
use AOI21X1  _1366_
timestamp 1727136778
transform -1 0 5010 0 1 8610
box -36 -24 336 816
use AOI22X1  _1367_
timestamp 1727136778
transform 1 0 4230 0 -1 8610
box -42 -24 396 816
use NOR2X1  _1368_
timestamp 1727136778
transform 1 0 6390 0 -1 8610
box -36 -24 276 816
use NAND3X1  _1369_
timestamp 1727136778
transform 1 0 8850 0 -1 8610
box -36 -24 336 816
use AOI21X1  _1370_
timestamp 1727136778
transform 1 0 6870 0 1 8610
box -36 -24 336 816
use INVX1  _1371_
timestamp 1727136778
transform 1 0 7590 0 -1 8610
box -36 -24 216 816
use NAND2X1  _1372_
timestamp 1727136778
transform -1 0 4110 0 -1 13290
box -36 -24 276 816
use OAI21X1  _1373_
timestamp 1727136778
transform 1 0 2970 0 -1 13290
box -36 -24 336 816
use INVX1  _1374_
timestamp 1727136778
transform -1 0 1770 0 1 14850
box -36 -24 216 816
use AOI21X1  _1375_
timestamp 1727136778
transform -1 0 1350 0 1 13290
box -36 -24 336 816
use NAND2X1  _1376_
timestamp 1727136778
transform -1 0 4110 0 1 16410
box -36 -24 276 816
use INVX1  _1377_
timestamp 1727136778
transform -1 0 2850 0 1 16410
box -36 -24 216 816
use NOR2X1  _1378_
timestamp 1727136778
transform -1 0 3810 0 1 14850
box -36 -24 276 816
use OAI21X1  _1379_
timestamp 1727136778
transform -1 0 3390 0 1 14850
box -36 -24 336 816
use NAND2X1  _1380_
timestamp 1727136778
transform -1 0 3750 0 1 16410
box -36 -24 276 816
use OR2X2  _1381_
timestamp 1727136778
transform -1 0 3330 0 1 16410
box -36 -24 336 816
use NAND3X1  _1382_
timestamp 1727136778
transform -1 0 2490 0 1 16410
box -36 -24 336 816
use AND2X2  _1383_
timestamp 1727136778
transform -1 0 3330 0 -1 17970
box -36 -24 336 819
use NOR2X1  _1384_
timestamp 1727136778
transform -1 0 3750 0 -1 17970
box -36 -24 276 816
use OAI21X1  _1385_
timestamp 1727136778
transform -1 0 2850 0 -1 17970
box -36 -24 336 816
use NAND2X1  _1386_
timestamp 1727136778
transform -1 0 930 0 -1 17970
box -36 -24 276 816
use OR2X2  _1387_
timestamp 1727136778
transform 1 0 1950 0 -1 13290
box -36 -24 336 816
use NAND2X1  _1388_
timestamp 1727136778
transform 1 0 4830 0 -1 16410
box -36 -24 276 816
use NAND2X1  _1389_
timestamp 1727136778
transform -1 0 5670 0 1 14850
box -36 -24 276 816
use NAND2X1  _1390_
timestamp 1727136778
transform -1 0 5310 0 1 14850
box -36 -24 276 816
use AOI22X1  _1391_
timestamp 1727136778
transform -1 0 4890 0 1 14850
box -42 -24 396 816
use INVX1  _1392_
timestamp 1727136778
transform 1 0 6150 0 -1 16410
box -36 -24 216 816
use OAI21X1  _1393_
timestamp 1727136778
transform 1 0 5730 0 -1 16410
box -36 -24 336 816
use XNOR2X1  _1394_
timestamp 1727153789
transform 1 0 4230 0 -1 16410
box -36 -24 456 816
use AOI21X1  _1395_
timestamp 1727136778
transform 1 0 1290 0 1 16410
box -36 -24 336 816
use NAND3X1  _1396_
timestamp 1727136778
transform -1 0 2070 0 1 16410
box -36 -24 336 816
use INVX1  _1397_
timestamp 1727136778
transform -1 0 390 0 1 17970
box -36 -24 216 816
use OAI21X1  _1398_
timestamp 1727136778
transform -1 0 1290 0 1 17970
box -36 -24 336 816
use AND2X2  _1399_
timestamp 1727136778
transform -1 0 2370 0 -1 17970
box -36 -24 336 819
use NAND2X1  _1400_
timestamp 1727136778
transform -1 0 1170 0 1 16410
box -36 -24 276 816
use INVX1  _1401_
timestamp 1727136778
transform -1 0 330 0 1 16410
box -36 -24 216 816
use NAND2X1  _1402_
timestamp 1727136778
transform -1 0 750 0 1 16410
box -36 -24 276 816
use NAND3X1  _1403_
timestamp 1727136778
transform 1 0 1110 0 -1 17970
box -36 -24 336 816
use NAND3X1  _1404_
timestamp 1727136778
transform -1 0 1770 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1405_
timestamp 1727136778
transform 1 0 1110 0 -1 14850
box -36 -24 336 816
use AOI22X1  _1406_
timestamp 1727136778
transform -1 0 570 0 -1 17970
box -42 -24 396 816
use OR2X2  _1407_
timestamp 1727136778
transform -1 0 510 0 -1 16410
box -36 -24 336 816
use NAND2X1  _1408_
timestamp 1727136778
transform -1 0 1350 0 -1 16410
box -36 -24 276 816
use AOI21X1  _1409_
timestamp 1727136778
transform -1 0 990 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1410_
timestamp 1727136778
transform 1 0 690 0 1 14850
box -36 -24 336 816
use NAND3X1  _1411_
timestamp 1727136778
transform -1 0 1410 0 1 14850
box -36 -24 336 816
use NAND3X1  _1412_
timestamp 1727136778
transform 1 0 1950 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1413_
timestamp 1727136778
transform -1 0 510 0 1 14850
box -36 -24 336 816
use NAND3X1  _1414_
timestamp 1727136778
transform -1 0 2190 0 1 14850
box -36 -24 336 816
use NAND2X1  _1415_
timestamp 1727136778
transform -1 0 4170 0 1 11730
box -36 -24 276 816
use NAND3X1  _1416_
timestamp 1727136778
transform 1 0 5790 0 1 10170
box -36 -24 336 816
use AOI21X1  _1417_
timestamp 1727136778
transform 1 0 3210 0 -1 11730
box -36 -24 336 816
use OAI21X1  _1418_
timestamp 1727136778
transform -1 0 3990 0 -1 11730
box -36 -24 336 816
use NAND3X1  _1419_
timestamp 1727136778
transform 1 0 4170 0 -1 11730
box -36 -24 336 816
use NAND2X1  _1420_
timestamp 1727136778
transform -1 0 7650 0 1 10170
box -36 -24 276 816
use AOI21X1  _1421_
timestamp 1727136778
transform -1 0 7710 0 1 7050
box -36 -24 336 816
use NAND2X1  _1422_
timestamp 1727136778
transform 1 0 8430 0 -1 8610
box -36 -24 276 816
use OAI21X1  _1423_
timestamp 1727136778
transform -1 0 8130 0 1 7050
box -36 -24 336 816
use INVX1  _1424_
timestamp 1727136778
transform 1 0 8670 0 -1 7050
box -36 -24 216 816
use NOR2X1  _1425_
timestamp 1727136778
transform -1 0 9270 0 -1 7050
box -36 -24 276 816
use OAI21X1  _1426_
timestamp 1727136778
transform 1 0 9390 0 -1 7050
box -36 -24 336 816
use NOR2X1  _1427_
timestamp 1727136778
transform 1 0 13890 0 -1 8610
box -36 -24 276 816
use NOR2X1  _1428_
timestamp 1727136778
transform -1 0 13170 0 1 7050
box -36 -24 276 816
use AOI21X1  _1429_
timestamp 1727136778
transform 1 0 13110 0 1 3930
box -36 -24 336 816
use OAI21X1  _1430_
timestamp 1727136778
transform 1 0 13530 0 1 3930
box -36 -24 336 816
use NOR2X1  _1431_
timestamp 1727136778
transform -1 0 14430 0 1 7050
box -36 -24 276 816
use NOR2X1  _1432_
timestamp 1727136778
transform 1 0 14310 0 -1 7050
box -36 -24 276 816
use AOI22X1  _1433_
timestamp 1727136778
transform -1 0 13410 0 -1 7050
box -42 -24 396 816
use OAI21X1  _1434_
timestamp 1727136778
transform 1 0 14010 0 1 3930
box -36 -24 336 816
use INVX1  _1435_
timestamp 1727136778
transform 1 0 17910 0 -1 2370
box -36 -24 216 816
use INVX1  _1436_
timestamp 1727136778
transform -1 0 17490 0 1 8610
box -36 -24 216 816
use OAI21X1  _1437_
timestamp 1727136778
transform -1 0 11970 0 -1 8610
box -36 -24 336 816
use INVX1  _1438_
timestamp 1727136778
transform 1 0 8070 0 -1 10170
box -36 -24 216 816
use OAI21X1  _1439_
timestamp 1727136778
transform 1 0 3870 0 -1 17970
box -36 -24 336 816
use INVX1  _1440_
timestamp 1727136778
transform -1 0 3810 0 1 17970
box -36 -24 216 816
use AOI21X1  _1441_
timestamp 1727136778
transform 1 0 1590 0 -1 17970
box -36 -24 336 816
use NAND2X1  _1442_
timestamp 1727136778
transform 1 0 5490 0 1 16410
box -36 -24 276 816
use INVX1  _1443_
timestamp 1727136778
transform -1 0 6450 0 -1 17970
box -36 -24 216 816
use NOR2X1  _1444_
timestamp 1727136778
transform -1 0 4530 0 1 16410
box -36 -24 276 816
use OAI22X1  _1445_
timestamp 1727136778
transform -1 0 5550 0 -1 16410
box -36 -24 396 816
use NAND2X1  _1446_
timestamp 1727136778
transform 1 0 4710 0 1 16410
box -36 -24 276 816
use NOR2X1  _1447_
timestamp 1727136778
transform 1 0 5130 0 1 16410
box -36 -24 276 816
use INVX1  _1448_
timestamp 1727136778
transform 1 0 5430 0 -1 17970
box -36 -24 216 816
use NAND3X1  _1449_
timestamp 1727136778
transform -1 0 6090 0 -1 17970
box -36 -24 336 816
use INVX1  _1450_
timestamp 1727136778
transform -1 0 4890 0 -1 17970
box -36 -24 216 816
use OAI21X1  _1451_
timestamp 1727136778
transform 1 0 5010 0 -1 17970
box -36 -24 336 816
use NAND2X1  _1452_
timestamp 1727136778
transform 1 0 5790 0 -1 14850
box -36 -24 276 816
use NAND2X1  _1453_
timestamp 1727136778
transform 1 0 6330 0 1 14850
box -36 -24 276 816
use OR2X2  _1454_
timestamp 1727136778
transform 1 0 5850 0 1 14850
box -36 -24 336 816
use INVX1  _1455_
timestamp 1727136778
transform 1 0 8670 0 -1 16410
box -36 -24 216 816
use OAI21X1  _1456_
timestamp 1727136778
transform -1 0 6810 0 -1 16410
box -36 -24 336 816
use AND2X2  _1457_
timestamp 1727136778
transform -1 0 6210 0 1 16410
box -36 -24 336 819
use AOI21X1  _1458_
timestamp 1727136778
transform -1 0 5130 0 1 17970
box -36 -24 336 816
use INVX1  _1459_
timestamp 1727136778
transform -1 0 1650 0 1 17970
box -36 -24 216 816
use NAND3X1  _1460_
timestamp 1727136778
transform 1 0 5310 0 1 17970
box -36 -24 336 816
use NAND3X1  _1461_
timestamp 1727136778
transform 1 0 2250 0 1 17970
box -36 -24 336 816
use OAI21X1  _1462_
timestamp 1727136778
transform -1 0 870 0 1 17970
box -36 -24 336 816
use INVX1  _1463_
timestamp 1727136778
transform -1 0 4530 0 -1 17970
box -36 -24 216 816
use OAI21X1  _1464_
timestamp 1727136778
transform -1 0 2970 0 1 17970
box -36 -24 336 816
use NAND3X1  _1465_
timestamp 1727136778
transform -1 0 3450 0 1 17970
box -36 -24 336 816
use NAND3X1  _1466_
timestamp 1727136778
transform -1 0 2130 0 1 17970
box -36 -24 336 816
use OAI21X1  _1467_
timestamp 1727136778
transform -1 0 4230 0 1 17970
box -36 -24 336 816
use NAND3X1  _1468_
timestamp 1727136778
transform 1 0 4410 0 1 17970
box -36 -24 336 816
use NAND2X1  _1469_
timestamp 1727136778
transform -1 0 3630 0 -1 16410
box -36 -24 276 816
use NAND3X1  _1470_
timestamp 1727136778
transform -1 0 2970 0 1 14850
box -36 -24 336 816
use AOI21X1  _1471_
timestamp 1727136778
transform 1 0 2430 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1472_
timestamp 1727136778
transform 1 0 2910 0 -1 16410
box -36 -24 336 816
use NAND3X1  _1473_
timestamp 1727136778
transform 1 0 3750 0 -1 16410
box -36 -24 336 816
use NAND2X1  _1474_
timestamp 1727136778
transform 1 0 8430 0 -1 10170
box -36 -24 276 816
use NOR3X1  _1475_
timestamp 1727136778
transform 1 0 8310 0 1 7050
box -36 -24 576 819
use AOI21X1  _1476_
timestamp 1727136778
transform 1 0 9030 0 1 7050
box -36 -24 336 816
use INVX1  _1477_
timestamp 1727136778
transform 1 0 9450 0 1 7050
box -36 -24 216 816
use OAI21X1  _1478_
timestamp 1727136778
transform 1 0 9810 0 1 7050
box -36 -24 336 816
use OAI21X1  _1479_
timestamp 1727136778
transform 1 0 10650 0 1 7050
box -36 -24 336 816
use NAND2X1  _1480_
timestamp 1727136778
transform -1 0 12930 0 -1 3930
box -36 -24 276 816
use NAND2X1  _1481_
timestamp 1727136778
transform -1 0 13350 0 -1 3930
box -36 -24 276 816
use NAND2X1  _1482_
timestamp 1727136778
transform 1 0 14010 0 1 2370
box -36 -24 276 816
use NAND2X1  _1483_
timestamp 1727136778
transform 1 0 16170 0 1 2370
box -36 -24 276 816
use OAI21X1  _1484_
timestamp 1727136778
transform -1 0 16890 0 1 2370
box -36 -24 336 816
use AOI21X1  _1485_
timestamp 1727136778
transform 1 0 16590 0 -1 2370
box -36 -24 336 816
use AOI22X1  _1486_
timestamp 1727136778
transform -1 0 17370 0 -1 2370
box -42 -24 396 816
use INVX1  _1487_
timestamp 1727136778
transform 1 0 17550 0 -1 2370
box -36 -24 216 816
use OAI21X1  _1488_
timestamp 1727136778
transform 1 0 6630 0 -1 17970
box -36 -24 336 816
use INVX1  _1489_
timestamp 1727136778
transform 1 0 7050 0 -1 17970
box -36 -24 216 816
use INVX1  _1490_
timestamp 1727136778
transform -1 0 7290 0 1 14850
box -36 -24 216 816
use NAND2X1  _1491_
timestamp 1727136778
transform -1 0 8910 0 1 16410
box -36 -24 276 816
use OAI21X1  _1492_
timestamp 1727136778
transform -1 0 6630 0 1 16410
box -36 -24 336 816
use OAI21X1  _1493_
timestamp 1727136778
transform -1 0 7110 0 1 16410
box -36 -24 336 816
use OR2X2  _1494_
timestamp 1727136778
transform 1 0 7770 0 1 16410
box -36 -24 336 816
use INVX1  _1495_
timestamp 1727136778
transform 1 0 8970 0 -1 16410
box -36 -24 216 816
use OAI21X1  _1496_
timestamp 1727136778
transform 1 0 7290 0 1 16410
box -36 -24 336 816
use NAND2X1  _1497_
timestamp 1727136778
transform 1 0 7890 0 -1 16410
box -36 -24 276 816
use OAI21X1  _1498_
timestamp 1727136778
transform 1 0 8250 0 -1 16410
box -36 -24 336 816
use INVX1  _1499_
timestamp 1727136778
transform 1 0 6750 0 1 14850
box -36 -24 216 816
use NAND3X1  _1500_
timestamp 1727136778
transform 1 0 7410 0 -1 16410
box -36 -24 336 816
use NAND2X1  _1501_
timestamp 1727136778
transform 1 0 8250 0 1 16410
box -36 -24 276 816
use NOR2X1  _1502_
timestamp 1727136778
transform 1 0 8250 0 -1 17970
box -36 -24 276 816
use NAND2X1  _1503_
timestamp 1727136778
transform 1 0 8430 0 1 17970
box -36 -24 276 816
use INVX1  _1504_
timestamp 1727136778
transform 1 0 8670 0 -1 17970
box -36 -24 216 816
use OAI21X1  _1505_
timestamp 1727136778
transform -1 0 7650 0 -1 17970
box -36 -24 336 816
use OR2X2  _1506_
timestamp 1727136778
transform -1 0 8250 0 1 17970
box -36 -24 336 816
use NAND3X1  _1507_
timestamp 1727136778
transform -1 0 7770 0 1 17970
box -36 -24 336 816
use NAND2X1  _1508_
timestamp 1727136778
transform -1 0 6870 0 1 17970
box -36 -24 276 816
use NAND3X1  _1509_
timestamp 1727136778
transform 1 0 6210 0 1 17970
box -36 -24 336 816
use NAND2X1  _1510_
timestamp 1727136778
transform -1 0 6030 0 1 17970
box -36 -24 276 816
use NAND3X1  _1511_
timestamp 1727136778
transform 1 0 6990 0 1 17970
box -36 -24 336 816
use NAND2X1  _1512_
timestamp 1727136778
transform -1 0 8430 0 1 10170
box -36 -24 276 816
use NOR2X1  _1513_
timestamp 1727136778
transform 1 0 10050 0 1 8610
box -36 -24 276 816
use NOR2X1  _1514_
timestamp 1727136778
transform -1 0 9390 0 1 8610
box -36 -24 276 816
use NAND3X1  _1515_
timestamp 1727136778
transform 1 0 9570 0 1 8610
box -36 -24 336 816
use NAND2X1  _1516_
timestamp 1727136778
transform -1 0 7890 0 -1 10170
box -36 -24 276 816
use AOI22X1  _1517_
timestamp 1727136778
transform 1 0 8670 0 1 8610
box -42 -24 396 816
use AOI21X1  _1518_
timestamp 1727136778
transform -1 0 9990 0 -1 10170
box -36 -24 336 816
use NAND2X1  _1519_
timestamp 1727136778
transform 1 0 8850 0 -1 10170
box -36 -24 276 816
use OAI21X1  _1520_
timestamp 1727136778
transform 1 0 9210 0 -1 10170
box -36 -24 336 816
use AOI21X1  _1521_
timestamp 1727136778
transform 1 0 7770 0 1 8610
box -36 -24 336 816
use OAI21X1  _1522_
timestamp 1727136778
transform 1 0 8250 0 1 8610
box -36 -24 336 816
use AOI22X1  _1523_
timestamp 1727136778
transform 1 0 8610 0 1 10170
box -42 -24 396 816
use OAI21X1  _1524_
timestamp 1727136778
transform 1 0 9930 0 1 10170
box -36 -24 336 816
use OR2X2  _1525_
timestamp 1727136778
transform -1 0 16770 0 1 8610
box -36 -24 336 816
use NAND3X1  _1526_
timestamp 1727136778
transform -1 0 15270 0 1 7050
box -36 -24 336 816
use INVX1  _1527_
timestamp 1727136778
transform 1 0 13470 0 -1 2370
box -36 -24 216 816
use OAI21X1  _1528_
timestamp 1727136778
transform 1 0 13050 0 -1 2370
box -36 -24 336 816
use NAND2X1  _1529_
timestamp 1727136778
transform 1 0 13830 0 -1 2370
box -36 -24 276 816
use NAND2X1  _1530_
timestamp 1727136778
transform -1 0 14790 0 1 7050
box -36 -24 276 816
use OAI21X1  _1531_
timestamp 1727136778
transform -1 0 15570 0 1 2370
box -36 -24 336 816
use AOI21X1  _1532_
timestamp 1727136778
transform 1 0 15750 0 1 2370
box -36 -24 336 816
use AOI22X1  _1533_
timestamp 1727136778
transform -1 0 16410 0 -1 2370
box -42 -24 396 816
use INVX1  _1534_
timestamp 1727136778
transform -1 0 15690 0 1 810
box -36 -24 216 816
use INVX1  _1535_
timestamp 1727136778
transform -1 0 11490 0 -1 8610
box -36 -24 216 816
use NAND2X1  _1536_
timestamp 1727136778
transform 1 0 9570 0 1 10170
box -36 -24 276 816
use INVX1  _1537_
timestamp 1727136778
transform 1 0 8490 0 1 11730
box -36 -24 216 816
use AOI21X1  _1538_
timestamp 1727136778
transform 1 0 7830 0 -1 17970
box -36 -24 336 816
use OAI21X1  _1539_
timestamp 1727136778
transform 1 0 6930 0 -1 16410
box -36 -24 336 816
use NOR2X1  _1540_
timestamp 1727136778
transform -1 0 8190 0 1 14850
box -36 -24 276 816
use NAND3X1  _1541_
timestamp 1727136778
transform -1 0 8730 0 -1 14850
box -36 -24 336 816
use OAI22X1  _1542_
timestamp 1727136778
transform -1 0 7770 0 1 14850
box -36 -24 396 816
use NAND2X1  _1543_
timestamp 1727136778
transform 1 0 8010 0 -1 14850
box -36 -24 276 816
use XNOR2X1  _1544_
timestamp 1727153789
transform 1 0 7410 0 -1 14850
box -36 -24 456 816
use XOR2X1  _1545_
timestamp 1727152697
transform -1 0 7830 0 1 13290
box -36 -24 453 816
use XOR2X1  _1546_
timestamp 1727152697
transform -1 0 7950 0 -1 13290
box -36 -24 453 816
use NOR2X1  _1547_
timestamp 1727136778
transform -1 0 8310 0 -1 11730
box -36 -24 276 816
use OAI21X1  _1548_
timestamp 1727136778
transform -1 0 9450 0 1 10170
box -36 -24 336 816
use OAI21X1  _1549_
timestamp 1727136778
transform -1 0 8730 0 -1 11730
box -36 -24 336 816
use NAND3X1  _1550_
timestamp 1727136778
transform 1 0 10470 0 1 8610
box -36 -24 336 816
use AOI21X1  _1551_
timestamp 1727136778
transform 1 0 11790 0 1 810
box -36 -24 336 816
use OAI21X1  _1552_
timestamp 1727136778
transform 1 0 12570 0 1 810
box -36 -24 336 816
use INVX1  _1553_
timestamp 1727136778
transform -1 0 15390 0 1 5490
box -36 -24 216 816
use AOI21X1  _1554_
timestamp 1727136778
transform 1 0 15750 0 -1 3930
box -36 -24 336 816
use AOI21X1  _1555_
timestamp 1727136778
transform 1 0 15630 0 -1 2370
box -36 -24 336 816
use AOI22X1  _1556_
timestamp 1727136778
transform -1 0 15330 0 1 810
box -42 -24 396 816
use INVX1  _1557_
timestamp 1727136778
transform -1 0 14790 0 1 810
box -36 -24 216 816
use NAND3X1  _1558_
timestamp 1727136778
transform 1 0 7590 0 -1 11730
box -36 -24 336 816
use INVX1  _1559_
timestamp 1727136778
transform 1 0 10650 0 -1 10170
box -36 -24 216 816
use NAND3X1  _1560_
timestamp 1727136778
transform 1 0 11010 0 -1 10170
box -36 -24 336 816
use NAND2X1  _1561_
timestamp 1727136778
transform -1 0 8310 0 1 11730
box -36 -24 276 816
use OAI21X1  _1562_
timestamp 1727136778
transform 1 0 8130 0 -1 13290
box -36 -24 336 816
use INVX1  _1563_
timestamp 1727136778
transform 1 0 11190 0 1 10170
box -36 -24 216 816
use INVX1  _1564_
timestamp 1727136778
transform -1 0 6330 0 -1 14850
box -36 -24 216 816
use NAND2X1  _1565_
timestamp 1727136778
transform -1 0 6750 0 -1 14850
box -36 -24 276 816
use OAI21X1  _1566_
timestamp 1727136778
transform -1 0 7230 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1567_
timestamp 1727136778
transform 1 0 8730 0 1 13290
box -36 -24 336 816
use XOR2X1  _1568_
timestamp 1727152697
transform 1 0 10050 0 1 13290
box -36 -24 453 816
use NAND3X1  _1569_
timestamp 1727136778
transform 1 0 11910 0 -1 10170
box -36 -24 336 816
use AOI21X1  _1570_
timestamp 1727136778
transform 1 0 10170 0 -1 10170
box -36 -24 336 816
use INVX1  _1571_
timestamp 1727136778
transform -1 0 11010 0 1 10170
box -36 -24 216 816
use OAI21X1  _1572_
timestamp 1727136778
transform 1 0 10410 0 1 10170
box -36 -24 336 816
use NAND3X1  _1573_
timestamp 1727136778
transform 1 0 12390 0 -1 10170
box -36 -24 336 816
use NAND2X1  _1574_
timestamp 1727136778
transform -1 0 12390 0 -1 810
box -36 -24 276 816
use NOR2X1  _1575_
timestamp 1727136778
transform 1 0 13050 0 -1 810
box -36 -24 276 816
use AOI21X1  _1576_
timestamp 1727136778
transform 1 0 12570 0 -1 810
box -36 -24 336 816
use OAI21X1  _1577_
timestamp 1727136778
transform 1 0 13410 0 -1 810
box -36 -24 336 816
use NOR2X1  _1578_
timestamp 1727136778
transform 1 0 17190 0 -1 10170
box -36 -24 276 816
use NOR2X1  _1579_
timestamp 1727136778
transform -1 0 15630 0 -1 7050
box -36 -24 276 816
use AOI21X1  _1580_
timestamp 1727136778
transform -1 0 15510 0 -1 2370
box -36 -24 336 816
use AOI22X1  _1581_
timestamp 1727136778
transform 1 0 14730 0 -1 2370
box -42 -24 396 816
use INVX1  _1582_
timestamp 1727136778
transform -1 0 13710 0 1 810
box -36 -24 216 816
use AOI21X1  _1583_
timestamp 1727136778
transform -1 0 11730 0 -1 10170
box -36 -24 336 816
use NAND3X1  _1584_
timestamp 1727136778
transform 1 0 8910 0 -1 14850
box -36 -24 336 816
use NAND2X1  _1585_
timestamp 1727136778
transform 1 0 9390 0 -1 14850
box -36 -24 276 816
use OAI21X1  _1586_
timestamp 1727136778
transform 1 0 10890 0 1 8610
box -36 -24 336 816
use NAND2X1  _1587_
timestamp 1727136778
transform 1 0 7710 0 -1 810
box -36 -24 276 816
use XNOR2X1  _1588_
timestamp 1727153789
transform -1 0 12030 0 -1 810
box -36 -24 456 816
use NAND2X1  _1589_
timestamp 1727136778
transform 1 0 14850 0 1 2370
box -36 -24 276 816
use OAI21X1  _1590_
timestamp 1727136778
transform 1 0 14430 0 1 2370
box -36 -24 336 816
use AOI21X1  _1591_
timestamp 1727136778
transform -1 0 14550 0 -1 2370
box -36 -24 336 816
use AOI22X1  _1592_
timestamp 1727136778
transform -1 0 13350 0 1 810
box -42 -24 396 816
use NAND2X1  _1593_
timestamp 1727136778
transform -1 0 13290 0 -1 8610
box -36 -24 276 816
use OAI21X1  _1594_
timestamp 1727136778
transform 1 0 12990 0 1 8610
box -36 -24 336 816
use NAND2X1  _1595_
timestamp 1727136778
transform 1 0 12030 0 1 11730
box -36 -24 276 816
use OAI21X1  _1596_
timestamp 1727136778
transform -1 0 12690 0 1 11730
box -36 -24 336 816
use NAND2X1  _1597_
timestamp 1727136778
transform 1 0 12090 0 1 8610
box -36 -24 276 816
use OAI21X1  _1598_
timestamp 1727136778
transform -1 0 12810 0 1 8610
box -36 -24 336 816
use NAND2X1  _1599_
timestamp 1727136778
transform -1 0 11910 0 -1 11730
box -36 -24 276 816
use OAI21X1  _1600_
timestamp 1727136778
transform -1 0 12390 0 -1 11730
box -36 -24 336 816
use NAND2X1  _1601_
timestamp 1727136778
transform 1 0 9990 0 1 11730
box -36 -24 276 816
use OAI21X1  _1602_
timestamp 1727136778
transform -1 0 10290 0 -1 13290
box -36 -24 336 816
use NAND2X1  _1603_
timestamp 1727136778
transform 1 0 8910 0 -1 11730
box -36 -24 276 816
use OAI21X1  _1604_
timestamp 1727136778
transform -1 0 9630 0 -1 11730
box -36 -24 336 816
use NAND2X1  _1605_
timestamp 1727136778
transform -1 0 13650 0 1 10170
box -36 -24 276 816
use OAI21X1  _1606_
timestamp 1727136778
transform -1 0 15810 0 -1 10170
box -36 -24 336 816
use NAND2X1  _1607_
timestamp 1727136778
transform 1 0 13350 0 1 7050
box -36 -24 276 816
use OAI21X1  _1608_
timestamp 1727136778
transform -1 0 14010 0 1 7050
box -36 -24 336 816
use DFFPOSX1  _1609_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726828622
transform -1 0 14370 0 1 10170
box -39 -24 759 816
use DFFPOSX1  _1610_
timestamp 1726828622
transform -1 0 10950 0 1 11730
box -39 -24 759 816
use DFFPOSX1  _1611_
timestamp 1726828622
transform -1 0 14730 0 1 8610
box -39 -24 759 816
use DFFPOSX1  _1612_
timestamp 1726828622
transform -1 0 11850 0 -1 13290
box -39 -24 759 816
use DFFPOSX1  _1613_
timestamp 1726828622
transform -1 0 9870 0 -1 13290
box -39 -24 759 816
use DFFPOSX1  _1614_
timestamp 1726828622
transform -1 0 10350 0 -1 11730
box -39 -24 759 816
use DFFPOSX1  _1615_
timestamp 1726828622
transform -1 0 15810 0 1 10170
box -39 -24 759 816
use DFFPOSX1  _1616_
timestamp 1726828622
transform 1 0 14490 0 -1 8610
box -39 -24 759 816
use DFFPOSX1  _1617_
timestamp 1726828622
transform -1 0 15210 0 -1 5490
box -39 -24 759 816
use DFFPOSX1  _1618_
timestamp 1726828622
transform -1 0 11610 0 -1 7050
box -39 -24 759 816
use DFFPOSX1  _1619_
timestamp 1726828622
transform -1 0 14790 0 -1 3930
box -39 -24 759 816
use DFFPOSX1  _1620_
timestamp 1726828622
transform 1 0 16410 0 1 810
box -39 -24 759 816
use DFFPOSX1  _1621_
timestamp 1726828622
transform -1 0 16410 0 1 810
box -39 -24 759 816
use DFFPOSX1  _1622_
timestamp 1726828622
transform 1 0 15270 0 -1 810
box -39 -24 759 816
use DFFPOSX1  _1623_
timestamp 1726828622
transform 1 0 14130 0 -1 810
box -39 -24 759 816
use DFFPOSX1  _1624_
timestamp 1726828622
transform -1 0 14430 0 1 810
box -39 -24 759 816
use DFFPOSX1  _1625_
timestamp 1726828622
transform -1 0 14010 0 1 8610
box -39 -24 759 816
use DFFPOSX1  _1626_
timestamp 1726828622
transform -1 0 13110 0 -1 11730
box -39 -24 759 816
use DFFPOSX1  _1627_
timestamp 1726828622
transform -1 0 11910 0 1 8610
box -39 -24 759 816
use DFFPOSX1  _1628_
timestamp 1726828622
transform -1 0 12510 0 1 10170
box -39 -24 759 816
use DFFPOSX1  _1629_
timestamp 1726828622
transform -1 0 9150 0 -1 13290
box -39 -24 759 816
use DFFPOSX1  _1630_
timestamp 1726828622
transform -1 0 9810 0 1 11730
box -39 -24 759 816
use DFFPOSX1  _1631_
timestamp 1726828622
transform -1 0 15090 0 1 10170
box -39 -24 759 816
use DFFPOSX1  _1632_
timestamp 1726828622
transform -1 0 14130 0 -1 7050
box -39 -24 759 816
use DFFSR  _1633_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727133863
transform -1 0 17790 0 1 3930
box -36 -24 1476 819
use DFFSR  _1634_
timestamp 1727133863
transform -1 0 18210 0 -1 3930
box -36 -24 1476 819
use DFFSR  _1635_
timestamp 1727133863
transform -1 0 18150 0 -1 5490
box -36 -24 1476 819
use INVX1  _1636_
timestamp 1727136778
transform -1 0 17910 0 -1 16410
box -36 -24 216 816
use INVX4  _1637_
timestamp 1727136778
transform 1 0 17790 0 1 17970
box -36 -24 276 816
use OAI21X1  _1638_
timestamp 1727136778
transform -1 0 16350 0 -1 16410
box -36 -24 336 816
use NOR2X1  _1639_
timestamp 1727136778
transform 1 0 15690 0 -1 16410
box -36 -24 276 816
use INVX1  _1640_
timestamp 1727136778
transform 1 0 15690 0 1 16410
box -36 -24 216 816
use INVX2  _1641_
timestamp 1727136778
transform -1 0 11430 0 1 16410
box -36 -24 216 816
use NAND2X1  _1642_
timestamp 1727136778
transform -1 0 9750 0 1 16410
box -36 -24 276 816
use INVX2  _1643_
timestamp 1727136778
transform -1 0 9210 0 -1 17970
box -36 -24 216 816
use NAND2X1  _1644_
timestamp 1727136778
transform -1 0 11850 0 1 16410
box -36 -24 276 816
use NAND2X1  _1645_
timestamp 1727136778
transform -1 0 13410 0 -1 16410
box -36 -24 276 816
use AOI22X1  _1646_
timestamp 1727136778
transform -1 0 12690 0 -1 16410
box -42 -24 396 816
use INVX2  _1647_
timestamp 1727136778
transform 1 0 9570 0 1 17970
box -36 -24 216 816
use INVX1  _1648_
timestamp 1727136778
transform 1 0 17370 0 -1 16410
box -36 -24 216 816
use INVX1  _1649_
timestamp 1727136778
transform -1 0 13050 0 -1 16410
box -36 -24 216 816
use OAI21X1  _1650_
timestamp 1727136778
transform -1 0 13650 0 1 16410
box -36 -24 336 816
use NAND2X1  _1651_
timestamp 1727136778
transform 1 0 12930 0 1 16410
box -36 -24 276 816
use NAND2X1  _1652_
timestamp 1727136778
transform -1 0 11130 0 1 16410
box -36 -24 276 816
use OAI21X1  _1653_
timestamp 1727136778
transform 1 0 12510 0 1 16410
box -36 -24 336 816
use OAI21X1  _1654_
timestamp 1727136778
transform 1 0 17430 0 1 16410
box -36 -24 336 816
use AOI21X1  _1655_
timestamp 1727136778
transform -1 0 17310 0 1 16410
box -36 -24 336 816
use NOR2X1  _1656_
timestamp 1727136778
transform 1 0 17850 0 -1 17970
box -36 -24 276 816
use OAI21X1  _1657_
timestamp 1727136778
transform 1 0 17370 0 -1 17970
box -36 -24 336 816
use OAI21X1  _1658_
timestamp 1727136778
transform 1 0 16950 0 -1 17970
box -36 -24 336 816
use XOR2X1  _1659_
timestamp 1727152697
transform -1 0 16470 0 1 16410
box -36 -24 453 816
use NOR2X1  _1660_
timestamp 1727136778
transform -1 0 16770 0 -1 17970
box -36 -24 276 816
use OAI21X1  _1661_
timestamp 1727136778
transform 1 0 16110 0 -1 17970
box -36 -24 336 816
use NAND2X1  _1662_
timestamp 1727136778
transform -1 0 10650 0 1 17970
box -36 -24 276 816
use NAND3X1  _1663_
timestamp 1727136778
transform -1 0 10170 0 1 16410
box -36 -24 336 816
use AOI22X1  _1664_
timestamp 1727136778
transform -1 0 10710 0 1 16410
box -42 -24 396 816
use INVX1  _1665_
timestamp 1727136778
transform -1 0 11130 0 -1 13290
box -36 -24 216 816
use NOR2X1  _1666_
timestamp 1727136778
transform -1 0 11730 0 1 13290
box -36 -24 276 816
use OAI21X1  _1667_
timestamp 1727136778
transform 1 0 11550 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1668_
timestamp 1727136778
transform 1 0 11190 0 -1 17970
box -36 -24 336 816
use OAI21X1  _1669_
timestamp 1727136778
transform -1 0 12450 0 -1 17970
box -36 -24 336 816
use AOI21X1  _1670_
timestamp 1727136778
transform 1 0 12570 0 -1 17970
box -36 -24 336 816
use INVX1  _1671_
timestamp 1727136778
transform 1 0 15750 0 1 17970
box -36 -24 216 816
use OAI21X1  _1672_
timestamp 1727136778
transform -1 0 17310 0 1 17970
box -36 -24 336 816
use MUX2X1  _1673_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 16470 0 1 17970
box -36 -24 393 816
use NAND2X1  _1674_
timestamp 1727136778
transform -1 0 16350 0 1 17970
box -36 -24 276 816
use INVX1  _1675_
timestamp 1727136778
transform -1 0 16830 0 1 16410
box -36 -24 216 816
use OAI21X1  _1676_
timestamp 1727136778
transform 1 0 16470 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1677_
timestamp 1727136778
transform -1 0 14970 0 1 16410
box -36 -24 336 816
use MUX2X1  _1678_
timestamp 1727136778
transform -1 0 15150 0 -1 16410
box -36 -24 393 816
use NAND2X1  _1679_
timestamp 1727136778
transform -1 0 13770 0 -1 16410
box -36 -24 276 816
use NAND2X1  _1680_
timestamp 1727136778
transform 1 0 13950 0 -1 16410
box -36 -24 276 816
use AOI21X1  _1681_
timestamp 1727136778
transform -1 0 12330 0 1 16410
box -36 -24 336 816
use NAND2X1  _1682_
timestamp 1727136778
transform 1 0 13770 0 1 16410
box -36 -24 276 816
use NAND3X1  _1683_
timestamp 1727136778
transform 1 0 14190 0 1 16410
box -36 -24 336 816
use AOI22X1  _1684_
timestamp 1727136778
transform 1 0 15150 0 1 16410
box -42 -24 396 816
use OAI21X1  _1685_
timestamp 1727136778
transform -1 0 12810 0 1 17970
box -36 -24 336 816
use OAI21X1  _1686_
timestamp 1727136778
transform 1 0 12990 0 1 17970
box -36 -24 336 816
use NAND2X1  _1687_
timestamp 1727136778
transform -1 0 15570 0 -1 17970
box -36 -24 276 816
use NAND2X1  _1688_
timestamp 1727136778
transform 1 0 15690 0 -1 17970
box -36 -24 276 816
use INVX1  _1689_
timestamp 1727136778
transform 1 0 14730 0 -1 7050
box -36 -24 216 816
use NOR2X1  _1690_
timestamp 1727136778
transform 1 0 15330 0 1 17970
box -36 -24 276 816
use OAI21X1  _1691_
timestamp 1727136778
transform -1 0 15150 0 1 17970
box -36 -24 336 816
use NAND2X1  _1692_
timestamp 1727136778
transform 1 0 10770 0 -1 17970
box -36 -24 276 816
use NAND3X1  _1693_
timestamp 1727136778
transform 1 0 9390 0 -1 17970
box -36 -24 336 816
use AOI22X1  _1694_
timestamp 1727136778
transform -1 0 10230 0 -1 17970
box -42 -24 396 816
use INVX1  _1695_
timestamp 1727136778
transform -1 0 8970 0 1 17970
box -36 -24 216 816
use NOR2X1  _1696_
timestamp 1727136778
transform -1 0 9390 0 1 17970
box -36 -24 276 816
use OAI21X1  _1697_
timestamp 1727136778
transform -1 0 10230 0 1 17970
box -36 -24 336 816
use OAI21X1  _1698_
timestamp 1727136778
transform 1 0 10350 0 -1 17970
box -36 -24 336 816
use OAI21X1  _1699_
timestamp 1727136778
transform -1 0 11970 0 -1 17970
box -36 -24 336 816
use AOI21X1  _1700_
timestamp 1727136778
transform -1 0 12030 0 1 17970
box -36 -24 336 816
use OAI21X1  _1701_
timestamp 1727136778
transform -1 0 11070 0 1 17970
box -36 -24 336 816
use OAI21X1  _1702_
timestamp 1727136778
transform 1 0 11250 0 1 17970
box -36 -24 336 816
use XOR2X1  _1703_
timestamp 1727152697
transform -1 0 14190 0 1 17970
box -36 -24 453 816
use INVX1  _1704_
timestamp 1727136778
transform -1 0 14550 0 -1 11730
box -36 -24 216 816
use INVX1  _1705_
timestamp 1727136778
transform 1 0 12210 0 1 17970
box -36 -24 216 816
use OAI21X1  _1706_
timestamp 1727136778
transform -1 0 13350 0 -1 17970
box -36 -24 336 816
use INVX1  _1707_
timestamp 1727136778
transform -1 0 13590 0 1 17970
box -36 -24 216 816
use AOI22X1  _1708_
timestamp 1727136778
transform 1 0 13530 0 -1 17970
box -42 -24 396 816
use NAND2X1  _1709_
timestamp 1727136778
transform -1 0 11250 0 -1 14850
box -36 -24 276 816
use AND2X2  _1710_
timestamp 1727136778
transform -1 0 11910 0 1 14850
box -36 -24 336 819
use NAND2X1  _1711_
timestamp 1727136778
transform -1 0 10950 0 1 14850
box -36 -24 276 816
use AOI22X1  _1712_
timestamp 1727136778
transform -1 0 11490 0 1 14850
box -42 -24 396 816
use OAI21X1  _1713_
timestamp 1727136778
transform -1 0 10530 0 1 14850
box -36 -24 336 816
use OAI21X1  _1714_
timestamp 1727136778
transform 1 0 11370 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1715_
timestamp 1727136778
transform -1 0 12150 0 -1 14850
box -36 -24 336 816
use AOI21X1  _1716_
timestamp 1727136778
transform 1 0 12330 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1717_
timestamp 1727136778
transform -1 0 13590 0 1 13290
box -36 -24 336 816
use OAI21X1  _1718_
timestamp 1727136778
transform 1 0 13770 0 1 13290
box -36 -24 336 816
use XOR2X1  _1719_
timestamp 1727152697
transform 1 0 14250 0 1 13290
box -36 -24 453 816
use XNOR2X1  _1720_
timestamp 1727153789
transform 1 0 12750 0 -1 13290
box -36 -24 456 816
use NAND2X1  _1721_
timestamp 1727136778
transform 1 0 14070 0 -1 17970
box -36 -24 276 816
use NAND3X1  _1722_
timestamp 1727136778
transform 1 0 14370 0 1 17970
box -36 -24 336 816
use NAND3X1  _1723_
timestamp 1727136778
transform 1 0 14430 0 -1 17970
box -36 -24 336 816
use NAND2X1  _1724_
timestamp 1727136778
transform -1 0 14670 0 1 11730
box -36 -24 276 816
use OAI21X1  _1725_
timestamp 1727136778
transform 1 0 13350 0 -1 13290
box -36 -24 336 816
use INVX1  _1726_
timestamp 1727136778
transform -1 0 12990 0 1 11730
box -36 -24 216 816
use OAI21X1  _1727_
timestamp 1727136778
transform -1 0 13470 0 1 11730
box -36 -24 336 816
use NAND2X1  _1728_
timestamp 1727136778
transform -1 0 9330 0 1 16410
box -36 -24 276 816
use AND2X2  _1729_
timestamp 1727136778
transform 1 0 9270 0 -1 16410
box -36 -24 336 819
use NAND2X1  _1730_
timestamp 1727136778
transform -1 0 9990 0 -1 16410
box -36 -24 276 816
use AOI22X1  _1731_
timestamp 1727136778
transform -1 0 10530 0 -1 16410
box -42 -24 396 816
use OAI21X1  _1732_
timestamp 1727136778
transform 1 0 10650 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1733_
timestamp 1727136778
transform 1 0 11130 0 -1 16410
box -36 -24 336 816
use OAI21X1  _1734_
timestamp 1727136778
transform 1 0 14970 0 -1 14850
box -36 -24 336 816
use AOI21X1  _1735_
timestamp 1727136778
transform 1 0 14790 0 1 13290
box -36 -24 336 816
use OAI21X1  _1736_
timestamp 1727136778
transform -1 0 16050 0 1 13290
box -36 -24 336 816
use OAI21X1  _1737_
timestamp 1727136778
transform 1 0 15270 0 1 13290
box -36 -24 336 816
use INVX1  _1738_
timestamp 1727136778
transform 1 0 15390 0 1 11730
box -36 -24 216 816
use XOR2X1  _1739_
timestamp 1727152697
transform 1 0 14790 0 1 11730
box -36 -24 453 816
use INVX1  _1740_
timestamp 1727136778
transform -1 0 15690 0 -1 13290
box -36 -24 216 816
use AOI21X1  _1741_
timestamp 1727136778
transform 1 0 15750 0 1 11730
box -36 -24 336 816
use NAND2X1  _1742_
timestamp 1727136778
transform 1 0 10590 0 -1 14850
box -36 -24 276 816
use AND2X2  _1743_
timestamp 1727136778
transform -1 0 8670 0 1 14850
box -36 -24 336 819
use NAND2X1  _1744_
timestamp 1727136778
transform -1 0 9090 0 1 14850
box -36 -24 276 816
use AOI22X1  _1745_
timestamp 1727136778
transform -1 0 10050 0 1 14850
box -42 -24 396 816
use OAI21X1  _1746_
timestamp 1727136778
transform 1 0 9270 0 1 14850
box -36 -24 336 816
use OAI21X1  _1747_
timestamp 1727136778
transform 1 0 10170 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1748_
timestamp 1727136778
transform -1 0 15570 0 1 14850
box -36 -24 336 816
use AOI21X1  _1749_
timestamp 1727136778
transform 1 0 15750 0 1 14850
box -36 -24 336 816
use OAI21X1  _1750_
timestamp 1727136778
transform 1 0 16410 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1751_
timestamp 1727136778
transform 1 0 16170 0 1 13290
box -36 -24 336 816
use INVX1  _1752_
timestamp 1727136778
transform -1 0 16050 0 -1 13290
box -36 -24 216 816
use XOR2X1  _1753_
timestamp 1727152697
transform 1 0 16230 0 1 11730
box -36 -24 453 816
use INVX1  _1754_
timestamp 1727136778
transform 1 0 15510 0 1 5490
box -36 -24 216 816
use OAI21X1  _1755_
timestamp 1727136778
transform 1 0 16230 0 -1 13290
box -36 -24 336 816
use INVX1  _1756_
timestamp 1727136778
transform 1 0 14610 0 -1 14850
box -36 -24 216 816
use AND2X2  _1757_
timestamp 1727136778
transform -1 0 13470 0 -1 14850
box -36 -24 336 819
use NAND2X1  _1758_
timestamp 1727136778
transform 1 0 12810 0 -1 14850
box -36 -24 276 816
use AOI22X1  _1759_
timestamp 1727136778
transform 1 0 12090 0 1 14850
box -42 -24 396 816
use OAI21X1  _1760_
timestamp 1727136778
transform 1 0 13650 0 -1 14850
box -36 -24 336 816
use OAI22X1  _1761_
timestamp 1727136778
transform -1 0 14430 0 -1 14850
box -36 -24 396 816
use OAI21X1  _1762_
timestamp 1727136778
transform -1 0 15750 0 -1 14850
box -36 -24 336 816
use AOI21X1  _1763_
timestamp 1727136778
transform 1 0 15930 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1764_
timestamp 1727136778
transform 1 0 16830 0 -1 14850
box -36 -24 336 816
use OAI21X1  _1765_
timestamp 1727136778
transform 1 0 17310 0 -1 14850
box -36 -24 336 816
use NAND2X1  _1766_
timestamp 1727136778
transform 1 0 17610 0 -1 11730
box -36 -24 276 816
use INVX1  _1767_
timestamp 1727136778
transform 1 0 14730 0 -1 13290
box -36 -24 216 816
use AOI21X1  _1768_
timestamp 1727136778
transform -1 0 14610 0 -1 13290
box -36 -24 336 816
use AOI21X1  _1769_
timestamp 1727136778
transform -1 0 14130 0 -1 13290
box -36 -24 336 816
use OAI21X1  _1770_
timestamp 1727136778
transform -1 0 15330 0 -1 13290
box -36 -24 336 816
use OR2X2  _1771_
timestamp 1727136778
transform 1 0 16650 0 1 13290
box -36 -24 336 816
use AOI22X1  _1772_
timestamp 1727136778
transform 1 0 16710 0 -1 13290
box -42 -24 396 816
use INVX1  _1773_
timestamp 1727136778
transform -1 0 17610 0 1 17970
box -36 -24 216 816
use NAND2X1  _1774_
timestamp 1727136778
transform -1 0 17070 0 1 11730
box -36 -24 276 816
use NAND2X1  _1775_
timestamp 1727136778
transform -1 0 17430 0 -1 11730
box -36 -24 276 816
use OAI21X1  _1776_
timestamp 1727136778
transform 1 0 17190 0 -1 13290
box -36 -24 336 816
use NAND2X1  _1777_
timestamp 1727136778
transform 1 0 14910 0 1 14850
box -36 -24 276 816
use AND2X2  _1778_
timestamp 1727136778
transform 1 0 13530 0 1 14850
box -36 -24 336 819
use NAND2X1  _1779_
timestamp 1727136778
transform 1 0 13110 0 1 14850
box -36 -24 276 816
use AOI22X1  _1780_
timestamp 1727136778
transform 1 0 12630 0 1 14850
box -42 -24 396 816
use OAI21X1  _1781_
timestamp 1727136778
transform 1 0 14010 0 1 14850
box -36 -24 336 816
use OAI21X1  _1782_
timestamp 1727136778
transform 1 0 14430 0 1 14850
box -36 -24 336 816
use OAI21X1  _1783_
timestamp 1727136778
transform 1 0 16950 0 -1 16410
box -36 -24 336 816
use AOI21X1  _1784_
timestamp 1727136778
transform 1 0 16530 0 1 14850
box -36 -24 336 816
use OAI21X1  _1785_
timestamp 1727136778
transform -1 0 17790 0 1 14850
box -36 -24 336 816
use OAI21X1  _1786_
timestamp 1727136778
transform 1 0 17910 0 1 14850
box -36 -24 336 816
use NAND2X1  _1787_
timestamp 1727136778
transform -1 0 17970 0 -1 810
box -36 -24 276 816
use NAND2X1  _1788_
timestamp 1727136778
transform 1 0 17250 0 1 11730
box -36 -24 276 816
use INVX1  _1789_
timestamp 1727136778
transform 1 0 18030 0 -1 13290
box -36 -24 216 816
use NAND3X1  _1790_
timestamp 1727136778
transform 1 0 18090 0 1 11730
box -36 -24 336 816
use NAND2X1  _1791_
timestamp 1727136778
transform 1 0 18030 0 1 7050
box -36 -24 276 816
use NOR2X1  _1792_
timestamp 1727136778
transform 1 0 14010 0 1 11730
box -36 -24 276 816
use NAND2X1  _1793_
timestamp 1727136778
transform 1 0 13650 0 1 11730
box -36 -24 276 816
use NOR2X1  _1794_
timestamp 1727136778
transform 1 0 14730 0 -1 11730
box -36 -24 276 816
use NAND3X1  _1795_
timestamp 1727136778
transform -1 0 17010 0 -1 11730
box -36 -24 336 816
use NOR2X1  _1796_
timestamp 1727136778
transform 1 0 16350 0 -1 11730
box -36 -24 276 816
use AND2X2  _1797_
timestamp 1727136778
transform -1 0 15450 0 -1 11730
box -36 -24 336 819
use NAND3X1  _1798_
timestamp 1727136778
transform -1 0 17910 0 1 11730
box -36 -24 336 816
use NAND2X1  _1799_
timestamp 1727136778
transform -1 0 17910 0 -1 13290
box -36 -24 276 816
use NAND2X1  _1800_
timestamp 1727136778
transform -1 0 17850 0 1 10170
box -36 -24 276 816
use NAND2X1  _1801_
timestamp 1727136778
transform 1 0 16290 0 1 10170
box -36 -24 276 816
use NOR2X1  _1802_
timestamp 1727136778
transform 1 0 14370 0 -1 16410
box -36 -24 276 816
use OAI21X1  _1803_
timestamp 1727136778
transform 1 0 17730 0 1 810
box -36 -24 336 816
use NOR2X1  _1804_
timestamp 1727136778
transform -1 0 17910 0 1 13290
box -36 -24 276 816
use AOI21X1  _1805_
timestamp 1727136778
transform 1 0 18090 0 1 13290
box -36 -24 336 816
use XOR2X1  _1806_
timestamp 1727152697
transform -1 0 17550 0 1 13290
box -36 -24 453 816
use OAI21X1  _1807_
timestamp 1727136778
transform 1 0 17130 0 1 10170
box -36 -24 336 816
use NAND3X1  _1808_
timestamp 1727136778
transform 1 0 16650 0 1 10170
box -36 -24 336 816
use AOI21X1  _1809_
timestamp 1727136778
transform 1 0 17010 0 1 14850
box -36 -24 336 816
use XOR2X1  _1810_
timestamp 1727152697
transform 1 0 17790 0 -1 14850
box -36 -24 453 816
use NAND3X1  _1811_
timestamp 1727136778
transform 1 0 17250 0 1 810
box -36 -24 336 816
use INVX1  _1812_
timestamp 1727136778
transform 1 0 18030 0 -1 11730
box -36 -24 216 816
use NAND3X1  _1813_
timestamp 1727136778
transform -1 0 18330 0 1 10170
box -36 -24 336 816
use NAND2X1  _1814_
timestamp 1727136778
transform -1 0 18270 0 -1 10170
box -36 -24 276 816
use NAND3X1  _1815_
timestamp 1727136778
transform 1 0 17610 0 -1 10170
box -36 -24 336 816
use NAND3X1  _1816_
timestamp 1727136778
transform -1 0 18330 0 1 8610
box -36 -24 336 816
use NAND2X1  _1817_
timestamp 1727136778
transform -1 0 17850 0 1 8610
box -36 -24 276 816
use BUFX2  _1818_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 10110 0 -1 7050
box -36 -24 276 816
use BUFX2  _1819_
timestamp 1727136778
transform -1 0 8070 0 -1 7050
box -36 -24 276 816
use BUFX2  _1820_
timestamp 1727136778
transform -1 0 14070 0 -1 3930
box -36 -24 276 816
use BUFX2  _1821_
timestamp 1727136778
transform -1 0 17190 0 -1 810
box -36 -24 276 816
use BUFX2  _1822_
timestamp 1727136778
transform 1 0 16530 0 -1 810
box -36 -24 276 816
use BUFX2  _1823_
timestamp 1727136778
transform 1 0 16110 0 -1 810
box -36 -24 276 816
use BUFX2  _1824_
timestamp 1727136778
transform 1 0 15030 0 -1 810
box -36 -24 276 816
use BUFX2  _1825_
timestamp 1727136778
transform 1 0 13890 0 -1 810
box -36 -24 276 816
use BUFX2  _1826_
timestamp 1727136778
transform 1 0 17310 0 -1 810
box -36 -24 276 816
use BUFX2  BUFX2_insert0
timestamp 1727136778
transform 1 0 11910 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert1
timestamp 1727136778
transform -1 0 6930 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert2
timestamp 1727136778
transform -1 0 7230 0 1 7050
box -36 -24 276 816
use BUFX2  BUFX2_insert3
timestamp 1727136778
transform -1 0 7110 0 -1 11730
box -36 -24 276 816
use BUFX2  BUFX2_insert4
timestamp 1727136778
transform -1 0 13530 0 -1 11730
box -36 -24 276 816
use BUFX2  BUFX2_insert5
timestamp 1727136778
transform -1 0 11550 0 -1 11730
box -36 -24 276 816
use BUFX2  BUFX2_insert6
timestamp 1727136778
transform -1 0 8490 0 -1 7050
box -36 -24 276 816
use BUFX2  BUFX2_insert7
timestamp 1727136778
transform -1 0 10530 0 -1 7050
box -36 -24 276 816
use BUFX2  BUFX2_insert13
timestamp 1727136778
transform 1 0 15690 0 1 8610
box -36 -24 276 816
use BUFX2  BUFX2_insert14
timestamp 1727136778
transform -1 0 11790 0 1 10170
box -36 -24 276 816
use BUFX2  BUFX2_insert15
timestamp 1727136778
transform -1 0 13290 0 1 10170
box -36 -24 276 816
use BUFX2  BUFX2_insert16
timestamp 1727136778
transform -1 0 12390 0 -1 8610
box -36 -24 276 816
use BUFX2  BUFX2_insert17
timestamp 1727136778
transform 1 0 7710 0 1 11730
box -36 -24 276 816
use BUFX2  BUFX2_insert18
timestamp 1727136778
transform -1 0 7290 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert19
timestamp 1727136778
transform 1 0 9210 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert20
timestamp 1727136778
transform -1 0 7590 0 1 8610
box -36 -24 276 816
use BUFX2  BUFX2_insert21
timestamp 1727136778
transform 1 0 16050 0 1 8610
box -36 -24 276 816
use BUFX2  BUFX2_insert22
timestamp 1727136778
transform -1 0 12930 0 1 10170
box -36 -24 276 816
use BUFX2  BUFX2_insert23
timestamp 1727136778
transform 1 0 12870 0 -1 10170
box -36 -24 276 816
use BUFX2  BUFX2_insert24
timestamp 1727136778
transform 1 0 15930 0 -1 10170
box -36 -24 276 816
use BUFX2  BUFX2_insert25
timestamp 1727136778
transform -1 0 7350 0 -1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert26
timestamp 1727136778
transform -1 0 8250 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert27
timestamp 1727136778
transform -1 0 7470 0 -1 11730
box -36 -24 276 816
use BUFX2  BUFX2_insert28
timestamp 1727136778
transform 1 0 9630 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert29
timestamp 1727136778
transform -1 0 6870 0 1 7050
box -36 -24 276 816
use BUFX2  BUFX2_insert30
timestamp 1727136778
transform 1 0 10230 0 1 7050
box -36 -24 276 816
use BUFX2  BUFX2_insert31
timestamp 1727136778
transform -1 0 6930 0 -1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert32
timestamp 1727136778
transform 1 0 10650 0 1 13290
box -36 -24 276 816
use BUFX2  BUFX2_insert33
timestamp 1727136778
transform -1 0 15510 0 -1 16410
box -36 -24 276 816
use BUFX2  BUFX2_insert34
timestamp 1727136778
transform -1 0 18330 0 -1 16410
box -36 -24 276 816
use BUFX2  BUFX2_insert35
timestamp 1727136778
transform -1 0 15150 0 -1 17970
box -36 -24 276 816
use BUFX2  BUFX2_insert36
timestamp 1727136778
transform -1 0 18150 0 1 16410
box -36 -24 276 816
use CLKBUF1  CLKBUF1_insert8 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 14250 0 -1 11730
box -36 -24 636 816
use CLKBUF1  CLKBUF1_insert9
timestamp 1727136778
transform -1 0 15510 0 1 8610
box -36 -24 636 816
use CLKBUF1  CLKBUF1_insert10
timestamp 1727136778
transform -1 0 18090 0 1 2370
box -36 -24 636 816
use CLKBUF1  CLKBUF1_insert11
timestamp 1727136778
transform -1 0 16170 0 -1 11730
box -36 -24 636 816
use CLKBUF1  CLKBUF1_insert12
timestamp 1727136778
transform -1 0 15570 0 -1 3930
box -36 -24 636 816
use FILL  FILL89850x150 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1700315010
transform -1 0 18030 0 -1 810
box -36 -24 96 816
use FILL  FILL90150x150
timestamp 1700315010
transform -1 0 18090 0 -1 810
box -36 -24 96 816
use FILL  FILL90150x4050
timestamp 1700315010
transform 1 0 18030 0 1 810
box -36 -24 96 816
use FILL  FILL90150x89850
timestamp 1700315010
transform 1 0 18030 0 1 17970
box -36 -24 96 816
use FILL  FILL90450x150
timestamp 1700315010
transform -1 0 18150 0 -1 810
box -36 -24 96 816
use FILL  FILL90450x4050
timestamp 1700315010
transform 1 0 18090 0 1 810
box -36 -24 96 816
use FILL  FILL90450x7950
timestamp 1700315010
transform -1 0 18150 0 -1 2370
box -36 -24 96 816
use FILL  FILL90450x11850
timestamp 1700315010
transform 1 0 18090 0 1 2370
box -36 -24 96 816
use FILL  FILL90450x27450
timestamp 1700315010
transform 1 0 18090 0 1 5490
box -36 -24 96 816
use FILL  FILL90450x31350
timestamp 1700315010
transform -1 0 18150 0 -1 7050
box -36 -24 96 816
use FILL  FILL90450x85950
timestamp 1700315010
transform -1 0 18150 0 -1 17970
box -36 -24 96 816
use FILL  FILL90450x89850
timestamp 1700315010
transform 1 0 18090 0 1 17970
box -36 -24 96 816
use FILL  FILL90750x150
timestamp 1700315010
transform -1 0 18210 0 -1 810
box -36 -24 96 816
use FILL  FILL90750x4050
timestamp 1700315010
transform 1 0 18150 0 1 810
box -36 -24 96 816
use FILL  FILL90750x7950
timestamp 1700315010
transform -1 0 18210 0 -1 2370
box -36 -24 96 816
use FILL  FILL90750x11850
timestamp 1700315010
transform 1 0 18150 0 1 2370
box -36 -24 96 816
use FILL  FILL90750x19650
timestamp 1700315010
transform 1 0 18150 0 1 3930
box -36 -24 96 816
use FILL  FILL90750x23550
timestamp 1700315010
transform -1 0 18210 0 -1 5490
box -36 -24 96 816
use FILL  FILL90750x27450
timestamp 1700315010
transform 1 0 18150 0 1 5490
box -36 -24 96 816
use FILL  FILL90750x31350
timestamp 1700315010
transform -1 0 18210 0 -1 7050
box -36 -24 96 816
use FILL  FILL90750x39150
timestamp 1700315010
transform -1 0 18210 0 -1 8610
box -36 -24 96 816
use FILL  FILL90750x82050
timestamp 1700315010
transform 1 0 18150 0 1 16410
box -36 -24 96 816
use FILL  FILL90750x85950
timestamp 1700315010
transform -1 0 18210 0 -1 17970
box -36 -24 96 816
use FILL  FILL90750x89850
timestamp 1700315010
transform 1 0 18150 0 1 17970
box -36 -24 96 816
use FILL  FILL91050x150
timestamp 1700315010
transform -1 0 18270 0 -1 810
box -36 -24 96 816
use FILL  FILL91050x4050
timestamp 1700315010
transform 1 0 18210 0 1 810
box -36 -24 96 816
use FILL  FILL91050x7950
timestamp 1700315010
transform -1 0 18270 0 -1 2370
box -36 -24 96 816
use FILL  FILL91050x11850
timestamp 1700315010
transform 1 0 18210 0 1 2370
box -36 -24 96 816
use FILL  FILL91050x15750
timestamp 1700315010
transform -1 0 18270 0 -1 3930
box -36 -24 96 816
use FILL  FILL91050x19650
timestamp 1700315010
transform 1 0 18210 0 1 3930
box -36 -24 96 816
use FILL  FILL91050x23550
timestamp 1700315010
transform -1 0 18270 0 -1 5490
box -36 -24 96 816
use FILL  FILL91050x27450
timestamp 1700315010
transform 1 0 18210 0 1 5490
box -36 -24 96 816
use FILL  FILL91050x31350
timestamp 1700315010
transform -1 0 18270 0 -1 7050
box -36 -24 96 816
use FILL  FILL91050x39150
timestamp 1700315010
transform -1 0 18270 0 -1 8610
box -36 -24 96 816
use FILL  FILL91050x54750
timestamp 1700315010
transform -1 0 18270 0 -1 11730
box -36 -24 96 816
use FILL  FILL91050x62550
timestamp 1700315010
transform -1 0 18270 0 -1 13290
box -36 -24 96 816
use FILL  FILL91050x70350
timestamp 1700315010
transform -1 0 18270 0 -1 14850
box -36 -24 96 816
use FILL  FILL91050x74250
timestamp 1700315010
transform 1 0 18210 0 1 14850
box -36 -24 96 816
use FILL  FILL91050x82050
timestamp 1700315010
transform 1 0 18210 0 1 16410
box -36 -24 96 816
use FILL  FILL91050x85950
timestamp 1700315010
transform -1 0 18270 0 -1 17970
box -36 -24 96 816
use FILL  FILL91050x89850
timestamp 1700315010
transform 1 0 18210 0 1 17970
box -36 -24 96 816
use FILL  FILL91350x150
timestamp 1700315010
transform -1 0 18330 0 -1 810
box -36 -24 96 816
use FILL  FILL91350x4050
timestamp 1700315010
transform 1 0 18270 0 1 810
box -36 -24 96 816
use FILL  FILL91350x7950
timestamp 1700315010
transform -1 0 18330 0 -1 2370
box -36 -24 96 816
use FILL  FILL91350x11850
timestamp 1700315010
transform 1 0 18270 0 1 2370
box -36 -24 96 816
use FILL  FILL91350x15750
timestamp 1700315010
transform -1 0 18330 0 -1 3930
box -36 -24 96 816
use FILL  FILL91350x19650
timestamp 1700315010
transform 1 0 18270 0 1 3930
box -36 -24 96 816
use FILL  FILL91350x23550
timestamp 1700315010
transform -1 0 18330 0 -1 5490
box -36 -24 96 816
use FILL  FILL91350x27450
timestamp 1700315010
transform 1 0 18270 0 1 5490
box -36 -24 96 816
use FILL  FILL91350x31350
timestamp 1700315010
transform -1 0 18330 0 -1 7050
box -36 -24 96 816
use FILL  FILL91350x35250
timestamp 1700315010
transform 1 0 18270 0 1 7050
box -36 -24 96 816
use FILL  FILL91350x39150
timestamp 1700315010
transform -1 0 18330 0 -1 8610
box -36 -24 96 816
use FILL  FILL91350x46950
timestamp 1700315010
transform -1 0 18330 0 -1 10170
box -36 -24 96 816
use FILL  FILL91350x54750
timestamp 1700315010
transform -1 0 18330 0 -1 11730
box -36 -24 96 816
use FILL  FILL91350x62550
timestamp 1700315010
transform -1 0 18330 0 -1 13290
box -36 -24 96 816
use FILL  FILL91350x70350
timestamp 1700315010
transform -1 0 18330 0 -1 14850
box -36 -24 96 816
use FILL  FILL91350x74250
timestamp 1700315010
transform 1 0 18270 0 1 14850
box -36 -24 96 816
use FILL  FILL91350x82050
timestamp 1700315010
transform 1 0 18270 0 1 16410
box -36 -24 96 816
use FILL  FILL91350x85950
timestamp 1700315010
transform -1 0 18330 0 -1 17970
box -36 -24 96 816
use FILL  FILL91350x89850
timestamp 1700315010
transform 1 0 18270 0 1 17970
box -36 -24 96 816
use FILL  FILL91650x150
timestamp 1700315010
transform -1 0 18390 0 -1 810
box -36 -24 96 816
use FILL  FILL91650x4050
timestamp 1700315010
transform 1 0 18330 0 1 810
box -36 -24 96 816
use FILL  FILL91650x7950
timestamp 1700315010
transform -1 0 18390 0 -1 2370
box -36 -24 96 816
use FILL  FILL91650x11850
timestamp 1700315010
transform 1 0 18330 0 1 2370
box -36 -24 96 816
use FILL  FILL91650x15750
timestamp 1700315010
transform -1 0 18390 0 -1 3930
box -36 -24 96 816
use FILL  FILL91650x19650
timestamp 1700315010
transform 1 0 18330 0 1 3930
box -36 -24 96 816
use FILL  FILL91650x23550
timestamp 1700315010
transform -1 0 18390 0 -1 5490
box -36 -24 96 816
use FILL  FILL91650x27450
timestamp 1700315010
transform 1 0 18330 0 1 5490
box -36 -24 96 816
use FILL  FILL91650x31350
timestamp 1700315010
transform -1 0 18390 0 -1 7050
box -36 -24 96 816
use FILL  FILL91650x35250
timestamp 1700315010
transform 1 0 18330 0 1 7050
box -36 -24 96 816
use FILL  FILL91650x39150
timestamp 1700315010
transform -1 0 18390 0 -1 8610
box -36 -24 96 816
use FILL  FILL91650x43050
timestamp 1700315010
transform 1 0 18330 0 1 8610
box -36 -24 96 816
use FILL  FILL91650x46950
timestamp 1700315010
transform -1 0 18390 0 -1 10170
box -36 -24 96 816
use FILL  FILL91650x50850
timestamp 1700315010
transform 1 0 18330 0 1 10170
box -36 -24 96 816
use FILL  FILL91650x54750
timestamp 1700315010
transform -1 0 18390 0 -1 11730
box -36 -24 96 816
use FILL  FILL91650x62550
timestamp 1700315010
transform -1 0 18390 0 -1 13290
box -36 -24 96 816
use FILL  FILL91650x70350
timestamp 1700315010
transform -1 0 18390 0 -1 14850
box -36 -24 96 816
use FILL  FILL91650x74250
timestamp 1700315010
transform 1 0 18330 0 1 14850
box -36 -24 96 816
use FILL  FILL91650x78150
timestamp 1700315010
transform -1 0 18390 0 -1 16410
box -36 -24 96 816
use FILL  FILL91650x82050
timestamp 1700315010
transform 1 0 18330 0 1 16410
box -36 -24 96 816
use FILL  FILL91650x85950
timestamp 1700315010
transform -1 0 18390 0 -1 17970
box -36 -24 96 816
use FILL  FILL91650x89850
timestamp 1700315010
transform 1 0 18330 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__889_
timestamp 1700315010
transform 1 0 15990 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__890_
timestamp 1700315010
transform -1 0 14850 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__891_
timestamp 1700315010
transform -1 0 15270 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__892_
timestamp 1700315010
transform 1 0 16050 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__893_
timestamp 1700315010
transform -1 0 15630 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__894_
timestamp 1700315010
transform 1 0 16410 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__895_
timestamp 1700315010
transform -1 0 15690 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__896_
timestamp 1700315010
transform -1 0 15270 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__897_
timestamp 1700315010
transform 1 0 15270 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__898_
timestamp 1700315010
transform -1 0 16410 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__899_
timestamp 1700315010
transform 1 0 15690 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__900_
timestamp 1700315010
transform -1 0 17490 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__901_
timestamp 1700315010
transform -1 0 17070 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__902_
timestamp 1700315010
transform 1 0 17310 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__903_
timestamp 1700315010
transform 1 0 14610 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__904_
timestamp 1700315010
transform -1 0 15990 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__905_
timestamp 1700315010
transform -1 0 17010 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__906_
timestamp 1700315010
transform -1 0 12570 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__907_
timestamp 1700315010
transform 1 0 14910 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__908_
timestamp 1700315010
transform 1 0 17790 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__909_
timestamp 1700315010
transform 1 0 16710 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__910_
timestamp 1700315010
transform 1 0 16530 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__911_
timestamp 1700315010
transform 1 0 16170 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__912_
timestamp 1700315010
transform 1 0 17190 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__913_
timestamp 1700315010
transform -1 0 16650 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__914_
timestamp 1700315010
transform -1 0 15690 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__915_
timestamp 1700315010
transform 1 0 15630 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__916_
timestamp 1700315010
transform -1 0 16830 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__917_
timestamp 1700315010
transform 1 0 17430 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__918_
timestamp 1700315010
transform -1 0 16110 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__919_
timestamp 1700315010
transform 1 0 16110 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__920_
timestamp 1700315010
transform -1 0 16650 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__921_
timestamp 1700315010
transform 1 0 16890 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__922_
timestamp 1700315010
transform 1 0 16050 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__923_
timestamp 1700315010
transform 1 0 17670 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__924_
timestamp 1700315010
transform 1 0 17610 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__925_
timestamp 1700315010
transform -1 0 17850 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__926_
timestamp 1700315010
transform -1 0 12930 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__927_
timestamp 1700315010
transform 1 0 14490 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__928_
timestamp 1700315010
transform 1 0 14010 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__929_
timestamp 1700315010
transform 1 0 12570 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__930_
timestamp 1700315010
transform 1 0 10950 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__931_
timestamp 1700315010
transform -1 0 11430 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__932_
timestamp 1700315010
transform 1 0 12330 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__933_
timestamp 1700315010
transform -1 0 13170 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__934_
timestamp 1700315010
transform 1 0 13530 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__935_
timestamp 1700315010
transform -1 0 16110 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__936_
timestamp 1700315010
transform 1 0 12150 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__937_
timestamp 1700315010
transform -1 0 11910 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__938_
timestamp 1700315010
transform -1 0 11910 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__939_
timestamp 1700315010
transform 1 0 10890 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__940_
timestamp 1700315010
transform 1 0 10290 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__941_
timestamp 1700315010
transform -1 0 9690 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__942_
timestamp 1700315010
transform 1 0 10830 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__943_
timestamp 1700315010
transform 1 0 10350 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__944_
timestamp 1700315010
transform -1 0 15870 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__945_
timestamp 1700315010
transform 1 0 16650 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__946_
timestamp 1700315010
transform 1 0 16170 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__947_
timestamp 1700315010
transform 1 0 16890 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__948_
timestamp 1700315010
transform 1 0 15690 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__949_
timestamp 1700315010
transform 1 0 15210 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__950_
timestamp 1700315010
transform -1 0 13890 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__951_
timestamp 1700315010
transform 1 0 11670 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__952_
timestamp 1700315010
transform 1 0 6930 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__953_
timestamp 1700315010
transform 1 0 7830 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__954_
timestamp 1700315010
transform -1 0 7410 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__955_
timestamp 1700315010
transform 1 0 8190 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__956_
timestamp 1700315010
transform 1 0 9450 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__957_
timestamp 1700315010
transform 1 0 10410 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__958_
timestamp 1700315010
transform 1 0 10770 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__959_
timestamp 1700315010
transform 1 0 10770 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__960_
timestamp 1700315010
transform 1 0 9450 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__961_
timestamp 1700315010
transform -1 0 10350 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__962_
timestamp 1700315010
transform 1 0 11250 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__963_
timestamp 1700315010
transform 1 0 8670 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__964_
timestamp 1700315010
transform -1 0 7890 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__965_
timestamp 1700315010
transform 1 0 7410 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__966_
timestamp 1700315010
transform 1 0 9930 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__967_
timestamp 1700315010
transform -1 0 8730 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__968_
timestamp 1700315010
transform 1 0 7650 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__969_
timestamp 1700315010
transform -1 0 8250 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__970_
timestamp 1700315010
transform 1 0 9030 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__971_
timestamp 1700315010
transform 1 0 9030 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__972_
timestamp 1700315010
transform -1 0 9510 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__973_
timestamp 1700315010
transform 1 0 9030 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__974_
timestamp 1700315010
transform -1 0 10410 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__975_
timestamp 1700315010
transform 1 0 9090 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__976_
timestamp 1700315010
transform 1 0 7770 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__977_
timestamp 1700315010
transform 1 0 6270 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__978_
timestamp 1700315010
transform 1 0 7410 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__979_
timestamp 1700315010
transform 1 0 6210 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__980_
timestamp 1700315010
transform 1 0 8610 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__981_
timestamp 1700315010
transform 1 0 10830 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__982_
timestamp 1700315010
transform -1 0 10350 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__983_
timestamp 1700315010
transform -1 0 8190 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__984_
timestamp 1700315010
transform -1 0 7230 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__985_
timestamp 1700315010
transform -1 0 6990 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__986_
timestamp 1700315010
transform -1 0 5130 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__987_
timestamp 1700315010
transform -1 0 4710 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__988_
timestamp 1700315010
transform -1 0 4050 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__989_
timestamp 1700315010
transform -1 0 5370 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__990_
timestamp 1700315010
transform 1 0 5490 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__991_
timestamp 1700315010
transform 1 0 7110 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__992_
timestamp 1700315010
transform -1 0 7110 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__993_
timestamp 1700315010
transform 1 0 5970 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__994_
timestamp 1700315010
transform 1 0 7710 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__995_
timestamp 1700315010
transform -1 0 8310 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__996_
timestamp 1700315010
transform 1 0 5010 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__997_
timestamp 1700315010
transform -1 0 4230 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__998_
timestamp 1700315010
transform 1 0 4770 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__999_
timestamp 1700315010
transform 1 0 6510 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1000_
timestamp 1700315010
transform 1 0 6630 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1001_
timestamp 1700315010
transform 1 0 8250 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1002_
timestamp 1700315010
transform 1 0 6930 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1003_
timestamp 1700315010
transform -1 0 8790 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1004_
timestamp 1700315010
transform 1 0 7350 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1005_
timestamp 1700315010
transform -1 0 6930 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1006_
timestamp 1700315010
transform 1 0 6030 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1007_
timestamp 1700315010
transform -1 0 4950 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1008_
timestamp 1700315010
transform 1 0 5250 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1009_
timestamp 1700315010
transform -1 0 5790 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1010_
timestamp 1700315010
transform 1 0 6870 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1011_
timestamp 1700315010
transform -1 0 6570 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1012_
timestamp 1700315010
transform -1 0 4350 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1013_
timestamp 1700315010
transform -1 0 7350 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1014_
timestamp 1700315010
transform -1 0 6510 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1015_
timestamp 1700315010
transform -1 0 6090 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1016_
timestamp 1700315010
transform -1 0 6150 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1017_
timestamp 1700315010
transform 1 0 6510 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1018_
timestamp 1700315010
transform -1 0 7050 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1019_
timestamp 1700315010
transform -1 0 5250 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1020_
timestamp 1700315010
transform -1 0 4470 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1021_
timestamp 1700315010
transform -1 0 4230 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1022_
timestamp 1700315010
transform -1 0 4110 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1023_
timestamp 1700315010
transform 1 0 3330 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1024_
timestamp 1700315010
transform 1 0 4410 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1025_
timestamp 1700315010
transform 1 0 4290 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1026_
timestamp 1700315010
transform 1 0 3690 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1027_
timestamp 1700315010
transform 1 0 4410 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1028_
timestamp 1700315010
transform 1 0 3090 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1029_
timestamp 1700315010
transform -1 0 2670 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1030_
timestamp 1700315010
transform -1 0 4710 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1031_
timestamp 1700315010
transform 1 0 3810 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1032_
timestamp 1700315010
transform -1 0 3630 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1033_
timestamp 1700315010
transform -1 0 3150 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1034_
timestamp 1700315010
transform -1 0 4890 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1035_
timestamp 1700315010
transform -1 0 3210 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1036_
timestamp 1700315010
transform -1 0 3450 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1037_
timestamp 1700315010
transform -1 0 3090 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1038_
timestamp 1700315010
transform 1 0 4830 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1039_
timestamp 1700315010
transform -1 0 3930 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1040_
timestamp 1700315010
transform -1 0 6090 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1041_
timestamp 1700315010
transform -1 0 7890 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1042_
timestamp 1700315010
transform 1 0 5610 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1043_
timestamp 1700315010
transform 1 0 6810 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1044_
timestamp 1700315010
transform 1 0 6690 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1045_
timestamp 1700315010
transform 1 0 6210 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1046_
timestamp 1700315010
transform -1 0 4770 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1047_
timestamp 1700315010
transform 1 0 5190 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1048_
timestamp 1700315010
transform -1 0 5790 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1049_
timestamp 1700315010
transform -1 0 4290 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1050_
timestamp 1700315010
transform 1 0 4410 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1051_
timestamp 1700315010
transform -1 0 2010 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1052_
timestamp 1700315010
transform 1 0 3510 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1053_
timestamp 1700315010
transform 1 0 3570 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1054_
timestamp 1700315010
transform -1 0 4050 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1055_
timestamp 1700315010
transform -1 0 2790 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1056_
timestamp 1700315010
transform 1 0 2910 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1057_
timestamp 1700315010
transform -1 0 5670 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1058_
timestamp 1700315010
transform 1 0 3690 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1059_
timestamp 1700315010
transform 1 0 3210 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1060_
timestamp 1700315010
transform -1 0 3450 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1061_
timestamp 1700315010
transform -1 0 8730 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1062_
timestamp 1700315010
transform -1 0 5670 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1063_
timestamp 1700315010
transform 1 0 6450 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1064_
timestamp 1700315010
transform 1 0 4050 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1065_
timestamp 1700315010
transform -1 0 2730 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1066_
timestamp 1700315010
transform 1 0 3030 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1067_
timestamp 1700315010
transform 1 0 3810 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1068_
timestamp 1700315010
transform -1 0 2490 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1069_
timestamp 1700315010
transform 1 0 3630 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1070_
timestamp 1700315010
transform 1 0 5790 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1071_
timestamp 1700315010
transform 1 0 4650 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1072_
timestamp 1700315010
transform -1 0 570 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1073_
timestamp 1700315010
transform -1 0 2790 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1074_
timestamp 1700315010
transform -1 0 2310 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1075_
timestamp 1700315010
transform -1 0 2310 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1076_
timestamp 1700315010
transform -1 0 2850 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1077_
timestamp 1700315010
transform 1 0 3270 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1078_
timestamp 1700315010
transform -1 0 1410 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1079_
timestamp 1700315010
transform -1 0 2610 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1080_
timestamp 1700315010
transform -1 0 2490 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1081_
timestamp 1700315010
transform -1 0 570 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1082_
timestamp 1700315010
transform -1 0 3030 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1083_
timestamp 1700315010
transform -1 0 2190 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1084_
timestamp 1700315010
transform -1 0 1050 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1085_
timestamp 1700315010
transform -1 0 990 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1086_
timestamp 1700315010
transform 1 0 1950 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1087_
timestamp 1700315010
transform 1 0 1470 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1088_
timestamp 1700315010
transform -1 0 1830 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1089_
timestamp 1700315010
transform 1 0 5790 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1090_
timestamp 1700315010
transform 1 0 4590 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1091_
timestamp 1700315010
transform -1 0 5610 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1092_
timestamp 1700315010
transform -1 0 6030 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1093_
timestamp 1700315010
transform 1 0 5550 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1094_
timestamp 1700315010
transform 1 0 6450 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1095_
timestamp 1700315010
transform -1 0 5490 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1096_
timestamp 1700315010
transform -1 0 5010 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1097_
timestamp 1700315010
transform -1 0 4710 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1098_
timestamp 1700315010
transform -1 0 5130 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1099_
timestamp 1700315010
transform -1 0 4230 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1100_
timestamp 1700315010
transform -1 0 90 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1101_
timestamp 1700315010
transform -1 0 90 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1102_
timestamp 1700315010
transform -1 0 2730 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1103_
timestamp 1700315010
transform 1 0 1770 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1104_
timestamp 1700315010
transform 1 0 1350 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1105_
timestamp 1700315010
transform 1 0 450 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1106_
timestamp 1700315010
transform -1 0 90 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1107_
timestamp 1700315010
transform 1 0 510 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1108_
timestamp 1700315010
transform 1 0 2550 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1109_
timestamp 1700315010
transform -1 0 990 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1110_
timestamp 1700315010
transform -1 0 570 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1111_
timestamp 1700315010
transform -1 0 90 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1112_
timestamp 1700315010
transform -1 0 6030 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1113_
timestamp 1700315010
transform 1 0 1350 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1114_
timestamp 1700315010
transform -1 0 5250 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1115_
timestamp 1700315010
transform -1 0 1470 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1116_
timestamp 1700315010
transform -1 0 1830 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1117_
timestamp 1700315010
transform 1 0 2190 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1118_
timestamp 1700315010
transform -1 0 990 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1119_
timestamp 1700315010
transform 1 0 1410 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1120_
timestamp 1700315010
transform 1 0 1350 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1121_
timestamp 1700315010
transform 1 0 2610 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1122_
timestamp 1700315010
transform -1 0 2190 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1123_
timestamp 1700315010
transform -1 0 1890 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1124_
timestamp 1700315010
transform 1 0 1470 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1125_
timestamp 1700315010
transform 1 0 510 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1126_
timestamp 1700315010
transform -1 0 90 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1127_
timestamp 1700315010
transform 1 0 1650 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1128_
timestamp 1700315010
transform -1 0 930 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1129_
timestamp 1700315010
transform -1 0 570 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1130_
timestamp 1700315010
transform 1 0 990 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1131_
timestamp 1700315010
transform -1 0 990 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1132_
timestamp 1700315010
transform -1 0 2370 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1133_
timestamp 1700315010
transform -1 0 90 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1134_
timestamp 1700315010
transform -1 0 570 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1135_
timestamp 1700315010
transform 1 0 510 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1136_
timestamp 1700315010
transform -1 0 870 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1137_
timestamp 1700315010
transform -1 0 90 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1138_
timestamp 1700315010
transform 1 0 1410 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1139_
timestamp 1700315010
transform 1 0 1710 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1140_
timestamp 1700315010
transform 1 0 5310 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1141_
timestamp 1700315010
transform 1 0 6750 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1142_
timestamp 1700315010
transform 1 0 7470 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1143_
timestamp 1700315010
transform 1 0 9870 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1144_
timestamp 1700315010
transform 1 0 10890 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1145_
timestamp 1700315010
transform 1 0 8970 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1146_
timestamp 1700315010
transform -1 0 9990 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1147_
timestamp 1700315010
transform -1 0 8670 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1148_
timestamp 1700315010
transform 1 0 9450 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1149_
timestamp 1700315010
transform -1 0 9510 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1150_
timestamp 1700315010
transform 1 0 8370 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1151_
timestamp 1700315010
transform 1 0 9930 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1152_
timestamp 1700315010
transform -1 0 9450 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1153_
timestamp 1700315010
transform 1 0 6990 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1154_
timestamp 1700315010
transform 1 0 7470 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1155_
timestamp 1700315010
transform 1 0 7890 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1156_
timestamp 1700315010
transform -1 0 7890 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1157_
timestamp 1700315010
transform -1 0 3270 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1158_
timestamp 1700315010
transform 1 0 3450 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1159_
timestamp 1700315010
transform -1 0 5130 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1160_
timestamp 1700315010
transform 1 0 1290 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1161_
timestamp 1700315010
transform 1 0 2190 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1162_
timestamp 1700315010
transform 1 0 3930 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1163_
timestamp 1700315010
transform 1 0 9870 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1164_
timestamp 1700315010
transform 1 0 11190 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1165_
timestamp 1700315010
transform -1 0 11670 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1166_
timestamp 1700315010
transform 1 0 12390 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1167_
timestamp 1700315010
transform 1 0 12810 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1168_
timestamp 1700315010
transform -1 0 10350 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1169_
timestamp 1700315010
transform 1 0 11970 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1170_
timestamp 1700315010
transform 1 0 10410 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1171_
timestamp 1700315010
transform 1 0 12090 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1172_
timestamp 1700315010
transform 1 0 11670 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1173_
timestamp 1700315010
transform 1 0 12090 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1174_
timestamp 1700315010
transform 1 0 10710 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1175_
timestamp 1700315010
transform -1 0 11250 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1176_
timestamp 1700315010
transform 1 0 10890 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1177_
timestamp 1700315010
transform -1 0 8910 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1178_
timestamp 1700315010
transform -1 0 8850 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1179_
timestamp 1700315010
transform 1 0 9990 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1180_
timestamp 1700315010
transform 1 0 6270 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1181_
timestamp 1700315010
transform 1 0 9810 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1182_
timestamp 1700315010
transform -1 0 11850 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1183_
timestamp 1700315010
transform 1 0 11310 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1184_
timestamp 1700315010
transform -1 0 10890 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1185_
timestamp 1700315010
transform -1 0 11250 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1186_
timestamp 1700315010
transform 1 0 12030 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1187_
timestamp 1700315010
transform -1 0 9930 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1188_
timestamp 1700315010
transform -1 0 13290 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1189_
timestamp 1700315010
transform 1 0 11190 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1190_
timestamp 1700315010
transform 1 0 11550 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1191_
timestamp 1700315010
transform -1 0 12570 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1192_
timestamp 1700315010
transform 1 0 13350 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1193_
timestamp 1700315010
transform 1 0 12990 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1194_
timestamp 1700315010
transform 1 0 12570 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1195_
timestamp 1700315010
transform 1 0 13350 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1196_
timestamp 1700315010
transform 1 0 11670 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1197_
timestamp 1700315010
transform -1 0 12210 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1198_
timestamp 1700315010
transform 1 0 9270 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1199_
timestamp 1700315010
transform 1 0 8310 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1200_
timestamp 1700315010
transform 1 0 10410 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1201_
timestamp 1700315010
transform -1 0 11250 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1202_
timestamp 1700315010
transform 1 0 12090 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1203_
timestamp 1700315010
transform 1 0 10530 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1204_
timestamp 1700315010
transform -1 0 11070 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1205_
timestamp 1700315010
transform 1 0 7950 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1206_
timestamp 1700315010
transform -1 0 90 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1207_
timestamp 1700315010
transform 1 0 2250 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1208_
timestamp 1700315010
transform -1 0 90 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1209_
timestamp 1700315010
transform 1 0 7050 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1210_
timestamp 1700315010
transform -1 0 4590 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1211_
timestamp 1700315010
transform -1 0 6450 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1212_
timestamp 1700315010
transform 1 0 5430 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1213_
timestamp 1700315010
transform 1 0 6210 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1214_
timestamp 1700315010
transform 1 0 6570 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1215_
timestamp 1700315010
transform -1 0 4110 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1216_
timestamp 1700315010
transform -1 0 5850 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1217_
timestamp 1700315010
transform 1 0 5910 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1218_
timestamp 1700315010
transform -1 0 5370 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1219_
timestamp 1700315010
transform 1 0 3630 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1220_
timestamp 1700315010
transform -1 0 570 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1221_
timestamp 1700315010
transform -1 0 4530 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1222_
timestamp 1700315010
transform -1 0 5670 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1223_
timestamp 1700315010
transform 1 0 5310 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1224_
timestamp 1700315010
transform -1 0 6270 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1225_
timestamp 1700315010
transform 1 0 5730 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1226_
timestamp 1700315010
transform -1 0 4950 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1227_
timestamp 1700315010
transform 1 0 4650 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1228_
timestamp 1700315010
transform 1 0 5850 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1229_
timestamp 1700315010
transform 1 0 6630 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1230_
timestamp 1700315010
transform 1 0 5490 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1231_
timestamp 1700315010
transform -1 0 5070 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1232_
timestamp 1700315010
transform 1 0 2250 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1233_
timestamp 1700315010
transform 1 0 870 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1234_
timestamp 1700315010
transform 1 0 3270 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1235_
timestamp 1700315010
transform 1 0 2730 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1236_
timestamp 1700315010
transform -1 0 810 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1237_
timestamp 1700315010
transform 1 0 1650 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1238_
timestamp 1700315010
transform 1 0 2190 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1239_
timestamp 1700315010
transform -1 0 1470 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1240_
timestamp 1700315010
transform -1 0 1230 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1241_
timestamp 1700315010
transform -1 0 630 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1242_
timestamp 1700315010
transform 1 0 1830 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1243_
timestamp 1700315010
transform 1 0 990 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1244_
timestamp 1700315010
transform 1 0 510 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1245_
timestamp 1700315010
transform -1 0 570 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1246_
timestamp 1700315010
transform -1 0 90 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1247_
timestamp 1700315010
transform -1 0 90 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1248_
timestamp 1700315010
transform 1 0 1650 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1249_
timestamp 1700315010
transform 1 0 30 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1250_
timestamp 1700315010
transform -1 0 570 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1251_
timestamp 1700315010
transform -1 0 3270 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1252_
timestamp 1700315010
transform 1 0 1350 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1253_
timestamp 1700315010
transform 1 0 30 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1254_
timestamp 1700315010
transform -1 0 1890 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1255_
timestamp 1700315010
transform -1 0 90 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1256_
timestamp 1700315010
transform 1 0 930 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1257_
timestamp 1700315010
transform -1 0 2790 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1258_
timestamp 1700315010
transform 1 0 990 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1259_
timestamp 1700315010
transform -1 0 2430 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1260_
timestamp 1700315010
transform -1 0 2430 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1261_
timestamp 1700315010
transform 1 0 2790 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1262_
timestamp 1700315010
transform 1 0 510 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1263_
timestamp 1700315010
transform -1 0 2010 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1264_
timestamp 1700315010
transform 1 0 1410 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1265_
timestamp 1700315010
transform -1 0 1950 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1266_
timestamp 1700315010
transform -1 0 1890 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1267_
timestamp 1700315010
transform -1 0 1050 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1268_
timestamp 1700315010
transform 1 0 3150 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1269_
timestamp 1700315010
transform 1 0 3630 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1270_
timestamp 1700315010
transform 1 0 6990 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1271_
timestamp 1700315010
transform -1 0 9210 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1272_
timestamp 1700315010
transform 1 0 14910 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1273_
timestamp 1700315010
transform -1 0 14190 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1274_
timestamp 1700315010
transform 1 0 12390 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1275_
timestamp 1700315010
transform 1 0 11790 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1276_
timestamp 1700315010
transform -1 0 13350 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1277_
timestamp 1700315010
transform 1 0 12270 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1278_
timestamp 1700315010
transform 1 0 14190 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1279_
timestamp 1700315010
transform 1 0 14070 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1280_
timestamp 1700315010
transform -1 0 10590 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1281_
timestamp 1700315010
transform -1 0 11490 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1282_
timestamp 1700315010
transform -1 0 12150 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1283_
timestamp 1700315010
transform -1 0 11010 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1284_
timestamp 1700315010
transform -1 0 4890 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1285_
timestamp 1700315010
transform -1 0 9750 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1286_
timestamp 1700315010
transform -1 0 4470 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1287_
timestamp 1700315010
transform 1 0 5610 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1288_
timestamp 1700315010
transform 1 0 8910 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1289_
timestamp 1700315010
transform 1 0 8430 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1290_
timestamp 1700315010
transform -1 0 9390 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1291_
timestamp 1700315010
transform -1 0 7110 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1292_
timestamp 1700315010
transform -1 0 6690 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1293_
timestamp 1700315010
transform -1 0 7830 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1294_
timestamp 1700315010
transform 1 0 3690 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1295_
timestamp 1700315010
transform 1 0 3270 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1296_
timestamp 1700315010
transform -1 0 4890 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1297_
timestamp 1700315010
transform 1 0 4770 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1298_
timestamp 1700315010
transform 1 0 930 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1299_
timestamp 1700315010
transform 1 0 2250 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1300_
timestamp 1700315010
transform -1 0 4770 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1301_
timestamp 1700315010
transform 1 0 6090 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1302_
timestamp 1700315010
transform -1 0 5670 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1303_
timestamp 1700315010
transform -1 0 6150 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1304_
timestamp 1700315010
transform -1 0 5190 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1305_
timestamp 1700315010
transform -1 0 4170 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1306_
timestamp 1700315010
transform 1 0 2250 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1307_
timestamp 1700315010
transform 1 0 990 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1308_
timestamp 1700315010
transform -1 0 90 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1309_
timestamp 1700315010
transform 1 0 3870 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1310_
timestamp 1700315010
transform 1 0 4770 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1311_
timestamp 1700315010
transform 1 0 3210 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1312_
timestamp 1700315010
transform -1 0 5190 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1313_
timestamp 1700315010
transform -1 0 3990 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1314_
timestamp 1700315010
transform -1 0 3630 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1315_
timestamp 1700315010
transform 1 0 3810 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1316_
timestamp 1700315010
transform -1 0 2250 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1317_
timestamp 1700315010
transform 1 0 2790 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1318_
timestamp 1700315010
transform 1 0 8250 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1319_
timestamp 1700315010
transform -1 0 6090 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1320_
timestamp 1700315010
transform -1 0 5250 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1321_
timestamp 1700315010
transform -1 0 4770 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1322_
timestamp 1700315010
transform -1 0 3390 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1323_
timestamp 1700315010
transform -1 0 4350 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1324_
timestamp 1700315010
transform -1 0 2370 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1325_
timestamp 1700315010
transform -1 0 2970 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1326_
timestamp 1700315010
transform -1 0 1950 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1327_
timestamp 1700315010
transform -1 0 90 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1328_
timestamp 1700315010
transform -1 0 90 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1329_
timestamp 1700315010
transform 1 0 1830 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1330_
timestamp 1700315010
transform -1 0 1410 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1331_
timestamp 1700315010
transform 1 0 450 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1332_
timestamp 1700315010
transform 1 0 1350 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1333_
timestamp 1700315010
transform 1 0 2310 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1334_
timestamp 1700315010
transform 1 0 1410 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1335_
timestamp 1700315010
transform -1 0 90 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1336_
timestamp 1700315010
transform 1 0 1350 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1337_
timestamp 1700315010
transform 1 0 3270 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1338_
timestamp 1700315010
transform 1 0 30 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1339_
timestamp 1700315010
transform 1 0 2070 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1340_
timestamp 1700315010
transform 1 0 1830 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1341_
timestamp 1700315010
transform 1 0 390 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1342_
timestamp 1700315010
transform -1 0 510 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1343_
timestamp 1700315010
transform 1 0 870 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1344_
timestamp 1700315010
transform -1 0 2550 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1345_
timestamp 1700315010
transform -1 0 4410 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1346_
timestamp 1700315010
transform 1 0 2610 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1347_
timestamp 1700315010
transform 1 0 2970 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1348_
timestamp 1700315010
transform -1 0 3990 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1349_
timestamp 1700315010
transform -1 0 4110 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1350_
timestamp 1700315010
transform 1 0 1470 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1351_
timestamp 1700315010
transform 1 0 2850 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1352_
timestamp 1700315010
transform 1 0 5130 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1353_
timestamp 1700315010
transform -1 0 3510 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1354_
timestamp 1700315010
transform 1 0 5010 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1355_
timestamp 1700315010
transform -1 0 6390 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1356_
timestamp 1700315010
transform 1 0 9750 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1357_
timestamp 1700315010
transform 1 0 10230 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1358_
timestamp 1700315010
transform 1 0 10650 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1359_
timestamp 1700315010
transform 1 0 13590 0 -1 5490
box -36 -24 96 816
use FILL  FILL_0__1360_
timestamp 1700315010
transform 1 0 13410 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1361_
timestamp 1700315010
transform -1 0 12570 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1362_
timestamp 1700315010
transform 1 0 12930 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1363_
timestamp 1700315010
transform -1 0 12090 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1364_
timestamp 1700315010
transform 1 0 11610 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1365_
timestamp 1700315010
transform -1 0 14370 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1366_
timestamp 1700315010
transform -1 0 4590 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1367_
timestamp 1700315010
transform 1 0 4110 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1368_
timestamp 1700315010
transform 1 0 6210 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1369_
timestamp 1700315010
transform 1 0 8670 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1370_
timestamp 1700315010
transform 1 0 6750 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1371_
timestamp 1700315010
transform 1 0 7410 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1372_
timestamp 1700315010
transform -1 0 3750 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1373_
timestamp 1700315010
transform 1 0 2850 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1374_
timestamp 1700315010
transform -1 0 1470 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1375_
timestamp 1700315010
transform -1 0 930 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1376_
timestamp 1700315010
transform -1 0 3810 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1377_
timestamp 1700315010
transform -1 0 2550 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1378_
timestamp 1700315010
transform -1 0 3450 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1379_
timestamp 1700315010
transform -1 0 3030 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1380_
timestamp 1700315010
transform -1 0 3390 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1381_
timestamp 1700315010
transform -1 0 2910 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1382_
timestamp 1700315010
transform -1 0 2130 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1383_
timestamp 1700315010
transform -1 0 2910 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1384_
timestamp 1700315010
transform -1 0 3390 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1385_
timestamp 1700315010
transform -1 0 2430 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1386_
timestamp 1700315010
transform -1 0 630 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1387_
timestamp 1700315010
transform 1 0 1770 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1388_
timestamp 1700315010
transform 1 0 4650 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1389_
timestamp 1700315010
transform -1 0 5370 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1390_
timestamp 1700315010
transform -1 0 4950 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1391_
timestamp 1700315010
transform -1 0 4410 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1392_
timestamp 1700315010
transform 1 0 6030 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1393_
timestamp 1700315010
transform 1 0 5550 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1394_
timestamp 1700315010
transform 1 0 4050 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1395_
timestamp 1700315010
transform 1 0 1170 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1396_
timestamp 1700315010
transform -1 0 1650 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1397_
timestamp 1700315010
transform -1 0 90 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1398_
timestamp 1700315010
transform -1 0 930 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1399_
timestamp 1700315010
transform -1 0 1950 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1400_
timestamp 1700315010
transform -1 0 810 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1401_
timestamp 1700315010
transform -1 0 90 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1402_
timestamp 1700315010
transform -1 0 390 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1403_
timestamp 1700315010
transform 1 0 930 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1404_
timestamp 1700315010
transform -1 0 1410 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1405_
timestamp 1700315010
transform 1 0 930 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1406_
timestamp 1700315010
transform -1 0 90 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1407_
timestamp 1700315010
transform -1 0 90 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1408_
timestamp 1700315010
transform -1 0 1050 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1409_
timestamp 1700315010
transform -1 0 570 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1410_
timestamp 1700315010
transform 1 0 510 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1411_
timestamp 1700315010
transform -1 0 1050 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1412_
timestamp 1700315010
transform 1 0 1770 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1413_
timestamp 1700315010
transform -1 0 90 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1414_
timestamp 1700315010
transform -1 0 1830 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1415_
timestamp 1700315010
transform -1 0 3810 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1416_
timestamp 1700315010
transform 1 0 5610 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1417_
timestamp 1700315010
transform 1 0 3090 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1418_
timestamp 1700315010
transform -1 0 3570 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1419_
timestamp 1700315010
transform 1 0 3990 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1420_
timestamp 1700315010
transform -1 0 7350 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1421_
timestamp 1700315010
transform -1 0 7290 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1422_
timestamp 1700315010
transform 1 0 8250 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1423_
timestamp 1700315010
transform -1 0 7770 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1424_
timestamp 1700315010
transform 1 0 8490 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1425_
timestamp 1700315010
transform -1 0 8910 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1426_
timestamp 1700315010
transform 1 0 9270 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1427_
timestamp 1700315010
transform 1 0 13710 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1428_
timestamp 1700315010
transform -1 0 12810 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1429_
timestamp 1700315010
transform 1 0 12930 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1430_
timestamp 1700315010
transform 1 0 13410 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1431_
timestamp 1700315010
transform -1 0 14070 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1432_
timestamp 1700315010
transform 1 0 14130 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1433_
timestamp 1700315010
transform -1 0 12990 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1434_
timestamp 1700315010
transform 1 0 13830 0 1 3930
box -36 -24 96 816
use FILL  FILL_0__1435_
timestamp 1700315010
transform 1 0 17730 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1436_
timestamp 1700315010
transform -1 0 17250 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1437_
timestamp 1700315010
transform -1 0 11550 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1438_
timestamp 1700315010
transform 1 0 7890 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1439_
timestamp 1700315010
transform 1 0 3750 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1440_
timestamp 1700315010
transform -1 0 3510 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1441_
timestamp 1700315010
transform 1 0 1410 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1442_
timestamp 1700315010
transform 1 0 5370 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1443_
timestamp 1700315010
transform -1 0 6150 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1444_
timestamp 1700315010
transform -1 0 4170 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1445_
timestamp 1700315010
transform -1 0 5130 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1446_
timestamp 1700315010
transform 1 0 4530 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1447_
timestamp 1700315010
transform 1 0 4950 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1448_
timestamp 1700315010
transform 1 0 5310 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1449_
timestamp 1700315010
transform -1 0 5670 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1450_
timestamp 1700315010
transform -1 0 4590 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1451_
timestamp 1700315010
transform 1 0 4890 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1452_
timestamp 1700315010
transform 1 0 5610 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1453_
timestamp 1700315010
transform 1 0 6150 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1454_
timestamp 1700315010
transform 1 0 5670 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1455_
timestamp 1700315010
transform 1 0 8550 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1456_
timestamp 1700315010
transform -1 0 6390 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1457_
timestamp 1700315010
transform -1 0 5790 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1458_
timestamp 1700315010
transform -1 0 4770 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1459_
timestamp 1700315010
transform -1 0 1350 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1460_
timestamp 1700315010
transform 1 0 5130 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1461_
timestamp 1700315010
transform 1 0 2130 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1462_
timestamp 1700315010
transform -1 0 450 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1463_
timestamp 1700315010
transform -1 0 4230 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1464_
timestamp 1700315010
transform -1 0 2610 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1465_
timestamp 1700315010
transform -1 0 3030 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1466_
timestamp 1700315010
transform -1 0 1710 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1467_
timestamp 1700315010
transform -1 0 3870 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1468_
timestamp 1700315010
transform 1 0 4230 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1469_
timestamp 1700315010
transform -1 0 3270 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1470_
timestamp 1700315010
transform -1 0 2610 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1471_
timestamp 1700315010
transform 1 0 2250 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1472_
timestamp 1700315010
transform 1 0 2730 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1473_
timestamp 1700315010
transform 1 0 3630 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1474_
timestamp 1700315010
transform 1 0 8250 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1475_
timestamp 1700315010
transform 1 0 8130 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1476_
timestamp 1700315010
transform 1 0 8850 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1477_
timestamp 1700315010
transform 1 0 9330 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1478_
timestamp 1700315010
transform 1 0 9630 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1479_
timestamp 1700315010
transform 1 0 10470 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1480_
timestamp 1700315010
transform -1 0 12630 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1481_
timestamp 1700315010
transform -1 0 12990 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1482_
timestamp 1700315010
transform 1 0 13830 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1483_
timestamp 1700315010
transform 1 0 16050 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1484_
timestamp 1700315010
transform -1 0 16470 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1485_
timestamp 1700315010
transform 1 0 16410 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1486_
timestamp 1700315010
transform -1 0 16950 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1487_
timestamp 1700315010
transform 1 0 17370 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1488_
timestamp 1700315010
transform 1 0 6450 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1489_
timestamp 1700315010
transform 1 0 6930 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1490_
timestamp 1700315010
transform -1 0 6990 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1491_
timestamp 1700315010
transform -1 0 8550 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1492_
timestamp 1700315010
transform -1 0 6270 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1493_
timestamp 1700315010
transform -1 0 6690 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1494_
timestamp 1700315010
transform 1 0 7590 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1495_
timestamp 1700315010
transform 1 0 8850 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1496_
timestamp 1700315010
transform 1 0 7110 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1497_
timestamp 1700315010
transform 1 0 7710 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1498_
timestamp 1700315010
transform 1 0 8130 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1499_
timestamp 1700315010
transform 1 0 6570 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1500_
timestamp 1700315010
transform 1 0 7230 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1501_
timestamp 1700315010
transform 1 0 8070 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1502_
timestamp 1700315010
transform 1 0 8130 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1503_
timestamp 1700315010
transform 1 0 8250 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1504_
timestamp 1700315010
transform 1 0 8490 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1505_
timestamp 1700315010
transform -1 0 7290 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1506_
timestamp 1700315010
transform -1 0 7830 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1507_
timestamp 1700315010
transform -1 0 7350 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1508_
timestamp 1700315010
transform -1 0 6570 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1509_
timestamp 1700315010
transform 1 0 6030 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1510_
timestamp 1700315010
transform -1 0 5670 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1511_
timestamp 1700315010
transform 1 0 6870 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1512_
timestamp 1700315010
transform -1 0 8070 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1513_
timestamp 1700315010
transform 1 0 9870 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1514_
timestamp 1700315010
transform -1 0 9090 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1515_
timestamp 1700315010
transform 1 0 9390 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1516_
timestamp 1700315010
transform -1 0 7530 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1517_
timestamp 1700315010
transform 1 0 8550 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1518_
timestamp 1700315010
transform -1 0 9570 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1519_
timestamp 1700315010
transform 1 0 8670 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1520_
timestamp 1700315010
transform 1 0 9090 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1521_
timestamp 1700315010
transform 1 0 7590 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1522_
timestamp 1700315010
transform 1 0 8070 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1523_
timestamp 1700315010
transform 1 0 8430 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1524_
timestamp 1700315010
transform 1 0 9810 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1525_
timestamp 1700315010
transform -1 0 16350 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1526_
timestamp 1700315010
transform -1 0 14850 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1527_
timestamp 1700315010
transform 1 0 13350 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1528_
timestamp 1700315010
transform 1 0 12870 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1529_
timestamp 1700315010
transform 1 0 13650 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1530_
timestamp 1700315010
transform -1 0 14490 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1531_
timestamp 1700315010
transform -1 0 15150 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1532_
timestamp 1700315010
transform 1 0 15570 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1533_
timestamp 1700315010
transform -1 0 15990 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1534_
timestamp 1700315010
transform -1 0 15390 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1535_
timestamp 1700315010
transform -1 0 11190 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1536_
timestamp 1700315010
transform 1 0 9450 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1537_
timestamp 1700315010
transform 1 0 8310 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1538_
timestamp 1700315010
transform 1 0 7650 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1539_
timestamp 1700315010
transform 1 0 6810 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1540_
timestamp 1700315010
transform -1 0 7830 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1541_
timestamp 1700315010
transform -1 0 8310 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1542_
timestamp 1700315010
transform -1 0 7350 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1543_
timestamp 1700315010
transform 1 0 7830 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1544_
timestamp 1700315010
transform 1 0 7230 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1545_
timestamp 1700315010
transform -1 0 7350 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1546_
timestamp 1700315010
transform -1 0 7410 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1547_
timestamp 1700315010
transform -1 0 7950 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1548_
timestamp 1700315010
transform -1 0 9030 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1549_
timestamp 1700315010
transform -1 0 8370 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1550_
timestamp 1700315010
transform 1 0 10290 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1551_
timestamp 1700315010
transform 1 0 11610 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1552_
timestamp 1700315010
transform 1 0 12450 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1553_
timestamp 1700315010
transform -1 0 15090 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1554_
timestamp 1700315010
transform 1 0 15570 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1555_
timestamp 1700315010
transform 1 0 15510 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1556_
timestamp 1700315010
transform -1 0 14850 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1557_
timestamp 1700315010
transform -1 0 14490 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1558_
timestamp 1700315010
transform 1 0 7470 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1559_
timestamp 1700315010
transform 1 0 10470 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1560_
timestamp 1700315010
transform 1 0 10830 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1561_
timestamp 1700315010
transform -1 0 8010 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1562_
timestamp 1700315010
transform 1 0 7950 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1563_
timestamp 1700315010
transform 1 0 11010 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1564_
timestamp 1700315010
transform -1 0 6090 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1565_
timestamp 1700315010
transform -1 0 6390 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1566_
timestamp 1700315010
transform -1 0 6810 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1567_
timestamp 1700315010
transform 1 0 8610 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1568_
timestamp 1700315010
transform 1 0 9870 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1569_
timestamp 1700315010
transform 1 0 11730 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1570_
timestamp 1700315010
transform 1 0 9990 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1571_
timestamp 1700315010
transform -1 0 10770 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1572_
timestamp 1700315010
transform 1 0 10230 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1573_
timestamp 1700315010
transform 1 0 12210 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1574_
timestamp 1700315010
transform -1 0 12090 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1575_
timestamp 1700315010
transform 1 0 12870 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1576_
timestamp 1700315010
transform 1 0 12390 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1577_
timestamp 1700315010
transform 1 0 13290 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1578_
timestamp 1700315010
transform 1 0 17010 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1579_
timestamp 1700315010
transform -1 0 15270 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1580_
timestamp 1700315010
transform -1 0 15150 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1581_
timestamp 1700315010
transform 1 0 14550 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1582_
timestamp 1700315010
transform -1 0 13410 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1583_
timestamp 1700315010
transform -1 0 11370 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1584_
timestamp 1700315010
transform 1 0 8730 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1585_
timestamp 1700315010
transform 1 0 9210 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1586_
timestamp 1700315010
transform 1 0 10770 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1587_
timestamp 1700315010
transform 1 0 7530 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1588_
timestamp 1700315010
transform -1 0 11490 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1589_
timestamp 1700315010
transform 1 0 14730 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1590_
timestamp 1700315010
transform 1 0 14250 0 1 2370
box -36 -24 96 816
use FILL  FILL_0__1591_
timestamp 1700315010
transform -1 0 14130 0 -1 2370
box -36 -24 96 816
use FILL  FILL_0__1592_
timestamp 1700315010
transform -1 0 12930 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1593_
timestamp 1700315010
transform -1 0 12930 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0__1594_
timestamp 1700315010
transform 1 0 12810 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1595_
timestamp 1700315010
transform 1 0 11850 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1596_
timestamp 1700315010
transform -1 0 12330 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1597_
timestamp 1700315010
transform 1 0 11910 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1598_
timestamp 1700315010
transform -1 0 12390 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1599_
timestamp 1700315010
transform -1 0 11610 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1600_
timestamp 1700315010
transform -1 0 11970 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1601_
timestamp 1700315010
transform 1 0 9810 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1602_
timestamp 1700315010
transform -1 0 9930 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1603_
timestamp 1700315010
transform 1 0 8730 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1604_
timestamp 1700315010
transform -1 0 9210 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1605_
timestamp 1700315010
transform -1 0 13350 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1606_
timestamp 1700315010
transform -1 0 15390 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1607_
timestamp 1700315010
transform 1 0 13170 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1608_
timestamp 1700315010
transform -1 0 13650 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1636_
timestamp 1700315010
transform -1 0 17610 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1637_
timestamp 1700315010
transform 1 0 17610 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1638_
timestamp 1700315010
transform -1 0 15990 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1639_
timestamp 1700315010
transform 1 0 15510 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1640_
timestamp 1700315010
transform 1 0 15510 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1641_
timestamp 1700315010
transform -1 0 11190 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1642_
timestamp 1700315010
transform -1 0 9390 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1643_
timestamp 1700315010
transform -1 0 8910 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1644_
timestamp 1700315010
transform -1 0 11490 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1645_
timestamp 1700315010
transform -1 0 13110 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1646_
timestamp 1700315010
transform -1 0 12210 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1647_
timestamp 1700315010
transform 1 0 9390 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1648_
timestamp 1700315010
transform 1 0 17250 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1649_
timestamp 1700315010
transform -1 0 12750 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1650_
timestamp 1700315010
transform -1 0 13230 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1651_
timestamp 1700315010
transform 1 0 12810 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1652_
timestamp 1700315010
transform -1 0 10770 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1653_
timestamp 1700315010
transform 1 0 12330 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1654_
timestamp 1700315010
transform 1 0 17310 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1655_
timestamp 1700315010
transform -1 0 16890 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1656_
timestamp 1700315010
transform 1 0 17670 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1657_
timestamp 1700315010
transform 1 0 17250 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1658_
timestamp 1700315010
transform 1 0 16770 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1659_
timestamp 1700315010
transform -1 0 15930 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1660_
timestamp 1700315010
transform -1 0 16470 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1661_
timestamp 1700315010
transform 1 0 15930 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1662_
timestamp 1700315010
transform -1 0 10290 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1663_
timestamp 1700315010
transform -1 0 9810 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1664_
timestamp 1700315010
transform -1 0 10230 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1665_
timestamp 1700315010
transform -1 0 10830 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1666_
timestamp 1700315010
transform -1 0 11370 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1667_
timestamp 1700315010
transform 1 0 11430 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1668_
timestamp 1700315010
transform 1 0 11010 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1669_
timestamp 1700315010
transform -1 0 12030 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1670_
timestamp 1700315010
transform 1 0 12450 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1671_
timestamp 1700315010
transform 1 0 15570 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1672_
timestamp 1700315010
transform -1 0 16890 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1673_
timestamp 1700315010
transform 1 0 16350 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1674_
timestamp 1700315010
transform -1 0 15990 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1675_
timestamp 1700315010
transform -1 0 16530 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1676_
timestamp 1700315010
transform 1 0 16350 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1677_
timestamp 1700315010
transform -1 0 14550 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1678_
timestamp 1700315010
transform -1 0 14670 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1679_
timestamp 1700315010
transform -1 0 13470 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1680_
timestamp 1700315010
transform 1 0 13770 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1681_
timestamp 1700315010
transform -1 0 11910 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1682_
timestamp 1700315010
transform 1 0 13650 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1683_
timestamp 1700315010
transform 1 0 14010 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1684_
timestamp 1700315010
transform 1 0 14970 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1685_
timestamp 1700315010
transform -1 0 12450 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1686_
timestamp 1700315010
transform 1 0 12810 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1687_
timestamp 1700315010
transform -1 0 15210 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1688_
timestamp 1700315010
transform 1 0 15570 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1689_
timestamp 1700315010
transform 1 0 14550 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1690_
timestamp 1700315010
transform 1 0 15150 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1691_
timestamp 1700315010
transform -1 0 14730 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1692_
timestamp 1700315010
transform 1 0 10650 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1693_
timestamp 1700315010
transform 1 0 9210 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1694_
timestamp 1700315010
transform -1 0 9750 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1695_
timestamp 1700315010
transform -1 0 8730 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1696_
timestamp 1700315010
transform -1 0 9030 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1697_
timestamp 1700315010
transform -1 0 9810 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1698_
timestamp 1700315010
transform 1 0 10230 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1699_
timestamp 1700315010
transform -1 0 11550 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1700_
timestamp 1700315010
transform -1 0 11610 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1701_
timestamp 1700315010
transform -1 0 10710 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1702_
timestamp 1700315010
transform 1 0 11070 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1703_
timestamp 1700315010
transform -1 0 13650 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1704_
timestamp 1700315010
transform -1 0 14310 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1705_
timestamp 1700315010
transform 1 0 12030 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1706_
timestamp 1700315010
transform -1 0 12930 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1707_
timestamp 1700315010
transform -1 0 13350 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1708_
timestamp 1700315010
transform 1 0 13350 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1709_
timestamp 1700315010
transform -1 0 10890 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1710_
timestamp 1700315010
transform -1 0 11550 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1711_
timestamp 1700315010
transform -1 0 10590 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1712_
timestamp 1700315010
transform -1 0 11010 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1713_
timestamp 1700315010
transform -1 0 10110 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1714_
timestamp 1700315010
transform 1 0 11250 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1715_
timestamp 1700315010
transform -1 0 11730 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1716_
timestamp 1700315010
transform 1 0 12150 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1717_
timestamp 1700315010
transform -1 0 13230 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1718_
timestamp 1700315010
transform 1 0 13590 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1719_
timestamp 1700315010
transform 1 0 14070 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1720_
timestamp 1700315010
transform 1 0 12630 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1721_
timestamp 1700315010
transform 1 0 13890 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1722_
timestamp 1700315010
transform 1 0 14190 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1723_
timestamp 1700315010
transform 1 0 14310 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0__1724_
timestamp 1700315010
transform -1 0 14310 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1725_
timestamp 1700315010
transform 1 0 13170 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1726_
timestamp 1700315010
transform -1 0 12750 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1727_
timestamp 1700315010
transform -1 0 13050 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1728_
timestamp 1700315010
transform -1 0 8970 0 1 16410
box -36 -24 96 816
use FILL  FILL_0__1729_
timestamp 1700315010
transform 1 0 9150 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1730_
timestamp 1700315010
transform -1 0 9630 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1731_
timestamp 1700315010
transform -1 0 10050 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1732_
timestamp 1700315010
transform 1 0 10530 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1733_
timestamp 1700315010
transform 1 0 10950 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1734_
timestamp 1700315010
transform 1 0 14790 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1735_
timestamp 1700315010
transform 1 0 14670 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1736_
timestamp 1700315010
transform -1 0 15630 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1737_
timestamp 1700315010
transform 1 0 15090 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1738_
timestamp 1700315010
transform 1 0 15210 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1739_
timestamp 1700315010
transform 1 0 14670 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1740_
timestamp 1700315010
transform -1 0 15390 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1741_
timestamp 1700315010
transform 1 0 15570 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1742_
timestamp 1700315010
transform 1 0 10470 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1743_
timestamp 1700315010
transform -1 0 8250 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1744_
timestamp 1700315010
transform -1 0 8730 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1745_
timestamp 1700315010
transform -1 0 9630 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1746_
timestamp 1700315010
transform 1 0 9090 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1747_
timestamp 1700315010
transform 1 0 9990 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1748_
timestamp 1700315010
transform -1 0 15210 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1749_
timestamp 1700315010
transform 1 0 15570 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1750_
timestamp 1700315010
transform 1 0 16230 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1751_
timestamp 1700315010
transform 1 0 16050 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1752_
timestamp 1700315010
transform -1 0 15750 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1753_
timestamp 1700315010
transform 1 0 16050 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1754_
timestamp 1700315010
transform 1 0 15390 0 1 5490
box -36 -24 96 816
use FILL  FILL_0__1755_
timestamp 1700315010
transform 1 0 16050 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1756_
timestamp 1700315010
transform 1 0 14430 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1757_
timestamp 1700315010
transform -1 0 13110 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1758_
timestamp 1700315010
transform 1 0 12630 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1759_
timestamp 1700315010
transform 1 0 11910 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1760_
timestamp 1700315010
transform 1 0 13470 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1761_
timestamp 1700315010
transform -1 0 14010 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1762_
timestamp 1700315010
transform -1 0 15330 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1763_
timestamp 1700315010
transform 1 0 15750 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1764_
timestamp 1700315010
transform 1 0 16710 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1765_
timestamp 1700315010
transform 1 0 17130 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1766_
timestamp 1700315010
transform 1 0 17430 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1767_
timestamp 1700315010
transform 1 0 14610 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1768_
timestamp 1700315010
transform -1 0 14190 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1769_
timestamp 1700315010
transform -1 0 13710 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1770_
timestamp 1700315010
transform -1 0 14970 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1771_
timestamp 1700315010
transform 1 0 16470 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1772_
timestamp 1700315010
transform 1 0 16530 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1773_
timestamp 1700315010
transform -1 0 17370 0 1 17970
box -36 -24 96 816
use FILL  FILL_0__1774_
timestamp 1700315010
transform -1 0 16710 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1775_
timestamp 1700315010
transform -1 0 17070 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1776_
timestamp 1700315010
transform 1 0 17070 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1777_
timestamp 1700315010
transform 1 0 14730 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1778_
timestamp 1700315010
transform 1 0 13350 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1779_
timestamp 1700315010
transform 1 0 12990 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1780_
timestamp 1700315010
transform 1 0 12450 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1781_
timestamp 1700315010
transform 1 0 13830 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1782_
timestamp 1700315010
transform 1 0 14310 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1783_
timestamp 1700315010
transform 1 0 16770 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1784_
timestamp 1700315010
transform 1 0 16350 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1785_
timestamp 1700315010
transform -1 0 17370 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1786_
timestamp 1700315010
transform 1 0 17790 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1787_
timestamp 1700315010
transform -1 0 17610 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1788_
timestamp 1700315010
transform 1 0 17070 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1789_
timestamp 1700315010
transform 1 0 17910 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1790_
timestamp 1700315010
transform 1 0 17910 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1791_
timestamp 1700315010
transform 1 0 17850 0 1 7050
box -36 -24 96 816
use FILL  FILL_0__1792_
timestamp 1700315010
transform 1 0 13890 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1793_
timestamp 1700315010
transform 1 0 13470 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1794_
timestamp 1700315010
transform 1 0 14550 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1795_
timestamp 1700315010
transform -1 0 16650 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1796_
timestamp 1700315010
transform 1 0 16170 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1797_
timestamp 1700315010
transform -1 0 15030 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1798_
timestamp 1700315010
transform -1 0 17550 0 1 11730
box -36 -24 96 816
use FILL  FILL_0__1799_
timestamp 1700315010
transform -1 0 17550 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0__1800_
timestamp 1700315010
transform -1 0 17490 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1801_
timestamp 1700315010
transform 1 0 16170 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1802_
timestamp 1700315010
transform 1 0 14190 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0__1803_
timestamp 1700315010
transform 1 0 17550 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1804_
timestamp 1700315010
transform -1 0 17610 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1805_
timestamp 1700315010
transform 1 0 17910 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1806_
timestamp 1700315010
transform -1 0 17010 0 1 13290
box -36 -24 96 816
use FILL  FILL_0__1807_
timestamp 1700315010
transform 1 0 16950 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1808_
timestamp 1700315010
transform 1 0 16530 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1809_
timestamp 1700315010
transform 1 0 16830 0 1 14850
box -36 -24 96 816
use FILL  FILL_0__1810_
timestamp 1700315010
transform 1 0 17610 0 -1 14850
box -36 -24 96 816
use FILL  FILL_0__1811_
timestamp 1700315010
transform 1 0 17130 0 1 810
box -36 -24 96 816
use FILL  FILL_0__1812_
timestamp 1700315010
transform 1 0 17850 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0__1813_
timestamp 1700315010
transform -1 0 17910 0 1 10170
box -36 -24 96 816
use FILL  FILL_0__1814_
timestamp 1700315010
transform -1 0 17970 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1815_
timestamp 1700315010
transform 1 0 17430 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0__1816_
timestamp 1700315010
transform -1 0 17910 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1817_
timestamp 1700315010
transform -1 0 17550 0 1 8610
box -36 -24 96 816
use FILL  FILL_0__1818_
timestamp 1700315010
transform -1 0 9750 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1819_
timestamp 1700315010
transform -1 0 7710 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0__1820_
timestamp 1700315010
transform -1 0 13770 0 -1 3930
box -36 -24 96 816
use FILL  FILL_0__1821_
timestamp 1700315010
transform -1 0 16830 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1822_
timestamp 1700315010
transform 1 0 16350 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1823_
timestamp 1700315010
transform 1 0 15990 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1824_
timestamp 1700315010
transform 1 0 14850 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1825_
timestamp 1700315010
transform 1 0 13710 0 -1 810
box -36 -24 96 816
use FILL  FILL_0__1826_
timestamp 1700315010
transform 1 0 17190 0 -1 810
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert0
timestamp 1700315010
transform 1 0 11730 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert1
timestamp 1700315010
transform -1 0 6570 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert2
timestamp 1700315010
transform -1 0 6930 0 1 7050
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert3
timestamp 1700315010
transform -1 0 6750 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert4
timestamp 1700315010
transform -1 0 13170 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert5
timestamp 1700315010
transform -1 0 11250 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert6
timestamp 1700315010
transform -1 0 8130 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert7
timestamp 1700315010
transform -1 0 10170 0 -1 7050
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert13
timestamp 1700315010
transform 1 0 15510 0 1 8610
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert14
timestamp 1700315010
transform -1 0 11430 0 1 10170
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert15
timestamp 1700315010
transform -1 0 12990 0 1 10170
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert16
timestamp 1700315010
transform -1 0 12030 0 -1 8610
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert17
timestamp 1700315010
transform 1 0 7530 0 1 11730
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert18
timestamp 1700315010
transform -1 0 6990 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert19
timestamp 1700315010
transform 1 0 9030 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert20
timestamp 1700315010
transform -1 0 7230 0 1 8610
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert21
timestamp 1700315010
transform 1 0 15930 0 1 8610
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert22
timestamp 1700315010
transform -1 0 12570 0 1 10170
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert23
timestamp 1700315010
transform 1 0 12690 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert24
timestamp 1700315010
transform 1 0 15810 0 -1 10170
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert25
timestamp 1700315010
transform -1 0 6990 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert26
timestamp 1700315010
transform -1 0 7890 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert27
timestamp 1700315010
transform -1 0 7170 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert28
timestamp 1700315010
transform 1 0 9450 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert29
timestamp 1700315010
transform -1 0 6510 0 1 7050
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert30
timestamp 1700315010
transform 1 0 10110 0 1 7050
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert31
timestamp 1700315010
transform -1 0 6570 0 -1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert32
timestamp 1700315010
transform 1 0 10470 0 1 13290
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert33
timestamp 1700315010
transform -1 0 15210 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert34
timestamp 1700315010
transform -1 0 17970 0 -1 16410
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert35
timestamp 1700315010
transform -1 0 14790 0 -1 17970
box -36 -24 96 816
use FILL  FILL_0_BUFX2_insert36
timestamp 1700315010
transform -1 0 17790 0 1 16410
box -36 -24 96 816
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1700315010
transform -1 0 13590 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 14790 0 1 8610
box -36 -24 96 816
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 17370 0 1 2370
box -36 -24 96 816
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1700315010
transform -1 0 15510 0 -1 11730
box -36 -24 96 816
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 14850 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__889_
timestamp 1700315010
transform 1 0 16050 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__890_
timestamp 1700315010
transform -1 0 14910 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__891_
timestamp 1700315010
transform -1 0 15330 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__892_
timestamp 1700315010
transform 1 0 16110 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__893_
timestamp 1700315010
transform -1 0 15690 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__894_
timestamp 1700315010
transform 1 0 16470 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__895_
timestamp 1700315010
transform -1 0 15750 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__896_
timestamp 1700315010
transform -1 0 15330 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__897_
timestamp 1700315010
transform 1 0 15330 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__898_
timestamp 1700315010
transform -1 0 16470 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__899_
timestamp 1700315010
transform 1 0 15750 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__900_
timestamp 1700315010
transform -1 0 17550 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__901_
timestamp 1700315010
transform -1 0 17130 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__902_
timestamp 1700315010
transform 1 0 17370 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__903_
timestamp 1700315010
transform 1 0 14670 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__904_
timestamp 1700315010
transform -1 0 16050 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__905_
timestamp 1700315010
transform -1 0 17070 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__906_
timestamp 1700315010
transform -1 0 12630 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__907_
timestamp 1700315010
transform 1 0 14970 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__908_
timestamp 1700315010
transform 1 0 17850 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__909_
timestamp 1700315010
transform 1 0 16770 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__910_
timestamp 1700315010
transform 1 0 16590 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__911_
timestamp 1700315010
transform 1 0 16230 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__912_
timestamp 1700315010
transform 1 0 17250 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__913_
timestamp 1700315010
transform -1 0 16710 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__914_
timestamp 1700315010
transform -1 0 15750 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__915_
timestamp 1700315010
transform 1 0 15690 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__916_
timestamp 1700315010
transform -1 0 16890 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__917_
timestamp 1700315010
transform 1 0 17490 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__918_
timestamp 1700315010
transform -1 0 16170 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__919_
timestamp 1700315010
transform 1 0 16170 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__920_
timestamp 1700315010
transform -1 0 16710 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__921_
timestamp 1700315010
transform 1 0 16950 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__922_
timestamp 1700315010
transform 1 0 16110 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__923_
timestamp 1700315010
transform 1 0 17730 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__924_
timestamp 1700315010
transform 1 0 17670 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__925_
timestamp 1700315010
transform -1 0 17910 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__926_
timestamp 1700315010
transform -1 0 12990 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__927_
timestamp 1700315010
transform 1 0 14550 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__928_
timestamp 1700315010
transform 1 0 14070 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__929_
timestamp 1700315010
transform 1 0 12630 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__930_
timestamp 1700315010
transform 1 0 11010 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__931_
timestamp 1700315010
transform -1 0 11490 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__932_
timestamp 1700315010
transform 1 0 12390 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__933_
timestamp 1700315010
transform -1 0 13230 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__934_
timestamp 1700315010
transform 1 0 13590 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__935_
timestamp 1700315010
transform -1 0 16170 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__936_
timestamp 1700315010
transform 1 0 12210 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__937_
timestamp 1700315010
transform -1 0 11970 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__938_
timestamp 1700315010
transform -1 0 11970 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__939_
timestamp 1700315010
transform 1 0 10950 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__940_
timestamp 1700315010
transform 1 0 10350 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__941_
timestamp 1700315010
transform -1 0 9750 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__942_
timestamp 1700315010
transform 1 0 10890 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__943_
timestamp 1700315010
transform 1 0 10410 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__944_
timestamp 1700315010
transform -1 0 15930 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__945_
timestamp 1700315010
transform 1 0 16710 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__946_
timestamp 1700315010
transform 1 0 16230 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__947_
timestamp 1700315010
transform 1 0 16950 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__948_
timestamp 1700315010
transform 1 0 15750 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__949_
timestamp 1700315010
transform 1 0 15270 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__950_
timestamp 1700315010
transform -1 0 13950 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__951_
timestamp 1700315010
transform 1 0 11730 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__952_
timestamp 1700315010
transform 1 0 6990 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__953_
timestamp 1700315010
transform 1 0 7890 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__954_
timestamp 1700315010
transform -1 0 7470 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__955_
timestamp 1700315010
transform 1 0 8250 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__956_
timestamp 1700315010
transform 1 0 9510 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__957_
timestamp 1700315010
transform 1 0 10470 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__958_
timestamp 1700315010
transform 1 0 10830 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__959_
timestamp 1700315010
transform 1 0 10830 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__960_
timestamp 1700315010
transform 1 0 9510 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__961_
timestamp 1700315010
transform -1 0 10410 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__962_
timestamp 1700315010
transform 1 0 11310 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__963_
timestamp 1700315010
transform 1 0 8730 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__964_
timestamp 1700315010
transform -1 0 7950 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__965_
timestamp 1700315010
transform 1 0 7470 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__966_
timestamp 1700315010
transform 1 0 9990 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__967_
timestamp 1700315010
transform -1 0 8790 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__968_
timestamp 1700315010
transform 1 0 7710 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__969_
timestamp 1700315010
transform -1 0 8310 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__970_
timestamp 1700315010
transform 1 0 9090 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__971_
timestamp 1700315010
transform 1 0 9090 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__972_
timestamp 1700315010
transform -1 0 9570 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__973_
timestamp 1700315010
transform 1 0 9090 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__974_
timestamp 1700315010
transform -1 0 10470 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__975_
timestamp 1700315010
transform 1 0 9150 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__976_
timestamp 1700315010
transform 1 0 7830 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__977_
timestamp 1700315010
transform 1 0 6330 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__978_
timestamp 1700315010
transform 1 0 7470 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__979_
timestamp 1700315010
transform 1 0 6270 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__980_
timestamp 1700315010
transform 1 0 8670 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__981_
timestamp 1700315010
transform 1 0 10890 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__982_
timestamp 1700315010
transform -1 0 10410 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__983_
timestamp 1700315010
transform -1 0 8250 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__984_
timestamp 1700315010
transform -1 0 7290 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__985_
timestamp 1700315010
transform -1 0 7050 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__986_
timestamp 1700315010
transform -1 0 5190 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__987_
timestamp 1700315010
transform -1 0 4770 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__988_
timestamp 1700315010
transform -1 0 4110 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__989_
timestamp 1700315010
transform -1 0 5430 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__990_
timestamp 1700315010
transform 1 0 5550 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__991_
timestamp 1700315010
transform 1 0 7170 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__992_
timestamp 1700315010
transform -1 0 7170 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__993_
timestamp 1700315010
transform 1 0 6030 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__994_
timestamp 1700315010
transform 1 0 7770 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__995_
timestamp 1700315010
transform -1 0 8370 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__996_
timestamp 1700315010
transform 1 0 5070 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__997_
timestamp 1700315010
transform -1 0 4290 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__998_
timestamp 1700315010
transform 1 0 4830 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__999_
timestamp 1700315010
transform 1 0 6570 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1000_
timestamp 1700315010
transform 1 0 6690 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1001_
timestamp 1700315010
transform 1 0 8310 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1002_
timestamp 1700315010
transform 1 0 6990 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1003_
timestamp 1700315010
transform -1 0 8850 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1004_
timestamp 1700315010
transform 1 0 7410 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1005_
timestamp 1700315010
transform -1 0 6990 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1006_
timestamp 1700315010
transform 1 0 6090 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1007_
timestamp 1700315010
transform -1 0 5010 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1008_
timestamp 1700315010
transform 1 0 5310 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1009_
timestamp 1700315010
transform -1 0 5850 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1010_
timestamp 1700315010
transform 1 0 6930 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1011_
timestamp 1700315010
transform -1 0 6630 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1012_
timestamp 1700315010
transform -1 0 4410 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1013_
timestamp 1700315010
transform -1 0 7410 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1014_
timestamp 1700315010
transform -1 0 6570 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1015_
timestamp 1700315010
transform -1 0 6150 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1016_
timestamp 1700315010
transform -1 0 6210 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1017_
timestamp 1700315010
transform 1 0 6570 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1018_
timestamp 1700315010
transform -1 0 7110 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1019_
timestamp 1700315010
transform -1 0 5310 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1020_
timestamp 1700315010
transform -1 0 4530 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1021_
timestamp 1700315010
transform -1 0 4290 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1022_
timestamp 1700315010
transform -1 0 4170 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1023_
timestamp 1700315010
transform 1 0 3390 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1024_
timestamp 1700315010
transform 1 0 4470 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1025_
timestamp 1700315010
transform 1 0 4350 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1026_
timestamp 1700315010
transform 1 0 3750 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1027_
timestamp 1700315010
transform 1 0 4470 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1028_
timestamp 1700315010
transform 1 0 3150 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1029_
timestamp 1700315010
transform -1 0 2730 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1030_
timestamp 1700315010
transform -1 0 4770 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1031_
timestamp 1700315010
transform 1 0 3870 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1032_
timestamp 1700315010
transform -1 0 3690 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1033_
timestamp 1700315010
transform -1 0 3210 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1034_
timestamp 1700315010
transform -1 0 4950 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1035_
timestamp 1700315010
transform -1 0 3270 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1036_
timestamp 1700315010
transform -1 0 3510 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1037_
timestamp 1700315010
transform -1 0 3150 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1038_
timestamp 1700315010
transform 1 0 4890 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1039_
timestamp 1700315010
transform -1 0 3990 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1040_
timestamp 1700315010
transform -1 0 6150 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1041_
timestamp 1700315010
transform -1 0 7950 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1042_
timestamp 1700315010
transform 1 0 5670 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1043_
timestamp 1700315010
transform 1 0 6870 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1044_
timestamp 1700315010
transform 1 0 6750 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1045_
timestamp 1700315010
transform 1 0 6270 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1046_
timestamp 1700315010
transform -1 0 4830 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1047_
timestamp 1700315010
transform 1 0 5250 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1048_
timestamp 1700315010
transform -1 0 5850 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1049_
timestamp 1700315010
transform -1 0 4350 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1050_
timestamp 1700315010
transform 1 0 4470 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1051_
timestamp 1700315010
transform -1 0 2070 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1052_
timestamp 1700315010
transform 1 0 3570 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1053_
timestamp 1700315010
transform 1 0 3630 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1054_
timestamp 1700315010
transform -1 0 4110 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1055_
timestamp 1700315010
transform -1 0 2850 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1056_
timestamp 1700315010
transform 1 0 2970 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1057_
timestamp 1700315010
transform -1 0 5730 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1058_
timestamp 1700315010
transform 1 0 3750 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1059_
timestamp 1700315010
transform 1 0 3270 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1060_
timestamp 1700315010
transform -1 0 3510 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1061_
timestamp 1700315010
transform -1 0 8790 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1062_
timestamp 1700315010
transform -1 0 5730 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1063_
timestamp 1700315010
transform 1 0 6510 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1064_
timestamp 1700315010
transform 1 0 4110 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1065_
timestamp 1700315010
transform -1 0 2790 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1066_
timestamp 1700315010
transform 1 0 3090 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1067_
timestamp 1700315010
transform 1 0 3870 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1068_
timestamp 1700315010
transform -1 0 2550 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1069_
timestamp 1700315010
transform 1 0 3690 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1070_
timestamp 1700315010
transform 1 0 5850 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1071_
timestamp 1700315010
transform 1 0 4710 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1072_
timestamp 1700315010
transform -1 0 630 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1073_
timestamp 1700315010
transform -1 0 2850 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1074_
timestamp 1700315010
transform -1 0 2370 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1075_
timestamp 1700315010
transform -1 0 2370 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1076_
timestamp 1700315010
transform -1 0 2910 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1077_
timestamp 1700315010
transform 1 0 3330 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1078_
timestamp 1700315010
transform -1 0 1470 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1079_
timestamp 1700315010
transform -1 0 2670 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1080_
timestamp 1700315010
transform -1 0 2550 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1081_
timestamp 1700315010
transform -1 0 630 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1082_
timestamp 1700315010
transform -1 0 3090 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1083_
timestamp 1700315010
transform -1 0 2250 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1084_
timestamp 1700315010
transform -1 0 1110 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1085_
timestamp 1700315010
transform -1 0 1050 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1086_
timestamp 1700315010
transform 1 0 2010 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1087_
timestamp 1700315010
transform 1 0 1530 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1088_
timestamp 1700315010
transform -1 0 1890 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1089_
timestamp 1700315010
transform 1 0 5850 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1090_
timestamp 1700315010
transform 1 0 4650 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1091_
timestamp 1700315010
transform -1 0 5670 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1092_
timestamp 1700315010
transform -1 0 6090 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1093_
timestamp 1700315010
transform 1 0 5610 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1094_
timestamp 1700315010
transform 1 0 6510 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1095_
timestamp 1700315010
transform -1 0 5550 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1096_
timestamp 1700315010
transform -1 0 5070 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1097_
timestamp 1700315010
transform -1 0 4770 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1098_
timestamp 1700315010
transform -1 0 5190 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1099_
timestamp 1700315010
transform -1 0 4290 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1100_
timestamp 1700315010
transform -1 0 150 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1101_
timestamp 1700315010
transform -1 0 150 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1102_
timestamp 1700315010
transform -1 0 2790 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1103_
timestamp 1700315010
transform 1 0 1830 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1104_
timestamp 1700315010
transform 1 0 1410 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1105_
timestamp 1700315010
transform 1 0 510 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1106_
timestamp 1700315010
transform -1 0 150 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1107_
timestamp 1700315010
transform 1 0 570 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1108_
timestamp 1700315010
transform 1 0 2610 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1109_
timestamp 1700315010
transform -1 0 1050 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1110_
timestamp 1700315010
transform -1 0 630 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1111_
timestamp 1700315010
transform -1 0 150 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1112_
timestamp 1700315010
transform -1 0 6090 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1113_
timestamp 1700315010
transform 1 0 1410 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1114_
timestamp 1700315010
transform -1 0 5310 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1115_
timestamp 1700315010
transform -1 0 1530 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1116_
timestamp 1700315010
transform -1 0 1890 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1117_
timestamp 1700315010
transform 1 0 2250 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1118_
timestamp 1700315010
transform -1 0 1050 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1119_
timestamp 1700315010
transform 1 0 1470 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1120_
timestamp 1700315010
transform 1 0 1410 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1121_
timestamp 1700315010
transform 1 0 2670 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1122_
timestamp 1700315010
transform -1 0 2250 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1123_
timestamp 1700315010
transform -1 0 1950 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1124_
timestamp 1700315010
transform 1 0 1530 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1125_
timestamp 1700315010
transform 1 0 570 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1126_
timestamp 1700315010
transform -1 0 150 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1127_
timestamp 1700315010
transform 1 0 1710 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1128_
timestamp 1700315010
transform -1 0 990 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1129_
timestamp 1700315010
transform -1 0 630 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1130_
timestamp 1700315010
transform 1 0 1050 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1131_
timestamp 1700315010
transform -1 0 1050 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1132_
timestamp 1700315010
transform -1 0 2430 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1133_
timestamp 1700315010
transform -1 0 150 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1134_
timestamp 1700315010
transform -1 0 630 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1135_
timestamp 1700315010
transform 1 0 570 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1136_
timestamp 1700315010
transform -1 0 930 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1137_
timestamp 1700315010
transform -1 0 150 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1138_
timestamp 1700315010
transform 1 0 1470 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1139_
timestamp 1700315010
transform 1 0 1770 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1140_
timestamp 1700315010
transform 1 0 5370 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1141_
timestamp 1700315010
transform 1 0 6810 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1142_
timestamp 1700315010
transform 1 0 7530 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1143_
timestamp 1700315010
transform 1 0 9930 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1144_
timestamp 1700315010
transform 1 0 10950 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1145_
timestamp 1700315010
transform 1 0 9030 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1146_
timestamp 1700315010
transform -1 0 10050 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1147_
timestamp 1700315010
transform -1 0 8730 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1148_
timestamp 1700315010
transform 1 0 9510 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1149_
timestamp 1700315010
transform -1 0 9570 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1150_
timestamp 1700315010
transform 1 0 8430 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1151_
timestamp 1700315010
transform 1 0 9990 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1152_
timestamp 1700315010
transform -1 0 9510 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1153_
timestamp 1700315010
transform 1 0 7050 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1154_
timestamp 1700315010
transform 1 0 7530 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1155_
timestamp 1700315010
transform 1 0 7950 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1156_
timestamp 1700315010
transform -1 0 7950 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1157_
timestamp 1700315010
transform -1 0 3330 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1158_
timestamp 1700315010
transform 1 0 3510 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1159_
timestamp 1700315010
transform -1 0 5190 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1160_
timestamp 1700315010
transform 1 0 1350 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1161_
timestamp 1700315010
transform 1 0 2250 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1162_
timestamp 1700315010
transform 1 0 3990 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1163_
timestamp 1700315010
transform 1 0 9930 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1164_
timestamp 1700315010
transform 1 0 11250 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1165_
timestamp 1700315010
transform -1 0 11730 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1166_
timestamp 1700315010
transform 1 0 12450 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1167_
timestamp 1700315010
transform 1 0 12870 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1168_
timestamp 1700315010
transform -1 0 10410 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1169_
timestamp 1700315010
transform 1 0 12030 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1170_
timestamp 1700315010
transform 1 0 10470 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1171_
timestamp 1700315010
transform 1 0 12150 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1172_
timestamp 1700315010
transform 1 0 11730 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1173_
timestamp 1700315010
transform 1 0 12150 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1174_
timestamp 1700315010
transform 1 0 10770 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1175_
timestamp 1700315010
transform -1 0 11310 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1176_
timestamp 1700315010
transform 1 0 10950 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1177_
timestamp 1700315010
transform -1 0 8970 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1178_
timestamp 1700315010
transform -1 0 8910 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1179_
timestamp 1700315010
transform 1 0 10050 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1180_
timestamp 1700315010
transform 1 0 6330 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1181_
timestamp 1700315010
transform 1 0 9870 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1182_
timestamp 1700315010
transform -1 0 11910 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1183_
timestamp 1700315010
transform 1 0 11370 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1184_
timestamp 1700315010
transform -1 0 10950 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1185_
timestamp 1700315010
transform -1 0 11310 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1186_
timestamp 1700315010
transform 1 0 12090 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1187_
timestamp 1700315010
transform -1 0 9990 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1188_
timestamp 1700315010
transform -1 0 13350 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1189_
timestamp 1700315010
transform 1 0 11250 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1190_
timestamp 1700315010
transform 1 0 11610 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1191_
timestamp 1700315010
transform -1 0 12630 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1192_
timestamp 1700315010
transform 1 0 13410 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1193_
timestamp 1700315010
transform 1 0 13050 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1194_
timestamp 1700315010
transform 1 0 12630 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1195_
timestamp 1700315010
transform 1 0 13410 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1196_
timestamp 1700315010
transform 1 0 11730 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1197_
timestamp 1700315010
transform -1 0 12270 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1198_
timestamp 1700315010
transform 1 0 9330 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1199_
timestamp 1700315010
transform 1 0 8370 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1200_
timestamp 1700315010
transform 1 0 10470 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1201_
timestamp 1700315010
transform -1 0 11310 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1202_
timestamp 1700315010
transform 1 0 12150 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1203_
timestamp 1700315010
transform 1 0 10590 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1204_
timestamp 1700315010
transform -1 0 11130 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1205_
timestamp 1700315010
transform 1 0 8010 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1206_
timestamp 1700315010
transform -1 0 150 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1207_
timestamp 1700315010
transform 1 0 2310 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1208_
timestamp 1700315010
transform -1 0 150 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1209_
timestamp 1700315010
transform 1 0 7110 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1210_
timestamp 1700315010
transform -1 0 4650 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1211_
timestamp 1700315010
transform -1 0 6510 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1212_
timestamp 1700315010
transform 1 0 5490 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1213_
timestamp 1700315010
transform 1 0 6270 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1214_
timestamp 1700315010
transform 1 0 6630 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1215_
timestamp 1700315010
transform -1 0 4170 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1216_
timestamp 1700315010
transform -1 0 5910 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1217_
timestamp 1700315010
transform 1 0 5970 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1218_
timestamp 1700315010
transform -1 0 5430 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1219_
timestamp 1700315010
transform 1 0 3690 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1220_
timestamp 1700315010
transform -1 0 630 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1221_
timestamp 1700315010
transform -1 0 4590 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1222_
timestamp 1700315010
transform -1 0 5730 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1223_
timestamp 1700315010
transform 1 0 5370 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1224_
timestamp 1700315010
transform -1 0 6330 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1225_
timestamp 1700315010
transform 1 0 5790 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1226_
timestamp 1700315010
transform -1 0 5010 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1227_
timestamp 1700315010
transform 1 0 4710 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1228_
timestamp 1700315010
transform 1 0 5910 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1229_
timestamp 1700315010
transform 1 0 6690 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1230_
timestamp 1700315010
transform 1 0 5550 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1231_
timestamp 1700315010
transform -1 0 5130 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1232_
timestamp 1700315010
transform 1 0 2310 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1233_
timestamp 1700315010
transform 1 0 930 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1234_
timestamp 1700315010
transform 1 0 3330 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1235_
timestamp 1700315010
transform 1 0 2790 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1236_
timestamp 1700315010
transform -1 0 870 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1237_
timestamp 1700315010
transform 1 0 1710 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1238_
timestamp 1700315010
transform 1 0 2250 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1239_
timestamp 1700315010
transform -1 0 1530 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1240_
timestamp 1700315010
transform -1 0 1290 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1241_
timestamp 1700315010
transform -1 0 690 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1242_
timestamp 1700315010
transform 1 0 1890 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1243_
timestamp 1700315010
transform 1 0 1050 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1244_
timestamp 1700315010
transform 1 0 570 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1245_
timestamp 1700315010
transform -1 0 630 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1246_
timestamp 1700315010
transform -1 0 150 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1247_
timestamp 1700315010
transform -1 0 150 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1248_
timestamp 1700315010
transform 1 0 1710 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1249_
timestamp 1700315010
transform 1 0 90 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1250_
timestamp 1700315010
transform -1 0 630 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1251_
timestamp 1700315010
transform -1 0 3330 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1252_
timestamp 1700315010
transform 1 0 1410 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1253_
timestamp 1700315010
transform 1 0 90 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1254_
timestamp 1700315010
transform -1 0 1950 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1255_
timestamp 1700315010
transform -1 0 150 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1256_
timestamp 1700315010
transform 1 0 990 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1257_
timestamp 1700315010
transform -1 0 2850 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1258_
timestamp 1700315010
transform 1 0 1050 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1259_
timestamp 1700315010
transform -1 0 2490 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1260_
timestamp 1700315010
transform -1 0 2490 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1261_
timestamp 1700315010
transform 1 0 2850 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1262_
timestamp 1700315010
transform 1 0 570 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1263_
timestamp 1700315010
transform -1 0 2070 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1264_
timestamp 1700315010
transform 1 0 1470 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1265_
timestamp 1700315010
transform -1 0 2010 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1266_
timestamp 1700315010
transform -1 0 1950 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1267_
timestamp 1700315010
transform -1 0 1110 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1268_
timestamp 1700315010
transform 1 0 3210 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1269_
timestamp 1700315010
transform 1 0 3690 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1270_
timestamp 1700315010
transform 1 0 7050 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1271_
timestamp 1700315010
transform -1 0 9270 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1272_
timestamp 1700315010
transform 1 0 14970 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1273_
timestamp 1700315010
transform -1 0 14250 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1274_
timestamp 1700315010
transform 1 0 12450 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1275_
timestamp 1700315010
transform 1 0 11850 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1276_
timestamp 1700315010
transform -1 0 13410 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1277_
timestamp 1700315010
transform 1 0 12330 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1278_
timestamp 1700315010
transform 1 0 14250 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1279_
timestamp 1700315010
transform 1 0 14130 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1280_
timestamp 1700315010
transform -1 0 10650 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1281_
timestamp 1700315010
transform -1 0 11550 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1282_
timestamp 1700315010
transform -1 0 12210 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1283_
timestamp 1700315010
transform -1 0 11070 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1284_
timestamp 1700315010
transform -1 0 4950 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1285_
timestamp 1700315010
transform -1 0 9810 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1286_
timestamp 1700315010
transform -1 0 4530 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1287_
timestamp 1700315010
transform 1 0 5670 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1288_
timestamp 1700315010
transform 1 0 8970 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1289_
timestamp 1700315010
transform 1 0 8490 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1290_
timestamp 1700315010
transform -1 0 9450 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1291_
timestamp 1700315010
transform -1 0 7170 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1292_
timestamp 1700315010
transform -1 0 6750 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1293_
timestamp 1700315010
transform -1 0 7890 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1294_
timestamp 1700315010
transform 1 0 3750 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1295_
timestamp 1700315010
transform 1 0 3330 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1296_
timestamp 1700315010
transform -1 0 4950 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1297_
timestamp 1700315010
transform 1 0 4830 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1298_
timestamp 1700315010
transform 1 0 990 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1299_
timestamp 1700315010
transform 1 0 2310 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1300_
timestamp 1700315010
transform -1 0 4830 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1301_
timestamp 1700315010
transform 1 0 6150 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1302_
timestamp 1700315010
transform -1 0 5730 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1303_
timestamp 1700315010
transform -1 0 6210 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1304_
timestamp 1700315010
transform -1 0 5250 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1305_
timestamp 1700315010
transform -1 0 4230 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1306_
timestamp 1700315010
transform 1 0 2310 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1307_
timestamp 1700315010
transform 1 0 1050 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1308_
timestamp 1700315010
transform -1 0 150 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1309_
timestamp 1700315010
transform 1 0 3930 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1310_
timestamp 1700315010
transform 1 0 4830 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1311_
timestamp 1700315010
transform 1 0 3270 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1312_
timestamp 1700315010
transform -1 0 5250 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1313_
timestamp 1700315010
transform -1 0 4050 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1314_
timestamp 1700315010
transform -1 0 3690 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1315_
timestamp 1700315010
transform 1 0 3870 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1316_
timestamp 1700315010
transform -1 0 2310 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1317_
timestamp 1700315010
transform 1 0 2850 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1318_
timestamp 1700315010
transform 1 0 8310 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1319_
timestamp 1700315010
transform -1 0 6150 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1320_
timestamp 1700315010
transform -1 0 5310 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1321_
timestamp 1700315010
transform -1 0 4830 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1322_
timestamp 1700315010
transform -1 0 3450 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1323_
timestamp 1700315010
transform -1 0 4410 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1324_
timestamp 1700315010
transform -1 0 2430 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1325_
timestamp 1700315010
transform -1 0 3030 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1326_
timestamp 1700315010
transform -1 0 2010 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1327_
timestamp 1700315010
transform -1 0 150 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1328_
timestamp 1700315010
transform -1 0 150 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1329_
timestamp 1700315010
transform 1 0 1890 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1330_
timestamp 1700315010
transform -1 0 1470 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1331_
timestamp 1700315010
transform 1 0 510 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1332_
timestamp 1700315010
transform 1 0 1410 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1333_
timestamp 1700315010
transform 1 0 2370 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1334_
timestamp 1700315010
transform 1 0 1470 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1335_
timestamp 1700315010
transform -1 0 150 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1336_
timestamp 1700315010
transform 1 0 1410 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1337_
timestamp 1700315010
transform 1 0 3330 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1338_
timestamp 1700315010
transform 1 0 90 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1339_
timestamp 1700315010
transform 1 0 2130 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1340_
timestamp 1700315010
transform 1 0 1890 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1341_
timestamp 1700315010
transform 1 0 450 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1342_
timestamp 1700315010
transform -1 0 570 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1343_
timestamp 1700315010
transform 1 0 930 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1344_
timestamp 1700315010
transform -1 0 2610 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1345_
timestamp 1700315010
transform -1 0 4470 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1346_
timestamp 1700315010
transform 1 0 2670 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1347_
timestamp 1700315010
transform 1 0 3030 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1348_
timestamp 1700315010
transform -1 0 4050 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1349_
timestamp 1700315010
transform -1 0 4170 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1350_
timestamp 1700315010
transform 1 0 1530 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1351_
timestamp 1700315010
transform 1 0 2910 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1352_
timestamp 1700315010
transform 1 0 5190 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1353_
timestamp 1700315010
transform -1 0 3570 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1354_
timestamp 1700315010
transform 1 0 5070 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1355_
timestamp 1700315010
transform -1 0 6450 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1356_
timestamp 1700315010
transform 1 0 9810 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1357_
timestamp 1700315010
transform 1 0 10290 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1358_
timestamp 1700315010
transform 1 0 10710 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1359_
timestamp 1700315010
transform 1 0 13650 0 -1 5490
box -36 -24 96 816
use FILL  FILL_1__1360_
timestamp 1700315010
transform 1 0 13470 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1361_
timestamp 1700315010
transform -1 0 12630 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1362_
timestamp 1700315010
transform 1 0 12990 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1363_
timestamp 1700315010
transform -1 0 12150 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1364_
timestamp 1700315010
transform 1 0 11670 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1365_
timestamp 1700315010
transform -1 0 14430 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1366_
timestamp 1700315010
transform -1 0 4650 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1367_
timestamp 1700315010
transform 1 0 4170 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1368_
timestamp 1700315010
transform 1 0 6270 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1369_
timestamp 1700315010
transform 1 0 8730 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1370_
timestamp 1700315010
transform 1 0 6810 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1371_
timestamp 1700315010
transform 1 0 7470 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1372_
timestamp 1700315010
transform -1 0 3810 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1373_
timestamp 1700315010
transform 1 0 2910 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1374_
timestamp 1700315010
transform -1 0 1530 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1375_
timestamp 1700315010
transform -1 0 990 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1376_
timestamp 1700315010
transform -1 0 3870 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1377_
timestamp 1700315010
transform -1 0 2610 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1378_
timestamp 1700315010
transform -1 0 3510 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1379_
timestamp 1700315010
transform -1 0 3090 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1380_
timestamp 1700315010
transform -1 0 3450 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1381_
timestamp 1700315010
transform -1 0 2970 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1382_
timestamp 1700315010
transform -1 0 2190 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1383_
timestamp 1700315010
transform -1 0 2970 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1384_
timestamp 1700315010
transform -1 0 3450 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1385_
timestamp 1700315010
transform -1 0 2490 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1386_
timestamp 1700315010
transform -1 0 690 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1387_
timestamp 1700315010
transform 1 0 1830 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1388_
timestamp 1700315010
transform 1 0 4710 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1389_
timestamp 1700315010
transform -1 0 5430 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1390_
timestamp 1700315010
transform -1 0 5010 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1391_
timestamp 1700315010
transform -1 0 4470 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1392_
timestamp 1700315010
transform 1 0 6090 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1393_
timestamp 1700315010
transform 1 0 5610 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1394_
timestamp 1700315010
transform 1 0 4110 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1395_
timestamp 1700315010
transform 1 0 1230 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1396_
timestamp 1700315010
transform -1 0 1710 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1397_
timestamp 1700315010
transform -1 0 150 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1398_
timestamp 1700315010
transform -1 0 990 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1399_
timestamp 1700315010
transform -1 0 2010 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1400_
timestamp 1700315010
transform -1 0 870 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1401_
timestamp 1700315010
transform -1 0 150 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1402_
timestamp 1700315010
transform -1 0 450 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1403_
timestamp 1700315010
transform 1 0 990 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1404_
timestamp 1700315010
transform -1 0 1470 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1405_
timestamp 1700315010
transform 1 0 990 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1406_
timestamp 1700315010
transform -1 0 150 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1407_
timestamp 1700315010
transform -1 0 150 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1408_
timestamp 1700315010
transform -1 0 1110 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1409_
timestamp 1700315010
transform -1 0 630 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1410_
timestamp 1700315010
transform 1 0 570 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1411_
timestamp 1700315010
transform -1 0 1110 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1412_
timestamp 1700315010
transform 1 0 1830 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1413_
timestamp 1700315010
transform -1 0 150 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1414_
timestamp 1700315010
transform -1 0 1890 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1415_
timestamp 1700315010
transform -1 0 3870 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1416_
timestamp 1700315010
transform 1 0 5670 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1417_
timestamp 1700315010
transform 1 0 3150 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1418_
timestamp 1700315010
transform -1 0 3630 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1419_
timestamp 1700315010
transform 1 0 4050 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1420_
timestamp 1700315010
transform -1 0 7410 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1421_
timestamp 1700315010
transform -1 0 7350 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1422_
timestamp 1700315010
transform 1 0 8310 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1423_
timestamp 1700315010
transform -1 0 7830 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1424_
timestamp 1700315010
transform 1 0 8550 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1425_
timestamp 1700315010
transform -1 0 8970 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1426_
timestamp 1700315010
transform 1 0 9330 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1427_
timestamp 1700315010
transform 1 0 13770 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1428_
timestamp 1700315010
transform -1 0 12870 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1429_
timestamp 1700315010
transform 1 0 12990 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1430_
timestamp 1700315010
transform 1 0 13470 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1431_
timestamp 1700315010
transform -1 0 14130 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1432_
timestamp 1700315010
transform 1 0 14190 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1433_
timestamp 1700315010
transform -1 0 13050 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1434_
timestamp 1700315010
transform 1 0 13890 0 1 3930
box -36 -24 96 816
use FILL  FILL_1__1435_
timestamp 1700315010
transform 1 0 17790 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1436_
timestamp 1700315010
transform -1 0 17310 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1437_
timestamp 1700315010
transform -1 0 11610 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1438_
timestamp 1700315010
transform 1 0 7950 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1439_
timestamp 1700315010
transform 1 0 3810 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1440_
timestamp 1700315010
transform -1 0 3570 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1441_
timestamp 1700315010
transform 1 0 1470 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1442_
timestamp 1700315010
transform 1 0 5430 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1443_
timestamp 1700315010
transform -1 0 6210 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1444_
timestamp 1700315010
transform -1 0 4230 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1445_
timestamp 1700315010
transform -1 0 5190 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1446_
timestamp 1700315010
transform 1 0 4590 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1447_
timestamp 1700315010
transform 1 0 5010 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1448_
timestamp 1700315010
transform 1 0 5370 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1449_
timestamp 1700315010
transform -1 0 5730 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1450_
timestamp 1700315010
transform -1 0 4650 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1451_
timestamp 1700315010
transform 1 0 4950 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1452_
timestamp 1700315010
transform 1 0 5670 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1453_
timestamp 1700315010
transform 1 0 6210 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1454_
timestamp 1700315010
transform 1 0 5730 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1455_
timestamp 1700315010
transform 1 0 8610 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1456_
timestamp 1700315010
transform -1 0 6450 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1457_
timestamp 1700315010
transform -1 0 5850 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1458_
timestamp 1700315010
transform -1 0 4830 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1459_
timestamp 1700315010
transform -1 0 1410 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1460_
timestamp 1700315010
transform 1 0 5190 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1461_
timestamp 1700315010
transform 1 0 2190 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1462_
timestamp 1700315010
transform -1 0 510 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1463_
timestamp 1700315010
transform -1 0 4290 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1464_
timestamp 1700315010
transform -1 0 2670 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1465_
timestamp 1700315010
transform -1 0 3090 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1466_
timestamp 1700315010
transform -1 0 1770 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1467_
timestamp 1700315010
transform -1 0 3930 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1468_
timestamp 1700315010
transform 1 0 4290 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1469_
timestamp 1700315010
transform -1 0 3330 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1470_
timestamp 1700315010
transform -1 0 2670 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1471_
timestamp 1700315010
transform 1 0 2310 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1472_
timestamp 1700315010
transform 1 0 2790 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1473_
timestamp 1700315010
transform 1 0 3690 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1474_
timestamp 1700315010
transform 1 0 8310 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1475_
timestamp 1700315010
transform 1 0 8190 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1476_
timestamp 1700315010
transform 1 0 8910 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1477_
timestamp 1700315010
transform 1 0 9390 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1478_
timestamp 1700315010
transform 1 0 9690 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1479_
timestamp 1700315010
transform 1 0 10530 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1480_
timestamp 1700315010
transform -1 0 12690 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1481_
timestamp 1700315010
transform -1 0 13050 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1482_
timestamp 1700315010
transform 1 0 13890 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1483_
timestamp 1700315010
transform 1 0 16110 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1484_
timestamp 1700315010
transform -1 0 16530 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1485_
timestamp 1700315010
transform 1 0 16470 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1486_
timestamp 1700315010
transform -1 0 17010 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1487_
timestamp 1700315010
transform 1 0 17430 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1488_
timestamp 1700315010
transform 1 0 6510 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1489_
timestamp 1700315010
transform 1 0 6990 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1490_
timestamp 1700315010
transform -1 0 7050 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1491_
timestamp 1700315010
transform -1 0 8610 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1492_
timestamp 1700315010
transform -1 0 6330 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1493_
timestamp 1700315010
transform -1 0 6750 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1494_
timestamp 1700315010
transform 1 0 7650 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1495_
timestamp 1700315010
transform 1 0 8910 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1496_
timestamp 1700315010
transform 1 0 7170 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1497_
timestamp 1700315010
transform 1 0 7770 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1498_
timestamp 1700315010
transform 1 0 8190 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1499_
timestamp 1700315010
transform 1 0 6630 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1500_
timestamp 1700315010
transform 1 0 7290 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1501_
timestamp 1700315010
transform 1 0 8130 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1502_
timestamp 1700315010
transform 1 0 8190 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1503_
timestamp 1700315010
transform 1 0 8310 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1504_
timestamp 1700315010
transform 1 0 8550 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1505_
timestamp 1700315010
transform -1 0 7350 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1506_
timestamp 1700315010
transform -1 0 7890 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1507_
timestamp 1700315010
transform -1 0 7410 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1508_
timestamp 1700315010
transform -1 0 6630 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1509_
timestamp 1700315010
transform 1 0 6090 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1510_
timestamp 1700315010
transform -1 0 5730 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1511_
timestamp 1700315010
transform 1 0 6930 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1512_
timestamp 1700315010
transform -1 0 8130 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1513_
timestamp 1700315010
transform 1 0 9930 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1514_
timestamp 1700315010
transform -1 0 9150 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1515_
timestamp 1700315010
transform 1 0 9450 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1516_
timestamp 1700315010
transform -1 0 7590 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1517_
timestamp 1700315010
transform 1 0 8610 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1518_
timestamp 1700315010
transform -1 0 9630 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1519_
timestamp 1700315010
transform 1 0 8730 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1520_
timestamp 1700315010
transform 1 0 9150 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1521_
timestamp 1700315010
transform 1 0 7650 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1522_
timestamp 1700315010
transform 1 0 8130 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1523_
timestamp 1700315010
transform 1 0 8490 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1524_
timestamp 1700315010
transform 1 0 9870 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1525_
timestamp 1700315010
transform -1 0 16410 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1526_
timestamp 1700315010
transform -1 0 14910 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1527_
timestamp 1700315010
transform 1 0 13410 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1528_
timestamp 1700315010
transform 1 0 12930 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1529_
timestamp 1700315010
transform 1 0 13710 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1530_
timestamp 1700315010
transform -1 0 14550 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1531_
timestamp 1700315010
transform -1 0 15210 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1532_
timestamp 1700315010
transform 1 0 15630 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1533_
timestamp 1700315010
transform -1 0 16050 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1534_
timestamp 1700315010
transform -1 0 15450 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1535_
timestamp 1700315010
transform -1 0 11250 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1536_
timestamp 1700315010
transform 1 0 9510 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1537_
timestamp 1700315010
transform 1 0 8370 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1538_
timestamp 1700315010
transform 1 0 7710 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1539_
timestamp 1700315010
transform 1 0 6870 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1540_
timestamp 1700315010
transform -1 0 7890 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1541_
timestamp 1700315010
transform -1 0 8370 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1542_
timestamp 1700315010
transform -1 0 7410 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1543_
timestamp 1700315010
transform 1 0 7890 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1544_
timestamp 1700315010
transform 1 0 7290 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1545_
timestamp 1700315010
transform -1 0 7410 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1546_
timestamp 1700315010
transform -1 0 7470 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1547_
timestamp 1700315010
transform -1 0 8010 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1548_
timestamp 1700315010
transform -1 0 9090 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1549_
timestamp 1700315010
transform -1 0 8430 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1550_
timestamp 1700315010
transform 1 0 10350 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1551_
timestamp 1700315010
transform 1 0 11670 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1552_
timestamp 1700315010
transform 1 0 12510 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1553_
timestamp 1700315010
transform -1 0 15150 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1554_
timestamp 1700315010
transform 1 0 15630 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1555_
timestamp 1700315010
transform 1 0 15570 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1556_
timestamp 1700315010
transform -1 0 14910 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1557_
timestamp 1700315010
transform -1 0 14550 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1558_
timestamp 1700315010
transform 1 0 7530 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1559_
timestamp 1700315010
transform 1 0 10530 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1560_
timestamp 1700315010
transform 1 0 10890 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1561_
timestamp 1700315010
transform -1 0 8070 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1562_
timestamp 1700315010
transform 1 0 8010 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1563_
timestamp 1700315010
transform 1 0 11070 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1564_
timestamp 1700315010
transform -1 0 6150 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1565_
timestamp 1700315010
transform -1 0 6450 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1566_
timestamp 1700315010
transform -1 0 6870 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1567_
timestamp 1700315010
transform 1 0 8670 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1568_
timestamp 1700315010
transform 1 0 9930 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1569_
timestamp 1700315010
transform 1 0 11790 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1570_
timestamp 1700315010
transform 1 0 10050 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1571_
timestamp 1700315010
transform -1 0 10830 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1572_
timestamp 1700315010
transform 1 0 10290 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1573_
timestamp 1700315010
transform 1 0 12270 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1574_
timestamp 1700315010
transform -1 0 12150 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1575_
timestamp 1700315010
transform 1 0 12930 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1576_
timestamp 1700315010
transform 1 0 12450 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1577_
timestamp 1700315010
transform 1 0 13350 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1578_
timestamp 1700315010
transform 1 0 17070 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1579_
timestamp 1700315010
transform -1 0 15330 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1580_
timestamp 1700315010
transform -1 0 15210 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1581_
timestamp 1700315010
transform 1 0 14610 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1582_
timestamp 1700315010
transform -1 0 13470 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1583_
timestamp 1700315010
transform -1 0 11430 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1584_
timestamp 1700315010
transform 1 0 8790 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1585_
timestamp 1700315010
transform 1 0 9270 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1586_
timestamp 1700315010
transform 1 0 10830 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1587_
timestamp 1700315010
transform 1 0 7590 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1588_
timestamp 1700315010
transform -1 0 11550 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1589_
timestamp 1700315010
transform 1 0 14790 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1590_
timestamp 1700315010
transform 1 0 14310 0 1 2370
box -36 -24 96 816
use FILL  FILL_1__1591_
timestamp 1700315010
transform -1 0 14190 0 -1 2370
box -36 -24 96 816
use FILL  FILL_1__1592_
timestamp 1700315010
transform -1 0 12990 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1593_
timestamp 1700315010
transform -1 0 12990 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1__1594_
timestamp 1700315010
transform 1 0 12870 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1595_
timestamp 1700315010
transform 1 0 11910 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1596_
timestamp 1700315010
transform -1 0 12390 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1597_
timestamp 1700315010
transform 1 0 11970 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1598_
timestamp 1700315010
transform -1 0 12450 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1599_
timestamp 1700315010
transform -1 0 11670 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1600_
timestamp 1700315010
transform -1 0 12030 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1601_
timestamp 1700315010
transform 1 0 9870 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1602_
timestamp 1700315010
transform -1 0 9990 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1603_
timestamp 1700315010
transform 1 0 8790 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1604_
timestamp 1700315010
transform -1 0 9270 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1605_
timestamp 1700315010
transform -1 0 13410 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1606_
timestamp 1700315010
transform -1 0 15450 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1607_
timestamp 1700315010
transform 1 0 13230 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1608_
timestamp 1700315010
transform -1 0 13710 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1636_
timestamp 1700315010
transform -1 0 17670 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1637_
timestamp 1700315010
transform 1 0 17670 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1638_
timestamp 1700315010
transform -1 0 16050 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1639_
timestamp 1700315010
transform 1 0 15570 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1640_
timestamp 1700315010
transform 1 0 15570 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1641_
timestamp 1700315010
transform -1 0 11250 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1642_
timestamp 1700315010
transform -1 0 9450 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1643_
timestamp 1700315010
transform -1 0 8970 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1644_
timestamp 1700315010
transform -1 0 11550 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1645_
timestamp 1700315010
transform -1 0 13170 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1646_
timestamp 1700315010
transform -1 0 12270 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1647_
timestamp 1700315010
transform 1 0 9450 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1648_
timestamp 1700315010
transform 1 0 17310 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1649_
timestamp 1700315010
transform -1 0 12810 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1650_
timestamp 1700315010
transform -1 0 13290 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1651_
timestamp 1700315010
transform 1 0 12870 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1652_
timestamp 1700315010
transform -1 0 10830 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1653_
timestamp 1700315010
transform 1 0 12390 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1654_
timestamp 1700315010
transform 1 0 17370 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1655_
timestamp 1700315010
transform -1 0 16950 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1656_
timestamp 1700315010
transform 1 0 17730 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1657_
timestamp 1700315010
transform 1 0 17310 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1658_
timestamp 1700315010
transform 1 0 16830 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1659_
timestamp 1700315010
transform -1 0 15990 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1660_
timestamp 1700315010
transform -1 0 16530 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1661_
timestamp 1700315010
transform 1 0 15990 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1662_
timestamp 1700315010
transform -1 0 10350 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1663_
timestamp 1700315010
transform -1 0 9870 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1664_
timestamp 1700315010
transform -1 0 10290 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1665_
timestamp 1700315010
transform -1 0 10890 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1666_
timestamp 1700315010
transform -1 0 11430 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1667_
timestamp 1700315010
transform 1 0 11490 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1668_
timestamp 1700315010
transform 1 0 11070 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1669_
timestamp 1700315010
transform -1 0 12090 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1670_
timestamp 1700315010
transform 1 0 12510 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1671_
timestamp 1700315010
transform 1 0 15630 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1672_
timestamp 1700315010
transform -1 0 16950 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1673_
timestamp 1700315010
transform 1 0 16410 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1674_
timestamp 1700315010
transform -1 0 16050 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1675_
timestamp 1700315010
transform -1 0 16590 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1676_
timestamp 1700315010
transform 1 0 16410 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1677_
timestamp 1700315010
transform -1 0 14610 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1678_
timestamp 1700315010
transform -1 0 14730 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1679_
timestamp 1700315010
transform -1 0 13530 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1680_
timestamp 1700315010
transform 1 0 13830 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1681_
timestamp 1700315010
transform -1 0 11970 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1682_
timestamp 1700315010
transform 1 0 13710 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1683_
timestamp 1700315010
transform 1 0 14070 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1684_
timestamp 1700315010
transform 1 0 15030 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1685_
timestamp 1700315010
transform -1 0 12510 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1686_
timestamp 1700315010
transform 1 0 12870 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1687_
timestamp 1700315010
transform -1 0 15270 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1688_
timestamp 1700315010
transform 1 0 15630 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1689_
timestamp 1700315010
transform 1 0 14610 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1690_
timestamp 1700315010
transform 1 0 15210 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1691_
timestamp 1700315010
transform -1 0 14790 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1692_
timestamp 1700315010
transform 1 0 10710 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1693_
timestamp 1700315010
transform 1 0 9270 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1694_
timestamp 1700315010
transform -1 0 9810 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1695_
timestamp 1700315010
transform -1 0 8790 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1696_
timestamp 1700315010
transform -1 0 9090 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1697_
timestamp 1700315010
transform -1 0 9870 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1698_
timestamp 1700315010
transform 1 0 10290 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1699_
timestamp 1700315010
transform -1 0 11610 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1700_
timestamp 1700315010
transform -1 0 11670 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1701_
timestamp 1700315010
transform -1 0 10770 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1702_
timestamp 1700315010
transform 1 0 11130 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1703_
timestamp 1700315010
transform -1 0 13710 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1704_
timestamp 1700315010
transform -1 0 14370 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1705_
timestamp 1700315010
transform 1 0 12090 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1706_
timestamp 1700315010
transform -1 0 12990 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1707_
timestamp 1700315010
transform -1 0 13410 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1708_
timestamp 1700315010
transform 1 0 13410 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1709_
timestamp 1700315010
transform -1 0 10950 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1710_
timestamp 1700315010
transform -1 0 11610 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1711_
timestamp 1700315010
transform -1 0 10650 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1712_
timestamp 1700315010
transform -1 0 11070 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1713_
timestamp 1700315010
transform -1 0 10170 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1714_
timestamp 1700315010
transform 1 0 11310 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1715_
timestamp 1700315010
transform -1 0 11790 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1716_
timestamp 1700315010
transform 1 0 12210 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1717_
timestamp 1700315010
transform -1 0 13290 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1718_
timestamp 1700315010
transform 1 0 13650 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1719_
timestamp 1700315010
transform 1 0 14130 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1720_
timestamp 1700315010
transform 1 0 12690 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1721_
timestamp 1700315010
transform 1 0 13950 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1722_
timestamp 1700315010
transform 1 0 14250 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1723_
timestamp 1700315010
transform 1 0 14370 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1__1724_
timestamp 1700315010
transform -1 0 14370 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1725_
timestamp 1700315010
transform 1 0 13230 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1726_
timestamp 1700315010
transform -1 0 12810 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1727_
timestamp 1700315010
transform -1 0 13110 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1728_
timestamp 1700315010
transform -1 0 9030 0 1 16410
box -36 -24 96 816
use FILL  FILL_1__1729_
timestamp 1700315010
transform 1 0 9210 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1730_
timestamp 1700315010
transform -1 0 9690 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1731_
timestamp 1700315010
transform -1 0 10110 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1732_
timestamp 1700315010
transform 1 0 10590 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1733_
timestamp 1700315010
transform 1 0 11010 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1734_
timestamp 1700315010
transform 1 0 14850 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1735_
timestamp 1700315010
transform 1 0 14730 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1736_
timestamp 1700315010
transform -1 0 15690 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1737_
timestamp 1700315010
transform 1 0 15150 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1738_
timestamp 1700315010
transform 1 0 15270 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1739_
timestamp 1700315010
transform 1 0 14730 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1740_
timestamp 1700315010
transform -1 0 15450 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1741_
timestamp 1700315010
transform 1 0 15630 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1742_
timestamp 1700315010
transform 1 0 10530 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1743_
timestamp 1700315010
transform -1 0 8310 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1744_
timestamp 1700315010
transform -1 0 8790 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1745_
timestamp 1700315010
transform -1 0 9690 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1746_
timestamp 1700315010
transform 1 0 9150 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1747_
timestamp 1700315010
transform 1 0 10050 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1748_
timestamp 1700315010
transform -1 0 15270 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1749_
timestamp 1700315010
transform 1 0 15630 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1750_
timestamp 1700315010
transform 1 0 16290 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1751_
timestamp 1700315010
transform 1 0 16110 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1752_
timestamp 1700315010
transform -1 0 15810 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1753_
timestamp 1700315010
transform 1 0 16110 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1754_
timestamp 1700315010
transform 1 0 15450 0 1 5490
box -36 -24 96 816
use FILL  FILL_1__1755_
timestamp 1700315010
transform 1 0 16110 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1756_
timestamp 1700315010
transform 1 0 14490 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1757_
timestamp 1700315010
transform -1 0 13170 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1758_
timestamp 1700315010
transform 1 0 12690 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1759_
timestamp 1700315010
transform 1 0 11970 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1760_
timestamp 1700315010
transform 1 0 13530 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1761_
timestamp 1700315010
transform -1 0 14070 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1762_
timestamp 1700315010
transform -1 0 15390 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1763_
timestamp 1700315010
transform 1 0 15810 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1764_
timestamp 1700315010
transform 1 0 16770 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1765_
timestamp 1700315010
transform 1 0 17190 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1766_
timestamp 1700315010
transform 1 0 17490 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1767_
timestamp 1700315010
transform 1 0 14670 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1768_
timestamp 1700315010
transform -1 0 14250 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1769_
timestamp 1700315010
transform -1 0 13770 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1770_
timestamp 1700315010
transform -1 0 15030 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1771_
timestamp 1700315010
transform 1 0 16530 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1772_
timestamp 1700315010
transform 1 0 16590 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1773_
timestamp 1700315010
transform -1 0 17430 0 1 17970
box -36 -24 96 816
use FILL  FILL_1__1774_
timestamp 1700315010
transform -1 0 16770 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1775_
timestamp 1700315010
transform -1 0 17130 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1776_
timestamp 1700315010
transform 1 0 17130 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1777_
timestamp 1700315010
transform 1 0 14790 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1778_
timestamp 1700315010
transform 1 0 13410 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1779_
timestamp 1700315010
transform 1 0 13050 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1780_
timestamp 1700315010
transform 1 0 12510 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1781_
timestamp 1700315010
transform 1 0 13890 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1782_
timestamp 1700315010
transform 1 0 14370 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1783_
timestamp 1700315010
transform 1 0 16830 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1784_
timestamp 1700315010
transform 1 0 16410 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1785_
timestamp 1700315010
transform -1 0 17430 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1786_
timestamp 1700315010
transform 1 0 17850 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1787_
timestamp 1700315010
transform -1 0 17670 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1788_
timestamp 1700315010
transform 1 0 17130 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1789_
timestamp 1700315010
transform 1 0 17970 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1790_
timestamp 1700315010
transform 1 0 17970 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1791_
timestamp 1700315010
transform 1 0 17910 0 1 7050
box -36 -24 96 816
use FILL  FILL_1__1792_
timestamp 1700315010
transform 1 0 13950 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1793_
timestamp 1700315010
transform 1 0 13530 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1794_
timestamp 1700315010
transform 1 0 14610 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1795_
timestamp 1700315010
transform -1 0 16710 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1796_
timestamp 1700315010
transform 1 0 16230 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1797_
timestamp 1700315010
transform -1 0 15090 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1798_
timestamp 1700315010
transform -1 0 17610 0 1 11730
box -36 -24 96 816
use FILL  FILL_1__1799_
timestamp 1700315010
transform -1 0 17610 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1__1800_
timestamp 1700315010
transform -1 0 17550 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1801_
timestamp 1700315010
transform 1 0 16230 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1802_
timestamp 1700315010
transform 1 0 14250 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1__1803_
timestamp 1700315010
transform 1 0 17610 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1804_
timestamp 1700315010
transform -1 0 17670 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1805_
timestamp 1700315010
transform 1 0 17970 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1806_
timestamp 1700315010
transform -1 0 17070 0 1 13290
box -36 -24 96 816
use FILL  FILL_1__1807_
timestamp 1700315010
transform 1 0 17010 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1808_
timestamp 1700315010
transform 1 0 16590 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1809_
timestamp 1700315010
transform 1 0 16890 0 1 14850
box -36 -24 96 816
use FILL  FILL_1__1810_
timestamp 1700315010
transform 1 0 17670 0 -1 14850
box -36 -24 96 816
use FILL  FILL_1__1811_
timestamp 1700315010
transform 1 0 17190 0 1 810
box -36 -24 96 816
use FILL  FILL_1__1812_
timestamp 1700315010
transform 1 0 17910 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1__1813_
timestamp 1700315010
transform -1 0 17970 0 1 10170
box -36 -24 96 816
use FILL  FILL_1__1814_
timestamp 1700315010
transform -1 0 18030 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1815_
timestamp 1700315010
transform 1 0 17490 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1__1816_
timestamp 1700315010
transform -1 0 17970 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1817_
timestamp 1700315010
transform -1 0 17610 0 1 8610
box -36 -24 96 816
use FILL  FILL_1__1818_
timestamp 1700315010
transform -1 0 9810 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1819_
timestamp 1700315010
transform -1 0 7770 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1__1820_
timestamp 1700315010
transform -1 0 13830 0 -1 3930
box -36 -24 96 816
use FILL  FILL_1__1821_
timestamp 1700315010
transform -1 0 16890 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1822_
timestamp 1700315010
transform 1 0 16410 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1823_
timestamp 1700315010
transform 1 0 16050 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1824_
timestamp 1700315010
transform 1 0 14910 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1825_
timestamp 1700315010
transform 1 0 13770 0 -1 810
box -36 -24 96 816
use FILL  FILL_1__1826_
timestamp 1700315010
transform 1 0 17250 0 -1 810
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert0
timestamp 1700315010
transform 1 0 11790 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert1
timestamp 1700315010
transform -1 0 6630 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert2
timestamp 1700315010
transform -1 0 6990 0 1 7050
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert3
timestamp 1700315010
transform -1 0 6810 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert4
timestamp 1700315010
transform -1 0 13230 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert5
timestamp 1700315010
transform -1 0 11310 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert6
timestamp 1700315010
transform -1 0 8190 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert7
timestamp 1700315010
transform -1 0 10230 0 -1 7050
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert13
timestamp 1700315010
transform 1 0 15570 0 1 8610
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert14
timestamp 1700315010
transform -1 0 11490 0 1 10170
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert15
timestamp 1700315010
transform -1 0 13050 0 1 10170
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert16
timestamp 1700315010
transform -1 0 12090 0 -1 8610
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert17
timestamp 1700315010
transform 1 0 7590 0 1 11730
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert18
timestamp 1700315010
transform -1 0 7050 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert19
timestamp 1700315010
transform 1 0 9090 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert20
timestamp 1700315010
transform -1 0 7290 0 1 8610
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert21
timestamp 1700315010
transform 1 0 15990 0 1 8610
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert22
timestamp 1700315010
transform -1 0 12630 0 1 10170
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert23
timestamp 1700315010
transform 1 0 12750 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert24
timestamp 1700315010
transform 1 0 15870 0 -1 10170
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert25
timestamp 1700315010
transform -1 0 7050 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert26
timestamp 1700315010
transform -1 0 7950 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert27
timestamp 1700315010
transform -1 0 7230 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert28
timestamp 1700315010
transform 1 0 9510 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert29
timestamp 1700315010
transform -1 0 6570 0 1 7050
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert30
timestamp 1700315010
transform 1 0 10170 0 1 7050
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert31
timestamp 1700315010
transform -1 0 6630 0 -1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert32
timestamp 1700315010
transform 1 0 10530 0 1 13290
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert33
timestamp 1700315010
transform -1 0 15270 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert34
timestamp 1700315010
transform -1 0 18030 0 -1 16410
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert35
timestamp 1700315010
transform -1 0 14850 0 -1 17970
box -36 -24 96 816
use FILL  FILL_1_BUFX2_insert36
timestamp 1700315010
transform -1 0 17850 0 1 16410
box -36 -24 96 816
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1700315010
transform -1 0 13650 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 14850 0 1 8610
box -36 -24 96 816
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 17430 0 1 2370
box -36 -24 96 816
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1700315010
transform -1 0 15570 0 -1 11730
box -36 -24 96 816
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 14910 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__889_
timestamp 1700315010
transform 1 0 16110 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__890_
timestamp 1700315010
transform -1 0 14970 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__892_
timestamp 1700315010
transform 1 0 16170 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__893_
timestamp 1700315010
transform -1 0 15750 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__894_
timestamp 1700315010
transform 1 0 16530 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__896_
timestamp 1700315010
transform -1 0 15390 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__897_
timestamp 1700315010
transform 1 0 15390 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__899_
timestamp 1700315010
transform 1 0 15810 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__900_
timestamp 1700315010
transform -1 0 17610 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__902_
timestamp 1700315010
transform 1 0 17430 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__903_
timestamp 1700315010
transform 1 0 14730 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__905_
timestamp 1700315010
transform -1 0 17130 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__906_
timestamp 1700315010
transform -1 0 12690 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__908_
timestamp 1700315010
transform 1 0 17910 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__909_
timestamp 1700315010
transform 1 0 16830 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__911_
timestamp 1700315010
transform 1 0 16290 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__912_
timestamp 1700315010
transform 1 0 17310 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__914_
timestamp 1700315010
transform -1 0 15810 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__915_
timestamp 1700315010
transform 1 0 15750 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__916_
timestamp 1700315010
transform -1 0 16950 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__918_
timestamp 1700315010
transform -1 0 16230 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__919_
timestamp 1700315010
transform 1 0 16230 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__921_
timestamp 1700315010
transform 1 0 17010 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__922_
timestamp 1700315010
transform 1 0 16170 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__924_
timestamp 1700315010
transform 1 0 17730 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__925_
timestamp 1700315010
transform -1 0 17970 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__927_
timestamp 1700315010
transform 1 0 14610 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__928_
timestamp 1700315010
transform 1 0 14130 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__930_
timestamp 1700315010
transform 1 0 11070 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__931_
timestamp 1700315010
transform -1 0 11550 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__933_
timestamp 1700315010
transform -1 0 13290 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__934_
timestamp 1700315010
transform 1 0 13650 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__936_
timestamp 1700315010
transform 1 0 12270 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__937_
timestamp 1700315010
transform -1 0 12030 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__939_
timestamp 1700315010
transform 1 0 11010 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__940_
timestamp 1700315010
transform 1 0 10410 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__941_
timestamp 1700315010
transform -1 0 9810 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__943_
timestamp 1700315010
transform 1 0 10470 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__944_
timestamp 1700315010
transform -1 0 15990 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__946_
timestamp 1700315010
transform 1 0 16290 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__947_
timestamp 1700315010
transform 1 0 17010 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__949_
timestamp 1700315010
transform 1 0 15330 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__950_
timestamp 1700315010
transform -1 0 14010 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__952_
timestamp 1700315010
transform 1 0 7050 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__953_
timestamp 1700315010
transform 1 0 7950 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__955_
timestamp 1700315010
transform 1 0 8310 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__956_
timestamp 1700315010
transform 1 0 9570 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__958_
timestamp 1700315010
transform 1 0 10890 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__959_
timestamp 1700315010
transform 1 0 10890 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__961_
timestamp 1700315010
transform -1 0 10470 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__962_
timestamp 1700315010
transform 1 0 11370 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__963_
timestamp 1700315010
transform 1 0 8790 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__965_
timestamp 1700315010
transform 1 0 7530 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__966_
timestamp 1700315010
transform 1 0 10050 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__968_
timestamp 1700315010
transform 1 0 7770 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__969_
timestamp 1700315010
transform -1 0 8370 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__971_
timestamp 1700315010
transform 1 0 9150 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__972_
timestamp 1700315010
transform -1 0 9630 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__974_
timestamp 1700315010
transform -1 0 10530 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__975_
timestamp 1700315010
transform 1 0 9210 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__977_
timestamp 1700315010
transform 1 0 6390 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__978_
timestamp 1700315010
transform 1 0 7530 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__980_
timestamp 1700315010
transform 1 0 8730 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__981_
timestamp 1700315010
transform 1 0 10950 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__983_
timestamp 1700315010
transform -1 0 8310 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__984_
timestamp 1700315010
transform -1 0 7350 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__985_
timestamp 1700315010
transform -1 0 7110 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__987_
timestamp 1700315010
transform -1 0 4830 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__988_
timestamp 1700315010
transform -1 0 4170 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__990_
timestamp 1700315010
transform 1 0 5610 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__991_
timestamp 1700315010
transform 1 0 7230 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__993_
timestamp 1700315010
transform 1 0 6090 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__994_
timestamp 1700315010
transform 1 0 7830 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__996_
timestamp 1700315010
transform 1 0 5130 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__997_
timestamp 1700315010
transform -1 0 4350 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__999_
timestamp 1700315010
transform 1 0 6630 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1001_
timestamp 1700315010
transform 1 0 8370 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1002_
timestamp 1700315010
transform 1 0 7050 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1004_
timestamp 1700315010
transform 1 0 7470 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1005_
timestamp 1700315010
transform -1 0 7050 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1007_
timestamp 1700315010
transform -1 0 5070 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1008_
timestamp 1700315010
transform 1 0 5370 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1009_
timestamp 1700315010
transform -1 0 5910 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1011_
timestamp 1700315010
transform -1 0 6690 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1012_
timestamp 1700315010
transform -1 0 4470 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1014_
timestamp 1700315010
transform -1 0 6630 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1015_
timestamp 1700315010
transform -1 0 6210 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1017_
timestamp 1700315010
transform 1 0 6630 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1018_
timestamp 1700315010
transform -1 0 7170 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1020_
timestamp 1700315010
transform -1 0 4590 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1021_
timestamp 1700315010
transform -1 0 4350 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1023_
timestamp 1700315010
transform 1 0 3450 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1024_
timestamp 1700315010
transform 1 0 4530 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1026_
timestamp 1700315010
transform 1 0 3810 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1027_
timestamp 1700315010
transform 1 0 4530 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1029_
timestamp 1700315010
transform -1 0 2790 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1030_
timestamp 1700315010
transform -1 0 4830 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1032_
timestamp 1700315010
transform -1 0 3750 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1033_
timestamp 1700315010
transform -1 0 3270 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1034_
timestamp 1700315010
transform -1 0 5010 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1036_
timestamp 1700315010
transform -1 0 3570 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1037_
timestamp 1700315010
transform -1 0 3210 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1039_
timestamp 1700315010
transform -1 0 4050 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1040_
timestamp 1700315010
transform -1 0 6210 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1042_
timestamp 1700315010
transform 1 0 5730 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1043_
timestamp 1700315010
transform 1 0 6930 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1045_
timestamp 1700315010
transform 1 0 6330 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1046_
timestamp 1700315010
transform -1 0 4890 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1048_
timestamp 1700315010
transform -1 0 5910 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1049_
timestamp 1700315010
transform -1 0 4410 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1051_
timestamp 1700315010
transform -1 0 2130 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1052_
timestamp 1700315010
transform 1 0 3630 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1054_
timestamp 1700315010
transform -1 0 4170 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1055_
timestamp 1700315010
transform -1 0 2910 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1056_
timestamp 1700315010
transform 1 0 3030 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1058_
timestamp 1700315010
transform 1 0 3810 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1059_
timestamp 1700315010
transform 1 0 3330 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1061_
timestamp 1700315010
transform -1 0 8850 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1062_
timestamp 1700315010
transform -1 0 5790 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1064_
timestamp 1700315010
transform 1 0 4170 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1065_
timestamp 1700315010
transform -1 0 2850 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1067_
timestamp 1700315010
transform 1 0 3930 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1068_
timestamp 1700315010
transform -1 0 2610 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1070_
timestamp 1700315010
transform 1 0 5910 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1071_
timestamp 1700315010
transform 1 0 4770 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1073_
timestamp 1700315010
transform -1 0 2910 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1074_
timestamp 1700315010
transform -1 0 2430 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1076_
timestamp 1700315010
transform -1 0 2970 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1077_
timestamp 1700315010
transform 1 0 3390 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1079_
timestamp 1700315010
transform -1 0 2730 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1080_
timestamp 1700315010
transform -1 0 2610 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1081_
timestamp 1700315010
transform -1 0 690 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1083_
timestamp 1700315010
transform -1 0 2310 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1084_
timestamp 1700315010
transform -1 0 1170 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1086_
timestamp 1700315010
transform 1 0 2070 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1087_
timestamp 1700315010
transform 1 0 1590 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1089_
timestamp 1700315010
transform 1 0 5910 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1090_
timestamp 1700315010
transform 1 0 4710 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1092_
timestamp 1700315010
transform -1 0 6150 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1093_
timestamp 1700315010
transform 1 0 5670 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1095_
timestamp 1700315010
transform -1 0 5610 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1096_
timestamp 1700315010
transform -1 0 5130 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1098_
timestamp 1700315010
transform -1 0 5250 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1099_
timestamp 1700315010
transform -1 0 4350 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1101_
timestamp 1700315010
transform -1 0 210 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1102_
timestamp 1700315010
transform -1 0 2850 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1103_
timestamp 1700315010
transform 1 0 1890 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1105_
timestamp 1700315010
transform 1 0 570 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1106_
timestamp 1700315010
transform -1 0 210 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1108_
timestamp 1700315010
transform 1 0 2670 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1109_
timestamp 1700315010
transform -1 0 1110 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1111_
timestamp 1700315010
transform -1 0 210 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1112_
timestamp 1700315010
transform -1 0 6150 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1114_
timestamp 1700315010
transform -1 0 5370 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1115_
timestamp 1700315010
transform -1 0 1590 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1117_
timestamp 1700315010
transform 1 0 2310 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1118_
timestamp 1700315010
transform -1 0 1110 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1120_
timestamp 1700315010
transform 1 0 1470 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1121_
timestamp 1700315010
transform 1 0 2730 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1123_
timestamp 1700315010
transform -1 0 2010 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1124_
timestamp 1700315010
transform 1 0 1590 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1126_
timestamp 1700315010
transform -1 0 210 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1127_
timestamp 1700315010
transform 1 0 1770 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1128_
timestamp 1700315010
transform -1 0 1050 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1130_
timestamp 1700315010
transform 1 0 1110 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1131_
timestamp 1700315010
transform -1 0 1110 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1133_
timestamp 1700315010
transform -1 0 210 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1134_
timestamp 1700315010
transform -1 0 690 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1136_
timestamp 1700315010
transform -1 0 990 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1137_
timestamp 1700315010
transform -1 0 210 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1139_
timestamp 1700315010
transform 1 0 1830 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1140_
timestamp 1700315010
transform 1 0 5430 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1142_
timestamp 1700315010
transform 1 0 7590 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1143_
timestamp 1700315010
transform 1 0 9990 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1145_
timestamp 1700315010
transform 1 0 9090 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1146_
timestamp 1700315010
transform -1 0 10110 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1148_
timestamp 1700315010
transform 1 0 9570 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1149_
timestamp 1700315010
transform -1 0 9630 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1150_
timestamp 1700315010
transform 1 0 8490 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1152_
timestamp 1700315010
transform -1 0 9570 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1153_
timestamp 1700315010
transform 1 0 7110 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1155_
timestamp 1700315010
transform 1 0 8010 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1156_
timestamp 1700315010
transform -1 0 8010 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1158_
timestamp 1700315010
transform 1 0 3570 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1159_
timestamp 1700315010
transform -1 0 5250 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1161_
timestamp 1700315010
transform 1 0 2310 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1162_
timestamp 1700315010
transform 1 0 4050 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1164_
timestamp 1700315010
transform 1 0 11310 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1165_
timestamp 1700315010
transform -1 0 11790 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1167_
timestamp 1700315010
transform 1 0 12930 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1168_
timestamp 1700315010
transform -1 0 10470 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1170_
timestamp 1700315010
transform 1 0 10530 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1171_
timestamp 1700315010
transform 1 0 12210 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1173_
timestamp 1700315010
transform 1 0 12210 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1174_
timestamp 1700315010
transform 1 0 10830 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1175_
timestamp 1700315010
transform -1 0 11370 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1177_
timestamp 1700315010
transform -1 0 9030 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1178_
timestamp 1700315010
transform -1 0 8970 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1180_
timestamp 1700315010
transform 1 0 6390 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1181_
timestamp 1700315010
transform 1 0 9930 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1183_
timestamp 1700315010
transform 1 0 11430 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1184_
timestamp 1700315010
transform -1 0 11010 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1186_
timestamp 1700315010
transform 1 0 12150 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1187_
timestamp 1700315010
transform -1 0 10050 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1189_
timestamp 1700315010
transform 1 0 11310 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1190_
timestamp 1700315010
transform 1 0 11670 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1192_
timestamp 1700315010
transform 1 0 13470 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1193_
timestamp 1700315010
transform 1 0 13110 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1195_
timestamp 1700315010
transform 1 0 13470 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1196_
timestamp 1700315010
transform 1 0 11790 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1197_
timestamp 1700315010
transform -1 0 12330 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1199_
timestamp 1700315010
transform 1 0 8430 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1200_
timestamp 1700315010
transform 1 0 10530 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1202_
timestamp 1700315010
transform 1 0 12210 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1203_
timestamp 1700315010
transform 1 0 10650 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1205_
timestamp 1700315010
transform 1 0 8070 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1206_
timestamp 1700315010
transform -1 0 210 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1208_
timestamp 1700315010
transform -1 0 210 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1209_
timestamp 1700315010
transform 1 0 7170 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1211_
timestamp 1700315010
transform -1 0 6570 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1212_
timestamp 1700315010
transform 1 0 5550 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1214_
timestamp 1700315010
transform 1 0 6690 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1215_
timestamp 1700315010
transform -1 0 4230 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1217_
timestamp 1700315010
transform 1 0 6030 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1218_
timestamp 1700315010
transform -1 0 5490 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1219_
timestamp 1700315010
transform 1 0 3750 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1221_
timestamp 1700315010
transform -1 0 4650 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1222_
timestamp 1700315010
transform -1 0 5790 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1224_
timestamp 1700315010
transform -1 0 6390 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1225_
timestamp 1700315010
transform 1 0 5850 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1227_
timestamp 1700315010
transform 1 0 4770 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1228_
timestamp 1700315010
transform 1 0 5970 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1230_
timestamp 1700315010
transform 1 0 5610 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1231_
timestamp 1700315010
transform -1 0 5190 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1233_
timestamp 1700315010
transform 1 0 990 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1234_
timestamp 1700315010
transform 1 0 3390 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1236_
timestamp 1700315010
transform -1 0 930 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1237_
timestamp 1700315010
transform 1 0 1770 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1239_
timestamp 1700315010
transform -1 0 1590 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1240_
timestamp 1700315010
transform -1 0 1350 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1242_
timestamp 1700315010
transform 1 0 1950 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1243_
timestamp 1700315010
transform 1 0 1110 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1244_
timestamp 1700315010
transform 1 0 630 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1246_
timestamp 1700315010
transform -1 0 210 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1247_
timestamp 1700315010
transform -1 0 210 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1249_
timestamp 1700315010
transform 1 0 150 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1250_
timestamp 1700315010
transform -1 0 690 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1252_
timestamp 1700315010
transform 1 0 1470 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1253_
timestamp 1700315010
transform 1 0 150 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1255_
timestamp 1700315010
transform -1 0 210 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1256_
timestamp 1700315010
transform 1 0 1050 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1258_
timestamp 1700315010
transform 1 0 1110 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1259_
timestamp 1700315010
transform -1 0 2550 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1261_
timestamp 1700315010
transform 1 0 2910 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1262_
timestamp 1700315010
transform 1 0 630 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1264_
timestamp 1700315010
transform 1 0 1530 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1265_
timestamp 1700315010
transform -1 0 2070 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1266_
timestamp 1700315010
transform -1 0 2010 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1268_
timestamp 1700315010
transform 1 0 3270 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1269_
timestamp 1700315010
transform 1 0 3750 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1271_
timestamp 1700315010
transform -1 0 9330 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1272_
timestamp 1700315010
transform 1 0 15030 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1274_
timestamp 1700315010
transform 1 0 12510 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1275_
timestamp 1700315010
transform 1 0 11910 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1277_
timestamp 1700315010
transform 1 0 12390 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1278_
timestamp 1700315010
transform 1 0 14310 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1280_
timestamp 1700315010
transform -1 0 10710 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1281_
timestamp 1700315010
transform -1 0 11610 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1283_
timestamp 1700315010
transform -1 0 11130 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1284_
timestamp 1700315010
transform -1 0 5010 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1286_
timestamp 1700315010
transform -1 0 4590 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1287_
timestamp 1700315010
transform 1 0 5730 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1289_
timestamp 1700315010
transform 1 0 8550 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1290_
timestamp 1700315010
transform -1 0 9510 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1291_
timestamp 1700315010
transform -1 0 7230 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1293_
timestamp 1700315010
transform -1 0 7950 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1294_
timestamp 1700315010
transform 1 0 3810 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1296_
timestamp 1700315010
transform -1 0 5010 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1297_
timestamp 1700315010
transform 1 0 4890 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1299_
timestamp 1700315010
transform 1 0 2370 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1300_
timestamp 1700315010
transform -1 0 4890 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1302_
timestamp 1700315010
transform -1 0 5790 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1303_
timestamp 1700315010
transform -1 0 6270 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1305_
timestamp 1700315010
transform -1 0 4290 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1306_
timestamp 1700315010
transform 1 0 2370 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1308_
timestamp 1700315010
transform -1 0 210 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1309_
timestamp 1700315010
transform 1 0 3990 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1311_
timestamp 1700315010
transform 1 0 3330 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1312_
timestamp 1700315010
transform -1 0 5310 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1313_
timestamp 1700315010
transform -1 0 4110 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1315_
timestamp 1700315010
transform 1 0 3930 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1316_
timestamp 1700315010
transform -1 0 2370 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1318_
timestamp 1700315010
transform 1 0 8370 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1319_
timestamp 1700315010
transform -1 0 6210 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1321_
timestamp 1700315010
transform -1 0 4890 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1322_
timestamp 1700315010
transform -1 0 3510 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1324_
timestamp 1700315010
transform -1 0 2490 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1325_
timestamp 1700315010
transform -1 0 3090 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1327_
timestamp 1700315010
transform -1 0 210 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1328_
timestamp 1700315010
transform -1 0 210 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1330_
timestamp 1700315010
transform -1 0 1530 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1331_
timestamp 1700315010
transform 1 0 570 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1333_
timestamp 1700315010
transform 1 0 2430 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1334_
timestamp 1700315010
transform 1 0 1530 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1336_
timestamp 1700315010
transform 1 0 1470 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1337_
timestamp 1700315010
transform 1 0 3390 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1338_
timestamp 1700315010
transform 1 0 150 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1340_
timestamp 1700315010
transform 1 0 1950 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1341_
timestamp 1700315010
transform 1 0 510 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1343_
timestamp 1700315010
transform 1 0 990 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1344_
timestamp 1700315010
transform -1 0 2670 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1346_
timestamp 1700315010
transform 1 0 2730 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1347_
timestamp 1700315010
transform 1 0 3090 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1349_
timestamp 1700315010
transform -1 0 4230 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1350_
timestamp 1700315010
transform 1 0 1590 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1352_
timestamp 1700315010
transform 1 0 5250 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1353_
timestamp 1700315010
transform -1 0 3630 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1355_
timestamp 1700315010
transform -1 0 6510 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1356_
timestamp 1700315010
transform 1 0 9870 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1358_
timestamp 1700315010
transform 1 0 10770 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1359_
timestamp 1700315010
transform 1 0 13710 0 -1 5490
box -36 -24 96 816
use FILL  FILL_2__1360_
timestamp 1700315010
transform 1 0 13530 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1362_
timestamp 1700315010
transform 1 0 13050 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1363_
timestamp 1700315010
transform -1 0 12210 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1365_
timestamp 1700315010
transform -1 0 14490 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1366_
timestamp 1700315010
transform -1 0 4710 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1368_
timestamp 1700315010
transform 1 0 6330 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1369_
timestamp 1700315010
transform 1 0 8790 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1371_
timestamp 1700315010
transform 1 0 7530 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1372_
timestamp 1700315010
transform -1 0 3870 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1374_
timestamp 1700315010
transform -1 0 1590 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1375_
timestamp 1700315010
transform -1 0 1050 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1377_
timestamp 1700315010
transform -1 0 2670 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1378_
timestamp 1700315010
transform -1 0 3570 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1380_
timestamp 1700315010
transform -1 0 3510 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1381_
timestamp 1700315010
transform -1 0 3030 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1383_
timestamp 1700315010
transform -1 0 3030 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1384_
timestamp 1700315010
transform -1 0 3510 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1385_
timestamp 1700315010
transform -1 0 2550 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1387_
timestamp 1700315010
transform 1 0 1890 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1388_
timestamp 1700315010
transform 1 0 4770 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1390_
timestamp 1700315010
transform -1 0 5070 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1391_
timestamp 1700315010
transform -1 0 4530 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1393_
timestamp 1700315010
transform 1 0 5670 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1394_
timestamp 1700315010
transform 1 0 4170 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1396_
timestamp 1700315010
transform -1 0 1770 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1397_
timestamp 1700315010
transform -1 0 210 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1399_
timestamp 1700315010
transform -1 0 2070 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1400_
timestamp 1700315010
transform -1 0 930 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1402_
timestamp 1700315010
transform -1 0 510 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1403_
timestamp 1700315010
transform 1 0 1050 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1405_
timestamp 1700315010
transform 1 0 1050 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1406_
timestamp 1700315010
transform -1 0 210 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1407_
timestamp 1700315010
transform -1 0 210 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1409_
timestamp 1700315010
transform -1 0 690 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1410_
timestamp 1700315010
transform 1 0 630 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1412_
timestamp 1700315010
transform 1 0 1890 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1413_
timestamp 1700315010
transform -1 0 210 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1415_
timestamp 1700315010
transform -1 0 3930 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1416_
timestamp 1700315010
transform 1 0 5730 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1418_
timestamp 1700315010
transform -1 0 3690 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1419_
timestamp 1700315010
transform 1 0 4110 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1421_
timestamp 1700315010
transform -1 0 7410 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1422_
timestamp 1700315010
transform 1 0 8370 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1424_
timestamp 1700315010
transform 1 0 8610 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1425_
timestamp 1700315010
transform -1 0 9030 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1427_
timestamp 1700315010
transform 1 0 13830 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1428_
timestamp 1700315010
transform -1 0 12930 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1429_
timestamp 1700315010
transform 1 0 13050 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1431_
timestamp 1700315010
transform -1 0 14190 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1432_
timestamp 1700315010
transform 1 0 14250 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1434_
timestamp 1700315010
transform 1 0 13950 0 1 3930
box -36 -24 96 816
use FILL  FILL_2__1435_
timestamp 1700315010
transform 1 0 17850 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1437_
timestamp 1700315010
transform -1 0 11670 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1438_
timestamp 1700315010
transform 1 0 8010 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1440_
timestamp 1700315010
transform -1 0 3630 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1441_
timestamp 1700315010
transform 1 0 1530 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1443_
timestamp 1700315010
transform -1 0 6270 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1444_
timestamp 1700315010
transform -1 0 4290 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1446_
timestamp 1700315010
transform 1 0 4650 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1447_
timestamp 1700315010
transform 1 0 5070 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1449_
timestamp 1700315010
transform -1 0 5790 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1450_
timestamp 1700315010
transform -1 0 4710 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1452_
timestamp 1700315010
transform 1 0 5730 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1453_
timestamp 1700315010
transform 1 0 6270 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1454_
timestamp 1700315010
transform 1 0 5790 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1456_
timestamp 1700315010
transform -1 0 6510 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1457_
timestamp 1700315010
transform -1 0 5910 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1459_
timestamp 1700315010
transform -1 0 1470 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1460_
timestamp 1700315010
transform 1 0 5250 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1462_
timestamp 1700315010
transform -1 0 570 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1463_
timestamp 1700315010
transform -1 0 4350 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1465_
timestamp 1700315010
transform -1 0 3150 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1466_
timestamp 1700315010
transform -1 0 1830 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1468_
timestamp 1700315010
transform 1 0 4350 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1469_
timestamp 1700315010
transform -1 0 3390 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1471_
timestamp 1700315010
transform 1 0 2370 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1472_
timestamp 1700315010
transform 1 0 2850 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1474_
timestamp 1700315010
transform 1 0 8370 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1475_
timestamp 1700315010
transform 1 0 8250 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1476_
timestamp 1700315010
transform 1 0 8970 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1478_
timestamp 1700315010
transform 1 0 9750 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1479_
timestamp 1700315010
transform 1 0 10590 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1481_
timestamp 1700315010
transform -1 0 13110 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1482_
timestamp 1700315010
transform 1 0 13950 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1484_
timestamp 1700315010
transform -1 0 16590 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1485_
timestamp 1700315010
transform 1 0 16530 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1487_
timestamp 1700315010
transform 1 0 17490 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1488_
timestamp 1700315010
transform 1 0 6570 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1490_
timestamp 1700315010
transform -1 0 7110 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1491_
timestamp 1700315010
transform -1 0 8670 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1493_
timestamp 1700315010
transform -1 0 6810 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1494_
timestamp 1700315010
transform 1 0 7710 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1496_
timestamp 1700315010
transform 1 0 7230 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1497_
timestamp 1700315010
transform 1 0 7830 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1499_
timestamp 1700315010
transform 1 0 6690 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1500_
timestamp 1700315010
transform 1 0 7350 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1501_
timestamp 1700315010
transform 1 0 8190 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1503_
timestamp 1700315010
transform 1 0 8370 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1504_
timestamp 1700315010
transform 1 0 8610 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1506_
timestamp 1700315010
transform -1 0 7950 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1507_
timestamp 1700315010
transform -1 0 7470 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1509_
timestamp 1700315010
transform 1 0 6150 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1510_
timestamp 1700315010
transform -1 0 5790 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1512_
timestamp 1700315010
transform -1 0 8190 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1513_
timestamp 1700315010
transform 1 0 9990 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1515_
timestamp 1700315010
transform 1 0 9510 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1516_
timestamp 1700315010
transform -1 0 7650 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1518_
timestamp 1700315010
transform -1 0 9690 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1519_
timestamp 1700315010
transform 1 0 8790 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1521_
timestamp 1700315010
transform 1 0 7710 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1522_
timestamp 1700315010
transform 1 0 8190 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1523_
timestamp 1700315010
transform 1 0 8550 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1525_
timestamp 1700315010
transform -1 0 16470 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1526_
timestamp 1700315010
transform -1 0 14970 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1528_
timestamp 1700315010
transform 1 0 12990 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1529_
timestamp 1700315010
transform 1 0 13770 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1531_
timestamp 1700315010
transform -1 0 15270 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1532_
timestamp 1700315010
transform 1 0 15690 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1534_
timestamp 1700315010
transform -1 0 15510 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1535_
timestamp 1700315010
transform -1 0 11310 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1537_
timestamp 1700315010
transform 1 0 8430 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1538_
timestamp 1700315010
transform 1 0 7770 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1540_
timestamp 1700315010
transform -1 0 7950 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1541_
timestamp 1700315010
transform -1 0 8430 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1543_
timestamp 1700315010
transform 1 0 7950 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1544_
timestamp 1700315010
transform 1 0 7350 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1546_
timestamp 1700315010
transform -1 0 7530 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1547_
timestamp 1700315010
transform -1 0 8070 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1548_
timestamp 1700315010
transform -1 0 9150 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1550_
timestamp 1700315010
transform 1 0 10410 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1551_
timestamp 1700315010
transform 1 0 11730 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1553_
timestamp 1700315010
transform -1 0 15210 0 1 5490
box -36 -24 96 816
use FILL  FILL_2__1554_
timestamp 1700315010
transform 1 0 15690 0 -1 3930
box -36 -24 96 816
use FILL  FILL_2__1556_
timestamp 1700315010
transform -1 0 14970 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1557_
timestamp 1700315010
transform -1 0 14610 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1559_
timestamp 1700315010
transform 1 0 10590 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1560_
timestamp 1700315010
transform 1 0 10950 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1562_
timestamp 1700315010
transform 1 0 8070 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1563_
timestamp 1700315010
transform 1 0 11130 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1565_
timestamp 1700315010
transform -1 0 6510 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1566_
timestamp 1700315010
transform -1 0 6930 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1568_
timestamp 1700315010
transform 1 0 9990 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1569_
timestamp 1700315010
transform 1 0 11850 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1570_
timestamp 1700315010
transform 1 0 10110 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1572_
timestamp 1700315010
transform 1 0 10350 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1573_
timestamp 1700315010
transform 1 0 12330 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1575_
timestamp 1700315010
transform 1 0 12990 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1576_
timestamp 1700315010
transform 1 0 12510 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1578_
timestamp 1700315010
transform 1 0 17130 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1579_
timestamp 1700315010
transform -1 0 15390 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1581_
timestamp 1700315010
transform 1 0 14670 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1582_
timestamp 1700315010
transform -1 0 13530 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1584_
timestamp 1700315010
transform 1 0 8850 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1585_
timestamp 1700315010
transform 1 0 9330 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1587_
timestamp 1700315010
transform 1 0 7650 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1588_
timestamp 1700315010
transform -1 0 11610 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1590_
timestamp 1700315010
transform 1 0 14370 0 1 2370
box -36 -24 96 816
use FILL  FILL_2__1591_
timestamp 1700315010
transform -1 0 14250 0 -1 2370
box -36 -24 96 816
use FILL  FILL_2__1593_
timestamp 1700315010
transform -1 0 13050 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2__1594_
timestamp 1700315010
transform 1 0 12930 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1595_
timestamp 1700315010
transform 1 0 11970 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1597_
timestamp 1700315010
transform 1 0 12030 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1598_
timestamp 1700315010
transform -1 0 12510 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1600_
timestamp 1700315010
transform -1 0 12090 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1601_
timestamp 1700315010
transform 1 0 9930 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1603_
timestamp 1700315010
transform 1 0 8850 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1604_
timestamp 1700315010
transform -1 0 9330 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1606_
timestamp 1700315010
transform -1 0 15510 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1607_
timestamp 1700315010
transform 1 0 13290 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1636_
timestamp 1700315010
transform -1 0 17730 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1637_
timestamp 1700315010
transform 1 0 17730 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1639_
timestamp 1700315010
transform 1 0 15630 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1640_
timestamp 1700315010
transform 1 0 15630 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1642_
timestamp 1700315010
transform -1 0 9510 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1643_
timestamp 1700315010
transform -1 0 9030 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1644_
timestamp 1700315010
transform -1 0 11610 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1646_
timestamp 1700315010
transform -1 0 12330 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1647_
timestamp 1700315010
transform 1 0 9510 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1649_
timestamp 1700315010
transform -1 0 12870 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1650_
timestamp 1700315010
transform -1 0 13350 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1652_
timestamp 1700315010
transform -1 0 10890 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1653_
timestamp 1700315010
transform 1 0 12450 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1655_
timestamp 1700315010
transform -1 0 17010 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1656_
timestamp 1700315010
transform 1 0 17790 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1658_
timestamp 1700315010
transform 1 0 16890 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1659_
timestamp 1700315010
transform -1 0 16050 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1661_
timestamp 1700315010
transform 1 0 16050 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1662_
timestamp 1700315010
transform -1 0 10410 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1664_
timestamp 1700315010
transform -1 0 10350 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1665_
timestamp 1700315010
transform -1 0 10950 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1666_
timestamp 1700315010
transform -1 0 11490 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1668_
timestamp 1700315010
transform 1 0 11130 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1669_
timestamp 1700315010
transform -1 0 12150 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1671_
timestamp 1700315010
transform 1 0 15690 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1672_
timestamp 1700315010
transform -1 0 17010 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1674_
timestamp 1700315010
transform -1 0 16110 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1675_
timestamp 1700315010
transform -1 0 16650 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1677_
timestamp 1700315010
transform -1 0 14670 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1678_
timestamp 1700315010
transform -1 0 14790 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1680_
timestamp 1700315010
transform 1 0 13890 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1681_
timestamp 1700315010
transform -1 0 12030 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1683_
timestamp 1700315010
transform 1 0 14130 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1684_
timestamp 1700315010
transform 1 0 15090 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1686_
timestamp 1700315010
transform 1 0 12930 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1687_
timestamp 1700315010
transform -1 0 15330 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1689_
timestamp 1700315010
transform 1 0 14670 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1690_
timestamp 1700315010
transform 1 0 15270 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1691_
timestamp 1700315010
transform -1 0 14850 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1693_
timestamp 1700315010
transform 1 0 9330 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1694_
timestamp 1700315010
transform -1 0 9870 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1696_
timestamp 1700315010
transform -1 0 9150 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1697_
timestamp 1700315010
transform -1 0 9930 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1699_
timestamp 1700315010
transform -1 0 11670 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1700_
timestamp 1700315010
transform -1 0 11730 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1702_
timestamp 1700315010
transform 1 0 11190 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1703_
timestamp 1700315010
transform -1 0 13770 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1705_
timestamp 1700315010
transform 1 0 12150 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1706_
timestamp 1700315010
transform -1 0 13050 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1708_
timestamp 1700315010
transform 1 0 13470 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1709_
timestamp 1700315010
transform -1 0 11010 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1711_
timestamp 1700315010
transform -1 0 10710 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1712_
timestamp 1700315010
transform -1 0 11130 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1713_
timestamp 1700315010
transform -1 0 10230 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1715_
timestamp 1700315010
transform -1 0 11850 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1716_
timestamp 1700315010
transform 1 0 12270 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1718_
timestamp 1700315010
transform 1 0 13710 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1719_
timestamp 1700315010
transform 1 0 14190 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1721_
timestamp 1700315010
transform 1 0 14010 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2__1722_
timestamp 1700315010
transform 1 0 14310 0 1 17970
box -36 -24 96 816
use FILL  FILL_2__1724_
timestamp 1700315010
transform -1 0 14430 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1725_
timestamp 1700315010
transform 1 0 13290 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1727_
timestamp 1700315010
transform -1 0 13170 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1728_
timestamp 1700315010
transform -1 0 9090 0 1 16410
box -36 -24 96 816
use FILL  FILL_2__1730_
timestamp 1700315010
transform -1 0 9750 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1731_
timestamp 1700315010
transform -1 0 10170 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1733_
timestamp 1700315010
transform 1 0 11070 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1734_
timestamp 1700315010
transform 1 0 14910 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1736_
timestamp 1700315010
transform -1 0 15750 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1737_
timestamp 1700315010
transform 1 0 15210 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1738_
timestamp 1700315010
transform 1 0 15330 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1740_
timestamp 1700315010
transform -1 0 15510 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1741_
timestamp 1700315010
transform 1 0 15690 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1743_
timestamp 1700315010
transform -1 0 8370 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1744_
timestamp 1700315010
transform -1 0 8850 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1746_
timestamp 1700315010
transform 1 0 9210 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1747_
timestamp 1700315010
transform 1 0 10110 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1749_
timestamp 1700315010
transform 1 0 15690 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1750_
timestamp 1700315010
transform 1 0 16350 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1752_
timestamp 1700315010
transform -1 0 15870 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1753_
timestamp 1700315010
transform 1 0 16170 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1755_
timestamp 1700315010
transform 1 0 16170 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1756_
timestamp 1700315010
transform 1 0 14550 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1758_
timestamp 1700315010
transform 1 0 12750 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1759_
timestamp 1700315010
transform 1 0 12030 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1760_
timestamp 1700315010
transform 1 0 13590 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1762_
timestamp 1700315010
transform -1 0 15450 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1763_
timestamp 1700315010
transform 1 0 15870 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1765_
timestamp 1700315010
transform 1 0 17250 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1766_
timestamp 1700315010
transform 1 0 17550 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1768_
timestamp 1700315010
transform -1 0 14310 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1769_
timestamp 1700315010
transform -1 0 13830 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1771_
timestamp 1700315010
transform 1 0 16590 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1772_
timestamp 1700315010
transform 1 0 16650 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1774_
timestamp 1700315010
transform -1 0 16830 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1775_
timestamp 1700315010
transform -1 0 17190 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1777_
timestamp 1700315010
transform 1 0 14850 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1778_
timestamp 1700315010
transform 1 0 13470 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1780_
timestamp 1700315010
transform 1 0 12570 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1781_
timestamp 1700315010
transform 1 0 13950 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1783_
timestamp 1700315010
transform 1 0 16890 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1784_
timestamp 1700315010
transform 1 0 16470 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1785_
timestamp 1700315010
transform -1 0 17490 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1787_
timestamp 1700315010
transform -1 0 17730 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1788_
timestamp 1700315010
transform 1 0 17190 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1790_
timestamp 1700315010
transform 1 0 18030 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1791_
timestamp 1700315010
transform 1 0 17970 0 1 7050
box -36 -24 96 816
use FILL  FILL_2__1793_
timestamp 1700315010
transform 1 0 13590 0 1 11730
box -36 -24 96 816
use FILL  FILL_2__1794_
timestamp 1700315010
transform 1 0 14670 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1796_
timestamp 1700315010
transform 1 0 16290 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1797_
timestamp 1700315010
transform -1 0 15150 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1799_
timestamp 1700315010
transform -1 0 17670 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2__1800_
timestamp 1700315010
transform -1 0 17610 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1802_
timestamp 1700315010
transform 1 0 14310 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2__1803_
timestamp 1700315010
transform 1 0 17670 0 1 810
box -36 -24 96 816
use FILL  FILL_2__1805_
timestamp 1700315010
transform 1 0 18030 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1806_
timestamp 1700315010
transform -1 0 17130 0 1 13290
box -36 -24 96 816
use FILL  FILL_2__1807_
timestamp 1700315010
transform 1 0 17070 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1809_
timestamp 1700315010
transform 1 0 16950 0 1 14850
box -36 -24 96 816
use FILL  FILL_2__1810_
timestamp 1700315010
transform 1 0 17730 0 -1 14850
box -36 -24 96 816
use FILL  FILL_2__1812_
timestamp 1700315010
transform 1 0 17970 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2__1813_
timestamp 1700315010
transform -1 0 18030 0 1 10170
box -36 -24 96 816
use FILL  FILL_2__1815_
timestamp 1700315010
transform 1 0 17550 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2__1816_
timestamp 1700315010
transform -1 0 18030 0 1 8610
box -36 -24 96 816
use FILL  FILL_2__1818_
timestamp 1700315010
transform -1 0 9870 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1819_
timestamp 1700315010
transform -1 0 7830 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2__1821_
timestamp 1700315010
transform -1 0 16950 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1822_
timestamp 1700315010
transform 1 0 16470 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1824_
timestamp 1700315010
transform 1 0 14970 0 -1 810
box -36 -24 96 816
use FILL  FILL_2__1825_
timestamp 1700315010
transform 1 0 13830 0 -1 810
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert0
timestamp 1700315010
transform 1 0 11850 0 1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert1
timestamp 1700315010
transform -1 0 6690 0 1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert3
timestamp 1700315010
transform -1 0 6870 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert4
timestamp 1700315010
transform -1 0 13290 0 -1 11730
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert6
timestamp 1700315010
transform -1 0 8250 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert7
timestamp 1700315010
transform -1 0 10290 0 -1 7050
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert13
timestamp 1700315010
transform 1 0 15630 0 1 8610
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert14
timestamp 1700315010
transform -1 0 11550 0 1 10170
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert16
timestamp 1700315010
transform -1 0 12150 0 -1 8610
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert17
timestamp 1700315010
transform 1 0 7650 0 1 11730
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert19
timestamp 1700315010
transform 1 0 9150 0 1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert20
timestamp 1700315010
transform -1 0 7350 0 1 8610
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert22
timestamp 1700315010
transform -1 0 12690 0 1 10170
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert23
timestamp 1700315010
transform 1 0 12810 0 -1 10170
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert25
timestamp 1700315010
transform -1 0 7110 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert26
timestamp 1700315010
transform -1 0 8010 0 1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert28
timestamp 1700315010
transform 1 0 9570 0 1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert29
timestamp 1700315010
transform -1 0 6630 0 1 7050
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert31
timestamp 1700315010
transform -1 0 6690 0 -1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert32
timestamp 1700315010
transform 1 0 10590 0 1 13290
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert34
timestamp 1700315010
transform -1 0 18090 0 -1 16410
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert35
timestamp 1700315010
transform -1 0 14910 0 -1 17970
box -36 -24 96 816
use FILL  FILL_2_BUFX2_insert36
timestamp 1700315010
transform -1 0 17910 0 1 16410
box -36 -24 96 816
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 14910 0 1 8610
box -36 -24 96 816
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 17490 0 1 2370
box -36 -24 96 816
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 14970 0 -1 3930
box -36 -24 96 816
<< labels >>
flabel metal1 s 18429 6 18609 6 3 FreeSans 48 270 0 0 gnd
port 0 nsew
flabel metal1 s -189 6 -9 6 7 FreeSans 48 270 0 0 vdd
port 1 nsew
flabel metal2 s 10008 18888 10032 18912 3 FreeSans 48 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 14568 18888 14592 18912 3 FreeSans 48 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 14868 18888 14892 18912 3 FreeSans 48 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 15348 18888 15372 18912 3 FreeSans 48 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 17448 18888 17472 18912 3 FreeSans 48 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s 18528 16308 18552 16332 3 FreeSans 48 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal2 s 15108 -72 15132 -48 7 FreeSans 48 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 16188 -72 16212 -48 7 FreeSans 48 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 16608 -72 16632 -48 7 FreeSans 48 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 17028 -72 17052 -48 7 FreeSans 48 270 0 0 ACC_o[3]
port 14 nsew
flabel metal3 s -72 3528 -48 3552 7 FreeSans 48 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -72 6768 -48 6792 7 FreeSans 48 0 0 0 ACC_o[0]
port 17 nsew
flabel metal2 s 17388 -72 17412 -48 7 FreeSans 48 270 0 0 Done_o
port 18 nsew
flabel metal2 s 17568 18888 17592 18912 3 FreeSans 48 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s 18528 2748 18552 2772 3 FreeSans 48 0 0 0 clk
port 22 nsew
flabel metal3 s 18609 15828 18633 15852 3 FreeSans 48 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s 18609 15528 18633 15552 3 FreeSans 48 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal3 s 18609 4188 18633 4212 3 FreeSans 48 0 0 0 reset
port 23 nsew
flabel metal3 s -72 6588 -48 6612 7 FreeSans 48 0 0 0 ACC_o[1]
port 16 nsew
flabel metal2 s 13968 -72 13992 -48 7 FreeSans 48 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 18008 18888 18032 18912 3 FreeSans 48 90 0 0 LoadA_i
port 19 nsew
flabel metal2 s 17747 18888 17771 18912 3 FreeSans 48 90 0 0 LoadB_i
port 20 nsew
<< properties >>
string FIXED_BBOX -120 -120 18540 18900
<< end >>
