* NGSPICE file created from DFFSR.ext - technology: scmos

.subckt DFFSR D S R CLK Q vdd gnd
M1000 vdd S a_20_122# vdd pfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=5.4p ps=7.8u
M1001 vdd D a_114_12# vdd pfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=4.95p ps=7.8u
M1002 a_260_12# a_210_12# a_244_12# gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=10.8p ps=15.6u
M1003 a_20_122# a_46_54# vdd vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=5.4p ps=7.8u
M1004 a_226_12# S a_292_12# gnd nfet w=6u l=0.6u
+  ad=10.8p pd=15.6u as=3.6p ps=7.2u
M1005 a_226_12# a_244_12# vdd vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=5.4p ps=7.8u
M1006 a_20_12# R a_4_12# gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=10.8p ps=15.6u
M1007 vdd S a_226_12# vdd pfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=5.4p ps=7.8u
M1008 a_210_12# a_94_8# a_20_122# gnd nfet w=3u l=0.6u
+  ad=2.7p pd=4.8u as=4.5p ps=9u
M1009 gnd R a_260_12# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=3.6p ps=7.2u
M1010 gnd a_20_122# a_20_12# gnd nfet w=6u l=0.6u
+  ad=7.200001p pd=8.400001u as=3.6p ps=7.2u
M1011 a_20_122# S a_52_12# gnd nfet w=6u l=0.6u
+  ad=10.8p pd=15.6u as=3.6p ps=7.2u
M1012 gnd a_94_142# a_94_8# gnd nfet w=3u l=0.6u
+  ad=2.7p pd=4.8u as=4.5p ps=9u
M1013 vdd a_20_122# a_4_12# vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=5.4p ps=7.8u
M1014 a_94_142# CLK vdd vdd pfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=5.4p ps=7.8u
M1015 vdd R a_244_12# vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=5.4p ps=7.8u
M1016 a_226_12# a_94_8# a_210_12# vdd pfet w=3u l=0.6u
+  ad=4.5p pd=9u as=2.7p ps=4.8u
M1017 a_292_12# a_244_12# gnd gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=7.200001p ps=8.400001u
M1018 gnd a_244_12# Q gnd nfet w=3u l=0.6u
+  ad=4.5p pd=9u as=4.5p ps=9u
M1019 a_4_12# R vdd vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=9p ps=15.000001u
M1020 a_114_12# a_94_8# a_46_54# vdd pfet w=3u l=0.6u
+  ad=4.95p pd=7.8u as=2.7p ps=4.8u
M1021 vdd a_94_142# a_94_8# vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=9p ps=15.000001u
M1022 a_244_12# a_210_12# vdd vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=9p ps=15.000001u
M1023 a_210_12# a_94_142# a_20_122# vdd pfet w=3u l=0.6u
+  ad=2.7p pd=4.8u as=4.5p ps=9u
M1024 a_52_12# a_46_54# gnd gnd nfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=7.200001p ps=8.400001u
M1025 a_46_54# a_94_8# a_4_12# gnd nfet w=3u l=0.6u
+  ad=2.7p pd=4.8u as=4.5p ps=9u
M1026 a_226_12# a_94_142# a_210_12# gnd nfet w=3u l=0.6u
+  ad=4.5p pd=9u as=2.7p ps=4.8u
M1027 a_94_142# CLK gnd gnd nfet w=3u l=0.6u
+  ad=4.5p pd=9u as=2.7p ps=4.8u
M1028 vdd a_244_12# Q vdd pfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=9p ps=15.000001u
M1029 gnd D a_114_12# gnd nfet w=3u l=0.6u
+  ad=4.5p pd=9u as=2.7p ps=4.8u
M1030 a_114_12# a_94_142# a_46_54# gnd nfet w=3u l=0.6u
+  ad=2.7p pd=4.8u as=2.7p ps=4.8u
M1031 a_46_54# a_94_142# a_4_12# vdd pfet w=3u l=0.6u
+  ad=2.7p pd=4.8u as=4.5p ps=9u
.ends

