magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -60 -60 78 152
<< polysilicon >>
rect 1 85 17 91
rect 1 79 6 85
rect 12 79 17 85
rect 1 73 17 79
rect 1 67 6 73
rect 12 67 17 73
rect 1 61 17 67
rect 1 55 6 61
rect 12 55 17 61
rect 1 49 17 55
rect 1 43 6 49
rect 12 43 17 49
rect 1 37 17 43
rect 1 31 6 37
rect 12 31 17 37
rect 1 25 17 31
rect 1 19 6 25
rect 12 19 17 25
rect 1 13 17 19
rect 1 7 6 13
rect 12 7 17 13
rect 1 1 17 7
<< polycontact >>
rect 6 79 12 85
rect 6 67 12 73
rect 6 55 12 61
rect 6 43 12 49
rect 6 31 12 37
rect 6 19 12 25
rect 6 7 12 13
<< genericcontact >>
rect 6 79 12 85
rect 6 67 12 73
rect 6 55 12 61
rect 6 43 12 49
rect 6 31 12 37
rect 6 19 12 25
rect 6 7 12 13
<< metal1 >>
rect 0 85 18 92
rect 0 79 6 85
rect 12 79 18 85
rect 0 73 18 79
rect 0 67 6 73
rect 12 67 18 73
rect 0 61 18 67
rect 0 55 6 61
rect 12 55 18 61
rect 0 49 18 55
rect 0 43 6 49
rect 12 43 18 49
rect 0 37 18 43
rect 0 31 6 37
rect 12 31 18 37
rect 0 25 18 31
rect 0 19 6 25
rect 12 19 18 25
rect 0 13 18 19
rect 0 7 6 13
rect 12 7 18 13
rect 0 0 18 7
<< end >>
