magic
tech scmos
timestamp 1700409309
<< metal1 >>
rect 590 242 618 243
rect 583 241 621 242
rect 548 240 550 241
rect 578 240 623 241
rect 545 239 555 240
rect 574 239 624 240
rect 544 238 559 239
rect 569 238 626 239
rect 543 237 628 238
rect 542 236 629 237
rect 541 235 630 236
rect 541 234 632 235
rect 541 233 633 234
rect 541 232 555 233
rect 557 232 586 233
rect 599 232 634 233
rect 541 231 550 232
rect 563 231 586 232
rect 603 231 635 232
rect 542 230 549 231
rect 565 230 589 231
rect 607 230 636 231
rect 531 229 533 230
rect 543 229 546 230
rect 566 229 593 230
rect 613 229 637 230
rect 528 228 536 229
rect 567 228 596 229
rect 621 228 638 229
rect 527 227 538 228
rect 551 227 555 228
rect 568 227 599 228
rect 625 227 639 228
rect 526 226 539 227
rect 548 226 558 227
rect 568 226 602 227
rect 629 226 640 227
rect 525 225 540 226
rect 546 225 559 226
rect 568 225 607 226
rect 632 225 641 226
rect 524 224 541 225
rect 544 224 560 225
rect 568 224 618 225
rect 635 224 641 225
rect 523 222 561 224
rect 568 223 622 224
rect 638 223 642 224
rect 568 222 625 223
rect 640 222 642 223
rect 522 221 561 222
rect 521 220 561 221
rect 567 221 628 222
rect 567 220 631 221
rect 520 219 560 220
rect 566 219 633 220
rect 519 218 560 219
rect 567 218 636 219
rect 518 217 559 218
rect 569 217 639 218
rect 517 216 558 217
rect 570 216 597 217
rect 598 216 641 217
rect 516 215 557 216
rect 572 215 597 216
rect 601 215 643 216
rect 515 214 535 215
rect 537 214 556 215
rect 573 214 597 215
rect 604 214 645 215
rect 513 213 530 214
rect 536 213 555 214
rect 574 213 597 214
rect 606 213 647 214
rect 512 212 527 213
rect 534 212 554 213
rect 576 212 598 213
rect 609 212 647 213
rect 510 211 524 212
rect 533 211 553 212
rect 577 211 598 212
rect 611 211 648 212
rect 508 210 523 211
rect 531 210 552 211
rect 578 210 599 211
rect 614 210 649 211
rect 506 209 521 210
rect 529 209 552 210
rect 504 208 519 209
rect 502 207 518 208
rect 522 207 523 208
rect 528 207 552 209
rect 560 209 561 210
rect 565 209 566 210
rect 579 209 600 210
rect 619 209 649 210
rect 560 208 570 209
rect 580 208 601 209
rect 623 208 650 209
rect 500 206 523 207
rect 527 206 552 207
rect 499 205 523 206
rect 497 204 523 205
rect 526 205 552 206
rect 561 207 572 208
rect 581 207 602 208
rect 625 207 650 208
rect 561 205 573 207
rect 581 206 604 207
rect 627 206 650 207
rect 582 205 606 206
rect 629 205 651 206
rect 526 204 553 205
rect 496 203 524 204
rect 525 203 553 204
rect 495 201 553 203
rect 494 200 553 201
rect 562 204 574 205
rect 583 204 609 205
rect 631 204 651 205
rect 562 202 575 204
rect 584 203 612 204
rect 633 203 651 204
rect 584 202 616 203
rect 634 202 651 203
rect 562 200 576 202
rect 585 201 621 202
rect 636 201 652 202
rect 585 200 623 201
rect 637 200 652 201
rect 494 199 554 200
rect 494 198 503 199
rect 504 198 554 199
rect 495 197 501 198
rect 503 197 554 198
rect 496 196 498 197
rect 502 196 554 197
rect 501 195 554 196
rect 562 198 577 200
rect 586 199 625 200
rect 638 199 652 200
rect 586 198 627 199
rect 639 198 652 199
rect 562 196 578 198
rect 587 197 628 198
rect 641 197 652 198
rect 587 196 630 197
rect 642 196 652 197
rect 500 194 553 195
rect 499 192 553 194
rect 562 194 579 196
rect 588 195 631 196
rect 643 195 652 196
rect 588 194 632 195
rect 644 194 652 195
rect 562 192 580 194
rect 589 193 634 194
rect 590 192 635 193
rect 645 192 652 194
rect 498 190 552 192
rect 561 191 581 192
rect 592 191 636 192
rect 646 191 652 192
rect 498 189 551 190
rect 561 189 582 191
rect 594 190 637 191
rect 647 190 652 191
rect 597 189 638 190
rect 499 188 551 189
rect 560 188 583 189
rect 602 188 639 189
rect 648 188 652 190
rect 499 187 550 188
rect 560 187 585 188
rect 608 187 640 188
rect 500 186 549 187
rect 560 186 586 187
rect 611 186 641 187
rect 649 186 651 188
rect 500 185 521 186
rect 524 185 549 186
rect 559 185 589 186
rect 614 185 642 186
rect 501 184 520 185
rect 525 184 548 185
rect 559 184 592 185
rect 616 184 642 185
rect 502 183 519 184
rect 526 183 547 184
rect 503 182 516 183
rect 525 182 547 183
rect 558 183 597 184
rect 619 183 643 184
rect 558 182 602 183
rect 621 182 643 183
rect 524 181 546 182
rect 557 181 605 182
rect 623 181 643 182
rect 521 180 545 181
rect 557 180 608 181
rect 624 180 643 181
rect 516 179 545 180
rect 556 179 610 180
rect 625 179 644 180
rect 507 178 544 179
rect 556 178 612 179
rect 626 178 644 179
rect 506 177 543 178
rect 555 177 614 178
rect 627 177 644 178
rect 505 176 543 177
rect 554 176 616 177
rect 628 176 644 177
rect 505 175 542 176
rect 553 175 617 176
rect 629 175 644 176
rect 505 174 541 175
rect 553 174 618 175
rect 506 173 540 174
rect 552 173 619 174
rect 630 173 644 175
rect 506 172 539 173
rect 551 172 620 173
rect 0 154 111 172
rect 131 171 244 172
rect 261 171 369 172
rect 130 154 245 171
rect 261 170 371 171
rect 261 169 373 170
rect 261 168 375 169
rect 261 167 376 168
rect 261 165 377 167
rect 261 164 378 165
rect 261 162 379 164
rect 261 157 380 162
rect 261 154 381 157
rect 0 153 35 154
rect 0 139 34 153
rect 0 138 110 139
rect 0 120 111 138
rect 0 119 35 120
rect 0 105 34 119
rect 0 98 111 105
rect 1 96 111 98
rect 2 94 111 96
rect 3 93 111 94
rect 4 91 111 93
rect 5 90 111 91
rect 7 89 111 90
rect 8 88 111 89
rect 11 87 111 88
rect 170 87 205 154
rect 261 87 296 154
rect 346 127 381 154
rect 307 126 308 127
rect 309 126 344 127
rect 345 126 380 127
rect 307 125 348 126
rect 308 124 349 125
rect 309 123 350 124
rect 310 122 351 123
rect 311 121 352 122
rect 312 120 353 121
rect 313 119 354 120
rect 314 118 355 119
rect 315 117 356 118
rect 316 116 357 117
rect 317 115 358 116
rect 318 114 359 115
rect 319 113 360 114
rect 320 112 361 113
rect 321 111 362 112
rect 322 110 363 111
rect 323 109 364 110
rect 324 108 365 109
rect 325 107 366 108
rect 326 106 367 107
rect 327 105 368 106
rect 328 104 369 105
rect 329 103 370 104
rect 330 102 371 103
rect 331 101 372 102
rect 332 100 373 101
rect 333 99 374 100
rect 334 98 375 99
rect 335 97 376 98
rect 336 96 377 97
rect 337 95 378 96
rect 338 94 379 95
rect 339 93 380 94
rect 340 92 381 93
rect 341 91 382 92
rect 342 90 383 91
rect 343 89 384 90
rect 344 88 385 89
rect 345 87 386 88
rect 406 87 440 172
rect 507 171 537 172
rect 550 171 580 172
rect 585 171 620 172
rect 631 171 644 173
rect 507 170 535 171
rect 549 170 579 171
rect 588 170 621 171
rect 508 169 533 170
rect 548 169 578 170
rect 590 169 622 170
rect 632 169 644 171
rect 509 168 531 169
rect 547 168 577 169
rect 591 168 622 169
rect 509 167 528 168
rect 545 167 577 168
rect 592 167 623 168
rect 633 167 643 169
rect 510 166 526 167
rect 544 166 576 167
rect 593 166 623 167
rect 510 165 522 166
rect 542 165 576 166
rect 594 165 623 166
rect 634 165 643 167
rect 510 164 519 165
rect 540 164 576 165
rect 595 164 623 165
rect 511 163 516 164
rect 538 163 575 164
rect 596 163 623 164
rect 635 164 643 165
rect 536 162 575 163
rect 584 162 585 163
rect 597 162 624 163
rect 635 162 642 164
rect 534 161 575 162
rect 583 161 586 162
rect 597 161 623 162
rect 531 160 574 161
rect 583 160 587 161
rect 529 159 574 160
rect 582 159 587 160
rect 598 159 623 161
rect 636 161 642 162
rect 636 159 641 161
rect 527 158 573 159
rect 582 158 588 159
rect 525 157 573 158
rect 523 156 572 157
rect 581 156 589 158
rect 599 157 623 159
rect 637 157 640 159
rect 521 155 572 156
rect 520 154 571 155
rect 580 154 590 156
rect 599 155 622 157
rect 637 156 639 157
rect 637 155 638 156
rect 600 154 621 155
rect 519 153 570 154
rect 518 152 570 153
rect 517 151 569 152
rect 579 151 591 154
rect 600 153 620 154
rect 600 151 619 153
rect 516 150 568 151
rect 515 149 567 150
rect 578 149 592 151
rect 515 148 566 149
rect 577 148 592 149
rect 514 147 565 148
rect 514 146 564 147
rect 576 146 592 148
rect 601 150 618 151
rect 601 149 617 150
rect 601 148 616 149
rect 629 148 630 149
rect 601 147 614 148
rect 628 147 631 148
rect 601 146 613 147
rect 627 146 631 147
rect 513 145 563 146
rect 575 145 593 146
rect 513 144 562 145
rect 512 143 561 144
rect 574 143 593 145
rect 512 142 560 143
rect 573 142 593 143
rect 512 141 558 142
rect 572 141 593 142
rect 601 145 611 146
rect 626 145 631 146
rect 601 144 610 145
rect 625 144 631 145
rect 601 143 608 144
rect 624 143 631 144
rect 601 142 606 143
rect 623 142 631 143
rect 601 141 604 142
rect 622 141 631 142
rect 512 140 557 141
rect 571 140 593 141
rect 620 140 631 141
rect 511 139 555 140
rect 570 139 593 140
rect 619 139 631 140
rect 511 138 553 139
rect 568 138 593 139
rect 617 138 631 139
rect 511 137 552 138
rect 567 137 593 138
rect 616 137 631 138
rect 511 136 549 137
rect 566 136 592 137
rect 614 136 631 137
rect 511 135 547 136
rect 564 135 592 136
rect 612 135 631 136
rect 511 134 545 135
rect 562 134 592 135
rect 611 134 631 135
rect 511 133 543 134
rect 561 133 592 134
rect 609 133 631 134
rect 511 132 540 133
rect 559 132 592 133
rect 606 132 631 133
rect 511 131 538 132
rect 557 131 591 132
rect 604 131 631 132
rect 512 130 537 131
rect 555 130 591 131
rect 601 130 630 131
rect 512 129 535 130
rect 553 129 591 130
rect 598 129 630 130
rect 512 128 534 129
rect 551 128 591 129
rect 594 128 630 129
rect 512 127 533 128
rect 549 127 630 128
rect 512 126 532 127
rect 548 126 629 127
rect 513 125 531 126
rect 546 125 629 126
rect 513 123 530 125
rect 545 124 629 125
rect 543 123 628 124
rect 514 121 529 123
rect 542 122 628 123
rect 541 121 628 122
rect 515 119 528 121
rect 540 120 627 121
rect 539 119 571 120
rect 573 119 627 120
rect 516 117 528 119
rect 538 118 569 119
rect 573 118 626 119
rect 537 117 568 118
rect 572 117 626 118
rect 517 115 527 117
rect 536 116 566 117
rect 572 116 625 117
rect 536 115 565 116
rect 518 114 527 115
rect 519 112 527 114
rect 535 114 563 115
rect 571 114 624 116
rect 535 113 562 114
rect 570 113 623 114
rect 520 111 527 112
rect 534 112 560 113
rect 569 112 622 113
rect 534 111 559 112
rect 568 111 622 112
rect 521 110 526 111
rect 522 109 526 110
rect 523 108 526 109
rect 533 110 558 111
rect 568 110 591 111
rect 593 110 621 111
rect 533 109 557 110
rect 567 109 590 110
rect 592 109 620 110
rect 533 108 556 109
rect 566 108 589 109
rect 592 108 619 109
rect 524 107 526 108
rect 525 106 526 107
rect 532 107 555 108
rect 565 107 587 108
rect 532 106 554 107
rect 565 106 586 107
rect 591 106 618 108
rect 532 104 553 106
rect 564 105 585 106
rect 591 105 617 106
rect 564 104 584 105
rect 591 104 616 105
rect 531 103 552 104
rect 563 103 584 104
rect 590 103 615 104
rect 531 101 551 103
rect 563 102 583 103
rect 590 102 614 103
rect 531 99 550 101
rect 562 100 582 102
rect 590 101 612 102
rect 590 100 611 101
rect 532 98 550 99
rect 561 99 581 100
rect 590 99 610 100
rect 532 96 549 98
rect 561 96 580 99
rect 590 98 609 99
rect 589 97 608 98
rect 589 96 606 97
rect 533 94 549 96
rect 534 93 549 94
rect 535 92 549 93
rect 536 90 549 92
rect 537 89 549 90
rect 539 88 549 89
rect 540 87 549 88
rect 15 86 110 87
rect 171 86 204 87
rect 346 86 387 87
rect 407 86 440 87
rect 541 86 549 87
rect 347 85 388 86
rect 543 85 549 86
rect 348 84 389 85
rect 544 84 549 85
rect 560 93 579 96
rect 589 95 605 96
rect 589 94 604 95
rect 589 93 602 94
rect 560 88 578 93
rect 589 92 601 93
rect 589 91 600 92
rect 589 90 599 91
rect 590 89 598 90
rect 590 88 597 89
rect 349 83 390 84
rect 545 83 550 84
rect 560 83 577 88
rect 590 86 596 88
rect 590 85 595 86
rect 590 84 594 85
rect 350 82 391 83
rect 546 82 550 83
rect 351 81 392 82
rect 548 81 550 82
rect 549 80 550 81
rect 561 80 577 83
rect 591 83 594 84
rect 591 81 593 83
rect 591 80 592 81
rect 562 79 577 80
rect 562 78 578 79
rect 563 76 578 78
rect 564 75 578 76
rect 565 74 578 75
rect 566 73 578 74
rect 567 72 579 73
rect 568 71 579 72
rect 569 70 579 71
rect 570 69 580 70
rect 571 68 580 69
rect 572 67 580 68
rect 574 66 581 67
rect 8 65 20 66
rect 29 65 33 66
rect 132 65 136 66
rect 8 62 21 65
rect 8 61 20 62
rect 3 55 26 60
rect 29 54 34 65
rect 56 59 84 64
rect 78 56 84 59
rect 106 58 125 63
rect 112 57 118 58
rect 131 57 136 65
rect 180 65 184 66
rect 155 61 175 62
rect 155 57 176 61
rect 113 56 118 57
rect 125 56 136 57
rect 162 56 168 57
rect 35 54 37 55
rect 11 53 18 54
rect 8 52 21 53
rect 6 51 22 52
rect 5 50 23 51
rect 5 49 24 50
rect 4 48 11 49
rect 18 48 24 49
rect 4 45 10 48
rect 19 46 24 48
rect 29 49 38 54
rect 78 53 83 56
rect 112 55 118 56
rect 112 53 119 55
rect 77 50 83 53
rect 111 52 120 53
rect 124 52 136 56
rect 163 54 168 56
rect 111 51 121 52
rect 110 50 122 51
rect 19 45 25 46
rect 4 44 11 45
rect 17 44 24 45
rect 5 43 24 44
rect 6 42 23 43
rect 7 41 22 42
rect 9 40 20 41
rect 8 37 13 38
rect 29 37 34 49
rect 52 46 88 50
rect 109 49 123 50
rect 108 48 115 49
rect 116 48 124 49
rect 106 47 115 48
rect 117 47 126 48
rect 105 46 114 47
rect 118 46 126 47
rect 53 45 88 46
rect 103 45 113 46
rect 119 45 126 46
rect 67 39 72 45
rect 104 44 112 45
rect 120 44 125 45
rect 105 43 110 44
rect 122 43 124 44
rect 106 42 109 43
rect 8 32 14 37
rect 29 36 33 37
rect 56 34 84 39
rect 8 31 34 32
rect 8 27 35 31
rect 79 26 84 34
rect 110 32 115 40
rect 131 37 136 52
rect 162 51 168 54
rect 180 51 185 65
rect 208 61 235 65
rect 264 64 268 65
rect 264 61 269 64
rect 208 60 214 61
rect 232 60 233 61
rect 208 59 213 60
rect 208 58 234 59
rect 208 55 235 58
rect 263 56 269 61
rect 208 54 214 55
rect 263 54 270 56
rect 208 53 213 54
rect 262 53 270 54
rect 208 52 214 53
rect 261 52 271 53
rect 162 48 169 51
rect 161 47 169 48
rect 180 50 186 51
rect 188 50 189 51
rect 161 46 170 47
rect 160 45 170 46
rect 180 45 190 50
rect 208 48 235 52
rect 261 51 272 52
rect 260 50 273 51
rect 259 49 266 50
rect 267 49 274 50
rect 258 48 265 49
rect 267 48 275 49
rect 218 46 224 48
rect 257 47 264 48
rect 268 47 277 48
rect 255 46 264 47
rect 269 46 278 47
rect 204 45 238 46
rect 254 45 263 46
rect 270 45 278 46
rect 160 44 171 45
rect 159 43 171 44
rect 159 42 165 43
rect 158 41 165 42
rect 166 42 172 43
rect 166 41 173 42
rect 157 40 164 41
rect 167 40 174 41
rect 156 39 163 40
rect 155 38 163 39
rect 168 39 175 40
rect 168 38 176 39
rect 154 37 162 38
rect 169 37 177 38
rect 153 36 161 37
rect 170 36 176 37
rect 153 35 160 36
rect 171 35 176 36
rect 154 34 159 35
rect 173 34 175 35
rect 155 33 158 34
rect 110 27 137 32
rect 180 26 185 45
rect 203 41 239 45
rect 254 44 262 45
rect 272 44 277 45
rect 255 43 260 44
rect 273 43 276 44
rect 256 42 259 43
rect 257 41 258 42
rect 261 39 265 40
rect 213 38 229 39
rect 210 37 232 38
rect 209 36 233 37
rect 208 35 235 36
rect 207 34 216 35
rect 226 34 235 35
rect 207 31 213 34
rect 229 33 236 34
rect 230 32 236 33
rect 229 31 236 32
rect 261 32 266 39
rect 282 37 287 66
rect 316 64 317 65
rect 311 63 320 64
rect 310 62 322 63
rect 309 61 323 62
rect 332 61 337 66
rect 413 65 424 66
rect 412 64 425 65
rect 308 60 337 61
rect 307 59 315 60
rect 316 59 337 60
rect 358 59 386 64
rect 411 63 426 64
rect 410 62 427 63
rect 307 58 313 59
rect 319 58 337 59
rect 306 57 312 58
rect 306 52 311 57
rect 320 56 337 58
rect 320 55 326 56
rect 321 53 326 55
rect 332 53 337 56
rect 306 50 312 52
rect 320 51 337 53
rect 380 55 386 59
rect 409 61 416 62
rect 421 61 428 62
rect 409 60 415 61
rect 422 60 428 61
rect 409 57 414 60
rect 423 57 428 60
rect 409 56 416 57
rect 421 56 428 57
rect 409 55 427 56
rect 380 51 385 55
rect 410 54 427 55
rect 411 53 426 54
rect 413 52 424 53
rect 416 51 422 52
rect 319 50 337 51
rect 307 49 313 50
rect 318 49 337 50
rect 307 48 337 49
rect 308 47 324 48
rect 309 46 323 47
rect 310 45 321 46
rect 312 44 319 45
rect 311 32 316 40
rect 332 37 337 48
rect 379 50 385 51
rect 430 50 432 51
rect 379 47 384 50
rect 354 43 390 47
rect 406 46 432 50
rect 406 45 430 46
rect 355 42 390 43
rect 414 44 420 45
rect 261 31 287 32
rect 207 30 215 31
rect 227 30 235 31
rect 208 29 235 30
rect 209 28 234 29
rect 210 27 233 28
rect 261 27 288 31
rect 311 27 338 32
rect 212 26 230 27
rect 369 26 374 42
rect 414 38 419 44
rect 426 43 427 44
rect 428 43 432 44
rect 433 43 438 66
rect 576 65 581 66
rect 577 64 581 65
rect 579 63 582 64
rect 471 45 481 47
rect 484 45 493 47
rect 496 45 506 47
rect 510 45 518 47
rect 521 45 531 47
rect 536 45 545 47
rect 547 45 554 47
rect 563 45 571 47
rect 582 46 593 47
rect 579 45 585 46
rect 588 45 594 46
rect 607 45 617 47
rect 621 45 631 47
rect 636 45 652 47
rect 657 45 674 47
rect 473 44 479 45
rect 486 44 490 45
rect 498 44 504 45
rect 425 39 438 43
rect 412 32 417 37
rect 433 36 438 39
rect 474 36 478 44
rect 486 43 488 44
rect 499 43 504 44
rect 512 44 515 45
rect 523 44 529 45
rect 538 44 543 45
rect 550 44 555 45
rect 512 43 514 44
rect 485 42 487 43
rect 484 41 486 42
rect 500 41 505 43
rect 511 42 514 43
rect 511 41 513 42
rect 483 40 485 41
rect 482 39 484 40
rect 501 39 506 41
rect 510 39 512 41
rect 481 38 483 39
rect 502 38 507 39
rect 480 37 483 38
rect 503 37 507 38
rect 509 37 511 39
rect 479 36 484 37
rect 503 36 510 37
rect 474 35 485 36
rect 412 27 439 32
rect 474 27 478 35
rect 479 34 485 35
rect 504 35 510 36
rect 480 33 486 34
rect 481 32 487 33
rect 482 31 487 32
rect 482 30 488 31
rect 483 29 489 30
rect 484 28 490 29
rect 484 27 491 28
rect 473 26 479 27
rect 485 26 492 27
rect 504 26 509 35
rect 523 32 528 44
rect 524 31 528 32
rect 524 28 529 31
rect 539 30 542 44
rect 550 43 556 44
rect 550 42 557 43
rect 550 41 558 42
rect 566 41 569 45
rect 578 44 583 45
rect 590 44 594 45
rect 609 44 615 45
rect 623 44 629 45
rect 577 43 581 44
rect 591 43 594 44
rect 576 42 581 43
rect 592 42 594 43
rect 575 41 580 42
rect 538 28 541 30
rect 525 27 530 28
rect 537 27 541 28
rect 550 28 552 41
rect 553 40 559 41
rect 553 39 560 40
rect 554 38 561 39
rect 555 37 561 38
rect 556 36 562 37
rect 557 35 563 36
rect 558 34 564 35
rect 559 33 565 34
rect 559 32 566 33
rect 567 32 568 41
rect 574 38 579 41
rect 593 40 594 42
rect 610 43 615 44
rect 573 33 579 38
rect 610 37 614 43
rect 624 37 629 44
rect 610 35 629 37
rect 586 34 596 35
rect 587 33 595 34
rect 560 31 568 32
rect 561 30 568 31
rect 574 31 579 33
rect 589 32 594 33
rect 574 30 580 31
rect 562 29 568 30
rect 563 28 568 29
rect 575 29 580 30
rect 575 28 581 29
rect 525 26 532 27
rect 536 26 540 27
rect 550 26 553 28
rect 564 26 568 28
rect 576 27 581 28
rect 590 27 594 32
rect 610 27 614 35
rect 577 26 583 27
rect 217 25 226 26
rect 471 24 481 26
rect 486 24 494 26
rect 502 25 512 26
rect 526 25 539 26
rect 548 25 555 26
rect 565 25 568 26
rect 579 25 585 26
rect 589 25 594 27
rect 609 26 615 27
rect 624 26 629 35
rect 638 37 643 45
rect 649 44 652 45
rect 650 43 652 44
rect 651 41 652 43
rect 649 37 650 39
rect 638 35 650 37
rect 638 26 643 35
rect 648 34 650 35
rect 649 32 650 34
rect 660 37 665 45
rect 671 44 674 45
rect 672 41 674 44
rect 671 38 672 39
rect 670 37 672 38
rect 660 35 672 37
rect 652 28 654 30
rect 651 27 654 28
rect 650 26 653 27
rect 660 26 665 35
rect 670 33 672 35
rect 671 32 672 33
rect 674 29 676 30
rect 673 27 675 29
rect 672 26 675 27
rect 501 24 513 25
rect 528 24 538 25
rect 547 24 556 25
rect 566 24 568 25
rect 581 24 593 25
rect 607 24 617 26
rect 621 24 631 26
rect 635 24 653 26
rect 657 25 675 26
rect 657 24 674 25
rect 14 18 16 19
rect 121 18 122 19
rect 148 18 149 19
rect 359 18 360 19
rect 4 15 12 17
rect 4 11 7 15
rect 4 8 11 11
rect 4 5 7 8
rect 4 4 11 5
rect 4 2 12 4
rect 13 2 16 18
rect 21 13 23 14
rect 30 13 33 14
rect 36 13 39 16
rect 69 15 72 18
rect 46 13 47 14
rect 51 13 54 14
rect 63 13 65 14
rect 77 13 79 14
rect 84 13 86 14
rect 96 13 99 14
rect 108 13 110 14
rect 117 13 118 14
rect 120 13 123 18
rect 128 15 138 17
rect 131 14 135 15
rect 19 12 25 13
rect 29 12 41 13
rect 18 11 25 12
rect 28 11 41 12
rect 42 11 48 13
rect 50 12 56 13
rect 49 11 56 12
rect 59 11 67 13
rect 18 10 21 11
rect 18 9 20 10
rect 23 9 26 11
rect 18 6 26 9
rect 27 10 31 11
rect 18 5 20 6
rect 27 5 30 10
rect 18 4 21 5
rect 24 4 25 5
rect 28 4 31 5
rect 33 4 34 5
rect 18 3 26 4
rect 28 3 34 4
rect 36 4 39 11
rect 42 10 52 11
rect 36 3 41 4
rect 19 2 25 3
rect 29 2 34 3
rect 37 2 41 3
rect 42 2 45 10
rect 48 5 51 10
rect 54 9 57 11
rect 55 7 57 9
rect 54 5 57 7
rect 48 4 52 5
rect 53 4 57 5
rect 49 3 56 4
rect 50 2 55 3
rect 59 2 62 11
rect 64 10 67 11
rect 65 2 67 10
rect 69 2 72 13
rect 75 12 80 13
rect 82 12 88 13
rect 95 12 101 13
rect 104 12 111 13
rect 115 12 123 13
rect 74 11 80 12
rect 81 11 88 12
rect 94 11 102 12
rect 74 8 77 11
rect 81 9 84 11
rect 94 10 96 11
rect 99 9 102 11
rect 81 8 86 9
rect 95 8 102 9
rect 74 7 76 8
rect 82 7 87 8
rect 94 7 102 8
rect 74 5 77 7
rect 84 6 88 7
rect 94 6 97 7
rect 74 4 78 5
rect 79 4 80 5
rect 82 4 83 5
rect 85 4 88 6
rect 93 5 96 6
rect 99 5 102 7
rect 74 3 88 4
rect 94 4 97 5
rect 98 4 102 5
rect 94 3 102 4
rect 75 2 87 3
rect 95 2 102 3
rect 104 11 112 12
rect 104 9 107 11
rect 104 2 106 9
rect 109 2 112 11
rect 114 11 123 12
rect 114 8 117 11
rect 119 9 123 11
rect 114 7 116 8
rect 114 5 117 7
rect 120 6 123 9
rect 114 4 118 5
rect 119 4 123 6
rect 114 3 123 4
rect 115 2 123 3
rect 132 2 135 14
rect 140 13 142 14
rect 138 12 144 13
rect 137 11 144 12
rect 137 10 140 11
rect 137 9 139 10
rect 142 9 145 11
rect 136 6 145 9
rect 137 5 139 6
rect 137 4 140 5
rect 143 4 145 5
rect 137 3 145 4
rect 138 2 144 3
rect 147 2 149 18
rect 231 15 233 18
rect 254 15 256 16
rect 259 15 262 18
rect 297 16 305 17
rect 297 15 306 16
rect 154 13 156 14
rect 164 13 166 14
rect 172 13 174 14
rect 183 13 185 14
rect 188 13 190 14
rect 198 13 200 14
rect 204 13 206 14
rect 224 13 227 14
rect 238 13 241 14
rect 245 13 248 14
rect 253 13 256 15
rect 297 14 301 15
rect 302 14 306 15
rect 267 13 270 14
rect 279 13 281 14
rect 287 13 290 14
rect 152 12 158 13
rect 162 12 167 13
rect 170 12 176 13
rect 179 12 186 13
rect 187 12 192 13
rect 152 11 159 12
rect 151 9 154 11
rect 156 10 159 11
rect 161 11 167 12
rect 169 11 177 12
rect 161 10 164 11
rect 168 10 172 11
rect 157 9 159 10
rect 151 6 159 9
rect 160 6 163 10
rect 151 5 154 6
rect 160 5 164 6
rect 168 5 171 10
rect 174 9 177 11
rect 179 11 192 12
rect 175 6 178 9
rect 151 4 155 5
rect 157 4 159 5
rect 152 3 159 4
rect 161 4 165 5
rect 166 4 167 5
rect 168 4 172 5
rect 174 4 177 6
rect 161 3 167 4
rect 169 3 177 4
rect 153 2 159 3
rect 162 2 167 3
rect 170 2 176 3
rect 179 2 182 11
rect 184 10 188 11
rect 189 10 192 11
rect 184 2 187 10
rect 190 2 192 10
rect 194 11 207 13
rect 194 10 198 11
rect 194 2 197 10
rect 199 9 203 11
rect 200 2 202 9
rect 205 2 208 11
rect 210 5 212 13
rect 215 5 218 13
rect 210 4 213 5
rect 214 4 218 5
rect 210 3 218 4
rect 211 2 218 3
rect 220 11 228 13
rect 220 10 224 11
rect 225 10 229 11
rect 220 2 223 10
rect 226 2 229 10
rect 231 2 233 13
rect 237 12 242 13
rect 236 11 242 12
rect 243 11 250 13
rect 252 11 258 13
rect 235 10 239 11
rect 244 10 245 11
rect 235 5 238 10
rect 248 9 251 11
rect 244 8 251 9
rect 243 7 251 8
rect 243 6 246 7
rect 242 5 245 6
rect 248 5 251 7
rect 235 4 239 5
rect 241 4 242 5
rect 236 3 242 4
rect 237 2 242 3
rect 243 4 246 5
rect 247 4 251 5
rect 253 5 256 11
rect 253 4 257 5
rect 243 2 251 4
rect 254 2 258 4
rect 259 2 262 13
rect 265 12 271 13
rect 275 12 282 13
rect 265 11 272 12
rect 275 11 283 12
rect 285 11 291 13
rect 297 11 300 14
rect 303 11 306 14
rect 311 13 313 14
rect 319 13 322 14
rect 328 13 330 14
rect 337 13 340 14
rect 348 13 349 14
rect 353 13 356 14
rect 358 13 361 18
rect 363 13 364 14
rect 309 12 315 13
rect 318 12 323 13
rect 326 12 332 13
rect 308 11 315 12
rect 317 11 323 12
rect 325 11 333 12
rect 264 9 267 11
rect 269 10 273 11
rect 264 6 266 9
rect 264 5 267 6
rect 270 5 273 10
rect 274 9 278 11
rect 275 6 277 9
rect 264 4 268 5
rect 269 4 273 5
rect 274 4 277 6
rect 265 3 272 4
rect 266 2 271 3
rect 275 2 277 4
rect 280 2 283 11
rect 284 9 288 11
rect 285 8 290 9
rect 297 8 305 11
rect 308 10 311 11
rect 308 9 310 10
rect 313 9 316 11
rect 285 7 291 8
rect 287 6 291 7
rect 285 4 286 5
rect 288 4 291 6
rect 285 3 291 4
rect 285 2 290 3
rect 297 2 300 8
rect 302 7 305 8
rect 302 6 306 7
rect 307 6 316 9
rect 317 9 320 11
rect 325 10 328 11
rect 330 10 333 11
rect 335 11 342 13
rect 335 10 336 11
rect 339 10 342 11
rect 325 9 327 10
rect 331 9 333 10
rect 340 9 342 10
rect 317 8 322 9
rect 318 7 323 8
rect 320 6 324 7
rect 303 3 306 6
rect 308 5 310 6
rect 321 5 324 6
rect 308 4 311 5
rect 314 4 316 5
rect 308 3 316 4
rect 317 4 318 5
rect 320 4 324 5
rect 325 6 333 9
rect 336 8 342 9
rect 335 7 342 8
rect 325 4 328 6
rect 331 4 333 5
rect 304 2 307 3
rect 309 2 315 3
rect 317 2 323 4
rect 325 3 333 4
rect 334 4 337 7
rect 340 5 342 7
rect 339 4 342 5
rect 334 3 342 4
rect 344 11 350 13
rect 352 12 357 13
rect 351 11 357 12
rect 358 11 366 13
rect 344 10 349 11
rect 350 10 354 11
rect 358 10 362 11
rect 344 9 348 10
rect 326 2 333 3
rect 335 2 343 3
rect 344 2 347 9
rect 350 5 353 10
rect 350 4 354 5
rect 356 4 357 5
rect 351 3 357 4
rect 352 2 357 3
rect 358 2 361 10
rect 364 2 367 11
rect 373 2 376 17
rect 383 13 385 14
rect 391 13 394 14
rect 397 13 400 16
rect 403 15 406 18
rect 409 14 411 16
rect 408 13 411 14
rect 426 14 428 16
rect 594 14 597 15
rect 612 14 613 15
rect 621 14 622 15
rect 426 13 429 14
rect 434 13 437 14
rect 511 13 514 14
rect 378 12 386 13
rect 389 12 394 13
rect 378 11 387 12
rect 378 10 382 11
rect 378 2 381 10
rect 384 2 387 11
rect 388 11 394 12
rect 395 11 402 13
rect 388 10 391 11
rect 388 9 392 10
rect 388 8 394 9
rect 389 7 395 8
rect 391 6 395 7
rect 389 4 390 5
rect 392 4 395 6
rect 388 3 395 4
rect 397 4 400 11
rect 397 3 402 4
rect 388 2 394 3
rect 398 2 402 3
rect 403 2 406 13
rect 407 11 413 13
rect 409 5 411 11
rect 415 5 417 13
rect 420 5 423 13
rect 424 11 430 13
rect 433 12 438 13
rect 432 11 439 12
rect 409 4 412 5
rect 415 4 418 5
rect 419 4 423 5
rect 409 2 414 4
rect 415 3 423 4
rect 426 6 428 11
rect 432 10 434 11
rect 431 9 434 10
rect 437 10 439 11
rect 437 9 440 10
rect 431 6 440 9
rect 512 6 514 13
rect 519 12 521 14
rect 526 13 529 14
rect 534 13 536 14
rect 527 12 530 13
rect 426 4 429 6
rect 431 5 434 6
rect 512 5 515 6
rect 519 5 520 12
rect 527 11 531 12
rect 527 5 528 11
rect 529 10 532 11
rect 530 9 533 10
rect 530 8 534 9
rect 535 8 536 13
rect 531 7 536 8
rect 532 6 536 7
rect 533 5 536 6
rect 432 4 435 5
rect 438 4 439 5
rect 513 4 516 5
rect 517 4 519 5
rect 526 4 528 5
rect 534 4 536 5
rect 542 4 545 14
rect 551 12 554 14
rect 552 11 554 12
rect 558 12 560 14
rect 552 10 555 11
rect 558 10 559 12
rect 566 10 569 14
rect 571 13 573 14
rect 572 12 573 13
rect 579 13 582 14
rect 583 13 586 14
rect 593 13 594 14
rect 571 10 572 11
rect 553 9 555 10
rect 553 7 556 9
rect 557 7 558 10
rect 566 9 572 10
rect 554 5 557 7
rect 426 3 431 4
rect 432 3 439 4
rect 514 3 518 4
rect 535 3 536 4
rect 555 3 556 5
rect 566 4 569 9
rect 571 8 572 9
rect 579 9 581 13
rect 584 10 586 13
rect 592 11 594 13
rect 597 12 598 14
rect 592 10 595 11
rect 583 9 586 10
rect 593 9 597 10
rect 579 8 585 9
rect 594 8 598 9
rect 573 5 574 7
rect 572 4 574 5
rect 579 5 581 8
rect 583 7 585 8
rect 596 7 599 8
rect 583 6 586 7
rect 584 5 586 6
rect 592 5 593 6
rect 597 5 599 7
rect 579 4 582 5
rect 584 4 587 5
rect 592 4 594 5
rect 596 4 598 5
rect 604 4 607 14
rect 612 13 614 14
rect 612 11 613 13
rect 616 5 618 14
rect 620 13 622 14
rect 621 12 622 13
rect 627 12 630 14
rect 628 11 630 12
rect 633 13 635 14
rect 633 11 634 13
rect 629 10 631 11
rect 632 10 633 11
rect 629 9 633 10
rect 630 5 632 9
rect 615 4 618 5
rect 629 4 632 5
rect 586 3 588 4
rect 593 3 596 4
rect 416 2 423 3
rect 427 2 431 3
rect 433 2 439 3
<< metal2 >>
rect 591 241 619 242
rect 584 240 622 241
rect 549 239 551 240
rect 579 239 624 240
rect 546 238 556 239
rect 575 238 625 239
rect 545 237 560 238
rect 570 237 627 238
rect 544 236 629 237
rect 543 235 630 236
rect 542 234 631 235
rect 542 233 633 234
rect 542 232 634 233
rect 542 231 556 232
rect 558 231 587 232
rect 600 231 635 232
rect 542 230 551 231
rect 564 230 587 231
rect 604 230 636 231
rect 543 229 550 230
rect 566 229 590 230
rect 608 229 637 230
rect 532 228 534 229
rect 544 228 547 229
rect 567 228 594 229
rect 614 228 638 229
rect 529 227 537 228
rect 568 227 597 228
rect 622 227 639 228
rect 528 226 539 227
rect 552 226 556 227
rect 569 226 600 227
rect 626 226 640 227
rect 527 225 540 226
rect 549 225 559 226
rect 569 225 603 226
rect 630 225 641 226
rect 526 224 541 225
rect 547 224 560 225
rect 569 224 608 225
rect 633 224 642 225
rect 525 223 542 224
rect 545 223 561 224
rect 569 223 619 224
rect 636 223 642 224
rect 524 221 562 223
rect 569 222 623 223
rect 639 222 643 223
rect 569 221 626 222
rect 641 221 643 222
rect 523 220 562 221
rect 522 219 562 220
rect 568 220 629 221
rect 568 219 632 220
rect 521 218 561 219
rect 567 218 634 219
rect 520 217 561 218
rect 568 217 637 218
rect 519 216 560 217
rect 570 216 640 217
rect 518 215 559 216
rect 571 215 598 216
rect 599 215 642 216
rect 517 214 558 215
rect 573 214 598 215
rect 602 214 644 215
rect 516 213 536 214
rect 538 213 557 214
rect 574 213 598 214
rect 605 213 646 214
rect 514 212 531 213
rect 537 212 556 213
rect 575 212 598 213
rect 607 212 648 213
rect 513 211 528 212
rect 535 211 555 212
rect 577 211 599 212
rect 610 211 648 212
rect 511 210 525 211
rect 534 210 554 211
rect 578 210 599 211
rect 612 210 649 211
rect 509 209 524 210
rect 532 209 553 210
rect 579 209 600 210
rect 615 209 650 210
rect 507 208 522 209
rect 530 208 553 209
rect 505 207 520 208
rect 503 206 519 207
rect 523 206 524 207
rect 529 206 553 208
rect 561 208 562 209
rect 566 208 567 209
rect 580 208 601 209
rect 620 208 650 209
rect 561 207 571 208
rect 581 207 602 208
rect 624 207 651 208
rect 501 205 524 206
rect 528 205 553 206
rect 500 204 524 205
rect 498 203 524 204
rect 527 204 553 205
rect 562 206 573 207
rect 582 206 603 207
rect 626 206 651 207
rect 562 204 574 206
rect 582 205 605 206
rect 628 205 651 206
rect 583 204 607 205
rect 630 204 652 205
rect 527 203 554 204
rect 497 202 525 203
rect 526 202 554 203
rect 496 200 554 202
rect 495 199 554 200
rect 563 203 575 204
rect 584 203 610 204
rect 632 203 652 204
rect 563 201 576 203
rect 585 202 613 203
rect 634 202 652 203
rect 585 201 617 202
rect 635 201 652 202
rect 563 199 577 201
rect 586 200 622 201
rect 637 200 653 201
rect 586 199 624 200
rect 638 199 653 200
rect 495 198 555 199
rect 495 197 504 198
rect 505 197 555 198
rect 496 196 502 197
rect 504 196 555 197
rect 497 195 499 196
rect 503 195 555 196
rect 502 194 555 195
rect 563 197 578 199
rect 587 198 626 199
rect 639 198 653 199
rect 587 197 628 198
rect 640 197 653 198
rect 563 195 579 197
rect 588 196 629 197
rect 642 196 653 197
rect 588 195 631 196
rect 643 195 653 196
rect 501 193 554 194
rect 500 191 554 193
rect 563 193 580 195
rect 589 194 632 195
rect 644 194 653 195
rect 589 193 633 194
rect 645 193 653 194
rect 563 191 581 193
rect 590 192 635 193
rect 591 191 636 192
rect 646 191 653 193
rect 499 189 553 191
rect 562 190 582 191
rect 593 190 637 191
rect 647 190 653 191
rect 499 188 552 189
rect 562 188 583 190
rect 595 189 638 190
rect 648 189 653 190
rect 598 188 639 189
rect 500 187 552 188
rect 561 187 584 188
rect 603 187 640 188
rect 649 187 653 189
rect 500 186 551 187
rect 561 186 586 187
rect 609 186 641 187
rect 501 185 550 186
rect 561 185 587 186
rect 612 185 642 186
rect 650 185 652 187
rect 501 184 522 185
rect 525 184 550 185
rect 560 184 590 185
rect 615 184 643 185
rect 502 183 521 184
rect 526 183 549 184
rect 560 183 593 184
rect 617 183 643 184
rect 503 182 520 183
rect 527 182 548 183
rect 504 181 517 182
rect 526 181 548 182
rect 559 182 598 183
rect 620 182 644 183
rect 559 181 603 182
rect 622 181 644 182
rect 525 180 547 181
rect 558 180 606 181
rect 624 180 644 181
rect 522 179 546 180
rect 558 179 609 180
rect 625 179 644 180
rect 517 178 546 179
rect 557 178 611 179
rect 626 178 645 179
rect 508 177 545 178
rect 557 177 613 178
rect 627 177 645 178
rect 507 176 544 177
rect 556 176 615 177
rect 628 176 645 177
rect 506 175 544 176
rect 555 175 617 176
rect 629 175 645 176
rect 506 174 543 175
rect 554 174 618 175
rect 630 174 645 175
rect 506 173 542 174
rect 554 173 619 174
rect 507 172 541 173
rect 553 172 620 173
rect 631 172 645 174
rect 507 171 540 172
rect 552 171 621 172
rect 1 153 112 171
rect 132 170 245 171
rect 262 170 370 171
rect 131 153 246 170
rect 262 169 372 170
rect 262 168 374 169
rect 262 167 376 168
rect 262 166 377 167
rect 262 164 378 166
rect 262 163 379 164
rect 262 161 380 163
rect 262 156 381 161
rect 262 153 382 156
rect 1 152 36 153
rect 1 138 35 152
rect 1 137 111 138
rect 1 119 112 137
rect 1 118 36 119
rect 1 104 35 118
rect 1 97 112 104
rect 2 95 112 97
rect 3 93 112 95
rect 4 92 112 93
rect 5 90 112 92
rect 6 89 112 90
rect 8 88 112 89
rect 9 87 112 88
rect 12 86 112 87
rect 171 86 206 153
rect 262 86 297 153
rect 347 126 382 153
rect 308 125 309 126
rect 310 125 345 126
rect 346 125 381 126
rect 308 124 349 125
rect 309 123 350 124
rect 310 122 351 123
rect 311 121 352 122
rect 312 120 353 121
rect 313 119 354 120
rect 314 118 355 119
rect 315 117 356 118
rect 316 116 357 117
rect 317 115 358 116
rect 318 114 359 115
rect 319 113 360 114
rect 320 112 361 113
rect 321 111 362 112
rect 322 110 363 111
rect 323 109 364 110
rect 324 108 365 109
rect 325 107 366 108
rect 326 106 367 107
rect 327 105 368 106
rect 328 104 369 105
rect 329 103 370 104
rect 330 102 371 103
rect 331 101 372 102
rect 332 100 373 101
rect 333 99 374 100
rect 334 98 375 99
rect 335 97 376 98
rect 336 96 377 97
rect 337 95 378 96
rect 338 94 379 95
rect 339 93 380 94
rect 340 92 381 93
rect 341 91 382 92
rect 342 90 383 91
rect 343 89 384 90
rect 344 88 385 89
rect 345 87 386 88
rect 346 86 387 87
rect 407 86 441 171
rect 508 170 538 171
rect 551 170 581 171
rect 586 170 621 171
rect 632 170 645 172
rect 508 169 536 170
rect 550 169 580 170
rect 589 169 622 170
rect 509 168 534 169
rect 549 168 579 169
rect 591 168 623 169
rect 633 168 645 170
rect 510 167 532 168
rect 548 167 578 168
rect 592 167 623 168
rect 510 166 529 167
rect 546 166 578 167
rect 593 166 624 167
rect 634 166 644 168
rect 511 165 527 166
rect 545 165 577 166
rect 594 165 624 166
rect 511 164 523 165
rect 543 164 577 165
rect 595 164 624 165
rect 635 164 644 166
rect 511 163 520 164
rect 541 163 577 164
rect 596 163 624 164
rect 512 162 517 163
rect 539 162 576 163
rect 597 162 624 163
rect 636 163 644 164
rect 537 161 576 162
rect 585 161 586 162
rect 598 161 625 162
rect 636 161 643 163
rect 535 160 576 161
rect 584 160 587 161
rect 598 160 624 161
rect 532 159 575 160
rect 584 159 588 160
rect 530 158 575 159
rect 583 158 588 159
rect 599 158 624 160
rect 637 160 643 161
rect 637 158 642 160
rect 528 157 574 158
rect 583 157 589 158
rect 526 156 574 157
rect 524 155 573 156
rect 582 155 590 157
rect 600 156 624 158
rect 638 156 641 158
rect 522 154 573 155
rect 521 153 572 154
rect 581 153 591 155
rect 600 154 623 156
rect 638 155 640 156
rect 638 154 639 155
rect 601 153 622 154
rect 520 152 571 153
rect 519 151 571 152
rect 518 150 570 151
rect 580 150 592 153
rect 601 152 621 153
rect 601 150 620 152
rect 517 149 569 150
rect 516 148 568 149
rect 579 148 593 150
rect 516 147 567 148
rect 578 147 593 148
rect 515 146 566 147
rect 515 145 565 146
rect 577 145 593 147
rect 602 149 619 150
rect 602 148 618 149
rect 602 147 617 148
rect 630 147 631 148
rect 602 146 615 147
rect 629 146 632 147
rect 602 145 614 146
rect 628 145 632 146
rect 514 144 564 145
rect 576 144 594 145
rect 514 143 563 144
rect 513 142 562 143
rect 575 142 594 144
rect 513 141 561 142
rect 574 141 594 142
rect 513 140 559 141
rect 573 140 594 141
rect 602 144 612 145
rect 627 144 632 145
rect 602 143 611 144
rect 626 143 632 144
rect 602 142 609 143
rect 625 142 632 143
rect 602 141 607 142
rect 624 141 632 142
rect 602 140 605 141
rect 623 140 632 141
rect 513 139 558 140
rect 572 139 594 140
rect 621 139 632 140
rect 512 138 556 139
rect 571 138 594 139
rect 620 138 632 139
rect 512 137 554 138
rect 569 137 594 138
rect 618 137 632 138
rect 512 136 553 137
rect 568 136 594 137
rect 617 136 632 137
rect 512 135 550 136
rect 567 135 593 136
rect 615 135 632 136
rect 512 134 548 135
rect 565 134 593 135
rect 613 134 632 135
rect 512 133 546 134
rect 563 133 593 134
rect 612 133 632 134
rect 512 132 544 133
rect 562 132 593 133
rect 610 132 632 133
rect 512 131 541 132
rect 560 131 593 132
rect 607 131 632 132
rect 512 130 539 131
rect 558 130 592 131
rect 605 130 632 131
rect 513 129 538 130
rect 556 129 592 130
rect 602 129 631 130
rect 513 128 536 129
rect 554 128 592 129
rect 599 128 631 129
rect 513 127 535 128
rect 552 127 592 128
rect 595 127 631 128
rect 513 126 534 127
rect 550 126 631 127
rect 513 125 533 126
rect 549 125 630 126
rect 514 124 532 125
rect 547 124 630 125
rect 514 122 531 124
rect 546 123 630 124
rect 544 122 629 123
rect 515 120 530 122
rect 543 121 629 122
rect 542 120 629 121
rect 516 118 529 120
rect 541 119 628 120
rect 540 118 572 119
rect 574 118 628 119
rect 517 116 529 118
rect 539 117 570 118
rect 574 117 627 118
rect 538 116 569 117
rect 573 116 627 117
rect 518 114 528 116
rect 537 115 567 116
rect 573 115 626 116
rect 537 114 566 115
rect 519 113 528 114
rect 520 111 528 113
rect 536 113 564 114
rect 572 113 625 115
rect 536 112 563 113
rect 571 112 624 113
rect 521 110 528 111
rect 535 111 561 112
rect 570 111 623 112
rect 535 110 560 111
rect 569 110 623 111
rect 522 109 527 110
rect 523 108 527 109
rect 524 107 527 108
rect 534 109 559 110
rect 569 109 592 110
rect 594 109 622 110
rect 534 108 558 109
rect 568 108 591 109
rect 593 108 621 109
rect 534 107 557 108
rect 567 107 590 108
rect 593 107 620 108
rect 525 106 527 107
rect 526 105 527 106
rect 533 106 556 107
rect 566 106 588 107
rect 533 105 555 106
rect 566 105 587 106
rect 592 105 619 107
rect 533 103 554 105
rect 565 104 586 105
rect 592 104 618 105
rect 565 103 585 104
rect 592 103 617 104
rect 532 102 553 103
rect 564 102 585 103
rect 591 102 616 103
rect 532 100 552 102
rect 564 101 584 102
rect 591 101 615 102
rect 532 98 551 100
rect 563 99 583 101
rect 591 100 613 101
rect 591 99 612 100
rect 533 97 551 98
rect 562 98 582 99
rect 591 98 611 99
rect 533 95 550 97
rect 562 95 581 98
rect 591 97 610 98
rect 590 96 609 97
rect 590 95 607 96
rect 534 93 550 95
rect 535 92 550 93
rect 536 91 550 92
rect 537 89 550 91
rect 538 88 550 89
rect 540 87 550 88
rect 541 86 550 87
rect 16 85 111 86
rect 172 85 205 86
rect 347 85 388 86
rect 408 85 441 86
rect 542 85 550 86
rect 348 84 389 85
rect 544 84 550 85
rect 349 83 390 84
rect 545 83 550 84
rect 561 92 580 95
rect 590 94 606 95
rect 590 93 605 94
rect 590 92 603 93
rect 561 87 579 92
rect 590 91 602 92
rect 590 90 601 91
rect 590 89 600 90
rect 591 88 599 89
rect 591 87 598 88
rect 350 82 391 83
rect 546 82 551 83
rect 561 82 578 87
rect 591 85 597 87
rect 591 84 596 85
rect 591 83 595 84
rect 351 81 392 82
rect 547 81 551 82
rect 352 80 393 81
rect 549 80 551 81
rect 550 79 551 80
rect 562 79 578 82
rect 592 82 595 83
rect 592 80 594 82
rect 592 79 593 80
rect 563 78 578 79
rect 563 77 579 78
rect 564 75 579 77
rect 565 74 579 75
rect 566 73 579 74
rect 567 72 579 73
rect 568 71 580 72
rect 569 70 580 71
rect 570 69 580 70
rect 571 68 581 69
rect 572 67 581 68
rect 573 66 581 67
rect 575 65 582 66
rect 9 64 21 65
rect 30 64 34 65
rect 133 64 137 65
rect 9 61 22 64
rect 9 60 21 61
rect 4 54 27 59
rect 30 53 35 64
rect 57 58 85 63
rect 79 55 85 58
rect 107 57 126 62
rect 113 56 119 57
rect 132 56 137 64
rect 181 64 185 65
rect 156 60 176 61
rect 156 56 177 60
rect 114 55 119 56
rect 126 55 137 56
rect 163 55 169 56
rect 36 53 38 54
rect 12 52 19 53
rect 9 51 22 52
rect 7 50 23 51
rect 6 49 24 50
rect 6 48 25 49
rect 5 47 12 48
rect 19 47 25 48
rect 5 44 11 47
rect 20 45 25 47
rect 30 48 39 53
rect 79 52 84 55
rect 113 54 119 55
rect 113 52 120 54
rect 78 49 84 52
rect 112 51 121 52
rect 125 51 137 55
rect 164 53 169 55
rect 112 50 122 51
rect 111 49 123 50
rect 20 44 26 45
rect 5 43 12 44
rect 18 43 25 44
rect 6 42 25 43
rect 7 41 24 42
rect 8 40 23 41
rect 10 39 21 40
rect 9 36 14 37
rect 30 36 35 48
rect 53 45 89 49
rect 110 48 124 49
rect 109 47 116 48
rect 117 47 125 48
rect 107 46 116 47
rect 118 46 127 47
rect 106 45 115 46
rect 119 45 127 46
rect 54 44 89 45
rect 104 44 114 45
rect 120 44 127 45
rect 68 38 73 44
rect 105 43 113 44
rect 121 43 126 44
rect 106 42 111 43
rect 123 42 125 43
rect 107 41 110 42
rect 9 31 15 36
rect 30 35 34 36
rect 57 33 85 38
rect 9 30 35 31
rect 9 26 36 30
rect 80 25 85 33
rect 111 31 116 39
rect 132 36 137 51
rect 163 50 169 53
rect 181 50 186 64
rect 209 60 236 64
rect 265 63 269 64
rect 265 60 270 63
rect 209 59 215 60
rect 233 59 234 60
rect 209 58 214 59
rect 209 57 235 58
rect 209 54 236 57
rect 264 55 270 60
rect 209 53 215 54
rect 264 53 271 55
rect 209 52 214 53
rect 263 52 271 53
rect 209 51 215 52
rect 262 51 272 52
rect 163 47 170 50
rect 162 46 170 47
rect 181 49 187 50
rect 189 49 190 50
rect 162 45 171 46
rect 161 44 171 45
rect 181 44 191 49
rect 209 47 236 51
rect 262 50 273 51
rect 261 49 274 50
rect 260 48 267 49
rect 268 48 275 49
rect 259 47 266 48
rect 268 47 276 48
rect 219 45 225 47
rect 258 46 265 47
rect 269 46 278 47
rect 256 45 265 46
rect 270 45 279 46
rect 205 44 239 45
rect 255 44 264 45
rect 271 44 279 45
rect 161 43 172 44
rect 160 42 172 43
rect 160 41 166 42
rect 159 40 166 41
rect 167 41 173 42
rect 167 40 174 41
rect 158 39 165 40
rect 168 39 175 40
rect 157 38 164 39
rect 156 37 164 38
rect 169 38 176 39
rect 169 37 177 38
rect 155 36 163 37
rect 170 36 178 37
rect 154 35 162 36
rect 171 35 177 36
rect 154 34 161 35
rect 172 34 177 35
rect 155 33 160 34
rect 174 33 176 34
rect 156 32 159 33
rect 111 26 138 31
rect 181 25 186 44
rect 204 40 240 44
rect 255 43 263 44
rect 273 43 278 44
rect 256 42 261 43
rect 274 42 277 43
rect 257 41 260 42
rect 258 40 259 41
rect 262 38 266 39
rect 214 37 230 38
rect 211 36 233 37
rect 210 35 234 36
rect 209 34 236 35
rect 208 33 217 34
rect 227 33 236 34
rect 208 30 214 33
rect 230 32 237 33
rect 231 31 237 32
rect 230 30 237 31
rect 262 31 267 38
rect 283 36 288 65
rect 317 63 318 64
rect 312 62 321 63
rect 311 61 323 62
rect 310 60 324 61
rect 333 60 338 65
rect 414 64 425 65
rect 413 63 426 64
rect 309 59 338 60
rect 308 58 316 59
rect 317 58 338 59
rect 359 58 387 63
rect 412 62 427 63
rect 411 61 428 62
rect 308 57 314 58
rect 320 57 338 58
rect 307 56 313 57
rect 307 51 312 56
rect 321 55 338 57
rect 321 54 327 55
rect 322 52 327 54
rect 333 52 338 55
rect 307 49 313 51
rect 321 50 338 52
rect 381 54 387 58
rect 410 60 417 61
rect 422 60 429 61
rect 410 59 416 60
rect 423 59 429 60
rect 410 56 415 59
rect 424 56 429 59
rect 410 55 417 56
rect 422 55 429 56
rect 410 54 428 55
rect 381 50 386 54
rect 411 53 428 54
rect 412 52 427 53
rect 414 51 425 52
rect 417 50 423 51
rect 320 49 338 50
rect 308 48 314 49
rect 319 48 338 49
rect 308 47 338 48
rect 309 46 325 47
rect 310 45 324 46
rect 311 44 322 45
rect 313 43 320 44
rect 312 31 317 39
rect 333 36 338 47
rect 380 49 386 50
rect 431 49 433 50
rect 380 46 385 49
rect 355 42 391 46
rect 407 45 433 49
rect 407 44 431 45
rect 356 41 391 42
rect 415 43 421 44
rect 262 30 288 31
rect 208 29 216 30
rect 228 29 236 30
rect 209 28 236 29
rect 210 27 235 28
rect 211 26 234 27
rect 262 26 289 30
rect 312 26 339 31
rect 213 25 231 26
rect 370 25 375 41
rect 415 37 420 43
rect 427 42 428 43
rect 429 42 433 43
rect 434 42 439 65
rect 577 64 582 65
rect 578 63 582 64
rect 580 62 583 63
rect 472 44 482 46
rect 485 44 494 46
rect 497 44 507 46
rect 511 44 519 46
rect 522 44 532 46
rect 537 44 546 46
rect 548 44 555 46
rect 564 44 572 46
rect 583 45 594 46
rect 580 44 586 45
rect 589 44 595 45
rect 608 44 618 46
rect 622 44 632 46
rect 637 44 653 46
rect 658 44 675 46
rect 474 43 480 44
rect 487 43 491 44
rect 499 43 505 44
rect 426 38 439 42
rect 413 31 418 36
rect 434 35 439 38
rect 475 35 479 43
rect 487 42 489 43
rect 500 42 505 43
rect 513 43 516 44
rect 524 43 530 44
rect 539 43 544 44
rect 551 43 556 44
rect 513 42 515 43
rect 486 41 488 42
rect 485 40 487 41
rect 501 40 506 42
rect 512 41 515 42
rect 512 40 514 41
rect 484 39 486 40
rect 483 38 485 39
rect 502 38 507 40
rect 511 38 513 40
rect 482 37 484 38
rect 503 37 508 38
rect 481 36 484 37
rect 504 36 508 37
rect 510 36 512 38
rect 480 35 485 36
rect 504 35 511 36
rect 475 34 486 35
rect 413 26 440 31
rect 475 26 479 34
rect 480 33 486 34
rect 505 34 511 35
rect 481 32 487 33
rect 482 31 488 32
rect 483 30 488 31
rect 483 29 489 30
rect 484 28 490 29
rect 485 27 491 28
rect 485 26 492 27
rect 474 25 480 26
rect 486 25 493 26
rect 505 25 510 34
rect 524 31 529 43
rect 525 30 529 31
rect 525 27 530 30
rect 540 29 543 43
rect 551 42 557 43
rect 551 41 558 42
rect 551 40 559 41
rect 567 40 570 44
rect 579 43 584 44
rect 591 43 595 44
rect 610 43 616 44
rect 624 43 630 44
rect 578 42 582 43
rect 592 42 595 43
rect 577 41 582 42
rect 593 41 595 42
rect 576 40 581 41
rect 539 27 542 29
rect 526 26 531 27
rect 538 26 542 27
rect 551 27 553 40
rect 554 39 560 40
rect 554 38 561 39
rect 555 37 562 38
rect 556 36 562 37
rect 557 35 563 36
rect 558 34 564 35
rect 559 33 565 34
rect 560 32 566 33
rect 560 31 567 32
rect 568 31 569 40
rect 575 37 580 40
rect 594 39 595 41
rect 611 42 616 43
rect 574 32 580 37
rect 611 36 615 42
rect 625 36 630 43
rect 611 34 630 36
rect 587 33 597 34
rect 588 32 596 33
rect 561 30 569 31
rect 562 29 569 30
rect 575 30 580 32
rect 590 31 595 32
rect 575 29 581 30
rect 563 28 569 29
rect 564 27 569 28
rect 576 28 581 29
rect 576 27 582 28
rect 526 25 533 26
rect 537 25 541 26
rect 551 25 554 27
rect 565 25 569 27
rect 577 26 582 27
rect 591 26 595 31
rect 611 26 615 34
rect 578 25 584 26
rect 218 24 227 25
rect 472 23 482 25
rect 487 23 495 25
rect 503 24 513 25
rect 527 24 540 25
rect 549 24 556 25
rect 566 24 569 25
rect 580 24 586 25
rect 590 24 595 26
rect 610 25 616 26
rect 625 25 630 34
rect 639 36 644 44
rect 650 43 653 44
rect 651 42 653 43
rect 652 40 653 42
rect 650 36 651 38
rect 639 34 651 36
rect 639 25 644 34
rect 649 33 651 34
rect 650 31 651 33
rect 661 36 666 44
rect 672 43 675 44
rect 673 40 675 43
rect 672 37 673 38
rect 671 36 673 37
rect 661 34 673 36
rect 653 27 655 29
rect 652 26 655 27
rect 651 25 654 26
rect 661 25 666 34
rect 671 32 673 34
rect 672 31 673 32
rect 675 28 677 29
rect 674 26 676 28
rect 673 25 676 26
rect 502 23 514 24
rect 529 23 539 24
rect 548 23 557 24
rect 567 23 569 24
rect 582 23 594 24
rect 608 23 618 25
rect 622 23 632 25
rect 636 23 654 25
rect 658 24 676 25
rect 658 23 675 24
rect 15 17 17 18
rect 122 17 123 18
rect 149 17 150 18
rect 360 17 361 18
rect 5 14 13 16
rect 5 10 8 14
rect 5 7 12 10
rect 5 4 8 7
rect 5 3 12 4
rect 5 1 13 3
rect 14 1 17 17
rect 22 12 24 13
rect 31 12 34 13
rect 37 12 40 15
rect 70 14 73 17
rect 47 12 48 13
rect 52 12 55 13
rect 64 12 66 13
rect 78 12 80 13
rect 85 12 87 13
rect 97 12 100 13
rect 109 12 111 13
rect 118 12 119 13
rect 121 12 124 17
rect 129 14 139 16
rect 132 13 136 14
rect 20 11 26 12
rect 30 11 42 12
rect 19 10 26 11
rect 29 10 42 11
rect 43 10 49 12
rect 51 11 57 12
rect 50 10 57 11
rect 60 10 68 12
rect 19 9 22 10
rect 19 8 21 9
rect 24 8 27 10
rect 19 5 27 8
rect 28 9 32 10
rect 19 4 21 5
rect 28 4 31 9
rect 19 3 22 4
rect 25 3 26 4
rect 29 3 32 4
rect 34 3 35 4
rect 19 2 27 3
rect 29 2 35 3
rect 37 3 40 10
rect 43 9 53 10
rect 37 2 42 3
rect 20 1 26 2
rect 30 1 35 2
rect 38 1 42 2
rect 43 1 46 9
rect 49 4 52 9
rect 55 8 58 10
rect 56 6 58 8
rect 55 4 58 6
rect 49 3 53 4
rect 54 3 58 4
rect 50 2 57 3
rect 51 1 56 2
rect 60 1 63 10
rect 65 9 68 10
rect 66 1 68 9
rect 70 1 73 12
rect 76 11 81 12
rect 83 11 89 12
rect 96 11 102 12
rect 105 11 112 12
rect 116 11 124 12
rect 75 10 81 11
rect 82 10 89 11
rect 95 10 103 11
rect 75 7 78 10
rect 82 8 85 10
rect 95 9 97 10
rect 100 8 103 10
rect 82 7 87 8
rect 96 7 103 8
rect 75 6 77 7
rect 83 6 88 7
rect 95 6 103 7
rect 75 4 78 6
rect 85 5 89 6
rect 95 5 98 6
rect 75 3 79 4
rect 80 3 81 4
rect 83 3 84 4
rect 86 3 89 5
rect 94 4 97 5
rect 100 4 103 6
rect 75 2 89 3
rect 95 3 98 4
rect 99 3 103 4
rect 95 2 103 3
rect 76 1 88 2
rect 96 1 103 2
rect 105 10 113 11
rect 105 8 108 10
rect 105 1 107 8
rect 110 1 113 10
rect 115 10 124 11
rect 115 7 118 10
rect 120 8 124 10
rect 115 6 117 7
rect 115 4 118 6
rect 121 5 124 8
rect 115 3 119 4
rect 120 3 124 5
rect 115 2 124 3
rect 116 1 124 2
rect 133 1 136 13
rect 141 12 143 13
rect 139 11 145 12
rect 138 10 145 11
rect 138 9 141 10
rect 138 8 140 9
rect 143 8 146 10
rect 137 5 146 8
rect 138 4 140 5
rect 138 3 141 4
rect 144 3 146 4
rect 138 2 146 3
rect 139 1 145 2
rect 148 1 150 17
rect 232 14 234 17
rect 255 14 257 15
rect 260 14 263 17
rect 298 15 306 16
rect 298 14 307 15
rect 155 12 157 13
rect 165 12 167 13
rect 173 12 175 13
rect 184 12 186 13
rect 189 12 191 13
rect 199 12 201 13
rect 205 12 207 13
rect 225 12 228 13
rect 239 12 242 13
rect 246 12 249 13
rect 254 12 257 14
rect 298 13 302 14
rect 303 13 307 14
rect 268 12 271 13
rect 280 12 282 13
rect 288 12 291 13
rect 153 11 159 12
rect 163 11 168 12
rect 171 11 177 12
rect 180 11 187 12
rect 188 11 193 12
rect 153 10 160 11
rect 152 8 155 10
rect 157 9 160 10
rect 162 10 168 11
rect 170 10 178 11
rect 162 9 165 10
rect 169 9 173 10
rect 158 8 160 9
rect 152 5 160 8
rect 161 5 164 9
rect 152 4 155 5
rect 161 4 165 5
rect 169 4 172 9
rect 175 8 178 10
rect 180 10 193 11
rect 176 5 179 8
rect 152 3 156 4
rect 158 3 160 4
rect 153 2 160 3
rect 162 3 166 4
rect 167 3 168 4
rect 169 3 173 4
rect 175 3 178 5
rect 162 2 168 3
rect 170 2 178 3
rect 154 1 160 2
rect 163 1 168 2
rect 171 1 177 2
rect 180 1 183 10
rect 185 9 189 10
rect 190 9 193 10
rect 185 1 188 9
rect 191 1 193 9
rect 195 10 208 12
rect 195 9 199 10
rect 195 1 198 9
rect 200 8 204 10
rect 201 1 203 8
rect 206 1 209 10
rect 211 4 213 12
rect 216 4 219 12
rect 211 3 214 4
rect 215 3 219 4
rect 211 2 219 3
rect 212 1 219 2
rect 221 10 229 12
rect 221 9 225 10
rect 226 9 230 10
rect 221 1 224 9
rect 227 1 230 9
rect 232 1 234 12
rect 238 11 243 12
rect 237 10 243 11
rect 244 10 251 12
rect 253 10 259 12
rect 236 9 240 10
rect 245 9 246 10
rect 236 4 239 9
rect 249 8 252 10
rect 245 7 252 8
rect 244 6 252 7
rect 244 5 247 6
rect 243 4 246 5
rect 249 4 252 6
rect 236 3 240 4
rect 242 3 243 4
rect 237 2 243 3
rect 238 1 243 2
rect 244 3 247 4
rect 248 3 252 4
rect 254 4 257 10
rect 254 3 258 4
rect 244 1 252 3
rect 255 1 259 3
rect 260 1 263 12
rect 266 11 272 12
rect 276 11 283 12
rect 266 10 273 11
rect 276 10 284 11
rect 286 10 292 12
rect 298 10 301 13
rect 304 10 307 13
rect 312 12 314 13
rect 320 12 323 13
rect 329 12 331 13
rect 338 12 341 13
rect 349 12 350 13
rect 354 12 357 13
rect 359 12 362 17
rect 364 12 365 13
rect 310 11 316 12
rect 319 11 324 12
rect 327 11 333 12
rect 309 10 316 11
rect 318 10 324 11
rect 326 10 334 11
rect 265 8 268 10
rect 270 9 274 10
rect 265 5 267 8
rect 265 4 268 5
rect 271 4 274 9
rect 275 8 279 10
rect 276 5 278 8
rect 265 3 269 4
rect 270 3 274 4
rect 275 3 278 5
rect 266 2 273 3
rect 267 1 272 2
rect 276 1 278 3
rect 281 1 284 10
rect 285 8 289 10
rect 286 7 291 8
rect 298 7 306 10
rect 309 9 312 10
rect 309 8 311 9
rect 314 8 317 10
rect 286 6 292 7
rect 288 5 292 6
rect 286 3 287 4
rect 289 3 292 5
rect 286 2 292 3
rect 286 1 291 2
rect 298 1 301 7
rect 303 6 306 7
rect 303 5 307 6
rect 308 5 317 8
rect 318 8 321 10
rect 326 9 329 10
rect 331 9 334 10
rect 336 10 343 12
rect 336 9 337 10
rect 340 9 343 10
rect 326 8 328 9
rect 332 8 334 9
rect 341 8 343 9
rect 318 7 323 8
rect 319 6 324 7
rect 321 5 325 6
rect 304 2 307 5
rect 309 4 311 5
rect 322 4 325 5
rect 309 3 312 4
rect 315 3 317 4
rect 309 2 317 3
rect 318 3 319 4
rect 321 3 325 4
rect 326 5 334 8
rect 337 7 343 8
rect 336 6 343 7
rect 326 3 329 5
rect 332 3 334 4
rect 305 1 308 2
rect 310 1 316 2
rect 318 1 324 3
rect 326 2 334 3
rect 335 3 338 6
rect 341 4 343 6
rect 340 3 343 4
rect 335 2 343 3
rect 345 10 351 12
rect 353 11 358 12
rect 352 10 358 11
rect 359 10 367 12
rect 345 9 350 10
rect 351 9 355 10
rect 359 9 363 10
rect 345 8 349 9
rect 327 1 334 2
rect 336 1 344 2
rect 345 1 348 8
rect 351 4 354 9
rect 351 3 355 4
rect 357 3 358 4
rect 352 2 358 3
rect 353 1 358 2
rect 359 1 362 9
rect 365 1 368 10
rect 374 1 377 16
rect 384 12 386 13
rect 392 12 395 13
rect 398 12 401 15
rect 404 14 407 17
rect 410 13 412 15
rect 409 12 412 13
rect 427 13 429 15
rect 595 13 598 14
rect 613 13 614 14
rect 622 13 623 14
rect 427 12 430 13
rect 435 12 438 13
rect 512 12 515 13
rect 379 11 387 12
rect 390 11 395 12
rect 379 10 388 11
rect 379 9 383 10
rect 379 1 382 9
rect 385 1 388 10
rect 389 10 395 11
rect 396 10 403 12
rect 389 9 392 10
rect 389 8 393 9
rect 389 7 395 8
rect 390 6 396 7
rect 392 5 396 6
rect 390 3 391 4
rect 393 3 396 5
rect 389 2 396 3
rect 398 3 401 10
rect 398 2 403 3
rect 389 1 395 2
rect 399 1 403 2
rect 404 1 407 12
rect 408 10 414 12
rect 410 4 412 10
rect 416 4 418 12
rect 421 4 424 12
rect 425 10 431 12
rect 434 11 439 12
rect 433 10 440 11
rect 410 3 413 4
rect 416 3 419 4
rect 420 3 424 4
rect 410 1 415 3
rect 416 2 424 3
rect 427 5 429 10
rect 433 9 435 10
rect 432 8 435 9
rect 438 9 440 10
rect 438 8 441 9
rect 432 5 441 8
rect 513 5 515 12
rect 520 11 522 13
rect 527 12 530 13
rect 535 12 537 13
rect 528 11 531 12
rect 427 3 430 5
rect 432 4 435 5
rect 513 4 516 5
rect 520 4 521 11
rect 528 10 532 11
rect 528 4 529 10
rect 530 9 533 10
rect 531 8 534 9
rect 531 7 535 8
rect 536 7 537 12
rect 532 6 537 7
rect 533 5 537 6
rect 534 4 537 5
rect 433 3 436 4
rect 439 3 440 4
rect 514 3 517 4
rect 518 3 520 4
rect 527 3 529 4
rect 535 3 537 4
rect 543 3 546 13
rect 552 11 555 13
rect 553 10 555 11
rect 559 11 561 13
rect 553 9 556 10
rect 559 9 560 11
rect 567 9 570 13
rect 572 12 574 13
rect 573 11 574 12
rect 580 12 583 13
rect 584 12 587 13
rect 594 12 595 13
rect 572 9 573 10
rect 554 8 556 9
rect 554 6 557 8
rect 558 6 559 9
rect 567 8 573 9
rect 555 4 558 6
rect 427 2 432 3
rect 433 2 440 3
rect 515 2 519 3
rect 536 2 537 3
rect 556 2 557 4
rect 567 3 570 8
rect 572 7 573 8
rect 580 8 582 12
rect 585 9 587 12
rect 593 10 595 12
rect 598 11 599 13
rect 593 9 596 10
rect 584 8 587 9
rect 594 8 598 9
rect 580 7 586 8
rect 595 7 599 8
rect 574 4 575 6
rect 573 3 575 4
rect 580 4 582 7
rect 584 6 586 7
rect 597 6 600 7
rect 584 5 587 6
rect 585 4 587 5
rect 593 4 594 5
rect 598 4 600 6
rect 580 3 583 4
rect 585 3 588 4
rect 593 3 595 4
rect 597 3 599 4
rect 605 3 608 13
rect 613 12 615 13
rect 613 10 614 12
rect 617 4 619 13
rect 621 12 623 13
rect 622 11 623 12
rect 628 11 631 13
rect 629 10 631 11
rect 634 12 636 13
rect 634 10 635 12
rect 630 9 632 10
rect 633 9 634 10
rect 630 8 634 9
rect 631 4 633 8
rect 616 3 619 4
rect 630 3 633 4
rect 587 2 589 3
rect 594 2 597 3
rect 417 1 424 2
rect 428 1 432 2
rect 434 1 440 2
<< metal3 >>
rect 592 240 620 241
rect 585 239 623 240
rect 550 238 552 239
rect 580 238 625 239
rect 547 237 557 238
rect 576 237 626 238
rect 546 236 561 237
rect 571 236 628 237
rect 545 235 630 236
rect 544 234 631 235
rect 543 233 632 234
rect 543 232 634 233
rect 543 231 635 232
rect 543 230 557 231
rect 559 230 588 231
rect 601 230 636 231
rect 543 229 552 230
rect 565 229 588 230
rect 605 229 637 230
rect 544 228 551 229
rect 567 228 591 229
rect 609 228 638 229
rect 533 227 535 228
rect 545 227 548 228
rect 568 227 595 228
rect 615 227 639 228
rect 530 226 538 227
rect 569 226 598 227
rect 623 226 640 227
rect 529 225 540 226
rect 553 225 557 226
rect 570 225 601 226
rect 627 225 641 226
rect 528 224 541 225
rect 550 224 560 225
rect 570 224 604 225
rect 631 224 642 225
rect 527 223 542 224
rect 548 223 561 224
rect 570 223 609 224
rect 634 223 643 224
rect 526 222 543 223
rect 546 222 562 223
rect 570 222 620 223
rect 637 222 643 223
rect 525 220 563 222
rect 570 221 624 222
rect 640 221 644 222
rect 570 220 627 221
rect 642 220 644 221
rect 524 219 563 220
rect 523 218 563 219
rect 569 219 630 220
rect 569 218 633 219
rect 522 217 562 218
rect 568 217 635 218
rect 521 216 562 217
rect 569 216 638 217
rect 520 215 561 216
rect 571 215 641 216
rect 519 214 560 215
rect 572 214 599 215
rect 600 214 643 215
rect 518 213 559 214
rect 574 213 599 214
rect 603 213 645 214
rect 517 212 537 213
rect 539 212 558 213
rect 575 212 599 213
rect 606 212 647 213
rect 515 211 532 212
rect 538 211 557 212
rect 576 211 599 212
rect 608 211 649 212
rect 514 210 529 211
rect 536 210 556 211
rect 578 210 600 211
rect 611 210 649 211
rect 512 209 526 210
rect 535 209 555 210
rect 579 209 600 210
rect 613 209 650 210
rect 510 208 525 209
rect 533 208 554 209
rect 580 208 601 209
rect 616 208 651 209
rect 508 207 523 208
rect 531 207 554 208
rect 506 206 521 207
rect 504 205 520 206
rect 524 205 525 206
rect 530 205 554 207
rect 562 207 563 208
rect 567 207 568 208
rect 581 207 602 208
rect 621 207 651 208
rect 562 206 572 207
rect 582 206 603 207
rect 625 206 652 207
rect 502 204 525 205
rect 529 204 554 205
rect 501 203 525 204
rect 499 202 525 203
rect 528 203 554 204
rect 563 205 574 206
rect 583 205 604 206
rect 627 205 652 206
rect 563 203 575 205
rect 583 204 606 205
rect 629 204 652 205
rect 584 203 608 204
rect 631 203 653 204
rect 528 202 555 203
rect 498 201 526 202
rect 527 201 555 202
rect 497 199 555 201
rect 496 198 555 199
rect 564 202 576 203
rect 585 202 611 203
rect 633 202 653 203
rect 564 200 577 202
rect 586 201 614 202
rect 635 201 653 202
rect 586 200 618 201
rect 636 200 653 201
rect 564 198 578 200
rect 587 199 623 200
rect 638 199 654 200
rect 587 198 625 199
rect 639 198 654 199
rect 496 197 556 198
rect 496 196 505 197
rect 506 196 556 197
rect 497 195 503 196
rect 505 195 556 196
rect 498 194 500 195
rect 504 194 556 195
rect 503 193 556 194
rect 564 196 579 198
rect 588 197 627 198
rect 640 197 654 198
rect 588 196 629 197
rect 641 196 654 197
rect 564 194 580 196
rect 589 195 630 196
rect 643 195 654 196
rect 589 194 632 195
rect 644 194 654 195
rect 502 192 555 193
rect 501 190 555 192
rect 564 192 581 194
rect 590 193 633 194
rect 645 193 654 194
rect 590 192 634 193
rect 646 192 654 193
rect 564 190 582 192
rect 591 191 636 192
rect 592 190 637 191
rect 647 190 654 192
rect 500 188 554 190
rect 563 189 583 190
rect 594 189 638 190
rect 648 189 654 190
rect 500 187 553 188
rect 563 187 584 189
rect 596 188 639 189
rect 649 188 654 189
rect 599 187 640 188
rect 501 186 553 187
rect 562 186 585 187
rect 604 186 641 187
rect 650 186 654 188
rect 501 185 552 186
rect 562 185 587 186
rect 610 185 642 186
rect 502 184 551 185
rect 562 184 588 185
rect 613 184 643 185
rect 651 184 653 186
rect 502 183 523 184
rect 526 183 551 184
rect 561 183 591 184
rect 616 183 644 184
rect 503 182 522 183
rect 527 182 550 183
rect 561 182 594 183
rect 618 182 644 183
rect 504 181 521 182
rect 528 181 549 182
rect 505 180 518 181
rect 527 180 549 181
rect 560 181 599 182
rect 621 181 645 182
rect 560 180 604 181
rect 623 180 645 181
rect 526 179 548 180
rect 559 179 607 180
rect 625 179 645 180
rect 523 178 547 179
rect 559 178 610 179
rect 626 178 645 179
rect 518 177 547 178
rect 558 177 612 178
rect 627 177 646 178
rect 509 176 546 177
rect 558 176 614 177
rect 628 176 646 177
rect 508 175 545 176
rect 557 175 616 176
rect 629 175 646 176
rect 507 174 545 175
rect 556 174 618 175
rect 630 174 646 175
rect 507 173 544 174
rect 555 173 619 174
rect 631 173 646 174
rect 507 172 543 173
rect 555 172 620 173
rect 508 171 542 172
rect 554 171 621 172
rect 632 171 646 173
rect 508 170 541 171
rect 553 170 622 171
rect 2 152 113 170
rect 133 169 246 170
rect 263 169 371 170
rect 132 152 247 169
rect 263 168 373 169
rect 263 167 375 168
rect 263 166 377 167
rect 263 165 378 166
rect 263 163 379 165
rect 263 162 380 163
rect 263 160 381 162
rect 263 155 382 160
rect 263 152 383 155
rect 2 151 37 152
rect 2 137 36 151
rect 2 136 112 137
rect 2 118 113 136
rect 2 117 37 118
rect 2 103 36 117
rect 2 96 113 103
rect 3 94 113 96
rect 4 92 113 94
rect 5 91 113 92
rect 6 89 113 91
rect 7 88 113 89
rect 9 87 113 88
rect 10 86 113 87
rect 13 85 113 86
rect 172 85 207 152
rect 263 85 298 152
rect 348 125 383 152
rect 309 124 310 125
rect 311 124 346 125
rect 347 124 382 125
rect 309 123 350 124
rect 310 122 351 123
rect 311 121 352 122
rect 312 120 353 121
rect 313 119 354 120
rect 314 118 355 119
rect 315 117 356 118
rect 316 116 357 117
rect 317 115 358 116
rect 318 114 359 115
rect 319 113 360 114
rect 320 112 361 113
rect 321 111 362 112
rect 322 110 363 111
rect 323 109 364 110
rect 324 108 365 109
rect 325 107 366 108
rect 326 106 367 107
rect 327 105 368 106
rect 328 104 369 105
rect 329 103 370 104
rect 330 102 371 103
rect 331 101 372 102
rect 332 100 373 101
rect 333 99 374 100
rect 334 98 375 99
rect 335 97 376 98
rect 336 96 377 97
rect 337 95 378 96
rect 338 94 379 95
rect 339 93 380 94
rect 340 92 381 93
rect 341 91 382 92
rect 342 90 383 91
rect 343 89 384 90
rect 344 88 385 89
rect 345 87 386 88
rect 346 86 387 87
rect 347 85 388 86
rect 408 85 442 170
rect 509 169 539 170
rect 552 169 582 170
rect 587 169 622 170
rect 633 169 646 171
rect 509 168 537 169
rect 551 168 581 169
rect 590 168 623 169
rect 510 167 535 168
rect 550 167 580 168
rect 592 167 624 168
rect 634 167 646 169
rect 511 166 533 167
rect 549 166 579 167
rect 593 166 624 167
rect 511 165 530 166
rect 547 165 579 166
rect 594 165 625 166
rect 635 165 645 167
rect 512 164 528 165
rect 546 164 578 165
rect 595 164 625 165
rect 512 163 524 164
rect 544 163 578 164
rect 596 163 625 164
rect 636 163 645 165
rect 512 162 521 163
rect 542 162 578 163
rect 597 162 625 163
rect 513 161 518 162
rect 540 161 577 162
rect 598 161 625 162
rect 637 162 645 163
rect 538 160 577 161
rect 586 160 587 161
rect 599 160 626 161
rect 637 160 644 162
rect 536 159 577 160
rect 585 159 588 160
rect 599 159 625 160
rect 533 158 576 159
rect 585 158 589 159
rect 531 157 576 158
rect 584 157 589 158
rect 600 157 625 159
rect 638 159 644 160
rect 638 157 643 159
rect 529 156 575 157
rect 584 156 590 157
rect 527 155 575 156
rect 525 154 574 155
rect 583 154 591 156
rect 601 155 625 157
rect 639 155 642 157
rect 523 153 574 154
rect 522 152 573 153
rect 582 152 592 154
rect 601 153 624 155
rect 639 154 641 155
rect 639 153 640 154
rect 602 152 623 153
rect 521 151 572 152
rect 520 150 572 151
rect 519 149 571 150
rect 581 149 593 152
rect 602 151 622 152
rect 602 149 621 151
rect 518 148 570 149
rect 517 147 569 148
rect 580 147 594 149
rect 517 146 568 147
rect 579 146 594 147
rect 516 145 567 146
rect 516 144 566 145
rect 578 144 594 146
rect 603 148 620 149
rect 603 147 619 148
rect 603 146 618 147
rect 631 146 632 147
rect 603 145 616 146
rect 630 145 633 146
rect 603 144 615 145
rect 629 144 633 145
rect 515 143 565 144
rect 577 143 595 144
rect 515 142 564 143
rect 514 141 563 142
rect 576 141 595 143
rect 514 140 562 141
rect 575 140 595 141
rect 514 139 560 140
rect 574 139 595 140
rect 603 143 613 144
rect 628 143 633 144
rect 603 142 612 143
rect 627 142 633 143
rect 603 141 610 142
rect 626 141 633 142
rect 603 140 608 141
rect 625 140 633 141
rect 603 139 606 140
rect 624 139 633 140
rect 514 138 559 139
rect 573 138 595 139
rect 622 138 633 139
rect 513 137 557 138
rect 572 137 595 138
rect 621 137 633 138
rect 513 136 555 137
rect 570 136 595 137
rect 619 136 633 137
rect 513 135 554 136
rect 569 135 595 136
rect 618 135 633 136
rect 513 134 551 135
rect 568 134 594 135
rect 616 134 633 135
rect 513 133 549 134
rect 566 133 594 134
rect 614 133 633 134
rect 513 132 547 133
rect 564 132 594 133
rect 613 132 633 133
rect 513 131 545 132
rect 563 131 594 132
rect 611 131 633 132
rect 513 130 542 131
rect 561 130 594 131
rect 608 130 633 131
rect 513 129 540 130
rect 559 129 593 130
rect 606 129 633 130
rect 514 128 539 129
rect 557 128 593 129
rect 603 128 632 129
rect 514 127 537 128
rect 555 127 593 128
rect 600 127 632 128
rect 514 126 536 127
rect 553 126 593 127
rect 596 126 632 127
rect 514 125 535 126
rect 551 125 632 126
rect 514 124 534 125
rect 550 124 631 125
rect 515 123 533 124
rect 548 123 631 124
rect 515 121 532 123
rect 547 122 631 123
rect 545 121 630 122
rect 516 119 531 121
rect 544 120 630 121
rect 543 119 630 120
rect 517 117 530 119
rect 542 118 629 119
rect 541 117 573 118
rect 575 117 629 118
rect 518 115 530 117
rect 540 116 571 117
rect 575 116 628 117
rect 539 115 570 116
rect 574 115 628 116
rect 519 113 529 115
rect 538 114 568 115
rect 574 114 627 115
rect 538 113 567 114
rect 520 112 529 113
rect 521 110 529 112
rect 537 112 565 113
rect 573 112 626 114
rect 537 111 564 112
rect 572 111 625 112
rect 522 109 529 110
rect 536 110 562 111
rect 571 110 624 111
rect 536 109 561 110
rect 570 109 624 110
rect 523 108 528 109
rect 524 107 528 108
rect 525 106 528 107
rect 535 108 560 109
rect 570 108 593 109
rect 595 108 623 109
rect 535 107 559 108
rect 569 107 592 108
rect 594 107 622 108
rect 535 106 558 107
rect 568 106 591 107
rect 594 106 621 107
rect 526 105 528 106
rect 527 104 528 105
rect 534 105 557 106
rect 567 105 589 106
rect 534 104 556 105
rect 567 104 588 105
rect 593 104 620 106
rect 534 102 555 104
rect 566 103 587 104
rect 593 103 619 104
rect 566 102 586 103
rect 593 102 618 103
rect 533 101 554 102
rect 565 101 586 102
rect 592 101 617 102
rect 533 99 553 101
rect 565 100 585 101
rect 592 100 616 101
rect 533 97 552 99
rect 564 98 584 100
rect 592 99 614 100
rect 592 98 613 99
rect 534 96 552 97
rect 563 97 583 98
rect 592 97 612 98
rect 534 94 551 96
rect 563 94 582 97
rect 592 96 611 97
rect 591 95 610 96
rect 591 94 608 95
rect 535 92 551 94
rect 536 91 551 92
rect 537 90 551 91
rect 538 88 551 90
rect 539 87 551 88
rect 541 86 551 87
rect 542 85 551 86
rect 17 84 112 85
rect 173 84 206 85
rect 348 84 389 85
rect 409 84 442 85
rect 543 84 551 85
rect 349 83 390 84
rect 545 83 551 84
rect 350 82 391 83
rect 546 82 551 83
rect 562 91 581 94
rect 591 93 607 94
rect 591 92 606 93
rect 591 91 604 92
rect 562 86 580 91
rect 591 90 603 91
rect 591 89 602 90
rect 591 88 601 89
rect 592 87 600 88
rect 592 86 599 87
rect 351 81 392 82
rect 547 81 552 82
rect 562 81 579 86
rect 592 84 598 86
rect 592 83 597 84
rect 592 82 596 83
rect 352 80 393 81
rect 548 80 552 81
rect 353 79 394 80
rect 550 79 552 80
rect 551 78 552 79
rect 563 78 579 81
rect 593 81 596 82
rect 593 79 595 81
rect 593 78 594 79
rect 564 77 579 78
rect 564 76 580 77
rect 565 74 580 76
rect 566 73 580 74
rect 567 72 580 73
rect 568 71 580 72
rect 569 70 581 71
rect 570 69 581 70
rect 571 68 581 69
rect 572 67 582 68
rect 573 66 582 67
rect 574 65 582 66
rect 576 64 583 65
rect 10 63 22 64
rect 31 63 35 64
rect 134 63 138 64
rect 10 60 23 63
rect 10 59 22 60
rect 5 53 28 58
rect 31 52 36 63
rect 58 57 86 62
rect 80 54 86 57
rect 108 56 127 61
rect 114 55 120 56
rect 133 55 138 63
rect 182 63 186 64
rect 157 59 177 60
rect 157 55 178 59
rect 115 54 120 55
rect 127 54 138 55
rect 164 54 170 55
rect 37 52 39 53
rect 13 51 20 52
rect 10 50 23 51
rect 8 49 24 50
rect 7 48 25 49
rect 7 47 26 48
rect 6 46 13 47
rect 20 46 26 47
rect 6 43 12 46
rect 21 44 26 46
rect 31 47 40 52
rect 80 51 85 54
rect 114 53 120 54
rect 114 51 121 53
rect 79 48 85 51
rect 113 50 122 51
rect 126 50 138 54
rect 165 52 170 54
rect 113 49 123 50
rect 112 48 124 49
rect 21 43 27 44
rect 6 42 13 43
rect 19 42 26 43
rect 7 41 26 42
rect 8 40 25 41
rect 9 39 24 40
rect 11 38 22 39
rect 10 35 15 36
rect 31 35 36 47
rect 54 44 90 48
rect 111 47 125 48
rect 110 46 117 47
rect 118 46 126 47
rect 108 45 117 46
rect 119 45 128 46
rect 107 44 116 45
rect 120 44 128 45
rect 55 43 90 44
rect 105 43 115 44
rect 121 43 128 44
rect 69 37 74 43
rect 106 42 114 43
rect 122 42 127 43
rect 107 41 112 42
rect 124 41 126 42
rect 108 40 111 41
rect 10 30 16 35
rect 31 34 35 35
rect 58 32 86 37
rect 10 29 36 30
rect 10 25 37 29
rect 81 24 86 32
rect 112 30 117 38
rect 133 35 138 50
rect 164 49 170 52
rect 182 49 187 63
rect 210 59 237 63
rect 266 62 270 63
rect 266 59 271 62
rect 210 58 216 59
rect 234 58 235 59
rect 210 57 215 58
rect 210 56 236 57
rect 210 53 237 56
rect 265 54 271 59
rect 210 52 216 53
rect 265 52 272 54
rect 210 51 215 52
rect 264 51 272 52
rect 210 50 216 51
rect 263 50 273 51
rect 164 46 171 49
rect 163 45 171 46
rect 182 48 188 49
rect 190 48 191 49
rect 163 44 172 45
rect 162 43 172 44
rect 182 43 192 48
rect 210 46 237 50
rect 263 49 274 50
rect 262 48 275 49
rect 261 47 268 48
rect 269 47 276 48
rect 260 46 267 47
rect 269 46 277 47
rect 220 44 226 46
rect 259 45 266 46
rect 270 45 279 46
rect 257 44 266 45
rect 271 44 280 45
rect 206 43 240 44
rect 256 43 265 44
rect 272 43 280 44
rect 162 42 173 43
rect 161 41 173 42
rect 161 40 167 41
rect 160 39 167 40
rect 168 40 174 41
rect 168 39 175 40
rect 159 38 166 39
rect 169 38 176 39
rect 158 37 165 38
rect 157 36 165 37
rect 170 37 177 38
rect 170 36 178 37
rect 156 35 164 36
rect 171 35 179 36
rect 155 34 163 35
rect 172 34 178 35
rect 155 33 162 34
rect 173 33 178 34
rect 156 32 161 33
rect 175 32 177 33
rect 157 31 160 32
rect 112 25 139 30
rect 182 24 187 43
rect 205 39 241 43
rect 256 42 264 43
rect 274 42 279 43
rect 257 41 262 42
rect 275 41 278 42
rect 258 40 261 41
rect 259 39 260 40
rect 263 37 267 38
rect 215 36 231 37
rect 212 35 234 36
rect 211 34 235 35
rect 210 33 237 34
rect 209 32 218 33
rect 228 32 237 33
rect 209 29 215 32
rect 231 31 238 32
rect 232 30 238 31
rect 231 29 238 30
rect 263 30 268 37
rect 284 35 289 64
rect 318 62 319 63
rect 313 61 322 62
rect 312 60 324 61
rect 311 59 325 60
rect 334 59 339 64
rect 415 63 426 64
rect 414 62 427 63
rect 310 58 339 59
rect 309 57 317 58
rect 318 57 339 58
rect 360 57 388 62
rect 413 61 428 62
rect 412 60 429 61
rect 309 56 315 57
rect 321 56 339 57
rect 308 55 314 56
rect 308 50 313 55
rect 322 54 339 56
rect 322 53 328 54
rect 323 51 328 53
rect 334 51 339 54
rect 308 48 314 50
rect 322 49 339 51
rect 382 53 388 57
rect 411 59 418 60
rect 423 59 430 60
rect 411 58 417 59
rect 424 58 430 59
rect 411 55 416 58
rect 425 55 430 58
rect 411 54 418 55
rect 423 54 430 55
rect 411 53 429 54
rect 382 49 387 53
rect 412 52 429 53
rect 413 51 428 52
rect 415 50 426 51
rect 418 49 424 50
rect 321 48 339 49
rect 309 47 315 48
rect 320 47 339 48
rect 309 46 339 47
rect 310 45 326 46
rect 311 44 325 45
rect 312 43 323 44
rect 314 42 321 43
rect 313 30 318 38
rect 334 35 339 46
rect 381 48 387 49
rect 432 48 434 49
rect 381 45 386 48
rect 356 41 392 45
rect 408 44 434 48
rect 408 43 432 44
rect 357 40 392 41
rect 416 42 422 43
rect 263 29 289 30
rect 209 28 217 29
rect 229 28 237 29
rect 210 27 237 28
rect 211 26 236 27
rect 212 25 235 26
rect 263 25 290 29
rect 313 25 340 30
rect 214 24 232 25
rect 371 24 376 40
rect 416 36 421 42
rect 428 41 429 42
rect 430 41 434 42
rect 435 41 440 64
rect 578 63 583 64
rect 579 62 583 63
rect 581 61 584 62
rect 473 43 483 45
rect 486 43 495 45
rect 498 43 508 45
rect 512 43 520 45
rect 523 43 533 45
rect 538 43 547 45
rect 549 43 556 45
rect 565 43 573 45
rect 584 44 595 45
rect 581 43 587 44
rect 590 43 596 44
rect 609 43 619 45
rect 623 43 633 45
rect 638 43 654 45
rect 659 43 676 45
rect 475 42 481 43
rect 488 42 492 43
rect 500 42 506 43
rect 427 37 440 41
rect 414 30 419 35
rect 435 34 440 37
rect 476 34 480 42
rect 488 41 490 42
rect 501 41 506 42
rect 514 42 517 43
rect 525 42 531 43
rect 540 42 545 43
rect 552 42 557 43
rect 514 41 516 42
rect 487 40 489 41
rect 486 39 488 40
rect 502 39 507 41
rect 513 40 516 41
rect 513 39 515 40
rect 485 38 487 39
rect 484 37 486 38
rect 503 37 508 39
rect 512 37 514 39
rect 483 36 485 37
rect 504 36 509 37
rect 482 35 485 36
rect 505 35 509 36
rect 511 35 513 37
rect 481 34 486 35
rect 505 34 512 35
rect 476 33 487 34
rect 414 25 441 30
rect 476 25 480 33
rect 481 32 487 33
rect 506 33 512 34
rect 482 31 488 32
rect 483 30 489 31
rect 484 29 489 30
rect 484 28 490 29
rect 485 27 491 28
rect 486 26 492 27
rect 486 25 493 26
rect 475 24 481 25
rect 487 24 494 25
rect 506 24 511 33
rect 525 30 530 42
rect 526 29 530 30
rect 526 26 531 29
rect 541 28 544 42
rect 552 41 558 42
rect 552 40 559 41
rect 552 39 560 40
rect 568 39 571 43
rect 580 42 585 43
rect 592 42 596 43
rect 611 42 617 43
rect 625 42 631 43
rect 579 41 583 42
rect 593 41 596 42
rect 578 40 583 41
rect 594 40 596 41
rect 577 39 582 40
rect 540 26 543 28
rect 527 25 532 26
rect 539 25 543 26
rect 552 26 554 39
rect 555 38 561 39
rect 555 37 562 38
rect 556 36 563 37
rect 557 35 563 36
rect 558 34 564 35
rect 559 33 565 34
rect 560 32 566 33
rect 561 31 567 32
rect 561 30 568 31
rect 569 30 570 39
rect 576 36 581 39
rect 595 38 596 40
rect 612 41 617 42
rect 575 31 581 36
rect 612 35 616 41
rect 626 35 631 42
rect 612 33 631 35
rect 588 32 598 33
rect 589 31 597 32
rect 562 29 570 30
rect 563 28 570 29
rect 576 29 581 31
rect 591 30 596 31
rect 576 28 582 29
rect 564 27 570 28
rect 565 26 570 27
rect 577 27 582 28
rect 577 26 583 27
rect 527 24 534 25
rect 538 24 542 25
rect 552 24 555 26
rect 566 24 570 26
rect 578 25 583 26
rect 592 25 596 30
rect 612 25 616 33
rect 579 24 585 25
rect 219 23 228 24
rect 473 22 483 24
rect 488 22 496 24
rect 504 23 514 24
rect 528 23 541 24
rect 550 23 557 24
rect 567 23 570 24
rect 581 23 587 24
rect 591 23 596 25
rect 611 24 617 25
rect 626 24 631 33
rect 640 35 645 43
rect 651 42 654 43
rect 652 41 654 42
rect 653 39 654 41
rect 651 35 652 37
rect 640 33 652 35
rect 640 24 645 33
rect 650 32 652 33
rect 651 30 652 32
rect 662 35 667 43
rect 673 42 676 43
rect 674 39 676 42
rect 673 36 674 37
rect 672 35 674 36
rect 662 33 674 35
rect 654 26 656 28
rect 653 25 656 26
rect 652 24 655 25
rect 662 24 667 33
rect 672 31 674 33
rect 673 30 674 31
rect 676 27 678 28
rect 675 25 677 27
rect 674 24 677 25
rect 503 22 515 23
rect 530 22 540 23
rect 549 22 558 23
rect 568 22 570 23
rect 583 22 595 23
rect 609 22 619 24
rect 623 22 633 24
rect 637 22 655 24
rect 659 23 677 24
rect 659 22 676 23
rect 16 16 18 17
rect 123 16 124 17
rect 150 16 151 17
rect 361 16 362 17
rect 6 13 14 15
rect 6 9 9 13
rect 6 6 13 9
rect 6 3 9 6
rect 6 2 13 3
rect 6 0 14 2
rect 15 0 18 16
rect 23 11 25 12
rect 32 11 35 12
rect 38 11 41 14
rect 71 13 74 16
rect 48 11 49 12
rect 53 11 56 12
rect 65 11 67 12
rect 79 11 81 12
rect 86 11 88 12
rect 98 11 101 12
rect 110 11 112 12
rect 119 11 120 12
rect 122 11 125 16
rect 130 13 140 15
rect 133 12 137 13
rect 21 10 27 11
rect 31 10 43 11
rect 20 9 27 10
rect 30 9 43 10
rect 44 9 50 11
rect 52 10 58 11
rect 51 9 58 10
rect 61 9 69 11
rect 20 8 23 9
rect 20 7 22 8
rect 25 7 28 9
rect 20 4 28 7
rect 29 8 33 9
rect 20 3 22 4
rect 29 3 32 8
rect 20 2 23 3
rect 26 2 27 3
rect 30 2 33 3
rect 35 2 36 3
rect 20 1 28 2
rect 30 1 36 2
rect 38 2 41 9
rect 44 8 54 9
rect 38 1 43 2
rect 21 0 27 1
rect 31 0 36 1
rect 39 0 43 1
rect 44 0 47 8
rect 50 3 53 8
rect 56 7 59 9
rect 57 5 59 7
rect 56 3 59 5
rect 50 2 54 3
rect 55 2 59 3
rect 51 1 58 2
rect 52 0 57 1
rect 61 0 64 9
rect 66 8 69 9
rect 67 0 69 8
rect 71 0 74 11
rect 77 10 82 11
rect 84 10 90 11
rect 97 10 103 11
rect 106 10 113 11
rect 117 10 125 11
rect 76 9 82 10
rect 83 9 90 10
rect 96 9 104 10
rect 76 6 79 9
rect 83 7 86 9
rect 96 8 98 9
rect 101 7 104 9
rect 83 6 88 7
rect 97 6 104 7
rect 76 5 78 6
rect 84 5 89 6
rect 96 5 104 6
rect 76 3 79 5
rect 86 4 90 5
rect 96 4 99 5
rect 76 2 80 3
rect 81 2 82 3
rect 84 2 85 3
rect 87 2 90 4
rect 95 3 98 4
rect 101 3 104 5
rect 76 1 90 2
rect 96 2 99 3
rect 100 2 104 3
rect 96 1 104 2
rect 77 0 89 1
rect 97 0 104 1
rect 106 9 114 10
rect 106 7 109 9
rect 106 0 108 7
rect 111 0 114 9
rect 116 9 125 10
rect 116 6 119 9
rect 121 7 125 9
rect 116 5 118 6
rect 116 3 119 5
rect 122 4 125 7
rect 116 2 120 3
rect 121 2 125 4
rect 116 1 125 2
rect 117 0 125 1
rect 134 0 137 12
rect 142 11 144 12
rect 140 10 146 11
rect 139 9 146 10
rect 139 8 142 9
rect 139 7 141 8
rect 144 7 147 9
rect 138 4 147 7
rect 139 3 141 4
rect 139 2 142 3
rect 145 2 147 3
rect 139 1 147 2
rect 140 0 146 1
rect 149 0 151 16
rect 233 13 235 16
rect 256 13 258 14
rect 261 13 264 16
rect 299 14 307 15
rect 299 13 308 14
rect 156 11 158 12
rect 166 11 168 12
rect 174 11 176 12
rect 185 11 187 12
rect 190 11 192 12
rect 200 11 202 12
rect 206 11 208 12
rect 226 11 229 12
rect 240 11 243 12
rect 247 11 250 12
rect 255 11 258 13
rect 299 12 303 13
rect 304 12 308 13
rect 269 11 272 12
rect 281 11 283 12
rect 289 11 292 12
rect 154 10 160 11
rect 164 10 169 11
rect 172 10 178 11
rect 181 10 188 11
rect 189 10 194 11
rect 154 9 161 10
rect 153 7 156 9
rect 158 8 161 9
rect 163 9 169 10
rect 171 9 179 10
rect 163 8 166 9
rect 170 8 174 9
rect 159 7 161 8
rect 153 4 161 7
rect 162 4 165 8
rect 153 3 156 4
rect 162 3 166 4
rect 170 3 173 8
rect 176 7 179 9
rect 181 9 194 10
rect 177 4 180 7
rect 153 2 157 3
rect 159 2 161 3
rect 154 1 161 2
rect 163 2 167 3
rect 168 2 169 3
rect 170 2 174 3
rect 176 2 179 4
rect 163 1 169 2
rect 171 1 179 2
rect 155 0 161 1
rect 164 0 169 1
rect 172 0 178 1
rect 181 0 184 9
rect 186 8 190 9
rect 191 8 194 9
rect 186 0 189 8
rect 192 0 194 8
rect 196 9 209 11
rect 196 8 200 9
rect 196 0 199 8
rect 201 7 205 9
rect 202 0 204 7
rect 207 0 210 9
rect 212 3 214 11
rect 217 3 220 11
rect 212 2 215 3
rect 216 2 220 3
rect 212 1 220 2
rect 213 0 220 1
rect 222 9 230 11
rect 222 8 226 9
rect 227 8 231 9
rect 222 0 225 8
rect 228 0 231 8
rect 233 0 235 11
rect 239 10 244 11
rect 238 9 244 10
rect 245 9 252 11
rect 254 9 260 11
rect 237 8 241 9
rect 246 8 247 9
rect 237 3 240 8
rect 250 7 253 9
rect 246 6 253 7
rect 245 5 253 6
rect 245 4 248 5
rect 244 3 247 4
rect 250 3 253 5
rect 237 2 241 3
rect 243 2 244 3
rect 238 1 244 2
rect 239 0 244 1
rect 245 2 248 3
rect 249 2 253 3
rect 255 3 258 9
rect 255 2 259 3
rect 245 0 253 2
rect 256 0 260 2
rect 261 0 264 11
rect 267 10 273 11
rect 277 10 284 11
rect 267 9 274 10
rect 277 9 285 10
rect 287 9 293 11
rect 299 9 302 12
rect 305 9 308 12
rect 313 11 315 12
rect 321 11 324 12
rect 330 11 332 12
rect 339 11 342 12
rect 350 11 351 12
rect 355 11 358 12
rect 360 11 363 16
rect 365 11 366 12
rect 311 10 317 11
rect 320 10 325 11
rect 328 10 334 11
rect 310 9 317 10
rect 319 9 325 10
rect 327 9 335 10
rect 266 7 269 9
rect 271 8 275 9
rect 266 4 268 7
rect 266 3 269 4
rect 272 3 275 8
rect 276 7 280 9
rect 277 4 279 7
rect 266 2 270 3
rect 271 2 275 3
rect 276 2 279 4
rect 267 1 274 2
rect 268 0 273 1
rect 277 0 279 2
rect 282 0 285 9
rect 286 7 290 9
rect 287 6 292 7
rect 299 6 307 9
rect 310 8 313 9
rect 310 7 312 8
rect 315 7 318 9
rect 287 5 293 6
rect 289 4 293 5
rect 287 2 288 3
rect 290 2 293 4
rect 287 1 293 2
rect 287 0 292 1
rect 299 0 302 6
rect 304 5 307 6
rect 304 4 308 5
rect 309 4 318 7
rect 319 7 322 9
rect 327 8 330 9
rect 332 8 335 9
rect 337 9 344 11
rect 337 8 338 9
rect 341 8 344 9
rect 327 7 329 8
rect 333 7 335 8
rect 342 7 344 8
rect 319 6 324 7
rect 320 5 325 6
rect 322 4 326 5
rect 305 1 308 4
rect 310 3 312 4
rect 323 3 326 4
rect 310 2 313 3
rect 316 2 318 3
rect 310 1 318 2
rect 319 2 320 3
rect 322 2 326 3
rect 327 4 335 7
rect 338 6 344 7
rect 337 5 344 6
rect 327 2 330 4
rect 333 2 335 3
rect 306 0 309 1
rect 311 0 317 1
rect 319 0 325 2
rect 327 1 335 2
rect 336 2 339 5
rect 342 3 344 5
rect 341 2 344 3
rect 336 1 344 2
rect 346 9 352 11
rect 354 10 359 11
rect 353 9 359 10
rect 360 9 368 11
rect 346 8 351 9
rect 352 8 356 9
rect 360 8 364 9
rect 346 7 350 8
rect 328 0 335 1
rect 337 0 345 1
rect 346 0 349 7
rect 352 3 355 8
rect 352 2 356 3
rect 358 2 359 3
rect 353 1 359 2
rect 354 0 359 1
rect 360 0 363 8
rect 366 0 369 9
rect 375 0 378 15
rect 385 11 387 12
rect 393 11 396 12
rect 399 11 402 14
rect 405 13 408 16
rect 411 12 413 14
rect 410 11 413 12
rect 428 12 430 14
rect 596 12 599 13
rect 614 12 615 13
rect 623 12 624 13
rect 428 11 431 12
rect 436 11 439 12
rect 513 11 516 12
rect 380 10 388 11
rect 391 10 396 11
rect 380 9 389 10
rect 380 8 384 9
rect 380 0 383 8
rect 386 0 389 9
rect 390 9 396 10
rect 397 9 404 11
rect 390 8 393 9
rect 390 7 394 8
rect 390 6 396 7
rect 391 5 397 6
rect 393 4 397 5
rect 391 2 392 3
rect 394 2 397 4
rect 390 1 397 2
rect 399 2 402 9
rect 399 1 404 2
rect 390 0 396 1
rect 400 0 404 1
rect 405 0 408 11
rect 409 9 415 11
rect 411 3 413 9
rect 417 3 419 11
rect 422 3 425 11
rect 426 9 432 11
rect 435 10 440 11
rect 434 9 441 10
rect 411 2 414 3
rect 417 2 420 3
rect 421 2 425 3
rect 411 0 416 2
rect 417 1 425 2
rect 428 4 430 9
rect 434 8 436 9
rect 433 7 436 8
rect 439 8 441 9
rect 439 7 442 8
rect 433 4 442 7
rect 514 4 516 11
rect 521 10 523 12
rect 528 11 531 12
rect 536 11 538 12
rect 529 10 532 11
rect 428 2 431 4
rect 433 3 436 4
rect 514 3 517 4
rect 521 3 522 10
rect 529 9 533 10
rect 529 3 530 9
rect 531 8 534 9
rect 532 7 535 8
rect 532 6 536 7
rect 537 6 538 11
rect 533 5 538 6
rect 534 4 538 5
rect 535 3 538 4
rect 434 2 437 3
rect 440 2 441 3
rect 515 2 518 3
rect 519 2 521 3
rect 528 2 530 3
rect 536 2 538 3
rect 544 2 547 12
rect 553 10 556 12
rect 554 9 556 10
rect 560 10 562 12
rect 554 8 557 9
rect 560 8 561 10
rect 568 8 571 12
rect 573 11 575 12
rect 574 10 575 11
rect 581 11 584 12
rect 585 11 588 12
rect 595 11 596 12
rect 573 8 574 9
rect 555 7 557 8
rect 555 5 558 7
rect 559 5 560 8
rect 568 7 574 8
rect 556 3 559 5
rect 428 1 433 2
rect 434 1 441 2
rect 516 1 520 2
rect 537 1 538 2
rect 557 1 558 3
rect 568 2 571 7
rect 573 6 574 7
rect 581 7 583 11
rect 586 8 588 11
rect 594 9 596 11
rect 599 10 600 12
rect 594 8 597 9
rect 585 7 588 8
rect 595 7 599 8
rect 581 6 587 7
rect 596 6 600 7
rect 575 3 576 5
rect 574 2 576 3
rect 581 3 583 6
rect 585 5 587 6
rect 598 5 601 6
rect 585 4 588 5
rect 586 3 588 4
rect 594 3 595 4
rect 599 3 601 5
rect 581 2 584 3
rect 586 2 589 3
rect 594 2 596 3
rect 598 2 600 3
rect 606 2 609 12
rect 614 11 616 12
rect 614 9 615 11
rect 618 3 620 12
rect 622 11 624 12
rect 623 10 624 11
rect 629 10 632 12
rect 630 9 632 10
rect 635 11 637 12
rect 635 9 636 11
rect 631 8 633 9
rect 634 8 635 9
rect 631 7 635 8
rect 632 3 634 7
rect 617 2 620 3
rect 631 2 634 3
rect 588 1 590 2
rect 595 1 598 2
rect 418 0 425 1
rect 429 0 433 1
rect 435 0 441 1
<< end >>
